
module compare_N16384_CC4 ( clk, rst, x, y, g, e );
  input [4095:0] x;
  input [4095:0] y;
  input clk, rst;
  output g, e;
  wire   ebreg, n4, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626,
         n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
         n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
         n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,
         n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
         n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666,
         n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674,
         n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
         n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
         n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706,
         n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
         n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,
         n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
         n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,
         n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746,
         n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
         n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,
         n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770,
         n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778,
         n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786,
         n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794,
         n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802,
         n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810,
         n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818,
         n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826,
         n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834,
         n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842,
         n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850,
         n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858,
         n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866,
         n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874,
         n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882,
         n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890,
         n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898,
         n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906,
         n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914,
         n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922,
         n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930,
         n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938,
         n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946,
         n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954,
         n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962,
         n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970,
         n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978,
         n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986,
         n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994,
         n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002,
         n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010,
         n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
         n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,
         n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034,
         n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,
         n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050,
         n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058,
         n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066,
         n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
         n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082,
         n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,
         n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,
         n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106,
         n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114,
         n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122,
         n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130,
         n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
         n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146,
         n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154,
         n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,
         n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170,
         n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178,
         n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186,
         n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194,
         n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202,
         n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
         n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218,
         n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226,
         n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
         n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242,
         n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250,
         n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258,
         n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266,
         n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274,
         n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282,
         n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290,
         n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298,
         n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
         n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314,
         n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322,
         n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330,
         n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
         n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346,
         n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354,
         n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,
         n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370,
         n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
         n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386,
         n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394,
         n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402,
         n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
         n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,
         n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,
         n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,
         n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442,
         n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
         n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458,
         n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466,
         n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,
         n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
         n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490,
         n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
         n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
         n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
         n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
         n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538,
         n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546,
         n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
         n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562,
         n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,
         n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
         n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,
         n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
         n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602,
         n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610,
         n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618,
         n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626,
         n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634,
         n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642,
         n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650,
         n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658,
         n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
         n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674,
         n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682,
         n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690,
         n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
         n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706,
         n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714,
         n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722,
         n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730,
         n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,
         n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746,
         n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754,
         n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762,
         n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770,
         n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778,
         n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786,
         n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794,
         n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802,
         n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,
         n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818,
         n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826,
         n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834,
         n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842,
         n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850,
         n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858,
         n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866,
         n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874,
         n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,
         n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890,
         n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898,
         n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906,
         n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914,
         n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922,
         n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930,
         n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938,
         n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946,
         n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,
         n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962,
         n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970,
         n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978,
         n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986,
         n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994,
         n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002,
         n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010,
         n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018,
         n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
         n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034,
         n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042,
         n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050,
         n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058,
         n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
         n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074,
         n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082,
         n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090,
         n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
         n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106,
         n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114,
         n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122,
         n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130,
         n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,
         n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,
         n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
         n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
         n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
         n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178,
         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,
         n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194,
         n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,
         n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,
         n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218,
         n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
         n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234,
         n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
         n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250,
         n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258,
         n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266,
         n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
         n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282,
         n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290,
         n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
         n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306,
         n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314,
         n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322,
         n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330,
         n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338,
         n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346,
         n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
         n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362,
         n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,
         n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378,
         n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386,
         n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394,
         n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402,
         n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410,
         n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418,
         n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426,
         n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434,
         n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,
         n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450,
         n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458,
         n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466,
         n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474,
         n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482,
         n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490,
         n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498,
         n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506,
         n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514,
         n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522,
         n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530,
         n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538,
         n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546,
         n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554,
         n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562,
         n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570,
         n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578,
         n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586,
         n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594,
         n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602,
         n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610,
         n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618,
         n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626,
         n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634,
         n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642,
         n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650,
         n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658,
         n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666,
         n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674,
         n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682,
         n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690,
         n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698,
         n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706,
         n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714,
         n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722,
         n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730,
         n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738,
         n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746,
         n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754,
         n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762,
         n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770,
         n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778,
         n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786,
         n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794,
         n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802,
         n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810,
         n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818,
         n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826,
         n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834,
         n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842,
         n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850,
         n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858,
         n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866,
         n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874,
         n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882,
         n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890,
         n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898,
         n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906,
         n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914,
         n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922,
         n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930,
         n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938,
         n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946,
         n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954,
         n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962,
         n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970,
         n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978,
         n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986,
         n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994,
         n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002,
         n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010,
         n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018,
         n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026,
         n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034,
         n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042,
         n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050,
         n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058,
         n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066,
         n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074,
         n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082,
         n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090,
         n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098,
         n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106,
         n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114,
         n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122,
         n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130,
         n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138,
         n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146,
         n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154,
         n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162,
         n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170,
         n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178,
         n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186,
         n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194,
         n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202,
         n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210,
         n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218,
         n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226,
         n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234,
         n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242,
         n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250,
         n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258,
         n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266,
         n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274,
         n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282,
         n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290,
         n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298,
         n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306,
         n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314,
         n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322,
         n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330,
         n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338,
         n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346,
         n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354,
         n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362,
         n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370,
         n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378,
         n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386,
         n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394,
         n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402,
         n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410,
         n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418,
         n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426,
         n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434,
         n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442,
         n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450,
         n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458,
         n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466,
         n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474,
         n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482,
         n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490,
         n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498,
         n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506,
         n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514,
         n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522,
         n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530,
         n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538,
         n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546,
         n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554,
         n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562,
         n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570,
         n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578,
         n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586,
         n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594,
         n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602,
         n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610,
         n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618,
         n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626,
         n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634,
         n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642,
         n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650,
         n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658,
         n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666,
         n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674,
         n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682,
         n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690,
         n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698,
         n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706,
         n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714,
         n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722,
         n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730,
         n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738,
         n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746,
         n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754,
         n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762,
         n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770,
         n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778,
         n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786,
         n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794,
         n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802,
         n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810,
         n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818,
         n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826,
         n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834,
         n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842,
         n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850,
         n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858,
         n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866,
         n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874,
         n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882,
         n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890,
         n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898,
         n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906,
         n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914,
         n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922,
         n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930,
         n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938,
         n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946,
         n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954,
         n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962,
         n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970,
         n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978,
         n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986,
         n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994,
         n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002,
         n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010,
         n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018,
         n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026,
         n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034,
         n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042,
         n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050,
         n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058,
         n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066,
         n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074,
         n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082,
         n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090,
         n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098,
         n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106,
         n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114,
         n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122,
         n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130,
         n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138,
         n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146,
         n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154,
         n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162,
         n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170,
         n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178,
         n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186,
         n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194,
         n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202,
         n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210,
         n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218,
         n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226,
         n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234,
         n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242,
         n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250,
         n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258,
         n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266,
         n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274,
         n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282,
         n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290,
         n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298,
         n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306,
         n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314,
         n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322,
         n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330,
         n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338,
         n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346,
         n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354,
         n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362,
         n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370,
         n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378,
         n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386,
         n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394,
         n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402,
         n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410,
         n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418,
         n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426,
         n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434,
         n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442,
         n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450,
         n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458,
         n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466,
         n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474,
         n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482,
         n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490,
         n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498,
         n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506,
         n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514,
         n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522,
         n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530,
         n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538,
         n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546,
         n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554,
         n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562,
         n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570,
         n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578,
         n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586,
         n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594,
         n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602,
         n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610,
         n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618,
         n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626,
         n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634,
         n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642,
         n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650,
         n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658,
         n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666,
         n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674,
         n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682,
         n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690,
         n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698,
         n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706,
         n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714,
         n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
         n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730,
         n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738,
         n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746,
         n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754,
         n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762,
         n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770,
         n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778,
         n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786,
         n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794,
         n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802,
         n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810,
         n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818,
         n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826,
         n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834,
         n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842,
         n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850,
         n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858,
         n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866,
         n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874,
         n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882,
         n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890,
         n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898,
         n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906,
         n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914,
         n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922,
         n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930,
         n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
         n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946,
         n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954,
         n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962,
         n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970,
         n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978,
         n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986,
         n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994,
         n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002,
         n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010,
         n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018,
         n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026,
         n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034,
         n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042,
         n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050,
         n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058,
         n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066,
         n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074,
         n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082,
         n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090,
         n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098,
         n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106,
         n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114,
         n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122,
         n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130,
         n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138,
         n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146,
         n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154,
         n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162,
         n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170,
         n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178,
         n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186,
         n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194,
         n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202,
         n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210,
         n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218,
         n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226,
         n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234,
         n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242,
         n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250,
         n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258,
         n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266,
         n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274,
         n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282,
         n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290,
         n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298,
         n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306,
         n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314,
         n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322,
         n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330,
         n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338,
         n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346,
         n21347, n21348, n21349, n21350, n21351, n21352, n21353, n21354,
         n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362,
         n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370,
         n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378,
         n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386,
         n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394,
         n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402,
         n21403, n21404, n21405, n21406, n21407, n21408, n21409, n21410,
         n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418,
         n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426,
         n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434,
         n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442,
         n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450,
         n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458,
         n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466,
         n21467, n21468, n21469, n21470, n21471, n21472, n21473, n21474,
         n21475, n21476, n21477, n21478, n21479, n21480, n21481, n21482,
         n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490,
         n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498,
         n21499, n21500, n21501, n21502, n21503, n21504, n21505, n21506,
         n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514,
         n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522,
         n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530,
         n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538,
         n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546,
         n21547, n21548, n21549, n21550, n21551, n21552, n21553, n21554,
         n21555, n21556, n21557, n21558, n21559, n21560, n21561, n21562,
         n21563, n21564, n21565, n21566, n21567, n21568, n21569, n21570,
         n21571, n21572, n21573, n21574, n21575, n21576, n21577, n21578,
         n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586,
         n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594,
         n21595, n21596, n21597, n21598, n21599, n21600, n21601, n21602,
         n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610,
         n21611, n21612, n21613, n21614, n21615, n21616, n21617, n21618,
         n21619, n21620, n21621, n21622, n21623, n21624, n21625, n21626,
         n21627, n21628, n21629, n21630, n21631, n21632, n21633, n21634,
         n21635, n21636, n21637, n21638, n21639, n21640, n21641, n21642,
         n21643, n21644, n21645, n21646, n21647, n21648, n21649, n21650,
         n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658,
         n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666,
         n21667, n21668, n21669, n21670, n21671, n21672, n21673, n21674,
         n21675, n21676, n21677, n21678, n21679, n21680, n21681, n21682,
         n21683, n21684, n21685, n21686, n21687, n21688, n21689, n21690,
         n21691, n21692, n21693, n21694, n21695, n21696, n21697, n21698,
         n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706,
         n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21714,
         n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722,
         n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730,
         n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738,
         n21739, n21740, n21741, n21742, n21743, n21744, n21745, n21746,
         n21747, n21748, n21749, n21750, n21751, n21752, n21753, n21754,
         n21755, n21756, n21757, n21758, n21759, n21760, n21761, n21762,
         n21763, n21764, n21765, n21766, n21767, n21768, n21769, n21770,
         n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778,
         n21779, n21780, n21781, n21782, n21783, n21784, n21785, n21786,
         n21787, n21788, n21789, n21790, n21791, n21792, n21793, n21794,
         n21795, n21796, n21797, n21798, n21799, n21800, n21801, n21802,
         n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810,
         n21811, n21812, n21813, n21814, n21815, n21816, n21817, n21818,
         n21819, n21820, n21821, n21822, n21823, n21824, n21825, n21826,
         n21827, n21828, n21829, n21830, n21831, n21832, n21833, n21834,
         n21835, n21836, n21837, n21838, n21839, n21840, n21841, n21842,
         n21843, n21844, n21845, n21846, n21847, n21848, n21849, n21850,
         n21851, n21852, n21853, n21854, n21855, n21856, n21857, n21858,
         n21859, n21860, n21861, n21862, n21863, n21864, n21865, n21866,
         n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21874,
         n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882,
         n21883, n21884, n21885, n21886, n21887, n21888, n21889, n21890,
         n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21898,
         n21899, n21900, n21901, n21902, n21903, n21904, n21905, n21906,
         n21907, n21908, n21909, n21910, n21911, n21912, n21913, n21914,
         n21915, n21916, n21917, n21918, n21919, n21920, n21921, n21922,
         n21923, n21924, n21925, n21926, n21927, n21928, n21929, n21930,
         n21931, n21932, n21933, n21934, n21935, n21936, n21937, n21938,
         n21939, n21940, n21941, n21942, n21943, n21944, n21945, n21946,
         n21947, n21948, n21949, n21950, n21951, n21952, n21953, n21954,
         n21955, n21956, n21957, n21958, n21959, n21960, n21961, n21962,
         n21963, n21964, n21965, n21966, n21967, n21968, n21969, n21970,
         n21971, n21972, n21973, n21974, n21975, n21976, n21977, n21978,
         n21979, n21980, n21981, n21982, n21983, n21984, n21985, n21986,
         n21987, n21988, n21989, n21990, n21991, n21992, n21993, n21994,
         n21995, n21996, n21997, n21998, n21999, n22000, n22001, n22002,
         n22003, n22004, n22005, n22006, n22007, n22008, n22009, n22010,
         n22011, n22012, n22013, n22014, n22015, n22016, n22017, n22018,
         n22019, n22020, n22021, n22022, n22023, n22024, n22025, n22026,
         n22027, n22028, n22029, n22030, n22031, n22032, n22033, n22034,
         n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042,
         n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050,
         n22051, n22052, n22053, n22054, n22055, n22056, n22057, n22058,
         n22059, n22060, n22061, n22062, n22063, n22064, n22065, n22066,
         n22067, n22068, n22069, n22070, n22071, n22072, n22073, n22074,
         n22075, n22076, n22077, n22078, n22079, n22080, n22081, n22082,
         n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090,
         n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098,
         n22099, n22100, n22101, n22102, n22103, n22104, n22105, n22106,
         n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114,
         n22115, n22116, n22117, n22118, n22119, n22120, n22121, n22122,
         n22123, n22124, n22125, n22126, n22127, n22128, n22129, n22130,
         n22131, n22132, n22133, n22134, n22135, n22136, n22137, n22138,
         n22139, n22140, n22141, n22142, n22143, n22144, n22145, n22146,
         n22147, n22148, n22149, n22150, n22151, n22152, n22153, n22154,
         n22155, n22156, n22157, n22158, n22159, n22160, n22161, n22162,
         n22163, n22164, n22165, n22166, n22167, n22168, n22169, n22170,
         n22171, n22172, n22173, n22174, n22175, n22176, n22177, n22178,
         n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22186,
         n22187, n22188, n22189, n22190, n22191, n22192, n22193, n22194,
         n22195, n22196, n22197, n22198, n22199, n22200, n22201, n22202,
         n22203, n22204, n22205, n22206, n22207, n22208, n22209, n22210,
         n22211, n22212, n22213, n22214, n22215, n22216, n22217, n22218,
         n22219, n22220, n22221, n22222, n22223, n22224, n22225, n22226,
         n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22234,
         n22235, n22236, n22237, n22238, n22239, n22240, n22241, n22242,
         n22243, n22244, n22245, n22246, n22247, n22248, n22249, n22250,
         n22251, n22252, n22253, n22254, n22255, n22256, n22257, n22258,
         n22259, n22260, n22261, n22262, n22263, n22264, n22265, n22266,
         n22267, n22268, n22269, n22270, n22271, n22272, n22273, n22274,
         n22275, n22276, n22277, n22278, n22279, n22280, n22281, n22282,
         n22283, n22284, n22285, n22286, n22287, n22288, n22289, n22290,
         n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298,
         n22299, n22300, n22301, n22302, n22303, n22304, n22305, n22306,
         n22307, n22308, n22309, n22310, n22311, n22312, n22313, n22314,
         n22315, n22316, n22317, n22318, n22319, n22320, n22321, n22322,
         n22323, n22324, n22325, n22326, n22327, n22328, n22329, n22330,
         n22331, n22332, n22333, n22334, n22335, n22336, n22337, n22338,
         n22339, n22340, n22341, n22342, n22343, n22344, n22345, n22346,
         n22347, n22348, n22349, n22350, n22351, n22352, n22353, n22354,
         n22355, n22356, n22357, n22358, n22359, n22360, n22361, n22362,
         n22363, n22364, n22365, n22366, n22367, n22368, n22369, n22370,
         n22371, n22372, n22373, n22374, n22375, n22376, n22377, n22378,
         n22379, n22380, n22381, n22382, n22383, n22384, n22385, n22386,
         n22387, n22388, n22389, n22390, n22391, n22392, n22393, n22394,
         n22395, n22396, n22397, n22398, n22399, n22400, n22401, n22402,
         n22403, n22404, n22405, n22406, n22407, n22408, n22409, n22410,
         n22411, n22412, n22413, n22414, n22415, n22416, n22417, n22418,
         n22419, n22420, n22421, n22422, n22423, n22424, n22425, n22426,
         n22427, n22428, n22429, n22430, n22431, n22432, n22433, n22434,
         n22435, n22436, n22437, n22438, n22439, n22440, n22441, n22442,
         n22443, n22444, n22445, n22446, n22447, n22448, n22449, n22450,
         n22451, n22452, n22453, n22454, n22455, n22456, n22457, n22458,
         n22459, n22460, n22461, n22462, n22463, n22464, n22465, n22466,
         n22467, n22468, n22469, n22470, n22471, n22472, n22473, n22474,
         n22475, n22476, n22477, n22478, n22479, n22480, n22481, n22482,
         n22483, n22484, n22485, n22486, n22487, n22488, n22489, n22490,
         n22491, n22492, n22493, n22494, n22495, n22496, n22497, n22498,
         n22499, n22500, n22501, n22502, n22503, n22504, n22505, n22506,
         n22507, n22508, n22509, n22510, n22511, n22512, n22513, n22514,
         n22515, n22516, n22517, n22518, n22519, n22520, n22521, n22522,
         n22523, n22524, n22525, n22526, n22527, n22528, n22529, n22530,
         n22531, n22532, n22533, n22534, n22535, n22536, n22537, n22538,
         n22539, n22540, n22541, n22542, n22543, n22544, n22545, n22546,
         n22547, n22548, n22549, n22550, n22551, n22552, n22553, n22554,
         n22555, n22556, n22557, n22558, n22559, n22560, n22561, n22562,
         n22563, n22564, n22565, n22566, n22567, n22568, n22569, n22570,
         n22571, n22572, n22573, n22574, n22575, n22576, n22577, n22578,
         n22579, n22580, n22581, n22582, n22583, n22584, n22585, n22586,
         n22587, n22588, n22589, n22590, n22591, n22592, n22593, n22594,
         n22595, n22596, n22597, n22598, n22599, n22600, n22601, n22602,
         n22603, n22604, n22605, n22606, n22607, n22608, n22609, n22610,
         n22611, n22612, n22613, n22614, n22615, n22616, n22617, n22618,
         n22619, n22620, n22621, n22622, n22623, n22624, n22625, n22626,
         n22627, n22628, n22629, n22630, n22631, n22632, n22633, n22634,
         n22635, n22636, n22637, n22638, n22639, n22640, n22641, n22642,
         n22643, n22644, n22645, n22646, n22647, n22648, n22649, n22650,
         n22651, n22652, n22653, n22654, n22655, n22656, n22657, n22658,
         n22659, n22660, n22661, n22662, n22663, n22664, n22665, n22666,
         n22667, n22668, n22669, n22670, n22671, n22672, n22673, n22674,
         n22675, n22676, n22677, n22678, n22679, n22680, n22681, n22682,
         n22683, n22684, n22685, n22686, n22687, n22688, n22689, n22690,
         n22691, n22692, n22693, n22694, n22695, n22696, n22697, n22698,
         n22699, n22700, n22701, n22702, n22703, n22704, n22705, n22706,
         n22707, n22708, n22709, n22710, n22711, n22712, n22713, n22714,
         n22715, n22716, n22717, n22718, n22719, n22720, n22721, n22722,
         n22723, n22724, n22725, n22726, n22727, n22728, n22729, n22730,
         n22731, n22732, n22733, n22734, n22735, n22736, n22737, n22738,
         n22739, n22740, n22741, n22742, n22743, n22744, n22745, n22746,
         n22747, n22748, n22749, n22750, n22751, n22752, n22753, n22754,
         n22755, n22756, n22757, n22758, n22759, n22760, n22761, n22762,
         n22763, n22764, n22765, n22766, n22767, n22768, n22769, n22770,
         n22771, n22772, n22773, n22774, n22775, n22776, n22777, n22778,
         n22779, n22780, n22781, n22782, n22783, n22784, n22785, n22786,
         n22787, n22788, n22789, n22790, n22791, n22792, n22793, n22794,
         n22795, n22796, n22797, n22798, n22799, n22800, n22801, n22802,
         n22803, n22804, n22805, n22806, n22807, n22808, n22809, n22810,
         n22811, n22812, n22813, n22814, n22815, n22816, n22817, n22818,
         n22819, n22820, n22821, n22822, n22823, n22824, n22825, n22826,
         n22827, n22828, n22829, n22830, n22831, n22832, n22833, n22834,
         n22835, n22836, n22837, n22838, n22839, n22840, n22841, n22842,
         n22843, n22844, n22845, n22846, n22847, n22848, n22849, n22850,
         n22851, n22852, n22853, n22854, n22855, n22856, n22857, n22858,
         n22859, n22860, n22861, n22862, n22863, n22864, n22865, n22866,
         n22867, n22868, n22869, n22870, n22871, n22872, n22873, n22874,
         n22875, n22876, n22877, n22878, n22879, n22880, n22881, n22882,
         n22883, n22884, n22885, n22886, n22887, n22888, n22889, n22890,
         n22891, n22892, n22893, n22894, n22895, n22896, n22897, n22898,
         n22899, n22900, n22901, n22902, n22903, n22904, n22905, n22906,
         n22907, n22908, n22909, n22910, n22911, n22912, n22913, n22914,
         n22915, n22916, n22917, n22918, n22919, n22920, n22921, n22922,
         n22923, n22924, n22925, n22926, n22927, n22928, n22929, n22930,
         n22931, n22932, n22933, n22934, n22935, n22936, n22937, n22938,
         n22939, n22940, n22941, n22942, n22943, n22944, n22945, n22946,
         n22947, n22948, n22949, n22950, n22951, n22952, n22953, n22954,
         n22955, n22956, n22957, n22958, n22959, n22960, n22961, n22962,
         n22963, n22964, n22965, n22966, n22967, n22968, n22969, n22970,
         n22971, n22972, n22973, n22974, n22975, n22976, n22977, n22978,
         n22979, n22980, n22981, n22982, n22983, n22984, n22985, n22986,
         n22987, n22988, n22989, n22990, n22991, n22992, n22993, n22994,
         n22995, n22996, n22997, n22998, n22999, n23000, n23001, n23002,
         n23003, n23004, n23005, n23006, n23007, n23008, n23009, n23010,
         n23011, n23012, n23013, n23014, n23015, n23016, n23017, n23018,
         n23019, n23020, n23021, n23022, n23023, n23024, n23025, n23026,
         n23027, n23028, n23029, n23030, n23031, n23032, n23033, n23034,
         n23035, n23036, n23037, n23038, n23039, n23040, n23041, n23042,
         n23043, n23044, n23045, n23046, n23047, n23048, n23049, n23050,
         n23051, n23052, n23053, n23054, n23055, n23056, n23057, n23058,
         n23059, n23060, n23061, n23062, n23063, n23064, n23065, n23066,
         n23067, n23068, n23069, n23070, n23071, n23072, n23073, n23074,
         n23075, n23076, n23077, n23078, n23079, n23080, n23081, n23082,
         n23083, n23084, n23085, n23086, n23087, n23088, n23089, n23090,
         n23091, n23092, n23093, n23094, n23095, n23096, n23097, n23098,
         n23099, n23100, n23101, n23102, n23103, n23104, n23105, n23106,
         n23107, n23108, n23109, n23110, n23111, n23112, n23113, n23114,
         n23115, n23116, n23117, n23118, n23119, n23120, n23121, n23122,
         n23123, n23124, n23125, n23126, n23127, n23128, n23129, n23130,
         n23131, n23132, n23133, n23134, n23135, n23136, n23137, n23138,
         n23139, n23140, n23141, n23142, n23143, n23144, n23145, n23146,
         n23147, n23148, n23149, n23150, n23151, n23152, n23153, n23154,
         n23155, n23156, n23157, n23158, n23159, n23160, n23161, n23162,
         n23163, n23164, n23165, n23166, n23167, n23168, n23169, n23170,
         n23171, n23172, n23173, n23174, n23175, n23176, n23177, n23178,
         n23179, n23180, n23181, n23182, n23183, n23184, n23185, n23186,
         n23187, n23188, n23189, n23190, n23191, n23192, n23193, n23194,
         n23195, n23196, n23197, n23198, n23199, n23200, n23201, n23202,
         n23203, n23204, n23205, n23206, n23207, n23208, n23209, n23210,
         n23211, n23212, n23213, n23214, n23215, n23216, n23217, n23218,
         n23219, n23220, n23221, n23222, n23223, n23224, n23225, n23226,
         n23227, n23228, n23229, n23230, n23231, n23232, n23233, n23234,
         n23235, n23236, n23237, n23238, n23239, n23240, n23241, n23242,
         n23243, n23244, n23245, n23246, n23247, n23248, n23249, n23250,
         n23251, n23252, n23253, n23254, n23255, n23256, n23257, n23258,
         n23259, n23260, n23261, n23262, n23263, n23264, n23265, n23266,
         n23267, n23268, n23269, n23270, n23271, n23272, n23273, n23274,
         n23275, n23276, n23277, n23278, n23279, n23280, n23281, n23282,
         n23283, n23284, n23285, n23286, n23287, n23288, n23289, n23290,
         n23291, n23292, n23293, n23294, n23295, n23296, n23297, n23298,
         n23299, n23300, n23301, n23302, n23303, n23304, n23305, n23306,
         n23307, n23308, n23309, n23310, n23311, n23312, n23313, n23314,
         n23315, n23316, n23317, n23318, n23319, n23320, n23321, n23322,
         n23323, n23324, n23325, n23326, n23327, n23328, n23329, n23330,
         n23331, n23332, n23333, n23334, n23335, n23336, n23337, n23338,
         n23339, n23340, n23341, n23342, n23343, n23344, n23345, n23346,
         n23347, n23348, n23349, n23350, n23351, n23352, n23353, n23354,
         n23355, n23356, n23357, n23358, n23359, n23360, n23361, n23362,
         n23363, n23364, n23365, n23366, n23367, n23368, n23369, n23370,
         n23371, n23372, n23373, n23374, n23375, n23376, n23377, n23378,
         n23379, n23380, n23381, n23382, n23383, n23384, n23385, n23386,
         n23387, n23388, n23389, n23390, n23391, n23392, n23393, n23394,
         n23395, n23396, n23397, n23398, n23399, n23400, n23401, n23402,
         n23403, n23404, n23405, n23406, n23407, n23408, n23409, n23410,
         n23411, n23412, n23413, n23414, n23415, n23416, n23417, n23418,
         n23419, n23420, n23421, n23422, n23423, n23424, n23425, n23426,
         n23427, n23428, n23429, n23430, n23431, n23432, n23433, n23434,
         n23435, n23436, n23437, n23438, n23439, n23440, n23441, n23442,
         n23443, n23444, n23445, n23446, n23447, n23448, n23449, n23450,
         n23451, n23452, n23453, n23454, n23455, n23456, n23457, n23458,
         n23459, n23460, n23461, n23462, n23463, n23464, n23465, n23466,
         n23467, n23468, n23469, n23470, n23471, n23472, n23473, n23474,
         n23475, n23476, n23477, n23478, n23479, n23480, n23481, n23482,
         n23483, n23484, n23485, n23486, n23487, n23488, n23489, n23490,
         n23491, n23492, n23493, n23494, n23495, n23496, n23497, n23498,
         n23499, n23500, n23501, n23502, n23503, n23504, n23505, n23506,
         n23507, n23508, n23509, n23510, n23511, n23512, n23513, n23514,
         n23515, n23516, n23517, n23518, n23519, n23520, n23521, n23522,
         n23523, n23524, n23525, n23526, n23527, n23528, n23529, n23530,
         n23531, n23532, n23533, n23534, n23535, n23536, n23537, n23538,
         n23539, n23540, n23541, n23542, n23543, n23544, n23545, n23546,
         n23547, n23548, n23549, n23550, n23551, n23552, n23553, n23554,
         n23555, n23556, n23557, n23558, n23559, n23560, n23561, n23562,
         n23563, n23564, n23565, n23566, n23567, n23568, n23569, n23570,
         n23571, n23572, n23573, n23574, n23575, n23576, n23577, n23578,
         n23579, n23580, n23581, n23582, n23583, n23584, n23585, n23586,
         n23587, n23588, n23589, n23590, n23591, n23592, n23593, n23594,
         n23595, n23596, n23597, n23598, n23599, n23600, n23601, n23602,
         n23603, n23604, n23605, n23606, n23607, n23608, n23609, n23610,
         n23611, n23612, n23613, n23614, n23615, n23616, n23617, n23618,
         n23619, n23620, n23621, n23622, n23623, n23624, n23625, n23626,
         n23627, n23628, n23629, n23630, n23631, n23632, n23633, n23634,
         n23635, n23636, n23637, n23638, n23639, n23640, n23641, n23642,
         n23643, n23644, n23645, n23646, n23647, n23648, n23649, n23650,
         n23651, n23652, n23653, n23654, n23655, n23656, n23657, n23658,
         n23659, n23660, n23661, n23662, n23663, n23664, n23665, n23666,
         n23667, n23668, n23669, n23670, n23671, n23672, n23673, n23674,
         n23675, n23676, n23677, n23678, n23679, n23680, n23681, n23682,
         n23683, n23684, n23685, n23686, n23687, n23688, n23689, n23690,
         n23691, n23692, n23693, n23694, n23695, n23696, n23697, n23698,
         n23699, n23700, n23701, n23702, n23703, n23704, n23705, n23706,
         n23707, n23708, n23709, n23710, n23711, n23712, n23713, n23714,
         n23715, n23716, n23717, n23718, n23719, n23720, n23721, n23722,
         n23723, n23724, n23725, n23726, n23727, n23728, n23729, n23730,
         n23731, n23732, n23733, n23734, n23735, n23736, n23737, n23738,
         n23739, n23740, n23741, n23742, n23743, n23744, n23745, n23746,
         n23747, n23748, n23749, n23750, n23751, n23752, n23753, n23754,
         n23755, n23756, n23757, n23758, n23759, n23760, n23761, n23762,
         n23763, n23764, n23765, n23766, n23767, n23768, n23769, n23770,
         n23771, n23772, n23773, n23774, n23775, n23776, n23777, n23778,
         n23779, n23780, n23781, n23782, n23783, n23784, n23785, n23786,
         n23787, n23788, n23789, n23790, n23791, n23792, n23793, n23794,
         n23795, n23796, n23797, n23798, n23799, n23800, n23801, n23802,
         n23803, n23804, n23805, n23806, n23807, n23808, n23809, n23810,
         n23811, n23812, n23813, n23814, n23815, n23816, n23817, n23818,
         n23819, n23820, n23821, n23822, n23823, n23824, n23825, n23826,
         n23827, n23828, n23829, n23830, n23831, n23832, n23833, n23834,
         n23835, n23836, n23837, n23838, n23839, n23840, n23841, n23842,
         n23843, n23844, n23845, n23846, n23847, n23848, n23849, n23850,
         n23851, n23852, n23853, n23854, n23855, n23856, n23857, n23858,
         n23859, n23860, n23861, n23862, n23863, n23864, n23865, n23866,
         n23867, n23868, n23869, n23870, n23871, n23872, n23873, n23874,
         n23875, n23876, n23877, n23878, n23879, n23880, n23881, n23882,
         n23883, n23884, n23885, n23886, n23887, n23888, n23889, n23890,
         n23891, n23892, n23893, n23894, n23895, n23896, n23897, n23898,
         n23899, n23900, n23901, n23902, n23903, n23904, n23905, n23906,
         n23907, n23908, n23909, n23910, n23911, n23912, n23913, n23914,
         n23915, n23916, n23917, n23918, n23919, n23920, n23921, n23922,
         n23923, n23924, n23925, n23926, n23927, n23928, n23929, n23930,
         n23931, n23932, n23933, n23934, n23935, n23936, n23937, n23938,
         n23939, n23940, n23941, n23942, n23943, n23944, n23945, n23946,
         n23947, n23948, n23949, n23950, n23951, n23952, n23953, n23954,
         n23955, n23956, n23957, n23958, n23959, n23960, n23961, n23962,
         n23963, n23964, n23965, n23966, n23967, n23968, n23969, n23970,
         n23971, n23972, n23973, n23974, n23975, n23976, n23977, n23978,
         n23979, n23980, n23981, n23982, n23983, n23984, n23985, n23986,
         n23987, n23988, n23989, n23990, n23991, n23992, n23993, n23994,
         n23995, n23996, n23997, n23998, n23999, n24000, n24001, n24002,
         n24003, n24004, n24005, n24006, n24007, n24008, n24009, n24010,
         n24011, n24012, n24013, n24014, n24015, n24016, n24017, n24018,
         n24019, n24020, n24021, n24022, n24023, n24024, n24025, n24026,
         n24027, n24028, n24029, n24030, n24031, n24032, n24033, n24034,
         n24035, n24036, n24037, n24038, n24039, n24040, n24041, n24042,
         n24043, n24044, n24045, n24046, n24047, n24048, n24049, n24050,
         n24051, n24052, n24053, n24054, n24055, n24056, n24057, n24058,
         n24059, n24060, n24061, n24062, n24063, n24064, n24065, n24066,
         n24067, n24068, n24069, n24070, n24071, n24072, n24073, n24074,
         n24075, n24076, n24077, n24078, n24079, n24080, n24081, n24082,
         n24083, n24084, n24085, n24086, n24087, n24088, n24089, n24090,
         n24091, n24092, n24093, n24094, n24095, n24096, n24097, n24098,
         n24099, n24100, n24101, n24102, n24103, n24104, n24105, n24106,
         n24107, n24108, n24109, n24110, n24111, n24112, n24113, n24114,
         n24115, n24116, n24117, n24118, n24119, n24120, n24121, n24122,
         n24123, n24124, n24125, n24126, n24127, n24128, n24129, n24130,
         n24131, n24132, n24133, n24134, n24135, n24136, n24137, n24138,
         n24139, n24140, n24141, n24142, n24143, n24144, n24145, n24146,
         n24147, n24148, n24149, n24150, n24151, n24152, n24153, n24154,
         n24155, n24156, n24157, n24158, n24159, n24160, n24161, n24162,
         n24163, n24164, n24165, n24166, n24167, n24168, n24169, n24170,
         n24171, n24172, n24173, n24174, n24175, n24176, n24177, n24178,
         n24179, n24180, n24181, n24182, n24183, n24184, n24185, n24186,
         n24187, n24188, n24189, n24190, n24191, n24192, n24193, n24194,
         n24195, n24196, n24197, n24198, n24199, n24200, n24201, n24202,
         n24203, n24204, n24205, n24206, n24207, n24208, n24209, n24210,
         n24211, n24212, n24213, n24214, n24215, n24216, n24217, n24218,
         n24219, n24220, n24221, n24222, n24223, n24224, n24225, n24226,
         n24227, n24228, n24229, n24230, n24231, n24232, n24233, n24234,
         n24235, n24236, n24237, n24238, n24239, n24240, n24241, n24242,
         n24243, n24244, n24245, n24246, n24247, n24248, n24249, n24250,
         n24251, n24252, n24253, n24254, n24255, n24256, n24257, n24258,
         n24259, n24260, n24261, n24262, n24263, n24264, n24265, n24266,
         n24267, n24268, n24269, n24270, n24271, n24272, n24273, n24274,
         n24275, n24276, n24277, n24278, n24279, n24280, n24281, n24282,
         n24283, n24284, n24285, n24286, n24287, n24288, n24289, n24290,
         n24291, n24292, n24293, n24294, n24295, n24296, n24297, n24298,
         n24299, n24300, n24301, n24302, n24303, n24304, n24305, n24306,
         n24307, n24308, n24309, n24310, n24311, n24312, n24313, n24314,
         n24315, n24316, n24317, n24318, n24319, n24320, n24321, n24322,
         n24323, n24324, n24325, n24326, n24327, n24328, n24329, n24330,
         n24331, n24332, n24333, n24334, n24335, n24336, n24337, n24338,
         n24339, n24340, n24341, n24342, n24343, n24344, n24345, n24346,
         n24347, n24348, n24349, n24350, n24351, n24352, n24353, n24354,
         n24355, n24356, n24357, n24358, n24359, n24360, n24361, n24362,
         n24363, n24364, n24365, n24366, n24367, n24368, n24369, n24370,
         n24371, n24372, n24373, n24374, n24375, n24376, n24377, n24378,
         n24379, n24380, n24381, n24382, n24383, n24384, n24385, n24386,
         n24387, n24388, n24389, n24390, n24391, n24392, n24393, n24394,
         n24395, n24396, n24397, n24398, n24399, n24400, n24401, n24402,
         n24403, n24404, n24405, n24406, n24407, n24408, n24409, n24410,
         n24411, n24412, n24413, n24414, n24415, n24416, n24417, n24418,
         n24419, n24420, n24421, n24422, n24423, n24424, n24425, n24426,
         n24427, n24428, n24429, n24430, n24431, n24432, n24433, n24434,
         n24435, n24436, n24437, n24438, n24439, n24440, n24441, n24442,
         n24443, n24444, n24445, n24446, n24447, n24448, n24449, n24450,
         n24451, n24452, n24453, n24454, n24455, n24456, n24457, n24458,
         n24459, n24460, n24461, n24462, n24463, n24464, n24465, n24466,
         n24467, n24468, n24469, n24470, n24471, n24472, n24473, n24474,
         n24475, n24476, n24477, n24478, n24479, n24480, n24481, n24482,
         n24483, n24484, n24485, n24486, n24487, n24488, n24489, n24490,
         n24491, n24492, n24493, n24494, n24495, n24496, n24497, n24498,
         n24499, n24500, n24501, n24502, n24503, n24504, n24505, n24506,
         n24507, n24508, n24509, n24510, n24511, n24512, n24513, n24514,
         n24515, n24516, n24517, n24518, n24519, n24520, n24521, n24522,
         n24523, n24524, n24525, n24526, n24527, n24528, n24529, n24530,
         n24531, n24532, n24533, n24534, n24535, n24536, n24537, n24538,
         n24539, n24540, n24541, n24542, n24543, n24544, n24545, n24546,
         n24547, n24548, n24549, n24550, n24551, n24552, n24553, n24554,
         n24555, n24556, n24557, n24558, n24559, n24560, n24561, n24562,
         n24563, n24564, n24565, n24566, n24567, n24568, n24569, n24570,
         n24571, n24572, n24573, n24574, n24575, n24576, n24577, n24578,
         n24579, n24580, n24581, n24582, n24583, n24584, n24585, n24586,
         n24587, n24588, n24589, n24590, n24591, n24592, n24593, n24594,
         n24595, n24596, n24597, n24598, n24599, n24600, n24601, n24602,
         n24603, n24604, n24605, n24606, n24607, n24608, n24609, n24610,
         n24611, n24612, n24613, n24614, n24615, n24616, n24617, n24618,
         n24619, n24620, n24621, n24622, n24623, n24624, n24625, n24626,
         n24627, n24628, n24629, n24630, n24631, n24632, n24633, n24634,
         n24635, n24636, n24637, n24638, n24639, n24640, n24641, n24642,
         n24643, n24644, n24645, n24646, n24647, n24648, n24649, n24650,
         n24651, n24652, n24653, n24654, n24655, n24656, n24657, n24658,
         n24659, n24660, n24661, n24662, n24663, n24664, n24665, n24666,
         n24667, n24668, n24669, n24670, n24671, n24672, n24673, n24674,
         n24675, n24676, n24677, n24678, n24679, n24680, n24681, n24682,
         n24683, n24684, n24685, n24686, n24687, n24688, n24689, n24690,
         n24691, n24692, n24693, n24694, n24695, n24696, n24697, n24698,
         n24699, n24700, n24701, n24702, n24703, n24704, n24705, n24706,
         n24707, n24708, n24709, n24710, n24711, n24712, n24713, n24714,
         n24715, n24716, n24717, n24718, n24719, n24720, n24721, n24722,
         n24723, n24724, n24725, n24726, n24727, n24728, n24729, n24730,
         n24731, n24732, n24733, n24734, n24735, n24736, n24737, n24738,
         n24739, n24740, n24741, n24742, n24743, n24744, n24745, n24746,
         n24747, n24748, n24749, n24750, n24751, n24752, n24753, n24754,
         n24755, n24756, n24757, n24758, n24759, n24760, n24761, n24762,
         n24763, n24764, n24765, n24766, n24767, n24768, n24769, n24770,
         n24771, n24772, n24773, n24774, n24775, n24776, n24777, n24778,
         n24779, n24780, n24781, n24782, n24783, n24784, n24785, n24786,
         n24787, n24788, n24789, n24790, n24791, n24792, n24793, n24794,
         n24795, n24796, n24797, n24798, n24799, n24800, n24801, n24802,
         n24803, n24804, n24805, n24806, n24807, n24808, n24809, n24810,
         n24811, n24812, n24813, n24814, n24815, n24816, n24817, n24818,
         n24819, n24820, n24821, n24822, n24823, n24824, n24825, n24826,
         n24827, n24828, n24829, n24830, n24831, n24832, n24833, n24834,
         n24835, n24836, n24837, n24838, n24839, n24840, n24841, n24842,
         n24843, n24844, n24845, n24846, n24847, n24848, n24849, n24850,
         n24851, n24852, n24853, n24854, n24855, n24856, n24857, n24858,
         n24859, n24860, n24861, n24862, n24863, n24864, n24865, n24866,
         n24867, n24868, n24869, n24870, n24871, n24872, n24873, n24874,
         n24875, n24876, n24877, n24878, n24879, n24880, n24881, n24882,
         n24883, n24884, n24885, n24886, n24887, n24888, n24889, n24890,
         n24891, n24892, n24893, n24894, n24895, n24896, n24897, n24898,
         n24899, n24900, n24901, n24902, n24903, n24904, n24905, n24906,
         n24907, n24908, n24909, n24910, n24911, n24912, n24913, n24914,
         n24915, n24916, n24917, n24918, n24919, n24920, n24921, n24922,
         n24923, n24924, n24925, n24926, n24927, n24928, n24929, n24930,
         n24931, n24932, n24933, n24934, n24935, n24936, n24937, n24938,
         n24939, n24940, n24941, n24942, n24943, n24944, n24945, n24946,
         n24947, n24948, n24949, n24950, n24951, n24952, n24953, n24954,
         n24955, n24956, n24957, n24958, n24959, n24960, n24961, n24962,
         n24963, n24964, n24965, n24966, n24967, n24968, n24969, n24970,
         n24971, n24972, n24973, n24974, n24975, n24976, n24977, n24978,
         n24979, n24980, n24981, n24982, n24983, n24984, n24985, n24986,
         n24987, n24988, n24989, n24990, n24991, n24992, n24993, n24994,
         n24995, n24996, n24997, n24998, n24999, n25000, n25001, n25002,
         n25003, n25004, n25005, n25006, n25007, n25008, n25009, n25010,
         n25011, n25012, n25013, n25014, n25015, n25016, n25017, n25018,
         n25019, n25020, n25021, n25022, n25023, n25024, n25025, n25026,
         n25027, n25028, n25029, n25030, n25031, n25032, n25033, n25034,
         n25035, n25036, n25037, n25038, n25039, n25040, n25041, n25042,
         n25043, n25044, n25045, n25046, n25047, n25048, n25049, n25050,
         n25051, n25052, n25053, n25054, n25055, n25056, n25057, n25058,
         n25059, n25060, n25061, n25062, n25063, n25064, n25065, n25066,
         n25067, n25068, n25069, n25070, n25071, n25072, n25073, n25074,
         n25075, n25076, n25077, n25078, n25079, n25080, n25081, n25082,
         n25083, n25084, n25085, n25086, n25087, n25088, n25089, n25090,
         n25091, n25092, n25093, n25094, n25095, n25096, n25097, n25098,
         n25099, n25100, n25101, n25102, n25103, n25104, n25105, n25106,
         n25107, n25108, n25109, n25110, n25111, n25112, n25113, n25114,
         n25115, n25116, n25117, n25118, n25119, n25120, n25121, n25122,
         n25123, n25124, n25125, n25126, n25127, n25128, n25129, n25130,
         n25131, n25132, n25133, n25134, n25135, n25136, n25137, n25138,
         n25139, n25140, n25141, n25142, n25143, n25144, n25145, n25146,
         n25147, n25148, n25149, n25150, n25151, n25152, n25153, n25154,
         n25155, n25156, n25157, n25158, n25159, n25160, n25161, n25162,
         n25163, n25164, n25165, n25166, n25167, n25168, n25169, n25170,
         n25171, n25172, n25173, n25174, n25175, n25176, n25177, n25178,
         n25179, n25180, n25181, n25182, n25183, n25184, n25185, n25186,
         n25187, n25188, n25189, n25190, n25191, n25192, n25193, n25194,
         n25195, n25196, n25197, n25198, n25199, n25200, n25201, n25202,
         n25203, n25204, n25205, n25206, n25207, n25208, n25209, n25210,
         n25211, n25212, n25213, n25214, n25215, n25216, n25217, n25218,
         n25219, n25220, n25221, n25222, n25223, n25224, n25225, n25226,
         n25227, n25228, n25229, n25230, n25231, n25232, n25233, n25234,
         n25235, n25236, n25237, n25238, n25239, n25240, n25241, n25242,
         n25243, n25244, n25245, n25246, n25247, n25248, n25249, n25250,
         n25251, n25252, n25253, n25254, n25255, n25256, n25257, n25258,
         n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266,
         n25267, n25268, n25269, n25270, n25271, n25272, n25273, n25274,
         n25275, n25276, n25277, n25278, n25279, n25280, n25281, n25282,
         n25283, n25284, n25285, n25286, n25287, n25288, n25289, n25290,
         n25291, n25292, n25293, n25294, n25295, n25296, n25297, n25298,
         n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25306,
         n25307, n25308, n25309, n25310, n25311, n25312, n25313, n25314,
         n25315, n25316, n25317, n25318, n25319, n25320, n25321, n25322,
         n25323, n25324, n25325, n25326, n25327, n25328, n25329, n25330,
         n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338,
         n25339, n25340, n25341, n25342, n25343, n25344, n25345, n25346,
         n25347, n25348, n25349, n25350, n25351, n25352, n25353, n25354,
         n25355, n25356, n25357, n25358, n25359, n25360, n25361, n25362,
         n25363, n25364, n25365, n25366, n25367, n25368, n25369, n25370,
         n25371, n25372, n25373, n25374, n25375, n25376, n25377, n25378,
         n25379, n25380, n25381, n25382, n25383, n25384, n25385, n25386,
         n25387, n25388, n25389, n25390, n25391, n25392, n25393, n25394,
         n25395, n25396, n25397, n25398, n25399, n25400, n25401, n25402,
         n25403, n25404, n25405, n25406, n25407, n25408, n25409, n25410,
         n25411, n25412, n25413, n25414, n25415, n25416, n25417, n25418,
         n25419, n25420, n25421, n25422, n25423, n25424, n25425, n25426,
         n25427, n25428, n25429, n25430, n25431, n25432, n25433, n25434,
         n25435, n25436, n25437, n25438, n25439, n25440, n25441, n25442,
         n25443, n25444, n25445, n25446, n25447, n25448, n25449, n25450,
         n25451, n25452, n25453, n25454, n25455, n25456, n25457, n25458,
         n25459, n25460, n25461, n25462, n25463, n25464, n25465, n25466,
         n25467, n25468, n25469, n25470, n25471, n25472, n25473, n25474,
         n25475, n25476, n25477, n25478, n25479, n25480, n25481, n25482,
         n25483, n25484, n25485, n25486, n25487, n25488, n25489, n25490,
         n25491, n25492, n25493, n25494, n25495, n25496, n25497, n25498,
         n25499, n25500, n25501, n25502, n25503, n25504, n25505, n25506,
         n25507, n25508, n25509, n25510, n25511, n25512, n25513, n25514,
         n25515, n25516, n25517, n25518, n25519, n25520, n25521, n25522,
         n25523, n25524, n25525, n25526, n25527, n25528, n25529, n25530,
         n25531, n25532, n25533, n25534, n25535, n25536, n25537, n25538,
         n25539, n25540, n25541, n25542, n25543, n25544, n25545, n25546,
         n25547, n25548, n25549, n25550, n25551, n25552, n25553, n25554,
         n25555, n25556, n25557, n25558, n25559, n25560, n25561, n25562,
         n25563, n25564, n25565, n25566, n25567, n25568, n25569, n25570,
         n25571, n25572, n25573, n25574, n25575, n25576, n25577, n25578,
         n25579, n25580, n25581, n25582, n25583, n25584, n25585, n25586,
         n25587, n25588, n25589, n25590, n25591, n25592, n25593, n25594,
         n25595, n25596, n25597, n25598, n25599, n25600, n25601, n25602,
         n25603, n25604, n25605, n25606, n25607, n25608, n25609, n25610,
         n25611, n25612, n25613, n25614, n25615, n25616, n25617, n25618,
         n25619, n25620, n25621, n25622, n25623, n25624, n25625, n25626,
         n25627, n25628, n25629, n25630, n25631, n25632, n25633, n25634,
         n25635, n25636, n25637, n25638, n25639, n25640, n25641, n25642,
         n25643, n25644, n25645, n25646, n25647, n25648, n25649, n25650,
         n25651, n25652, n25653, n25654, n25655, n25656, n25657, n25658,
         n25659, n25660, n25661, n25662, n25663, n25664, n25665, n25666,
         n25667, n25668, n25669, n25670, n25671, n25672, n25673, n25674,
         n25675, n25676, n25677, n25678, n25679, n25680, n25681, n25682,
         n25683, n25684, n25685, n25686, n25687, n25688, n25689, n25690,
         n25691, n25692, n25693, n25694, n25695, n25696, n25697, n25698,
         n25699, n25700, n25701, n25702, n25703, n25704, n25705, n25706,
         n25707, n25708, n25709, n25710, n25711, n25712, n25713, n25714,
         n25715, n25716, n25717, n25718, n25719, n25720, n25721, n25722,
         n25723, n25724, n25725, n25726, n25727, n25728, n25729, n25730,
         n25731, n25732, n25733, n25734, n25735, n25736, n25737, n25738,
         n25739, n25740, n25741, n25742, n25743, n25744, n25745, n25746,
         n25747, n25748, n25749, n25750, n25751, n25752, n25753, n25754,
         n25755, n25756, n25757, n25758, n25759, n25760, n25761, n25762,
         n25763, n25764, n25765, n25766, n25767, n25768, n25769, n25770,
         n25771, n25772, n25773, n25774, n25775, n25776, n25777, n25778,
         n25779, n25780, n25781, n25782, n25783, n25784, n25785, n25786,
         n25787, n25788, n25789, n25790, n25791, n25792, n25793, n25794,
         n25795, n25796, n25797, n25798, n25799, n25800, n25801, n25802,
         n25803, n25804, n25805, n25806, n25807, n25808, n25809, n25810,
         n25811, n25812, n25813, n25814, n25815, n25816, n25817, n25818,
         n25819, n25820, n25821, n25822, n25823, n25824, n25825, n25826,
         n25827, n25828, n25829, n25830, n25831, n25832, n25833, n25834,
         n25835, n25836, n25837, n25838, n25839, n25840, n25841, n25842,
         n25843, n25844, n25845, n25846, n25847, n25848, n25849, n25850,
         n25851, n25852, n25853, n25854, n25855, n25856, n25857, n25858,
         n25859, n25860, n25861, n25862, n25863, n25864, n25865, n25866,
         n25867, n25868, n25869, n25870, n25871, n25872, n25873, n25874,
         n25875, n25876, n25877, n25878, n25879, n25880, n25881, n25882,
         n25883, n25884, n25885, n25886, n25887, n25888, n25889, n25890,
         n25891, n25892, n25893, n25894, n25895, n25896, n25897, n25898,
         n25899, n25900, n25901, n25902, n25903, n25904, n25905, n25906,
         n25907, n25908, n25909, n25910, n25911, n25912, n25913, n25914,
         n25915, n25916, n25917, n25918, n25919, n25920, n25921, n25922,
         n25923, n25924, n25925, n25926, n25927, n25928, n25929, n25930,
         n25931, n25932, n25933, n25934, n25935, n25936, n25937, n25938,
         n25939, n25940, n25941, n25942, n25943, n25944, n25945, n25946,
         n25947, n25948, n25949, n25950, n25951, n25952, n25953, n25954,
         n25955, n25956, n25957, n25958, n25959, n25960, n25961, n25962,
         n25963, n25964, n25965, n25966, n25967, n25968, n25969, n25970,
         n25971, n25972, n25973, n25974, n25975, n25976, n25977, n25978,
         n25979, n25980, n25981, n25982, n25983, n25984, n25985, n25986,
         n25987, n25988, n25989, n25990, n25991, n25992, n25993, n25994,
         n25995, n25996, n25997, n25998, n25999, n26000, n26001, n26002,
         n26003, n26004, n26005, n26006, n26007, n26008, n26009, n26010,
         n26011, n26012, n26013, n26014, n26015, n26016, n26017, n26018,
         n26019, n26020, n26021, n26022, n26023, n26024, n26025, n26026,
         n26027, n26028, n26029, n26030, n26031, n26032, n26033, n26034,
         n26035, n26036, n26037, n26038, n26039, n26040, n26041, n26042,
         n26043, n26044, n26045, n26046, n26047, n26048, n26049, n26050,
         n26051, n26052, n26053, n26054, n26055, n26056, n26057, n26058,
         n26059, n26060, n26061, n26062, n26063, n26064, n26065, n26066,
         n26067, n26068, n26069, n26070, n26071, n26072, n26073, n26074,
         n26075, n26076, n26077, n26078, n26079, n26080, n26081, n26082,
         n26083, n26084, n26085, n26086, n26087, n26088, n26089, n26090,
         n26091, n26092, n26093, n26094, n26095, n26096, n26097, n26098,
         n26099, n26100, n26101, n26102, n26103, n26104, n26105, n26106,
         n26107, n26108, n26109, n26110, n26111, n26112, n26113, n26114,
         n26115, n26116, n26117, n26118, n26119, n26120, n26121, n26122,
         n26123, n26124, n26125, n26126, n26127, n26128, n26129, n26130,
         n26131, n26132, n26133, n26134, n26135, n26136, n26137, n26138,
         n26139, n26140, n26141, n26142, n26143, n26144, n26145, n26146,
         n26147, n26148, n26149, n26150, n26151, n26152, n26153, n26154,
         n26155, n26156, n26157, n26158, n26159, n26160, n26161, n26162,
         n26163, n26164, n26165, n26166, n26167, n26168, n26169, n26170,
         n26171, n26172, n26173, n26174, n26175, n26176, n26177, n26178,
         n26179, n26180, n26181, n26182, n26183, n26184, n26185, n26186,
         n26187, n26188, n26189, n26190, n26191, n26192, n26193, n26194,
         n26195, n26196, n26197, n26198, n26199, n26200, n26201, n26202,
         n26203, n26204, n26205, n26206, n26207, n26208, n26209, n26210,
         n26211, n26212, n26213, n26214, n26215, n26216, n26217, n26218,
         n26219, n26220, n26221, n26222, n26223, n26224, n26225, n26226,
         n26227, n26228, n26229, n26230, n26231, n26232, n26233, n26234,
         n26235, n26236, n26237, n26238, n26239, n26240, n26241, n26242,
         n26243, n26244, n26245, n26246, n26247, n26248, n26249, n26250,
         n26251, n26252, n26253, n26254, n26255, n26256, n26257, n26258,
         n26259, n26260, n26261, n26262, n26263, n26264, n26265, n26266,
         n26267, n26268, n26269, n26270, n26271, n26272, n26273, n26274,
         n26275, n26276, n26277, n26278, n26279, n26280, n26281, n26282,
         n26283, n26284, n26285, n26286, n26287, n26288, n26289, n26290,
         n26291, n26292, n26293, n26294, n26295, n26296, n26297, n26298,
         n26299, n26300, n26301, n26302, n26303, n26304, n26305, n26306,
         n26307, n26308, n26309, n26310, n26311, n26312, n26313, n26314,
         n26315, n26316, n26317, n26318, n26319, n26320, n26321, n26322,
         n26323, n26324, n26325, n26326, n26327, n26328, n26329, n26330,
         n26331, n26332, n26333, n26334, n26335, n26336, n26337, n26338,
         n26339, n26340, n26341, n26342, n26343, n26344, n26345, n26346,
         n26347, n26348, n26349, n26350, n26351, n26352, n26353, n26354,
         n26355, n26356, n26357, n26358, n26359, n26360, n26361, n26362,
         n26363, n26364, n26365, n26366, n26367, n26368, n26369, n26370,
         n26371, n26372, n26373, n26374, n26375, n26376, n26377, n26378,
         n26379, n26380, n26381, n26382, n26383, n26384, n26385, n26386,
         n26387, n26388, n26389, n26390, n26391, n26392, n26393, n26394,
         n26395, n26396, n26397, n26398, n26399, n26400, n26401, n26402,
         n26403, n26404, n26405, n26406, n26407, n26408, n26409, n26410,
         n26411, n26412, n26413, n26414, n26415, n26416, n26417, n26418,
         n26419, n26420, n26421, n26422, n26423, n26424, n26425, n26426,
         n26427, n26428, n26429, n26430, n26431, n26432, n26433, n26434,
         n26435, n26436, n26437, n26438, n26439, n26440, n26441, n26442,
         n26443, n26444, n26445, n26446, n26447, n26448, n26449, n26450,
         n26451, n26452, n26453, n26454, n26455, n26456, n26457, n26458,
         n26459, n26460, n26461, n26462, n26463, n26464, n26465, n26466,
         n26467, n26468, n26469, n26470, n26471, n26472, n26473, n26474,
         n26475, n26476, n26477, n26478, n26479, n26480, n26481, n26482,
         n26483, n26484, n26485, n26486, n26487, n26488, n26489, n26490,
         n26491, n26492, n26493, n26494, n26495, n26496, n26497, n26498,
         n26499, n26500, n26501, n26502, n26503, n26504, n26505, n26506,
         n26507, n26508, n26509, n26510, n26511, n26512, n26513, n26514,
         n26515, n26516, n26517, n26518, n26519, n26520, n26521, n26522,
         n26523, n26524, n26525, n26526, n26527, n26528, n26529, n26530,
         n26531, n26532, n26533, n26534, n26535, n26536, n26537, n26538,
         n26539, n26540, n26541, n26542, n26543, n26544, n26545, n26546,
         n26547, n26548, n26549, n26550, n26551, n26552, n26553, n26554,
         n26555, n26556, n26557, n26558, n26559, n26560, n26561, n26562,
         n26563, n26564, n26565, n26566, n26567, n26568, n26569, n26570,
         n26571, n26572, n26573, n26574, n26575, n26576, n26577, n26578,
         n26579, n26580, n26581, n26582, n26583, n26584, n26585, n26586,
         n26587, n26588, n26589, n26590, n26591, n26592, n26593, n26594,
         n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602,
         n26603, n26604, n26605, n26606, n26607, n26608, n26609, n26610,
         n26611, n26612, n26613, n26614, n26615, n26616, n26617, n26618,
         n26619, n26620, n26621, n26622, n26623, n26624, n26625, n26626,
         n26627, n26628, n26629, n26630, n26631, n26632, n26633, n26634,
         n26635, n26636, n26637, n26638, n26639, n26640, n26641, n26642,
         n26643, n26644, n26645, n26646, n26647, n26648, n26649, n26650,
         n26651, n26652, n26653, n26654, n26655, n26656, n26657, n26658,
         n26659, n26660, n26661, n26662, n26663, n26664, n26665, n26666,
         n26667, n26668, n26669, n26670, n26671, n26672, n26673, n26674,
         n26675, n26676, n26677, n26678, n26679, n26680, n26681, n26682,
         n26683, n26684, n26685, n26686, n26687, n26688, n26689, n26690,
         n26691, n26692, n26693, n26694, n26695, n26696, n26697, n26698,
         n26699, n26700, n26701, n26702, n26703, n26704, n26705, n26706,
         n26707, n26708, n26709, n26710, n26711, n26712, n26713, n26714,
         n26715, n26716, n26717, n26718, n26719, n26720, n26721, n26722,
         n26723, n26724, n26725, n26726, n26727, n26728, n26729, n26730,
         n26731, n26732, n26733, n26734, n26735, n26736, n26737, n26738,
         n26739, n26740, n26741, n26742, n26743, n26744, n26745, n26746,
         n26747, n26748, n26749, n26750, n26751, n26752, n26753, n26754,
         n26755, n26756, n26757, n26758, n26759, n26760, n26761, n26762,
         n26763, n26764, n26765, n26766, n26767, n26768, n26769, n26770,
         n26771, n26772, n26773, n26774, n26775, n26776, n26777, n26778,
         n26779, n26780, n26781, n26782, n26783, n26784, n26785, n26786,
         n26787, n26788, n26789, n26790, n26791, n26792, n26793, n26794,
         n26795, n26796, n26797, n26798, n26799, n26800, n26801, n26802,
         n26803, n26804, n26805, n26806, n26807, n26808, n26809, n26810,
         n26811, n26812, n26813, n26814, n26815, n26816, n26817, n26818,
         n26819, n26820, n26821, n26822, n26823, n26824, n26825, n26826,
         n26827, n26828, n26829, n26830, n26831, n26832, n26833, n26834,
         n26835, n26836, n26837, n26838, n26839, n26840, n26841, n26842,
         n26843, n26844, n26845, n26846, n26847, n26848, n26849, n26850,
         n26851, n26852, n26853, n26854, n26855, n26856, n26857, n26858,
         n26859, n26860, n26861, n26862, n26863, n26864, n26865, n26866,
         n26867, n26868, n26869, n26870, n26871, n26872, n26873, n26874,
         n26875, n26876, n26877, n26878, n26879, n26880, n26881, n26882,
         n26883, n26884, n26885, n26886, n26887, n26888, n26889, n26890,
         n26891, n26892, n26893, n26894, n26895, n26896, n26897, n26898,
         n26899, n26900, n26901, n26902, n26903, n26904, n26905, n26906,
         n26907, n26908, n26909, n26910, n26911, n26912, n26913, n26914,
         n26915, n26916, n26917, n26918, n26919, n26920, n26921, n26922,
         n26923, n26924, n26925, n26926, n26927, n26928, n26929, n26930,
         n26931, n26932, n26933, n26934, n26935, n26936, n26937, n26938,
         n26939, n26940, n26941, n26942, n26943, n26944, n26945, n26946,
         n26947, n26948, n26949, n26950, n26951, n26952, n26953, n26954,
         n26955, n26956, n26957, n26958, n26959, n26960, n26961, n26962,
         n26963, n26964, n26965, n26966, n26967, n26968, n26969, n26970,
         n26971, n26972, n26973, n26974, n26975, n26976, n26977, n26978,
         n26979, n26980, n26981, n26982, n26983, n26984, n26985, n26986,
         n26987, n26988, n26989, n26990, n26991, n26992, n26993, n26994,
         n26995, n26996, n26997, n26998, n26999, n27000, n27001, n27002,
         n27003, n27004, n27005, n27006, n27007, n27008, n27009, n27010,
         n27011, n27012, n27013, n27014, n27015, n27016, n27017, n27018,
         n27019, n27020, n27021, n27022, n27023, n27024, n27025, n27026,
         n27027, n27028, n27029, n27030, n27031, n27032, n27033, n27034,
         n27035, n27036, n27037, n27038, n27039, n27040, n27041, n27042,
         n27043, n27044, n27045, n27046, n27047, n27048, n27049, n27050,
         n27051, n27052, n27053, n27054, n27055, n27056, n27057, n27058,
         n27059, n27060, n27061, n27062, n27063, n27064, n27065, n27066,
         n27067, n27068, n27069, n27070, n27071, n27072, n27073, n27074,
         n27075, n27076, n27077, n27078, n27079, n27080, n27081, n27082,
         n27083, n27084, n27085, n27086, n27087, n27088, n27089, n27090,
         n27091, n27092, n27093, n27094, n27095, n27096, n27097, n27098,
         n27099, n27100, n27101, n27102, n27103, n27104, n27105, n27106,
         n27107, n27108, n27109, n27110, n27111, n27112, n27113, n27114,
         n27115, n27116, n27117, n27118, n27119, n27120, n27121, n27122,
         n27123, n27124, n27125, n27126, n27127, n27128, n27129, n27130,
         n27131, n27132, n27133, n27134, n27135, n27136, n27137, n27138,
         n27139, n27140, n27141, n27142, n27143, n27144, n27145, n27146,
         n27147, n27148, n27149, n27150, n27151, n27152, n27153, n27154,
         n27155, n27156, n27157, n27158, n27159, n27160, n27161, n27162,
         n27163, n27164, n27165, n27166, n27167, n27168, n27169, n27170,
         n27171, n27172, n27173, n27174, n27175, n27176, n27177, n27178,
         n27179, n27180, n27181, n27182, n27183, n27184, n27185, n27186,
         n27187, n27188, n27189, n27190, n27191, n27192, n27193, n27194,
         n27195, n27196, n27197, n27198, n27199, n27200, n27201, n27202,
         n27203, n27204, n27205, n27206, n27207, n27208, n27209, n27210,
         n27211, n27212, n27213, n27214, n27215, n27216, n27217, n27218,
         n27219, n27220, n27221, n27222, n27223, n27224, n27225, n27226,
         n27227, n27228, n27229, n27230, n27231, n27232, n27233, n27234,
         n27235, n27236, n27237, n27238, n27239, n27240, n27241, n27242,
         n27243, n27244, n27245, n27246, n27247, n27248, n27249, n27250,
         n27251, n27252, n27253, n27254, n27255, n27256, n27257, n27258,
         n27259, n27260, n27261, n27262, n27263, n27264, n27265, n27266,
         n27267, n27268, n27269, n27270, n27271, n27272, n27273, n27274,
         n27275, n27276, n27277, n27278, n27279, n27280, n27281, n27282,
         n27283, n27284, n27285, n27286, n27287, n27288, n27289, n27290,
         n27291, n27292, n27293, n27294, n27295, n27296, n27297, n27298,
         n27299, n27300, n27301, n27302, n27303, n27304, n27305, n27306,
         n27307, n27308, n27309, n27310, n27311, n27312, n27313, n27314,
         n27315, n27316, n27317, n27318, n27319, n27320, n27321, n27322,
         n27323, n27324, n27325, n27326, n27327, n27328, n27329, n27330,
         n27331, n27332, n27333, n27334, n27335, n27336, n27337, n27338,
         n27339, n27340, n27341, n27342, n27343, n27344, n27345, n27346,
         n27347, n27348, n27349, n27350, n27351, n27352, n27353, n27354,
         n27355, n27356, n27357, n27358, n27359, n27360, n27361, n27362,
         n27363, n27364, n27365, n27366, n27367, n27368, n27369, n27370,
         n27371, n27372, n27373, n27374, n27375, n27376, n27377, n27378,
         n27379, n27380, n27381, n27382, n27383, n27384, n27385, n27386,
         n27387, n27388, n27389, n27390, n27391, n27392, n27393, n27394,
         n27395, n27396, n27397, n27398, n27399, n27400, n27401, n27402,
         n27403, n27404, n27405, n27406, n27407, n27408, n27409, n27410,
         n27411, n27412, n27413, n27414, n27415, n27416, n27417, n27418,
         n27419, n27420, n27421, n27422, n27423, n27424, n27425, n27426,
         n27427, n27428, n27429, n27430, n27431, n27432, n27433, n27434,
         n27435, n27436, n27437, n27438, n27439, n27440, n27441, n27442,
         n27443, n27444, n27445, n27446, n27447, n27448, n27449, n27450,
         n27451, n27452, n27453, n27454, n27455, n27456, n27457, n27458,
         n27459, n27460, n27461, n27462, n27463, n27464, n27465, n27466,
         n27467, n27468, n27469, n27470, n27471, n27472, n27473, n27474,
         n27475, n27476, n27477, n27478, n27479, n27480, n27481, n27482,
         n27483, n27484, n27485, n27486, n27487, n27488, n27489, n27490,
         n27491, n27492, n27493, n27494, n27495, n27496, n27497, n27498,
         n27499, n27500, n27501, n27502, n27503, n27504, n27505, n27506,
         n27507, n27508, n27509, n27510, n27511, n27512, n27513, n27514,
         n27515, n27516, n27517, n27518, n27519, n27520, n27521, n27522,
         n27523, n27524, n27525, n27526, n27527, n27528, n27529, n27530,
         n27531, n27532, n27533, n27534, n27535, n27536, n27537, n27538,
         n27539, n27540, n27541, n27542, n27543, n27544, n27545, n27546,
         n27547, n27548, n27549, n27550, n27551, n27552, n27553, n27554,
         n27555, n27556, n27557, n27558, n27559, n27560, n27561, n27562,
         n27563, n27564, n27565, n27566, n27567, n27568, n27569, n27570,
         n27571, n27572, n27573, n27574, n27575, n27576, n27577, n27578,
         n27579, n27580, n27581, n27582, n27583, n27584, n27585, n27586,
         n27587, n27588, n27589, n27590, n27591, n27592, n27593, n27594,
         n27595, n27596, n27597, n27598, n27599, n27600, n27601, n27602,
         n27603, n27604, n27605, n27606, n27607, n27608, n27609, n27610,
         n27611, n27612, n27613, n27614, n27615, n27616, n27617, n27618,
         n27619, n27620, n27621, n27622, n27623, n27624, n27625, n27626,
         n27627, n27628, n27629, n27630, n27631, n27632, n27633, n27634,
         n27635, n27636, n27637, n27638, n27639, n27640, n27641, n27642,
         n27643, n27644, n27645, n27646, n27647, n27648, n27649, n27650,
         n27651, n27652, n27653, n27654, n27655, n27656, n27657, n27658,
         n27659, n27660, n27661, n27662, n27663, n27664, n27665, n27666,
         n27667, n27668, n27669, n27670, n27671, n27672, n27673, n27674,
         n27675, n27676, n27677, n27678, n27679, n27680, n27681, n27682,
         n27683, n27684, n27685, n27686, n27687, n27688, n27689, n27690,
         n27691, n27692, n27693, n27694, n27695, n27696, n27697, n27698,
         n27699, n27700, n27701, n27702, n27703, n27704, n27705, n27706,
         n27707, n27708, n27709, n27710, n27711, n27712, n27713, n27714,
         n27715, n27716, n27717, n27718, n27719, n27720, n27721, n27722,
         n27723, n27724, n27725, n27726, n27727, n27728, n27729, n27730,
         n27731, n27732, n27733, n27734, n27735, n27736, n27737, n27738,
         n27739, n27740, n27741, n27742, n27743, n27744, n27745, n27746,
         n27747, n27748, n27749, n27750, n27751, n27752, n27753, n27754,
         n27755, n27756, n27757, n27758, n27759, n27760, n27761, n27762,
         n27763, n27764, n27765, n27766, n27767, n27768, n27769, n27770,
         n27771, n27772, n27773, n27774, n27775, n27776, n27777, n27778,
         n27779, n27780, n27781, n27782, n27783, n27784, n27785, n27786,
         n27787, n27788, n27789, n27790, n27791, n27792, n27793, n27794,
         n27795, n27796, n27797, n27798, n27799, n27800, n27801, n27802,
         n27803, n27804, n27805, n27806, n27807, n27808, n27809, n27810,
         n27811, n27812, n27813, n27814, n27815, n27816, n27817, n27818,
         n27819, n27820, n27821, n27822, n27823, n27824, n27825, n27826,
         n27827, n27828, n27829, n27830, n27831, n27832, n27833, n27834,
         n27835, n27836, n27837, n27838, n27839, n27840, n27841, n27842,
         n27843, n27844, n27845, n27846, n27847, n27848, n27849, n27850,
         n27851, n27852, n27853, n27854, n27855, n27856, n27857, n27858,
         n27859, n27860, n27861, n27862, n27863, n27864, n27865, n27866,
         n27867, n27868, n27869, n27870, n27871, n27872, n27873, n27874,
         n27875, n27876, n27877, n27878, n27879, n27880, n27881, n27882,
         n27883, n27884, n27885, n27886, n27887, n27888, n27889, n27890,
         n27891, n27892, n27893, n27894, n27895, n27896, n27897, n27898,
         n27899, n27900, n27901, n27902, n27903, n27904, n27905, n27906,
         n27907, n27908, n27909, n27910, n27911, n27912, n27913, n27914,
         n27915, n27916, n27917, n27918, n27919, n27920, n27921, n27922,
         n27923, n27924, n27925, n27926, n27927, n27928, n27929, n27930,
         n27931, n27932, n27933, n27934, n27935, n27936, n27937, n27938,
         n27939, n27940, n27941, n27942, n27943, n27944, n27945, n27946,
         n27947, n27948, n27949, n27950, n27951, n27952, n27953, n27954,
         n27955, n27956, n27957, n27958, n27959, n27960, n27961, n27962,
         n27963, n27964, n27965, n27966, n27967, n27968, n27969, n27970,
         n27971, n27972, n27973, n27974, n27975, n27976, n27977, n27978,
         n27979, n27980, n27981, n27982, n27983, n27984, n27985, n27986,
         n27987, n27988, n27989, n27990, n27991, n27992, n27993, n27994,
         n27995, n27996, n27997, n27998, n27999, n28000, n28001, n28002,
         n28003, n28004, n28005, n28006, n28007, n28008, n28009, n28010,
         n28011, n28012, n28013, n28014, n28015, n28016, n28017, n28018,
         n28019, n28020, n28021, n28022, n28023, n28024, n28025, n28026,
         n28027, n28028, n28029, n28030, n28031, n28032, n28033, n28034,
         n28035, n28036, n28037, n28038, n28039, n28040, n28041, n28042,
         n28043, n28044, n28045, n28046, n28047, n28048, n28049, n28050,
         n28051, n28052, n28053, n28054, n28055, n28056, n28057, n28058,
         n28059, n28060, n28061, n28062, n28063, n28064, n28065, n28066,
         n28067, n28068, n28069, n28070, n28071, n28072, n28073, n28074,
         n28075, n28076, n28077, n28078, n28079, n28080, n28081, n28082,
         n28083, n28084, n28085, n28086, n28087, n28088, n28089, n28090,
         n28091, n28092, n28093, n28094, n28095, n28096, n28097, n28098,
         n28099, n28100, n28101, n28102, n28103, n28104, n28105, n28106,
         n28107, n28108, n28109, n28110, n28111, n28112, n28113, n28114,
         n28115, n28116, n28117, n28118, n28119, n28120, n28121, n28122,
         n28123, n28124, n28125, n28126, n28127, n28128, n28129, n28130,
         n28131, n28132, n28133, n28134, n28135, n28136, n28137, n28138,
         n28139, n28140, n28141, n28142, n28143, n28144, n28145, n28146,
         n28147, n28148, n28149, n28150, n28151, n28152, n28153, n28154,
         n28155, n28156, n28157, n28158, n28159, n28160, n28161, n28162,
         n28163, n28164, n28165, n28166, n28167, n28168, n28169, n28170,
         n28171, n28172, n28173, n28174, n28175, n28176, n28177, n28178,
         n28179, n28180, n28181, n28182, n28183, n28184, n28185, n28186,
         n28187, n28188, n28189, n28190, n28191, n28192, n28193, n28194,
         n28195, n28196, n28197, n28198, n28199, n28200, n28201, n28202,
         n28203, n28204, n28205, n28206, n28207, n28208, n28209, n28210,
         n28211, n28212, n28213, n28214, n28215, n28216, n28217, n28218,
         n28219, n28220, n28221, n28222, n28223, n28224, n28225, n28226,
         n28227, n28228, n28229, n28230, n28231, n28232, n28233, n28234,
         n28235, n28236, n28237, n28238, n28239, n28240, n28241, n28242,
         n28243, n28244, n28245, n28246, n28247, n28248, n28249, n28250,
         n28251, n28252, n28253, n28254, n28255, n28256, n28257, n28258,
         n28259, n28260, n28261, n28262, n28263, n28264, n28265, n28266,
         n28267, n28268, n28269, n28270, n28271, n28272, n28273, n28274,
         n28275, n28276, n28277, n28278, n28279, n28280, n28281, n28282,
         n28283, n28284, n28285, n28286, n28287, n28288, n28289, n28290,
         n28291, n28292, n28293, n28294, n28295, n28296, n28297, n28298,
         n28299, n28300, n28301, n28302, n28303, n28304, n28305, n28306,
         n28307, n28308, n28309, n28310, n28311, n28312, n28313, n28314,
         n28315, n28316, n28317, n28318, n28319, n28320, n28321, n28322,
         n28323, n28324, n28325, n28326, n28327, n28328, n28329, n28330,
         n28331, n28332, n28333, n28334, n28335, n28336, n28337, n28338,
         n28339, n28340, n28341, n28342, n28343, n28344, n28345, n28346,
         n28347, n28348, n28349, n28350, n28351, n28352, n28353, n28354,
         n28355, n28356, n28357, n28358, n28359, n28360, n28361, n28362,
         n28363, n28364, n28365, n28366, n28367, n28368, n28369, n28370,
         n28371, n28372, n28373, n28374, n28375, n28376, n28377, n28378,
         n28379, n28380, n28381, n28382, n28383, n28384, n28385, n28386,
         n28387, n28388, n28389, n28390, n28391, n28392, n28393, n28394,
         n28395, n28396, n28397, n28398, n28399, n28400, n28401, n28402,
         n28403, n28404, n28405, n28406, n28407, n28408, n28409, n28410,
         n28411, n28412, n28413, n28414, n28415, n28416, n28417, n28418,
         n28419, n28420, n28421, n28422, n28423, n28424, n28425, n28426,
         n28427, n28428, n28429, n28430, n28431, n28432, n28433, n28434,
         n28435, n28436, n28437, n28438, n28439, n28440, n28441, n28442,
         n28443, n28444, n28445, n28446, n28447, n28448, n28449, n28450,
         n28451, n28452, n28453, n28454, n28455, n28456, n28457, n28458,
         n28459, n28460, n28461, n28462, n28463, n28464, n28465, n28466,
         n28467, n28468, n28469, n28470, n28471, n28472, n28473, n28474,
         n28475, n28476, n28477, n28478, n28479, n28480, n28481, n28482,
         n28483, n28484, n28485, n28486, n28487, n28488, n28489, n28490,
         n28491, n28492, n28493, n28494, n28495, n28496, n28497, n28498,
         n28499, n28500, n28501, n28502, n28503, n28504, n28505, n28506,
         n28507, n28508, n28509, n28510, n28511, n28512, n28513, n28514,
         n28515, n28516, n28517, n28518, n28519, n28520, n28521, n28522,
         n28523, n28524, n28525, n28526, n28527, n28528, n28529, n28530,
         n28531, n28532, n28533, n28534, n28535, n28536, n28537, n28538,
         n28539, n28540, n28541, n28542, n28543, n28544, n28545, n28546,
         n28547, n28548, n28549, n28550, n28551, n28552, n28553, n28554,
         n28555, n28556, n28557, n28558, n28559, n28560, n28561, n28562,
         n28563, n28564, n28565, n28566, n28567, n28568, n28569, n28570,
         n28571, n28572, n28573, n28574, n28575, n28576, n28577, n28578,
         n28579, n28580, n28581, n28582, n28583, n28584, n28585, n28586,
         n28587, n28588, n28589, n28590, n28591, n28592, n28593, n28594,
         n28595, n28596, n28597, n28598, n28599, n28600, n28601, n28602,
         n28603, n28604, n28605, n28606, n28607, n28608, n28609, n28610,
         n28611, n28612, n28613, n28614, n28615, n28616, n28617, n28618,
         n28619, n28620, n28621, n28622, n28623, n28624, n28625, n28626,
         n28627, n28628, n28629, n28630, n28631, n28632, n28633, n28634,
         n28635, n28636, n28637, n28638, n28639, n28640, n28641, n28642,
         n28643, n28644, n28645, n28646, n28647, n28648, n28649, n28650,
         n28651, n28652, n28653, n28654, n28655, n28656, n28657, n28658,
         n28659, n28660, n28661, n28662, n28663, n28664, n28665, n28666,
         n28667, n28668, n28669, n28670, n28671, n28672, n28673, n28674,
         n28675, n28676, n28677, n28678, n28679, n28680, n28681, n28682,
         n28683, n28684, n28685, n28686, n28687, n28688, n28689, n28690,
         n28691, n28692, n28693, n28694, n28695, n28696, n28697, n28698,
         n28699, n28700, n28701, n28702, n28703, n28704, n28705, n28706,
         n28707, n28708, n28709, n28710, n28711, n28712, n28713, n28714,
         n28715, n28716, n28717, n28718, n28719, n28720, n28721, n28722,
         n28723, n28724, n28725, n28726, n28727, n28728, n28729, n28730,
         n28731, n28732, n28733, n28734, n28735, n28736, n28737, n28738,
         n28739, n28740, n28741, n28742, n28743, n28744, n28745, n28746,
         n28747, n28748, n28749, n28750, n28751, n28752, n28753, n28754,
         n28755, n28756, n28757, n28758, n28759, n28760, n28761, n28762,
         n28763, n28764, n28765, n28766, n28767, n28768, n28769, n28770,
         n28771, n28772, n28773;

  DFF ebreg_reg ( .D(n5), .CLK(clk), .RST(rst), .Q(ebreg) );
  DFF greg_reg ( .D(n4), .CLK(clk), .RST(rst), .Q(g) );
  XNOR U10 ( .A(y[3121]), .B(x[3121]), .Z(n8) );
  XNOR U11 ( .A(x[3120]), .B(y[3120]), .Z(n9) );
  ANDN U12 ( .B(n11589), .A(n11586), .Z(n10) );
  XNOR U13 ( .A(y[3117]), .B(x[3117]), .Z(n11) );
  XNOR U14 ( .A(x[3116]), .B(y[3116]), .Z(n12) );
  NAND U15 ( .A(n9924), .B(n9923), .Z(n13) );
  AND U16 ( .A(n9925), .B(n13), .Z(n14) );
  NANDN U17 ( .A(n11591), .B(n14), .Z(n15) );
  NANDN U18 ( .A(n11593), .B(n15), .Z(n16) );
  NAND U19 ( .A(n12), .B(n16), .Z(n17) );
  NAND U20 ( .A(n17), .B(n11588), .Z(n18) );
  NAND U21 ( .A(n11), .B(n18), .Z(n19) );
  NAND U22 ( .A(n10), .B(n19), .Z(n20) );
  ANDN U23 ( .B(n20), .A(n18353), .Z(n21) );
  NANDN U24 ( .A(n11585), .B(n21), .Z(n22) );
  NANDN U25 ( .A(n11587), .B(n22), .Z(n23) );
  NAND U26 ( .A(n9), .B(n23), .Z(n24) );
  NAND U27 ( .A(n24), .B(n11582), .Z(n25) );
  NAND U28 ( .A(n8), .B(n25), .Z(n9926) );
  XNOR U29 ( .A(x[3166]), .B(y[3166]), .Z(n26) );
  XNOR U30 ( .A(y[3165]), .B(x[3165]), .Z(n27) );
  ANDN U31 ( .B(n11544), .A(n11539), .Z(n28) );
  XNOR U32 ( .A(x[3162]), .B(y[3162]), .Z(n29) );
  XNOR U33 ( .A(y[3161]), .B(x[3161]), .Z(n30) );
  NAND U34 ( .A(n9986), .B(n9985), .Z(n31) );
  AND U35 ( .A(n9987), .B(n31), .Z(n32) );
  NANDN U36 ( .A(n11546), .B(n32), .Z(n33) );
  NANDN U37 ( .A(n18420), .B(n33), .Z(n34) );
  NAND U38 ( .A(n30), .B(n34), .Z(n35) );
  NAND U39 ( .A(n35), .B(n11543), .Z(n36) );
  NAND U40 ( .A(n29), .B(n36), .Z(n37) );
  NAND U41 ( .A(n28), .B(n37), .Z(n38) );
  ANDN U42 ( .B(n38), .A(n11541), .Z(n39) );
  NANDN U43 ( .A(n18426), .B(n39), .Z(n40) );
  NANDN U44 ( .A(n11540), .B(n40), .Z(n41) );
  NAND U45 ( .A(n27), .B(n41), .Z(n42) );
  NAND U46 ( .A(n42), .B(n11537), .Z(n43) );
  NAND U47 ( .A(n26), .B(n43), .Z(n9988) );
  XNOR U48 ( .A(y[3190]), .B(x[3190]), .Z(n44) );
  NOR U49 ( .A(n18469), .B(n11510), .Z(n45) );
  NANDN U50 ( .A(n11511), .B(n11514), .Z(n46) );
  XNOR U51 ( .A(x[3187]), .B(y[3187]), .Z(n47) );
  XNOR U52 ( .A(y[3186]), .B(x[3186]), .Z(n48) );
  ANDN U53 ( .B(n9994), .A(n11515), .Z(n49) );
  NAND U54 ( .A(n9993), .B(n9992), .Z(n50) );
  AND U55 ( .A(n18461), .B(n50), .Z(n51) );
  NANDN U56 ( .A(n11517), .B(n51), .Z(n52) );
  NAND U57 ( .A(n49), .B(n52), .Z(n53) );
  NANDN U58 ( .A(n11518), .B(n53), .Z(n54) );
  NAND U59 ( .A(n48), .B(n54), .Z(n55) );
  NAND U60 ( .A(n55), .B(n11513), .Z(n56) );
  NAND U61 ( .A(n47), .B(n56), .Z(n57) );
  NANDN U62 ( .A(n46), .B(n57), .Z(n58) );
  NAND U63 ( .A(n45), .B(n58), .Z(n59) );
  NANDN U64 ( .A(n11512), .B(n59), .Z(n60) );
  NAND U65 ( .A(n44), .B(n60), .Z(n61) );
  NAND U66 ( .A(n61), .B(n11507), .Z(n9995) );
  XNOR U67 ( .A(y[3214]), .B(x[3214]), .Z(n62) );
  NOR U68 ( .A(n18509), .B(n11480), .Z(n63) );
  NANDN U69 ( .A(n18512), .B(n11482), .Z(n64) );
  XNOR U70 ( .A(x[3211]), .B(y[3211]), .Z(n65) );
  XNOR U71 ( .A(y[3210]), .B(x[3210]), .Z(n66) );
  ANDN U72 ( .B(n10003), .A(n11484), .Z(n67) );
  NAND U73 ( .A(n10002), .B(n10001), .Z(n68) );
  AND U74 ( .A(n11488), .B(n68), .Z(n69) );
  NANDN U75 ( .A(n11485), .B(n69), .Z(n70) );
  NAND U76 ( .A(n67), .B(n70), .Z(n71) );
  NANDN U77 ( .A(n11486), .B(n71), .Z(n72) );
  NAND U78 ( .A(n66), .B(n72), .Z(n73) );
  NAND U79 ( .A(n73), .B(n11481), .Z(n74) );
  NAND U80 ( .A(n65), .B(n74), .Z(n75) );
  NANDN U81 ( .A(n64), .B(n75), .Z(n76) );
  NAND U82 ( .A(n63), .B(n76), .Z(n77) );
  NANDN U83 ( .A(n18513), .B(n77), .Z(n78) );
  NAND U84 ( .A(n62), .B(n78), .Z(n79) );
  NAND U85 ( .A(n79), .B(n11477), .Z(n10004) );
  XNOR U86 ( .A(y[3238]), .B(x[3238]), .Z(n80) );
  NOR U87 ( .A(n11449), .B(n18553), .Z(n81) );
  NANDN U88 ( .A(n11447), .B(n11452), .Z(n82) );
  XNOR U89 ( .A(x[3235]), .B(y[3235]), .Z(n83) );
  XNOR U90 ( .A(y[3234]), .B(x[3234]), .Z(n84) );
  ANDN U91 ( .B(n10012), .A(n11454), .Z(n85) );
  NAND U92 ( .A(n10011), .B(n10010), .Z(n86) );
  AND U93 ( .A(n11456), .B(n86), .Z(n87) );
  NANDN U94 ( .A(n18546), .B(n87), .Z(n88) );
  NAND U95 ( .A(n85), .B(n88), .Z(n89) );
  NANDN U96 ( .A(n18547), .B(n89), .Z(n90) );
  NAND U97 ( .A(n84), .B(n90), .Z(n91) );
  NAND U98 ( .A(n91), .B(n11451), .Z(n92) );
  NAND U99 ( .A(n83), .B(n92), .Z(n93) );
  NANDN U100 ( .A(n82), .B(n93), .Z(n94) );
  NAND U101 ( .A(n81), .B(n94), .Z(n95) );
  NANDN U102 ( .A(n11448), .B(n95), .Z(n96) );
  NAND U103 ( .A(n80), .B(n96), .Z(n97) );
  NAND U104 ( .A(n97), .B(n11445), .Z(n10013) );
  NAND U105 ( .A(n10017), .B(n10016), .Z(n98) );
  AND U106 ( .A(n11425), .B(n98), .Z(n99) );
  NANDN U107 ( .A(n11421), .B(n11426), .Z(n100) );
  XNOR U108 ( .A(y[3255]), .B(x[3255]), .Z(n101) );
  NANDN U109 ( .A(n99), .B(n101), .Z(n102) );
  NANDN U110 ( .A(n100), .B(n102), .Z(n103) );
  NOR U111 ( .A(n18587), .B(n11423), .Z(n104) );
  NAND U112 ( .A(n104), .B(n103), .Z(n105) );
  NANDN U113 ( .A(n11422), .B(n105), .Z(n106) );
  XNOR U114 ( .A(y[3258]), .B(x[3258]), .Z(n107) );
  NAND U115 ( .A(n107), .B(n106), .Z(n108) );
  AND U116 ( .A(n11420), .B(n108), .Z(n109) );
  NAND U117 ( .A(n109), .B(n11416), .Z(n110) );
  ANDN U118 ( .B(n110), .A(n11417), .Z(n111) );
  XNOR U119 ( .A(x[3259]), .B(n109), .Z(n112) );
  AND U120 ( .A(y[3259]), .B(n112), .Z(n113) );
  NANDN U121 ( .A(n113), .B(n111), .Z(n114) );
  NANDN U122 ( .A(n26977), .B(n114), .Z(n115) );
  NAND U123 ( .A(n115), .B(n26978), .Z(n10020) );
  NANDN U124 ( .A(n11394), .B(n11397), .Z(n116) );
  XNOR U125 ( .A(y[3284]), .B(x[3284]), .Z(n117) );
  XNOR U126 ( .A(x[3283]), .B(y[3283]), .Z(n118) );
  XOR U127 ( .A(y[3280]), .B(n11402), .Z(n119) );
  ANDN U128 ( .B(n10029), .A(n18624), .Z(n120) );
  NAND U129 ( .A(n119), .B(n120), .Z(n121) );
  NAND U130 ( .A(y[3280]), .B(n11402), .Z(n122) );
  AND U131 ( .A(n121), .B(n122), .Z(n123) );
  XNOR U132 ( .A(x[3281]), .B(y[3281]), .Z(n124) );
  NANDN U133 ( .A(n123), .B(n124), .Z(n125) );
  NAND U134 ( .A(n125), .B(n11398), .Z(n126) );
  XNOR U135 ( .A(x[3282]), .B(n126), .Z(n127) );
  NANDN U136 ( .A(y[3282]), .B(n127), .Z(n128) );
  NANDN U137 ( .A(n126), .B(x[3282]), .Z(n129) );
  AND U138 ( .A(n128), .B(n129), .Z(n130) );
  NAND U139 ( .A(n118), .B(n130), .Z(n131) );
  NAND U140 ( .A(n131), .B(n11396), .Z(n132) );
  NAND U141 ( .A(n117), .B(n132), .Z(n133) );
  NANDN U142 ( .A(n116), .B(n133), .Z(n10030) );
  NANDN U143 ( .A(n11367), .B(n11368), .Z(n134) );
  XNOR U144 ( .A(y[3302]), .B(x[3302]), .Z(n135) );
  XNOR U145 ( .A(x[3301]), .B(y[3301]), .Z(n136) );
  NAND U146 ( .A(y[3300]), .B(n11372), .Z(n137) );
  XOR U147 ( .A(n11372), .B(y[3300]), .Z(n138) );
  XNOR U148 ( .A(x[3299]), .B(y[3299]), .Z(n139) );
  XNOR U149 ( .A(x[3298]), .B(y[3298]), .Z(n140) );
  NANDN U150 ( .A(n18652), .B(n10032), .Z(n141) );
  NAND U151 ( .A(n140), .B(n141), .Z(n142) );
  NANDN U152 ( .A(y[3298]), .B(x[3298]), .Z(n143) );
  AND U153 ( .A(n142), .B(n143), .Z(n144) );
  NAND U154 ( .A(n139), .B(n144), .Z(n145) );
  NAND U155 ( .A(n145), .B(n11373), .Z(n146) );
  NAND U156 ( .A(n138), .B(n146), .Z(n147) );
  NAND U157 ( .A(n137), .B(n147), .Z(n148) );
  NAND U158 ( .A(n136), .B(n148), .Z(n149) );
  NAND U159 ( .A(n149), .B(n11369), .Z(n150) );
  NAND U160 ( .A(n135), .B(n150), .Z(n151) );
  NANDN U161 ( .A(n134), .B(n151), .Z(n10033) );
  ANDN U162 ( .B(n11331), .A(n27122), .Z(n152) );
  NAND U163 ( .A(n10059), .B(n10058), .Z(n153) );
  AND U164 ( .A(n152), .B(n153), .Z(n154) );
  ANDN U165 ( .B(n10063), .A(n154), .Z(n155) );
  NAND U166 ( .A(n155), .B(n27124), .Z(n156) );
  ANDN U167 ( .B(n156), .A(n27126), .Z(n157) );
  NANDN U168 ( .A(n157), .B(n27128), .Z(n158) );
  ANDN U169 ( .B(n158), .A(n11328), .Z(n159) );
  XNOR U170 ( .A(y[3337]), .B(x[3337]), .Z(n160) );
  NAND U171 ( .A(n160), .B(n159), .Z(n161) );
  AND U172 ( .A(n11325), .B(n161), .Z(n162) );
  OR U173 ( .A(n11324), .B(n162), .Z(n163) );
  AND U174 ( .A(n27138), .B(n163), .Z(n164) );
  ANDN U175 ( .B(n18724), .A(n11323), .Z(n165) );
  NANDN U176 ( .A(n11326), .B(n164), .Z(n166) );
  AND U177 ( .A(n165), .B(n166), .Z(n167) );
  NOR U178 ( .A(n167), .B(n18727), .Z(n168) );
  NANDN U179 ( .A(n27137), .B(n168), .Z(n169) );
  ANDN U180 ( .B(n169), .A(n11321), .Z(n10066) );
  NOR U181 ( .A(n18842), .B(n11249), .Z(n170) );
  NAND U182 ( .A(n10100), .B(n10099), .Z(n171) );
  AND U183 ( .A(n11257), .B(n171), .Z(n172) );
  NANDN U184 ( .A(n11255), .B(n11258), .Z(n173) );
  XNOR U185 ( .A(y[3399]), .B(x[3399]), .Z(n174) );
  NANDN U186 ( .A(n172), .B(n174), .Z(n175) );
  NANDN U187 ( .A(n173), .B(n175), .Z(n176) );
  NOR U188 ( .A(n18834), .B(n11254), .Z(n177) );
  NAND U189 ( .A(n177), .B(n176), .Z(n178) );
  NANDN U190 ( .A(n11256), .B(n178), .Z(n179) );
  XNOR U191 ( .A(y[3402]), .B(x[3402]), .Z(n180) );
  NAND U192 ( .A(n180), .B(n179), .Z(n181) );
  NAND U193 ( .A(n181), .B(n18839), .Z(n182) );
  NANDN U194 ( .A(n11251), .B(n18840), .Z(n183) );
  XNOR U195 ( .A(x[3403]), .B(y[3403]), .Z(n184) );
  NAND U196 ( .A(n184), .B(n182), .Z(n185) );
  NANDN U197 ( .A(n183), .B(n185), .Z(n186) );
  NAND U198 ( .A(n170), .B(n186), .Z(n10101) );
  XOR U199 ( .A(x[3433]), .B(n11213), .Z(n187) );
  NANDN U200 ( .A(n10127), .B(n187), .Z(n188) );
  NAND U201 ( .A(x[3433]), .B(n11213), .Z(n189) );
  AND U202 ( .A(n188), .B(n189), .Z(n190) );
  XNOR U203 ( .A(x[3434]), .B(y[3434]), .Z(n191) );
  AND U204 ( .A(n190), .B(n191), .Z(n192) );
  NOR U205 ( .A(n192), .B(n18901), .Z(n193) );
  NAND U206 ( .A(n193), .B(n18898), .Z(n194) );
  ANDN U207 ( .B(n194), .A(n11212), .Z(n195) );
  NANDN U208 ( .A(n11209), .B(n18902), .Z(n196) );
  XNOR U209 ( .A(x[3436]), .B(y[3436]), .Z(n197) );
  NAND U210 ( .A(n197), .B(n195), .Z(n198) );
  NANDN U211 ( .A(n196), .B(n198), .Z(n199) );
  NOR U212 ( .A(n18904), .B(n18909), .Z(n200) );
  NAND U213 ( .A(n200), .B(n199), .Z(n201) );
  NANDN U214 ( .A(n11210), .B(n201), .Z(n202) );
  XNOR U215 ( .A(x[3439]), .B(y[3439]), .Z(n203) );
  NAND U216 ( .A(n203), .B(n202), .Z(n204) );
  NAND U217 ( .A(n204), .B(n11207), .Z(n10128) );
  XNOR U218 ( .A(x[3463]), .B(y[3463]), .Z(n205) );
  NOR U219 ( .A(n18954), .B(n11186), .Z(n206) );
  NANDN U220 ( .A(n11187), .B(n11190), .Z(n207) );
  XNOR U221 ( .A(y[3460]), .B(x[3460]), .Z(n208) );
  XNOR U222 ( .A(x[3459]), .B(y[3459]), .Z(n209) );
  ANDN U223 ( .B(n10135), .A(n18951), .Z(n210) );
  NAND U224 ( .A(n10134), .B(n10133), .Z(n211) );
  AND U225 ( .A(n18944), .B(n211), .Z(n212) );
  NANDN U226 ( .A(n11191), .B(n212), .Z(n213) );
  NAND U227 ( .A(n210), .B(n213), .Z(n214) );
  NANDN U228 ( .A(n11192), .B(n214), .Z(n215) );
  NAND U229 ( .A(n209), .B(n215), .Z(n216) );
  NAND U230 ( .A(n216), .B(n11189), .Z(n217) );
  NAND U231 ( .A(n208), .B(n217), .Z(n218) );
  NANDN U232 ( .A(n207), .B(n218), .Z(n219) );
  NAND U233 ( .A(n206), .B(n219), .Z(n220) );
  NANDN U234 ( .A(n11188), .B(n220), .Z(n221) );
  NAND U235 ( .A(n205), .B(n221), .Z(n222) );
  NAND U236 ( .A(n222), .B(n18959), .Z(n10136) );
  NANDN U237 ( .A(n12547), .B(n22476), .Z(n223) );
  AND U238 ( .A(n6789), .B(n223), .Z(n224) );
  NANDN U239 ( .A(n12548), .B(n6782), .Z(n225) );
  NAND U240 ( .A(n225), .B(n22465), .Z(n226) );
  NAND U241 ( .A(n226), .B(n22466), .Z(n227) );
  NAND U242 ( .A(n227), .B(n22468), .Z(n228) );
  NAND U243 ( .A(n228), .B(n22470), .Z(n229) );
  ANDN U244 ( .B(n229), .A(n12546), .Z(n230) );
  NANDN U245 ( .A(n230), .B(n22475), .Z(n231) );
  NANDN U246 ( .A(n224), .B(n231), .Z(n232) );
  NANDN U247 ( .A(n22479), .B(n232), .Z(n233) );
  NAND U248 ( .A(n233), .B(n22480), .Z(n234) );
  AND U249 ( .A(n22482), .B(n234), .Z(n235) );
  NANDN U250 ( .A(n12543), .B(n235), .Z(n236) );
  NAND U251 ( .A(n236), .B(n22484), .Z(n237) );
  NANDN U252 ( .A(n237), .B(x[1319]), .Z(n238) );
  XNOR U253 ( .A(n237), .B(x[1319]), .Z(n239) );
  NAND U254 ( .A(n239), .B(n12542), .Z(n240) );
  NAND U255 ( .A(n238), .B(n240), .Z(n6791) );
  AND U256 ( .A(n16683), .B(n8835), .Z(n241) );
  NAND U257 ( .A(n241), .B(n24803), .Z(n242) );
  AND U258 ( .A(n24806), .B(n242), .Z(n243) );
  NANDN U259 ( .A(n12067), .B(n243), .Z(n244) );
  NAND U260 ( .A(n244), .B(n24807), .Z(n245) );
  ANDN U261 ( .B(n245), .A(n24810), .Z(n246) );
  ANDN U262 ( .B(n24813), .A(n16700), .Z(n247) );
  NANDN U263 ( .A(n246), .B(n24811), .Z(n248) );
  AND U264 ( .A(n247), .B(n248), .Z(n249) );
  NANDN U265 ( .A(n249), .B(n24815), .Z(n250) );
  ANDN U266 ( .B(n250), .A(n16703), .Z(n251) );
  OR U267 ( .A(n16699), .B(n8837), .Z(n252) );
  NAND U268 ( .A(n252), .B(n251), .Z(n253) );
  AND U269 ( .A(n24819), .B(n253), .Z(n254) );
  OR U270 ( .A(n24822), .B(n254), .Z(n255) );
  ANDN U271 ( .B(n255), .A(n24824), .Z(n256) );
  NANDN U272 ( .A(n256), .B(n24826), .Z(n257) );
  NAND U273 ( .A(n257), .B(n24827), .Z(n258) );
  NAND U274 ( .A(n258), .B(n24829), .Z(n8847) );
  NAND U275 ( .A(n25369), .B(n9228), .Z(n259) );
  NANDN U276 ( .A(n25372), .B(n259), .Z(n260) );
  ANDN U277 ( .B(n260), .A(n25373), .Z(n261) );
  NOR U278 ( .A(n261), .B(n11949), .Z(n262) );
  NAND U279 ( .A(n262), .B(n25375), .Z(n263) );
  NAND U280 ( .A(n263), .B(n25377), .Z(n264) );
  ANDN U281 ( .B(n20244), .A(n11952), .Z(n265) );
  NAND U282 ( .A(n265), .B(n264), .Z(n266) );
  NAND U283 ( .A(n266), .B(n25381), .Z(n267) );
  NAND U284 ( .A(n267), .B(n25383), .Z(n268) );
  NAND U285 ( .A(n268), .B(n25385), .Z(n269) );
  AND U286 ( .A(n25387), .B(n269), .Z(n270) );
  OR U287 ( .A(n25389), .B(n270), .Z(n271) );
  NAND U288 ( .A(n271), .B(n25391), .Z(n272) );
  NANDN U289 ( .A(n25394), .B(n272), .Z(n273) );
  NAND U290 ( .A(n273), .B(n25395), .Z(n274) );
  AND U291 ( .A(n25397), .B(n274), .Z(n275) );
  NANDN U292 ( .A(n17247), .B(n275), .Z(n276) );
  NAND U293 ( .A(n276), .B(n25399), .Z(n9231) );
  NAND U294 ( .A(n15523), .B(n15524), .Z(n277) );
  NAND U295 ( .A(n277), .B(n23466), .Z(n278) );
  NAND U296 ( .A(n278), .B(n23468), .Z(n279) );
  NAND U297 ( .A(n279), .B(n15525), .Z(n280) );
  NANDN U298 ( .A(n23472), .B(n280), .Z(n281) );
  AND U299 ( .A(n15526), .B(n281), .Z(n282) );
  NANDN U300 ( .A(n23473), .B(n282), .Z(n283) );
  NAND U301 ( .A(n283), .B(n23476), .Z(n284) );
  AND U302 ( .A(n15527), .B(n284), .Z(n285) );
  NANDN U303 ( .A(n285), .B(n23480), .Z(n286) );
  NAND U304 ( .A(n286), .B(n23482), .Z(n287) );
  NANDN U305 ( .A(n23485), .B(n287), .Z(n288) );
  NAND U306 ( .A(n288), .B(n23486), .Z(n289) );
  NAND U307 ( .A(n289), .B(n23489), .Z(n290) );
  ANDN U308 ( .B(n290), .A(n23491), .Z(n291) );
  OR U309 ( .A(n23493), .B(n291), .Z(n292) );
  NANDN U310 ( .A(n23495), .B(n292), .Z(n293) );
  NAND U311 ( .A(n293), .B(n23496), .Z(n294) );
  NANDN U312 ( .A(n23499), .B(n294), .Z(n15528) );
  ANDN U313 ( .B(n26394), .A(n18084), .Z(n9838) );
  NANDN U314 ( .A(n9920), .B(n9919), .Z(n295) );
  ANDN U315 ( .B(n295), .A(n11623), .Z(n296) );
  XNOR U316 ( .A(y[3099]), .B(x[3099]), .Z(n297) );
  NAND U317 ( .A(n297), .B(n296), .Z(n298) );
  ANDN U318 ( .B(n11621), .A(n11617), .Z(n299) );
  NAND U319 ( .A(n299), .B(n298), .Z(n300) );
  NANDN U320 ( .A(n11619), .B(n300), .Z(n301) );
  ANDN U321 ( .B(n11616), .A(n11614), .Z(n302) );
  XNOR U322 ( .A(y[3101]), .B(x[3101]), .Z(n303) );
  NANDN U323 ( .A(n301), .B(n303), .Z(n304) );
  AND U324 ( .A(n302), .B(n304), .Z(n305) );
  NOR U325 ( .A(n18333), .B(n11612), .Z(n306) );
  NANDN U326 ( .A(n305), .B(n306), .Z(n307) );
  ANDN U327 ( .B(n307), .A(n11615), .Z(n308) );
  XNOR U328 ( .A(y[3104]), .B(x[3104]), .Z(n309) );
  NANDN U329 ( .A(n308), .B(n309), .Z(n310) );
  AND U330 ( .A(n11610), .B(n310), .Z(n311) );
  XNOR U331 ( .A(x[3105]), .B(y[3105]), .Z(n312) );
  NANDN U332 ( .A(n311), .B(n312), .Z(n9921) );
  NAND U333 ( .A(n9952), .B(n26718), .Z(n313) );
  NANDN U334 ( .A(n26720), .B(n313), .Z(n314) );
  NAND U335 ( .A(n314), .B(n26722), .Z(n315) );
  NANDN U336 ( .A(n26724), .B(n315), .Z(n316) );
  NANDN U337 ( .A(n11566), .B(n316), .Z(n317) );
  ANDN U338 ( .B(n317), .A(n11565), .Z(n318) );
  XNOR U339 ( .A(y[3138]), .B(x[3138]), .Z(n319) );
  OR U340 ( .A(n11567), .B(n318), .Z(n320) );
  AND U341 ( .A(n319), .B(n320), .Z(n321) );
  XNOR U342 ( .A(x[3139]), .B(y[3139]), .Z(n322) );
  NANDN U343 ( .A(n321), .B(n18378), .Z(n323) );
  AND U344 ( .A(n322), .B(n323), .Z(n324) );
  NOR U345 ( .A(n324), .B(n11563), .Z(n325) );
  NAND U346 ( .A(n325), .B(n18379), .Z(n326) );
  NANDN U347 ( .A(n18381), .B(n326), .Z(n327) );
  NANDN U348 ( .A(n327), .B(x[3141]), .Z(n328) );
  XNOR U349 ( .A(n327), .B(x[3141]), .Z(n329) );
  NAND U350 ( .A(n329), .B(n11561), .Z(n330) );
  NAND U351 ( .A(n328), .B(n330), .Z(n9959) );
  NANDN U352 ( .A(n11535), .B(n11538), .Z(n331) );
  ANDN U353 ( .B(n9989), .A(n11534), .Z(n332) );
  NANDN U354 ( .A(n331), .B(n9988), .Z(n333) );
  AND U355 ( .A(n332), .B(n333), .Z(n334) );
  XNOR U356 ( .A(y[3169]), .B(x[3169]), .Z(n335) );
  OR U357 ( .A(n11536), .B(n334), .Z(n336) );
  NAND U358 ( .A(n335), .B(n336), .Z(n337) );
  XNOR U359 ( .A(x[3170]), .B(y[3170]), .Z(n338) );
  NAND U360 ( .A(n337), .B(n18435), .Z(n339) );
  NAND U361 ( .A(n338), .B(n339), .Z(n340) );
  ANDN U362 ( .B(n18436), .A(n11532), .Z(n341) );
  NAND U363 ( .A(n341), .B(n340), .Z(n342) );
  ANDN U364 ( .B(n342), .A(n18438), .Z(n343) );
  NANDN U365 ( .A(n11530), .B(n343), .Z(n344) );
  ANDN U366 ( .B(n26801), .A(n11531), .Z(n345) );
  NAND U367 ( .A(n345), .B(n344), .Z(n346) );
  NANDN U368 ( .A(n11529), .B(n346), .Z(n347) );
  NANDN U369 ( .A(n347), .B(n18443), .Z(n348) );
  ANDN U370 ( .B(n348), .A(n26800), .Z(n9990) );
  XNOR U371 ( .A(y[3198]), .B(x[3198]), .Z(n349) );
  NOR U372 ( .A(n11501), .B(n18485), .Z(n350) );
  NANDN U373 ( .A(n11499), .B(n11504), .Z(n351) );
  XNOR U374 ( .A(x[3195]), .B(y[3195]), .Z(n352) );
  XNOR U375 ( .A(y[3194]), .B(x[3194]), .Z(n353) );
  ANDN U376 ( .B(n9997), .A(n11506), .Z(n354) );
  NAND U377 ( .A(n9996), .B(n9995), .Z(n355) );
  AND U378 ( .A(n11508), .B(n355), .Z(n356) );
  NANDN U379 ( .A(n18478), .B(n356), .Z(n357) );
  NAND U380 ( .A(n354), .B(n357), .Z(n358) );
  NANDN U381 ( .A(n18479), .B(n358), .Z(n359) );
  NAND U382 ( .A(n353), .B(n359), .Z(n360) );
  NAND U383 ( .A(n360), .B(n11503), .Z(n361) );
  NAND U384 ( .A(n352), .B(n361), .Z(n362) );
  NANDN U385 ( .A(n351), .B(n362), .Z(n363) );
  NAND U386 ( .A(n350), .B(n363), .Z(n364) );
  NANDN U387 ( .A(n11500), .B(n364), .Z(n365) );
  NAND U388 ( .A(n349), .B(n365), .Z(n366) );
  NAND U389 ( .A(n366), .B(n11497), .Z(n9998) );
  XNOR U390 ( .A(y[3222]), .B(x[3222]), .Z(n367) );
  NOR U391 ( .A(n18523), .B(n11468), .Z(n368) );
  NANDN U392 ( .A(n11469), .B(n11472), .Z(n369) );
  XNOR U393 ( .A(x[3219]), .B(y[3219]), .Z(n370) );
  XNOR U394 ( .A(y[3218]), .B(x[3218]), .Z(n371) );
  ANDN U395 ( .B(n10006), .A(n18519), .Z(n372) );
  NAND U396 ( .A(n10005), .B(n10004), .Z(n373) );
  AND U397 ( .A(n11478), .B(n373), .Z(n374) );
  NANDN U398 ( .A(n11473), .B(n374), .Z(n375) );
  NAND U399 ( .A(n372), .B(n375), .Z(n376) );
  NANDN U400 ( .A(n11474), .B(n376), .Z(n377) );
  NAND U401 ( .A(n371), .B(n377), .Z(n378) );
  NAND U402 ( .A(n378), .B(n11471), .Z(n379) );
  NAND U403 ( .A(n370), .B(n379), .Z(n380) );
  NANDN U404 ( .A(n369), .B(n380), .Z(n381) );
  NAND U405 ( .A(n368), .B(n381), .Z(n382) );
  NANDN U406 ( .A(n11470), .B(n382), .Z(n383) );
  NAND U407 ( .A(n367), .B(n383), .Z(n384) );
  NAND U408 ( .A(n384), .B(n18528), .Z(n10007) );
  ANDN U409 ( .B(n11446), .A(n11443), .Z(n385) );
  NAND U410 ( .A(n10014), .B(n10013), .Z(n386) );
  AND U411 ( .A(n385), .B(n386), .Z(n387) );
  NOR U412 ( .A(n11442), .B(n18557), .Z(n388) );
  NANDN U413 ( .A(n387), .B(n388), .Z(n389) );
  ANDN U414 ( .B(n389), .A(n11444), .Z(n390) );
  XNOR U415 ( .A(y[3242]), .B(x[3242]), .Z(n391) );
  NANDN U416 ( .A(n390), .B(n391), .Z(n392) );
  AND U417 ( .A(n18562), .B(n392), .Z(n393) );
  ANDN U418 ( .B(n18563), .A(n11439), .Z(n394) );
  XNOR U419 ( .A(y[3243]), .B(x[3243]), .Z(n395) );
  NANDN U420 ( .A(n393), .B(n395), .Z(n396) );
  AND U421 ( .A(n394), .B(n396), .Z(n397) );
  NOR U422 ( .A(n11437), .B(n18565), .Z(n398) );
  NANDN U423 ( .A(n397), .B(n398), .Z(n399) );
  ANDN U424 ( .B(n399), .A(n11440), .Z(n400) );
  XNOR U425 ( .A(y[3246]), .B(x[3246]), .Z(n401) );
  NANDN U426 ( .A(n400), .B(n401), .Z(n10015) );
  ANDN U427 ( .B(n10020), .A(n11415), .Z(n402) );
  XNOR U428 ( .A(y[3263]), .B(x[3263]), .Z(n403) );
  AND U429 ( .A(n402), .B(n403), .Z(n404) );
  NOR U430 ( .A(n404), .B(n18596), .Z(n405) );
  NAND U431 ( .A(n405), .B(n18595), .Z(n406) );
  AND U432 ( .A(n26984), .B(n406), .Z(n407) );
  NANDN U433 ( .A(n407), .B(n26987), .Z(n408) );
  AND U434 ( .A(n26988), .B(n408), .Z(n409) );
  NANDN U435 ( .A(n409), .B(n26991), .Z(n410) );
  NANDN U436 ( .A(n18603), .B(n410), .Z(n411) );
  NAND U437 ( .A(n411), .B(n20231), .Z(n412) );
  ANDN U438 ( .B(n18606), .A(n18602), .Z(n413) );
  NAND U439 ( .A(n413), .B(n412), .Z(n414) );
  NANDN U440 ( .A(n20230), .B(n414), .Z(n415) );
  XNOR U441 ( .A(y[3271]), .B(x[3271]), .Z(n416) );
  NANDN U442 ( .A(n415), .B(n416), .Z(n417) );
  ANDN U443 ( .B(n11413), .A(n18612), .Z(n418) );
  NAND U444 ( .A(n418), .B(n417), .Z(n419) );
  NANDN U445 ( .A(n18609), .B(n419), .Z(n10028) );
  NANDN U446 ( .A(n11384), .B(n11388), .Z(n420) );
  XNOR U447 ( .A(y[3290]), .B(x[3290]), .Z(n421) );
  XNOR U448 ( .A(x[3289]), .B(y[3289]), .Z(n422) );
  XOR U449 ( .A(y[3286]), .B(n11393), .Z(n423) );
  ANDN U450 ( .B(n10030), .A(n18634), .Z(n424) );
  NAND U451 ( .A(n423), .B(n424), .Z(n425) );
  NAND U452 ( .A(y[3286]), .B(n11393), .Z(n426) );
  AND U453 ( .A(n425), .B(n426), .Z(n427) );
  XNOR U454 ( .A(x[3287]), .B(y[3287]), .Z(n428) );
  NANDN U455 ( .A(n427), .B(n428), .Z(n429) );
  NAND U456 ( .A(n429), .B(n18639), .Z(n430) );
  XNOR U457 ( .A(x[3288]), .B(n430), .Z(n431) );
  NANDN U458 ( .A(y[3288]), .B(n431), .Z(n432) );
  NANDN U459 ( .A(n430), .B(x[3288]), .Z(n433) );
  AND U460 ( .A(n432), .B(n433), .Z(n434) );
  NAND U461 ( .A(n422), .B(n434), .Z(n435) );
  NAND U462 ( .A(n435), .B(n11387), .Z(n436) );
  NAND U463 ( .A(n421), .B(n436), .Z(n437) );
  NANDN U464 ( .A(n420), .B(n437), .Z(n10031) );
  NANDN U465 ( .A(n18662), .B(n10033), .Z(n438) );
  XNOR U466 ( .A(x[3304]), .B(y[3304]), .Z(n439) );
  NAND U467 ( .A(n439), .B(n438), .Z(n440) );
  NANDN U468 ( .A(y[3304]), .B(x[3304]), .Z(n441) );
  AND U469 ( .A(n440), .B(n441), .Z(n442) );
  XNOR U470 ( .A(x[3305]), .B(y[3305]), .Z(n443) );
  NAND U471 ( .A(n443), .B(n442), .Z(n444) );
  NAND U472 ( .A(n444), .B(n11362), .Z(n445) );
  NAND U473 ( .A(y[3306]), .B(n11361), .Z(n446) );
  XOR U474 ( .A(n11361), .B(y[3306]), .Z(n447) );
  NAND U475 ( .A(n447), .B(n445), .Z(n448) );
  NAND U476 ( .A(n446), .B(n448), .Z(n449) );
  XNOR U477 ( .A(x[3307]), .B(y[3307]), .Z(n450) );
  NAND U478 ( .A(n450), .B(n449), .Z(n451) );
  NAND U479 ( .A(n451), .B(n18669), .Z(n452) );
  NANDN U480 ( .A(n11358), .B(n18670), .Z(n453) );
  XNOR U481 ( .A(y[3308]), .B(x[3308]), .Z(n454) );
  NAND U482 ( .A(n454), .B(n452), .Z(n455) );
  NANDN U483 ( .A(n453), .B(n455), .Z(n10034) );
  NANDN U484 ( .A(n11307), .B(n11312), .Z(n456) );
  XNOR U485 ( .A(x[3350]), .B(y[3350]), .Z(n457) );
  NAND U486 ( .A(n457), .B(n10069), .Z(n458) );
  NANDN U487 ( .A(n456), .B(n458), .Z(n459) );
  NOR U488 ( .A(n11309), .B(n18746), .Z(n460) );
  NAND U489 ( .A(n460), .B(n459), .Z(n461) );
  NANDN U490 ( .A(n11308), .B(n461), .Z(n462) );
  XNOR U491 ( .A(x[3353]), .B(y[3353]), .Z(n463) );
  NAND U492 ( .A(n463), .B(n462), .Z(n464) );
  NAND U493 ( .A(n464), .B(n11306), .Z(n465) );
  NAND U494 ( .A(n27172), .B(n11305), .Z(n466) );
  XNOR U495 ( .A(y[3354]), .B(x[3354]), .Z(n467) );
  NAND U496 ( .A(n467), .B(n465), .Z(n468) );
  NANDN U497 ( .A(n466), .B(n468), .Z(n469) );
  ANDN U498 ( .B(n18754), .A(n18750), .Z(n470) );
  NAND U499 ( .A(n470), .B(n469), .Z(n471) );
  NAND U500 ( .A(n471), .B(n27178), .Z(n472) );
  OR U501 ( .A(n27170), .B(n472), .Z(n473) );
  AND U502 ( .A(n18760), .B(n473), .Z(n10070) );
  NANDN U503 ( .A(n18823), .B(n11268), .Z(n474) );
  ANDN U504 ( .B(n10098), .A(n27244), .Z(n475) );
  XNOR U505 ( .A(x[3391]), .B(y[3391]), .Z(n476) );
  AND U506 ( .A(n475), .B(n476), .Z(n477) );
  NOR U507 ( .A(n18820), .B(n11266), .Z(n478) );
  OR U508 ( .A(n474), .B(n477), .Z(n479) );
  AND U509 ( .A(n478), .B(n479), .Z(n480) );
  XNOR U510 ( .A(x[3394]), .B(y[3394]), .Z(n481) );
  OR U511 ( .A(n18824), .B(n480), .Z(n482) );
  NAND U512 ( .A(n481), .B(n482), .Z(n483) );
  XNOR U513 ( .A(y[3395]), .B(x[3395]), .Z(n484) );
  NAND U514 ( .A(n483), .B(n11264), .Z(n485) );
  NAND U515 ( .A(n484), .B(n485), .Z(n486) );
  ANDN U516 ( .B(n11263), .A(n11259), .Z(n487) );
  NAND U517 ( .A(n487), .B(n486), .Z(n488) );
  ANDN U518 ( .B(n488), .A(n11261), .Z(n489) );
  NANDN U519 ( .A(n18830), .B(n489), .Z(n490) );
  NANDN U520 ( .A(n11260), .B(n490), .Z(n10099) );
  AND U521 ( .A(n10105), .B(n10104), .Z(n491) );
  XNOR U522 ( .A(x[3414]), .B(y[3414]), .Z(n492) );
  AND U523 ( .A(n491), .B(n492), .Z(n493) );
  NOR U524 ( .A(n493), .B(n11237), .Z(n494) );
  NAND U525 ( .A(n494), .B(n11240), .Z(n495) );
  NANDN U526 ( .A(n18862), .B(n495), .Z(n496) );
  NANDN U527 ( .A(n496), .B(y[3416]), .Z(n497) );
  XNOR U528 ( .A(n496), .B(y[3416]), .Z(n498) );
  NAND U529 ( .A(n498), .B(n11236), .Z(n499) );
  NAND U530 ( .A(n497), .B(n499), .Z(n500) );
  XNOR U531 ( .A(x[3417]), .B(y[3417]), .Z(n501) );
  NAND U532 ( .A(n501), .B(n500), .Z(n502) );
  NAND U533 ( .A(n502), .B(n18867), .Z(n503) );
  XNOR U534 ( .A(y[3418]), .B(x[3418]), .Z(n504) );
  AND U535 ( .A(n503), .B(n504), .Z(n505) );
  NOR U536 ( .A(n505), .B(n11233), .Z(n506) );
  NAND U537 ( .A(n506), .B(n18868), .Z(n507) );
  NANDN U538 ( .A(n18870), .B(n507), .Z(n10106) );
  XNOR U539 ( .A(x[3455]), .B(y[3455]), .Z(n508) );
  NOR U540 ( .A(n18936), .B(n11194), .Z(n509) );
  NANDN U541 ( .A(n18939), .B(n11196), .Z(n510) );
  XNOR U542 ( .A(y[3452]), .B(x[3452]), .Z(n511) );
  XNOR U543 ( .A(x[3451]), .B(y[3451]), .Z(n512) );
  ANDN U544 ( .B(n18929), .A(n18932), .Z(n513) );
  NAND U545 ( .A(n10132), .B(n10131), .Z(n514) );
  AND U546 ( .A(n11200), .B(n514), .Z(n515) );
  NANDN U547 ( .A(n11197), .B(n515), .Z(n516) );
  NAND U548 ( .A(n513), .B(n516), .Z(n517) );
  NANDN U549 ( .A(n11198), .B(n517), .Z(n518) );
  NAND U550 ( .A(n512), .B(n518), .Z(n519) );
  NAND U551 ( .A(n519), .B(n11195), .Z(n520) );
  NAND U552 ( .A(n511), .B(n520), .Z(n521) );
  NANDN U553 ( .A(n510), .B(n521), .Z(n522) );
  NAND U554 ( .A(n509), .B(n522), .Z(n523) );
  NANDN U555 ( .A(n18940), .B(n523), .Z(n524) );
  NAND U556 ( .A(n508), .B(n524), .Z(n525) );
  NAND U557 ( .A(n525), .B(n18943), .Z(n10133) );
  NAND U558 ( .A(n10139), .B(n10138), .Z(n526) );
  ANDN U559 ( .B(n526), .A(n18979), .Z(n527) );
  NANDN U560 ( .A(n11173), .B(n11177), .Z(n528) );
  XNOR U561 ( .A(y[3473]), .B(x[3473]), .Z(n529) );
  NAND U562 ( .A(n529), .B(n527), .Z(n530) );
  NANDN U563 ( .A(n528), .B(n530), .Z(n531) );
  ANDN U564 ( .B(n11176), .A(n11172), .Z(n532) );
  NAND U565 ( .A(n532), .B(n531), .Z(n533) );
  ANDN U566 ( .B(n533), .A(n11174), .Z(n534) );
  NANDN U567 ( .A(n534), .B(n18985), .Z(n535) );
  XOR U568 ( .A(n534), .B(y[3476]), .Z(n536) );
  NAND U569 ( .A(n536), .B(x[3476]), .Z(n537) );
  AND U570 ( .A(n535), .B(n537), .Z(n538) );
  ANDN U571 ( .B(n18990), .A(n18987), .Z(n539) );
  NANDN U572 ( .A(n538), .B(n27427), .Z(n540) );
  AND U573 ( .A(n539), .B(n540), .Z(n541) );
  NOR U574 ( .A(n541), .B(n18997), .Z(n542) );
  NANDN U575 ( .A(n27426), .B(n542), .Z(n543) );
  NANDN U576 ( .A(n18992), .B(n543), .Z(n10140) );
  OR U577 ( .A(n10924), .B(n19413), .Z(n10213) );
  NANDN U578 ( .A(n12957), .B(n4228), .Z(n544) );
  NANDN U579 ( .A(n12959), .B(n544), .Z(n545) );
  ANDN U580 ( .B(n545), .A(n12962), .Z(n546) );
  OR U581 ( .A(x[68]), .B(n546), .Z(n547) );
  XOR U582 ( .A(x[68]), .B(n546), .Z(n548) );
  NAND U583 ( .A(n548), .B(y[68]), .Z(n549) );
  NAND U584 ( .A(n547), .B(n549), .Z(n550) );
  AND U585 ( .A(n12964), .B(n550), .Z(n551) );
  OR U586 ( .A(n12970), .B(n551), .Z(n552) );
  NANDN U587 ( .A(n12972), .B(n552), .Z(n553) );
  ANDN U588 ( .B(n553), .A(n12973), .Z(n554) );
  OR U589 ( .A(n12976), .B(n554), .Z(n555) );
  NANDN U590 ( .A(n12978), .B(n555), .Z(n556) );
  ANDN U591 ( .B(n556), .A(n12980), .Z(n557) );
  OR U592 ( .A(n12982), .B(n557), .Z(n558) );
  NANDN U593 ( .A(n12984), .B(n558), .Z(n559) );
  ANDN U594 ( .B(n559), .A(n12985), .Z(n560) );
  OR U595 ( .A(n12988), .B(n560), .Z(n561) );
  ANDN U596 ( .B(n561), .A(n12990), .Z(n4233) );
  XNOR U597 ( .A(x[1320]), .B(y[1320]), .Z(n562) );
  NAND U598 ( .A(n562), .B(n6791), .Z(n563) );
  AND U599 ( .A(n12539), .B(n563), .Z(n564) );
  OR U600 ( .A(y[1321]), .B(n564), .Z(n565) );
  XOR U601 ( .A(n564), .B(y[1321]), .Z(n566) );
  NAND U602 ( .A(n566), .B(x[1321]), .Z(n567) );
  NAND U603 ( .A(n565), .B(n567), .Z(n568) );
  ANDN U604 ( .B(n568), .A(n12537), .Z(n569) );
  OR U605 ( .A(n22494), .B(n569), .Z(n570) );
  AND U606 ( .A(n22496), .B(n570), .Z(n571) );
  OR U607 ( .A(n22499), .B(n571), .Z(n572) );
  NANDN U608 ( .A(n14767), .B(n572), .Z(n573) );
  NAND U609 ( .A(n573), .B(n22502), .Z(n574) );
  OR U610 ( .A(n22504), .B(n14768), .Z(n575) );
  NAND U611 ( .A(n575), .B(n6796), .Z(n576) );
  AND U612 ( .A(n574), .B(n576), .Z(n577) );
  NOR U613 ( .A(n12535), .B(n12534), .Z(n578) );
  OR U614 ( .A(n14773), .B(n577), .Z(n579) );
  NAND U615 ( .A(n578), .B(n579), .Z(n6798) );
  XNOR U616 ( .A(y[1837]), .B(x[1837]), .Z(n580) );
  NAND U617 ( .A(n580), .B(n7934), .Z(n581) );
  AND U618 ( .A(n23625), .B(n12270), .Z(n582) );
  NAND U619 ( .A(n582), .B(n581), .Z(n583) );
  NANDN U620 ( .A(n12268), .B(n583), .Z(n584) );
  NAND U621 ( .A(n584), .B(n23630), .Z(n585) );
  AND U622 ( .A(n23633), .B(n585), .Z(n586) );
  NAND U623 ( .A(n586), .B(n23627), .Z(n587) );
  AND U624 ( .A(n23637), .B(n587), .Z(n588) );
  OR U625 ( .A(n15633), .B(n15629), .Z(n589) );
  AND U626 ( .A(n588), .B(n589), .Z(n590) );
  ANDN U627 ( .B(n23641), .A(n15639), .Z(n591) );
  NANDN U628 ( .A(n590), .B(n23639), .Z(n592) );
  AND U629 ( .A(n591), .B(n592), .Z(n593) );
  OR U630 ( .A(n23644), .B(n593), .Z(n594) );
  NANDN U631 ( .A(n15638), .B(n7935), .Z(n595) );
  AND U632 ( .A(n594), .B(n595), .Z(n596) );
  NANDN U633 ( .A(n15642), .B(n596), .Z(n7938) );
  OR U634 ( .A(n16035), .B(n16039), .Z(n597) );
  AND U635 ( .A(n8303), .B(n597), .Z(n598) );
  ANDN U636 ( .B(n8302), .A(n12197), .Z(n599) );
  NAND U637 ( .A(n599), .B(n24095), .Z(n600) );
  AND U638 ( .A(n24097), .B(n600), .Z(n601) );
  OR U639 ( .A(n24099), .B(n601), .Z(n602) );
  NAND U640 ( .A(n602), .B(n24101), .Z(n603) );
  ANDN U641 ( .B(n603), .A(n16036), .Z(n604) );
  NAND U642 ( .A(n604), .B(n24103), .Z(n605) );
  NAND U643 ( .A(n605), .B(n24105), .Z(n606) );
  ANDN U644 ( .B(n606), .A(n598), .Z(n607) );
  NANDN U645 ( .A(n607), .B(n24109), .Z(n608) );
  NAND U646 ( .A(n608), .B(n24112), .Z(n609) );
  NAND U647 ( .A(n609), .B(n24113), .Z(n610) );
  NAND U648 ( .A(n610), .B(n24115), .Z(n611) );
  NAND U649 ( .A(n611), .B(n24117), .Z(n612) );
  ANDN U650 ( .B(n612), .A(n24120), .Z(n613) );
  NANDN U651 ( .A(n613), .B(n24121), .Z(n614) );
  ANDN U652 ( .B(n614), .A(n24123), .Z(n8319) );
  NAND U653 ( .A(n9125), .B(n25189), .Z(n615) );
  NANDN U654 ( .A(n25192), .B(n615), .Z(n616) );
  AND U655 ( .A(n25193), .B(n616), .Z(n617) );
  OR U656 ( .A(n25196), .B(n617), .Z(n618) );
  NAND U657 ( .A(n618), .B(n25197), .Z(n619) );
  NANDN U658 ( .A(n25200), .B(n619), .Z(n620) );
  NANDN U659 ( .A(n25202), .B(n620), .Z(n621) );
  NAND U660 ( .A(n621), .B(n25203), .Z(n622) );
  ANDN U661 ( .B(n622), .A(n17066), .Z(n623) );
  NOR U662 ( .A(n623), .B(n25212), .Z(n624) );
  NANDN U663 ( .A(n25207), .B(n20246), .Z(n625) );
  NAND U664 ( .A(n624), .B(n625), .Z(n626) );
  AND U665 ( .A(n25215), .B(n626), .Z(n627) );
  NANDN U666 ( .A(n17071), .B(n17074), .Z(n628) );
  AND U667 ( .A(n627), .B(n628), .Z(n629) );
  NANDN U668 ( .A(n629), .B(n25218), .Z(n630) );
  NAND U669 ( .A(n630), .B(n25219), .Z(n631) );
  NAND U670 ( .A(n631), .B(n25222), .Z(n632) );
  AND U671 ( .A(n25223), .B(n632), .Z(n9131) );
  XOR U672 ( .A(y[2598]), .B(n17246), .Z(n633) );
  NANDN U673 ( .A(n9231), .B(n633), .Z(n634) );
  NAND U674 ( .A(y[2598]), .B(n17246), .Z(n635) );
  AND U675 ( .A(n634), .B(n635), .Z(n636) );
  XNOR U676 ( .A(x[2599]), .B(y[2599]), .Z(n637) );
  NANDN U677 ( .A(n636), .B(n637), .Z(n638) );
  AND U678 ( .A(n11942), .B(n638), .Z(n639) );
  ANDN U679 ( .B(n11943), .A(n11939), .Z(n640) );
  XNOR U680 ( .A(x[2600]), .B(y[2600]), .Z(n641) );
  NANDN U681 ( .A(n639), .B(n641), .Z(n642) );
  AND U682 ( .A(n640), .B(n642), .Z(n643) );
  NOR U683 ( .A(n643), .B(n11940), .Z(n644) );
  NAND U684 ( .A(n644), .B(n25411), .Z(n645) );
  ANDN U685 ( .B(n645), .A(n25414), .Z(n646) );
  NANDN U686 ( .A(n2802), .B(n11938), .Z(n647) );
  AND U687 ( .A(n646), .B(n647), .Z(n648) );
  NANDN U688 ( .A(n648), .B(n25415), .Z(n649) );
  NANDN U689 ( .A(n25418), .B(n649), .Z(n650) );
  NAND U690 ( .A(n650), .B(n25419), .Z(n9240) );
  NAND U691 ( .A(n9801), .B(n26238), .Z(n651) );
  ANDN U692 ( .B(n651), .A(n26240), .Z(n652) );
  ANDN U693 ( .B(n26244), .A(n17949), .Z(n653) );
  OR U694 ( .A(n26243), .B(n652), .Z(n654) );
  AND U695 ( .A(n653), .B(n654), .Z(n655) );
  ANDN U696 ( .B(n26252), .A(n17950), .Z(n656) );
  NOR U697 ( .A(n655), .B(n17953), .Z(n657) );
  NAND U698 ( .A(n657), .B(n26247), .Z(n658) );
  AND U699 ( .A(n656), .B(n658), .Z(n659) );
  NAND U700 ( .A(n17952), .B(n26254), .Z(n660) );
  NANDN U701 ( .A(n9803), .B(n660), .Z(n661) );
  NANDN U702 ( .A(n659), .B(n661), .Z(n662) );
  NAND U703 ( .A(n662), .B(n26256), .Z(n663) );
  NANDN U704 ( .A(n26258), .B(n663), .Z(n664) );
  AND U705 ( .A(n26260), .B(n664), .Z(n665) );
  NOR U706 ( .A(n11735), .B(n26262), .Z(n666) );
  NANDN U707 ( .A(n665), .B(n666), .Z(n667) );
  AND U708 ( .A(n26264), .B(n667), .Z(n9804) );
  ANDN U709 ( .B(n9837), .A(n26362), .Z(n668) );
  ANDN U710 ( .B(n26366), .A(n11706), .Z(n669) );
  OR U711 ( .A(n26365), .B(n668), .Z(n670) );
  NAND U712 ( .A(n669), .B(n670), .Z(n671) );
  ANDN U713 ( .B(n26368), .A(n18067), .Z(n672) );
  NAND U714 ( .A(n672), .B(n671), .Z(n673) );
  NAND U715 ( .A(n673), .B(n26374), .Z(n674) );
  ANDN U716 ( .B(n26377), .A(n18068), .Z(n675) );
  OR U717 ( .A(n11707), .B(n674), .Z(n676) );
  AND U718 ( .A(n675), .B(n676), .Z(n677) );
  NANDN U719 ( .A(n677), .B(n26378), .Z(n678) );
  ANDN U720 ( .B(n678), .A(n26381), .Z(n679) );
  ANDN U721 ( .B(n26384), .A(n11701), .Z(n680) );
  OR U722 ( .A(n26383), .B(n679), .Z(n681) );
  AND U723 ( .A(n680), .B(n681), .Z(n682) );
  NOR U724 ( .A(n682), .B(n18083), .Z(n683) );
  NAND U725 ( .A(n683), .B(n26386), .Z(n684) );
  AND U726 ( .A(n26392), .B(n684), .Z(n685) );
  ANDN U727 ( .B(n685), .A(n11700), .Z(n9839) );
  NAND U728 ( .A(n9844), .B(n9843), .Z(n686) );
  AND U729 ( .A(n26458), .B(n686), .Z(n687) );
  NANDN U730 ( .A(n18155), .B(n687), .Z(n688) );
  NAND U731 ( .A(n688), .B(n26464), .Z(n689) );
  AND U732 ( .A(n26466), .B(n18154), .Z(n690) );
  OR U733 ( .A(n11683), .B(n689), .Z(n691) );
  AND U734 ( .A(n690), .B(n691), .Z(n692) );
  NANDN U735 ( .A(n692), .B(n26468), .Z(n693) );
  ANDN U736 ( .B(n693), .A(n26470), .Z(n694) );
  ANDN U737 ( .B(n26474), .A(n18169), .Z(n695) );
  NANDN U738 ( .A(n694), .B(n26472), .Z(n696) );
  AND U739 ( .A(n695), .B(n696), .Z(n697) );
  NOR U740 ( .A(n697), .B(n18172), .Z(n698) );
  NAND U741 ( .A(n698), .B(n26476), .Z(n699) );
  AND U742 ( .A(n26482), .B(n699), .Z(n700) );
  ANDN U743 ( .B(n26485), .A(n18173), .Z(n701) );
  NANDN U744 ( .A(n18170), .B(n700), .Z(n702) );
  NAND U745 ( .A(n701), .B(n702), .Z(n703) );
  NAND U746 ( .A(n703), .B(n26486), .Z(n9846) );
  ANDN U747 ( .B(n26521), .A(n18213), .Z(n9849) );
  NOR U748 ( .A(n11652), .B(n11655), .Z(n704) );
  NAND U749 ( .A(n704), .B(n9873), .Z(n705) );
  AND U750 ( .A(n26583), .B(n705), .Z(n706) );
  NANDN U751 ( .A(x[3070]), .B(y[3070]), .Z(n707) );
  NANDN U752 ( .A(n11653), .B(n706), .Z(n708) );
  NAND U753 ( .A(n707), .B(n708), .Z(n709) );
  OR U754 ( .A(n11651), .B(n709), .Z(n710) );
  ANDN U755 ( .B(n710), .A(n18274), .Z(n711) );
  NAND U756 ( .A(y[3072]), .B(n11649), .Z(n712) );
  XOR U757 ( .A(n11649), .B(y[3072]), .Z(n713) );
  NAND U758 ( .A(n713), .B(n711), .Z(n714) );
  NAND U759 ( .A(n712), .B(n714), .Z(n715) );
  XNOR U760 ( .A(y[3073]), .B(x[3073]), .Z(n716) );
  NANDN U761 ( .A(n715), .B(n716), .Z(n717) );
  ANDN U762 ( .B(n18279), .A(n11646), .Z(n718) );
  NAND U763 ( .A(n718), .B(n717), .Z(n719) );
  NANDN U764 ( .A(n11648), .B(n719), .Z(n720) );
  XNOR U765 ( .A(y[3075]), .B(x[3075]), .Z(n721) );
  NANDN U766 ( .A(n720), .B(n721), .Z(n9874) );
  NAND U767 ( .A(n9922), .B(n9921), .Z(n722) );
  AND U768 ( .A(n11609), .B(n722), .Z(n723) );
  NANDN U769 ( .A(n11605), .B(n723), .Z(n724) );
  XNOR U770 ( .A(x[3108]), .B(y[3108]), .Z(n725) );
  NANDN U771 ( .A(n11607), .B(n724), .Z(n726) );
  NAND U772 ( .A(n725), .B(n726), .Z(n727) );
  XNOR U773 ( .A(y[3109]), .B(x[3109]), .Z(n728) );
  NAND U774 ( .A(n727), .B(n11602), .Z(n729) );
  NAND U775 ( .A(n728), .B(n729), .Z(n730) );
  ANDN U776 ( .B(n11603), .A(n11600), .Z(n731) );
  NAND U777 ( .A(n731), .B(n730), .Z(n732) );
  ANDN U778 ( .B(n732), .A(n18343), .Z(n733) );
  NANDN U779 ( .A(n11599), .B(n733), .Z(n734) );
  XNOR U780 ( .A(x[3112]), .B(y[3112]), .Z(n735) );
  NANDN U781 ( .A(n11601), .B(n734), .Z(n736) );
  NAND U782 ( .A(n735), .B(n736), .Z(n737) );
  XNOR U783 ( .A(y[3113]), .B(x[3113]), .Z(n738) );
  NAND U784 ( .A(n737), .B(n11596), .Z(n739) );
  NAND U785 ( .A(n738), .B(n739), .Z(n9923) );
  NOR U786 ( .A(n18359), .B(n11578), .Z(n9928) );
  NANDN U787 ( .A(x[1789]), .B(y[1789]), .Z(n12293) );
  NOR U788 ( .A(n9984), .B(n18400), .Z(n740) );
  NAND U789 ( .A(n740), .B(n18404), .Z(n741) );
  ANDN U790 ( .B(n741), .A(n20232), .Z(n742) );
  XNOR U791 ( .A(y[3153]), .B(x[3153]), .Z(n743) );
  AND U792 ( .A(n742), .B(n743), .Z(n744) );
  NOR U793 ( .A(n744), .B(n18410), .Z(n745) );
  NAND U794 ( .A(n745), .B(n11554), .Z(n746) );
  NANDN U795 ( .A(n18407), .B(n746), .Z(n747) );
  XNOR U796 ( .A(y[3155]), .B(x[3155]), .Z(n748) );
  NAND U797 ( .A(n748), .B(n747), .Z(n749) );
  NANDN U798 ( .A(x[3155]), .B(y[3155]), .Z(n750) );
  AND U799 ( .A(n749), .B(n750), .Z(n751) );
  XNOR U800 ( .A(x[3156]), .B(y[3156]), .Z(n752) );
  NANDN U801 ( .A(n751), .B(n752), .Z(n753) );
  ANDN U802 ( .B(n11552), .A(n11547), .Z(n754) );
  NAND U803 ( .A(n754), .B(n753), .Z(n755) );
  NANDN U804 ( .A(n11550), .B(n755), .Z(n756) );
  XNOR U805 ( .A(x[3158]), .B(y[3158]), .Z(n757) );
  NANDN U806 ( .A(n756), .B(n757), .Z(n9985) );
  XNOR U807 ( .A(y[3182]), .B(x[3182]), .Z(n758) );
  NOR U808 ( .A(n18455), .B(n11520), .Z(n759) );
  NANDN U809 ( .A(n11521), .B(n11524), .Z(n760) );
  XNOR U810 ( .A(x[3179]), .B(y[3179]), .Z(n761) );
  XNOR U811 ( .A(y[3178]), .B(x[3178]), .Z(n762) );
  ANDN U812 ( .B(n18448), .A(n18451), .Z(n763) );
  NAND U813 ( .A(n9991), .B(n9990), .Z(n764) );
  AND U814 ( .A(n11527), .B(n764), .Z(n765) );
  NANDN U815 ( .A(n11525), .B(n765), .Z(n766) );
  NAND U816 ( .A(n763), .B(n766), .Z(n767) );
  NANDN U817 ( .A(n11526), .B(n767), .Z(n768) );
  NAND U818 ( .A(n762), .B(n768), .Z(n769) );
  NAND U819 ( .A(n769), .B(n11523), .Z(n770) );
  NAND U820 ( .A(n761), .B(n770), .Z(n771) );
  NANDN U821 ( .A(n760), .B(n771), .Z(n772) );
  NAND U822 ( .A(n759), .B(n772), .Z(n773) );
  NANDN U823 ( .A(n11522), .B(n773), .Z(n774) );
  NAND U824 ( .A(n758), .B(n774), .Z(n775) );
  NAND U825 ( .A(n775), .B(n18460), .Z(n9992) );
  NANDN U826 ( .A(x[1901]), .B(y[1901]), .Z(n15770) );
  XNOR U827 ( .A(y[3206]), .B(x[3206]), .Z(n776) );
  NOR U828 ( .A(n18497), .B(n11489), .Z(n777) );
  NANDN U829 ( .A(n11491), .B(n18495), .Z(n778) );
  XNOR U830 ( .A(x[3203]), .B(y[3203]), .Z(n779) );
  XNOR U831 ( .A(y[3202]), .B(x[3202]), .Z(n780) );
  ANDN U832 ( .B(n10000), .A(n11494), .Z(n781) );
  NAND U833 ( .A(n9999), .B(n9998), .Z(n782) );
  AND U834 ( .A(n11498), .B(n782), .Z(n783) );
  NANDN U835 ( .A(n11495), .B(n783), .Z(n784) );
  NAND U836 ( .A(n781), .B(n784), .Z(n785) );
  NANDN U837 ( .A(n11496), .B(n785), .Z(n786) );
  NAND U838 ( .A(n780), .B(n786), .Z(n787) );
  NAND U839 ( .A(n787), .B(n18494), .Z(n788) );
  NAND U840 ( .A(n779), .B(n788), .Z(n789) );
  NANDN U841 ( .A(n778), .B(n789), .Z(n790) );
  NAND U842 ( .A(n777), .B(n790), .Z(n791) );
  NANDN U843 ( .A(n11492), .B(n791), .Z(n792) );
  NAND U844 ( .A(n776), .B(n792), .Z(n793) );
  NAND U845 ( .A(n793), .B(n11487), .Z(n10001) );
  XNOR U846 ( .A(y[3230]), .B(x[3230]), .Z(n794) );
  NOR U847 ( .A(n18537), .B(n11458), .Z(n795) );
  NANDN U848 ( .A(n11459), .B(n11462), .Z(n796) );
  XNOR U849 ( .A(x[3227]), .B(y[3227]), .Z(n797) );
  XNOR U850 ( .A(y[3226]), .B(x[3226]), .Z(n798) );
  ANDN U851 ( .B(n10009), .A(n11463), .Z(n799) );
  NAND U852 ( .A(n10008), .B(n10007), .Z(n800) );
  AND U853 ( .A(n18529), .B(n800), .Z(n801) );
  NANDN U854 ( .A(n11465), .B(n801), .Z(n802) );
  NAND U855 ( .A(n799), .B(n802), .Z(n803) );
  NANDN U856 ( .A(n11466), .B(n803), .Z(n804) );
  NAND U857 ( .A(n798), .B(n804), .Z(n805) );
  NAND U858 ( .A(n805), .B(n11461), .Z(n806) );
  NAND U859 ( .A(n797), .B(n806), .Z(n807) );
  NANDN U860 ( .A(n796), .B(n807), .Z(n808) );
  NAND U861 ( .A(n795), .B(n808), .Z(n809) );
  NANDN U862 ( .A(n11460), .B(n809), .Z(n810) );
  NAND U863 ( .A(n794), .B(n810), .Z(n811) );
  NAND U864 ( .A(n811), .B(n11455), .Z(n10010) );
  NANDN U865 ( .A(n11433), .B(n11436), .Z(n812) );
  XNOR U866 ( .A(x[3247]), .B(y[3247]), .Z(n813) );
  NAND U867 ( .A(n10015), .B(n11435), .Z(n814) );
  AND U868 ( .A(n813), .B(n814), .Z(n815) );
  NOR U869 ( .A(n18571), .B(n11432), .Z(n816) );
  OR U870 ( .A(n812), .B(n815), .Z(n817) );
  AND U871 ( .A(n816), .B(n817), .Z(n818) );
  XNOR U872 ( .A(x[3250]), .B(y[3250]), .Z(n819) );
  OR U873 ( .A(n11434), .B(n818), .Z(n820) );
  NAND U874 ( .A(n819), .B(n820), .Z(n821) );
  XNOR U875 ( .A(y[3251]), .B(x[3251]), .Z(n822) );
  NAND U876 ( .A(n821), .B(n11429), .Z(n823) );
  NAND U877 ( .A(n822), .B(n823), .Z(n824) );
  ANDN U878 ( .B(n11430), .A(n18580), .Z(n825) );
  NAND U879 ( .A(n825), .B(n824), .Z(n826) );
  ANDN U880 ( .B(n826), .A(n18577), .Z(n827) );
  NANDN U881 ( .A(n11428), .B(n827), .Z(n828) );
  NANDN U882 ( .A(n18581), .B(n828), .Z(n10016) );
  NANDN U883 ( .A(y[3273]), .B(n10027), .Z(n829) );
  NANDN U884 ( .A(n10028), .B(x[3273]), .Z(n830) );
  AND U885 ( .A(n829), .B(n830), .Z(n831) );
  XNOR U886 ( .A(x[3274]), .B(y[3274]), .Z(n832) );
  AND U887 ( .A(n831), .B(n832), .Z(n833) );
  NOR U888 ( .A(n833), .B(n11408), .Z(n834) );
  NAND U889 ( .A(n834), .B(n11411), .Z(n835) );
  ANDN U890 ( .B(n835), .A(n18616), .Z(n836) );
  NAND U891 ( .A(y[3276]), .B(n11407), .Z(n837) );
  XOR U892 ( .A(n11407), .B(y[3276]), .Z(n838) );
  NAND U893 ( .A(n838), .B(n836), .Z(n839) );
  NAND U894 ( .A(n837), .B(n839), .Z(n840) );
  XNOR U895 ( .A(x[3277]), .B(y[3277]), .Z(n841) );
  NAND U896 ( .A(n841), .B(n840), .Z(n842) );
  NAND U897 ( .A(n842), .B(n18621), .Z(n843) );
  NANDN U898 ( .A(n11404), .B(n18622), .Z(n844) );
  XNOR U899 ( .A(y[3278]), .B(x[3278]), .Z(n845) );
  NAND U900 ( .A(n845), .B(n843), .Z(n846) );
  NANDN U901 ( .A(n844), .B(n846), .Z(n10029) );
  NANDN U902 ( .A(n11385), .B(n10031), .Z(n847) );
  NANDN U903 ( .A(y[3292]), .B(x[3292]), .Z(n848) );
  XNOR U904 ( .A(y[3292]), .B(x[3292]), .Z(n849) );
  NAND U905 ( .A(n849), .B(n847), .Z(n850) );
  NAND U906 ( .A(n848), .B(n850), .Z(n851) );
  XNOR U907 ( .A(x[3293]), .B(y[3293]), .Z(n852) );
  NANDN U908 ( .A(n851), .B(n852), .Z(n853) );
  NAND U909 ( .A(n853), .B(n11381), .Z(n854) );
  XNOR U910 ( .A(x[3294]), .B(n854), .Z(n855) );
  NANDN U911 ( .A(y[3294]), .B(n855), .Z(n856) );
  NANDN U912 ( .A(n854), .B(x[3294]), .Z(n857) );
  AND U913 ( .A(n856), .B(n857), .Z(n858) );
  XNOR U914 ( .A(x[3295]), .B(y[3295]), .Z(n859) );
  NAND U915 ( .A(n859), .B(n858), .Z(n860) );
  NAND U916 ( .A(n860), .B(n11377), .Z(n861) );
  NANDN U917 ( .A(n18655), .B(n11378), .Z(n862) );
  XNOR U918 ( .A(y[3296]), .B(x[3296]), .Z(n863) );
  NAND U919 ( .A(n863), .B(n861), .Z(n864) );
  NANDN U920 ( .A(n862), .B(n864), .Z(n10032) );
  ANDN U921 ( .B(n10034), .A(n18672), .Z(n865) );
  XOR U922 ( .A(y[3310]), .B(n11356), .Z(n866) );
  NAND U923 ( .A(n866), .B(n865), .Z(n867) );
  NAND U924 ( .A(y[3310]), .B(n11356), .Z(n868) );
  AND U925 ( .A(n867), .B(n868), .Z(n869) );
  XNOR U926 ( .A(x[3311]), .B(y[3311]), .Z(n870) );
  NANDN U927 ( .A(n869), .B(n870), .Z(n871) );
  NAND U928 ( .A(n871), .B(n11352), .Z(n872) );
  XNOR U929 ( .A(x[3312]), .B(n872), .Z(n873) );
  NANDN U930 ( .A(y[3312]), .B(n873), .Z(n874) );
  NANDN U931 ( .A(n872), .B(x[3312]), .Z(n875) );
  AND U932 ( .A(n874), .B(n875), .Z(n876) );
  XNOR U933 ( .A(x[3313]), .B(y[3313]), .Z(n877) );
  NAND U934 ( .A(n877), .B(n876), .Z(n878) );
  NAND U935 ( .A(n878), .B(n11350), .Z(n879) );
  NANDN U936 ( .A(n11348), .B(n11351), .Z(n880) );
  XNOR U937 ( .A(y[3314]), .B(x[3314]), .Z(n881) );
  NAND U938 ( .A(n881), .B(n879), .Z(n882) );
  NANDN U939 ( .A(n880), .B(n882), .Z(n10035) );
  XNOR U940 ( .A(x[3349]), .B(y[3349]), .Z(n883) );
  NOR U941 ( .A(n18736), .B(n11314), .Z(n884) );
  NANDN U942 ( .A(n18739), .B(n11316), .Z(n885) );
  XNOR U943 ( .A(y[3346]), .B(x[3346]), .Z(n886) );
  XNOR U944 ( .A(x[3345]), .B(y[3345]), .Z(n887) );
  ANDN U945 ( .B(n10068), .A(n11318), .Z(n888) );
  NAND U946 ( .A(n10067), .B(n10066), .Z(n889) );
  AND U947 ( .A(n18728), .B(n889), .Z(n890) );
  NANDN U948 ( .A(n11319), .B(n890), .Z(n891) );
  NAND U949 ( .A(n888), .B(n891), .Z(n892) );
  NANDN U950 ( .A(n11320), .B(n892), .Z(n893) );
  NAND U951 ( .A(n887), .B(n893), .Z(n894) );
  NAND U952 ( .A(n894), .B(n11315), .Z(n895) );
  NAND U953 ( .A(n886), .B(n895), .Z(n896) );
  NANDN U954 ( .A(n885), .B(n896), .Z(n897) );
  NAND U955 ( .A(n884), .B(n897), .Z(n898) );
  NANDN U956 ( .A(n18740), .B(n898), .Z(n899) );
  NAND U957 ( .A(n883), .B(n899), .Z(n900) );
  NAND U958 ( .A(n900), .B(n11311), .Z(n10069) );
  NANDN U959 ( .A(n18773), .B(n10071), .Z(n901) );
  ANDN U960 ( .B(n901), .A(n27194), .Z(n902) );
  XNOR U961 ( .A(y[3367]), .B(x[3367]), .Z(n903) );
  NAND U962 ( .A(n903), .B(n902), .Z(n904) );
  ANDN U963 ( .B(n11296), .A(n18781), .Z(n905) );
  NAND U964 ( .A(n905), .B(n904), .Z(n906) );
  NANDN U965 ( .A(n11294), .B(n906), .Z(n907) );
  ANDN U966 ( .B(n18782), .A(n11291), .Z(n908) );
  XNOR U967 ( .A(y[3369]), .B(x[3369]), .Z(n909) );
  NANDN U968 ( .A(n907), .B(n909), .Z(n910) );
  AND U969 ( .A(n908), .B(n910), .Z(n911) );
  NOR U970 ( .A(n11289), .B(n18784), .Z(n912) );
  NANDN U971 ( .A(n911), .B(n912), .Z(n913) );
  ANDN U972 ( .B(n913), .A(n11292), .Z(n914) );
  XNOR U973 ( .A(y[3372]), .B(x[3372]), .Z(n915) );
  NANDN U974 ( .A(n914), .B(n915), .Z(n916) );
  AND U975 ( .A(n11287), .B(n916), .Z(n917) );
  XNOR U976 ( .A(x[3373]), .B(y[3373]), .Z(n918) );
  NANDN U977 ( .A(n917), .B(n918), .Z(n10072) );
  NANDN U978 ( .A(y[2360]), .B(x[2360]), .Z(n919) );
  ANDN U979 ( .B(n919), .A(n16716), .Z(n24833) );
  XNOR U980 ( .A(x[3406]), .B(y[3406]), .Z(n920) );
  NANDN U981 ( .A(n11252), .B(n10101), .Z(n921) );
  NAND U982 ( .A(n920), .B(n921), .Z(n922) );
  XNOR U983 ( .A(y[3407]), .B(x[3407]), .Z(n923) );
  NAND U984 ( .A(n922), .B(n11247), .Z(n924) );
  NAND U985 ( .A(n923), .B(n924), .Z(n925) );
  ANDN U986 ( .B(n11248), .A(n11246), .Z(n926) );
  NAND U987 ( .A(n926), .B(n925), .Z(n927) );
  AND U988 ( .A(n27288), .B(n927), .Z(n928) );
  NANDN U989 ( .A(n18848), .B(n928), .Z(n929) );
  ANDN U990 ( .B(n929), .A(n11245), .Z(n930) );
  XNOR U991 ( .A(x[3410]), .B(y[3410]), .Z(n931) );
  AND U992 ( .A(n930), .B(n931), .Z(n932) );
  ANDN U993 ( .B(n27286), .A(n932), .Z(n933) );
  XNOR U994 ( .A(x[3411]), .B(y[3411]), .Z(n934) );
  NAND U995 ( .A(n933), .B(n934), .Z(n935) );
  ANDN U996 ( .B(n11242), .A(n18858), .Z(n936) );
  NAND U997 ( .A(n936), .B(n935), .Z(n937) );
  NANDN U998 ( .A(n18855), .B(n937), .Z(n10103) );
  XOR U999 ( .A(y[3420]), .B(n11231), .Z(n938) );
  NANDN U1000 ( .A(n10106), .B(n938), .Z(n939) );
  NAND U1001 ( .A(y[3420]), .B(n11231), .Z(n940) );
  AND U1002 ( .A(n939), .B(n940), .Z(n941) );
  XNOR U1003 ( .A(x[3421]), .B(y[3421]), .Z(n942) );
  NANDN U1004 ( .A(n941), .B(n942), .Z(n943) );
  NAND U1005 ( .A(n943), .B(n11227), .Z(n944) );
  NANDN U1006 ( .A(n944), .B(x[3422]), .Z(n945) );
  XNOR U1007 ( .A(n944), .B(x[3422]), .Z(n946) );
  NANDN U1008 ( .A(y[3422]), .B(n946), .Z(n947) );
  NAND U1009 ( .A(n945), .B(n947), .Z(n948) );
  XNOR U1010 ( .A(x[3423]), .B(y[3423]), .Z(n949) );
  NANDN U1011 ( .A(n948), .B(n949), .Z(n950) );
  AND U1012 ( .A(n11225), .B(n950), .Z(n951) );
  XNOR U1013 ( .A(y[3424]), .B(x[3424]), .Z(n952) );
  NANDN U1014 ( .A(n951), .B(n952), .Z(n953) );
  ANDN U1015 ( .B(n11226), .A(n11223), .Z(n954) );
  NAND U1016 ( .A(n954), .B(n953), .Z(n955) );
  NANDN U1017 ( .A(n18880), .B(n955), .Z(n10107) );
  NANDN U1018 ( .A(x[2450]), .B(y[2450]), .Z(n956) );
  ANDN U1019 ( .B(n956), .A(n16937), .Z(n25057) );
  NAND U1020 ( .A(n10129), .B(n10128), .Z(n957) );
  AND U1021 ( .A(n11208), .B(n957), .Z(n958) );
  NANDN U1022 ( .A(n11205), .B(n958), .Z(n959) );
  ANDN U1023 ( .B(n10130), .A(n11204), .Z(n960) );
  NAND U1024 ( .A(n960), .B(n959), .Z(n961) );
  NANDN U1025 ( .A(n11206), .B(n961), .Z(n962) );
  XNOR U1026 ( .A(x[3443]), .B(y[3443]), .Z(n963) );
  NAND U1027 ( .A(n963), .B(n962), .Z(n964) );
  NAND U1028 ( .A(n964), .B(n18917), .Z(n965) );
  NANDN U1029 ( .A(n18923), .B(n18918), .Z(n966) );
  XNOR U1030 ( .A(y[3444]), .B(x[3444]), .Z(n967) );
  NAND U1031 ( .A(n967), .B(n965), .Z(n968) );
  NANDN U1032 ( .A(n966), .B(n968), .Z(n969) );
  NOR U1033 ( .A(n18920), .B(n11202), .Z(n970) );
  NAND U1034 ( .A(n970), .B(n969), .Z(n971) );
  NANDN U1035 ( .A(n18924), .B(n971), .Z(n972) );
  XNOR U1036 ( .A(x[3447]), .B(y[3447]), .Z(n973) );
  NAND U1037 ( .A(n973), .B(n972), .Z(n974) );
  NAND U1038 ( .A(n974), .B(n11199), .Z(n10131) );
  NAND U1039 ( .A(n10137), .B(n10136), .Z(n975) );
  AND U1040 ( .A(n18960), .B(n975), .Z(n976) );
  NANDN U1041 ( .A(n18965), .B(n976), .Z(n977) );
  NOR U1042 ( .A(n18962), .B(n11184), .Z(n978) );
  NAND U1043 ( .A(n978), .B(n977), .Z(n979) );
  NANDN U1044 ( .A(n18966), .B(n979), .Z(n980) );
  XNOR U1045 ( .A(x[3467]), .B(y[3467]), .Z(n981) );
  NAND U1046 ( .A(n981), .B(n980), .Z(n982) );
  NAND U1047 ( .A(n982), .B(n11182), .Z(n983) );
  NAND U1048 ( .A(n27410), .B(n11181), .Z(n984) );
  XNOR U1049 ( .A(y[3468]), .B(x[3468]), .Z(n985) );
  NAND U1050 ( .A(n985), .B(n983), .Z(n986) );
  NANDN U1051 ( .A(n984), .B(n986), .Z(n987) );
  ANDN U1052 ( .B(n987), .A(n18971), .Z(n988) );
  XNOR U1053 ( .A(x[3470]), .B(y[3470]), .Z(n989) );
  AND U1054 ( .A(n988), .B(n989), .Z(n990) );
  ANDN U1055 ( .B(n27408), .A(n990), .Z(n991) );
  XNOR U1056 ( .A(x[3471]), .B(y[3471]), .Z(n992) );
  NAND U1057 ( .A(n991), .B(n992), .Z(n10138) );
  NANDN U1058 ( .A(y[3486]), .B(x[3486]), .Z(n993) );
  XNOR U1059 ( .A(x[3486]), .B(y[3486]), .Z(n994) );
  NAND U1060 ( .A(n994), .B(n10141), .Z(n995) );
  NAND U1061 ( .A(n993), .B(n995), .Z(n996) );
  ANDN U1062 ( .B(n996), .A(n11160), .Z(n997) );
  OR U1063 ( .A(n11163), .B(n997), .Z(n998) );
  NANDN U1064 ( .A(n11161), .B(n998), .Z(n999) );
  NAND U1065 ( .A(n999), .B(n27450), .Z(n1000) );
  NAND U1066 ( .A(n1000), .B(n27452), .Z(n1001) );
  NAND U1067 ( .A(n1001), .B(n27455), .Z(n1002) );
  AND U1068 ( .A(n27456), .B(n1002), .Z(n1003) );
  NANDN U1069 ( .A(n1003), .B(n27459), .Z(n1004) );
  NANDN U1070 ( .A(n19018), .B(n1004), .Z(n1005) );
  NANDN U1071 ( .A(n11159), .B(n1005), .Z(n1006) );
  NANDN U1072 ( .A(n19019), .B(n1006), .Z(n1007) );
  NANDN U1073 ( .A(x[3495]), .B(y[3495]), .Z(n1008) );
  XNOR U1074 ( .A(x[3495]), .B(y[3495]), .Z(n1009) );
  NAND U1075 ( .A(n1009), .B(n1007), .Z(n1010) );
  NAND U1076 ( .A(n1008), .B(n1010), .Z(n10150) );
  NAND U1077 ( .A(y[3512]), .B(n11135), .Z(n1011) );
  ANDN U1078 ( .B(n1011), .A(n11134), .Z(n1012) );
  XOR U1079 ( .A(n11135), .B(y[3512]), .Z(n1013) );
  NANDN U1080 ( .A(n11137), .B(n10152), .Z(n1014) );
  ANDN U1081 ( .B(n1014), .A(n19048), .Z(n1015) );
  NAND U1082 ( .A(n1013), .B(n1015), .Z(n1016) );
  NAND U1083 ( .A(n1012), .B(n1016), .Z(n1017) );
  AND U1084 ( .A(n19053), .B(n1017), .Z(n1018) );
  NANDN U1085 ( .A(x[3514]), .B(n1018), .Z(n1019) );
  ANDN U1086 ( .B(n1019), .A(n11130), .Z(n1020) );
  XNOR U1087 ( .A(n1018), .B(x[3514]), .Z(n1021) );
  NAND U1088 ( .A(n1021), .B(y[3514]), .Z(n1022) );
  NAND U1089 ( .A(n1020), .B(n1022), .Z(n1023) );
  AND U1090 ( .A(n11132), .B(n1023), .Z(n1024) );
  NANDN U1091 ( .A(x[3516]), .B(n1024), .Z(n1025) );
  ANDN U1092 ( .B(n1025), .A(n19063), .Z(n1026) );
  XNOR U1093 ( .A(n1024), .B(x[3516]), .Z(n1027) );
  NAND U1094 ( .A(n1027), .B(y[3516]), .Z(n1028) );
  NAND U1095 ( .A(n1026), .B(n1028), .Z(n10153) );
  ANDN U1096 ( .B(n19094), .A(n19091), .Z(n1029) );
  NAND U1097 ( .A(n1029), .B(n10155), .Z(n1030) );
  NANDN U1098 ( .A(n27540), .B(n1030), .Z(n1031) );
  OR U1099 ( .A(n19101), .B(n1031), .Z(n1032) );
  ANDN U1100 ( .B(n1032), .A(n19096), .Z(n1033) );
  NAND U1101 ( .A(n19099), .B(y[3534]), .Z(n1034) );
  ANDN U1102 ( .B(n1034), .A(n11116), .Z(n1035) );
  XOR U1103 ( .A(y[3534]), .B(n19099), .Z(n1036) );
  NAND U1104 ( .A(n1036), .B(n1033), .Z(n1037) );
  NAND U1105 ( .A(n1035), .B(n1037), .Z(n1038) );
  ANDN U1106 ( .B(n1038), .A(n19103), .Z(n1039) );
  NANDN U1107 ( .A(x[3536]), .B(n1039), .Z(n1040) );
  ANDN U1108 ( .B(n1040), .A(n11114), .Z(n1041) );
  XNOR U1109 ( .A(n1039), .B(x[3536]), .Z(n1042) );
  NAND U1110 ( .A(n1042), .B(y[3536]), .Z(n1043) );
  NAND U1111 ( .A(n1041), .B(n1043), .Z(n1044) );
  NANDN U1112 ( .A(n19107), .B(n1044), .Z(n10157) );
  AND U1113 ( .A(n10159), .B(n10160), .Z(n1045) );
  NAND U1114 ( .A(n11091), .B(y[3552]), .Z(n1046) );
  ANDN U1115 ( .B(n1046), .A(n11090), .Z(n1047) );
  XOR U1116 ( .A(y[3552]), .B(n11091), .Z(n1048) );
  NAND U1117 ( .A(n1048), .B(n1045), .Z(n1049) );
  NAND U1118 ( .A(n1047), .B(n1049), .Z(n1050) );
  ANDN U1119 ( .B(n1050), .A(n19135), .Z(n1051) );
  NANDN U1120 ( .A(x[3554]), .B(n1051), .Z(n1052) );
  ANDN U1121 ( .B(n1052), .A(n11088), .Z(n1053) );
  XNOR U1122 ( .A(n1051), .B(x[3554]), .Z(n1054) );
  NAND U1123 ( .A(n1054), .B(y[3554]), .Z(n1055) );
  NAND U1124 ( .A(n1053), .B(n1055), .Z(n1056) );
  NANDN U1125 ( .A(n19139), .B(n1056), .Z(n1057) );
  NANDN U1126 ( .A(n1057), .B(y[3556]), .Z(n1058) );
  ANDN U1127 ( .B(n1058), .A(n11083), .Z(n1059) );
  XNOR U1128 ( .A(y[3556]), .B(n1057), .Z(n1060) );
  NAND U1129 ( .A(n1060), .B(n11086), .Z(n1061) );
  AND U1130 ( .A(n1059), .B(n1061), .Z(n10162) );
  NAND U1131 ( .A(n10166), .B(n10165), .Z(n1062) );
  AND U1132 ( .A(n19177), .B(n1062), .Z(n1063) );
  NANDN U1133 ( .A(n11062), .B(n1063), .Z(n1064) );
  ANDN U1134 ( .B(n10167), .A(n11060), .Z(n1065) );
  NAND U1135 ( .A(n1065), .B(n1064), .Z(n1066) );
  ANDN U1136 ( .B(n1066), .A(n11063), .Z(n1067) );
  NANDN U1137 ( .A(n11058), .B(n1067), .Z(n1068) );
  NOR U1138 ( .A(n11061), .B(n11057), .Z(n1069) );
  NAND U1139 ( .A(n1069), .B(n1068), .Z(n1070) );
  AND U1140 ( .A(n11059), .B(n1070), .Z(n1071) );
  OR U1141 ( .A(y[3580]), .B(n1071), .Z(n1072) );
  XOR U1142 ( .A(n1071), .B(y[3580]), .Z(n1073) );
  NAND U1143 ( .A(n1073), .B(x[3580]), .Z(n1074) );
  NAND U1144 ( .A(n1072), .B(n1074), .Z(n1075) );
  ANDN U1145 ( .B(n1075), .A(n11055), .Z(n1076) );
  NOR U1146 ( .A(n1076), .B(n19186), .Z(n1077) );
  NAND U1147 ( .A(n1077), .B(n11052), .Z(n1078) );
  ANDN U1148 ( .B(n1078), .A(n27653), .Z(n1079) );
  ANDN U1149 ( .B(n1079), .A(n11054), .Z(n10169) );
  NANDN U1150 ( .A(n11031), .B(n10173), .Z(n1080) );
  ANDN U1151 ( .B(n1080), .A(n27690), .Z(n1081) );
  NOR U1152 ( .A(n19222), .B(n11028), .Z(n1082) );
  NANDN U1153 ( .A(n11030), .B(n1081), .Z(n1083) );
  AND U1154 ( .A(n1082), .B(n1083), .Z(n1084) );
  NOR U1155 ( .A(n1084), .B(n27701), .Z(n1085) );
  NAND U1156 ( .A(n1085), .B(n11029), .Z(n1086) );
  ANDN U1157 ( .B(n1086), .A(n11026), .Z(n1087) );
  ANDN U1158 ( .B(n27708), .A(n27700), .Z(n1088) );
  NANDN U1159 ( .A(n11027), .B(n1087), .Z(n1089) );
  NAND U1160 ( .A(n1088), .B(n1089), .Z(n1090) );
  NAND U1161 ( .A(n1090), .B(n19233), .Z(n1091) );
  ANDN U1162 ( .B(n27707), .A(n19236), .Z(n1092) );
  OR U1163 ( .A(n19229), .B(n1091), .Z(n1093) );
  AND U1164 ( .A(n1092), .B(n1093), .Z(n1094) );
  NOR U1165 ( .A(n1094), .B(n11024), .Z(n1095) );
  NANDN U1166 ( .A(n19239), .B(n1095), .Z(n1096) );
  NANDN U1167 ( .A(n19237), .B(n1096), .Z(n10175) );
  ANDN U1168 ( .B(n19268), .A(n11006), .Z(n1097) );
  NAND U1169 ( .A(n10180), .B(n10179), .Z(n1098) );
  AND U1170 ( .A(n1097), .B(n1098), .Z(n1099) );
  NOR U1171 ( .A(n11007), .B(n11003), .Z(n1100) );
  NOR U1172 ( .A(n1099), .B(n11005), .Z(n1101) );
  NAND U1173 ( .A(n1101), .B(n10181), .Z(n1102) );
  AND U1174 ( .A(n1100), .B(n1102), .Z(n1103) );
  NOR U1175 ( .A(n27755), .B(n11004), .Z(n1104) );
  NANDN U1176 ( .A(n1103), .B(n1104), .Z(n1105) );
  ANDN U1177 ( .B(n1105), .A(n11001), .Z(n1106) );
  NOR U1178 ( .A(n19281), .B(n27754), .Z(n1107) );
  NANDN U1179 ( .A(n11002), .B(n1106), .Z(n1108) );
  NAND U1180 ( .A(n1107), .B(n1108), .Z(n1109) );
  NOR U1181 ( .A(n19285), .B(n19278), .Z(n1110) );
  NAND U1182 ( .A(n1110), .B(n1109), .Z(n1111) );
  AND U1183 ( .A(n20223), .B(n1111), .Z(n1112) );
  NANDN U1184 ( .A(n19282), .B(n1112), .Z(n10182) );
  NANDN U1185 ( .A(n10962), .B(n10965), .Z(n1113) );
  ANDN U1186 ( .B(n19353), .A(n10960), .Z(n1114) );
  NANDN U1187 ( .A(n1113), .B(n10208), .Z(n1115) );
  AND U1188 ( .A(n1114), .B(n1115), .Z(n1116) );
  NOR U1189 ( .A(n1116), .B(n19357), .Z(n1117) );
  NANDN U1190 ( .A(n10963), .B(n1117), .Z(n1118) );
  NANDN U1191 ( .A(n10961), .B(n1118), .Z(n1119) );
  OR U1192 ( .A(n10959), .B(n1119), .Z(n1120) );
  AND U1193 ( .A(n19358), .B(n1120), .Z(n1121) );
  NAND U1194 ( .A(n10957), .B(y[3670]), .Z(n1122) );
  ANDN U1195 ( .B(n1122), .A(n10956), .Z(n1123) );
  XOR U1196 ( .A(y[3670]), .B(n10957), .Z(n1124) );
  NAND U1197 ( .A(n1124), .B(n1121), .Z(n1125) );
  NAND U1198 ( .A(n1123), .B(n1125), .Z(n1126) );
  NAND U1199 ( .A(n1126), .B(n19362), .Z(n1127) );
  NANDN U1200 ( .A(y[3672]), .B(x[3672]), .Z(n1128) );
  XNOR U1201 ( .A(y[3672]), .B(x[3672]), .Z(n1129) );
  NAND U1202 ( .A(n1129), .B(n1127), .Z(n1130) );
  NAND U1203 ( .A(n1128), .B(n1130), .Z(n10209) );
  ANDN U1204 ( .B(n10211), .A(n19388), .Z(n1131) );
  NAND U1205 ( .A(y[3686]), .B(n19391), .Z(n1132) );
  ANDN U1206 ( .B(n1132), .A(n10939), .Z(n1133) );
  XOR U1207 ( .A(n19391), .B(y[3686]), .Z(n1134) );
  NAND U1208 ( .A(n1134), .B(n1131), .Z(n1135) );
  NAND U1209 ( .A(n1133), .B(n1135), .Z(n1136) );
  ANDN U1210 ( .B(n1136), .A(n19395), .Z(n1137) );
  NANDN U1211 ( .A(x[3688]), .B(n1137), .Z(n1138) );
  ANDN U1212 ( .B(n1138), .A(n10937), .Z(n1139) );
  XNOR U1213 ( .A(n1137), .B(x[3688]), .Z(n1140) );
  NAND U1214 ( .A(n1140), .B(y[3688]), .Z(n1141) );
  NAND U1215 ( .A(n1139), .B(n1141), .Z(n1142) );
  ANDN U1216 ( .B(n1142), .A(n19399), .Z(n1143) );
  XOR U1217 ( .A(y[3690]), .B(n10935), .Z(n1144) );
  NAND U1218 ( .A(n1144), .B(n1143), .Z(n1145) );
  NAND U1219 ( .A(y[3690]), .B(n10935), .Z(n1146) );
  AND U1220 ( .A(n1145), .B(n1146), .Z(n10212) );
  NANDN U1221 ( .A(n19439), .B(n10215), .Z(n1147) );
  NANDN U1222 ( .A(n19434), .B(n1147), .Z(n1148) );
  NANDN U1223 ( .A(n1148), .B(y[3706]), .Z(n1149) );
  ANDN U1224 ( .B(n1149), .A(n19446), .Z(n1150) );
  XNOR U1225 ( .A(n1148), .B(y[3706]), .Z(n1151) );
  NAND U1226 ( .A(n1151), .B(n19437), .Z(n1152) );
  NAND U1227 ( .A(n1150), .B(n1152), .Z(n1153) );
  ANDN U1228 ( .B(n1153), .A(n19441), .Z(n1154) );
  NAND U1229 ( .A(n19444), .B(y[3708]), .Z(n1155) );
  ANDN U1230 ( .B(n1155), .A(n19450), .Z(n1156) );
  XOR U1231 ( .A(y[3708]), .B(n19444), .Z(n1157) );
  NAND U1232 ( .A(n1157), .B(n1154), .Z(n1158) );
  AND U1233 ( .A(n1156), .B(n1158), .Z(n1159) );
  NOR U1234 ( .A(n10922), .B(n19453), .Z(n1160) );
  NANDN U1235 ( .A(n1159), .B(n1160), .Z(n1161) );
  ANDN U1236 ( .B(n1161), .A(n27937), .Z(n1162) );
  ANDN U1237 ( .B(n1162), .A(n19449), .Z(n10217) );
  NOR U1238 ( .A(n27977), .B(n27968), .Z(n1163) );
  NAND U1239 ( .A(n1163), .B(n10219), .Z(n1164) );
  ANDN U1240 ( .B(n1164), .A(n10907), .Z(n1165) );
  ANDN U1241 ( .B(n27975), .A(n10904), .Z(n1166) );
  NANDN U1242 ( .A(n19488), .B(n1165), .Z(n1167) );
  NAND U1243 ( .A(n1166), .B(n1167), .Z(n1168) );
  ANDN U1244 ( .B(n1168), .A(n10905), .Z(n1169) );
  NANDN U1245 ( .A(x[3730]), .B(n1169), .Z(n1170) );
  ANDN U1246 ( .B(n1170), .A(n10902), .Z(n1171) );
  XNOR U1247 ( .A(n1169), .B(x[3730]), .Z(n1172) );
  NAND U1248 ( .A(n1172), .B(y[3730]), .Z(n1173) );
  NAND U1249 ( .A(n1171), .B(n1173), .Z(n1174) );
  NANDN U1250 ( .A(n19495), .B(n1174), .Z(n1175) );
  NANDN U1251 ( .A(n1175), .B(y[3732]), .Z(n1176) );
  ANDN U1252 ( .B(n1176), .A(n10897), .Z(n1177) );
  XNOR U1253 ( .A(n1175), .B(y[3732]), .Z(n1178) );
  NAND U1254 ( .A(n1178), .B(n10900), .Z(n1179) );
  NAND U1255 ( .A(n1177), .B(n1179), .Z(n10220) );
  ANDN U1256 ( .B(n10223), .A(n19537), .Z(n1180) );
  NOR U1257 ( .A(n19535), .B(n19528), .Z(n1181) );
  NAND U1258 ( .A(n1181), .B(n10222), .Z(n1182) );
  AND U1259 ( .A(n1180), .B(n1182), .Z(n1183) );
  NOR U1260 ( .A(n10878), .B(n19534), .Z(n1184) );
  NANDN U1261 ( .A(n1183), .B(n1184), .Z(n1185) );
  ANDN U1262 ( .B(n1185), .A(n19538), .Z(n1186) );
  NAND U1263 ( .A(n10877), .B(x[3753]), .Z(n1187) );
  ANDN U1264 ( .B(n1187), .A(n19544), .Z(n1188) );
  XOR U1265 ( .A(x[3753]), .B(n10877), .Z(n1189) );
  NAND U1266 ( .A(n1189), .B(n1186), .Z(n1190) );
  NAND U1267 ( .A(n1188), .B(n1190), .Z(n1191) );
  ANDN U1268 ( .B(n1191), .A(n19541), .Z(n1192) );
  NANDN U1269 ( .A(y[3755]), .B(n1192), .Z(n1193) );
  ANDN U1270 ( .B(n1193), .A(n10875), .Z(n1194) );
  XNOR U1271 ( .A(n1192), .B(y[3755]), .Z(n1195) );
  NAND U1272 ( .A(n1195), .B(x[3755]), .Z(n1196) );
  NAND U1273 ( .A(n1194), .B(n1196), .Z(n10224) );
  NANDN U1274 ( .A(n10858), .B(n10228), .Z(n1197) );
  ANDN U1275 ( .B(n1197), .A(n10229), .Z(n1198) );
  NOR U1276 ( .A(n1198), .B(n10856), .Z(n1199) );
  NAND U1277 ( .A(n1199), .B(n28066), .Z(n1200) );
  ANDN U1278 ( .B(n1200), .A(n19580), .Z(n1201) );
  NANDN U1279 ( .A(x[3774]), .B(n1201), .Z(n1202) );
  ANDN U1280 ( .B(n1202), .A(n19586), .Z(n1203) );
  XNOR U1281 ( .A(n1201), .B(x[3774]), .Z(n1204) );
  NAND U1282 ( .A(n1204), .B(y[3774]), .Z(n1205) );
  NAND U1283 ( .A(n1203), .B(n1205), .Z(n1206) );
  NOR U1284 ( .A(n10854), .B(n19589), .Z(n1207) );
  NAND U1285 ( .A(n1207), .B(n1206), .Z(n1208) );
  NANDN U1286 ( .A(n28083), .B(n1208), .Z(n1209) );
  OR U1287 ( .A(n19585), .B(n1209), .Z(n1210) );
  ANDN U1288 ( .B(n1210), .A(n10852), .Z(n1211) );
  ANDN U1289 ( .B(n28081), .A(n10851), .Z(n1212) );
  NANDN U1290 ( .A(n19588), .B(n1211), .Z(n1213) );
  NAND U1291 ( .A(n1212), .B(n1213), .Z(n10230) );
  NOR U1292 ( .A(n20214), .B(n10838), .Z(n1214) );
  OR U1293 ( .A(n10233), .B(n10234), .Z(n1215) );
  AND U1294 ( .A(n1214), .B(n1215), .Z(n1216) );
  NOR U1295 ( .A(n10835), .B(n10837), .Z(n1217) );
  NANDN U1296 ( .A(n1216), .B(n1217), .Z(n1218) );
  AND U1297 ( .A(n28119), .B(n1218), .Z(n1219) );
  ANDN U1298 ( .B(n19629), .A(n10833), .Z(n1220) );
  NANDN U1299 ( .A(n20215), .B(n1219), .Z(n1221) );
  NAND U1300 ( .A(n1220), .B(n1221), .Z(n1222) );
  NOR U1301 ( .A(n10832), .B(n28118), .Z(n1223) );
  NAND U1302 ( .A(n1223), .B(n1222), .Z(n1224) );
  ANDN U1303 ( .B(n1224), .A(n19631), .Z(n1225) );
  NANDN U1304 ( .A(x[3798]), .B(n1225), .Z(n1226) );
  ANDN U1305 ( .B(n1226), .A(n10829), .Z(n1227) );
  XNOR U1306 ( .A(n1225), .B(x[3798]), .Z(n1228) );
  NAND U1307 ( .A(n1228), .B(y[3798]), .Z(n1229) );
  NAND U1308 ( .A(n1227), .B(n1229), .Z(n1230) );
  NANDN U1309 ( .A(n19635), .B(n1230), .Z(n10236) );
  AND U1310 ( .A(n10298), .B(n10299), .Z(n1231) );
  NANDN U1311 ( .A(x[3866]), .B(n1231), .Z(n1232) );
  ANDN U1312 ( .B(n1232), .A(n10743), .Z(n1233) );
  XNOR U1313 ( .A(n1231), .B(x[3866]), .Z(n1234) );
  NAND U1314 ( .A(n1234), .B(y[3866]), .Z(n1235) );
  NAND U1315 ( .A(n1233), .B(n1235), .Z(n1236) );
  ANDN U1316 ( .B(n1236), .A(n19751), .Z(n1237) );
  NAND U1317 ( .A(n10741), .B(y[3868]), .Z(n1238) );
  ANDN U1318 ( .B(n1238), .A(n19757), .Z(n1239) );
  XOR U1319 ( .A(y[3868]), .B(n10741), .Z(n1240) );
  NAND U1320 ( .A(n1240), .B(n1237), .Z(n1241) );
  NAND U1321 ( .A(n1239), .B(n1241), .Z(n1242) );
  ANDN U1322 ( .B(n1242), .A(n10739), .Z(n1243) );
  NANDN U1323 ( .A(x[3870]), .B(n1243), .Z(n1244) );
  ANDN U1324 ( .B(n1244), .A(n19764), .Z(n1245) );
  XNOR U1325 ( .A(n1243), .B(x[3870]), .Z(n1246) );
  NAND U1326 ( .A(n1246), .B(y[3870]), .Z(n1247) );
  NAND U1327 ( .A(n1245), .B(n1247), .Z(n10300) );
  NAND U1328 ( .A(n10324), .B(n10325), .Z(n1248) );
  ANDN U1329 ( .B(n1248), .A(n10702), .Z(n1249) );
  NANDN U1330 ( .A(n10701), .B(n1249), .Z(n1250) );
  AND U1331 ( .A(n28347), .B(n1250), .Z(n1251) );
  NANDN U1332 ( .A(y[3901]), .B(n1251), .Z(n1252) );
  ANDN U1333 ( .B(n1252), .A(n19822), .Z(n1253) );
  XNOR U1334 ( .A(n1251), .B(y[3901]), .Z(n1254) );
  NAND U1335 ( .A(n1254), .B(x[3901]), .Z(n1255) );
  NAND U1336 ( .A(n1253), .B(n1255), .Z(n1256) );
  ANDN U1337 ( .B(n28357), .A(n10700), .Z(n1257) );
  NAND U1338 ( .A(n1257), .B(n1256), .Z(n1258) );
  NANDN U1339 ( .A(n19821), .B(n1258), .Z(n1259) );
  ANDN U1340 ( .B(n28356), .A(n10695), .Z(n1260) );
  NANDN U1341 ( .A(n1259), .B(n10698), .Z(n1261) );
  AND U1342 ( .A(n1260), .B(n1261), .Z(n1262) );
  NOR U1343 ( .A(n19829), .B(n10696), .Z(n1263) );
  NANDN U1344 ( .A(n1262), .B(n1263), .Z(n1264) );
  AND U1345 ( .A(n20209), .B(n1264), .Z(n1265) );
  ANDN U1346 ( .B(n1265), .A(n10694), .Z(n10326) );
  NOR U1347 ( .A(n19910), .B(n10358), .Z(n1266) );
  XNOR U1348 ( .A(x[3950]), .B(y[3950]), .Z(n1267) );
  NAND U1349 ( .A(n1266), .B(n1267), .Z(n1268) );
  OR U1350 ( .A(n19916), .B(n10642), .Z(n1269) );
  ANDN U1351 ( .B(n28465), .A(n28456), .Z(n1270) );
  NAND U1352 ( .A(n1270), .B(n1268), .Z(n1271) );
  NANDN U1353 ( .A(n1269), .B(n1271), .Z(n1272) );
  OR U1354 ( .A(n10641), .B(n19922), .Z(n1273) );
  NOR U1355 ( .A(n28462), .B(n28470), .Z(n1274) );
  NAND U1356 ( .A(n1274), .B(n1272), .Z(n1275) );
  NANDN U1357 ( .A(n1273), .B(n1275), .Z(n1276) );
  NOR U1358 ( .A(n19927), .B(n28468), .Z(n1277) );
  NAND U1359 ( .A(n1277), .B(n1276), .Z(n1278) );
  NANDN U1360 ( .A(n10639), .B(n1278), .Z(n1279) );
  OR U1361 ( .A(n10637), .B(n1279), .Z(n1280) );
  AND U1362 ( .A(n28479), .B(n1280), .Z(n1281) );
  NOR U1363 ( .A(n19930), .B(n10636), .Z(n1282) );
  NANDN U1364 ( .A(n19926), .B(n1281), .Z(n1283) );
  NAND U1365 ( .A(n1282), .B(n1283), .Z(n10359) );
  NANDN U1366 ( .A(n10364), .B(x[3975]), .Z(n1284) );
  NANDN U1367 ( .A(y[3975]), .B(n10363), .Z(n1285) );
  NAND U1368 ( .A(n1284), .B(n1285), .Z(n1286) );
  OR U1369 ( .A(n10617), .B(n1286), .Z(n1287) );
  ANDN U1370 ( .B(n1287), .A(n19969), .Z(n1288) );
  NAND U1371 ( .A(n10616), .B(x[3977]), .Z(n1289) );
  ANDN U1372 ( .B(n1289), .A(n10614), .Z(n1290) );
  XOR U1373 ( .A(x[3977]), .B(n10616), .Z(n1291) );
  NAND U1374 ( .A(n1291), .B(n1288), .Z(n1292) );
  NAND U1375 ( .A(n1290), .B(n1292), .Z(n1293) );
  NANDN U1376 ( .A(n19973), .B(n1293), .Z(n1294) );
  NANDN U1377 ( .A(x[3979]), .B(y[3979]), .Z(n1295) );
  XNOR U1378 ( .A(x[3979]), .B(y[3979]), .Z(n1296) );
  NAND U1379 ( .A(n1296), .B(n1294), .Z(n1297) );
  NAND U1380 ( .A(n1295), .B(n1297), .Z(n1298) );
  ANDN U1381 ( .B(n28535), .A(n19978), .Z(n1299) );
  NANDN U1382 ( .A(n10613), .B(n1298), .Z(n1300) );
  NAND U1383 ( .A(n1299), .B(n1300), .Z(n10365) );
  NAND U1384 ( .A(n10546), .B(n10448), .Z(n1301) );
  NANDN U1385 ( .A(n10449), .B(y[4046]), .Z(n1302) );
  NAND U1386 ( .A(n1301), .B(n1302), .Z(n1303) );
  OR U1387 ( .A(n20106), .B(n1303), .Z(n1304) );
  ANDN U1388 ( .B(n1304), .A(n20103), .Z(n1305) );
  NANDN U1389 ( .A(x[4048]), .B(y[4048]), .Z(n1306) );
  ANDN U1390 ( .B(n1306), .A(n10543), .Z(n1307) );
  XNOR U1391 ( .A(x[4048]), .B(y[4048]), .Z(n1308) );
  NAND U1392 ( .A(n1308), .B(n1305), .Z(n1309) );
  AND U1393 ( .A(n1307), .B(n1309), .Z(n1310) );
  NOR U1394 ( .A(n10545), .B(n20112), .Z(n1311) );
  NANDN U1395 ( .A(n1310), .B(n1311), .Z(n1312) );
  ANDN U1396 ( .B(n1312), .A(n20200), .Z(n1313) );
  NOR U1397 ( .A(n20111), .B(n10541), .Z(n1314) );
  NANDN U1398 ( .A(n10542), .B(n1313), .Z(n1315) );
  NAND U1399 ( .A(n1314), .B(n1315), .Z(n1316) );
  ANDN U1400 ( .B(n1316), .A(n28690), .Z(n1317) );
  NANDN U1401 ( .A(n20201), .B(n1317), .Z(n10450) );
  NANDN U1402 ( .A(n6218), .B(n14341), .Z(n1318) );
  AND U1403 ( .A(n21908), .B(n1318), .Z(n1319) );
  XOR U1404 ( .A(x[1038]), .B(n6218), .Z(n1320) );
  NAND U1405 ( .A(n1320), .B(y[1038]), .Z(n1321) );
  AND U1406 ( .A(n1319), .B(n1321), .Z(n1322) );
  NOR U1407 ( .A(n21911), .B(n12699), .Z(n1323) );
  NANDN U1408 ( .A(n1322), .B(n1323), .Z(n1324) );
  AND U1409 ( .A(n21912), .B(n1324), .Z(n1325) );
  NOR U1410 ( .A(n1325), .B(n14354), .Z(n1326) );
  NAND U1411 ( .A(n1326), .B(n21914), .Z(n1327) );
  AND U1412 ( .A(n21916), .B(n1327), .Z(n1328) );
  NOR U1413 ( .A(n1328), .B(n14357), .Z(n1329) );
  OR U1414 ( .A(n6220), .B(n14353), .Z(n1330) );
  NAND U1415 ( .A(n1329), .B(n1330), .Z(n1331) );
  NAND U1416 ( .A(n1331), .B(n21920), .Z(n1332) );
  NANDN U1417 ( .A(n21923), .B(n1332), .Z(n1333) );
  AND U1418 ( .A(n21924), .B(n1333), .Z(n1334) );
  OR U1419 ( .A(n21927), .B(n1334), .Z(n1335) );
  ANDN U1420 ( .B(n1335), .A(n12696), .Z(n6231) );
  NANDN U1421 ( .A(n12645), .B(n6410), .Z(n1336) );
  NAND U1422 ( .A(n1336), .B(n22094), .Z(n1337) );
  NANDN U1423 ( .A(n22096), .B(n1337), .Z(n1338) );
  NAND U1424 ( .A(n1338), .B(n22098), .Z(n1339) );
  NANDN U1425 ( .A(n22100), .B(n1339), .Z(n1340) );
  ANDN U1426 ( .B(n1340), .A(n14479), .Z(n1341) );
  NANDN U1427 ( .A(y[1134]), .B(x[1134]), .Z(n1342) );
  XNOR U1428 ( .A(x[1134]), .B(y[1134]), .Z(n1343) );
  NAND U1429 ( .A(n1343), .B(n1341), .Z(n1344) );
  NAND U1430 ( .A(n1342), .B(n1344), .Z(n1345) );
  AND U1431 ( .A(n22106), .B(n1345), .Z(n1346) );
  NOR U1432 ( .A(n1346), .B(n14482), .Z(n1347) );
  NAND U1433 ( .A(n1347), .B(n22108), .Z(n1348) );
  AND U1434 ( .A(n22110), .B(n1348), .Z(n1349) );
  NOR U1435 ( .A(n1349), .B(n12640), .Z(n1350) );
  NAND U1436 ( .A(n1350), .B(n22113), .Z(n1351) );
  AND U1437 ( .A(n22114), .B(n1351), .Z(n1352) );
  OR U1438 ( .A(n12641), .B(n1352), .Z(n1353) );
  NAND U1439 ( .A(n1353), .B(n22118), .Z(n6421) );
  XNOR U1440 ( .A(x[1189]), .B(y[1189]), .Z(n1354) );
  NAND U1441 ( .A(n1354), .B(n6528), .Z(n1355) );
  NAND U1442 ( .A(n1355), .B(n12623), .Z(n1356) );
  NANDN U1443 ( .A(n14569), .B(n1356), .Z(n1357) );
  NAND U1444 ( .A(n1357), .B(n22214), .Z(n1358) );
  ANDN U1445 ( .B(n1358), .A(n22217), .Z(n1359) );
  NANDN U1446 ( .A(n1359), .B(n22218), .Z(n1360) );
  AND U1447 ( .A(n12621), .B(n1360), .Z(n1361) );
  NAND U1448 ( .A(x[1194]), .B(n14575), .Z(n1362) );
  XOR U1449 ( .A(n14575), .B(x[1194]), .Z(n1363) );
  NAND U1450 ( .A(n1363), .B(n1361), .Z(n1364) );
  NAND U1451 ( .A(n1362), .B(n1364), .Z(n1365) );
  AND U1452 ( .A(n22225), .B(n1365), .Z(n1366) );
  NOR U1453 ( .A(n1366), .B(n14576), .Z(n1367) );
  NAND U1454 ( .A(n1367), .B(n22226), .Z(n1368) );
  ANDN U1455 ( .B(n1368), .A(n22229), .Z(n1369) );
  NOR U1456 ( .A(n1369), .B(n14588), .Z(n1370) );
  NAND U1457 ( .A(n1370), .B(n22230), .Z(n1371) );
  ANDN U1458 ( .B(n1371), .A(n22232), .Z(n6537) );
  NAND U1459 ( .A(n7378), .B(n22991), .Z(n1372) );
  NAND U1460 ( .A(n1372), .B(n22993), .Z(n1373) );
  AND U1461 ( .A(n22995), .B(n1373), .Z(n1374) );
  OR U1462 ( .A(n12394), .B(n1374), .Z(n1375) );
  AND U1463 ( .A(n22999), .B(n1375), .Z(n1376) );
  NAND U1464 ( .A(n12393), .B(n23001), .Z(n1377) );
  NANDN U1465 ( .A(n7382), .B(n1377), .Z(n1378) );
  NANDN U1466 ( .A(n1376), .B(n1378), .Z(n1379) );
  NAND U1467 ( .A(n1379), .B(n23003), .Z(n1380) );
  NANDN U1468 ( .A(n23006), .B(n1380), .Z(n1381) );
  AND U1469 ( .A(n23007), .B(n1381), .Z(n1382) );
  NANDN U1470 ( .A(n12387), .B(n1382), .Z(n1383) );
  NAND U1471 ( .A(n1383), .B(n23010), .Z(n1384) );
  ANDN U1472 ( .B(n1384), .A(n12390), .Z(n1385) );
  NANDN U1473 ( .A(n7384), .B(n12386), .Z(n1386) );
  AND U1474 ( .A(n1385), .B(n1386), .Z(n1387) );
  NANDN U1475 ( .A(n1387), .B(n23014), .Z(n1388) );
  NAND U1476 ( .A(n1388), .B(n23015), .Z(n1389) );
  NAND U1477 ( .A(n1389), .B(n23018), .Z(n7394) );
  NAND U1478 ( .A(n8688), .B(n24591), .Z(n1390) );
  AND U1479 ( .A(n24592), .B(n1390), .Z(n1391) );
  NANDN U1480 ( .A(x[2252]), .B(n16500), .Z(n1392) );
  NAND U1481 ( .A(n1392), .B(n8693), .Z(n1393) );
  ANDN U1482 ( .B(n1393), .A(n1391), .Z(n1394) );
  NANDN U1483 ( .A(n1394), .B(n24596), .Z(n1395) );
  NANDN U1484 ( .A(n24598), .B(n1395), .Z(n1396) );
  NAND U1485 ( .A(n1396), .B(n24600), .Z(n1397) );
  NANDN U1486 ( .A(n24603), .B(n1397), .Z(n1398) );
  NAND U1487 ( .A(n1398), .B(n24604), .Z(n1399) );
  ANDN U1488 ( .B(n1399), .A(n24606), .Z(n1400) );
  NANDN U1489 ( .A(n1400), .B(n24608), .Z(n1401) );
  AND U1490 ( .A(n24610), .B(n1401), .Z(n1402) );
  OR U1491 ( .A(n24612), .B(n1402), .Z(n1403) );
  NAND U1492 ( .A(n1403), .B(n24614), .Z(n1404) );
  NAND U1493 ( .A(n1404), .B(n24616), .Z(n1405) );
  ANDN U1494 ( .B(n24618), .A(n16530), .Z(n1406) );
  NAND U1495 ( .A(n1406), .B(n1405), .Z(n1407) );
  NAND U1496 ( .A(n1407), .B(n24621), .Z(n8706) );
  AND U1497 ( .A(n24701), .B(n24697), .Z(n1408) );
  ANDN U1498 ( .B(n8776), .A(n16595), .Z(n1409) );
  NAND U1499 ( .A(n1409), .B(n24694), .Z(n1410) );
  AND U1500 ( .A(n1408), .B(n1410), .Z(n1411) );
  NOR U1501 ( .A(n1411), .B(n16596), .Z(n1412) );
  NAND U1502 ( .A(n1412), .B(n24702), .Z(n1413) );
  AND U1503 ( .A(n24705), .B(n1413), .Z(n1414) );
  NANDN U1504 ( .A(n1414), .B(n24706), .Z(n1415) );
  AND U1505 ( .A(n24708), .B(n1415), .Z(n1416) );
  NANDN U1506 ( .A(n1416), .B(n24710), .Z(n1417) );
  NAND U1507 ( .A(n1417), .B(n24713), .Z(n1418) );
  NAND U1508 ( .A(n1418), .B(n24716), .Z(n1419) );
  AND U1509 ( .A(n24719), .B(n1419), .Z(n1420) );
  OR U1510 ( .A(n12089), .B(n16616), .Z(n1421) );
  AND U1511 ( .A(n1420), .B(n1421), .Z(n1422) );
  NANDN U1512 ( .A(n1422), .B(n24722), .Z(n1423) );
  NANDN U1513 ( .A(n24724), .B(n1423), .Z(n1424) );
  NAND U1514 ( .A(n1424), .B(n24726), .Z(n1425) );
  NAND U1515 ( .A(n1425), .B(n24729), .Z(n8781) );
  AND U1516 ( .A(x[1328]), .B(n20288), .Z(n14773) );
  NANDN U1517 ( .A(n9156), .B(n25263), .Z(n1426) );
  NANDN U1518 ( .A(n25265), .B(n1426), .Z(n1427) );
  NAND U1519 ( .A(n1427), .B(n25267), .Z(n1428) );
  NANDN U1520 ( .A(n25269), .B(n1428), .Z(n1429) );
  NAND U1521 ( .A(n1429), .B(n25271), .Z(n1430) );
  ANDN U1522 ( .B(n1430), .A(n25274), .Z(n1431) );
  NOR U1523 ( .A(n1431), .B(n17127), .Z(n1432) );
  NAND U1524 ( .A(n1432), .B(n25275), .Z(n1433) );
  ANDN U1525 ( .B(n1433), .A(n25278), .Z(n1434) );
  NOR U1526 ( .A(n1434), .B(n17130), .Z(n1435) );
  NANDN U1527 ( .A(n17126), .B(n9163), .Z(n1436) );
  AND U1528 ( .A(n1435), .B(n1436), .Z(n1437) );
  NANDN U1529 ( .A(n1437), .B(n25282), .Z(n1438) );
  NAND U1530 ( .A(n1438), .B(n25283), .Z(n1439) );
  NANDN U1531 ( .A(n25285), .B(n1439), .Z(n1440) );
  NAND U1532 ( .A(n1440), .B(n25287), .Z(n1441) );
  AND U1533 ( .A(n25290), .B(n1441), .Z(n1442) );
  NANDN U1534 ( .A(n11965), .B(n1442), .Z(n1443) );
  AND U1535 ( .A(n25291), .B(n1443), .Z(n9166) );
  ANDN U1536 ( .B(n14158), .A(n14164), .Z(n21623) );
  NANDN U1537 ( .A(x[1304]), .B(y[1304]), .Z(n1444) );
  NANDN U1538 ( .A(n12554), .B(n1444), .Z(n12557) );
  AND U1539 ( .A(n25987), .B(n25982), .Z(n1445) );
  NANDN U1540 ( .A(n11802), .B(n9655), .Z(n1446) );
  AND U1541 ( .A(n1445), .B(n1446), .Z(n1447) );
  NOR U1542 ( .A(n1447), .B(n11803), .Z(n1448) );
  NAND U1543 ( .A(n1448), .B(n25988), .Z(n1449) );
  ANDN U1544 ( .B(n1449), .A(n25990), .Z(n1450) );
  NANDN U1545 ( .A(n1450), .B(n25992), .Z(n1451) );
  NANDN U1546 ( .A(n25994), .B(n1451), .Z(n1452) );
  NAND U1547 ( .A(n1452), .B(n25996), .Z(n1453) );
  ANDN U1548 ( .B(n25999), .A(n17734), .Z(n1454) );
  NAND U1549 ( .A(n1454), .B(n1453), .Z(n1455) );
  NAND U1550 ( .A(n1455), .B(n26000), .Z(n1456) );
  XNOR U1551 ( .A(y[2840]), .B(x[2840]), .Z(n1457) );
  NAND U1552 ( .A(n1457), .B(n1456), .Z(n1458) );
  NAND U1553 ( .A(n1458), .B(n17737), .Z(n1459) );
  NAND U1554 ( .A(n1459), .B(n26007), .Z(n1460) );
  AND U1555 ( .A(n26008), .B(n1460), .Z(n1461) );
  NANDN U1556 ( .A(n17736), .B(n1461), .Z(n1462) );
  ANDN U1557 ( .B(n1462), .A(n26010), .Z(n9662) );
  NAND U1558 ( .A(n9774), .B(n26172), .Z(n1463) );
  NAND U1559 ( .A(n1463), .B(n26175), .Z(n1464) );
  AND U1560 ( .A(n26176), .B(n1464), .Z(n1465) );
  OR U1561 ( .A(n26178), .B(n1465), .Z(n1466) );
  ANDN U1562 ( .B(n1466), .A(n17888), .Z(n1467) );
  NOR U1563 ( .A(n1467), .B(n26189), .Z(n1468) );
  OR U1564 ( .A(n26184), .B(n26182), .Z(n1469) );
  NAND U1565 ( .A(n1468), .B(n1469), .Z(n1470) );
  NOR U1566 ( .A(n11751), .B(n17892), .Z(n1471) );
  NAND U1567 ( .A(n1471), .B(n1470), .Z(n1472) );
  NAND U1568 ( .A(n1472), .B(n26193), .Z(n1473) );
  AND U1569 ( .A(n26198), .B(n11752), .Z(n1474) );
  XNOR U1570 ( .A(y[2917]), .B(x[2917]), .Z(n1475) );
  NANDN U1571 ( .A(n1473), .B(n1475), .Z(n1476) );
  AND U1572 ( .A(n1474), .B(n1476), .Z(n1477) );
  NOR U1573 ( .A(n1477), .B(n26201), .Z(n1478) );
  NANDN U1574 ( .A(n11750), .B(n1478), .Z(n1479) );
  NANDN U1575 ( .A(n26203), .B(n1479), .Z(n1480) );
  ANDN U1576 ( .B(n1480), .A(n26204), .Z(n9781) );
  NAND U1577 ( .A(n9833), .B(n9832), .Z(n1481) );
  AND U1578 ( .A(n26303), .B(n1481), .Z(n1482) );
  NANDN U1579 ( .A(n11726), .B(n1482), .Z(n1483) );
  ANDN U1580 ( .B(n26304), .A(n11725), .Z(n1484) );
  NAND U1581 ( .A(n1484), .B(n1483), .Z(n1485) );
  NAND U1582 ( .A(n1485), .B(n26306), .Z(n1486) );
  NAND U1583 ( .A(n1486), .B(n26308), .Z(n1487) );
  ANDN U1584 ( .B(n26312), .A(n11718), .Z(n1488) );
  NANDN U1585 ( .A(n26310), .B(n1487), .Z(n1489) );
  NAND U1586 ( .A(n1488), .B(n1489), .Z(n1490) );
  ANDN U1587 ( .B(n26314), .A(n18013), .Z(n1491) );
  NAND U1588 ( .A(n1491), .B(n1490), .Z(n1492) );
  NAND U1589 ( .A(n1492), .B(n26320), .Z(n1493) );
  ANDN U1590 ( .B(n26322), .A(n18014), .Z(n1494) );
  OR U1591 ( .A(n11719), .B(n1493), .Z(n1495) );
  AND U1592 ( .A(n1494), .B(n1495), .Z(n1496) );
  NANDN U1593 ( .A(n1496), .B(n26324), .Z(n1497) );
  NANDN U1594 ( .A(n26326), .B(n1497), .Z(n1498) );
  NANDN U1595 ( .A(n26329), .B(n1498), .Z(n9834) );
  NANDN U1596 ( .A(n9839), .B(n9838), .Z(n1499) );
  NAND U1597 ( .A(n1499), .B(n26396), .Z(n1500) );
  ANDN U1598 ( .B(n1500), .A(n26398), .Z(n1501) );
  ANDN U1599 ( .B(n26402), .A(n11698), .Z(n1502) );
  OR U1600 ( .A(n26401), .B(n1501), .Z(n1503) );
  AND U1601 ( .A(n1502), .B(n1503), .Z(n1504) );
  NOR U1602 ( .A(n1504), .B(n18102), .Z(n1505) );
  NAND U1603 ( .A(n1505), .B(n26404), .Z(n1506) );
  AND U1604 ( .A(n26410), .B(n1506), .Z(n1507) );
  ANDN U1605 ( .B(n26413), .A(n18103), .Z(n1508) );
  NANDN U1606 ( .A(n11697), .B(n1507), .Z(n1509) );
  NAND U1607 ( .A(n1508), .B(n1509), .Z(n1510) );
  NAND U1608 ( .A(n1510), .B(n26414), .Z(n1511) );
  NANDN U1609 ( .A(n26417), .B(n1511), .Z(n1512) );
  ANDN U1610 ( .B(n1512), .A(n26419), .Z(n1513) );
  NANDN U1611 ( .A(n18118), .B(n26422), .Z(n1514) );
  NOR U1612 ( .A(n1513), .B(n11691), .Z(n1515) );
  NAND U1613 ( .A(n1515), .B(n26420), .Z(n1516) );
  NANDN U1614 ( .A(n1514), .B(n1516), .Z(n9840) );
  ANDN U1615 ( .B(n9846), .A(n26489), .Z(n1517) );
  ANDN U1616 ( .B(n26492), .A(n11673), .Z(n1518) );
  OR U1617 ( .A(n26491), .B(n1517), .Z(n1519) );
  NAND U1618 ( .A(n1518), .B(n1519), .Z(n1520) );
  ANDN U1619 ( .B(n26494), .A(n18189), .Z(n1521) );
  NAND U1620 ( .A(n1521), .B(n1520), .Z(n1522) );
  NAND U1621 ( .A(n1522), .B(n26500), .Z(n1523) );
  NOR U1622 ( .A(n26503), .B(n18190), .Z(n1524) );
  OR U1623 ( .A(n11674), .B(n1523), .Z(n1525) );
  AND U1624 ( .A(n1524), .B(n1525), .Z(n1526) );
  OR U1625 ( .A(n26505), .B(n1526), .Z(n1527) );
  ANDN U1626 ( .B(n1527), .A(n26506), .Z(n1528) );
  ANDN U1627 ( .B(n26510), .A(n18209), .Z(n1529) );
  OR U1628 ( .A(n26509), .B(n1528), .Z(n1530) );
  AND U1629 ( .A(n1529), .B(n1530), .Z(n1531) );
  NOR U1630 ( .A(n1531), .B(n18212), .Z(n1532) );
  NAND U1631 ( .A(n1532), .B(n26512), .Z(n1533) );
  AND U1632 ( .A(n26518), .B(n1533), .Z(n1534) );
  ANDN U1633 ( .B(n1534), .A(n18210), .Z(n9850) );
  AND U1634 ( .A(n9874), .B(n11645), .Z(n1535) );
  NAND U1635 ( .A(n1535), .B(n26602), .Z(n1536) );
  AND U1636 ( .A(n18286), .B(n1536), .Z(n1537) );
  XNOR U1637 ( .A(x[3077]), .B(y[3077]), .Z(n1538) );
  NANDN U1638 ( .A(n11643), .B(n1538), .Z(n1539) );
  NAND U1639 ( .A(n1537), .B(n1539), .Z(n1540) );
  NAND U1640 ( .A(n1540), .B(n18285), .Z(n1541) );
  ANDN U1641 ( .B(n1541), .A(n18294), .Z(n1542) );
  XNOR U1642 ( .A(x[3078]), .B(n1540), .Z(n1543) );
  NAND U1643 ( .A(n1543), .B(y[3078]), .Z(n1544) );
  NAND U1644 ( .A(n1544), .B(n1542), .Z(n1545) );
  ANDN U1645 ( .B(n1545), .A(n18289), .Z(n1546) );
  XOR U1646 ( .A(y[3080]), .B(n18292), .Z(n1547) );
  NAND U1647 ( .A(n1547), .B(n1546), .Z(n1548) );
  NAND U1648 ( .A(y[3080]), .B(n18292), .Z(n1549) );
  AND U1649 ( .A(n1548), .B(n1549), .Z(n1550) );
  XNOR U1650 ( .A(x[3081]), .B(y[3081]), .Z(n1551) );
  NANDN U1651 ( .A(n1550), .B(n1551), .Z(n1552) );
  AND U1652 ( .A(n18297), .B(n1552), .Z(n9875) );
  NANDN U1653 ( .A(n15284), .B(n15280), .Z(n1553) );
  NANDN U1654 ( .A(n7579), .B(n1553), .Z(n1554) );
  AND U1655 ( .A(n7586), .B(n1554), .Z(n1555) );
  AND U1656 ( .A(n15287), .B(n1555), .Z(n23214) );
  NANDN U1657 ( .A(y[1711]), .B(x[1711]), .Z(n12319) );
  NANDN U1658 ( .A(x[1694]), .B(y[1694]), .Z(n1556) );
  NANDN U1659 ( .A(n15377), .B(n1556), .Z(n23287) );
  NOR U1660 ( .A(n18326), .B(n11620), .Z(n9919) );
  NANDN U1661 ( .A(x[1790]), .B(y[1790]), .Z(n12294) );
  NANDN U1662 ( .A(x[1859]), .B(y[1859]), .Z(n12256) );
  NANDN U1663 ( .A(x[1896]), .B(y[1896]), .Z(n1557) );
  NAND U1664 ( .A(n1557), .B(n15761), .Z(n23757) );
  NANDN U1665 ( .A(y[2059]), .B(x[2059]), .Z(n1558) );
  NAND U1666 ( .A(n1558), .B(n12188), .Z(n24141) );
  NANDN U1667 ( .A(y[2099]), .B(x[2099]), .Z(n1559) );
  NAND U1668 ( .A(n1559), .B(n12162), .Z(n24236) );
  NANDN U1669 ( .A(n16280), .B(n8513), .Z(n1560) );
  NAND U1670 ( .A(n1560), .B(n12147), .Z(n24359) );
  ANDN U1671 ( .B(n18694), .A(n18701), .Z(n1561) );
  NAND U1672 ( .A(n1561), .B(n10056), .Z(n1562) );
  AND U1673 ( .A(n10057), .B(n1562), .Z(n1563) );
  NANDN U1674 ( .A(n11339), .B(n1563), .Z(n1564) );
  ANDN U1675 ( .B(n27107), .A(n18700), .Z(n1565) );
  NAND U1676 ( .A(n1565), .B(n1564), .Z(n1566) );
  NANDN U1677 ( .A(n11338), .B(n1566), .Z(n1567) );
  NANDN U1678 ( .A(n1567), .B(n11337), .Z(n1568) );
  ANDN U1679 ( .B(n1568), .A(n27106), .Z(n1569) );
  NANDN U1680 ( .A(n18710), .B(n11336), .Z(n1570) );
  XNOR U1681 ( .A(y[3327]), .B(x[3327]), .Z(n1571) );
  NAND U1682 ( .A(n1571), .B(n1569), .Z(n1572) );
  NANDN U1683 ( .A(n1570), .B(n1572), .Z(n1573) );
  NOR U1684 ( .A(n18707), .B(n11334), .Z(n1574) );
  NAND U1685 ( .A(n1574), .B(n1573), .Z(n1575) );
  NANDN U1686 ( .A(n18711), .B(n1575), .Z(n1576) );
  XNOR U1687 ( .A(y[3330]), .B(x[3330]), .Z(n1577) );
  NAND U1688 ( .A(n1577), .B(n1576), .Z(n1578) );
  NAND U1689 ( .A(n1578), .B(n11332), .Z(n10058) );
  NANDN U1690 ( .A(n18756), .B(n10070), .Z(n1579) );
  ANDN U1691 ( .B(n1579), .A(n27176), .Z(n1580) );
  NANDN U1692 ( .A(n1580), .B(n18763), .Z(n1581) );
  XOR U1693 ( .A(n1580), .B(x[3359]), .Z(n1582) );
  NAND U1694 ( .A(n1582), .B(y[3359]), .Z(n1583) );
  NAND U1695 ( .A(n1581), .B(n1583), .Z(n1584) );
  NOR U1696 ( .A(n18764), .B(n11302), .Z(n1585) );
  NANDN U1697 ( .A(n18767), .B(n1584), .Z(n1586) );
  NAND U1698 ( .A(n1585), .B(n1586), .Z(n1587) );
  ANDN U1699 ( .B(n1587), .A(n18768), .Z(n1588) );
  XNOR U1700 ( .A(y[3362]), .B(x[3362]), .Z(n1589) );
  AND U1701 ( .A(n1588), .B(n1589), .Z(n1590) );
  NOR U1702 ( .A(n1590), .B(n11298), .Z(n1591) );
  NAND U1703 ( .A(n1591), .B(n11301), .Z(n1592) );
  ANDN U1704 ( .B(n1592), .A(n11300), .Z(n1593) );
  ANDN U1705 ( .B(n27195), .A(n11297), .Z(n1594) );
  NANDN U1706 ( .A(n18774), .B(n1593), .Z(n1595) );
  NAND U1707 ( .A(n1594), .B(n1595), .Z(n1596) );
  AND U1708 ( .A(n18777), .B(n1596), .Z(n10071) );
  NANDN U1709 ( .A(n11270), .B(n11271), .Z(n1597) );
  NAND U1710 ( .A(n10097), .B(n27230), .Z(n1598) );
  NANDN U1711 ( .A(n11275), .B(n1598), .Z(n1599) );
  NAND U1712 ( .A(n1599), .B(n11273), .Z(n1600) );
  ANDN U1713 ( .B(n1600), .A(n11272), .Z(n1601) );
  XNOR U1714 ( .A(x[3384]), .B(n1599), .Z(n1602) );
  NAND U1715 ( .A(n1602), .B(y[3384]), .Z(n1603) );
  NAND U1716 ( .A(n1603), .B(n1601), .Z(n1604) );
  ANDN U1717 ( .B(n1604), .A(n18805), .Z(n1605) );
  XNOR U1718 ( .A(y[3386]), .B(x[3386]), .Z(n1606) );
  AND U1719 ( .A(n1605), .B(n1606), .Z(n1607) );
  NOR U1720 ( .A(n18814), .B(n18809), .Z(n1608) );
  OR U1721 ( .A(n1597), .B(n1607), .Z(n1609) );
  AND U1722 ( .A(n1608), .B(n1609), .Z(n1610) );
  NOR U1723 ( .A(n1610), .B(n11269), .Z(n1611) );
  NAND U1724 ( .A(n1611), .B(n27245), .Z(n1612) );
  ANDN U1725 ( .B(n1612), .A(n18813), .Z(n1613) );
  XNOR U1726 ( .A(y[3390]), .B(x[3390]), .Z(n1614) );
  NAND U1727 ( .A(n1613), .B(n1614), .Z(n10098) );
  NANDN U1728 ( .A(n16728), .B(n8853), .Z(n1615) );
  NAND U1729 ( .A(n1615), .B(n12053), .Z(n24844) );
  NANDN U1730 ( .A(x[2391]), .B(y[2391]), .Z(n12040) );
  NANDN U1731 ( .A(x[2456]), .B(y[2456]), .Z(n1616) );
  AND U1732 ( .A(n12011), .B(n1616), .Z(n25073) );
  NANDN U1733 ( .A(n10140), .B(y[3480]), .Z(n1617) );
  ANDN U1734 ( .B(n1617), .A(n11170), .Z(n1618) );
  XNOR U1735 ( .A(y[3480]), .B(n10140), .Z(n1619) );
  NAND U1736 ( .A(n1619), .B(n18995), .Z(n1620) );
  NAND U1737 ( .A(n1618), .B(n1620), .Z(n1621) );
  ANDN U1738 ( .B(n1621), .A(n18999), .Z(n1622) );
  NANDN U1739 ( .A(x[3482]), .B(n1622), .Z(n1623) );
  ANDN U1740 ( .B(n1623), .A(n11168), .Z(n1624) );
  XNOR U1741 ( .A(n1622), .B(x[3482]), .Z(n1625) );
  NAND U1742 ( .A(n1625), .B(y[3482]), .Z(n1626) );
  NAND U1743 ( .A(n1624), .B(n1626), .Z(n1627) );
  ANDN U1744 ( .B(n1627), .A(n19003), .Z(n1628) );
  NAND U1745 ( .A(n11166), .B(y[3484]), .Z(n1629) );
  ANDN U1746 ( .B(n1629), .A(n11165), .Z(n1630) );
  XOR U1747 ( .A(y[3484]), .B(n11166), .Z(n1631) );
  NAND U1748 ( .A(n1631), .B(n1628), .Z(n1632) );
  NAND U1749 ( .A(n1630), .B(n1632), .Z(n1633) );
  NAND U1750 ( .A(n1633), .B(n19008), .Z(n10141) );
  NANDN U1751 ( .A(x[2584]), .B(y[2584]), .Z(n1634) );
  NAND U1752 ( .A(n1634), .B(n11953), .Z(n25373) );
  ANDN U1753 ( .B(n10151), .A(n11146), .Z(n1635) );
  NAND U1754 ( .A(n1635), .B(n11142), .Z(n1636) );
  ANDN U1755 ( .B(n1636), .A(n11145), .Z(n1637) );
  NANDN U1756 ( .A(n11140), .B(n11143), .Z(n1638) );
  XNOR U1757 ( .A(y[3505]), .B(x[3505]), .Z(n1639) );
  NAND U1758 ( .A(n1639), .B(n1637), .Z(n1640) );
  NANDN U1759 ( .A(n1638), .B(n1640), .Z(n1641) );
  NOR U1760 ( .A(n19041), .B(n19037), .Z(n1642) );
  NAND U1761 ( .A(n1642), .B(n1641), .Z(n1643) );
  ANDN U1762 ( .B(n1643), .A(n11141), .Z(n1644) );
  NANDN U1763 ( .A(n19044), .B(n1644), .Z(n1645) );
  NOR U1764 ( .A(n11139), .B(n19042), .Z(n1646) );
  NAND U1765 ( .A(n1646), .B(n1645), .Z(n1647) );
  NAND U1766 ( .A(n1647), .B(n19045), .Z(n1648) );
  NANDN U1767 ( .A(y[3510]), .B(x[3510]), .Z(n1649) );
  XNOR U1768 ( .A(y[3510]), .B(x[3510]), .Z(n1650) );
  NAND U1769 ( .A(n1650), .B(n1648), .Z(n1651) );
  NAND U1770 ( .A(n1649), .B(n1651), .Z(n10152) );
  NOR U1771 ( .A(n27522), .B(n19082), .Z(n1652) );
  NAND U1772 ( .A(n1652), .B(n10154), .Z(n1653) );
  ANDN U1773 ( .B(n1653), .A(n19077), .Z(n1654) );
  NAND U1774 ( .A(y[3526]), .B(n19080), .Z(n1655) );
  ANDN U1775 ( .B(n1655), .A(n11122), .Z(n1656) );
  XOR U1776 ( .A(n19080), .B(y[3526]), .Z(n1657) );
  NAND U1777 ( .A(n1657), .B(n1654), .Z(n1658) );
  NAND U1778 ( .A(n1656), .B(n1658), .Z(n1659) );
  ANDN U1779 ( .B(n1659), .A(n19084), .Z(n1660) );
  OR U1780 ( .A(y[3528]), .B(n1660), .Z(n1661) );
  XOR U1781 ( .A(n1660), .B(y[3528]), .Z(n1662) );
  NAND U1782 ( .A(n1662), .B(x[3528]), .Z(n1663) );
  NAND U1783 ( .A(n1661), .B(n1663), .Z(n1664) );
  ANDN U1784 ( .B(n1664), .A(n11118), .Z(n1665) );
  NOR U1785 ( .A(n1665), .B(n11120), .Z(n1666) );
  NAND U1786 ( .A(n1666), .B(n19090), .Z(n1667) );
  AND U1787 ( .A(n27541), .B(n1667), .Z(n1668) );
  NANDN U1788 ( .A(n11117), .B(n1668), .Z(n10155) );
  ANDN U1789 ( .B(n10158), .A(n19123), .Z(n1669) );
  NAND U1790 ( .A(y[3546]), .B(n11102), .Z(n1670) );
  ANDN U1791 ( .B(n1670), .A(n11099), .Z(n1671) );
  XOR U1792 ( .A(n11102), .B(y[3546]), .Z(n1672) );
  NAND U1793 ( .A(n1672), .B(n1669), .Z(n1673) );
  NAND U1794 ( .A(n1671), .B(n1673), .Z(n1674) );
  ANDN U1795 ( .B(n1674), .A(n11100), .Z(n1675) );
  NANDN U1796 ( .A(x[3548]), .B(n1675), .Z(n1676) );
  ANDN U1797 ( .B(n1676), .A(n11095), .Z(n1677) );
  XNOR U1798 ( .A(n1675), .B(x[3548]), .Z(n1678) );
  NAND U1799 ( .A(n1678), .B(y[3548]), .Z(n1679) );
  NAND U1800 ( .A(n1677), .B(n1679), .Z(n1680) );
  AND U1801 ( .A(n11097), .B(n1680), .Z(n1681) );
  NANDN U1802 ( .A(x[3550]), .B(n1681), .Z(n1682) );
  ANDN U1803 ( .B(n1682), .A(n11092), .Z(n1683) );
  XNOR U1804 ( .A(n1681), .B(x[3550]), .Z(n1684) );
  NAND U1805 ( .A(n1684), .B(y[3550]), .Z(n1685) );
  NAND U1806 ( .A(n1683), .B(n1685), .Z(n10159) );
  NAND U1807 ( .A(n11073), .B(n10163), .Z(n1686) );
  NANDN U1808 ( .A(n10164), .B(x[3567]), .Z(n1687) );
  NAND U1809 ( .A(n1686), .B(n1687), .Z(n1688) );
  OR U1810 ( .A(n11072), .B(n1688), .Z(n1689) );
  AND U1811 ( .A(n19165), .B(n1689), .Z(n1690) );
  NANDN U1812 ( .A(y[3569]), .B(x[3569]), .Z(n1691) );
  ANDN U1813 ( .B(n1691), .A(n11068), .Z(n1692) );
  XNOR U1814 ( .A(x[3569]), .B(y[3569]), .Z(n1693) );
  NAND U1815 ( .A(n1693), .B(n1690), .Z(n1694) );
  NAND U1816 ( .A(n1692), .B(n1694), .Z(n1695) );
  ANDN U1817 ( .B(n27628), .A(n11070), .Z(n1696) );
  NAND U1818 ( .A(n1696), .B(n1695), .Z(n1697) );
  NANDN U1819 ( .A(n11067), .B(n1697), .Z(n1698) );
  ANDN U1820 ( .B(n27626), .A(n19174), .Z(n1699) );
  NANDN U1821 ( .A(n1698), .B(n11066), .Z(n1700) );
  AND U1822 ( .A(n1699), .B(n1700), .Z(n1701) );
  NOR U1823 ( .A(n1701), .B(n19176), .Z(n1702) );
  NANDN U1824 ( .A(n11065), .B(n1702), .Z(n1703) );
  ANDN U1825 ( .B(n1703), .A(n19173), .Z(n10165) );
  ANDN U1826 ( .B(n10172), .A(n19209), .Z(n1704) );
  NANDN U1827 ( .A(x[3592]), .B(n10170), .Z(n1705) );
  NAND U1828 ( .A(n1704), .B(n1705), .Z(n1706) );
  ANDN U1829 ( .B(n1706), .A(n19204), .Z(n1707) );
  NAND U1830 ( .A(n19207), .B(y[3594]), .Z(n1708) );
  ANDN U1831 ( .B(n1708), .A(n11035), .Z(n1709) );
  XOR U1832 ( .A(y[3594]), .B(n19207), .Z(n1710) );
  NAND U1833 ( .A(n1710), .B(n1707), .Z(n1711) );
  NAND U1834 ( .A(n1709), .B(n1711), .Z(n1712) );
  NOR U1835 ( .A(n19214), .B(n11037), .Z(n1713) );
  NAND U1836 ( .A(n1713), .B(n1712), .Z(n1714) );
  NANDN U1837 ( .A(n27687), .B(n1714), .Z(n1715) );
  NOR U1838 ( .A(n11033), .B(n19213), .Z(n1716) );
  OR U1839 ( .A(n11034), .B(n1715), .Z(n1717) );
  AND U1840 ( .A(n1716), .B(n1717), .Z(n1718) );
  NOR U1841 ( .A(n1718), .B(n27684), .Z(n1719) );
  NAND U1842 ( .A(n1719), .B(n27692), .Z(n1720) );
  AND U1843 ( .A(n19220), .B(n1720), .Z(n10173) );
  ANDN U1844 ( .B(n10178), .A(n11013), .Z(n1721) );
  NANDN U1845 ( .A(y[3615]), .B(n10176), .Z(n1722) );
  NAND U1846 ( .A(n1721), .B(n1722), .Z(n1723) );
  ANDN U1847 ( .B(n1723), .A(n19252), .Z(n1724) );
  NAND U1848 ( .A(n11012), .B(x[3617]), .Z(n1725) );
  ANDN U1849 ( .B(n1725), .A(n19258), .Z(n1726) );
  XOR U1850 ( .A(x[3617]), .B(n11012), .Z(n1727) );
  NAND U1851 ( .A(n1727), .B(n1724), .Z(n1728) );
  NAND U1852 ( .A(n1726), .B(n1728), .Z(n1729) );
  ANDN U1853 ( .B(n27737), .A(n11011), .Z(n1730) );
  NAND U1854 ( .A(n1730), .B(n1729), .Z(n1731) );
  NANDN U1855 ( .A(n19257), .B(n1731), .Z(n1732) );
  ANDN U1856 ( .B(n27736), .A(n19264), .Z(n1733) );
  NANDN U1857 ( .A(n1732), .B(n19261), .Z(n1734) );
  AND U1858 ( .A(n1733), .B(n1734), .Z(n1735) );
  NOR U1859 ( .A(n11009), .B(n19267), .Z(n1736) );
  NANDN U1860 ( .A(n1735), .B(n1736), .Z(n1737) );
  ANDN U1861 ( .B(n1737), .A(n19265), .Z(n10179) );
  ANDN U1862 ( .B(n10185), .A(n10991), .Z(n1738) );
  NANDN U1863 ( .A(y[3639]), .B(n10183), .Z(n1739) );
  NAND U1864 ( .A(n1738), .B(n1739), .Z(n1740) );
  ANDN U1865 ( .B(n1740), .A(n19303), .Z(n1741) );
  NANDN U1866 ( .A(y[3641]), .B(n1741), .Z(n1742) );
  ANDN U1867 ( .B(n1742), .A(n10987), .Z(n1743) );
  XNOR U1868 ( .A(n1741), .B(y[3641]), .Z(n1744) );
  NAND U1869 ( .A(n1744), .B(x[3641]), .Z(n1745) );
  NAND U1870 ( .A(n1743), .B(n1745), .Z(n1746) );
  ANDN U1871 ( .B(n27789), .A(n10989), .Z(n1747) );
  NAND U1872 ( .A(n1747), .B(n1746), .Z(n1748) );
  NANDN U1873 ( .A(n10986), .B(n1748), .Z(n1749) );
  ANDN U1874 ( .B(n27788), .A(n19313), .Z(n1750) );
  NANDN U1875 ( .A(n1749), .B(n19309), .Z(n1751) );
  AND U1876 ( .A(n1750), .B(n1751), .Z(n1752) );
  NOR U1877 ( .A(n1752), .B(n19316), .Z(n1753) );
  NANDN U1878 ( .A(n10985), .B(n1753), .Z(n1754) );
  ANDN U1879 ( .B(n1754), .A(n19314), .Z(n10186) );
  NOR U1880 ( .A(n19332), .B(n10975), .Z(n10187) );
  NANDN U1881 ( .A(n10952), .B(n10209), .Z(n1755) );
  AND U1882 ( .A(n10954), .B(n1755), .Z(n1756) );
  NANDN U1883 ( .A(x[3674]), .B(y[3674]), .Z(n1757) );
  ANDN U1884 ( .B(n1757), .A(n19372), .Z(n1758) );
  XNOR U1885 ( .A(y[3674]), .B(x[3674]), .Z(n1759) );
  NAND U1886 ( .A(n1759), .B(n1756), .Z(n1760) );
  NAND U1887 ( .A(n1758), .B(n1760), .Z(n1761) );
  ANDN U1888 ( .B(n1761), .A(n19367), .Z(n1762) );
  NAND U1889 ( .A(n19370), .B(y[3676]), .Z(n1763) );
  ANDN U1890 ( .B(n1763), .A(n10950), .Z(n1764) );
  XOR U1891 ( .A(y[3676]), .B(n19370), .Z(n1765) );
  NAND U1892 ( .A(n1765), .B(n1762), .Z(n1766) );
  NAND U1893 ( .A(n1764), .B(n1766), .Z(n1767) );
  NANDN U1894 ( .A(n19374), .B(n1767), .Z(n1768) );
  NANDN U1895 ( .A(y[3678]), .B(x[3678]), .Z(n1769) );
  XNOR U1896 ( .A(y[3678]), .B(x[3678]), .Z(n1770) );
  NAND U1897 ( .A(n1770), .B(n1768), .Z(n1771) );
  NAND U1898 ( .A(n1769), .B(n1771), .Z(n10210) );
  NANDN U1899 ( .A(n10934), .B(n10212), .Z(n1772) );
  AND U1900 ( .A(n19404), .B(n1772), .Z(n1773) );
  NANDN U1901 ( .A(x[3692]), .B(y[3692]), .Z(n1774) );
  ANDN U1902 ( .B(n1774), .A(n10930), .Z(n1775) );
  XNOR U1903 ( .A(y[3692]), .B(x[3692]), .Z(n1776) );
  NAND U1904 ( .A(n1776), .B(n1773), .Z(n1777) );
  NAND U1905 ( .A(n1775), .B(n1777), .Z(n1778) );
  AND U1906 ( .A(n10932), .B(n1778), .Z(n1779) );
  NANDN U1907 ( .A(x[3694]), .B(n1779), .Z(n1780) );
  ANDN U1908 ( .B(n1780), .A(n10928), .Z(n1781) );
  XNOR U1909 ( .A(n1779), .B(x[3694]), .Z(n1782) );
  NAND U1910 ( .A(n1782), .B(y[3694]), .Z(n1783) );
  NAND U1911 ( .A(n1781), .B(n1783), .Z(n1784) );
  ANDN U1912 ( .B(n1784), .A(n19409), .Z(n1785) );
  OR U1913 ( .A(y[3696]), .B(n1785), .Z(n1786) );
  XOR U1914 ( .A(n1785), .B(y[3696]), .Z(n1787) );
  NAND U1915 ( .A(n1787), .B(x[3696]), .Z(n1788) );
  NAND U1916 ( .A(n1786), .B(n1788), .Z(n1789) );
  ANDN U1917 ( .B(n1789), .A(n10926), .Z(n10214) );
  NANDN U1918 ( .A(x[3083]), .B(y[3083]), .Z(n11637) );
  NOR U1919 ( .A(n27936), .B(n19462), .Z(n1790) );
  OR U1920 ( .A(n10216), .B(n10217), .Z(n1791) );
  NAND U1921 ( .A(n1790), .B(n1791), .Z(n1792) );
  ANDN U1922 ( .B(n1792), .A(n19457), .Z(n1793) );
  NAND U1923 ( .A(n19460), .B(y[3714]), .Z(n1794) );
  ANDN U1924 ( .B(n1794), .A(n10919), .Z(n1795) );
  XOR U1925 ( .A(y[3714]), .B(n19460), .Z(n1796) );
  NAND U1926 ( .A(n1796), .B(n1793), .Z(n1797) );
  NAND U1927 ( .A(n1795), .B(n1797), .Z(n1798) );
  NANDN U1928 ( .A(n19464), .B(n1798), .Z(n1799) );
  NANDN U1929 ( .A(y[3716]), .B(x[3716]), .Z(n1800) );
  XNOR U1930 ( .A(y[3716]), .B(x[3716]), .Z(n1801) );
  NAND U1931 ( .A(n1801), .B(n1799), .Z(n1802) );
  NAND U1932 ( .A(n1800), .B(n1802), .Z(n1803) );
  NOR U1933 ( .A(n10917), .B(n19471), .Z(n1804) );
  NANDN U1934 ( .A(n10915), .B(n1803), .Z(n1805) );
  NAND U1935 ( .A(n1804), .B(n1805), .Z(n10218) );
  NANDN U1936 ( .A(y[3112]), .B(x[3112]), .Z(n11596) );
  NANDN U1937 ( .A(y[3116]), .B(x[3116]), .Z(n11588) );
  NANDN U1938 ( .A(y[3124]), .B(x[3124]), .Z(n11576) );
  NANDN U1939 ( .A(y[3142]), .B(x[3142]), .Z(n11557) );
  NANDN U1940 ( .A(x[3161]), .B(y[3161]), .Z(n11543) );
  ANDN U1941 ( .B(n10220), .A(n10898), .Z(n1806) );
  NAND U1942 ( .A(y[3734]), .B(n10895), .Z(n1807) );
  ANDN U1943 ( .B(n1807), .A(n10894), .Z(n1808) );
  XOR U1944 ( .A(n10895), .B(y[3734]), .Z(n1809) );
  NAND U1945 ( .A(n1809), .B(n1806), .Z(n1810) );
  NAND U1946 ( .A(n1808), .B(n1810), .Z(n1811) );
  AND U1947 ( .A(n19502), .B(n1811), .Z(n1812) );
  OR U1948 ( .A(y[3736]), .B(n1812), .Z(n1813) );
  XOR U1949 ( .A(n1812), .B(y[3736]), .Z(n1814) );
  NAND U1950 ( .A(n1814), .B(x[3736]), .Z(n1815) );
  NAND U1951 ( .A(n1813), .B(n1815), .Z(n1816) );
  ANDN U1952 ( .B(n1816), .A(n10890), .Z(n1817) );
  NOR U1953 ( .A(n1817), .B(n10892), .Z(n1818) );
  NAND U1954 ( .A(n1818), .B(n19507), .Z(n1819) );
  ANDN U1955 ( .B(n1819), .A(n20220), .Z(n1820) );
  NOR U1956 ( .A(n19508), .B(n19510), .Z(n1821) );
  NANDN U1957 ( .A(n10889), .B(n1820), .Z(n1822) );
  NAND U1958 ( .A(n1821), .B(n1822), .Z(n1823) );
  ANDN U1959 ( .B(n1823), .A(n20221), .Z(n10221) );
  NANDN U1960 ( .A(y[3178]), .B(x[3178]), .Z(n11523) );
  NANDN U1961 ( .A(y[3190]), .B(x[3190]), .Z(n11507) );
  NANDN U1962 ( .A(y[3194]), .B(x[3194]), .Z(n11503) );
  NANDN U1963 ( .A(y[3202]), .B(x[3202]), .Z(n18494) );
  NANDN U1964 ( .A(y[3210]), .B(x[3210]), .Z(n11481) );
  NANDN U1965 ( .A(y[3218]), .B(x[3218]), .Z(n11471) );
  NAND U1966 ( .A(n10224), .B(n10225), .Z(n1824) );
  NANDN U1967 ( .A(n1824), .B(x[3757]), .Z(n1825) );
  ANDN U1968 ( .B(n1825), .A(n10873), .Z(n1826) );
  XNOR U1969 ( .A(n1824), .B(x[3757]), .Z(n1827) );
  NAND U1970 ( .A(n1827), .B(n10874), .Z(n1828) );
  NAND U1971 ( .A(n1826), .B(n1828), .Z(n1829) );
  ANDN U1972 ( .B(n1829), .A(n19551), .Z(n1830) );
  NAND U1973 ( .A(n10871), .B(x[3759]), .Z(n1831) );
  ANDN U1974 ( .B(n1831), .A(n10868), .Z(n1832) );
  XOR U1975 ( .A(x[3759]), .B(n10871), .Z(n1833) );
  NAND U1976 ( .A(n1833), .B(n1830), .Z(n1834) );
  NAND U1977 ( .A(n1832), .B(n1834), .Z(n1835) );
  ANDN U1978 ( .B(n1835), .A(n10869), .Z(n1836) );
  NANDN U1979 ( .A(y[3761]), .B(n1836), .Z(n1837) );
  ANDN U1980 ( .B(n1837), .A(n10866), .Z(n1838) );
  XNOR U1981 ( .A(n1836), .B(y[3761]), .Z(n1839) );
  NAND U1982 ( .A(n1839), .B(x[3761]), .Z(n1840) );
  NAND U1983 ( .A(n1838), .B(n1840), .Z(n10227) );
  NANDN U1984 ( .A(y[3230]), .B(x[3230]), .Z(n11455) );
  NANDN U1985 ( .A(y[3234]), .B(x[3234]), .Z(n11451) );
  NANDN U1986 ( .A(y[3250]), .B(x[3250]), .Z(n11429) );
  NANDN U1987 ( .A(y[3254]), .B(x[3254]), .Z(n11425) );
  NANDN U1988 ( .A(x[3281]), .B(y[3281]), .Z(n11398) );
  AND U1989 ( .A(n10230), .B(n10231), .Z(n1841) );
  NANDN U1990 ( .A(x[3780]), .B(n1841), .Z(n1842) );
  ANDN U1991 ( .B(n1842), .A(n10848), .Z(n1843) );
  XNOR U1992 ( .A(n1841), .B(x[3780]), .Z(n1844) );
  NAND U1993 ( .A(n1844), .B(y[3780]), .Z(n1845) );
  NAND U1994 ( .A(n1843), .B(n1845), .Z(n1846) );
  ANDN U1995 ( .B(n1846), .A(n19597), .Z(n1847) );
  NAND U1996 ( .A(n10847), .B(y[3782]), .Z(n1848) );
  ANDN U1997 ( .B(n1848), .A(n19606), .Z(n1849) );
  XOR U1998 ( .A(y[3782]), .B(n10847), .Z(n1850) );
  NAND U1999 ( .A(n1850), .B(n1847), .Z(n1851) );
  NAND U2000 ( .A(n1849), .B(n1851), .Z(n1852) );
  NANDN U2001 ( .A(n19601), .B(n1852), .Z(n1853) );
  NANDN U2002 ( .A(n1853), .B(y[3784]), .Z(n1854) );
  ANDN U2003 ( .B(n1854), .A(n10846), .Z(n1855) );
  XNOR U2004 ( .A(y[3784]), .B(n1853), .Z(n1856) );
  NAND U2005 ( .A(n1856), .B(n19604), .Z(n1857) );
  NAND U2006 ( .A(n1855), .B(n1857), .Z(n10232) );
  NANDN U2007 ( .A(x[3287]), .B(y[3287]), .Z(n18639) );
  NANDN U2008 ( .A(x[3293]), .B(y[3293]), .Z(n11381) );
  NANDN U2009 ( .A(x[3299]), .B(y[3299]), .Z(n11373) );
  NANDN U2010 ( .A(x[3307]), .B(y[3307]), .Z(n18669) );
  NANDN U2011 ( .A(x[3311]), .B(y[3311]), .Z(n11352) );
  NAND U2012 ( .A(n10828), .B(n10235), .Z(n1858) );
  NANDN U2013 ( .A(n10236), .B(y[3800]), .Z(n1859) );
  NAND U2014 ( .A(n1858), .B(n1859), .Z(n1860) );
  OR U2015 ( .A(n10827), .B(n1860), .Z(n1861) );
  ANDN U2016 ( .B(n1861), .A(n19639), .Z(n1862) );
  NAND U2017 ( .A(n10825), .B(y[3802]), .Z(n1863) );
  ANDN U2018 ( .B(n1863), .A(n10822), .Z(n1864) );
  XOR U2019 ( .A(y[3802]), .B(n10825), .Z(n1865) );
  NAND U2020 ( .A(n1865), .B(n1862), .Z(n1866) );
  NAND U2021 ( .A(n1864), .B(n1866), .Z(n1867) );
  ANDN U2022 ( .B(n1867), .A(n10823), .Z(n1868) );
  NANDN U2023 ( .A(x[3804]), .B(n1868), .Z(n1869) );
  ANDN U2024 ( .B(n1869), .A(n10820), .Z(n1870) );
  XNOR U2025 ( .A(n1868), .B(x[3804]), .Z(n1871) );
  NAND U2026 ( .A(n1871), .B(y[3804]), .Z(n1872) );
  NAND U2027 ( .A(n1870), .B(n1872), .Z(n1873) );
  NANDN U2028 ( .A(n19645), .B(n1873), .Z(n10237) );
  NANDN U2029 ( .A(x[3345]), .B(y[3345]), .Z(n11315) );
  NANDN U2030 ( .A(y[3402]), .B(x[3402]), .Z(n18839) );
  NANDN U2031 ( .A(x[3421]), .B(y[3421]), .Z(n11227) );
  NANDN U2032 ( .A(n10784), .B(n19698), .Z(n1874) );
  XNOR U2033 ( .A(y[3835]), .B(x[3835]), .Z(n1875) );
  AND U2034 ( .A(n10271), .B(n1875), .Z(n1876) );
  NOR U2035 ( .A(n19700), .B(n19704), .Z(n1877) );
  OR U2036 ( .A(n1874), .B(n1876), .Z(n1878) );
  AND U2037 ( .A(n1877), .B(n1878), .Z(n1879) );
  NOR U2038 ( .A(n1879), .B(n10785), .Z(n1880) );
  NANDN U2039 ( .A(n19707), .B(n1880), .Z(n1881) );
  NANDN U2040 ( .A(n19705), .B(n1881), .Z(n1882) );
  OR U2041 ( .A(n19712), .B(n1882), .Z(n1883) );
  NAND U2042 ( .A(n1883), .B(n19708), .Z(n1884) );
  NANDN U2043 ( .A(n1884), .B(y[3840]), .Z(n1885) );
  ANDN U2044 ( .B(n1885), .A(n10783), .Z(n1886) );
  XNOR U2045 ( .A(n1884), .B(y[3840]), .Z(n1887) );
  NAND U2046 ( .A(n1887), .B(n19710), .Z(n1888) );
  NAND U2047 ( .A(n1886), .B(n1888), .Z(n1889) );
  NANDN U2048 ( .A(n19714), .B(n1889), .Z(n10272) );
  NANDN U2049 ( .A(x[3443]), .B(y[3443]), .Z(n18917) );
  NANDN U2050 ( .A(x[3451]), .B(y[3451]), .Z(n11195) );
  NANDN U2051 ( .A(x[3459]), .B(y[3459]), .Z(n11189) );
  NAND U2052 ( .A(n10296), .B(n10758), .Z(n1890) );
  NANDN U2053 ( .A(n10297), .B(y[3858]), .Z(n1891) );
  NAND U2054 ( .A(n1890), .B(n1891), .Z(n1892) );
  NOR U2055 ( .A(n19743), .B(n10756), .Z(n1893) );
  OR U2056 ( .A(n10755), .B(n1892), .Z(n1894) );
  AND U2057 ( .A(n1893), .B(n1894), .Z(n1895) );
  NOR U2058 ( .A(n19742), .B(n10753), .Z(n1896) );
  NOR U2059 ( .A(n28267), .B(n10754), .Z(n1897) );
  NANDN U2060 ( .A(n1895), .B(n1897), .Z(n1898) );
  AND U2061 ( .A(n1896), .B(n1898), .Z(n1899) );
  NOR U2062 ( .A(n10750), .B(n28264), .Z(n1900) );
  NANDN U2063 ( .A(n1899), .B(n1900), .Z(n1901) );
  ANDN U2064 ( .B(n1901), .A(n10751), .Z(n1902) );
  NAND U2065 ( .A(y[3864]), .B(n10748), .Z(n1903) );
  ANDN U2066 ( .B(n1903), .A(n10745), .Z(n1904) );
  XOR U2067 ( .A(n10748), .B(y[3864]), .Z(n1905) );
  NAND U2068 ( .A(n1905), .B(n1902), .Z(n1906) );
  NAND U2069 ( .A(n1904), .B(n1906), .Z(n10298) );
  ANDN U2070 ( .B(n10302), .A(n19774), .Z(n1907) );
  NAND U2071 ( .A(y[3878]), .B(n10731), .Z(n1908) );
  ANDN U2072 ( .B(n1908), .A(n19781), .Z(n1909) );
  XOR U2073 ( .A(n10731), .B(y[3878]), .Z(n1910) );
  NAND U2074 ( .A(n1910), .B(n1907), .Z(n1911) );
  NAND U2075 ( .A(n1909), .B(n1911), .Z(n1912) );
  ANDN U2076 ( .B(n1912), .A(n19778), .Z(n1913) );
  NANDN U2077 ( .A(x[3880]), .B(n1913), .Z(n1914) );
  ANDN U2078 ( .B(n1914), .A(n10729), .Z(n1915) );
  XNOR U2079 ( .A(n1913), .B(x[3880]), .Z(n1916) );
  NAND U2080 ( .A(n1916), .B(y[3880]), .Z(n1917) );
  NAND U2081 ( .A(n1915), .B(n1917), .Z(n1918) );
  NANDN U2082 ( .A(n19784), .B(n1918), .Z(n1919) );
  NANDN U2083 ( .A(y[3882]), .B(x[3882]), .Z(n1920) );
  XNOR U2084 ( .A(y[3882]), .B(x[3882]), .Z(n1921) );
  NAND U2085 ( .A(n1921), .B(n1919), .Z(n1922) );
  NAND U2086 ( .A(n1920), .B(n1922), .Z(n10303) );
  NOR U2087 ( .A(n10326), .B(n19828), .Z(n1923) );
  NAND U2088 ( .A(n1923), .B(n10327), .Z(n1924) );
  NAND U2089 ( .A(n1924), .B(n28371), .Z(n1925) );
  XNOR U2090 ( .A(x[3910]), .B(y[3910]), .Z(n1926) );
  ANDN U2091 ( .B(n1926), .A(n10690), .Z(n1927) );
  OR U2092 ( .A(n20208), .B(n1925), .Z(n1928) );
  NAND U2093 ( .A(n1928), .B(n1927), .Z(n1929) );
  NANDN U2094 ( .A(n28370), .B(n1929), .Z(n1930) );
  NOR U2095 ( .A(n19840), .B(n10689), .Z(n1931) );
  OR U2096 ( .A(n10687), .B(n1930), .Z(n1932) );
  AND U2097 ( .A(n1931), .B(n1932), .Z(n1933) );
  NOR U2098 ( .A(n20206), .B(n10686), .Z(n1934) );
  NANDN U2099 ( .A(n1933), .B(n1934), .Z(n1935) );
  ANDN U2100 ( .B(n1935), .A(n10685), .Z(n1936) );
  NOR U2101 ( .A(n19849), .B(n20207), .Z(n1937) );
  NANDN U2102 ( .A(n19839), .B(n1936), .Z(n1938) );
  NAND U2103 ( .A(n1937), .B(n1938), .Z(n1939) );
  NANDN U2104 ( .A(n19844), .B(n1939), .Z(n10329) );
  ANDN U2105 ( .B(n10334), .A(n19871), .Z(n1940) );
  NANDN U2106 ( .A(x[3924]), .B(n10332), .Z(n1941) );
  AND U2107 ( .A(n1940), .B(n1941), .Z(n1942) );
  NOR U2108 ( .A(n10677), .B(n19874), .Z(n1943) );
  NANDN U2109 ( .A(n1942), .B(n1943), .Z(n1944) );
  ANDN U2110 ( .B(n1944), .A(n28409), .Z(n1945) );
  NOR U2111 ( .A(n10675), .B(n19873), .Z(n1946) );
  NANDN U2112 ( .A(n19870), .B(n1945), .Z(n1947) );
  NAND U2113 ( .A(n1946), .B(n1947), .Z(n1948) );
  ANDN U2114 ( .B(n1948), .A(n28408), .Z(n1949) );
  NOR U2115 ( .A(n19878), .B(n10672), .Z(n1950) );
  NANDN U2116 ( .A(n10674), .B(n1949), .Z(n1951) );
  NAND U2117 ( .A(n1950), .B(n1951), .Z(n1952) );
  ANDN U2118 ( .B(n10673), .A(n20203), .Z(n1953) );
  NAND U2119 ( .A(n1953), .B(n1952), .Z(n1954) );
  NANDN U2120 ( .A(n10670), .B(n1954), .Z(n1955) );
  OR U2121 ( .A(n10671), .B(n1955), .Z(n1956) );
  ANDN U2122 ( .B(n1956), .A(n19887), .Z(n10335) );
  ANDN U2123 ( .B(n28478), .A(n28486), .Z(n1957) );
  NAND U2124 ( .A(n1957), .B(n10359), .Z(n1958) );
  ANDN U2125 ( .B(n1958), .A(n10633), .Z(n1959) );
  NOR U2126 ( .A(n10630), .B(n28484), .Z(n1960) );
  NANDN U2127 ( .A(n10635), .B(n1959), .Z(n1961) );
  NAND U2128 ( .A(n1960), .B(n1961), .Z(n1962) );
  NANDN U2129 ( .A(n19940), .B(n10629), .Z(n1963) );
  NOR U2130 ( .A(n10627), .B(n10632), .Z(n1964) );
  NAND U2131 ( .A(n1964), .B(n1962), .Z(n1965) );
  NANDN U2132 ( .A(n1963), .B(n1965), .Z(n1966) );
  NOR U2133 ( .A(n19942), .B(n10628), .Z(n1967) );
  NAND U2134 ( .A(n1967), .B(n1966), .Z(n1968) );
  AND U2135 ( .A(n19939), .B(n1968), .Z(n1969) );
  NANDN U2136 ( .A(y[3965]), .B(n1969), .Z(n1970) );
  ANDN U2137 ( .B(n1970), .A(n10625), .Z(n1971) );
  XNOR U2138 ( .A(n1969), .B(y[3965]), .Z(n1972) );
  NAND U2139 ( .A(n1972), .B(x[3965]), .Z(n1973) );
  NAND U2140 ( .A(n1971), .B(n1973), .Z(n1974) );
  NANDN U2141 ( .A(n19945), .B(n1974), .Z(n10361) );
  ANDN U2142 ( .B(n28534), .A(n10607), .Z(n1975) );
  ANDN U2143 ( .B(n10365), .A(n10612), .Z(n1976) );
  NAND U2144 ( .A(n1976), .B(n10611), .Z(n1977) );
  AND U2145 ( .A(n1975), .B(n1977), .Z(n1978) );
  NOR U2146 ( .A(n1978), .B(n10610), .Z(n1979) );
  NANDN U2147 ( .A(n19985), .B(n1979), .Z(n1980) );
  NANDN U2148 ( .A(n10608), .B(n1980), .Z(n1981) );
  ANDN U2149 ( .B(n19986), .A(n10605), .Z(n1982) );
  XNOR U2150 ( .A(y[3985]), .B(x[3985]), .Z(n1983) );
  NANDN U2151 ( .A(n1981), .B(n1983), .Z(n1984) );
  AND U2152 ( .A(n1982), .B(n1984), .Z(n1985) );
  NOR U2153 ( .A(n10606), .B(n19995), .Z(n1986) );
  NOR U2154 ( .A(n1985), .B(n19992), .Z(n1987) );
  NAND U2155 ( .A(n1987), .B(n19989), .Z(n1988) );
  AND U2156 ( .A(n1986), .B(n1988), .Z(n1989) );
  NOR U2157 ( .A(n1989), .B(n19993), .Z(n1990) );
  NANDN U2158 ( .A(n10604), .B(n1990), .Z(n1991) );
  NAND U2159 ( .A(n1991), .B(n19996), .Z(n10367) );
  NANDN U2160 ( .A(n10556), .B(n10439), .Z(n1992) );
  ANDN U2161 ( .B(n10443), .A(n28640), .Z(n1993) );
  NANDN U2162 ( .A(n1992), .B(n28638), .Z(n1994) );
  AND U2163 ( .A(n1993), .B(n1994), .Z(n1995) );
  NANDN U2164 ( .A(n1995), .B(n28642), .Z(n1996) );
  ANDN U2165 ( .B(n1996), .A(n20069), .Z(n1997) );
  ANDN U2166 ( .B(n28651), .A(n20068), .Z(n1998) );
  OR U2167 ( .A(n10553), .B(n1997), .Z(n1999) );
  AND U2168 ( .A(n1998), .B(n1999), .Z(n2000) );
  XNOR U2169 ( .A(x[4036]), .B(y[4036]), .Z(n2001) );
  NANDN U2170 ( .A(n2000), .B(n2001), .Z(n2002) );
  AND U2171 ( .A(n28657), .B(n2002), .Z(n2003) );
  ANDN U2172 ( .B(n10551), .A(n20076), .Z(n2004) );
  NANDN U2173 ( .A(n28648), .B(n2003), .Z(n2005) );
  NAND U2174 ( .A(n2004), .B(n2005), .Z(n2006) );
  NOR U2175 ( .A(n20086), .B(n28654), .Z(n2007) );
  NAND U2176 ( .A(n2007), .B(n2006), .Z(n2008) );
  NANDN U2177 ( .A(n20081), .B(n2008), .Z(n10447) );
  NOR U2178 ( .A(n20117), .B(n10540), .Z(n2009) );
  NAND U2179 ( .A(n2009), .B(n10450), .Z(n2010) );
  NAND U2180 ( .A(n2010), .B(n28689), .Z(n2011) );
  OR U2181 ( .A(n10537), .B(n2011), .Z(n2012) );
  NANDN U2182 ( .A(n20120), .B(n2012), .Z(n2013) );
  NANDN U2183 ( .A(n2013), .B(y[4056]), .Z(n2014) );
  ANDN U2184 ( .B(n2014), .A(n10534), .Z(n2015) );
  XNOR U2185 ( .A(n2013), .B(y[4056]), .Z(n2016) );
  NAND U2186 ( .A(n2016), .B(n10536), .Z(n2017) );
  NAND U2187 ( .A(n2015), .B(n2017), .Z(n2018) );
  NANDN U2188 ( .A(n20124), .B(n2018), .Z(n2019) );
  NANDN U2189 ( .A(n2019), .B(y[4058]), .Z(n2020) );
  ANDN U2190 ( .B(n2020), .A(n20131), .Z(n2021) );
  XNOR U2191 ( .A(n2019), .B(y[4058]), .Z(n2022) );
  NAND U2192 ( .A(n2022), .B(n10533), .Z(n2023) );
  NAND U2193 ( .A(n2021), .B(n2023), .Z(n2024) );
  NANDN U2194 ( .A(n20128), .B(n2024), .Z(n10452) );
  NANDN U2195 ( .A(x[0]), .B(y[0]), .Z(n2025) );
  NAND U2196 ( .A(n2025), .B(n12793), .Z(n2026) );
  NANDN U2197 ( .A(n12796), .B(n2026), .Z(n2027) );
  ANDN U2198 ( .B(n2027), .A(n12798), .Z(n2028) );
  NANDN U2199 ( .A(y[3]), .B(x[3]), .Z(n2029) );
  AND U2200 ( .A(n12800), .B(n2029), .Z(n2030) );
  XNOR U2201 ( .A(x[3]), .B(y[3]), .Z(n2031) );
  NAND U2202 ( .A(n2031), .B(n2028), .Z(n2032) );
  NAND U2203 ( .A(n2030), .B(n2032), .Z(n2033) );
  NANDN U2204 ( .A(n12806), .B(n2033), .Z(n4132) );
  ANDN U2205 ( .B(y[97]), .A(n4257), .Z(n2034) );
  NAND U2206 ( .A(y[98]), .B(n12780), .Z(n2035) );
  AND U2207 ( .A(n4259), .B(n2035), .Z(n2036) );
  NANDN U2208 ( .A(n2034), .B(n2036), .Z(n2037) );
  ANDN U2209 ( .B(n12784), .A(n12779), .Z(n2038) );
  NAND U2210 ( .A(n2038), .B(n2037), .Z(n2039) );
  NANDN U2211 ( .A(n12781), .B(n2039), .Z(n2040) );
  NAND U2212 ( .A(n2040), .B(n13036), .Z(n2041) );
  NANDN U2213 ( .A(n13039), .B(n2041), .Z(n2042) );
  AND U2214 ( .A(n13040), .B(n2042), .Z(n2043) );
  OR U2215 ( .A(n13043), .B(n2043), .Z(n2044) );
  NAND U2216 ( .A(n2044), .B(n13044), .Z(n2045) );
  NANDN U2217 ( .A(n13046), .B(n2045), .Z(n2046) );
  NAND U2218 ( .A(n2046), .B(n13048), .Z(n2047) );
  NANDN U2219 ( .A(n13051), .B(n2047), .Z(n2048) );
  AND U2220 ( .A(n13052), .B(n2048), .Z(n2049) );
  OR U2221 ( .A(n13055), .B(n2049), .Z(n2050) );
  NAND U2222 ( .A(n2050), .B(n13056), .Z(n2051) );
  NANDN U2223 ( .A(n13058), .B(n2051), .Z(n4270) );
  OR U2224 ( .A(n4439), .B(n13256), .Z(n2052) );
  ANDN U2225 ( .B(n2052), .A(n13257), .Z(n2053) );
  OR U2226 ( .A(n13260), .B(n2053), .Z(n2054) );
  NANDN U2227 ( .A(n13262), .B(n2054), .Z(n2055) );
  ANDN U2228 ( .B(n2055), .A(n13263), .Z(n2056) );
  OR U2229 ( .A(x[216]), .B(n2056), .Z(n2057) );
  XOR U2230 ( .A(x[216]), .B(n2056), .Z(n2058) );
  NAND U2231 ( .A(n2058), .B(y[216]), .Z(n2059) );
  NAND U2232 ( .A(n2057), .B(n2059), .Z(n2060) );
  ANDN U2233 ( .B(n2060), .A(n13269), .Z(n2061) );
  OR U2234 ( .A(n13272), .B(n2061), .Z(n2062) );
  NANDN U2235 ( .A(n13274), .B(n2062), .Z(n2063) );
  ANDN U2236 ( .B(n2063), .A(n13276), .Z(n2064) );
  OR U2237 ( .A(n13278), .B(n2064), .Z(n2065) );
  NANDN U2238 ( .A(n13280), .B(n2065), .Z(n2066) );
  NANDN U2239 ( .A(n13281), .B(n2066), .Z(n2067) );
  NAND U2240 ( .A(n2067), .B(n13286), .Z(n2068) );
  AND U2241 ( .A(n13283), .B(n2068), .Z(n2069) );
  NANDN U2242 ( .A(n13290), .B(n2069), .Z(n2070) );
  ANDN U2243 ( .B(n2070), .A(n13285), .Z(n4443) );
  NANDN U2244 ( .A(n13718), .B(n5202), .Z(n2071) );
  AND U2245 ( .A(n20879), .B(n2071), .Z(n2072) );
  NOR U2246 ( .A(n2072), .B(n12749), .Z(n2073) );
  NAND U2247 ( .A(n2073), .B(n20880), .Z(n2074) );
  NANDN U2248 ( .A(n20887), .B(n2074), .Z(n2075) );
  NANDN U2249 ( .A(n12751), .B(n2075), .Z(n2076) );
  NAND U2250 ( .A(n2076), .B(n20891), .Z(n2077) );
  AND U2251 ( .A(n20892), .B(n2077), .Z(n2078) );
  NANDN U2252 ( .A(n2078), .B(n20894), .Z(n2079) );
  NAND U2253 ( .A(n2079), .B(n20896), .Z(n2080) );
  NAND U2254 ( .A(n2080), .B(n20898), .Z(n2081) );
  NAND U2255 ( .A(n2081), .B(n20900), .Z(n2082) );
  NAND U2256 ( .A(n2082), .B(n20903), .Z(n2083) );
  ANDN U2257 ( .B(n2083), .A(n20905), .Z(n2084) );
  NANDN U2258 ( .A(n2084), .B(n20906), .Z(n2085) );
  ANDN U2259 ( .B(n2085), .A(n20908), .Z(n2086) );
  NANDN U2260 ( .A(n2086), .B(n20910), .Z(n2087) );
  NAND U2261 ( .A(n2087), .B(n20912), .Z(n2088) );
  NAND U2262 ( .A(n2088), .B(n20914), .Z(n5228) );
  NANDN U2263 ( .A(n6573), .B(n22266), .Z(n2089) );
  NAND U2264 ( .A(n2089), .B(n22268), .Z(n2090) );
  NAND U2265 ( .A(n2090), .B(n22271), .Z(n2091) );
  NAND U2266 ( .A(n2091), .B(n22272), .Z(n2092) );
  NANDN U2267 ( .A(n22275), .B(n2092), .Z(n2093) );
  ANDN U2268 ( .B(n2093), .A(n14616), .Z(n2094) );
  OR U2269 ( .A(n12612), .B(n2094), .Z(n2095) );
  NANDN U2270 ( .A(n14617), .B(n2095), .Z(n2096) );
  ANDN U2271 ( .B(n2096), .A(n14622), .Z(n2097) );
  OR U2272 ( .A(n6583), .B(n14621), .Z(n2098) );
  ANDN U2273 ( .B(n2098), .A(n14625), .Z(n2099) );
  NANDN U2274 ( .A(n12615), .B(n2097), .Z(n2100) );
  NAND U2275 ( .A(n2100), .B(n22280), .Z(n2101) );
  AND U2276 ( .A(n2099), .B(n2101), .Z(n2102) );
  NANDN U2277 ( .A(n2102), .B(n22284), .Z(n2103) );
  ANDN U2278 ( .B(n2103), .A(n22286), .Z(n2104) );
  NANDN U2279 ( .A(n2104), .B(n22288), .Z(n2105) );
  NANDN U2280 ( .A(n22291), .B(n2105), .Z(n2106) );
  NANDN U2281 ( .A(n12610), .B(n2106), .Z(n6591) );
  NANDN U2282 ( .A(n14955), .B(n22766), .Z(n3147) );
  NANDN U2283 ( .A(x[22]), .B(y[22]), .Z(n12861) );
  NANDN U2284 ( .A(x[56]), .B(y[56]), .Z(n12936) );
  NANDN U2285 ( .A(y[883]), .B(x[883]), .Z(n2107) );
  NAND U2286 ( .A(n2107), .B(n21530), .Z(n14110) );
  OR U2287 ( .A(n20295), .B(n21680), .Z(n14198) );
  NANDN U2288 ( .A(x[286]), .B(y[286]), .Z(n2108) );
  ANDN U2289 ( .B(n2108), .A(n4547), .Z(n20307) );
  NANDN U2290 ( .A(n20292), .B(n21820), .Z(n2109) );
  NANDN U2291 ( .A(n6142), .B(n2109), .Z(n2110) );
  AND U2292 ( .A(n21828), .B(n2110), .Z(n14282) );
  NANDN U2293 ( .A(y[364]), .B(x[364]), .Z(n20474) );
  NANDN U2294 ( .A(x[426]), .B(y[426]), .Z(n2111) );
  NANDN U2295 ( .A(n3656), .B(n2111), .Z(n20600) );
  NANDN U2296 ( .A(y[452]), .B(x[452]), .Z(n2112) );
  NANDN U2297 ( .A(y[453]), .B(x[453]), .Z(n2113) );
  AND U2298 ( .A(n2112), .B(n2113), .Z(n2114) );
  NANDN U2299 ( .A(y[454]), .B(x[454]), .Z(n2115) );
  NANDN U2300 ( .A(y[455]), .B(x[455]), .Z(n2116) );
  AND U2301 ( .A(n2115), .B(n2116), .Z(n2117) );
  OR U2302 ( .A(n3644), .B(n2114), .Z(n2118) );
  NAND U2303 ( .A(n2117), .B(n2118), .Z(n20659) );
  NANDN U2304 ( .A(x[558]), .B(y[558]), .Z(n2119) );
  NANDN U2305 ( .A(n3576), .B(n2119), .Z(n13708) );
  NANDN U2306 ( .A(y[590]), .B(x[590]), .Z(n13745) );
  NANDN U2307 ( .A(x[750]), .B(y[750]), .Z(n2120) );
  ANDN U2308 ( .B(n2120), .A(n5590), .Z(n13946) );
  NANDN U2309 ( .A(x[922]), .B(y[922]), .Z(n2121) );
  ANDN U2310 ( .B(n2121), .A(n12717), .Z(n21629) );
  NANDN U2311 ( .A(y[990]), .B(x[990]), .Z(n2122) );
  ANDN U2312 ( .B(n2122), .A(n6117), .Z(n21796) );
  NANDN U2313 ( .A(y[1032]), .B(x[1032]), .Z(n12701) );
  NANDN U2314 ( .A(x[1022]), .B(y[1022]), .Z(n2123) );
  ANDN U2315 ( .B(n2123), .A(n12707), .Z(n21868) );
  NAND U2316 ( .A(n9326), .B(n9325), .Z(n2124) );
  NAND U2317 ( .A(n2124), .B(n11911), .Z(n2125) );
  NAND U2318 ( .A(n2125), .B(n25531), .Z(n2126) );
  ANDN U2319 ( .B(n11912), .A(n25534), .Z(n2127) );
  NAND U2320 ( .A(n2127), .B(n2126), .Z(n2128) );
  NANDN U2321 ( .A(n25536), .B(n2128), .Z(n2129) );
  NAND U2322 ( .A(n2129), .B(n25537), .Z(n2130) );
  AND U2323 ( .A(n25540), .B(n2130), .Z(n2131) );
  NANDN U2324 ( .A(n11909), .B(n2131), .Z(n2132) );
  AND U2325 ( .A(n25541), .B(n2132), .Z(n2133) );
  NANDN U2326 ( .A(n2133), .B(n11905), .Z(n2134) );
  XOR U2327 ( .A(n2133), .B(y[2658]), .Z(n2135) );
  NAND U2328 ( .A(n2135), .B(x[2658]), .Z(n2136) );
  AND U2329 ( .A(n2134), .B(n2136), .Z(n2137) );
  ANDN U2330 ( .B(n25549), .A(n11906), .Z(n2138) );
  NANDN U2331 ( .A(n2137), .B(n25548), .Z(n2139) );
  AND U2332 ( .A(n2138), .B(n2139), .Z(n2140) );
  NANDN U2333 ( .A(n2140), .B(n25551), .Z(n2141) );
  AND U2334 ( .A(n25553), .B(n2141), .Z(n9327) );
  NANDN U2335 ( .A(x[1062]), .B(y[1062]), .Z(n12682) );
  NANDN U2336 ( .A(x[1127]), .B(y[1127]), .Z(n14472) );
  NANDN U2337 ( .A(y[1188]), .B(x[1188]), .Z(n12624) );
  NANDN U2338 ( .A(x[1175]), .B(y[1175]), .Z(n14547) );
  NANDN U2339 ( .A(y[1246]), .B(x[1246]), .Z(n12597) );
  NANDN U2340 ( .A(y[1320]), .B(x[1320]), .Z(n12539) );
  NANDN U2341 ( .A(x[1307]), .B(y[1307]), .Z(n14744) );
  NANDN U2342 ( .A(y[1330]), .B(x[1330]), .Z(n12532) );
  ANDN U2343 ( .B(n9686), .A(n11792), .Z(n2142) );
  NAND U2344 ( .A(n2142), .B(n26044), .Z(n2143) );
  AND U2345 ( .A(n26046), .B(n2143), .Z(n2144) );
  NANDN U2346 ( .A(n2144), .B(n26050), .Z(n2145) );
  NAND U2347 ( .A(n2145), .B(n26052), .Z(n2146) );
  NAND U2348 ( .A(n2146), .B(n17769), .Z(n2147) );
  NAND U2349 ( .A(n2147), .B(n26056), .Z(n2148) );
  NAND U2350 ( .A(n2148), .B(n26058), .Z(n2149) );
  ANDN U2351 ( .B(n2149), .A(n17773), .Z(n2150) );
  ANDN U2352 ( .B(n26064), .A(n17774), .Z(n2151) );
  OR U2353 ( .A(n17776), .B(n2150), .Z(n2152) );
  AND U2354 ( .A(n2151), .B(n2152), .Z(n2153) );
  NOR U2355 ( .A(n2153), .B(n17777), .Z(n2154) );
  NAND U2356 ( .A(n2154), .B(n26066), .Z(n2155) );
  AND U2357 ( .A(n26068), .B(n2155), .Z(n2156) );
  OR U2358 ( .A(n26071), .B(n2156), .Z(n2157) );
  NAND U2359 ( .A(n2157), .B(n26072), .Z(n2158) );
  NANDN U2360 ( .A(n26074), .B(n2158), .Z(n2159) );
  NANDN U2361 ( .A(n11784), .B(n2159), .Z(n9696) );
  NANDN U2362 ( .A(y[1354]), .B(x[1354]), .Z(n12514) );
  NANDN U2363 ( .A(y[1428]), .B(x[1428]), .Z(n12476) );
  NANDN U2364 ( .A(x[1439]), .B(y[1439]), .Z(n14930) );
  NANDN U2365 ( .A(y[1907]), .B(x[1907]), .Z(n2160) );
  ANDN U2366 ( .B(n2160), .A(n23787), .Z(n15783) );
  NANDN U2367 ( .A(x[1487]), .B(y[1487]), .Z(n12438) );
  NANDN U2368 ( .A(x[1489]), .B(y[1489]), .Z(n12434) );
  NAND U2369 ( .A(n12220), .B(x[1960]), .Z(n2161) );
  AND U2370 ( .A(n23910), .B(n2161), .Z(n15872) );
  NAND U2371 ( .A(n9835), .B(n9834), .Z(n2162) );
  NAND U2372 ( .A(n2162), .B(n9836), .Z(n2163) );
  NAND U2373 ( .A(n2163), .B(n26338), .Z(n2164) );
  ANDN U2374 ( .B(n26341), .A(n18033), .Z(n2165) );
  OR U2375 ( .A(n11716), .B(n2164), .Z(n2166) );
  AND U2376 ( .A(n2165), .B(n2166), .Z(n2167) );
  NANDN U2377 ( .A(n2167), .B(n26342), .Z(n2168) );
  ANDN U2378 ( .B(n2168), .A(n26345), .Z(n2169) );
  ANDN U2379 ( .B(n26348), .A(n11709), .Z(n2170) );
  OR U2380 ( .A(n26347), .B(n2169), .Z(n2171) );
  AND U2381 ( .A(n2170), .B(n2171), .Z(n2172) );
  NOR U2382 ( .A(n2172), .B(n18048), .Z(n2173) );
  NAND U2383 ( .A(n2173), .B(n26350), .Z(n2174) );
  AND U2384 ( .A(n26356), .B(n2174), .Z(n2175) );
  ANDN U2385 ( .B(n26358), .A(n18049), .Z(n2176) );
  NANDN U2386 ( .A(n11710), .B(n2175), .Z(n2177) );
  NAND U2387 ( .A(n2176), .B(n2177), .Z(n2178) );
  NAND U2388 ( .A(n2178), .B(n26360), .Z(n9837) );
  NANDN U2389 ( .A(y[1546]), .B(x[1546]), .Z(n15096) );
  NANDN U2390 ( .A(x[1559]), .B(y[1559]), .Z(n15116) );
  ANDN U2391 ( .B(n26430), .A(n18119), .Z(n2179) );
  ANDN U2392 ( .B(n9840), .A(n11692), .Z(n2180) );
  NAND U2393 ( .A(n2180), .B(n26428), .Z(n2181) );
  AND U2394 ( .A(n2179), .B(n2181), .Z(n2182) );
  NANDN U2395 ( .A(n2182), .B(n26432), .Z(n2183) );
  ANDN U2396 ( .B(n2183), .A(n26434), .Z(n2184) );
  ANDN U2397 ( .B(n26438), .A(n11688), .Z(n2185) );
  OR U2398 ( .A(n26437), .B(n2184), .Z(n2186) );
  NAND U2399 ( .A(n2185), .B(n2186), .Z(n2187) );
  ANDN U2400 ( .B(n26440), .A(n18137), .Z(n2188) );
  NAND U2401 ( .A(n2188), .B(n2187), .Z(n2189) );
  NAND U2402 ( .A(n2189), .B(n26446), .Z(n2190) );
  ANDN U2403 ( .B(n26449), .A(n18138), .Z(n2191) );
  OR U2404 ( .A(n11689), .B(n2190), .Z(n2192) );
  AND U2405 ( .A(n2191), .B(n2192), .Z(n2193) );
  NANDN U2406 ( .A(n2193), .B(n26450), .Z(n2194) );
  NANDN U2407 ( .A(n26453), .B(n2194), .Z(n2195) );
  NAND U2408 ( .A(n2195), .B(n26454), .Z(n9843) );
  NANDN U2409 ( .A(x[1580]), .B(y[1580]), .Z(n2196) );
  NANDN U2410 ( .A(n12384), .B(n2196), .Z(n3116) );
  NANDN U2411 ( .A(y[1621]), .B(x[1621]), .Z(n12367) );
  NANDN U2412 ( .A(x[1607]), .B(y[1607]), .Z(n15180) );
  NANDN U2413 ( .A(n9850), .B(n9849), .Z(n2197) );
  NAND U2414 ( .A(n2197), .B(n26522), .Z(n2198) );
  ANDN U2415 ( .B(n2198), .A(n26525), .Z(n2199) );
  ANDN U2416 ( .B(n26528), .A(n11667), .Z(n2200) );
  OR U2417 ( .A(n26527), .B(n2199), .Z(n2201) );
  AND U2418 ( .A(n2200), .B(n2201), .Z(n2202) );
  NOR U2419 ( .A(n2202), .B(n18229), .Z(n2203) );
  NAND U2420 ( .A(n2203), .B(n26530), .Z(n2204) );
  AND U2421 ( .A(n26536), .B(n2204), .Z(n2205) );
  ANDN U2422 ( .B(n26538), .A(n18230), .Z(n2206) );
  NANDN U2423 ( .A(n11668), .B(n2205), .Z(n2207) );
  NAND U2424 ( .A(n2206), .B(n2207), .Z(n2208) );
  NAND U2425 ( .A(n2208), .B(n26540), .Z(n2209) );
  AND U2426 ( .A(n26543), .B(n2209), .Z(n2210) );
  NANDN U2427 ( .A(n26545), .B(n2210), .Z(n2211) );
  NAND U2428 ( .A(n2211), .B(n26546), .Z(n2212) );
  AND U2429 ( .A(n26549), .B(n2212), .Z(n2213) );
  NANDN U2430 ( .A(n18245), .B(n2213), .Z(n2214) );
  AND U2431 ( .A(n26550), .B(n2214), .Z(n9852) );
  NANDN U2432 ( .A(y[1667]), .B(x[1667]), .Z(n2215) );
  NAND U2433 ( .A(n2215), .B(n12349), .Z(n23221) );
  NANDN U2434 ( .A(x[1686]), .B(y[1686]), .Z(n2216) );
  NAND U2435 ( .A(n2216), .B(n15352), .Z(n23266) );
  NANDN U2436 ( .A(y[1712]), .B(x[1712]), .Z(n12316) );
  NANDN U2437 ( .A(x[1700]), .B(y[1700]), .Z(n2217) );
  ANDN U2438 ( .B(n2217), .A(n15394), .Z(n23299) );
  OR U2439 ( .A(x[1764]), .B(n15500), .Z(n2218) );
  NANDN U2440 ( .A(n12303), .B(n2218), .Z(n23436) );
  NANDN U2441 ( .A(x[1793]), .B(y[1793]), .Z(n2219) );
  NANDN U2442 ( .A(x[1792]), .B(y[1792]), .Z(n2220) );
  NAND U2443 ( .A(n2219), .B(n2220), .Z(n23500) );
  NANDN U2444 ( .A(y[1837]), .B(x[1837]), .Z(n12270) );
  NANDN U2445 ( .A(x[1814]), .B(y[1814]), .Z(n2221) );
  ANDN U2446 ( .B(n2221), .A(n12281), .Z(n23554) );
  NANDN U2447 ( .A(x[1856]), .B(y[1856]), .Z(n2222) );
  ANDN U2448 ( .B(n2222), .A(n12260), .Z(n23667) );
  NANDN U2449 ( .A(y[1877]), .B(x[1877]), .Z(n2223) );
  NAND U2450 ( .A(n2223), .B(n12251), .Z(n23715) );
  NANDN U2451 ( .A(x[1898]), .B(y[1898]), .Z(n2224) );
  ANDN U2452 ( .B(n2224), .A(n12239), .Z(n23761) );
  NANDN U2453 ( .A(y[1995]), .B(x[1995]), .Z(n2225) );
  ANDN U2454 ( .B(n2225), .A(n12206), .Z(n23999) );
  NANDN U2455 ( .A(x[2038]), .B(y[2038]), .Z(n2226) );
  ANDN U2456 ( .B(n2226), .A(n12191), .Z(n24101) );
  NANDN U2457 ( .A(y[2064]), .B(x[2064]), .Z(n2227) );
  ANDN U2458 ( .B(n2227), .A(n12185), .Z(n24154) );
  NANDN U2459 ( .A(x[2079]), .B(y[2079]), .Z(n2228) );
  ANDN U2460 ( .B(n2228), .A(n16115), .Z(n24189) );
  ANDN U2461 ( .B(n12164), .A(n16173), .Z(n24237) );
  NANDN U2462 ( .A(y[2155]), .B(x[2155]), .Z(n2229) );
  NAND U2463 ( .A(n2229), .B(n12146), .Z(n24361) );
  NANDN U2464 ( .A(x[2172]), .B(y[2172]), .Z(n2230) );
  NANDN U2465 ( .A(x[2173]), .B(y[2173]), .Z(n2231) );
  AND U2466 ( .A(n2230), .B(n2231), .Z(n24404) );
  NANDN U2467 ( .A(y[2248]), .B(x[2248]), .Z(n2232) );
  NANDN U2468 ( .A(y[2247]), .B(x[2247]), .Z(n2233) );
  NAND U2469 ( .A(n2232), .B(n2233), .Z(n24586) );
  NANDN U2470 ( .A(x[2316]), .B(y[2316]), .Z(n2234) );
  NAND U2471 ( .A(n2234), .B(n12080), .Z(n24743) );
  NANDN U2472 ( .A(y[2365]), .B(x[2365]), .Z(n2235) );
  ANDN U2473 ( .B(n2235), .A(n12052), .Z(n24845) );
  NANDN U2474 ( .A(y[2401]), .B(x[2401]), .Z(n2236) );
  ANDN U2475 ( .B(n2236), .A(n12034), .Z(n24934) );
  NANDN U2476 ( .A(y[2457]), .B(x[2457]), .Z(n2237) );
  ANDN U2477 ( .B(n2237), .A(n12010), .Z(n25076) );
  NANDN U2478 ( .A(x[2498]), .B(y[2498]), .Z(n17028) );
  NANDN U2479 ( .A(n17114), .B(n17108), .Z(n25257) );
  NANDN U2480 ( .A(x[2599]), .B(y[2599]), .Z(n11942) );
  NANDN U2481 ( .A(n11157), .B(n10150), .Z(n2238) );
  ANDN U2482 ( .B(n2238), .A(n19022), .Z(n2239) );
  NAND U2483 ( .A(n11155), .B(x[3497]), .Z(n2240) );
  ANDN U2484 ( .B(n2240), .A(n11154), .Z(n2241) );
  XOR U2485 ( .A(x[3497]), .B(n11155), .Z(n2242) );
  NAND U2486 ( .A(n2242), .B(n2239), .Z(n2243) );
  NAND U2487 ( .A(n2241), .B(n2243), .Z(n2244) );
  AND U2488 ( .A(n19027), .B(n2244), .Z(n2245) );
  OR U2489 ( .A(x[3499]), .B(n2245), .Z(n2246) );
  XOR U2490 ( .A(n2245), .B(x[3499]), .Z(n2247) );
  NAND U2491 ( .A(n2247), .B(y[3499]), .Z(n2248) );
  NAND U2492 ( .A(n2246), .B(n2248), .Z(n2249) );
  ANDN U2493 ( .B(n2249), .A(n11150), .Z(n2250) );
  NOR U2494 ( .A(n2250), .B(n11152), .Z(n2251) );
  NAND U2495 ( .A(n2251), .B(n27478), .Z(n2252) );
  ANDN U2496 ( .B(n2252), .A(n11149), .Z(n2253) );
  NAND U2497 ( .A(n2253), .B(n11148), .Z(n2254) );
  AND U2498 ( .A(n27476), .B(n2254), .Z(n2255) );
  NANDN U2499 ( .A(n11144), .B(n2255), .Z(n10151) );
  NANDN U2500 ( .A(y[2591]), .B(x[2591]), .Z(n2256) );
  ANDN U2501 ( .B(n2256), .A(n17227), .Z(n25387) );
  NANDN U2502 ( .A(n19058), .B(n10153), .Z(n2257) );
  NANDN U2503 ( .A(n2257), .B(y[3518]), .Z(n2258) );
  ANDN U2504 ( .B(n2258), .A(n11128), .Z(n2259) );
  XNOR U2505 ( .A(n2257), .B(y[3518]), .Z(n2260) );
  NAND U2506 ( .A(n2260), .B(n19061), .Z(n2261) );
  NAND U2507 ( .A(n2259), .B(n2261), .Z(n2262) );
  ANDN U2508 ( .B(n2262), .A(n19065), .Z(n2263) );
  OR U2509 ( .A(y[3520]), .B(n2263), .Z(n2264) );
  XOR U2510 ( .A(n2263), .B(y[3520]), .Z(n2265) );
  NAND U2511 ( .A(n2265), .B(x[3520]), .Z(n2266) );
  NAND U2512 ( .A(n2264), .B(n2266), .Z(n2267) );
  ANDN U2513 ( .B(n2267), .A(n11124), .Z(n2268) );
  NOR U2514 ( .A(n2268), .B(n11126), .Z(n2269) );
  NAND U2515 ( .A(n2269), .B(n19071), .Z(n2270) );
  AND U2516 ( .A(n27523), .B(n2270), .Z(n2271) );
  ANDN U2517 ( .B(n19075), .A(n19072), .Z(n2272) );
  NANDN U2518 ( .A(n11123), .B(n2271), .Z(n2273) );
  NAND U2519 ( .A(n2272), .B(n2273), .Z(n10154) );
  XNOR U2520 ( .A(x[3542]), .B(y[3542]), .Z(n2274) );
  ANDN U2521 ( .B(n2274), .A(n11109), .Z(n2275) );
  NAND U2522 ( .A(n10156), .B(n11112), .Z(n2276) );
  NANDN U2523 ( .A(n10157), .B(y[3538]), .Z(n2277) );
  AND U2524 ( .A(n2276), .B(n2277), .Z(n2278) );
  ANDN U2525 ( .B(n11108), .A(n19112), .Z(n2279) );
  NANDN U2526 ( .A(n11111), .B(n2278), .Z(n2280) );
  NAND U2527 ( .A(n2279), .B(n2280), .Z(n2281) );
  ANDN U2528 ( .B(n27564), .A(n11110), .Z(n2282) );
  NAND U2529 ( .A(n2282), .B(n2281), .Z(n2283) );
  NAND U2530 ( .A(n2283), .B(n2275), .Z(n2284) );
  ANDN U2531 ( .B(n27562), .A(n11106), .Z(n2285) );
  NAND U2532 ( .A(n2285), .B(n2284), .Z(n2286) );
  ANDN U2533 ( .B(n2286), .A(n19119), .Z(n2287) );
  NANDN U2534 ( .A(x[3544]), .B(n2287), .Z(n2288) );
  ANDN U2535 ( .B(n2288), .A(n11104), .Z(n2289) );
  XNOR U2536 ( .A(n2287), .B(x[3544]), .Z(n2290) );
  NAND U2537 ( .A(n2290), .B(y[3544]), .Z(n2291) );
  NAND U2538 ( .A(n2289), .B(n2291), .Z(n10158) );
  NANDN U2539 ( .A(y[2816]), .B(x[2816]), .Z(n2292) );
  ANDN U2540 ( .B(n2292), .A(n25939), .Z(n17680) );
  NANDN U2541 ( .A(y[2720]), .B(x[2720]), .Z(n2293) );
  NANDN U2542 ( .A(y[2719]), .B(x[2719]), .Z(n2294) );
  NAND U2543 ( .A(n2293), .B(n2294), .Z(n25697) );
  ANDN U2544 ( .B(n25973), .A(n25983), .Z(n17709) );
  OR U2545 ( .A(n10161), .B(n10162), .Z(n2295) );
  AND U2546 ( .A(n20225), .B(n2295), .Z(n2296) );
  ANDN U2547 ( .B(n19147), .A(n11081), .Z(n2297) );
  NANDN U2548 ( .A(n11082), .B(n2296), .Z(n2298) );
  AND U2549 ( .A(n2297), .B(n2298), .Z(n2299) );
  NOR U2550 ( .A(n2299), .B(n20224), .Z(n2300) );
  NAND U2551 ( .A(n2300), .B(n27605), .Z(n2301) );
  AND U2552 ( .A(n19153), .B(n2301), .Z(n2302) );
  NOR U2553 ( .A(n19156), .B(n27604), .Z(n2303) );
  NANDN U2554 ( .A(n19149), .B(n2302), .Z(n2304) );
  NAND U2555 ( .A(n2303), .B(n2304), .Z(n2305) );
  NANDN U2556 ( .A(n11078), .B(n2305), .Z(n2306) );
  NOR U2557 ( .A(n19157), .B(n19160), .Z(n2307) );
  OR U2558 ( .A(n11076), .B(n2306), .Z(n2308) );
  AND U2559 ( .A(n2307), .B(n2308), .Z(n2309) );
  NOR U2560 ( .A(n2309), .B(n11077), .Z(n2310) );
  NANDN U2561 ( .A(n11075), .B(n2310), .Z(n2311) );
  NANDN U2562 ( .A(n19161), .B(n2311), .Z(n10164) );
  NANDN U2563 ( .A(y[2745]), .B(x[2745]), .Z(n2312) );
  ANDN U2564 ( .B(n2312), .A(n11856), .Z(n25760) );
  NANDN U2565 ( .A(y[2767]), .B(x[2767]), .Z(n2313) );
  NAND U2566 ( .A(n2313), .B(n11831), .Z(n25817) );
  NOR U2567 ( .A(n11048), .B(n27652), .Z(n2314) );
  OR U2568 ( .A(n10168), .B(n10169), .Z(n2315) );
  AND U2569 ( .A(n2314), .B(n2315), .Z(n2316) );
  NOR U2570 ( .A(n11050), .B(n19196), .Z(n2317) );
  NANDN U2571 ( .A(n2316), .B(n2317), .Z(n2318) );
  ANDN U2572 ( .B(n2318), .A(n27662), .Z(n2319) );
  NOR U2573 ( .A(n11046), .B(n19195), .Z(n2320) );
  NANDN U2574 ( .A(n11047), .B(n2319), .Z(n2321) );
  NAND U2575 ( .A(n2320), .B(n2321), .Z(n2322) );
  NOR U2576 ( .A(n11043), .B(n27663), .Z(n2323) );
  NAND U2577 ( .A(n2323), .B(n2322), .Z(n2324) );
  ANDN U2578 ( .B(n2324), .A(n11044), .Z(n2325) );
  NANDN U2579 ( .A(x[3590]), .B(n2325), .Z(n2326) );
  ANDN U2580 ( .B(n2326), .A(n11039), .Z(n2327) );
  XNOR U2581 ( .A(n2325), .B(x[3590]), .Z(n2328) );
  NAND U2582 ( .A(n2328), .B(y[3590]), .Z(n2329) );
  NAND U2583 ( .A(n2327), .B(n2329), .Z(n2330) );
  NAND U2584 ( .A(n2330), .B(n11041), .Z(n10171) );
  NANDN U2585 ( .A(y[2840]), .B(x[2840]), .Z(n17737) );
  NANDN U2586 ( .A(n10175), .B(x[3609]), .Z(n2331) );
  NANDN U2587 ( .A(y[3609]), .B(n10174), .Z(n2332) );
  NAND U2588 ( .A(n2331), .B(n2332), .Z(n2333) );
  OR U2589 ( .A(n11023), .B(n2333), .Z(n2334) );
  NANDN U2590 ( .A(n19242), .B(n2334), .Z(n2335) );
  NANDN U2591 ( .A(n2335), .B(x[3611]), .Z(n2336) );
  ANDN U2592 ( .B(n2336), .A(n11018), .Z(n2337) );
  XNOR U2593 ( .A(n2335), .B(x[3611]), .Z(n2338) );
  NAND U2594 ( .A(n2338), .B(n11021), .Z(n2339) );
  NAND U2595 ( .A(n2337), .B(n2339), .Z(n2340) );
  ANDN U2596 ( .B(n2340), .A(n11019), .Z(n2341) );
  NANDN U2597 ( .A(y[3613]), .B(n2341), .Z(n2342) );
  ANDN U2598 ( .B(n2342), .A(n11016), .Z(n2343) );
  XNOR U2599 ( .A(n2341), .B(y[3613]), .Z(n2344) );
  NAND U2600 ( .A(n2344), .B(x[3613]), .Z(n2345) );
  NAND U2601 ( .A(n2343), .B(n2345), .Z(n2346) );
  NANDN U2602 ( .A(n19248), .B(n2346), .Z(n10177) );
  ANDN U2603 ( .B(n19288), .A(n19284), .Z(n2347) );
  NAND U2604 ( .A(n2347), .B(n10182), .Z(n2348) );
  ANDN U2605 ( .B(n2348), .A(n19291), .Z(n2349) );
  NOR U2606 ( .A(n19294), .B(n10999), .Z(n2350) );
  NANDN U2607 ( .A(n20222), .B(n2349), .Z(n2351) );
  NAND U2608 ( .A(n2350), .B(n2351), .Z(n2352) );
  NOR U2609 ( .A(n19292), .B(n19297), .Z(n2353) );
  NAND U2610 ( .A(n2353), .B(n2352), .Z(n2354) );
  NANDN U2611 ( .A(n19295), .B(n2354), .Z(n2355) );
  OR U2612 ( .A(n10998), .B(n2355), .Z(n2356) );
  NANDN U2613 ( .A(n19298), .B(n2356), .Z(n2357) );
  NANDN U2614 ( .A(n2357), .B(x[3637]), .Z(n2358) );
  ANDN U2615 ( .B(n2358), .A(n10993), .Z(n2359) );
  XNOR U2616 ( .A(n2357), .B(x[3637]), .Z(n2360) );
  NAND U2617 ( .A(n2360), .B(n10996), .Z(n2361) );
  NAND U2618 ( .A(n2359), .B(n2361), .Z(n2362) );
  NANDN U2619 ( .A(n10994), .B(n2362), .Z(n10184) );
  NAND U2620 ( .A(n17861), .B(x[2899]), .Z(n2363) );
  NANDN U2621 ( .A(y[2900]), .B(x[2900]), .Z(n2364) );
  AND U2622 ( .A(n2363), .B(n2364), .Z(n26152) );
  NAND U2623 ( .A(y[2920]), .B(n17901), .Z(n2365) );
  NANDN U2624 ( .A(x[2921]), .B(y[2921]), .Z(n2366) );
  NAND U2625 ( .A(n2365), .B(n2366), .Z(n26204) );
  NANDN U2626 ( .A(y[2952]), .B(x[2952]), .Z(n11729) );
  XNOR U2627 ( .A(y[3647]), .B(x[3647]), .Z(n2367) );
  NAND U2628 ( .A(n2367), .B(n10186), .Z(n2368) );
  ANDN U2629 ( .B(n19317), .A(n10982), .Z(n2369) );
  NAND U2630 ( .A(n2369), .B(n2368), .Z(n2370) );
  ANDN U2631 ( .B(n2370), .A(n10981), .Z(n2371) );
  NANDN U2632 ( .A(n19319), .B(n2371), .Z(n2372) );
  NOR U2633 ( .A(n10983), .B(n10979), .Z(n2373) );
  NAND U2634 ( .A(n2373), .B(n2372), .Z(n2374) );
  NAND U2635 ( .A(n2374), .B(n27807), .Z(n2375) );
  ANDN U2636 ( .B(n19326), .A(n10978), .Z(n2376) );
  OR U2637 ( .A(n10980), .B(n2375), .Z(n2377) );
  AND U2638 ( .A(n2376), .B(n2377), .Z(n2378) );
  NOR U2639 ( .A(n2378), .B(n27806), .Z(n2379) );
  NAND U2640 ( .A(n2379), .B(n27814), .Z(n2380) );
  AND U2641 ( .A(n19331), .B(n2380), .Z(n2381) );
  NOR U2642 ( .A(n19336), .B(n27812), .Z(n2382) );
  NANDN U2643 ( .A(n10976), .B(n2381), .Z(n2383) );
  NAND U2644 ( .A(n2382), .B(n2383), .Z(n10188) );
  NANDN U2645 ( .A(n10948), .B(n10210), .Z(n2384) );
  ANDN U2646 ( .B(n2384), .A(n19378), .Z(n2385) );
  NAND U2647 ( .A(y[3680]), .B(n10946), .Z(n2386) );
  ANDN U2648 ( .B(n2386), .A(n10945), .Z(n2387) );
  XOR U2649 ( .A(n10946), .B(y[3680]), .Z(n2388) );
  NAND U2650 ( .A(n2388), .B(n2385), .Z(n2389) );
  NAND U2651 ( .A(n2387), .B(n2389), .Z(n2390) );
  AND U2652 ( .A(n19383), .B(n2390), .Z(n2391) );
  NANDN U2653 ( .A(x[3682]), .B(n2391), .Z(n2392) );
  ANDN U2654 ( .B(n2392), .A(n10941), .Z(n2393) );
  XNOR U2655 ( .A(n2391), .B(x[3682]), .Z(n2394) );
  NAND U2656 ( .A(n2394), .B(y[3682]), .Z(n2395) );
  NAND U2657 ( .A(n2393), .B(n2395), .Z(n2396) );
  AND U2658 ( .A(n10943), .B(n2396), .Z(n2397) );
  NANDN U2659 ( .A(x[3684]), .B(n2397), .Z(n2398) );
  ANDN U2660 ( .B(n2398), .A(n19393), .Z(n2399) );
  XNOR U2661 ( .A(n2397), .B(x[3684]), .Z(n2400) );
  NAND U2662 ( .A(n2400), .B(y[3684]), .Z(n2401) );
  NAND U2663 ( .A(n2399), .B(n2401), .Z(n10211) );
  NOR U2664 ( .A(n27913), .B(n10925), .Z(n2402) );
  OR U2665 ( .A(n10213), .B(n10214), .Z(n2403) );
  NAND U2666 ( .A(n2402), .B(n2403), .Z(n2404) );
  NOR U2667 ( .A(n19418), .B(n10923), .Z(n2405) );
  NAND U2668 ( .A(n2405), .B(n2404), .Z(n2406) );
  NAND U2669 ( .A(n2406), .B(n27911), .Z(n2407) );
  OR U2670 ( .A(n19426), .B(n2407), .Z(n2408) );
  ANDN U2671 ( .B(n2408), .A(n19421), .Z(n2409) );
  NAND U2672 ( .A(n19424), .B(y[3702]), .Z(n2410) );
  ANDN U2673 ( .B(n2410), .A(n19431), .Z(n2411) );
  XOR U2674 ( .A(y[3702]), .B(n19424), .Z(n2412) );
  NAND U2675 ( .A(n2412), .B(n2409), .Z(n2413) );
  NAND U2676 ( .A(n2411), .B(n2413), .Z(n2414) );
  NANDN U2677 ( .A(n19428), .B(n2414), .Z(n2415) );
  NANDN U2678 ( .A(y[3704]), .B(x[3704]), .Z(n2416) );
  XNOR U2679 ( .A(y[3704]), .B(x[3704]), .Z(n2417) );
  NAND U2680 ( .A(n2417), .B(n2415), .Z(n2418) );
  NAND U2681 ( .A(n2416), .B(n2418), .Z(n10215) );
  NANDN U2682 ( .A(x[3081]), .B(y[3081]), .Z(n18297) );
  NANDN U2683 ( .A(x[3087]), .B(y[3087]), .Z(n11633) );
  NANDN U2684 ( .A(y[3104]), .B(x[3104]), .Z(n11610) );
  NANDN U2685 ( .A(y[3120]), .B(x[3120]), .Z(n11582) );
  NANDN U2686 ( .A(y[3108]), .B(x[3108]), .Z(n11602) );
  NOR U2687 ( .A(n27954), .B(n10914), .Z(n2419) );
  NAND U2688 ( .A(n2419), .B(n10218), .Z(n2420) );
  ANDN U2689 ( .B(n2420), .A(n10913), .Z(n2421) );
  NOR U2690 ( .A(n27955), .B(n10912), .Z(n2422) );
  NANDN U2691 ( .A(n19470), .B(n2421), .Z(n2423) );
  NAND U2692 ( .A(n2422), .B(n2423), .Z(n2424) );
  ANDN U2693 ( .B(n2424), .A(n19475), .Z(n2425) );
  OR U2694 ( .A(y[3722]), .B(n2425), .Z(n2426) );
  XOR U2695 ( .A(n2425), .B(y[3722]), .Z(n2427) );
  NAND U2696 ( .A(n2427), .B(x[3722]), .Z(n2428) );
  NAND U2697 ( .A(n2426), .B(n2428), .Z(n2429) );
  ANDN U2698 ( .B(n2429), .A(n19481), .Z(n2430) );
  NOR U2699 ( .A(n10910), .B(n19484), .Z(n2431) );
  NANDN U2700 ( .A(n2430), .B(n2431), .Z(n2432) );
  ANDN U2701 ( .B(n2432), .A(n27971), .Z(n2433) );
  NOR U2702 ( .A(n19483), .B(n10908), .Z(n2434) );
  NANDN U2703 ( .A(n19480), .B(n2433), .Z(n2435) );
  NAND U2704 ( .A(n2434), .B(n2435), .Z(n10219) );
  NANDN U2705 ( .A(y[3138]), .B(x[3138]), .Z(n18378) );
  NANDN U2706 ( .A(y[3128]), .B(x[3128]), .Z(n11569) );
  NANDN U2707 ( .A(y[3144]), .B(x[3144]), .Z(n11556) );
  NANDN U2708 ( .A(x[3165]), .B(y[3165]), .Z(n11537) );
  NANDN U2709 ( .A(x[3169]), .B(y[3169]), .Z(n18435) );
  NANDN U2710 ( .A(y[3182]), .B(x[3182]), .Z(n18460) );
  NANDN U2711 ( .A(n10886), .B(n10221), .Z(n2436) );
  ANDN U2712 ( .B(n2436), .A(n10887), .Z(n2437) );
  NANDN U2713 ( .A(x[3742]), .B(y[3742]), .Z(n2438) );
  ANDN U2714 ( .B(n2438), .A(n10884), .Z(n2439) );
  XNOR U2715 ( .A(y[3742]), .B(x[3742]), .Z(n2440) );
  NAND U2716 ( .A(n2440), .B(n2437), .Z(n2441) );
  NAND U2717 ( .A(n2439), .B(n2441), .Z(n2442) );
  ANDN U2718 ( .B(n19519), .A(n19515), .Z(n2443) );
  NAND U2719 ( .A(n2443), .B(n2442), .Z(n2444) );
  NANDN U2720 ( .A(n20219), .B(n2444), .Z(n2445) );
  NOR U2721 ( .A(n19520), .B(n19522), .Z(n2446) );
  OR U2722 ( .A(n10883), .B(n2445), .Z(n2447) );
  AND U2723 ( .A(n2446), .B(n2447), .Z(n2448) );
  NOR U2724 ( .A(n2448), .B(n20218), .Z(n2449) );
  NAND U2725 ( .A(n2449), .B(n28017), .Z(n2450) );
  ANDN U2726 ( .B(n2450), .A(n10880), .Z(n2451) );
  NOR U2727 ( .A(n28016), .B(n19531), .Z(n2452) );
  NANDN U2728 ( .A(n10881), .B(n2451), .Z(n2453) );
  NAND U2729 ( .A(n2452), .B(n2453), .Z(n10222) );
  NANDN U2730 ( .A(y[3198]), .B(x[3198]), .Z(n11497) );
  NANDN U2731 ( .A(y[3186]), .B(x[3186]), .Z(n11513) );
  NANDN U2732 ( .A(y[3214]), .B(x[3214]), .Z(n11477) );
  NANDN U2733 ( .A(y[3206]), .B(x[3206]), .Z(n11487) );
  NANDN U2734 ( .A(y[3222]), .B(x[3222]), .Z(n18528) );
  NANDN U2735 ( .A(y[3238]), .B(x[3238]), .Z(n11445) );
  NANDN U2736 ( .A(y[3226]), .B(x[3226]), .Z(n11461) );
  NANDN U2737 ( .A(y[3242]), .B(x[3242]), .Z(n18562) );
  NAND U2738 ( .A(n10226), .B(n10227), .Z(n2454) );
  ANDN U2739 ( .B(n2454), .A(n10865), .Z(n2455) );
  ANDN U2740 ( .B(n20216), .A(n19564), .Z(n2456) );
  NAND U2741 ( .A(n2455), .B(n10864), .Z(n2457) );
  AND U2742 ( .A(n2456), .B(n2457), .Z(n2458) );
  NOR U2743 ( .A(n2458), .B(n10863), .Z(n2459) );
  NANDN U2744 ( .A(n19567), .B(n2459), .Z(n2460) );
  ANDN U2745 ( .B(n2460), .A(n19565), .Z(n2461) );
  NANDN U2746 ( .A(n10860), .B(n19568), .Z(n2462) );
  XNOR U2747 ( .A(y[3767]), .B(x[3767]), .Z(n2463) );
  NAND U2748 ( .A(n2463), .B(n2461), .Z(n2464) );
  NANDN U2749 ( .A(n2462), .B(n2464), .Z(n2465) );
  OR U2750 ( .A(n10861), .B(n19576), .Z(n2466) );
  NOR U2751 ( .A(n10859), .B(n19570), .Z(n2467) );
  NAND U2752 ( .A(n2467), .B(n2465), .Z(n2468) );
  NANDN U2753 ( .A(n2466), .B(n2468), .Z(n2469) );
  AND U2754 ( .A(n28068), .B(n2469), .Z(n10228) );
  NANDN U2755 ( .A(y[3258]), .B(x[3258]), .Z(n11420) );
  NANDN U2756 ( .A(y[3246]), .B(x[3246]), .Z(n11435) );
  NANDN U2757 ( .A(x[3277]), .B(y[3277]), .Z(n18621) );
  NANDN U2758 ( .A(x[3283]), .B(y[3283]), .Z(n11396) );
  NANDN U2759 ( .A(x[3289]), .B(y[3289]), .Z(n11387) );
  NANDN U2760 ( .A(x[3295]), .B(y[3295]), .Z(n11377) );
  NANDN U2761 ( .A(x[3301]), .B(y[3301]), .Z(n11369) );
  ANDN U2762 ( .B(n10232), .A(n19608), .Z(n2470) );
  NANDN U2763 ( .A(x[3786]), .B(n2470), .Z(n2471) );
  ANDN U2764 ( .B(n2471), .A(n10843), .Z(n2472) );
  XNOR U2765 ( .A(n2470), .B(x[3786]), .Z(n2473) );
  NAND U2766 ( .A(n2473), .B(y[3786]), .Z(n2474) );
  NAND U2767 ( .A(n2472), .B(n2474), .Z(n2475) );
  ANDN U2768 ( .B(n2475), .A(n19612), .Z(n2476) );
  NANDN U2769 ( .A(x[3788]), .B(n2476), .Z(n2477) );
  ANDN U2770 ( .B(n2477), .A(n10842), .Z(n2478) );
  XNOR U2771 ( .A(n2476), .B(x[3788]), .Z(n2479) );
  NAND U2772 ( .A(n2479), .B(y[3788]), .Z(n2480) );
  NAND U2773 ( .A(n2478), .B(n2480), .Z(n2481) );
  AND U2774 ( .A(n19617), .B(n2481), .Z(n2482) );
  NAND U2775 ( .A(y[3790]), .B(n10840), .Z(n2483) );
  ANDN U2776 ( .B(n2483), .A(n10839), .Z(n2484) );
  XOR U2777 ( .A(n10840), .B(y[3790]), .Z(n2485) );
  NAND U2778 ( .A(n2485), .B(n2482), .Z(n2486) );
  AND U2779 ( .A(n2484), .B(n2486), .Z(n10234) );
  NANDN U2780 ( .A(x[3313]), .B(y[3313]), .Z(n11350) );
  NANDN U2781 ( .A(x[3317]), .B(y[3317]), .Z(n18688) );
  NANDN U2782 ( .A(x[3305]), .B(y[3305]), .Z(n11362) );
  NANDN U2783 ( .A(y[3330]), .B(x[3330]), .Z(n11332) );
  NANDN U2784 ( .A(x[3349]), .B(y[3349]), .Z(n11311) );
  NANDN U2785 ( .A(x[3353]), .B(y[3353]), .Z(n11306) );
  NANDN U2786 ( .A(n10237), .B(y[3806]), .Z(n2487) );
  NAND U2787 ( .A(n2487), .B(n10239), .Z(n2488) );
  NAND U2788 ( .A(n2488), .B(n10815), .Z(n2489) );
  ANDN U2789 ( .B(n2489), .A(n10817), .Z(n2490) );
  XNOR U2790 ( .A(x[3807]), .B(n2488), .Z(n2491) );
  NAND U2791 ( .A(n2491), .B(y[3807]), .Z(n2492) );
  NAND U2792 ( .A(n2492), .B(n2490), .Z(n2493) );
  NAND U2793 ( .A(n2493), .B(n28147), .Z(n2494) );
  NAND U2794 ( .A(n2494), .B(n28148), .Z(n2495) );
  ANDN U2795 ( .B(n2495), .A(n28150), .Z(n2496) );
  OR U2796 ( .A(n10814), .B(n2496), .Z(n2497) );
  NANDN U2797 ( .A(n19658), .B(n2497), .Z(n2498) );
  NAND U2798 ( .A(n2498), .B(n28158), .Z(n2499) );
  NOR U2799 ( .A(n19657), .B(n10812), .Z(n2500) );
  OR U2800 ( .A(n10813), .B(n2499), .Z(n2501) );
  AND U2801 ( .A(n2500), .B(n2501), .Z(n2502) );
  NOR U2802 ( .A(n2502), .B(n10811), .Z(n2503) );
  NAND U2803 ( .A(n2503), .B(n28156), .Z(n2504) );
  NANDN U2804 ( .A(n19662), .B(n2504), .Z(n10247) );
  NANDN U2805 ( .A(y[3372]), .B(x[3372]), .Z(n11287) );
  NANDN U2806 ( .A(y[3376]), .B(x[3376]), .Z(n11281) );
  NANDN U2807 ( .A(y[3394]), .B(x[3394]), .Z(n11264) );
  NANDN U2808 ( .A(y[3406]), .B(x[3406]), .Z(n11247) );
  NANDN U2809 ( .A(y[3398]), .B(x[3398]), .Z(n11257) );
  ANDN U2810 ( .B(n10270), .A(n20212), .Z(n2505) );
  NAND U2811 ( .A(n2505), .B(n10798), .Z(n2506) );
  NANDN U2812 ( .A(n10795), .B(n2506), .Z(n2507) );
  OR U2813 ( .A(n10796), .B(n2507), .Z(n2508) );
  AND U2814 ( .A(n20213), .B(n2508), .Z(n2509) );
  NANDN U2815 ( .A(y[3829]), .B(x[3829]), .Z(n2510) );
  ANDN U2816 ( .B(n2510), .A(n10790), .Z(n2511) );
  XNOR U2817 ( .A(x[3829]), .B(y[3829]), .Z(n2512) );
  NAND U2818 ( .A(n2512), .B(n2509), .Z(n2513) );
  NAND U2819 ( .A(n2511), .B(n2513), .Z(n2514) );
  ANDN U2820 ( .B(n28202), .A(n10792), .Z(n2515) );
  NAND U2821 ( .A(n2515), .B(n2514), .Z(n2516) );
  NANDN U2822 ( .A(n10789), .B(n2516), .Z(n2517) );
  ANDN U2823 ( .B(n28200), .A(n19694), .Z(n2518) );
  NANDN U2824 ( .A(n2517), .B(n10788), .Z(n2519) );
  AND U2825 ( .A(n2518), .B(n2519), .Z(n2520) );
  NOR U2826 ( .A(n19697), .B(n10787), .Z(n2521) );
  NANDN U2827 ( .A(n2520), .B(n2521), .Z(n2522) );
  ANDN U2828 ( .B(n2522), .A(n19695), .Z(n10271) );
  NANDN U2829 ( .A(x[3417]), .B(y[3417]), .Z(n18867) );
  NANDN U2830 ( .A(x[3423]), .B(y[3423]), .Z(n11225) );
  NANDN U2831 ( .A(x[3427]), .B(y[3427]), .Z(n18885) );
  NANDN U2832 ( .A(x[3439]), .B(y[3439]), .Z(n11207) );
  NANDN U2833 ( .A(x[3447]), .B(y[3447]), .Z(n11199) );
  NANDN U2834 ( .A(x[3463]), .B(y[3463]), .Z(n18959) );
  NANDN U2835 ( .A(x[3467]), .B(y[3467]), .Z(n11182) );
  NANDN U2836 ( .A(x[3455]), .B(y[3455]), .Z(n18943) );
  NOR U2837 ( .A(n19729), .B(n10770), .Z(n2523) );
  NAND U2838 ( .A(n2523), .B(n10295), .Z(n2524) );
  NANDN U2839 ( .A(n28242), .B(n2524), .Z(n2525) );
  OR U2840 ( .A(n10767), .B(n2525), .Z(n2526) );
  ANDN U2841 ( .B(n2526), .A(n10768), .Z(n2527) );
  NANDN U2842 ( .A(x[3854]), .B(y[3854]), .Z(n2528) );
  ANDN U2843 ( .B(n2528), .A(n10765), .Z(n2529) );
  XNOR U2844 ( .A(y[3854]), .B(x[3854]), .Z(n2530) );
  NAND U2845 ( .A(n2530), .B(n2527), .Z(n2531) );
  NAND U2846 ( .A(n2529), .B(n2531), .Z(n2532) );
  ANDN U2847 ( .B(n2532), .A(n19734), .Z(n2533) );
  NAND U2848 ( .A(n10763), .B(y[3856]), .Z(n2534) );
  ANDN U2849 ( .B(n2534), .A(n10760), .Z(n2535) );
  XOR U2850 ( .A(y[3856]), .B(n10763), .Z(n2536) );
  NAND U2851 ( .A(n2536), .B(n2533), .Z(n2537) );
  NAND U2852 ( .A(n2535), .B(n2537), .Z(n2538) );
  NANDN U2853 ( .A(n10761), .B(n2538), .Z(n10297) );
  AND U2854 ( .A(n10300), .B(n10301), .Z(n2539) );
  NAND U2855 ( .A(n19762), .B(y[3872]), .Z(n2540) );
  ANDN U2856 ( .B(n2540), .A(n10738), .Z(n2541) );
  XOR U2857 ( .A(y[3872]), .B(n19762), .Z(n2542) );
  NAND U2858 ( .A(n2542), .B(n2539), .Z(n2543) );
  NAND U2859 ( .A(n2541), .B(n2543), .Z(n2544) );
  ANDN U2860 ( .B(n2544), .A(n19766), .Z(n2545) );
  NANDN U2861 ( .A(x[3874]), .B(n2545), .Z(n2546) );
  ANDN U2862 ( .B(n2546), .A(n10735), .Z(n2547) );
  XNOR U2863 ( .A(n2545), .B(x[3874]), .Z(n2548) );
  NAND U2864 ( .A(n2548), .B(y[3874]), .Z(n2549) );
  NAND U2865 ( .A(n2547), .B(n2549), .Z(n2550) );
  NANDN U2866 ( .A(n19770), .B(n2550), .Z(n2551) );
  NANDN U2867 ( .A(n2551), .B(y[3876]), .Z(n2552) );
  ANDN U2868 ( .B(n2552), .A(n10732), .Z(n2553) );
  XNOR U2869 ( .A(n2551), .B(y[3876]), .Z(n2554) );
  NAND U2870 ( .A(n2554), .B(n10734), .Z(n2555) );
  NAND U2871 ( .A(n2553), .B(n2555), .Z(n10302) );
  NANDN U2872 ( .A(n10714), .B(n10323), .Z(n2556) );
  ANDN U2873 ( .B(n2556), .A(n28327), .Z(n2557) );
  NOR U2874 ( .A(n10712), .B(n10713), .Z(n2558) );
  NANDN U2875 ( .A(n10715), .B(n2557), .Z(n2559) );
  NAND U2876 ( .A(n2558), .B(n2559), .Z(n2560) );
  NOR U2877 ( .A(n28326), .B(n10710), .Z(n2561) );
  NAND U2878 ( .A(n2561), .B(n2560), .Z(n2562) );
  ANDN U2879 ( .B(n2562), .A(n19803), .Z(n2563) );
  NANDN U2880 ( .A(n2563), .B(n10707), .Z(n2564) );
  XOR U2881 ( .A(n2563), .B(y[3894]), .Z(n2565) );
  NAND U2882 ( .A(n2565), .B(x[3894]), .Z(n2566) );
  AND U2883 ( .A(n2564), .B(n2566), .Z(n2567) );
  NOR U2884 ( .A(n19808), .B(n10709), .Z(n2568) );
  OR U2885 ( .A(n20210), .B(n2567), .Z(n2569) );
  AND U2886 ( .A(n2568), .B(n2569), .Z(n2570) );
  NOR U2887 ( .A(n28341), .B(n20211), .Z(n2571) );
  NANDN U2888 ( .A(n2570), .B(n2571), .Z(n2572) );
  ANDN U2889 ( .B(n2572), .A(n10704), .Z(n2573) );
  NANDN U2890 ( .A(n10706), .B(n2573), .Z(n10324) );
  NAND U2891 ( .A(n10330), .B(n10331), .Z(n2574) );
  NOR U2892 ( .A(n10684), .B(n19854), .Z(n2575) );
  OR U2893 ( .A(n10682), .B(n2574), .Z(n2576) );
  AND U2894 ( .A(n2575), .B(n2576), .Z(n2577) );
  NOR U2895 ( .A(n10680), .B(n19853), .Z(n2578) );
  NOR U2896 ( .A(n20205), .B(n10681), .Z(n2579) );
  NANDN U2897 ( .A(n2577), .B(n2579), .Z(n2580) );
  AND U2898 ( .A(n2578), .B(n2580), .Z(n2581) );
  NOR U2899 ( .A(n2581), .B(n20204), .Z(n2582) );
  NANDN U2900 ( .A(n19863), .B(n2582), .Z(n2583) );
  NANDN U2901 ( .A(n19858), .B(n2583), .Z(n2584) );
  NANDN U2902 ( .A(n2584), .B(y[3922]), .Z(n2585) );
  ANDN U2903 ( .B(n2585), .A(n10679), .Z(n2586) );
  XNOR U2904 ( .A(n2584), .B(y[3922]), .Z(n2587) );
  NAND U2905 ( .A(n2587), .B(n19861), .Z(n2588) );
  NAND U2906 ( .A(n2586), .B(n2588), .Z(n2589) );
  NANDN U2907 ( .A(n19865), .B(n2589), .Z(n10333) );
  ANDN U2908 ( .B(n10357), .A(n10653), .Z(n2590) );
  NANDN U2909 ( .A(y[3941]), .B(n10355), .Z(n2591) );
  NAND U2910 ( .A(n2590), .B(n2591), .Z(n2592) );
  AND U2911 ( .A(n10655), .B(n2592), .Z(n2593) );
  NAND U2912 ( .A(n10651), .B(x[3943]), .Z(n2594) );
  ANDN U2913 ( .B(n2594), .A(n10650), .Z(n2595) );
  XOR U2914 ( .A(x[3943]), .B(n10651), .Z(n2596) );
  NAND U2915 ( .A(n2596), .B(n2593), .Z(n2597) );
  NAND U2916 ( .A(n2595), .B(n2597), .Z(n2598) );
  ANDN U2917 ( .B(n28448), .A(n19903), .Z(n2599) );
  NAND U2918 ( .A(n2599), .B(n2598), .Z(n2600) );
  NANDN U2919 ( .A(n10649), .B(n2600), .Z(n2601) );
  ANDN U2920 ( .B(n28447), .A(n10645), .Z(n2602) );
  NANDN U2921 ( .A(n2601), .B(n10648), .Z(n2603) );
  AND U2922 ( .A(n2602), .B(n2603), .Z(n2604) );
  NOR U2923 ( .A(n19911), .B(n10647), .Z(n2605) );
  NANDN U2924 ( .A(n2604), .B(n2605), .Z(n2606) );
  AND U2925 ( .A(n28457), .B(n2606), .Z(n2607) );
  ANDN U2926 ( .B(n2607), .A(n10644), .Z(n10358) );
  NAND U2927 ( .A(n10360), .B(n10624), .Z(n2608) );
  AND U2928 ( .A(n10362), .B(n2608), .Z(n2609) );
  NANDN U2929 ( .A(n19953), .B(n2609), .Z(n2610) );
  NOR U2930 ( .A(n28507), .B(n19949), .Z(n2611) );
  NAND U2931 ( .A(n2611), .B(n2610), .Z(n2612) );
  NANDN U2932 ( .A(n10623), .B(n2612), .Z(n2613) );
  NOR U2933 ( .A(n28514), .B(n28506), .Z(n2614) );
  OR U2934 ( .A(n19952), .B(n2613), .Z(n2615) );
  AND U2935 ( .A(n2614), .B(n2615), .Z(n2616) );
  NOR U2936 ( .A(n10622), .B(n19957), .Z(n2617) );
  NANDN U2937 ( .A(n2616), .B(n2617), .Z(n2618) );
  AND U2938 ( .A(n28513), .B(n2618), .Z(n2619) );
  NAND U2939 ( .A(n10619), .B(x[3973]), .Z(n2620) );
  ANDN U2940 ( .B(n2620), .A(n19966), .Z(n2621) );
  XOR U2941 ( .A(x[3973]), .B(n10619), .Z(n2622) );
  NAND U2942 ( .A(n2622), .B(n2619), .Z(n2623) );
  NAND U2943 ( .A(n2621), .B(n2623), .Z(n2624) );
  NANDN U2944 ( .A(n19963), .B(n2624), .Z(n10364) );
  ANDN U2945 ( .B(n10369), .A(n10601), .Z(n2625) );
  NAND U2946 ( .A(n2625), .B(n10368), .Z(n2626) );
  ANDN U2947 ( .B(n2626), .A(n19999), .Z(n2627) );
  NANDN U2948 ( .A(x[3992]), .B(n2627), .Z(n2628) );
  ANDN U2949 ( .B(n2628), .A(n10600), .Z(n2629) );
  XNOR U2950 ( .A(n2627), .B(x[3992]), .Z(n2630) );
  NAND U2951 ( .A(n2630), .B(y[3992]), .Z(n2631) );
  NAND U2952 ( .A(n2629), .B(n2631), .Z(n2632) );
  AND U2953 ( .A(n20004), .B(n2632), .Z(n2633) );
  NAND U2954 ( .A(n10598), .B(y[3994]), .Z(n2634) );
  ANDN U2955 ( .B(n2634), .A(n10597), .Z(n2635) );
  XOR U2956 ( .A(y[3994]), .B(n10598), .Z(n2636) );
  NAND U2957 ( .A(n2636), .B(n2633), .Z(n2637) );
  NAND U2958 ( .A(n2635), .B(n2637), .Z(n2638) );
  NAND U2959 ( .A(n2638), .B(n20008), .Z(n2639) );
  NANDN U2960 ( .A(y[3996]), .B(x[3996]), .Z(n2640) );
  XNOR U2961 ( .A(y[3996]), .B(x[3996]), .Z(n2641) );
  NAND U2962 ( .A(n2641), .B(n2639), .Z(n2642) );
  NAND U2963 ( .A(n2640), .B(n2642), .Z(n10370) );
  NANDN U2964 ( .A(n10418), .B(x[4015]), .Z(n2643) );
  ANDN U2965 ( .B(n2643), .A(n20039), .Z(n2644) );
  XNOR U2966 ( .A(x[4015]), .B(n10418), .Z(n2645) );
  NAND U2967 ( .A(n2645), .B(n10571), .Z(n2646) );
  NAND U2968 ( .A(n2644), .B(n2646), .Z(n2647) );
  AND U2969 ( .A(n20037), .B(n2647), .Z(n2648) );
  NANDN U2970 ( .A(y[4017]), .B(n2648), .Z(n2649) );
  ANDN U2971 ( .B(n2649), .A(n10569), .Z(n2650) );
  XNOR U2972 ( .A(n2648), .B(y[4017]), .Z(n2651) );
  NAND U2973 ( .A(n2651), .B(x[4017]), .Z(n2652) );
  NAND U2974 ( .A(n2650), .B(n2652), .Z(n2653) );
  ANDN U2975 ( .B(n2653), .A(n20042), .Z(n2654) );
  NAND U2976 ( .A(n10568), .B(x[4019]), .Z(n2655) );
  ANDN U2977 ( .B(n2655), .A(n20049), .Z(n2656) );
  XOR U2978 ( .A(x[4019]), .B(n10568), .Z(n2657) );
  NAND U2979 ( .A(n2657), .B(n2654), .Z(n2658) );
  NAND U2980 ( .A(n2656), .B(n2658), .Z(n2659) );
  NANDN U2981 ( .A(n20046), .B(n2659), .Z(n10419) );
  NAND U2982 ( .A(n20084), .B(n10446), .Z(n2660) );
  NANDN U2983 ( .A(n10447), .B(y[4040]), .Z(n2661) );
  NAND U2984 ( .A(n2660), .B(n2661), .Z(n2662) );
  OR U2985 ( .A(n10550), .B(n2662), .Z(n2663) );
  ANDN U2986 ( .B(n2663), .A(n20088), .Z(n2664) );
  NANDN U2987 ( .A(x[4042]), .B(y[4042]), .Z(n2665) );
  ANDN U2988 ( .B(n2665), .A(n20097), .Z(n2666) );
  XNOR U2989 ( .A(y[4042]), .B(x[4042]), .Z(n2667) );
  NAND U2990 ( .A(n2667), .B(n2664), .Z(n2668) );
  NAND U2991 ( .A(n2666), .B(n2668), .Z(n2669) );
  ANDN U2992 ( .B(n2669), .A(n20092), .Z(n2670) );
  NAND U2993 ( .A(n20095), .B(y[4044]), .Z(n2671) );
  ANDN U2994 ( .B(n2671), .A(n10547), .Z(n2672) );
  XOR U2995 ( .A(y[4044]), .B(n20095), .Z(n2673) );
  NAND U2996 ( .A(n2673), .B(n2670), .Z(n2674) );
  NAND U2997 ( .A(n2672), .B(n2674), .Z(n2675) );
  NANDN U2998 ( .A(n20099), .B(n2675), .Z(n10449) );
  ANDN U2999 ( .B(n10454), .A(n10531), .Z(n2676) );
  NAND U3000 ( .A(n2676), .B(n10453), .Z(n2677) );
  NANDN U3001 ( .A(n20134), .B(n2677), .Z(n2678) );
  NANDN U3002 ( .A(n2678), .B(y[4062]), .Z(n2679) );
  ANDN U3003 ( .B(n2679), .A(n20140), .Z(n2680) );
  XNOR U3004 ( .A(y[4062]), .B(n2678), .Z(n2681) );
  NAND U3005 ( .A(n2681), .B(n10530), .Z(n2682) );
  NAND U3006 ( .A(n2680), .B(n2682), .Z(n2683) );
  NOR U3007 ( .A(n10529), .B(n20143), .Z(n2684) );
  NAND U3008 ( .A(n2684), .B(n2683), .Z(n2685) );
  NAND U3009 ( .A(n2685), .B(n28716), .Z(n2686) );
  NOR U3010 ( .A(n10527), .B(n20142), .Z(n2687) );
  OR U3011 ( .A(n20139), .B(n2686), .Z(n2688) );
  AND U3012 ( .A(n2687), .B(n2688), .Z(n2689) );
  NOR U3013 ( .A(n2689), .B(n28714), .Z(n2690) );
  NANDN U3014 ( .A(n10525), .B(n2690), .Z(n2691) );
  NANDN U3015 ( .A(n20147), .B(n2691), .Z(n10456) );
  NANDN U3016 ( .A(y[4087]), .B(x[4087]), .Z(n28760) );
  IV U3017 ( .A(ebreg), .Z(e) );
  NANDN U3018 ( .A(x[4089]), .B(y[4089]), .Z(n2693) );
  NANDN U3019 ( .A(x[4090]), .B(y[4090]), .Z(n2692) );
  AND U3020 ( .A(n2693), .B(n2692), .Z(n2696) );
  NANDN U3021 ( .A(x[4091]), .B(y[4091]), .Z(n2695) );
  NANDN U3022 ( .A(x[4092]), .B(y[4092]), .Z(n2694) );
  NAND U3023 ( .A(n2695), .B(n2694), .Z(n20183) );
  ANDN U3024 ( .B(n2696), .A(n20183), .Z(n20181) );
  ANDN U3025 ( .B(y[4086]), .A(x[4086]), .Z(n20194) );
  ANDN U3026 ( .B(n20181), .A(n20194), .Z(n2709) );
  NANDN U3027 ( .A(x[4095]), .B(y[4095]), .Z(n20190) );
  NANDN U3028 ( .A(y[4089]), .B(x[4089]), .Z(n2698) );
  NANDN U3029 ( .A(y[4088]), .B(x[4088]), .Z(n2697) );
  AND U3030 ( .A(n2698), .B(n2697), .Z(n2701) );
  NANDN U3031 ( .A(y[4091]), .B(x[4091]), .Z(n2700) );
  NANDN U3032 ( .A(y[4090]), .B(x[4090]), .Z(n2699) );
  NAND U3033 ( .A(n2700), .B(n2699), .Z(n20182) );
  ANDN U3034 ( .B(n2701), .A(n20182), .Z(n2707) );
  NANDN U3035 ( .A(y[4093]), .B(x[4093]), .Z(n2703) );
  NANDN U3036 ( .A(y[4092]), .B(x[4092]), .Z(n2702) );
  NAND U3037 ( .A(n2703), .B(n2702), .Z(n20180) );
  NANDN U3038 ( .A(y[4094]), .B(x[4094]), .Z(n2705) );
  NANDN U3039 ( .A(y[4095]), .B(x[4095]), .Z(n2704) );
  NAND U3040 ( .A(n2705), .B(n2704), .Z(n20189) );
  NOR U3041 ( .A(n20180), .B(n20189), .Z(n2706) );
  NAND U3042 ( .A(n2707), .B(n2706), .Z(n28766) );
  ANDN U3043 ( .B(n20190), .A(n28766), .Z(n2708) );
  AND U3044 ( .A(n2709), .B(n2708), .Z(n2712) );
  IV U3045 ( .A(y[4084]), .Z(n2720) );
  NAND U3046 ( .A(n2720), .B(x[4084]), .Z(n2711) );
  NANDN U3047 ( .A(y[4085]), .B(x[4085]), .Z(n2710) );
  NAND U3048 ( .A(n2711), .B(n2710), .Z(n28756) );
  ANDN U3049 ( .B(n2712), .A(n28756), .Z(n2719) );
  NANDN U3050 ( .A(y[4086]), .B(x[4086]), .Z(n28761) );
  NANDN U3051 ( .A(x[4088]), .B(y[4088]), .Z(n20192) );
  AND U3052 ( .A(n28761), .B(n20192), .Z(n2714) );
  XNOR U3053 ( .A(x[4087]), .B(y[4087]), .Z(n2713) );
  AND U3054 ( .A(n2714), .B(n2713), .Z(n2717) );
  NANDN U3055 ( .A(x[4094]), .B(y[4094]), .Z(n2716) );
  NANDN U3056 ( .A(x[4093]), .B(y[4093]), .Z(n2715) );
  NAND U3057 ( .A(n2716), .B(n2715), .Z(n20187) );
  ANDN U3058 ( .B(n2717), .A(n20187), .Z(n2718) );
  AND U3059 ( .A(n2719), .B(n2718), .Z(n10499) );
  NOR U3060 ( .A(n2720), .B(x[4084]), .Z(n20196) );
  XOR U3061 ( .A(x[4082]), .B(y[4082]), .Z(n20171) );
  IV U3062 ( .A(y[4079]), .Z(n10505) );
  ANDN U3063 ( .B(x[4078]), .A(y[4078]), .Z(n10507) );
  IV U3064 ( .A(y[4077]), .Z(n10508) );
  ANDN U3065 ( .B(x[4076]), .A(y[4076]), .Z(n10510) );
  ANDN U3066 ( .B(x[4073]), .A(y[4073]), .Z(n10516) );
  ANDN U3067 ( .B(y[4073]), .A(x[4073]), .Z(n28734) );
  NANDN U3068 ( .A(x[4072]), .B(y[4072]), .Z(n10518) );
  NANDN U3069 ( .A(n28734), .B(n10518), .Z(n10467) );
  ANDN U3070 ( .B(x[4072]), .A(y[4072]), .Z(n10517) );
  ANDN U3071 ( .B(y[4071]), .A(x[4071]), .Z(n10519) );
  NANDN U3072 ( .A(y[4070]), .B(x[4070]), .Z(n10520) );
  XNOR U3073 ( .A(x[4070]), .B(y[4070]), .Z(n10461) );
  IV U3074 ( .A(x[4068]), .Z(n10524) );
  ANDN U3075 ( .B(x[4067]), .A(y[4067]), .Z(n20147) );
  ANDN U3076 ( .B(y[4067]), .A(x[4067]), .Z(n10525) );
  NANDN U3077 ( .A(x[4065]), .B(y[4065]), .Z(n28716) );
  IV U3078 ( .A(x[4062]), .Z(n10530) );
  ANDN U3079 ( .B(x[4061]), .A(y[4061]), .Z(n20134) );
  ANDN U3080 ( .B(y[4061]), .A(x[4061]), .Z(n10531) );
  ANDN U3081 ( .B(x[4059]), .A(y[4059]), .Z(n20128) );
  ANDN U3082 ( .B(y[4059]), .A(x[4059]), .Z(n20131) );
  IV U3083 ( .A(x[4058]), .Z(n10533) );
  ANDN U3084 ( .B(x[4057]), .A(y[4057]), .Z(n20124) );
  ANDN U3085 ( .B(y[4057]), .A(x[4057]), .Z(n10534) );
  IV U3086 ( .A(x[4056]), .Z(n10536) );
  ANDN U3087 ( .B(x[4055]), .A(y[4055]), .Z(n20120) );
  ANDN U3088 ( .B(y[4055]), .A(x[4055]), .Z(n10537) );
  NANDN U3089 ( .A(x[4054]), .B(y[4054]), .Z(n28689) );
  ANDN U3090 ( .B(x[4053]), .A(y[4053]), .Z(n10540) );
  ANDN U3091 ( .B(y[4052]), .A(x[4052]), .Z(n20201) );
  ANDN U3092 ( .B(x[4047]), .A(y[4047]), .Z(n20103) );
  ANDN U3093 ( .B(y[4047]), .A(x[4047]), .Z(n20106) );
  IV U3094 ( .A(x[4046]), .Z(n10546) );
  ANDN U3095 ( .B(x[4045]), .A(y[4045]), .Z(n20099) );
  ANDN U3096 ( .B(y[4045]), .A(x[4045]), .Z(n10547) );
  IV U3097 ( .A(x[4044]), .Z(n20095) );
  ANDN U3098 ( .B(x[4043]), .A(y[4043]), .Z(n20092) );
  ANDN U3099 ( .B(y[4043]), .A(x[4043]), .Z(n20097) );
  ANDN U3100 ( .B(x[4041]), .A(y[4041]), .Z(n20088) );
  ANDN U3101 ( .B(y[4041]), .A(x[4041]), .Z(n10550) );
  IV U3102 ( .A(x[4040]), .Z(n20084) );
  ANDN U3103 ( .B(x[4039]), .A(y[4039]), .Z(n20081) );
  ANDN U3104 ( .B(y[4039]), .A(x[4039]), .Z(n20086) );
  NANDN U3105 ( .A(x[4037]), .B(y[4037]), .Z(n28657) );
  ANDN U3106 ( .B(y[4033]), .A(x[4033]), .Z(n20069) );
  NANDN U3107 ( .A(y[4031]), .B(x[4031]), .Z(n10440) );
  NANDN U3108 ( .A(y[4030]), .B(x[4030]), .Z(n2721) );
  AND U3109 ( .A(n10440), .B(n2721), .Z(n28638) );
  ANDN U3110 ( .B(y[4029]), .A(x[4029]), .Z(n10555) );
  ANDN U3111 ( .B(x[4027]), .A(y[4027]), .Z(n10559) );
  XOR U3112 ( .A(x[4028]), .B(y[4028]), .Z(n10558) );
  OR U3113 ( .A(n10559), .B(n10558), .Z(n10436) );
  NANDN U3114 ( .A(y[4025]), .B(x[4025]), .Z(n10564) );
  ANDN U3115 ( .B(x[4026]), .A(y[4026]), .Z(n10560) );
  ANDN U3116 ( .B(n10564), .A(n10560), .Z(n10432) );
  XNOR U3117 ( .A(x[4025]), .B(y[4025]), .Z(n10430) );
  ANDN U3118 ( .B(x[4023]), .A(y[4023]), .Z(n20053) );
  ANDN U3119 ( .B(x[4022]), .A(y[4022]), .Z(n20054) );
  ANDN U3120 ( .B(y[4020]), .A(x[4020]), .Z(n20046) );
  ANDN U3121 ( .B(x[4020]), .A(y[4020]), .Z(n20049) );
  IV U3122 ( .A(y[4019]), .Z(n10568) );
  ANDN U3123 ( .B(y[4018]), .A(x[4018]), .Z(n20042) );
  ANDN U3124 ( .B(x[4018]), .A(y[4018]), .Z(n10569) );
  ANDN U3125 ( .B(x[4016]), .A(y[4016]), .Z(n20039) );
  IV U3126 ( .A(y[4015]), .Z(n10571) );
  ANDN U3127 ( .B(x[4014]), .A(y[4014]), .Z(n10573) );
  ANDN U3128 ( .B(x[4012]), .A(y[4012]), .Z(n10577) );
  ANDN U3129 ( .B(y[4011]), .A(x[4011]), .Z(n20031) );
  NANDN U3130 ( .A(y[4010]), .B(x[4010]), .Z(n10578) );
  XNOR U3131 ( .A(x[4010]), .B(y[4010]), .Z(n10406) );
  NANDN U3132 ( .A(x[4006]), .B(y[4006]), .Z(n2723) );
  NANDN U3133 ( .A(x[4005]), .B(y[4005]), .Z(n2722) );
  AND U3134 ( .A(n2723), .B(n2722), .Z(n28584) );
  ANDN U3135 ( .B(y[4004]), .A(x[4004]), .Z(n10583) );
  ANDN U3136 ( .B(x[4003]), .A(y[4003]), .Z(n10585) );
  ANDN U3137 ( .B(y[4001]), .A(x[4001]), .Z(n10587) );
  IV U3138 ( .A(x[4000]), .Z(n10588) );
  ANDN U3139 ( .B(y[3999]), .A(x[3999]), .Z(n10590) );
  IV U3140 ( .A(x[3998]), .Z(n10591) );
  ANDN U3141 ( .B(y[3997]), .A(x[3997]), .Z(n10593) );
  ANDN U3142 ( .B(y[3995]), .A(x[3995]), .Z(n10597) );
  IV U3143 ( .A(x[3994]), .Z(n10598) );
  ANDN U3144 ( .B(y[3993]), .A(x[3993]), .Z(n10600) );
  ANDN U3145 ( .B(x[3991]), .A(y[3991]), .Z(n19999) );
  ANDN U3146 ( .B(y[3991]), .A(x[3991]), .Z(n10601) );
  NANDN U3147 ( .A(y[3989]), .B(x[3989]), .Z(n19996) );
  ANDN U3148 ( .B(y[3989]), .A(x[3989]), .Z(n10604) );
  ANDN U3149 ( .B(x[3987]), .A(y[3987]), .Z(n10606) );
  ANDN U3150 ( .B(x[3988]), .A(y[3988]), .Z(n19995) );
  NANDN U3151 ( .A(y[3985]), .B(x[3985]), .Z(n19986) );
  ANDN U3152 ( .B(x[3986]), .A(y[3986]), .Z(n10605) );
  ANDN U3153 ( .B(x[3983]), .A(y[3983]), .Z(n10610) );
  ANDN U3154 ( .B(x[3984]), .A(y[3984]), .Z(n19985) );
  ANDN U3155 ( .B(x[3981]), .A(y[3981]), .Z(n10612) );
  ANDN U3156 ( .B(x[3980]), .A(y[3980]), .Z(n10613) );
  ANDN U3157 ( .B(y[3978]), .A(x[3978]), .Z(n19973) );
  ANDN U3158 ( .B(x[3978]), .A(y[3978]), .Z(n10614) );
  IV U3159 ( .A(y[3977]), .Z(n10616) );
  ANDN U3160 ( .B(y[3976]), .A(x[3976]), .Z(n19969) );
  ANDN U3161 ( .B(x[3976]), .A(y[3976]), .Z(n10617) );
  ANDN U3162 ( .B(y[3974]), .A(x[3974]), .Z(n19963) );
  ANDN U3163 ( .B(x[3974]), .A(y[3974]), .Z(n19966) );
  IV U3164 ( .A(y[3973]), .Z(n10619) );
  ANDN U3165 ( .B(x[3971]), .A(y[3971]), .Z(n19957) );
  ANDN U3166 ( .B(y[3970]), .A(x[3970]), .Z(n28506) );
  ANDN U3167 ( .B(x[3969]), .A(y[3969]), .Z(n19952) );
  IV U3168 ( .A(y[3967]), .Z(n10624) );
  ANDN U3169 ( .B(y[3966]), .A(x[3966]), .Z(n19945) );
  ANDN U3170 ( .B(x[3966]), .A(y[3966]), .Z(n10625) );
  ANDN U3171 ( .B(x[3964]), .A(y[3964]), .Z(n19942) );
  ANDN U3172 ( .B(y[3960]), .A(x[3960]), .Z(n28484) );
  ANDN U3173 ( .B(x[3959]), .A(y[3959]), .Z(n10635) );
  ANDN U3174 ( .B(y[3959]), .A(x[3959]), .Z(n28486) );
  NANDN U3175 ( .A(x[3958]), .B(y[3958]), .Z(n28478) );
  ANDN U3176 ( .B(y[3956]), .A(x[3956]), .Z(n19926) );
  ANDN U3177 ( .B(x[3956]), .A(y[3956]), .Z(n10637) );
  ANDN U3178 ( .B(y[3955]), .A(x[3955]), .Z(n19927) );
  NANDN U3179 ( .A(x[3951]), .B(y[3951]), .Z(n28465) );
  NANDN U3180 ( .A(x[3949]), .B(y[3949]), .Z(n28457) );
  ANDN U3181 ( .B(x[3947]), .A(y[3947]), .Z(n10647) );
  ANDN U3182 ( .B(x[3948]), .A(y[3948]), .Z(n19911) );
  ANDN U3183 ( .B(x[3945]), .A(y[3945]), .Z(n10649) );
  ANDN U3184 ( .B(x[3944]), .A(y[3944]), .Z(n10650) );
  ANDN U3185 ( .B(x[3942]), .A(y[3942]), .Z(n10653) );
  ANDN U3186 ( .B(x[3940]), .A(y[3940]), .Z(n10657) );
  IV U3187 ( .A(y[3939]), .Z(n10658) );
  ANDN U3188 ( .B(x[3938]), .A(y[3938]), .Z(n10660) );
  IV U3189 ( .A(y[3937]), .Z(n10661) );
  ANDN U3190 ( .B(x[3936]), .A(y[3936]), .Z(n10663) );
  ANDN U3191 ( .B(y[3932]), .A(x[3932]), .Z(n20202) );
  ANDN U3192 ( .B(x[3931]), .A(y[3931]), .Z(n10671) );
  ANDN U3193 ( .B(y[3931]), .A(x[3931]), .Z(n20203) );
  NANDN U3194 ( .A(x[3930]), .B(y[3930]), .Z(n10673) );
  ANDN U3195 ( .B(y[3929]), .A(x[3929]), .Z(n10674) );
  ANDN U3196 ( .B(y[3928]), .A(x[3928]), .Z(n28408) );
  ANDN U3197 ( .B(x[3927]), .A(y[3927]), .Z(n19873) );
  ANDN U3198 ( .B(y[3926]), .A(x[3926]), .Z(n19870) );
  ANDN U3199 ( .B(x[3923]), .A(y[3923]), .Z(n19865) );
  ANDN U3200 ( .B(y[3923]), .A(x[3923]), .Z(n10679) );
  IV U3201 ( .A(x[3922]), .Z(n19861) );
  ANDN U3202 ( .B(x[3921]), .A(y[3921]), .Z(n19858) );
  ANDN U3203 ( .B(y[3921]), .A(x[3921]), .Z(n19863) );
  IV U3204 ( .A(x[3916]), .Z(n19847) );
  ANDN U3205 ( .B(x[3915]), .A(y[3915]), .Z(n19844) );
  ANDN U3206 ( .B(y[3915]), .A(x[3915]), .Z(n19849) );
  ANDN U3207 ( .B(x[3913]), .A(y[3913]), .Z(n19839) );
  ANDN U3208 ( .B(y[3912]), .A(x[3912]), .Z(n10686) );
  NANDN U3209 ( .A(x[3909]), .B(y[3909]), .Z(n28371) );
  NANDN U3210 ( .A(x[3907]), .B(y[3907]), .Z(n20209) );
  ANDN U3211 ( .B(x[3905]), .A(y[3905]), .Z(n10696) );
  ANDN U3212 ( .B(x[3906]), .A(y[3906]), .Z(n19829) );
  ANDN U3213 ( .B(x[3903]), .A(y[3903]), .Z(n19821) );
  ANDN U3214 ( .B(x[3902]), .A(y[3902]), .Z(n19822) );
  ANDN U3215 ( .B(x[3899]), .A(y[3899]), .Z(n10702) );
  NANDN U3216 ( .A(x[3899]), .B(y[3899]), .Z(n28348) );
  ANDN U3217 ( .B(y[3898]), .A(x[3898]), .Z(n28340) );
  ANDN U3218 ( .B(n28348), .A(n28340), .Z(n10325) );
  ANDN U3219 ( .B(x[3897]), .A(y[3897]), .Z(n10706) );
  ANDN U3220 ( .B(y[3896]), .A(x[3896]), .Z(n20211) );
  ANDN U3221 ( .B(x[3895]), .A(y[3895]), .Z(n10709) );
  ANDN U3222 ( .B(y[3895]), .A(x[3895]), .Z(n20210) );
  ANDN U3223 ( .B(y[3892]), .A(x[3892]), .Z(n28326) );
  ANDN U3224 ( .B(y[3893]), .A(x[3893]), .Z(n10710) );
  ANDN U3225 ( .B(y[3890]), .A(x[3890]), .Z(n10715) );
  ANDN U3226 ( .B(y[3891]), .A(x[3891]), .Z(n28327) );
  ANDN U3227 ( .B(x[3890]), .A(y[3890]), .Z(n10714) );
  ANDN U3228 ( .B(y[3889]), .A(x[3889]), .Z(n10716) );
  IV U3229 ( .A(x[3888]), .Z(n10719) );
  ANDN U3230 ( .B(y[3887]), .A(x[3887]), .Z(n10721) );
  ANDN U3231 ( .B(y[3885]), .A(x[3885]), .Z(n10725) );
  IV U3232 ( .A(x[3884]), .Z(n10726) );
  ANDN U3233 ( .B(y[3883]), .A(x[3883]), .Z(n10728) );
  ANDN U3234 ( .B(x[3881]), .A(y[3881]), .Z(n19784) );
  ANDN U3235 ( .B(y[3881]), .A(x[3881]), .Z(n10729) );
  ANDN U3236 ( .B(x[3879]), .A(y[3879]), .Z(n19778) );
  ANDN U3237 ( .B(y[3879]), .A(x[3879]), .Z(n19781) );
  IV U3238 ( .A(x[3878]), .Z(n10731) );
  ANDN U3239 ( .B(x[3877]), .A(y[3877]), .Z(n19774) );
  ANDN U3240 ( .B(y[3877]), .A(x[3877]), .Z(n10732) );
  IV U3241 ( .A(x[3876]), .Z(n10734) );
  ANDN U3242 ( .B(x[3875]), .A(y[3875]), .Z(n19770) );
  ANDN U3243 ( .B(y[3875]), .A(x[3875]), .Z(n10735) );
  ANDN U3244 ( .B(x[3873]), .A(y[3873]), .Z(n19766) );
  ANDN U3245 ( .B(y[3873]), .A(x[3873]), .Z(n10738) );
  IV U3246 ( .A(x[3872]), .Z(n19762) );
  ANDN U3247 ( .B(x[3871]), .A(y[3871]), .Z(n19759) );
  IV U3248 ( .A(n19759), .Z(n10301) );
  ANDN U3249 ( .B(y[3871]), .A(x[3871]), .Z(n19764) );
  ANDN U3250 ( .B(x[3869]), .A(y[3869]), .Z(n10739) );
  ANDN U3251 ( .B(y[3869]), .A(x[3869]), .Z(n19757) );
  IV U3252 ( .A(x[3868]), .Z(n10741) );
  ANDN U3253 ( .B(x[3867]), .A(y[3867]), .Z(n19751) );
  ANDN U3254 ( .B(y[3867]), .A(x[3867]), .Z(n10743) );
  ANDN U3255 ( .B(x[3865]), .A(y[3865]), .Z(n10746) );
  IV U3256 ( .A(n10746), .Z(n10299) );
  ANDN U3257 ( .B(y[3865]), .A(x[3865]), .Z(n10745) );
  IV U3258 ( .A(x[3864]), .Z(n10748) );
  ANDN U3259 ( .B(x[3863]), .A(y[3863]), .Z(n10751) );
  ANDN U3260 ( .B(y[3863]), .A(x[3863]), .Z(n10750) );
  IV U3261 ( .A(x[3858]), .Z(n10758) );
  ANDN U3262 ( .B(x[3857]), .A(y[3857]), .Z(n10761) );
  ANDN U3263 ( .B(y[3857]), .A(x[3857]), .Z(n10760) );
  IV U3264 ( .A(x[3856]), .Z(n10763) );
  ANDN U3265 ( .B(x[3855]), .A(y[3855]), .Z(n19734) );
  ANDN U3266 ( .B(y[3855]), .A(x[3855]), .Z(n10765) );
  ANDN U3267 ( .B(x[3853]), .A(y[3853]), .Z(n10768) );
  ANDN U3268 ( .B(y[3853]), .A(x[3853]), .Z(n10767) );
  ANDN U3269 ( .B(x[3851]), .A(y[3851]), .Z(n10770) );
  XOR U3270 ( .A(x[3852]), .B(y[3852]), .Z(n19729) );
  NANDN U3271 ( .A(y[3849]), .B(x[3849]), .Z(n10774) );
  ANDN U3272 ( .B(x[3850]), .A(y[3850]), .Z(n10771) );
  ANDN U3273 ( .B(n10774), .A(n10771), .Z(n10292) );
  XNOR U3274 ( .A(x[3849]), .B(y[3849]), .Z(n10290) );
  NANDN U3275 ( .A(y[3847]), .B(x[3847]), .Z(n19722) );
  ANDN U3276 ( .B(x[3848]), .A(y[3848]), .Z(n10775) );
  ANDN U3277 ( .B(n19722), .A(n10775), .Z(n10287) );
  XNOR U3278 ( .A(x[3847]), .B(y[3847]), .Z(n10285) );
  ANDN U3279 ( .B(x[3846]), .A(y[3846]), .Z(n19723) );
  ANDN U3280 ( .B(y[3845]), .A(x[3845]), .Z(n10778) );
  NANDN U3281 ( .A(y[3845]), .B(x[3845]), .Z(n2725) );
  NANDN U3282 ( .A(y[3844]), .B(x[3844]), .Z(n2724) );
  NAND U3283 ( .A(n2725), .B(n2724), .Z(n28228) );
  ANDN U3284 ( .B(x[3841]), .A(y[3841]), .Z(n19714) );
  ANDN U3285 ( .B(y[3841]), .A(x[3841]), .Z(n10783) );
  IV U3286 ( .A(x[3840]), .Z(n19710) );
  NANDN U3287 ( .A(y[3839]), .B(x[3839]), .Z(n19708) );
  ANDN U3288 ( .B(y[3839]), .A(x[3839]), .Z(n19712) );
  ANDN U3289 ( .B(x[3837]), .A(y[3837]), .Z(n10785) );
  ANDN U3290 ( .B(x[3838]), .A(y[3838]), .Z(n19707) );
  NANDN U3291 ( .A(y[3835]), .B(x[3835]), .Z(n19698) );
  ANDN U3292 ( .B(x[3836]), .A(y[3836]), .Z(n10784) );
  ANDN U3293 ( .B(x[3833]), .A(y[3833]), .Z(n10787) );
  ANDN U3294 ( .B(x[3834]), .A(y[3834]), .Z(n19697) );
  ANDN U3295 ( .B(x[3831]), .A(y[3831]), .Z(n10789) );
  ANDN U3296 ( .B(x[3830]), .A(y[3830]), .Z(n10790) );
  ANDN U3297 ( .B(x[3827]), .A(y[3827]), .Z(n10796) );
  ANDN U3298 ( .B(y[3827]), .A(x[3827]), .Z(n20212) );
  NANDN U3299 ( .A(x[3826]), .B(y[3826]), .Z(n10798) );
  ANDN U3300 ( .B(x[3826]), .A(y[3826]), .Z(n10797) );
  ANDN U3301 ( .B(y[3824]), .A(x[3824]), .Z(n28182) );
  ANDN U3302 ( .B(x[3823]), .A(y[3823]), .Z(n10803) );
  NANDN U3303 ( .A(x[3823]), .B(y[3823]), .Z(n28183) );
  ANDN U3304 ( .B(y[3822]), .A(x[3822]), .Z(n28176) );
  ANDN U3305 ( .B(n28183), .A(n28176), .Z(n10263) );
  NANDN U3306 ( .A(x[3819]), .B(y[3819]), .Z(n28172) );
  IV U3307 ( .A(x[3816]), .Z(n10809) );
  ANDN U3308 ( .B(x[3815]), .A(y[3815]), .Z(n19662) );
  ANDN U3309 ( .B(y[3815]), .A(x[3815]), .Z(n10811) );
  NANDN U3310 ( .A(x[3814]), .B(y[3814]), .Z(n28156) );
  ANDN U3311 ( .B(x[3813]), .A(y[3813]), .Z(n19657) );
  ANDN U3312 ( .B(y[3812]), .A(x[3812]), .Z(n10813) );
  NANDN U3313 ( .A(x[3813]), .B(y[3813]), .Z(n28158) );
  ANDN U3314 ( .B(x[3812]), .A(y[3812]), .Z(n19658) );
  ANDN U3315 ( .B(y[3811]), .A(x[3811]), .Z(n10814) );
  ANDN U3316 ( .B(x[3805]), .A(y[3805]), .Z(n19645) );
  ANDN U3317 ( .B(y[3805]), .A(x[3805]), .Z(n10820) );
  ANDN U3318 ( .B(x[3803]), .A(y[3803]), .Z(n10823) );
  ANDN U3319 ( .B(y[3803]), .A(x[3803]), .Z(n10822) );
  IV U3320 ( .A(x[3802]), .Z(n10825) );
  ANDN U3321 ( .B(x[3801]), .A(y[3801]), .Z(n19639) );
  ANDN U3322 ( .B(y[3801]), .A(x[3801]), .Z(n10827) );
  IV U3323 ( .A(x[3800]), .Z(n10828) );
  ANDN U3324 ( .B(x[3799]), .A(y[3799]), .Z(n19635) );
  ANDN U3325 ( .B(y[3799]), .A(x[3799]), .Z(n10829) );
  ANDN U3326 ( .B(x[3797]), .A(y[3797]), .Z(n19631) );
  ANDN U3327 ( .B(y[3797]), .A(x[3797]), .Z(n10832) );
  ANDN U3328 ( .B(x[3795]), .A(y[3795]), .Z(n10833) );
  XNOR U3329 ( .A(x[3796]), .B(y[3796]), .Z(n19629) );
  ANDN U3330 ( .B(y[3794]), .A(x[3794]), .Z(n20215) );
  NANDN U3331 ( .A(x[3795]), .B(y[3795]), .Z(n28119) );
  IV U3332 ( .A(x[3790]), .Z(n10840) );
  ANDN U3333 ( .B(y[3789]), .A(x[3789]), .Z(n10842) );
  ANDN U3334 ( .B(x[3787]), .A(y[3787]), .Z(n19612) );
  ANDN U3335 ( .B(y[3787]), .A(x[3787]), .Z(n10843) );
  ANDN U3336 ( .B(x[3785]), .A(y[3785]), .Z(n19608) );
  ANDN U3337 ( .B(y[3785]), .A(x[3785]), .Z(n10846) );
  IV U3338 ( .A(x[3784]), .Z(n19604) );
  ANDN U3339 ( .B(x[3783]), .A(y[3783]), .Z(n19601) );
  ANDN U3340 ( .B(y[3783]), .A(x[3783]), .Z(n19606) );
  IV U3341 ( .A(x[3782]), .Z(n10847) );
  ANDN U3342 ( .B(x[3781]), .A(y[3781]), .Z(n19597) );
  ANDN U3343 ( .B(y[3781]), .A(x[3781]), .Z(n10848) );
  ANDN U3344 ( .B(x[3779]), .A(y[3779]), .Z(n19593) );
  IV U3345 ( .A(n19593), .Z(n10231) );
  ANDN U3346 ( .B(y[3779]), .A(x[3779]), .Z(n10851) );
  NANDN U3347 ( .A(x[3778]), .B(y[3778]), .Z(n28081) );
  ANDN U3348 ( .B(x[3777]), .A(y[3777]), .Z(n19588) );
  ANDN U3349 ( .B(y[3776]), .A(x[3776]), .Z(n19585) );
  ANDN U3350 ( .B(x[3773]), .A(y[3773]), .Z(n19580) );
  ANDN U3351 ( .B(y[3773]), .A(x[3773]), .Z(n10856) );
  NANDN U3352 ( .A(x[3772]), .B(y[3772]), .Z(n28066) );
  NANDN U3353 ( .A(x[3771]), .B(y[3771]), .Z(n28068) );
  ANDN U3354 ( .B(x[3769]), .A(y[3769]), .Z(n10861) );
  ANDN U3355 ( .B(x[3770]), .A(y[3770]), .Z(n19576) );
  NANDN U3356 ( .A(y[3767]), .B(x[3767]), .Z(n19568) );
  ANDN U3357 ( .B(x[3768]), .A(y[3768]), .Z(n10860) );
  ANDN U3358 ( .B(x[3765]), .A(y[3765]), .Z(n10863) );
  ANDN U3359 ( .B(x[3766]), .A(y[3766]), .Z(n19567) );
  ANDN U3360 ( .B(x[3763]), .A(y[3763]), .Z(n10865) );
  ANDN U3361 ( .B(x[3762]), .A(y[3762]), .Z(n10866) );
  ANDN U3362 ( .B(y[3760]), .A(x[3760]), .Z(n10869) );
  ANDN U3363 ( .B(x[3760]), .A(y[3760]), .Z(n10868) );
  IV U3364 ( .A(y[3759]), .Z(n10871) );
  ANDN U3365 ( .B(y[3758]), .A(x[3758]), .Z(n19551) );
  ANDN U3366 ( .B(x[3758]), .A(y[3758]), .Z(n10873) );
  IV U3367 ( .A(y[3757]), .Z(n10874) );
  ANDN U3368 ( .B(y[3756]), .A(x[3756]), .Z(n19547) );
  IV U3369 ( .A(n19547), .Z(n10225) );
  ANDN U3370 ( .B(x[3756]), .A(y[3756]), .Z(n10875) );
  ANDN U3371 ( .B(y[3754]), .A(x[3754]), .Z(n19541) );
  ANDN U3372 ( .B(x[3754]), .A(y[3754]), .Z(n19544) );
  IV U3373 ( .A(y[3753]), .Z(n10877) );
  ANDN U3374 ( .B(y[3752]), .A(x[3752]), .Z(n19538) );
  ANDN U3375 ( .B(x[3752]), .A(y[3752]), .Z(n10878) );
  ANDN U3376 ( .B(y[3748]), .A(x[3748]), .Z(n28016) );
  ANDN U3377 ( .B(x[3747]), .A(y[3747]), .Z(n10881) );
  NANDN U3378 ( .A(x[3747]), .B(y[3747]), .Z(n28017) );
  ANDN U3379 ( .B(y[3746]), .A(x[3746]), .Z(n20218) );
  ANDN U3380 ( .B(x[3741]), .A(y[3741]), .Z(n10887) );
  ANDN U3381 ( .B(y[3741]), .A(x[3741]), .Z(n10886) );
  ANDN U3382 ( .B(y[3735]), .A(x[3735]), .Z(n10894) );
  IV U3383 ( .A(x[3734]), .Z(n10895) );
  ANDN U3384 ( .B(x[3733]), .A(y[3733]), .Z(n10898) );
  ANDN U3385 ( .B(y[3733]), .A(x[3733]), .Z(n10897) );
  IV U3386 ( .A(x[3732]), .Z(n10900) );
  ANDN U3387 ( .B(x[3731]), .A(y[3731]), .Z(n19495) );
  ANDN U3388 ( .B(y[3731]), .A(x[3731]), .Z(n10902) );
  ANDN U3389 ( .B(x[3729]), .A(y[3729]), .Z(n10905) );
  ANDN U3390 ( .B(y[3729]), .A(x[3729]), .Z(n10904) );
  NANDN U3391 ( .A(x[3728]), .B(y[3728]), .Z(n27975) );
  ANDN U3392 ( .B(x[3727]), .A(y[3727]), .Z(n19488) );
  ANDN U3393 ( .B(y[3726]), .A(x[3726]), .Z(n27968) );
  ANDN U3394 ( .B(x[3721]), .A(y[3721]), .Z(n19475) );
  ANDN U3395 ( .B(y[3721]), .A(x[3721]), .Z(n10912) );
  ANDN U3396 ( .B(x[3719]), .A(y[3719]), .Z(n19470) );
  ANDN U3397 ( .B(y[3718]), .A(x[3718]), .Z(n10914) );
  ANDN U3398 ( .B(x[3715]), .A(y[3715]), .Z(n19464) );
  ANDN U3399 ( .B(y[3715]), .A(x[3715]), .Z(n10919) );
  IV U3400 ( .A(x[3714]), .Z(n19460) );
  ANDN U3401 ( .B(x[3713]), .A(y[3713]), .Z(n19457) );
  ANDN U3402 ( .B(y[3713]), .A(x[3713]), .Z(n19462) );
  IV U3403 ( .A(x[3708]), .Z(n19444) );
  ANDN U3404 ( .B(x[3707]), .A(y[3707]), .Z(n19441) );
  ANDN U3405 ( .B(y[3707]), .A(x[3707]), .Z(n19446) );
  IV U3406 ( .A(x[3706]), .Z(n19437) );
  ANDN U3407 ( .B(x[3705]), .A(y[3705]), .Z(n19434) );
  ANDN U3408 ( .B(y[3705]), .A(x[3705]), .Z(n19439) );
  ANDN U3409 ( .B(x[3703]), .A(y[3703]), .Z(n19428) );
  ANDN U3410 ( .B(y[3703]), .A(x[3703]), .Z(n19431) );
  IV U3411 ( .A(x[3702]), .Z(n19424) );
  ANDN U3412 ( .B(x[3701]), .A(y[3701]), .Z(n19421) );
  ANDN U3413 ( .B(y[3701]), .A(x[3701]), .Z(n19426) );
  NANDN U3414 ( .A(x[3700]), .B(y[3700]), .Z(n27911) );
  ANDN U3415 ( .B(x[3699]), .A(y[3699]), .Z(n10923) );
  ANDN U3416 ( .B(y[3698]), .A(x[3698]), .Z(n10925) );
  ANDN U3417 ( .B(x[3695]), .A(y[3695]), .Z(n19409) );
  ANDN U3418 ( .B(y[3695]), .A(x[3695]), .Z(n10928) );
  ANDN U3419 ( .B(y[3693]), .A(x[3693]), .Z(n10930) );
  ANDN U3420 ( .B(y[3691]), .A(x[3691]), .Z(n10934) );
  IV U3421 ( .A(x[3690]), .Z(n10935) );
  ANDN U3422 ( .B(x[3689]), .A(y[3689]), .Z(n19399) );
  ANDN U3423 ( .B(y[3689]), .A(x[3689]), .Z(n10937) );
  ANDN U3424 ( .B(x[3687]), .A(y[3687]), .Z(n19395) );
  ANDN U3425 ( .B(y[3687]), .A(x[3687]), .Z(n10939) );
  IV U3426 ( .A(x[3686]), .Z(n19391) );
  ANDN U3427 ( .B(x[3685]), .A(y[3685]), .Z(n19388) );
  ANDN U3428 ( .B(y[3685]), .A(x[3685]), .Z(n19393) );
  ANDN U3429 ( .B(y[3683]), .A(x[3683]), .Z(n10941) );
  ANDN U3430 ( .B(y[3681]), .A(x[3681]), .Z(n10945) );
  IV U3431 ( .A(x[3680]), .Z(n10946) );
  ANDN U3432 ( .B(x[3679]), .A(y[3679]), .Z(n19378) );
  ANDN U3433 ( .B(y[3679]), .A(x[3679]), .Z(n10948) );
  ANDN U3434 ( .B(x[3677]), .A(y[3677]), .Z(n19374) );
  ANDN U3435 ( .B(y[3677]), .A(x[3677]), .Z(n10950) );
  IV U3436 ( .A(x[3676]), .Z(n19370) );
  ANDN U3437 ( .B(x[3675]), .A(y[3675]), .Z(n19367) );
  ANDN U3438 ( .B(y[3675]), .A(x[3675]), .Z(n19372) );
  ANDN U3439 ( .B(y[3673]), .A(x[3673]), .Z(n10952) );
  ANDN U3440 ( .B(y[3671]), .A(x[3671]), .Z(n10956) );
  IV U3441 ( .A(x[3670]), .Z(n10957) );
  NANDN U3442 ( .A(y[3669]), .B(x[3669]), .Z(n19358) );
  ANDN U3443 ( .B(y[3669]), .A(x[3669]), .Z(n10959) );
  ANDN U3444 ( .B(x[3667]), .A(y[3667]), .Z(n10963) );
  ANDN U3445 ( .B(x[3668]), .A(y[3668]), .Z(n19357) );
  NANDN U3446 ( .A(y[3665]), .B(x[3665]), .Z(n10965) );
  ANDN U3447 ( .B(x[3666]), .A(y[3666]), .Z(n10962) );
  XNOR U3448 ( .A(x[3665]), .B(y[3665]), .Z(n10207) );
  IV U3449 ( .A(x[3664]), .Z(n19348) );
  NAND U3450 ( .A(n19348), .B(y[3664]), .Z(n27836) );
  NANDN U3451 ( .A(x[3663]), .B(y[3663]), .Z(n27838) );
  ANDN U3452 ( .B(x[3662]), .A(y[3662]), .Z(n10967) );
  ANDN U3453 ( .B(y[3661]), .A(x[3661]), .Z(n10969) );
  NANDN U3454 ( .A(y[3661]), .B(x[3661]), .Z(n2727) );
  NANDN U3455 ( .A(y[3660]), .B(x[3660]), .Z(n2726) );
  NAND U3456 ( .A(n2727), .B(n2726), .Z(n27830) );
  ANDN U3457 ( .B(y[3660]), .A(x[3660]), .Z(n10971) );
  ANDN U3458 ( .B(y[3658]), .A(x[3658]), .Z(n27822) );
  ANDN U3459 ( .B(x[3657]), .A(y[3657]), .Z(n10974) );
  XNOR U3460 ( .A(x[3658]), .B(y[3658]), .Z(n19341) );
  NANDN U3461 ( .A(x[3657]), .B(y[3657]), .Z(n27823) );
  NANDN U3462 ( .A(x[3656]), .B(y[3656]), .Z(n19335) );
  NAND U3463 ( .A(n27823), .B(n19335), .Z(n10190) );
  ANDN U3464 ( .B(y[3655]), .A(x[3655]), .Z(n19336) );
  ANDN U3465 ( .B(y[3654]), .A(x[3654]), .Z(n27812) );
  ANDN U3466 ( .B(x[3653]), .A(y[3653]), .Z(n10976) );
  XNOR U3467 ( .A(x[3654]), .B(y[3654]), .Z(n19331) );
  ANDN U3468 ( .B(y[3652]), .A(x[3652]), .Z(n27806) );
  NANDN U3469 ( .A(x[3653]), .B(y[3653]), .Z(n27814) );
  NANDN U3470 ( .A(x[3651]), .B(y[3651]), .Z(n27807) );
  ANDN U3471 ( .B(x[3649]), .A(y[3649]), .Z(n10983) );
  ANDN U3472 ( .B(x[3650]), .A(y[3650]), .Z(n10979) );
  NANDN U3473 ( .A(y[3647]), .B(x[3647]), .Z(n19317) );
  ANDN U3474 ( .B(x[3648]), .A(y[3648]), .Z(n10982) );
  ANDN U3475 ( .B(x[3645]), .A(y[3645]), .Z(n10985) );
  ANDN U3476 ( .B(x[3646]), .A(y[3646]), .Z(n19316) );
  ANDN U3477 ( .B(x[3643]), .A(y[3643]), .Z(n10986) );
  ANDN U3478 ( .B(x[3642]), .A(y[3642]), .Z(n10987) );
  ANDN U3479 ( .B(y[3640]), .A(x[3640]), .Z(n19303) );
  ANDN U3480 ( .B(x[3640]), .A(y[3640]), .Z(n10991) );
  ANDN U3481 ( .B(y[3638]), .A(x[3638]), .Z(n10994) );
  ANDN U3482 ( .B(x[3638]), .A(y[3638]), .Z(n10993) );
  IV U3483 ( .A(y[3637]), .Z(n10996) );
  ANDN U3484 ( .B(y[3636]), .A(x[3636]), .Z(n19298) );
  ANDN U3485 ( .B(x[3636]), .A(y[3636]), .Z(n10998) );
  ANDN U3486 ( .B(y[3632]), .A(x[3632]), .Z(n20222) );
  ANDN U3487 ( .B(x[3631]), .A(y[3631]), .Z(n19284) );
  XNOR U3488 ( .A(x[3632]), .B(y[3632]), .Z(n19288) );
  ANDN U3489 ( .B(y[3630]), .A(x[3630]), .Z(n19282) );
  NANDN U3490 ( .A(x[3631]), .B(y[3631]), .Z(n20223) );
  ANDN U3491 ( .B(y[3629]), .A(x[3629]), .Z(n19281) );
  ANDN U3492 ( .B(y[3628]), .A(x[3628]), .Z(n27754) );
  ANDN U3493 ( .B(x[3627]), .A(y[3627]), .Z(n11002) );
  ANDN U3494 ( .B(y[3626]), .A(x[3626]), .Z(n11004) );
  ANDN U3495 ( .B(x[3625]), .A(y[3625]), .Z(n11007) );
  ANDN U3496 ( .B(x[3626]), .A(y[3626]), .Z(n11003) );
  NANDN U3497 ( .A(y[3623]), .B(x[3623]), .Z(n19268) );
  ANDN U3498 ( .B(x[3624]), .A(y[3624]), .Z(n11006) );
  XNOR U3499 ( .A(x[3623]), .B(y[3623]), .Z(n10180) );
  ANDN U3500 ( .B(x[3621]), .A(y[3621]), .Z(n11009) );
  ANDN U3501 ( .B(x[3622]), .A(y[3622]), .Z(n19267) );
  ANDN U3502 ( .B(x[3619]), .A(y[3619]), .Z(n19257) );
  ANDN U3503 ( .B(x[3618]), .A(y[3618]), .Z(n19258) );
  ANDN U3504 ( .B(y[3616]), .A(x[3616]), .Z(n19252) );
  ANDN U3505 ( .B(x[3616]), .A(y[3616]), .Z(n11013) );
  ANDN U3506 ( .B(y[3614]), .A(x[3614]), .Z(n19248) );
  ANDN U3507 ( .B(x[3614]), .A(y[3614]), .Z(n11016) );
  ANDN U3508 ( .B(y[3612]), .A(x[3612]), .Z(n11019) );
  ANDN U3509 ( .B(x[3612]), .A(y[3612]), .Z(n11018) );
  IV U3510 ( .A(y[3611]), .Z(n11021) );
  ANDN U3511 ( .B(y[3610]), .A(x[3610]), .Z(n19242) );
  ANDN U3512 ( .B(x[3610]), .A(y[3610]), .Z(n11023) );
  ANDN U3513 ( .B(y[3608]), .A(x[3608]), .Z(n19237) );
  ANDN U3514 ( .B(x[3608]), .A(y[3608]), .Z(n19239) );
  XNOR U3515 ( .A(x[3606]), .B(y[3606]), .Z(n19233) );
  ANDN U3516 ( .B(y[3604]), .A(x[3604]), .Z(n27700) );
  NANDN U3517 ( .A(x[3605]), .B(y[3605]), .Z(n27708) );
  ANDN U3518 ( .B(x[3603]), .A(y[3603]), .Z(n11027) );
  ANDN U3519 ( .B(y[3603]), .A(x[3603]), .Z(n27701) );
  NANDN U3520 ( .A(x[3602]), .B(y[3602]), .Z(n11029) );
  ANDN U3521 ( .B(y[3601]), .A(x[3601]), .Z(n11030) );
  ANDN U3522 ( .B(y[3600]), .A(x[3600]), .Z(n27690) );
  ANDN U3523 ( .B(x[3599]), .A(y[3599]), .Z(n11031) );
  XNOR U3524 ( .A(x[3600]), .B(y[3600]), .Z(n19220) );
  ANDN U3525 ( .B(y[3598]), .A(x[3598]), .Z(n27684) );
  NANDN U3526 ( .A(x[3599]), .B(y[3599]), .Z(n27692) );
  IV U3527 ( .A(x[3594]), .Z(n19207) );
  ANDN U3528 ( .B(x[3593]), .A(y[3593]), .Z(n19204) );
  ANDN U3529 ( .B(y[3593]), .A(x[3593]), .Z(n19209) );
  ANDN U3530 ( .B(y[3591]), .A(x[3591]), .Z(n11039) );
  ANDN U3531 ( .B(x[3589]), .A(y[3589]), .Z(n11044) );
  ANDN U3532 ( .B(y[3589]), .A(x[3589]), .Z(n11043) );
  ANDN U3533 ( .B(x[3587]), .A(y[3587]), .Z(n19195) );
  ANDN U3534 ( .B(y[3586]), .A(x[3586]), .Z(n11047) );
  NANDN U3535 ( .A(y[3579]), .B(x[3579]), .Z(n11059) );
  ANDN U3536 ( .B(y[3579]), .A(x[3579]), .Z(n11057) );
  ANDN U3537 ( .B(x[3577]), .A(y[3577]), .Z(n11063) );
  ANDN U3538 ( .B(x[3578]), .A(y[3578]), .Z(n11058) );
  NANDN U3539 ( .A(y[3575]), .B(x[3575]), .Z(n19177) );
  ANDN U3540 ( .B(x[3576]), .A(y[3576]), .Z(n11062) );
  XNOR U3541 ( .A(x[3575]), .B(y[3575]), .Z(n10166) );
  ANDN U3542 ( .B(x[3573]), .A(y[3573]), .Z(n11065) );
  ANDN U3543 ( .B(x[3574]), .A(y[3574]), .Z(n19176) );
  ANDN U3544 ( .B(x[3571]), .A(y[3571]), .Z(n11067) );
  ANDN U3545 ( .B(x[3570]), .A(y[3570]), .Z(n11068) );
  ANDN U3546 ( .B(x[3568]), .A(y[3568]), .Z(n11072) );
  IV U3547 ( .A(y[3567]), .Z(n11073) );
  ANDN U3548 ( .B(y[3566]), .A(x[3566]), .Z(n19161) );
  ANDN U3549 ( .B(x[3566]), .A(y[3566]), .Z(n11075) );
  ANDN U3550 ( .B(y[3562]), .A(x[3562]), .Z(n27604) );
  ANDN U3551 ( .B(x[3561]), .A(y[3561]), .Z(n19149) );
  XNOR U3552 ( .A(x[3562]), .B(y[3562]), .Z(n19153) );
  NANDN U3553 ( .A(x[3561]), .B(y[3561]), .Z(n27605) );
  ANDN U3554 ( .B(y[3560]), .A(x[3560]), .Z(n20224) );
  NANDN U3555 ( .A(x[3559]), .B(y[3559]), .Z(n20225) );
  IV U3556 ( .A(x[3556]), .Z(n11086) );
  ANDN U3557 ( .B(x[3555]), .A(y[3555]), .Z(n19139) );
  ANDN U3558 ( .B(y[3555]), .A(x[3555]), .Z(n11088) );
  ANDN U3559 ( .B(x[3553]), .A(y[3553]), .Z(n19135) );
  ANDN U3560 ( .B(y[3553]), .A(x[3553]), .Z(n11090) );
  IV U3561 ( .A(x[3552]), .Z(n11091) );
  ANDN U3562 ( .B(x[3551]), .A(y[3551]), .Z(n19131) );
  IV U3563 ( .A(n19131), .Z(n10160) );
  ANDN U3564 ( .B(y[3551]), .A(x[3551]), .Z(n11092) );
  ANDN U3565 ( .B(y[3549]), .A(x[3549]), .Z(n11095) );
  ANDN U3566 ( .B(x[3547]), .A(y[3547]), .Z(n11100) );
  ANDN U3567 ( .B(y[3547]), .A(x[3547]), .Z(n11099) );
  IV U3568 ( .A(x[3546]), .Z(n11102) );
  ANDN U3569 ( .B(x[3545]), .A(y[3545]), .Z(n19123) );
  ANDN U3570 ( .B(y[3545]), .A(x[3545]), .Z(n11104) );
  ANDN U3571 ( .B(x[3543]), .A(y[3543]), .Z(n19119) );
  ANDN U3572 ( .B(y[3543]), .A(x[3543]), .Z(n11106) );
  IV U3573 ( .A(x[3542]), .Z(n11107) );
  NAND U3574 ( .A(n11107), .B(y[3542]), .Z(n27562) );
  NANDN U3575 ( .A(x[3541]), .B(y[3541]), .Z(n27564) );
  IV U3576 ( .A(x[3538]), .Z(n11112) );
  ANDN U3577 ( .B(x[3537]), .A(y[3537]), .Z(n19107) );
  ANDN U3578 ( .B(y[3537]), .A(x[3537]), .Z(n11114) );
  ANDN U3579 ( .B(x[3535]), .A(y[3535]), .Z(n19103) );
  ANDN U3580 ( .B(y[3535]), .A(x[3535]), .Z(n11116) );
  IV U3581 ( .A(x[3534]), .Z(n19099) );
  ANDN U3582 ( .B(x[3533]), .A(y[3533]), .Z(n19096) );
  ANDN U3583 ( .B(y[3533]), .A(x[3533]), .Z(n19101) );
  ANDN U3584 ( .B(x[3531]), .A(y[3531]), .Z(n19091) );
  XNOR U3585 ( .A(x[3532]), .B(y[3532]), .Z(n19094) );
  ANDN U3586 ( .B(y[3530]), .A(x[3530]), .Z(n11117) );
  NANDN U3587 ( .A(x[3531]), .B(y[3531]), .Z(n27541) );
  ANDN U3588 ( .B(x[3527]), .A(y[3527]), .Z(n19084) );
  ANDN U3589 ( .B(y[3527]), .A(x[3527]), .Z(n11122) );
  IV U3590 ( .A(x[3526]), .Z(n19080) );
  ANDN U3591 ( .B(x[3525]), .A(y[3525]), .Z(n19077) );
  ANDN U3592 ( .B(y[3525]), .A(x[3525]), .Z(n19082) );
  NANDN U3593 ( .A(x[3523]), .B(y[3523]), .Z(n27523) );
  ANDN U3594 ( .B(x[3519]), .A(y[3519]), .Z(n19065) );
  ANDN U3595 ( .B(y[3519]), .A(x[3519]), .Z(n11128) );
  IV U3596 ( .A(x[3518]), .Z(n19061) );
  ANDN U3597 ( .B(x[3517]), .A(y[3517]), .Z(n19058) );
  ANDN U3598 ( .B(y[3517]), .A(x[3517]), .Z(n19063) );
  ANDN U3599 ( .B(y[3515]), .A(x[3515]), .Z(n11130) );
  ANDN U3600 ( .B(y[3513]), .A(x[3513]), .Z(n11134) );
  IV U3601 ( .A(x[3512]), .Z(n11135) );
  ANDN U3602 ( .B(x[3511]), .A(y[3511]), .Z(n19048) );
  ANDN U3603 ( .B(y[3511]), .A(x[3511]), .Z(n11137) );
  NANDN U3604 ( .A(y[3509]), .B(x[3509]), .Z(n19045) );
  ANDN U3605 ( .B(y[3509]), .A(x[3509]), .Z(n11139) );
  ANDN U3606 ( .B(x[3507]), .A(y[3507]), .Z(n11141) );
  ANDN U3607 ( .B(x[3508]), .A(y[3508]), .Z(n19044) );
  NANDN U3608 ( .A(y[3505]), .B(x[3505]), .Z(n11143) );
  ANDN U3609 ( .B(x[3506]), .A(y[3506]), .Z(n11140) );
  ANDN U3610 ( .B(x[3503]), .A(y[3503]), .Z(n11146) );
  NANDN U3611 ( .A(y[3504]), .B(x[3504]), .Z(n11142) );
  ANDN U3612 ( .B(x[3501]), .A(y[3501]), .Z(n11149) );
  ANDN U3613 ( .B(x[3500]), .A(y[3500]), .Z(n11150) );
  ANDN U3614 ( .B(x[3498]), .A(y[3498]), .Z(n11154) );
  IV U3615 ( .A(y[3497]), .Z(n11155) );
  ANDN U3616 ( .B(y[3496]), .A(x[3496]), .Z(n19022) );
  ANDN U3617 ( .B(x[3496]), .A(y[3496]), .Z(n11157) );
  ANDN U3618 ( .B(y[3494]), .A(x[3494]), .Z(n19019) );
  ANDN U3619 ( .B(x[3494]), .A(y[3494]), .Z(n11159) );
  ANDN U3620 ( .B(y[3493]), .A(x[3493]), .Z(n19018) );
  NANDN U3621 ( .A(x[3490]), .B(y[3490]), .Z(n2729) );
  NANDN U3622 ( .A(x[3489]), .B(y[3489]), .Z(n2728) );
  AND U3623 ( .A(n2729), .B(n2728), .Z(n27452) );
  ANDN U3624 ( .B(y[3488]), .A(x[3488]), .Z(n11161) );
  ANDN U3625 ( .B(x[3487]), .A(y[3487]), .Z(n11163) );
  ANDN U3626 ( .B(y[3485]), .A(x[3485]), .Z(n11165) );
  IV U3627 ( .A(x[3484]), .Z(n11166) );
  ANDN U3628 ( .B(x[3483]), .A(y[3483]), .Z(n19003) );
  ANDN U3629 ( .B(y[3483]), .A(x[3483]), .Z(n11168) );
  ANDN U3630 ( .B(x[3481]), .A(y[3481]), .Z(n18999) );
  ANDN U3631 ( .B(y[3481]), .A(x[3481]), .Z(n11170) );
  IV U3632 ( .A(x[3480]), .Z(n18995) );
  ANDN U3633 ( .B(x[3479]), .A(y[3479]), .Z(n18992) );
  ANDN U3634 ( .B(y[3478]), .A(x[3478]), .Z(n27426) );
  ANDN U3635 ( .B(x[3477]), .A(y[3477]), .Z(n18987) );
  XNOR U3636 ( .A(x[3478]), .B(y[3478]), .Z(n18990) );
  NANDN U3637 ( .A(y[3473]), .B(x[3473]), .Z(n11177) );
  ANDN U3638 ( .B(x[3474]), .A(y[3474]), .Z(n11173) );
  NANDN U3639 ( .A(y[3471]), .B(x[3471]), .Z(n11179) );
  ANDN U3640 ( .B(x[3472]), .A(y[3472]), .Z(n11178) );
  ANDN U3641 ( .B(n11179), .A(n11178), .Z(n10139) );
  IV U3642 ( .A(x[3470]), .Z(n18974) );
  NAND U3643 ( .A(n18974), .B(y[3470]), .Z(n27408) );
  NANDN U3644 ( .A(x[3469]), .B(y[3469]), .Z(n27410) );
  NANDN U3645 ( .A(x[3468]), .B(y[3468]), .Z(n11181) );
  ANDN U3646 ( .B(y[3466]), .A(x[3466]), .Z(n18966) );
  NANDN U3647 ( .A(x[3464]), .B(y[3464]), .Z(n18960) );
  ANDN U3648 ( .B(y[3465]), .A(x[3465]), .Z(n18965) );
  XNOR U3649 ( .A(y[3464]), .B(x[3464]), .Z(n10137) );
  ANDN U3650 ( .B(y[3462]), .A(x[3462]), .Z(n11188) );
  NANDN U3651 ( .A(x[3460]), .B(y[3460]), .Z(n11190) );
  ANDN U3652 ( .B(y[3461]), .A(x[3461]), .Z(n11187) );
  ANDN U3653 ( .B(y[3458]), .A(x[3458]), .Z(n11192) );
  NANDN U3654 ( .A(x[3456]), .B(y[3456]), .Z(n18944) );
  ANDN U3655 ( .B(y[3457]), .A(x[3457]), .Z(n11191) );
  XNOR U3656 ( .A(y[3456]), .B(x[3456]), .Z(n10134) );
  ANDN U3657 ( .B(y[3454]), .A(x[3454]), .Z(n18940) );
  NANDN U3658 ( .A(x[3452]), .B(y[3452]), .Z(n11196) );
  ANDN U3659 ( .B(y[3453]), .A(x[3453]), .Z(n18939) );
  ANDN U3660 ( .B(y[3450]), .A(x[3450]), .Z(n11198) );
  NANDN U3661 ( .A(x[3448]), .B(y[3448]), .Z(n11200) );
  ANDN U3662 ( .B(y[3449]), .A(x[3449]), .Z(n11197) );
  XNOR U3663 ( .A(y[3448]), .B(x[3448]), .Z(n10132) );
  ANDN U3664 ( .B(y[3446]), .A(x[3446]), .Z(n18924) );
  NANDN U3665 ( .A(x[3444]), .B(y[3444]), .Z(n18918) );
  ANDN U3666 ( .B(y[3445]), .A(x[3445]), .Z(n18923) );
  ANDN U3667 ( .B(y[3442]), .A(x[3442]), .Z(n11206) );
  NANDN U3668 ( .A(x[3440]), .B(y[3440]), .Z(n11208) );
  ANDN U3669 ( .B(y[3441]), .A(x[3441]), .Z(n11205) );
  XNOR U3670 ( .A(y[3440]), .B(x[3440]), .Z(n10129) );
  ANDN U3671 ( .B(y[3438]), .A(x[3438]), .Z(n11210) );
  NANDN U3672 ( .A(x[3436]), .B(y[3436]), .Z(n18902) );
  ANDN U3673 ( .B(y[3437]), .A(x[3437]), .Z(n11209) );
  NANDN U3674 ( .A(x[3434]), .B(y[3434]), .Z(n18898) );
  ANDN U3675 ( .B(y[3435]), .A(x[3435]), .Z(n18901) );
  IV U3676 ( .A(y[3433]), .Z(n11213) );
  NANDN U3677 ( .A(x[3431]), .B(y[3431]), .Z(n20227) );
  NANDN U3678 ( .A(y[3429]), .B(x[3429]), .Z(n11219) );
  ANDN U3679 ( .B(x[3430]), .A(y[3430]), .Z(n18891) );
  ANDN U3680 ( .B(n11219), .A(n18891), .Z(n10121) );
  XNOR U3681 ( .A(x[3429]), .B(y[3429]), .Z(n10119) );
  XNOR U3682 ( .A(x[3427]), .B(y[3427]), .Z(n10112) );
  ANDN U3683 ( .B(x[3425]), .A(y[3425]), .Z(n18880) );
  NANDN U3684 ( .A(x[3424]), .B(y[3424]), .Z(n11226) );
  ANDN U3685 ( .B(y[3425]), .A(x[3425]), .Z(n11223) );
  ANDN U3686 ( .B(x[3419]), .A(y[3419]), .Z(n18870) );
  NANDN U3687 ( .A(x[3418]), .B(y[3418]), .Z(n18868) );
  ANDN U3688 ( .B(y[3419]), .A(x[3419]), .Z(n11233) );
  ANDN U3689 ( .B(x[3415]), .A(y[3415]), .Z(n18862) );
  NANDN U3690 ( .A(x[3414]), .B(y[3414]), .Z(n11240) );
  ANDN U3691 ( .B(y[3415]), .A(x[3415]), .Z(n11237) );
  ANDN U3692 ( .B(y[3412]), .A(x[3412]), .Z(n18855) );
  NANDN U3693 ( .A(y[3411]), .B(x[3411]), .Z(n11242) );
  ANDN U3694 ( .B(x[3412]), .A(y[3412]), .Z(n18858) );
  IV U3695 ( .A(x[3410]), .Z(n11243) );
  NAND U3696 ( .A(n11243), .B(y[3410]), .Z(n27286) );
  ANDN U3697 ( .B(x[3409]), .A(y[3409]), .Z(n11245) );
  NANDN U3698 ( .A(y[3407]), .B(x[3407]), .Z(n11248) );
  ANDN U3699 ( .B(x[3408]), .A(y[3408]), .Z(n11246) );
  ANDN U3700 ( .B(x[3405]), .A(y[3405]), .Z(n11252) );
  NANDN U3701 ( .A(y[3403]), .B(x[3403]), .Z(n18840) );
  ANDN U3702 ( .B(x[3404]), .A(y[3404]), .Z(n11251) );
  ANDN U3703 ( .B(x[3401]), .A(y[3401]), .Z(n11256) );
  NANDN U3704 ( .A(y[3399]), .B(x[3399]), .Z(n11258) );
  ANDN U3705 ( .B(x[3400]), .A(y[3400]), .Z(n11255) );
  XNOR U3706 ( .A(y[3398]), .B(x[3398]), .Z(n10100) );
  ANDN U3707 ( .B(x[3397]), .A(y[3397]), .Z(n11260) );
  NANDN U3708 ( .A(y[3395]), .B(x[3395]), .Z(n11263) );
  ANDN U3709 ( .B(x[3396]), .A(y[3396]), .Z(n11259) );
  ANDN U3710 ( .B(x[3393]), .A(y[3393]), .Z(n18824) );
  NANDN U3711 ( .A(y[3391]), .B(x[3391]), .Z(n11268) );
  ANDN U3712 ( .B(x[3392]), .A(y[3392]), .Z(n18823) );
  NANDN U3713 ( .A(x[3386]), .B(y[3386]), .Z(n11271) );
  ANDN U3714 ( .B(y[3387]), .A(x[3387]), .Z(n11270) );
  ANDN U3715 ( .B(y[3383]), .A(x[3383]), .Z(n11275) );
  NANDN U3716 ( .A(y[3383]), .B(x[3383]), .Z(n2731) );
  NANDN U3717 ( .A(y[3382]), .B(x[3382]), .Z(n2730) );
  AND U3718 ( .A(n2731), .B(n2730), .Z(n27230) );
  NANDN U3719 ( .A(x[3381]), .B(y[3381]), .Z(n11276) );
  ANDN U3720 ( .B(y[3382]), .A(x[3382]), .Z(n11277) );
  ANDN U3721 ( .B(n11276), .A(n11277), .Z(n10096) );
  XNOR U3722 ( .A(y[3381]), .B(x[3381]), .Z(n10094) );
  XNOR U3723 ( .A(y[3376]), .B(x[3376]), .Z(n10079) );
  ANDN U3724 ( .B(x[3375]), .A(y[3375]), .Z(n11286) );
  NANDN U3725 ( .A(y[3373]), .B(x[3373]), .Z(n11288) );
  ANDN U3726 ( .B(x[3374]), .A(y[3374]), .Z(n11285) );
  ANDN U3727 ( .B(n11288), .A(n11285), .Z(n10073) );
  ANDN U3728 ( .B(x[3371]), .A(y[3371]), .Z(n11292) );
  NANDN U3729 ( .A(y[3369]), .B(x[3369]), .Z(n18782) );
  ANDN U3730 ( .B(x[3370]), .A(y[3370]), .Z(n11291) );
  NANDN U3731 ( .A(y[3367]), .B(x[3367]), .Z(n11296) );
  ANDN U3732 ( .B(x[3368]), .A(y[3368]), .Z(n18781) );
  XNOR U3733 ( .A(y[3366]), .B(x[3366]), .Z(n18777) );
  ANDN U3734 ( .B(y[3364]), .A(x[3364]), .Z(n11297) );
  ANDN U3735 ( .B(x[3364]), .A(y[3364]), .Z(n18774) );
  NANDN U3736 ( .A(x[3362]), .B(y[3362]), .Z(n11301) );
  ANDN U3737 ( .B(y[3363]), .A(x[3363]), .Z(n11298) );
  ANDN U3738 ( .B(x[3357]), .A(y[3357]), .Z(n18756) );
  XNOR U3739 ( .A(x[3358]), .B(y[3358]), .Z(n18760) );
  ANDN U3740 ( .B(y[3356]), .A(x[3356]), .Z(n27170) );
  NANDN U3741 ( .A(x[3357]), .B(y[3357]), .Z(n27178) );
  NANDN U3742 ( .A(x[3355]), .B(y[3355]), .Z(n27172) );
  NANDN U3743 ( .A(x[3354]), .B(y[3354]), .Z(n11305) );
  ANDN U3744 ( .B(y[3352]), .A(x[3352]), .Z(n11308) );
  NANDN U3745 ( .A(x[3350]), .B(y[3350]), .Z(n11312) );
  ANDN U3746 ( .B(y[3351]), .A(x[3351]), .Z(n11307) );
  ANDN U3747 ( .B(y[3348]), .A(x[3348]), .Z(n18740) );
  NANDN U3748 ( .A(x[3346]), .B(y[3346]), .Z(n11316) );
  ANDN U3749 ( .B(y[3347]), .A(x[3347]), .Z(n18739) );
  ANDN U3750 ( .B(y[3344]), .A(x[3344]), .Z(n11320) );
  NANDN U3751 ( .A(x[3342]), .B(y[3342]), .Z(n18728) );
  ANDN U3752 ( .B(y[3343]), .A(x[3343]), .Z(n11319) );
  XNOR U3753 ( .A(y[3342]), .B(x[3342]), .Z(n10067) );
  ANDN U3754 ( .B(y[3341]), .A(x[3341]), .Z(n18727) );
  ANDN U3755 ( .B(y[3340]), .A(x[3340]), .Z(n27137) );
  ANDN U3756 ( .B(x[3339]), .A(y[3339]), .Z(n11323) );
  ANDN U3757 ( .B(y[3338]), .A(x[3338]), .Z(n11326) );
  ANDN U3758 ( .B(x[3338]), .A(y[3338]), .Z(n11324) );
  NANDN U3759 ( .A(x[3337]), .B(y[3337]), .Z(n11325) );
  NANDN U3760 ( .A(y[3335]), .B(x[3335]), .Z(n2733) );
  NANDN U3761 ( .A(y[3334]), .B(x[3334]), .Z(n2732) );
  NAND U3762 ( .A(n2733), .B(n2732), .Z(n27126) );
  NANDN U3763 ( .A(y[3331]), .B(x[3331]), .Z(n11331) );
  NANDN U3764 ( .A(y[3333]), .B(x[3333]), .Z(n10062) );
  NANDN U3765 ( .A(y[3332]), .B(x[3332]), .Z(n2734) );
  NAND U3766 ( .A(n10062), .B(n2734), .Z(n27122) );
  XNOR U3767 ( .A(x[3331]), .B(y[3331]), .Z(n10059) );
  ANDN U3768 ( .B(x[3329]), .A(y[3329]), .Z(n18711) );
  NANDN U3769 ( .A(y[3327]), .B(x[3327]), .Z(n11336) );
  ANDN U3770 ( .B(x[3328]), .A(y[3328]), .Z(n18710) );
  NANDN U3771 ( .A(x[3322]), .B(y[3322]), .Z(n18694) );
  ANDN U3772 ( .B(y[3323]), .A(x[3323]), .Z(n18701) );
  XNOR U3773 ( .A(y[3322]), .B(x[3322]), .Z(n10055) );
  NANDN U3774 ( .A(x[3320]), .B(y[3320]), .Z(n20228) );
  ANDN U3775 ( .B(y[3321]), .A(x[3321]), .Z(n18695) );
  ANDN U3776 ( .B(n20228), .A(n18695), .Z(n10052) );
  ANDN U3777 ( .B(x[3319]), .A(y[3319]), .Z(n11344) );
  XNOR U3778 ( .A(x[3320]), .B(y[3320]), .Z(n11342) );
  XNOR U3779 ( .A(x[3317]), .B(y[3317]), .Z(n10042) );
  ANDN U3780 ( .B(x[3315]), .A(y[3315]), .Z(n18682) );
  IV U3781 ( .A(n18682), .Z(n10036) );
  NANDN U3782 ( .A(x[3314]), .B(y[3314]), .Z(n11351) );
  ANDN U3783 ( .B(y[3315]), .A(x[3315]), .Z(n11348) );
  ANDN U3784 ( .B(x[3309]), .A(y[3309]), .Z(n18672) );
  NANDN U3785 ( .A(x[3308]), .B(y[3308]), .Z(n18670) );
  ANDN U3786 ( .B(y[3309]), .A(x[3309]), .Z(n11358) );
  ANDN U3787 ( .B(x[3303]), .A(y[3303]), .Z(n18662) );
  NANDN U3788 ( .A(x[3302]), .B(y[3302]), .Z(n11368) );
  ANDN U3789 ( .B(y[3303]), .A(x[3303]), .Z(n11367) );
  ANDN U3790 ( .B(x[3297]), .A(y[3297]), .Z(n18652) );
  NANDN U3791 ( .A(x[3296]), .B(y[3296]), .Z(n11378) );
  ANDN U3792 ( .B(y[3297]), .A(x[3297]), .Z(n18655) );
  ANDN U3793 ( .B(x[3291]), .A(y[3291]), .Z(n11385) );
  NANDN U3794 ( .A(x[3290]), .B(y[3290]), .Z(n11388) );
  ANDN U3795 ( .B(y[3291]), .A(x[3291]), .Z(n11384) );
  ANDN U3796 ( .B(x[3285]), .A(y[3285]), .Z(n18634) );
  NANDN U3797 ( .A(x[3284]), .B(y[3284]), .Z(n11397) );
  ANDN U3798 ( .B(y[3285]), .A(x[3285]), .Z(n11394) );
  ANDN U3799 ( .B(x[3279]), .A(y[3279]), .Z(n18624) );
  NANDN U3800 ( .A(x[3278]), .B(y[3278]), .Z(n18622) );
  ANDN U3801 ( .B(y[3279]), .A(x[3279]), .Z(n11404) );
  ANDN U3802 ( .B(x[3275]), .A(y[3275]), .Z(n18616) );
  NANDN U3803 ( .A(x[3274]), .B(y[3274]), .Z(n11411) );
  ANDN U3804 ( .B(y[3275]), .A(x[3275]), .Z(n11408) );
  ANDN U3805 ( .B(y[3272]), .A(x[3272]), .Z(n18609) );
  NANDN U3806 ( .A(y[3271]), .B(x[3271]), .Z(n11413) );
  ANDN U3807 ( .B(x[3272]), .A(y[3272]), .Z(n18612) );
  ANDN U3808 ( .B(x[3269]), .A(y[3269]), .Z(n18602) );
  XNOR U3809 ( .A(x[3270]), .B(y[3270]), .Z(n18606) );
  NANDN U3810 ( .A(y[3265]), .B(x[3265]), .Z(n2736) );
  NANDN U3811 ( .A(y[3264]), .B(x[3264]), .Z(n2735) );
  AND U3812 ( .A(n2736), .B(n2735), .Z(n26984) );
  NANDN U3813 ( .A(x[3263]), .B(y[3263]), .Z(n18595) );
  ANDN U3814 ( .B(y[3264]), .A(x[3264]), .Z(n18596) );
  NANDN U3815 ( .A(y[3261]), .B(x[3261]), .Z(n2738) );
  NANDN U3816 ( .A(y[3260]), .B(x[3260]), .Z(n2737) );
  NAND U3817 ( .A(n2738), .B(n2737), .Z(n26977) );
  ANDN U3818 ( .B(x[3257]), .A(y[3257]), .Z(n11422) );
  NANDN U3819 ( .A(y[3255]), .B(x[3255]), .Z(n11426) );
  ANDN U3820 ( .B(x[3256]), .A(y[3256]), .Z(n11421) );
  XNOR U3821 ( .A(y[3254]), .B(x[3254]), .Z(n10017) );
  ANDN U3822 ( .B(x[3253]), .A(y[3253]), .Z(n18581) );
  NANDN U3823 ( .A(y[3251]), .B(x[3251]), .Z(n11430) );
  ANDN U3824 ( .B(x[3252]), .A(y[3252]), .Z(n18580) );
  ANDN U3825 ( .B(x[3249]), .A(y[3249]), .Z(n11434) );
  NANDN U3826 ( .A(y[3247]), .B(x[3247]), .Z(n11436) );
  ANDN U3827 ( .B(x[3248]), .A(y[3248]), .Z(n11433) );
  ANDN U3828 ( .B(x[3245]), .A(y[3245]), .Z(n11440) );
  NANDN U3829 ( .A(y[3243]), .B(x[3243]), .Z(n18563) );
  ANDN U3830 ( .B(x[3244]), .A(y[3244]), .Z(n11439) );
  ANDN U3831 ( .B(x[3241]), .A(y[3241]), .Z(n11444) );
  NANDN U3832 ( .A(y[3239]), .B(x[3239]), .Z(n11446) );
  ANDN U3833 ( .B(x[3240]), .A(y[3240]), .Z(n11443) );
  XNOR U3834 ( .A(x[3239]), .B(y[3239]), .Z(n10014) );
  ANDN U3835 ( .B(x[3237]), .A(y[3237]), .Z(n11448) );
  NANDN U3836 ( .A(y[3235]), .B(x[3235]), .Z(n11452) );
  ANDN U3837 ( .B(x[3236]), .A(y[3236]), .Z(n11447) );
  ANDN U3838 ( .B(x[3233]), .A(y[3233]), .Z(n18547) );
  NANDN U3839 ( .A(y[3231]), .B(x[3231]), .Z(n11456) );
  ANDN U3840 ( .B(x[3232]), .A(y[3232]), .Z(n18546) );
  XNOR U3841 ( .A(x[3231]), .B(y[3231]), .Z(n10011) );
  ANDN U3842 ( .B(x[3229]), .A(y[3229]), .Z(n11460) );
  NANDN U3843 ( .A(y[3227]), .B(x[3227]), .Z(n11462) );
  ANDN U3844 ( .B(x[3228]), .A(y[3228]), .Z(n11459) );
  ANDN U3845 ( .B(x[3225]), .A(y[3225]), .Z(n11466) );
  NANDN U3846 ( .A(y[3223]), .B(x[3223]), .Z(n18529) );
  ANDN U3847 ( .B(x[3224]), .A(y[3224]), .Z(n11465) );
  XNOR U3848 ( .A(x[3223]), .B(y[3223]), .Z(n10008) );
  ANDN U3849 ( .B(x[3221]), .A(y[3221]), .Z(n11470) );
  NANDN U3850 ( .A(y[3219]), .B(x[3219]), .Z(n11472) );
  ANDN U3851 ( .B(x[3220]), .A(y[3220]), .Z(n11469) );
  ANDN U3852 ( .B(x[3217]), .A(y[3217]), .Z(n11474) );
  NANDN U3853 ( .A(y[3215]), .B(x[3215]), .Z(n11478) );
  ANDN U3854 ( .B(x[3216]), .A(y[3216]), .Z(n11473) );
  XNOR U3855 ( .A(x[3215]), .B(y[3215]), .Z(n10005) );
  ANDN U3856 ( .B(x[3213]), .A(y[3213]), .Z(n18513) );
  NANDN U3857 ( .A(y[3211]), .B(x[3211]), .Z(n11482) );
  ANDN U3858 ( .B(x[3212]), .A(y[3212]), .Z(n18512) );
  ANDN U3859 ( .B(x[3209]), .A(y[3209]), .Z(n11486) );
  NANDN U3860 ( .A(y[3207]), .B(x[3207]), .Z(n11488) );
  ANDN U3861 ( .B(x[3208]), .A(y[3208]), .Z(n11485) );
  XNOR U3862 ( .A(x[3207]), .B(y[3207]), .Z(n10002) );
  ANDN U3863 ( .B(x[3205]), .A(y[3205]), .Z(n11492) );
  NANDN U3864 ( .A(y[3203]), .B(x[3203]), .Z(n18495) );
  ANDN U3865 ( .B(x[3204]), .A(y[3204]), .Z(n11491) );
  ANDN U3866 ( .B(x[3201]), .A(y[3201]), .Z(n11496) );
  NANDN U3867 ( .A(y[3199]), .B(x[3199]), .Z(n11498) );
  ANDN U3868 ( .B(x[3200]), .A(y[3200]), .Z(n11495) );
  XNOR U3869 ( .A(x[3199]), .B(y[3199]), .Z(n9999) );
  ANDN U3870 ( .B(x[3197]), .A(y[3197]), .Z(n11500) );
  NANDN U3871 ( .A(y[3195]), .B(x[3195]), .Z(n11504) );
  ANDN U3872 ( .B(x[3196]), .A(y[3196]), .Z(n11499) );
  ANDN U3873 ( .B(x[3193]), .A(y[3193]), .Z(n18479) );
  NANDN U3874 ( .A(y[3191]), .B(x[3191]), .Z(n11508) );
  ANDN U3875 ( .B(x[3192]), .A(y[3192]), .Z(n18478) );
  XNOR U3876 ( .A(x[3191]), .B(y[3191]), .Z(n9996) );
  ANDN U3877 ( .B(x[3189]), .A(y[3189]), .Z(n11512) );
  NANDN U3878 ( .A(y[3187]), .B(x[3187]), .Z(n11514) );
  ANDN U3879 ( .B(x[3188]), .A(y[3188]), .Z(n11511) );
  ANDN U3880 ( .B(x[3185]), .A(y[3185]), .Z(n11518) );
  NANDN U3881 ( .A(y[3183]), .B(x[3183]), .Z(n18461) );
  ANDN U3882 ( .B(x[3184]), .A(y[3184]), .Z(n11517) );
  XNOR U3883 ( .A(x[3183]), .B(y[3183]), .Z(n9993) );
  ANDN U3884 ( .B(x[3181]), .A(y[3181]), .Z(n11522) );
  NANDN U3885 ( .A(y[3179]), .B(x[3179]), .Z(n11524) );
  ANDN U3886 ( .B(x[3180]), .A(y[3180]), .Z(n11521) );
  ANDN U3887 ( .B(x[3177]), .A(y[3177]), .Z(n11526) );
  NANDN U3888 ( .A(y[3175]), .B(x[3175]), .Z(n11527) );
  ANDN U3889 ( .B(x[3176]), .A(y[3176]), .Z(n11525) );
  XNOR U3890 ( .A(x[3175]), .B(y[3175]), .Z(n9991) );
  NANDN U3891 ( .A(x[3170]), .B(y[3170]), .Z(n18436) );
  ANDN U3892 ( .B(y[3171]), .A(x[3171]), .Z(n11532) );
  ANDN U3893 ( .B(y[3168]), .A(x[3168]), .Z(n11536) );
  NANDN U3894 ( .A(x[3166]), .B(y[3166]), .Z(n11538) );
  ANDN U3895 ( .B(y[3167]), .A(x[3167]), .Z(n11535) );
  ANDN U3896 ( .B(y[3164]), .A(x[3164]), .Z(n11540) );
  NANDN U3897 ( .A(x[3162]), .B(y[3162]), .Z(n11544) );
  ANDN U3898 ( .B(y[3163]), .A(x[3163]), .Z(n11539) );
  ANDN U3899 ( .B(y[3160]), .A(x[3160]), .Z(n18420) );
  NANDN U3900 ( .A(x[3158]), .B(y[3158]), .Z(n11548) );
  ANDN U3901 ( .B(y[3159]), .A(x[3159]), .Z(n18419) );
  ANDN U3902 ( .B(n11548), .A(n18419), .Z(n9986) );
  NANDN U3903 ( .A(x[3156]), .B(y[3156]), .Z(n11552) );
  ANDN U3904 ( .B(y[3157]), .A(x[3157]), .Z(n11547) );
  ANDN U3905 ( .B(y[3154]), .A(x[3154]), .Z(n18407) );
  NANDN U3906 ( .A(y[3153]), .B(x[3153]), .Z(n11554) );
  ANDN U3907 ( .B(x[3154]), .A(y[3154]), .Z(n18410) );
  ANDN U3908 ( .B(x[3151]), .A(y[3151]), .Z(n18400) );
  NANDN U3909 ( .A(x[3151]), .B(y[3151]), .Z(n20233) );
  ANDN U3910 ( .B(x[3150]), .A(y[3150]), .Z(n18401) );
  ANDN U3911 ( .B(y[3149]), .A(x[3149]), .Z(n18398) );
  NANDN U3912 ( .A(x[3148]), .B(y[3148]), .Z(n2740) );
  NANDN U3913 ( .A(x[3147]), .B(y[3147]), .Z(n2739) );
  NAND U3914 ( .A(n2740), .B(n2739), .Z(n26749) );
  NANDN U3915 ( .A(y[3145]), .B(x[3145]), .Z(n11555) );
  XNOR U3916 ( .A(x[3145]), .B(y[3145]), .Z(n9970) );
  XNOR U3917 ( .A(y[3144]), .B(x[3144]), .Z(n9967) );
  XNOR U3918 ( .A(y[3142]), .B(x[3142]), .Z(n9960) );
  ANDN U3919 ( .B(y[3140]), .A(x[3140]), .Z(n18381) );
  NANDN U3920 ( .A(y[3139]), .B(x[3139]), .Z(n18379) );
  ANDN U3921 ( .B(x[3140]), .A(y[3140]), .Z(n11563) );
  ANDN U3922 ( .B(x[3137]), .A(y[3137]), .Z(n11567) );
  ANDN U3923 ( .B(y[3137]), .A(x[3137]), .Z(n11565) );
  ANDN U3924 ( .B(x[3136]), .A(y[3136]), .Z(n11566) );
  NANDN U3925 ( .A(x[3132]), .B(y[3132]), .Z(n2742) );
  NANDN U3926 ( .A(x[3131]), .B(y[3131]), .Z(n2741) );
  NAND U3927 ( .A(n2742), .B(n2741), .Z(n26716) );
  NANDN U3928 ( .A(x[3130]), .B(y[3130]), .Z(n2744) );
  NANDN U3929 ( .A(x[3129]), .B(y[3129]), .Z(n2743) );
  NAND U3930 ( .A(n2744), .B(n2743), .Z(n26713) );
  ANDN U3931 ( .B(x[3129]), .A(y[3129]), .Z(n11568) );
  XNOR U3932 ( .A(y[3128]), .B(x[3128]), .Z(n9942) );
  ANDN U3933 ( .B(x[3127]), .A(y[3127]), .Z(n11573) );
  NANDN U3934 ( .A(y[3125]), .B(x[3125]), .Z(n11577) );
  ANDN U3935 ( .B(x[3126]), .A(y[3126]), .Z(n11572) );
  ANDN U3936 ( .B(n11577), .A(n11572), .Z(n9937) );
  XNOR U3937 ( .A(x[3125]), .B(y[3125]), .Z(n9935) );
  XNOR U3938 ( .A(y[3124]), .B(x[3124]), .Z(n9932) );
  ANDN U3939 ( .B(x[3123]), .A(y[3123]), .Z(n11581) );
  NANDN U3940 ( .A(y[3121]), .B(x[3121]), .Z(n11583) );
  ANDN U3941 ( .B(x[3122]), .A(y[3122]), .Z(n11580) );
  ANDN U3942 ( .B(n11583), .A(n11580), .Z(n9927) );
  ANDN U3943 ( .B(x[3119]), .A(y[3119]), .Z(n11587) );
  NANDN U3944 ( .A(y[3117]), .B(x[3117]), .Z(n11589) );
  ANDN U3945 ( .B(x[3118]), .A(y[3118]), .Z(n11586) );
  ANDN U3946 ( .B(x[3115]), .A(y[3115]), .Z(n11593) );
  NANDN U3947 ( .A(y[3113]), .B(x[3113]), .Z(n11597) );
  ANDN U3948 ( .B(x[3114]), .A(y[3114]), .Z(n11592) );
  ANDN U3949 ( .B(n11597), .A(n11592), .Z(n9924) );
  ANDN U3950 ( .B(x[3111]), .A(y[3111]), .Z(n11601) );
  NANDN U3951 ( .A(y[3109]), .B(x[3109]), .Z(n11603) );
  ANDN U3952 ( .B(x[3110]), .A(y[3110]), .Z(n11600) );
  ANDN U3953 ( .B(x[3107]), .A(y[3107]), .Z(n11607) );
  NANDN U3954 ( .A(y[3105]), .B(x[3105]), .Z(n11611) );
  ANDN U3955 ( .B(x[3106]), .A(y[3106]), .Z(n11606) );
  ANDN U3956 ( .B(n11611), .A(n11606), .Z(n9922) );
  ANDN U3957 ( .B(x[3103]), .A(y[3103]), .Z(n11615) );
  NANDN U3958 ( .A(y[3101]), .B(x[3101]), .Z(n11616) );
  ANDN U3959 ( .B(x[3102]), .A(y[3102]), .Z(n11614) );
  NANDN U3960 ( .A(y[3099]), .B(x[3099]), .Z(n11621) );
  ANDN U3961 ( .B(x[3100]), .A(y[3100]), .Z(n11617) );
  NANDN U3962 ( .A(x[3096]), .B(y[3096]), .Z(n11624) );
  ANDN U3963 ( .B(y[3097]), .A(x[3097]), .Z(n11622) );
  ANDN U3964 ( .B(n11624), .A(n11622), .Z(n9918) );
  XNOR U3965 ( .A(y[3096]), .B(x[3096]), .Z(n9916) );
  NANDN U3966 ( .A(x[3094]), .B(y[3094]), .Z(n26639) );
  ANDN U3967 ( .B(y[3095]), .A(x[3095]), .Z(n11625) );
  ANDN U3968 ( .B(n26639), .A(n11625), .Z(n9913) );
  ANDN U3969 ( .B(x[3093]), .A(y[3093]), .Z(n11628) );
  XOR U3970 ( .A(x[3094]), .B(y[3094]), .Z(n9910) );
  NANDN U3971 ( .A(x[3091]), .B(y[3091]), .Z(n26634) );
  NANDN U3972 ( .A(y[3089]), .B(x[3089]), .Z(n11631) );
  ANDN U3973 ( .B(x[3090]), .A(y[3090]), .Z(n18315) );
  ANDN U3974 ( .B(n11631), .A(n18315), .Z(n9901) );
  XNOR U3975 ( .A(x[3089]), .B(y[3089]), .Z(n9899) );
  XNOR U3976 ( .A(x[3087]), .B(y[3087]), .Z(n9892) );
  NANDN U3977 ( .A(x[3084]), .B(y[3084]), .Z(n11638) );
  ANDN U3978 ( .B(y[3085]), .A(x[3085]), .Z(n11636) );
  ANDN U3979 ( .B(n11638), .A(n11636), .Z(n9885) );
  XNOR U3980 ( .A(y[3084]), .B(x[3084]), .Z(n9883) );
  XNOR U3981 ( .A(x[3083]), .B(y[3083]), .Z(n9880) );
  ANDN U3982 ( .B(x[3079]), .A(y[3079]), .Z(n18289) );
  NANDN U3983 ( .A(x[3077]), .B(y[3077]), .Z(n18286) );
  NANDN U3984 ( .A(y[3077]), .B(x[3077]), .Z(n2746) );
  NANDN U3985 ( .A(y[3076]), .B(x[3076]), .Z(n2745) );
  AND U3986 ( .A(n2746), .B(n2745), .Z(n26602) );
  NANDN U3987 ( .A(y[3075]), .B(x[3075]), .Z(n11645) );
  NANDN U3988 ( .A(y[3073]), .B(x[3073]), .Z(n18279) );
  ANDN U3989 ( .B(x[3074]), .A(y[3074]), .Z(n11646) );
  IV U3990 ( .A(x[3072]), .Z(n11649) );
  ANDN U3991 ( .B(x[3071]), .A(y[3071]), .Z(n18274) );
  ANDN U3992 ( .B(y[3071]), .A(x[3071]), .Z(n11651) );
  XOR U3993 ( .A(y[3070]), .B(x[3070]), .Z(n11653) );
  NANDN U3994 ( .A(y[3069]), .B(x[3069]), .Z(n26583) );
  ANDN U3995 ( .B(y[3068]), .A(x[3068]), .Z(n11655) );
  ANDN U3996 ( .B(x[3068]), .A(y[3068]), .Z(n11654) );
  NANDN U3997 ( .A(y[3067]), .B(x[3067]), .Z(n26580) );
  NANDN U3998 ( .A(y[3066]), .B(x[3066]), .Z(n26576) );
  NANDN U3999 ( .A(x[3065]), .B(y[3065]), .Z(n26575) );
  NANDN U4000 ( .A(x[3064]), .B(y[3064]), .Z(n11660) );
  AND U4001 ( .A(n26575), .B(n11660), .Z(n9867) );
  XNOR U4002 ( .A(y[3064]), .B(x[3064]), .Z(n9865) );
  NANDN U4003 ( .A(y[3063]), .B(x[3063]), .Z(n26568) );
  NANDN U4004 ( .A(x[3062]), .B(y[3062]), .Z(n26566) );
  NANDN U4005 ( .A(y[3061]), .B(x[3061]), .Z(n18256) );
  NANDN U4006 ( .A(y[3062]), .B(x[3062]), .Z(n18261) );
  NAND U4007 ( .A(n18256), .B(n18261), .Z(n26565) );
  NANDN U4008 ( .A(x[3060]), .B(y[3060]), .Z(n2747) );
  ANDN U4009 ( .B(y[3061]), .A(x[3061]), .Z(n11662) );
  ANDN U4010 ( .B(n2747), .A(n11662), .Z(n26562) );
  ANDN U4011 ( .B(y[3058]), .A(x[3058]), .Z(n11664) );
  NANDN U4012 ( .A(x[3059]), .B(y[3059]), .Z(n26558) );
  NANDN U4013 ( .A(y[3058]), .B(x[3058]), .Z(n26557) );
  NANDN U4014 ( .A(y[3057]), .B(x[3057]), .Z(n18244) );
  AND U4015 ( .A(n26557), .B(n18244), .Z(n9855) );
  XNOR U4016 ( .A(x[3057]), .B(y[3057]), .Z(n9853) );
  NANDN U4017 ( .A(x[3056]), .B(y[3056]), .Z(n26550) );
  NANDN U4018 ( .A(y[3055]), .B(x[3055]), .Z(n26549) );
  NANDN U4019 ( .A(y[3053]), .B(x[3053]), .Z(n26543) );
  NANDN U4020 ( .A(x[3051]), .B(y[3051]), .Z(n26536) );
  NANDN U4021 ( .A(x[3048]), .B(y[3048]), .Z(n26528) );
  ANDN U4022 ( .B(y[3049]), .A(x[3049]), .Z(n11667) );
  NANDN U4023 ( .A(y[3047]), .B(x[3047]), .Z(n11671) );
  NANDN U4024 ( .A(y[3048]), .B(x[3048]), .Z(n18225) );
  NAND U4025 ( .A(n11671), .B(n18225), .Z(n26527) );
  NANDN U4026 ( .A(y[3044]), .B(x[3044]), .Z(n26518) );
  NANDN U4027 ( .A(y[3041]), .B(x[3041]), .Z(n26510) );
  ANDN U4028 ( .B(x[3042]), .A(y[3042]), .Z(n18209) );
  IV U4029 ( .A(x[3040]), .Z(n18202) );
  NAND U4030 ( .A(n18202), .B(y[3040]), .Z(n2748) );
  NANDN U4031 ( .A(x[3041]), .B(y[3041]), .Z(n11672) );
  NAND U4032 ( .A(n2748), .B(n11672), .Z(n26509) );
  NANDN U4033 ( .A(x[3038]), .B(y[3038]), .Z(n18193) );
  NANDN U4034 ( .A(x[3039]), .B(y[3039]), .Z(n2749) );
  NAND U4035 ( .A(n18193), .B(n2749), .Z(n26505) );
  NANDN U4036 ( .A(x[3037]), .B(y[3037]), .Z(n26500) );
  NANDN U4037 ( .A(x[3034]), .B(y[3034]), .Z(n26492) );
  ANDN U4038 ( .B(y[3035]), .A(x[3035]), .Z(n11673) );
  NANDN U4039 ( .A(y[3033]), .B(x[3033]), .Z(n11677) );
  NANDN U4040 ( .A(y[3034]), .B(x[3034]), .Z(n18185) );
  NAND U4041 ( .A(n11677), .B(n18185), .Z(n26491) );
  NANDN U4042 ( .A(y[3030]), .B(x[3030]), .Z(n26482) );
  NANDN U4043 ( .A(y[3027]), .B(x[3027]), .Z(n26474) );
  ANDN U4044 ( .B(x[3028]), .A(y[3028]), .Z(n18169) );
  NANDN U4045 ( .A(x[3023]), .B(y[3023]), .Z(n26464) );
  NANDN U4046 ( .A(x[3020]), .B(y[3020]), .Z(n26456) );
  ANDN U4047 ( .B(y[3021]), .A(x[3021]), .Z(n11682) );
  ANDN U4048 ( .B(n26456), .A(n11682), .Z(n9844) );
  NANDN U4049 ( .A(y[3016]), .B(x[3016]), .Z(n26446) );
  NANDN U4050 ( .A(y[3013]), .B(x[3013]), .Z(n26438) );
  ANDN U4051 ( .B(x[3014]), .A(y[3014]), .Z(n11688) );
  NANDN U4052 ( .A(x[3012]), .B(y[3012]), .Z(n18128) );
  NANDN U4053 ( .A(x[3013]), .B(y[3013]), .Z(n18134) );
  NAND U4054 ( .A(n18128), .B(n18134), .Z(n26437) );
  NANDN U4055 ( .A(x[3009]), .B(y[3009]), .Z(n26428) );
  NANDN U4056 ( .A(x[3006]), .B(y[3006]), .Z(n26420) );
  ANDN U4057 ( .B(y[3007]), .A(x[3007]), .Z(n11691) );
  NANDN U4058 ( .A(y[3005]), .B(x[3005]), .Z(n11695) );
  NANDN U4059 ( .A(y[3006]), .B(x[3006]), .Z(n18114) );
  NAND U4060 ( .A(n11695), .B(n18114), .Z(n26419) );
  NANDN U4061 ( .A(y[3002]), .B(x[3002]), .Z(n26410) );
  NANDN U4062 ( .A(y[2999]), .B(x[2999]), .Z(n26402) );
  ANDN U4063 ( .B(x[3000]), .A(y[3000]), .Z(n11698) );
  NANDN U4064 ( .A(x[2998]), .B(y[2998]), .Z(n18093) );
  NANDN U4065 ( .A(x[2999]), .B(y[2999]), .Z(n18099) );
  NAND U4066 ( .A(n18093), .B(n18099), .Z(n26401) );
  NANDN U4067 ( .A(x[2995]), .B(y[2995]), .Z(n26392) );
  NANDN U4068 ( .A(x[2992]), .B(y[2992]), .Z(n26384) );
  ANDN U4069 ( .B(y[2993]), .A(x[2993]), .Z(n11701) );
  NANDN U4070 ( .A(y[2991]), .B(x[2991]), .Z(n11704) );
  NANDN U4071 ( .A(y[2992]), .B(x[2992]), .Z(n18079) );
  NAND U4072 ( .A(n11704), .B(n18079), .Z(n26383) );
  NANDN U4073 ( .A(y[2988]), .B(x[2988]), .Z(n26374) );
  NANDN U4074 ( .A(y[2985]), .B(x[2985]), .Z(n26366) );
  ANDN U4075 ( .B(x[2986]), .A(y[2986]), .Z(n11706) );
  NANDN U4076 ( .A(x[2984]), .B(y[2984]), .Z(n18058) );
  NANDN U4077 ( .A(x[2985]), .B(y[2985]), .Z(n18064) );
  NAND U4078 ( .A(n18058), .B(n18064), .Z(n26365) );
  NANDN U4079 ( .A(x[2981]), .B(y[2981]), .Z(n26356) );
  NANDN U4080 ( .A(x[2978]), .B(y[2978]), .Z(n26348) );
  ANDN U4081 ( .B(y[2979]), .A(x[2979]), .Z(n11709) );
  NANDN U4082 ( .A(y[2977]), .B(x[2977]), .Z(n11713) );
  NANDN U4083 ( .A(y[2978]), .B(x[2978]), .Z(n18044) );
  NAND U4084 ( .A(n11713), .B(n18044), .Z(n26347) );
  NANDN U4085 ( .A(y[2974]), .B(x[2974]), .Z(n26338) );
  NANDN U4086 ( .A(y[2971]), .B(x[2971]), .Z(n26330) );
  ANDN U4087 ( .B(x[2972]), .A(y[2972]), .Z(n11715) );
  ANDN U4088 ( .B(n26330), .A(n11715), .Z(n9835) );
  NANDN U4089 ( .A(x[2970]), .B(y[2970]), .Z(n18023) );
  NANDN U4090 ( .A(x[2971]), .B(y[2971]), .Z(n18029) );
  NAND U4091 ( .A(n18023), .B(n18029), .Z(n26329) );
  NANDN U4092 ( .A(x[2967]), .B(y[2967]), .Z(n26320) );
  NANDN U4093 ( .A(x[2964]), .B(y[2964]), .Z(n26312) );
  ANDN U4094 ( .B(y[2965]), .A(x[2965]), .Z(n11718) );
  NANDN U4095 ( .A(y[2963]), .B(x[2963]), .Z(n11722) );
  NANDN U4096 ( .A(y[2964]), .B(x[2964]), .Z(n18009) );
  NAND U4097 ( .A(n11722), .B(n18009), .Z(n26310) );
  NANDN U4098 ( .A(x[2962]), .B(y[2962]), .Z(n18002) );
  ANDN U4099 ( .B(y[2963]), .A(x[2963]), .Z(n11720) );
  ANDN U4100 ( .B(n18002), .A(n11720), .Z(n26308) );
  ANDN U4101 ( .B(y[2960]), .A(x[2960]), .Z(n11725) );
  NANDN U4102 ( .A(x[2961]), .B(y[2961]), .Z(n26304) );
  NANDN U4103 ( .A(x[2958]), .B(y[2958]), .Z(n26296) );
  ANDN U4104 ( .B(y[2959]), .A(x[2959]), .Z(n11724) );
  ANDN U4105 ( .B(n26296), .A(n11724), .Z(n9833) );
  ANDN U4106 ( .B(x[2958]), .A(y[2958]), .Z(n11727) );
  NANDN U4107 ( .A(x[2956]), .B(y[2956]), .Z(n17990) );
  NANDN U4108 ( .A(x[2957]), .B(y[2957]), .Z(n17996) );
  NAND U4109 ( .A(n17990), .B(n17996), .Z(n26293) );
  XNOR U4110 ( .A(y[2952]), .B(x[2952]), .Z(n9822) );
  ANDN U4111 ( .B(y[2951]), .A(x[2951]), .Z(n17980) );
  NANDN U4112 ( .A(x[2950]), .B(y[2950]), .Z(n26277) );
  ANDN U4113 ( .B(y[2946]), .A(x[2946]), .Z(n11732) );
  NANDN U4114 ( .A(y[2946]), .B(x[2946]), .Z(n26270) );
  NANDN U4115 ( .A(y[2945]), .B(x[2945]), .Z(n11734) );
  AND U4116 ( .A(n26270), .B(n11734), .Z(n9807) );
  XNOR U4117 ( .A(x[2945]), .B(y[2945]), .Z(n9805) );
  NANDN U4118 ( .A(x[2944]), .B(y[2944]), .Z(n26264) );
  NANDN U4119 ( .A(y[2937]), .B(x[2937]), .Z(n26247) );
  ANDN U4120 ( .B(x[2938]), .A(y[2938]), .Z(n17953) );
  ANDN U4121 ( .B(y[2937]), .A(x[2937]), .Z(n17949) );
  NANDN U4122 ( .A(y[2935]), .B(x[2935]), .Z(n2750) );
  NANDN U4123 ( .A(y[2936]), .B(x[2936]), .Z(n11738) );
  NAND U4124 ( .A(n2750), .B(n11738), .Z(n26243) );
  NANDN U4125 ( .A(x[2934]), .B(y[2934]), .Z(n17936) );
  IV U4126 ( .A(x[2935]), .Z(n17943) );
  NAND U4127 ( .A(n17943), .B(y[2935]), .Z(n2751) );
  NAND U4128 ( .A(n17936), .B(n2751), .Z(n26240) );
  XNOR U4129 ( .A(x[2934]), .B(y[2934]), .Z(n2752) );
  ANDN U4130 ( .B(x[2933]), .A(y[2933]), .Z(n11739) );
  ANDN U4131 ( .B(n2752), .A(n11739), .Z(n26238) );
  ANDN U4132 ( .B(y[2932]), .A(x[2932]), .Z(n11741) );
  NANDN U4133 ( .A(y[2932]), .B(x[2932]), .Z(n26234) );
  NANDN U4134 ( .A(x[2930]), .B(y[2930]), .Z(n26228) );
  ANDN U4135 ( .B(y[2931]), .A(x[2931]), .Z(n11740) );
  ANDN U4136 ( .B(n26228), .A(n11740), .Z(n9796) );
  ANDN U4137 ( .B(y[2927]), .A(x[2927]), .Z(n11744) );
  NANDN U4138 ( .A(x[2926]), .B(y[2926]), .Z(n17917) );
  NANDN U4139 ( .A(n11744), .B(n17917), .Z(n26220) );
  ANDN U4140 ( .B(x[2925]), .A(y[2925]), .Z(n11747) );
  NANDN U4141 ( .A(y[2926]), .B(x[2926]), .Z(n26218) );
  NANDN U4142 ( .A(x[2925]), .B(y[2925]), .Z(n26217) );
  NANDN U4143 ( .A(x[2924]), .B(y[2924]), .Z(n17913) );
  AND U4144 ( .A(n26217), .B(n17913), .Z(n9788) );
  XNOR U4145 ( .A(y[2924]), .B(x[2924]), .Z(n9786) );
  NANDN U4146 ( .A(y[2923]), .B(x[2923]), .Z(n26210) );
  NANDN U4147 ( .A(x[2922]), .B(y[2922]), .Z(n26209) );
  NANDN U4148 ( .A(y[2919]), .B(x[2919]), .Z(n17898) );
  NANDN U4149 ( .A(y[2920]), .B(x[2920]), .Z(n2753) );
  NAND U4150 ( .A(n17898), .B(n2753), .Z(n26203) );
  ANDN U4151 ( .B(y[2918]), .A(x[2918]), .Z(n11750) );
  NANDN U4152 ( .A(y[2918]), .B(x[2918]), .Z(n26198) );
  NANDN U4153 ( .A(y[2917]), .B(x[2917]), .Z(n11752) );
  NANDN U4154 ( .A(x[2916]), .B(y[2916]), .Z(n26193) );
  ANDN U4155 ( .B(y[2911]), .A(x[2911]), .Z(n26178) );
  NANDN U4156 ( .A(y[2911]), .B(x[2911]), .Z(n2755) );
  NANDN U4157 ( .A(y[2910]), .B(x[2910]), .Z(n2754) );
  AND U4158 ( .A(n2755), .B(n2754), .Z(n26176) );
  ANDN U4159 ( .B(y[2904]), .A(x[2904]), .Z(n11759) );
  NANDN U4160 ( .A(y[2904]), .B(x[2904]), .Z(n26164) );
  NANDN U4161 ( .A(y[2903]), .B(x[2903]), .Z(n11761) );
  AND U4162 ( .A(n26164), .B(n11761), .Z(n9762) );
  XNOR U4163 ( .A(x[2903]), .B(y[2903]), .Z(n9760) );
  NANDN U4164 ( .A(x[2902]), .B(y[2902]), .Z(n26158) );
  NANDN U4165 ( .A(y[2901]), .B(x[2901]), .Z(n26156) );
  IV U4166 ( .A(y[2899]), .Z(n17861) );
  NANDN U4167 ( .A(x[2898]), .B(y[2898]), .Z(n17858) );
  NANDN U4168 ( .A(x[2899]), .B(y[2899]), .Z(n2756) );
  NAND U4169 ( .A(n17858), .B(n2756), .Z(n26150) );
  ANDN U4170 ( .B(x[2897]), .A(y[2897]), .Z(n11764) );
  NANDN U4171 ( .A(y[2898]), .B(x[2898]), .Z(n26148) );
  NANDN U4172 ( .A(x[2897]), .B(y[2897]), .Z(n26147) );
  NANDN U4173 ( .A(x[2896]), .B(y[2896]), .Z(n17853) );
  AND U4174 ( .A(n26147), .B(n17853), .Z(n9749) );
  XNOR U4175 ( .A(y[2896]), .B(x[2896]), .Z(n9747) );
  NANDN U4176 ( .A(y[2895]), .B(x[2895]), .Z(n26140) );
  NANDN U4177 ( .A(x[2894]), .B(y[2894]), .Z(n26139) );
  ANDN U4178 ( .B(y[2890]), .A(x[2890]), .Z(n11771) );
  NANDN U4179 ( .A(x[2891]), .B(y[2891]), .Z(n26131) );
  NANDN U4180 ( .A(y[2890]), .B(x[2890]), .Z(n26128) );
  NANDN U4181 ( .A(y[2889]), .B(x[2889]), .Z(n17839) );
  AND U4182 ( .A(n26128), .B(n17839), .Z(n9737) );
  XNOR U4183 ( .A(x[2889]), .B(y[2889]), .Z(n9735) );
  NANDN U4184 ( .A(x[2888]), .B(y[2888]), .Z(n26122) );
  NANDN U4185 ( .A(y[2887]), .B(x[2887]), .Z(n26120) );
  ANDN U4186 ( .B(x[2886]), .A(y[2886]), .Z(n17831) );
  NANDN U4187 ( .A(y[2885]), .B(x[2885]), .Z(n2757) );
  NANDN U4188 ( .A(n17831), .B(n2757), .Z(n9726) );
  NANDN U4189 ( .A(y[2884]), .B(x[2884]), .Z(n2758) );
  NANDN U4190 ( .A(n9726), .B(n2758), .Z(n26116) );
  NANDN U4191 ( .A(y[2881]), .B(x[2881]), .Z(n26108) );
  ANDN U4192 ( .B(x[2882]), .A(y[2882]), .Z(n11774) );
  ANDN U4193 ( .B(n26108), .A(n11774), .Z(n9720) );
  ANDN U4194 ( .B(y[2880]), .A(x[2880]), .Z(n26107) );
  ANDN U4195 ( .B(y[2881]), .A(x[2881]), .Z(n11776) );
  NANDN U4196 ( .A(y[2877]), .B(x[2877]), .Z(n17813) );
  NANDN U4197 ( .A(y[2878]), .B(x[2878]), .Z(n11778) );
  AND U4198 ( .A(n17813), .B(n11778), .Z(n26100) );
  NANDN U4199 ( .A(y[2876]), .B(x[2876]), .Z(n26096) );
  NANDN U4200 ( .A(x[2870]), .B(y[2870]), .Z(n11785) );
  NANDN U4201 ( .A(x[2871]), .B(y[2871]), .Z(n2759) );
  NAND U4202 ( .A(n11785), .B(n2759), .Z(n26082) );
  IV U4203 ( .A(x[2869]), .Z(n20234) );
  OR U4204 ( .A(y[2869]), .B(n20234), .Z(n17792) );
  ANDN U4205 ( .B(x[2870]), .A(y[2870]), .Z(n26080) );
  ANDN U4206 ( .B(n17792), .A(n26080), .Z(n9697) );
  ANDN U4207 ( .B(y[2869]), .A(x[2869]), .Z(n11784) );
  NANDN U4208 ( .A(y[2865]), .B(x[2865]), .Z(n17781) );
  NANDN U4209 ( .A(y[2866]), .B(x[2866]), .Z(n11787) );
  NAND U4210 ( .A(n17781), .B(n11787), .Z(n26071) );
  NANDN U4211 ( .A(x[2863]), .B(y[2863]), .Z(n26064) );
  ANDN U4212 ( .B(x[2862]), .A(y[2862]), .Z(n17776) );
  ANDN U4213 ( .B(y[2861]), .A(x[2861]), .Z(n17773) );
  NANDN U4214 ( .A(x[2858]), .B(y[2858]), .Z(n26052) );
  NANDN U4215 ( .A(y[2851]), .B(x[2851]), .Z(n11797) );
  NANDN U4216 ( .A(y[2852]), .B(x[2852]), .Z(n17760) );
  NAND U4217 ( .A(n11797), .B(n17760), .Z(n26033) );
  NANDN U4218 ( .A(x[2850]), .B(y[2850]), .Z(n17752) );
  NANDN U4219 ( .A(x[2851]), .B(y[2851]), .Z(n17757) );
  NAND U4220 ( .A(n17752), .B(n17757), .Z(n26031) );
  NANDN U4221 ( .A(y[2849]), .B(x[2849]), .Z(n17749) );
  NANDN U4222 ( .A(y[2850]), .B(x[2850]), .Z(n11796) );
  NAND U4223 ( .A(n17749), .B(n11796), .Z(n26028) );
  ANDN U4224 ( .B(y[2848]), .A(x[2848]), .Z(n11799) );
  ANDN U4225 ( .B(y[2847]), .A(x[2847]), .Z(n11798) );
  NANDN U4226 ( .A(x[2846]), .B(y[2846]), .Z(n26019) );
  NANDN U4227 ( .A(x[2841]), .B(y[2841]), .Z(n26007) );
  ANDN U4228 ( .B(y[2839]), .A(x[2839]), .Z(n17734) );
  NANDN U4229 ( .A(x[2838]), .B(y[2838]), .Z(n25999) );
  NANDN U4230 ( .A(x[2836]), .B(y[2836]), .Z(n11801) );
  NANDN U4231 ( .A(x[2837]), .B(y[2837]), .Z(n2760) );
  NAND U4232 ( .A(n11801), .B(n2760), .Z(n25994) );
  ANDN U4233 ( .B(x[2833]), .A(y[2833]), .Z(n11803) );
  NANDN U4234 ( .A(y[2834]), .B(x[2834]), .Z(n25988) );
  ANDN U4235 ( .B(y[2831]), .A(x[2831]), .Z(n17711) );
  NANDN U4236 ( .A(y[2830]), .B(x[2830]), .Z(n25973) );
  ANDN U4237 ( .B(x[2831]), .A(y[2831]), .Z(n25983) );
  NANDN U4238 ( .A(y[2829]), .B(x[2829]), .Z(n25974) );
  IV U4239 ( .A(y[2828]), .Z(n11804) );
  NAND U4240 ( .A(n11804), .B(x[2828]), .Z(n25966) );
  AND U4241 ( .A(n25974), .B(n25966), .Z(n9651) );
  XNOR U4242 ( .A(x[2828]), .B(y[2828]), .Z(n9649) );
  NANDN U4243 ( .A(x[2827]), .B(y[2827]), .Z(n25964) );
  NANDN U4244 ( .A(y[2825]), .B(x[2825]), .Z(n25958) );
  ANDN U4245 ( .B(y[2824]), .A(x[2824]), .Z(n25956) );
  NANDN U4246 ( .A(y[2822]), .B(x[2822]), .Z(n25950) );
  ANDN U4247 ( .B(y[2820]), .A(x[2820]), .Z(n11808) );
  ANDN U4248 ( .B(x[2820]), .A(y[2820]), .Z(n17688) );
  NANDN U4249 ( .A(x[2818]), .B(y[2818]), .Z(n25938) );
  ANDN U4250 ( .B(y[2819]), .A(x[2819]), .Z(n11807) );
  ANDN U4251 ( .B(n25938), .A(n11807), .Z(n9630) );
  ANDN U4252 ( .B(x[2818]), .A(y[2818]), .Z(n17684) );
  ANDN U4253 ( .B(x[2813]), .A(y[2813]), .Z(n9613) );
  NANDN U4254 ( .A(x[2812]), .B(y[2812]), .Z(n11809) );
  OR U4255 ( .A(n9613), .B(n11809), .Z(n9620) );
  NANDN U4256 ( .A(y[2809]), .B(x[2809]), .Z(n11818) );
  ANDN U4257 ( .B(x[2810]), .A(y[2810]), .Z(n11815) );
  ANDN U4258 ( .B(n11818), .A(n11815), .Z(n25917) );
  ANDN U4259 ( .B(y[2806]), .A(x[2806]), .Z(n11822) );
  NANDN U4260 ( .A(x[2807]), .B(y[2807]), .Z(n25911) );
  NANDN U4261 ( .A(y[2805]), .B(x[2805]), .Z(n11823) );
  ANDN U4262 ( .B(x[2806]), .A(y[2806]), .Z(n25909) );
  ANDN U4263 ( .B(n11823), .A(n25909), .Z(n9602) );
  XNOR U4264 ( .A(x[2805]), .B(y[2805]), .Z(n9600) );
  NANDN U4265 ( .A(x[2804]), .B(y[2804]), .Z(n25903) );
  NANDN U4266 ( .A(y[2803]), .B(x[2803]), .Z(n25901) );
  NANDN U4267 ( .A(x[2802]), .B(y[2802]), .Z(n17654) );
  NANDN U4268 ( .A(x[2803]), .B(y[2803]), .Z(n17660) );
  NAND U4269 ( .A(n17654), .B(n17660), .Z(n25900) );
  ANDN U4270 ( .B(x[2802]), .A(y[2802]), .Z(n11825) );
  ANDN U4271 ( .B(x[2801]), .A(y[2801]), .Z(n17650) );
  NOR U4272 ( .A(n11825), .B(n17650), .Z(n25897) );
  ANDN U4273 ( .B(x[2799]), .A(y[2799]), .Z(n11827) );
  NANDN U4274 ( .A(y[2800]), .B(x[2800]), .Z(n25893) );
  NANDN U4275 ( .A(x[2799]), .B(y[2799]), .Z(n25892) );
  NANDN U4276 ( .A(x[2798]), .B(y[2798]), .Z(n17643) );
  AND U4277 ( .A(n25892), .B(n17643), .Z(n9590) );
  XNOR U4278 ( .A(y[2798]), .B(x[2798]), .Z(n9588) );
  NANDN U4279 ( .A(y[2797]), .B(x[2797]), .Z(n25885) );
  NANDN U4280 ( .A(x[2796]), .B(y[2796]), .Z(n25884) );
  NANDN U4281 ( .A(y[2795]), .B(x[2795]), .Z(n17636) );
  NANDN U4282 ( .A(y[2796]), .B(x[2796]), .Z(n17640) );
  NAND U4283 ( .A(n17636), .B(n17640), .Z(n25881) );
  NANDN U4284 ( .A(x[2793]), .B(y[2793]), .Z(n25876) );
  NANDN U4285 ( .A(x[2790]), .B(y[2790]), .Z(n2762) );
  NANDN U4286 ( .A(x[2789]), .B(y[2789]), .Z(n2761) );
  NAND U4287 ( .A(n2762), .B(n2761), .Z(n25868) );
  NANDN U4288 ( .A(y[2780]), .B(x[2780]), .Z(n2764) );
  NANDN U4289 ( .A(y[2779]), .B(x[2779]), .Z(n2763) );
  AND U4290 ( .A(n2764), .B(n2763), .Z(n25842) );
  NANDN U4291 ( .A(x[2768]), .B(y[2768]), .Z(n11833) );
  NANDN U4292 ( .A(x[2769]), .B(y[2769]), .Z(n17597) );
  NAND U4293 ( .A(n11833), .B(n17597), .Z(n25819) );
  NANDN U4294 ( .A(y[2768]), .B(x[2768]), .Z(n11831) );
  IV U4295 ( .A(x[2766]), .Z(n11835) );
  NAND U4296 ( .A(n11835), .B(y[2766]), .Z(n17590) );
  IV U4297 ( .A(x[2767]), .Z(n11834) );
  NAND U4298 ( .A(n11834), .B(y[2767]), .Z(n11832) );
  NAND U4299 ( .A(n17590), .B(n11832), .Z(n25815) );
  ANDN U4300 ( .B(y[2764]), .A(x[2764]), .Z(n11838) );
  ANDN U4301 ( .B(y[2763]), .A(x[2763]), .Z(n11837) );
  NANDN U4302 ( .A(x[2762]), .B(y[2762]), .Z(n25803) );
  NANDN U4303 ( .A(x[2758]), .B(y[2758]), .Z(n11844) );
  NANDN U4304 ( .A(x[2759]), .B(y[2759]), .Z(n11841) );
  NAND U4305 ( .A(n11844), .B(n11841), .Z(n25795) );
  ANDN U4306 ( .B(x[2757]), .A(y[2757]), .Z(n11846) );
  NANDN U4307 ( .A(y[2758]), .B(x[2758]), .Z(n25792) );
  NANDN U4308 ( .A(x[2757]), .B(y[2757]), .Z(n25791) );
  NANDN U4309 ( .A(x[2756]), .B(y[2756]), .Z(n11847) );
  AND U4310 ( .A(n25791), .B(n11847), .Z(n9500) );
  XNOR U4311 ( .A(y[2756]), .B(x[2756]), .Z(n9498) );
  NANDN U4312 ( .A(y[2755]), .B(x[2755]), .Z(n25784) );
  NANDN U4313 ( .A(y[2754]), .B(x[2754]), .Z(n17565) );
  ANDN U4314 ( .B(x[2753]), .A(y[2753]), .Z(n11849) );
  ANDN U4315 ( .B(n17565), .A(n11849), .Z(n25780) );
  ANDN U4316 ( .B(y[2752]), .A(x[2752]), .Z(n11851) );
  NANDN U4317 ( .A(x[2753]), .B(y[2753]), .Z(n25778) );
  ANDN U4318 ( .B(x[2751]), .A(y[2751]), .Z(n11853) );
  ANDN U4319 ( .B(y[2751]), .A(x[2751]), .Z(n11850) );
  NANDN U4320 ( .A(y[2749]), .B(x[2749]), .Z(n17554) );
  ANDN U4321 ( .B(x[2750]), .A(y[2750]), .Z(n11852) );
  ANDN U4322 ( .B(n17554), .A(n11852), .Z(n9486) );
  XNOR U4323 ( .A(x[2749]), .B(y[2749]), .Z(n9484) );
  NANDN U4324 ( .A(x[2748]), .B(y[2748]), .Z(n25766) );
  NANDN U4325 ( .A(x[2746]), .B(y[2746]), .Z(n11858) );
  NANDN U4326 ( .A(x[2747]), .B(y[2747]), .Z(n17551) );
  AND U4327 ( .A(n11858), .B(n17551), .Z(n25762) );
  NANDN U4328 ( .A(y[2744]), .B(x[2744]), .Z(n25757) );
  NANDN U4329 ( .A(y[2743]), .B(x[2743]), .Z(n2766) );
  NANDN U4330 ( .A(y[2742]), .B(x[2742]), .Z(n2765) );
  NAND U4331 ( .A(n2766), .B(n2765), .Z(n25753) );
  NANDN U4332 ( .A(y[2741]), .B(x[2741]), .Z(n25748) );
  NANDN U4333 ( .A(y[2739]), .B(x[2739]), .Z(n2768) );
  XNOR U4334 ( .A(x[2740]), .B(y[2740]), .Z(n2767) );
  NAND U4335 ( .A(n2768), .B(n2767), .Z(n25744) );
  NANDN U4336 ( .A(x[2738]), .B(y[2738]), .Z(n17527) );
  IV U4337 ( .A(x[2739]), .Z(n17533) );
  NAND U4338 ( .A(n17533), .B(y[2739]), .Z(n2769) );
  NAND U4339 ( .A(n17527), .B(n2769), .Z(n25743) );
  NANDN U4340 ( .A(x[2734]), .B(y[2734]), .Z(n25730) );
  NANDN U4341 ( .A(y[2733]), .B(x[2733]), .Z(n25729) );
  NANDN U4342 ( .A(x[2732]), .B(y[2732]), .Z(n11868) );
  NANDN U4343 ( .A(x[2733]), .B(y[2733]), .Z(n17519) );
  NAND U4344 ( .A(n11868), .B(n17519), .Z(n25726) );
  ANDN U4345 ( .B(x[2729]), .A(y[2729]), .Z(n11871) );
  NANDN U4346 ( .A(y[2730]), .B(x[2730]), .Z(n25721) );
  NANDN U4347 ( .A(x[2729]), .B(y[2729]), .Z(n25718) );
  NANDN U4348 ( .A(x[2728]), .B(y[2728]), .Z(n17507) );
  AND U4349 ( .A(n25718), .B(n17507), .Z(n9448) );
  XNOR U4350 ( .A(y[2728]), .B(x[2728]), .Z(n9446) );
  NANDN U4351 ( .A(x[2726]), .B(y[2726]), .Z(n25710) );
  IV U4352 ( .A(x[2724]), .Z(n17495) );
  NAND U4353 ( .A(n17495), .B(y[2724]), .Z(n2770) );
  ANDN U4354 ( .B(y[2725]), .A(x[2725]), .Z(n11873) );
  ANDN U4355 ( .B(n2770), .A(n11873), .Z(n25706) );
  NANDN U4356 ( .A(y[2723]), .B(x[2723]), .Z(n17490) );
  NANDN U4357 ( .A(y[2724]), .B(x[2724]), .Z(n2771) );
  NAND U4358 ( .A(n17490), .B(n2771), .Z(n25705) );
  ANDN U4359 ( .B(x[2722]), .A(y[2722]), .Z(n17493) );
  NANDN U4360 ( .A(y[2721]), .B(x[2721]), .Z(n17486) );
  NANDN U4361 ( .A(n17493), .B(n17486), .Z(n2772) );
  ANDN U4362 ( .B(y[2722]), .A(x[2722]), .Z(n9434) );
  ANDN U4363 ( .B(n2772), .A(n9434), .Z(n25701) );
  ANDN U4364 ( .B(y[2717]), .A(x[2717]), .Z(n11874) );
  ANDN U4365 ( .B(y[2716]), .A(x[2716]), .Z(n17467) );
  NOR U4366 ( .A(n11874), .B(n17467), .Z(n25690) );
  ANDN U4367 ( .B(x[2715]), .A(y[2715]), .Z(n17464) );
  ANDN U4368 ( .B(x[2714]), .A(y[2714]), .Z(n17463) );
  NANDN U4369 ( .A(x[2712]), .B(y[2712]), .Z(n2774) );
  NANDN U4370 ( .A(x[2713]), .B(y[2713]), .Z(n2773) );
  NAND U4371 ( .A(n2774), .B(n2773), .Z(n11878) );
  XOR U4372 ( .A(x[2712]), .B(y[2712]), .Z(n11877) );
  NANDN U4373 ( .A(y[2711]), .B(x[2711]), .Z(n2775) );
  NANDN U4374 ( .A(n11877), .B(n2775), .Z(n9419) );
  ANDN U4375 ( .B(y[2711]), .A(x[2711]), .Z(n11876) );
  NANDN U4376 ( .A(x[2710]), .B(y[2710]), .Z(n11880) );
  NANDN U4377 ( .A(n11876), .B(n11880), .Z(n2776) );
  NANDN U4378 ( .A(n9419), .B(n2776), .Z(n2777) );
  NANDN U4379 ( .A(n11878), .B(n2777), .Z(n25683) );
  ANDN U4380 ( .B(x[2709]), .A(y[2709]), .Z(n11881) );
  NANDN U4381 ( .A(x[2708]), .B(y[2708]), .Z(n25674) );
  NANDN U4382 ( .A(x[2709]), .B(y[2709]), .Z(n25678) );
  AND U4383 ( .A(n25674), .B(n25678), .Z(n9417) );
  ANDN U4384 ( .B(x[2708]), .A(y[2708]), .Z(n11882) );
  NANDN U4385 ( .A(x[2702]), .B(y[2702]), .Z(n2779) );
  NANDN U4386 ( .A(x[2703]), .B(y[2703]), .Z(n2778) );
  NAND U4387 ( .A(n2779), .B(n2778), .Z(n25658) );
  XNOR U4388 ( .A(x[2702]), .B(y[2702]), .Z(n25656) );
  NANDN U4389 ( .A(x[2698]), .B(y[2698]), .Z(n25647) );
  NANDN U4390 ( .A(y[2697]), .B(x[2697]), .Z(n11885) );
  NANDN U4391 ( .A(y[2698]), .B(x[2698]), .Z(n17439) );
  NAND U4392 ( .A(n11885), .B(n17439), .Z(n25645) );
  ANDN U4393 ( .B(y[2694]), .A(x[2694]), .Z(n17426) );
  NANDN U4394 ( .A(x[2695]), .B(y[2695]), .Z(n25637) );
  NANDN U4395 ( .A(y[2691]), .B(x[2691]), .Z(n2781) );
  NANDN U4396 ( .A(y[2692]), .B(x[2692]), .Z(n2780) );
  AND U4397 ( .A(n2781), .B(n2780), .Z(n25628) );
  NANDN U4398 ( .A(y[2688]), .B(x[2688]), .Z(n25616) );
  IV U4399 ( .A(y[2687]), .Z(n25618) );
  NAND U4400 ( .A(n25618), .B(x[2687]), .Z(n2782) );
  AND U4401 ( .A(n25616), .B(n2782), .Z(n17417) );
  NANDN U4402 ( .A(x[2687]), .B(y[2687]), .Z(n2784) );
  NANDN U4403 ( .A(x[2686]), .B(y[2686]), .Z(n2783) );
  NAND U4404 ( .A(n2784), .B(n2783), .Z(n17415) );
  NANDN U4405 ( .A(x[2682]), .B(y[2682]), .Z(n2786) );
  NANDN U4406 ( .A(x[2683]), .B(y[2683]), .Z(n2785) );
  NAND U4407 ( .A(n2786), .B(n2785), .Z(n25603) );
  NANDN U4408 ( .A(y[2680]), .B(x[2680]), .Z(n25597) );
  NANDN U4409 ( .A(y[2679]), .B(x[2679]), .Z(n11888) );
  AND U4410 ( .A(n25597), .B(n11888), .Z(n9359) );
  XNOR U4411 ( .A(x[2679]), .B(y[2679]), .Z(n9357) );
  NANDN U4412 ( .A(x[2678]), .B(y[2678]), .Z(n25591) );
  NANDN U4413 ( .A(y[2677]), .B(x[2677]), .Z(n25589) );
  NANDN U4414 ( .A(y[2676]), .B(x[2676]), .Z(n11890) );
  NANDN U4415 ( .A(y[2675]), .B(x[2675]), .Z(n2787) );
  NAND U4416 ( .A(n11890), .B(n2787), .Z(n9348) );
  NANDN U4417 ( .A(y[2674]), .B(x[2674]), .Z(n2788) );
  NANDN U4418 ( .A(n9348), .B(n2788), .Z(n25585) );
  NANDN U4419 ( .A(y[2671]), .B(x[2671]), .Z(n25577) );
  ANDN U4420 ( .B(x[2672]), .A(y[2672]), .Z(n11893) );
  ANDN U4421 ( .B(n25577), .A(n11893), .Z(n9342) );
  ANDN U4422 ( .B(y[2671]), .A(x[2671]), .Z(n17388) );
  ANDN U4423 ( .B(y[2670]), .A(x[2670]), .Z(n25576) );
  ANDN U4424 ( .B(x[2668]), .A(y[2668]), .Z(n11895) );
  ANDN U4425 ( .B(x[2667]), .A(y[2667]), .Z(n17375) );
  NOR U4426 ( .A(n11895), .B(n17375), .Z(n25569) );
  ANDN U4427 ( .B(y[2666]), .A(x[2666]), .Z(n11898) );
  ANDN U4428 ( .B(x[2665]), .A(y[2665]), .Z(n11900) );
  NANDN U4429 ( .A(y[2666]), .B(x[2666]), .Z(n25565) );
  ANDN U4430 ( .B(x[2664]), .A(y[2664]), .Z(n11899) );
  NANDN U4431 ( .A(y[2663]), .B(x[2663]), .Z(n25557) );
  NANDN U4432 ( .A(y[2662]), .B(x[2662]), .Z(n17368) );
  ANDN U4433 ( .B(x[2661]), .A(y[2661]), .Z(n11903) );
  ANDN U4434 ( .B(n17368), .A(n11903), .Z(n25553) );
  NANDN U4435 ( .A(x[2659]), .B(y[2659]), .Z(n25548) );
  IV U4436 ( .A(y[2655]), .Z(n17351) );
  NAND U4437 ( .A(n17351), .B(x[2655]), .Z(n2789) );
  ANDN U4438 ( .B(x[2656]), .A(y[2656]), .Z(n11910) );
  ANDN U4439 ( .B(n2789), .A(n11910), .Z(n25537) );
  NANDN U4440 ( .A(x[2654]), .B(y[2654]), .Z(n17348) );
  NANDN U4441 ( .A(x[2655]), .B(y[2655]), .Z(n2790) );
  NAND U4442 ( .A(n17348), .B(n2790), .Z(n25536) );
  NANDN U4443 ( .A(x[2653]), .B(y[2653]), .Z(n25531) );
  NANDN U4444 ( .A(y[2652]), .B(x[2652]), .Z(n11911) );
  XNOR U4445 ( .A(x[2652]), .B(y[2652]), .Z(n9326) );
  NANDN U4446 ( .A(y[2645]), .B(x[2645]), .Z(n11915) );
  XNOR U4447 ( .A(x[2645]), .B(y[2645]), .Z(n9306) );
  ANDN U4448 ( .B(y[2643]), .A(x[2643]), .Z(n11918) );
  NANDN U4449 ( .A(x[2642]), .B(y[2642]), .Z(n25507) );
  NANDN U4450 ( .A(y[2641]), .B(x[2641]), .Z(n11921) );
  NANDN U4451 ( .A(y[2642]), .B(x[2642]), .Z(n17332) );
  NAND U4452 ( .A(n11921), .B(n17332), .Z(n25505) );
  NANDN U4453 ( .A(y[2638]), .B(x[2638]), .Z(n20241) );
  ANDN U4454 ( .B(x[2637]), .A(y[2637]), .Z(n11922) );
  ANDN U4455 ( .B(n20241), .A(n11922), .Z(n25495) );
  NANDN U4456 ( .A(x[2636]), .B(y[2636]), .Z(n25493) );
  NANDN U4457 ( .A(x[2637]), .B(y[2637]), .Z(n17319) );
  NAND U4458 ( .A(n25493), .B(n17319), .Z(n9293) );
  NANDN U4459 ( .A(y[2634]), .B(x[2634]), .Z(n2792) );
  NANDN U4460 ( .A(y[2633]), .B(x[2633]), .Z(n2791) );
  AND U4461 ( .A(n2792), .B(n2791), .Z(n25487) );
  NANDN U4462 ( .A(x[2632]), .B(y[2632]), .Z(n2794) );
  NANDN U4463 ( .A(x[2633]), .B(y[2633]), .Z(n2793) );
  NAND U4464 ( .A(n2794), .B(n2793), .Z(n25486) );
  XNOR U4465 ( .A(x[2632]), .B(y[2632]), .Z(n25483) );
  ANDN U4466 ( .B(y[2631]), .A(x[2631]), .Z(n11929) );
  ANDN U4467 ( .B(y[2629]), .A(x[2629]), .Z(n11925) );
  NANDN U4468 ( .A(x[2628]), .B(y[2628]), .Z(n25478) );
  NANDN U4469 ( .A(y[2625]), .B(x[2625]), .Z(n17295) );
  NANDN U4470 ( .A(y[2626]), .B(x[2626]), .Z(n17301) );
  NAND U4471 ( .A(n17295), .B(n17301), .Z(n25472) );
  NANDN U4472 ( .A(x[2624]), .B(y[2624]), .Z(n17292) );
  NANDN U4473 ( .A(x[2625]), .B(y[2625]), .Z(n11931) );
  NAND U4474 ( .A(n17292), .B(n11931), .Z(n25469) );
  ANDN U4475 ( .B(x[2623]), .A(y[2623]), .Z(n11934) );
  NANDN U4476 ( .A(y[2624]), .B(x[2624]), .Z(n25467) );
  NANDN U4477 ( .A(x[2622]), .B(y[2622]), .Z(n25462) );
  NANDN U4478 ( .A(x[2623]), .B(y[2623]), .Z(n25466) );
  AND U4479 ( .A(n25462), .B(n25466), .Z(n9269) );
  ANDN U4480 ( .B(x[2622]), .A(y[2622]), .Z(n11933) );
  ANDN U4481 ( .B(x[2618]), .A(y[2618]), .Z(n25447) );
  NANDN U4482 ( .A(x[2617]), .B(y[2617]), .Z(n25445) );
  NANDN U4483 ( .A(x[2614]), .B(y[2614]), .Z(n25438) );
  NANDN U4484 ( .A(y[2613]), .B(x[2613]), .Z(n2795) );
  NANDN U4485 ( .A(y[2614]), .B(x[2614]), .Z(n17276) );
  NAND U4486 ( .A(n2795), .B(n17276), .Z(n25435) );
  NANDN U4487 ( .A(x[2612]), .B(y[2612]), .Z(n2797) );
  NANDN U4488 ( .A(x[2613]), .B(y[2613]), .Z(n2796) );
  NAND U4489 ( .A(n2797), .B(n2796), .Z(n25433) );
  NANDN U4490 ( .A(x[2609]), .B(y[2609]), .Z(n2799) );
  NANDN U4491 ( .A(x[2610]), .B(y[2610]), .Z(n2798) );
  NAND U4492 ( .A(n2799), .B(n2798), .Z(n25425) );
  NANDN U4493 ( .A(x[2608]), .B(y[2608]), .Z(n2801) );
  NANDN U4494 ( .A(x[2607]), .B(y[2607]), .Z(n2800) );
  NAND U4495 ( .A(n2801), .B(n2800), .Z(n25421) );
  ANDN U4496 ( .B(x[2603]), .A(y[2603]), .Z(n2802) );
  ANDN U4497 ( .B(y[2602]), .A(x[2602]), .Z(n11938) );
  NANDN U4498 ( .A(y[2602]), .B(x[2602]), .Z(n2803) );
  ANDN U4499 ( .B(n2803), .A(n2802), .Z(n25411) );
  ANDN U4500 ( .B(x[2601]), .A(y[2601]), .Z(n11940) );
  NANDN U4501 ( .A(x[2600]), .B(y[2600]), .Z(n11943) );
  ANDN U4502 ( .B(y[2601]), .A(x[2601]), .Z(n11939) );
  ANDN U4503 ( .B(y[2597]), .A(x[2597]), .Z(n17247) );
  NANDN U4504 ( .A(x[2596]), .B(y[2596]), .Z(n25397) );
  NANDN U4505 ( .A(x[2595]), .B(y[2595]), .Z(n17234) );
  IV U4506 ( .A(x[2594]), .Z(n17235) );
  NAND U4507 ( .A(n17235), .B(y[2594]), .Z(n2804) );
  NAND U4508 ( .A(n17234), .B(n2804), .Z(n25394) );
  IV U4509 ( .A(y[2593]), .Z(n17228) );
  NAND U4510 ( .A(n17228), .B(x[2593]), .Z(n2806) );
  NANDN U4511 ( .A(y[2594]), .B(x[2594]), .Z(n2805) );
  AND U4512 ( .A(n2806), .B(n2805), .Z(n25391) );
  NANDN U4513 ( .A(x[2592]), .B(y[2592]), .Z(n11947) );
  NANDN U4514 ( .A(x[2593]), .B(y[2593]), .Z(n2807) );
  NAND U4515 ( .A(n11947), .B(n2807), .Z(n25389) );
  NANDN U4516 ( .A(x[2588]), .B(y[2588]), .Z(n17211) );
  NANDN U4517 ( .A(x[2589]), .B(y[2589]), .Z(n17218) );
  AND U4518 ( .A(n17211), .B(n17218), .Z(n25381) );
  NANDN U4519 ( .A(y[2585]), .B(x[2585]), .Z(n25375) );
  ANDN U4520 ( .B(x[2586]), .A(y[2586]), .Z(n11949) );
  NANDN U4521 ( .A(x[2585]), .B(y[2585]), .Z(n11953) );
  NANDN U4522 ( .A(y[2583]), .B(x[2583]), .Z(n17201) );
  NANDN U4523 ( .A(y[2584]), .B(x[2584]), .Z(n2808) );
  NAND U4524 ( .A(n17201), .B(n2808), .Z(n25372) );
  NANDN U4525 ( .A(x[2581]), .B(y[2581]), .Z(n25365) );
  ANDN U4526 ( .B(y[2580]), .A(x[2580]), .Z(n11955) );
  ANDN U4527 ( .B(n25365), .A(n11955), .Z(n9224) );
  ANDN U4528 ( .B(x[2580]), .A(y[2580]), .Z(n25363) );
  NANDN U4529 ( .A(x[2578]), .B(y[2578]), .Z(n25357) );
  NANDN U4530 ( .A(y[2575]), .B(x[2575]), .Z(n17179) );
  NANDN U4531 ( .A(y[2576]), .B(x[2576]), .Z(n2809) );
  NAND U4532 ( .A(n17179), .B(n2809), .Z(n25350) );
  NANDN U4533 ( .A(y[2574]), .B(x[2574]), .Z(n2811) );
  NANDN U4534 ( .A(y[2573]), .B(x[2573]), .Z(n2810) );
  AND U4535 ( .A(n2811), .B(n2810), .Z(n25344) );
  ANDN U4536 ( .B(y[2574]), .A(x[2574]), .Z(n25345) );
  NOR U4537 ( .A(n25344), .B(n25345), .Z(n17178) );
  NANDN U4538 ( .A(x[2567]), .B(y[2567]), .Z(n2813) );
  NANDN U4539 ( .A(x[2566]), .B(y[2566]), .Z(n2812) );
  NAND U4540 ( .A(n2813), .B(n2812), .Z(n25329) );
  NANDN U4541 ( .A(y[2566]), .B(x[2566]), .Z(n2815) );
  NANDN U4542 ( .A(y[2565]), .B(x[2565]), .Z(n2814) );
  AND U4543 ( .A(n2815), .B(n2814), .Z(n25327) );
  NANDN U4544 ( .A(y[2564]), .B(x[2564]), .Z(n2817) );
  NANDN U4545 ( .A(y[2563]), .B(x[2563]), .Z(n2816) );
  AND U4546 ( .A(n2817), .B(n2816), .Z(n25323) );
  NANDN U4547 ( .A(y[2562]), .B(x[2562]), .Z(n2819) );
  NANDN U4548 ( .A(y[2561]), .B(x[2561]), .Z(n2818) );
  AND U4549 ( .A(n2819), .B(n2818), .Z(n25319) );
  ANDN U4550 ( .B(y[2560]), .A(x[2560]), .Z(n11957) );
  ANDN U4551 ( .B(x[2558]), .A(y[2558]), .Z(n17158) );
  NANDN U4552 ( .A(y[2557]), .B(x[2557]), .Z(n25307) );
  NANDN U4553 ( .A(x[2556]), .B(y[2556]), .Z(n11960) );
  NANDN U4554 ( .A(x[2557]), .B(y[2557]), .Z(n17156) );
  NAND U4555 ( .A(n11960), .B(n17156), .Z(n25306) );
  NANDN U4556 ( .A(y[2555]), .B(x[2555]), .Z(n2820) );
  ANDN U4557 ( .B(x[2556]), .A(y[2556]), .Z(n11958) );
  ANDN U4558 ( .B(n2820), .A(n11958), .Z(n25303) );
  NANDN U4559 ( .A(x[2554]), .B(y[2554]), .Z(n17146) );
  NANDN U4560 ( .A(x[2555]), .B(y[2555]), .Z(n11959) );
  NAND U4561 ( .A(n17146), .B(n11959), .Z(n25301) );
  NANDN U4562 ( .A(x[2553]), .B(y[2553]), .Z(n25298) );
  ANDN U4563 ( .B(y[2551]), .A(x[2551]), .Z(n11965) );
  NANDN U4564 ( .A(x[2550]), .B(y[2550]), .Z(n25290) );
  ANDN U4565 ( .B(y[2548]), .A(x[2548]), .Z(n11967) );
  NANDN U4566 ( .A(x[2549]), .B(y[2549]), .Z(n17139) );
  NANDN U4567 ( .A(n11967), .B(n17139), .Z(n25285) );
  NANDN U4568 ( .A(x[2547]), .B(y[2547]), .Z(n25282) );
  NANDN U4569 ( .A(x[2546]), .B(y[2546]), .Z(n9163) );
  NANDN U4570 ( .A(x[2545]), .B(y[2545]), .Z(n2821) );
  NAND U4571 ( .A(n9163), .B(n2821), .Z(n17129) );
  NANDN U4572 ( .A(x[2544]), .B(y[2544]), .Z(n2822) );
  NANDN U4573 ( .A(n17129), .B(n2822), .Z(n25278) );
  ANDN U4574 ( .B(x[2544]), .A(y[2544]), .Z(n17127) );
  NANDN U4575 ( .A(x[2542]), .B(y[2542]), .Z(n2824) );
  NANDN U4576 ( .A(x[2543]), .B(y[2543]), .Z(n2823) );
  NAND U4577 ( .A(n2824), .B(n2823), .Z(n25274) );
  NANDN U4578 ( .A(x[2539]), .B(y[2539]), .Z(n2826) );
  NANDN U4579 ( .A(x[2538]), .B(y[2538]), .Z(n2825) );
  NAND U4580 ( .A(n2826), .B(n2825), .Z(n25265) );
  ANDN U4581 ( .B(y[2535]), .A(x[2535]), .Z(n17114) );
  NANDN U4582 ( .A(x[2534]), .B(y[2534]), .Z(n17108) );
  NANDN U4583 ( .A(x[2533]), .B(y[2533]), .Z(n25254) );
  NANDN U4584 ( .A(x[2531]), .B(y[2531]), .Z(n2828) );
  NANDN U4585 ( .A(x[2532]), .B(y[2532]), .Z(n2827) );
  NAND U4586 ( .A(n2828), .B(n2827), .Z(n25249) );
  ANDN U4587 ( .B(x[2531]), .A(y[2531]), .Z(n11970) );
  ANDN U4588 ( .B(x[2530]), .A(y[2530]), .Z(n11969) );
  NANDN U4589 ( .A(y[2529]), .B(x[2529]), .Z(n25243) );
  ANDN U4590 ( .B(x[2526]), .A(y[2526]), .Z(n11974) );
  ANDN U4591 ( .B(x[2525]), .A(y[2525]), .Z(n17088) );
  NOR U4592 ( .A(n11974), .B(n17088), .Z(n25235) );
  NANDN U4593 ( .A(y[2524]), .B(x[2524]), .Z(n25231) );
  NANDN U4594 ( .A(x[2523]), .B(y[2523]), .Z(n2830) );
  NANDN U4595 ( .A(x[2524]), .B(y[2524]), .Z(n2829) );
  NAND U4596 ( .A(n2830), .B(n2829), .Z(n25230) );
  XNOR U4597 ( .A(x[2523]), .B(y[2523]), .Z(n25227) );
  NANDN U4598 ( .A(y[2521]), .B(x[2521]), .Z(n2832) );
  NANDN U4599 ( .A(y[2522]), .B(x[2522]), .Z(n2831) );
  AND U4600 ( .A(n2832), .B(n2831), .Z(n25223) );
  NANDN U4601 ( .A(y[2518]), .B(x[2518]), .Z(n25215) );
  NANDN U4602 ( .A(y[2517]), .B(x[2517]), .Z(n25214) );
  NANDN U4603 ( .A(y[2516]), .B(x[2516]), .Z(n20245) );
  AND U4604 ( .A(n25214), .B(n20245), .Z(n17071) );
  NANDN U4605 ( .A(x[2517]), .B(y[2517]), .Z(n17074) );
  NANDN U4606 ( .A(x[2512]), .B(y[2512]), .Z(n2834) );
  NANDN U4607 ( .A(x[2511]), .B(y[2511]), .Z(n2833) );
  NAND U4608 ( .A(n2834), .B(n2833), .Z(n17060) );
  NANDN U4609 ( .A(x[2510]), .B(y[2510]), .Z(n11981) );
  NANDN U4610 ( .A(y[2511]), .B(x[2511]), .Z(n9127) );
  NANDN U4611 ( .A(n11981), .B(n9127), .Z(n2835) );
  NANDN U4612 ( .A(n17060), .B(n2835), .Z(n25200) );
  NANDN U4613 ( .A(x[2508]), .B(y[2508]), .Z(n11984) );
  NANDN U4614 ( .A(x[2509]), .B(y[2509]), .Z(n11980) );
  NAND U4615 ( .A(n11984), .B(n11980), .Z(n25196) );
  ANDN U4616 ( .B(y[2504]), .A(x[2504]), .Z(n11989) );
  NANDN U4617 ( .A(x[2505]), .B(y[2505]), .Z(n25188) );
  NANDN U4618 ( .A(y[2504]), .B(x[2504]), .Z(n25185) );
  NANDN U4619 ( .A(y[2503]), .B(x[2503]), .Z(n17040) );
  AND U4620 ( .A(n25185), .B(n17040), .Z(n9122) );
  XNOR U4621 ( .A(x[2503]), .B(y[2503]), .Z(n9120) );
  IV U4622 ( .A(x[2502]), .Z(n11990) );
  NANDN U4623 ( .A(x[2499]), .B(y[2499]), .Z(n17035) );
  NAND U4624 ( .A(n17028), .B(n17035), .Z(n25172) );
  ANDN U4625 ( .B(y[2495]), .A(x[2495]), .Z(n9100) );
  NANDN U4626 ( .A(x[2494]), .B(y[2494]), .Z(n2836) );
  NANDN U4627 ( .A(n9100), .B(n2836), .Z(n25164) );
  NANDN U4628 ( .A(x[2490]), .B(y[2490]), .Z(n2838) );
  NANDN U4629 ( .A(x[2489]), .B(y[2489]), .Z(n2837) );
  AND U4630 ( .A(n2838), .B(n2837), .Z(n25153) );
  ANDN U4631 ( .B(x[2489]), .A(y[2489]), .Z(n11995) );
  NANDN U4632 ( .A(y[2487]), .B(x[2487]), .Z(n25148) );
  ANDN U4633 ( .B(x[2488]), .A(y[2488]), .Z(n11994) );
  ANDN U4634 ( .B(n25148), .A(n11994), .Z(n9083) );
  NANDN U4635 ( .A(y[2485]), .B(x[2485]), .Z(n2839) );
  ANDN U4636 ( .B(x[2486]), .A(y[2486]), .Z(n11997) );
  ANDN U4637 ( .B(n2839), .A(n11997), .Z(n25143) );
  NANDN U4638 ( .A(y[2482]), .B(x[2482]), .Z(n25136) );
  NANDN U4639 ( .A(x[2480]), .B(y[2480]), .Z(n25129) );
  ANDN U4640 ( .B(y[2481]), .A(x[2481]), .Z(n11999) );
  ANDN U4641 ( .B(n25129), .A(n11999), .Z(n9069) );
  NANDN U4642 ( .A(x[2476]), .B(y[2476]), .Z(n16987) );
  ANDN U4643 ( .B(y[2477]), .A(x[2477]), .Z(n12004) );
  ANDN U4644 ( .B(n16987), .A(n12004), .Z(n25121) );
  ANDN U4645 ( .B(x[2475]), .A(y[2475]), .Z(n12006) );
  NANDN U4646 ( .A(x[2469]), .B(y[2469]), .Z(n2841) );
  NANDN U4647 ( .A(x[2468]), .B(y[2468]), .Z(n2840) );
  AND U4648 ( .A(n2841), .B(n2840), .Z(n25101) );
  NANDN U4649 ( .A(x[2464]), .B(y[2464]), .Z(n16968) );
  ANDN U4650 ( .B(y[2465]), .A(x[2465]), .Z(n16973) );
  ANDN U4651 ( .B(n16968), .A(n16973), .Z(n25093) );
  NANDN U4652 ( .A(x[2461]), .B(y[2461]), .Z(n2842) );
  ANDN U4653 ( .B(y[2462]), .A(x[2462]), .Z(n9030) );
  ANDN U4654 ( .B(n2842), .A(n9030), .Z(n25085) );
  IV U4655 ( .A(y[2460]), .Z(n16960) );
  ANDN U4656 ( .B(x[2459]), .A(y[2459]), .Z(n25080) );
  ANDN U4657 ( .B(y[2459]), .A(x[2459]), .Z(n12009) );
  NANDN U4658 ( .A(x[2455]), .B(y[2455]), .Z(n25069) );
  ANDN U4659 ( .B(y[2454]), .A(x[2454]), .Z(n16943) );
  ANDN U4660 ( .B(n25069), .A(n16943), .Z(n9017) );
  ANDN U4661 ( .B(x[2454]), .A(y[2454]), .Z(n25067) );
  NANDN U4662 ( .A(x[2452]), .B(y[2452]), .Z(n25061) );
  NANDN U4663 ( .A(y[2451]), .B(x[2451]), .Z(n12015) );
  NANDN U4664 ( .A(y[2452]), .B(x[2452]), .Z(n16941) );
  NAND U4665 ( .A(n12015), .B(n16941), .Z(n25060) );
  NANDN U4666 ( .A(y[2449]), .B(x[2449]), .Z(n2843) );
  IV U4667 ( .A(y[2450]), .Z(n12016) );
  NAND U4668 ( .A(n12016), .B(x[2450]), .Z(n12014) );
  NAND U4669 ( .A(n2843), .B(n12014), .Z(n25055) );
  NANDN U4670 ( .A(x[2448]), .B(y[2448]), .Z(n16926) );
  NANDN U4671 ( .A(x[2449]), .B(y[2449]), .Z(n2844) );
  AND U4672 ( .A(n16926), .B(n2844), .Z(n25053) );
  ANDN U4673 ( .B(x[2447]), .A(y[2447]), .Z(n12020) );
  ANDN U4674 ( .B(x[2448]), .A(y[2448]), .Z(n25052) );
  ANDN U4675 ( .B(x[2446]), .A(y[2446]), .Z(n12017) );
  NANDN U4676 ( .A(y[2445]), .B(x[2445]), .Z(n25045) );
  NANDN U4677 ( .A(y[2443]), .B(x[2443]), .Z(n16916) );
  NANDN U4678 ( .A(y[2444]), .B(x[2444]), .Z(n2845) );
  AND U4679 ( .A(n16916), .B(n2845), .Z(n25041) );
  NANDN U4680 ( .A(x[2442]), .B(y[2442]), .Z(n2847) );
  NANDN U4681 ( .A(x[2443]), .B(y[2443]), .Z(n2846) );
  NAND U4682 ( .A(n2847), .B(n2846), .Z(n25040) );
  ANDN U4683 ( .B(y[2439]), .A(x[2439]), .Z(n12023) );
  NANDN U4684 ( .A(x[2438]), .B(y[2438]), .Z(n2848) );
  ANDN U4685 ( .B(y[2437]), .A(x[2437]), .Z(n25025) );
  ANDN U4686 ( .B(n2848), .A(n25025), .Z(n16905) );
  NANDN U4687 ( .A(x[2432]), .B(y[2432]), .Z(n25011) );
  ANDN U4688 ( .B(y[2433]), .A(x[2433]), .Z(n16899) );
  ANDN U4689 ( .B(n25011), .A(n16899), .Z(n8979) );
  NANDN U4690 ( .A(y[2431]), .B(x[2431]), .Z(n25009) );
  NANDN U4691 ( .A(y[2432]), .B(x[2432]), .Z(n25013) );
  NAND U4692 ( .A(n25009), .B(n25013), .Z(n16893) );
  NANDN U4693 ( .A(y[2427]), .B(x[2427]), .Z(n24997) );
  ANDN U4694 ( .B(x[2428]), .A(y[2428]), .Z(n16884) );
  IV U4695 ( .A(n16884), .Z(n25001) );
  AND U4696 ( .A(n24997), .B(n25001), .Z(n8970) );
  NANDN U4697 ( .A(x[2427]), .B(y[2427]), .Z(n24999) );
  NANDN U4698 ( .A(x[2426]), .B(y[2426]), .Z(n24993) );
  NAND U4699 ( .A(n24999), .B(n24993), .Z(n16879) );
  ANDN U4700 ( .B(x[2426]), .A(y[2426]), .Z(n24995) );
  ANDN U4701 ( .B(x[2425]), .A(y[2425]), .Z(n24992) );
  NOR U4702 ( .A(n24995), .B(n24992), .Z(n16877) );
  NANDN U4703 ( .A(y[2424]), .B(x[2424]), .Z(n2850) );
  NANDN U4704 ( .A(y[2423]), .B(x[2423]), .Z(n2849) );
  NAND U4705 ( .A(n2850), .B(n2849), .Z(n24987) );
  ANDN U4706 ( .B(y[2421]), .A(x[2421]), .Z(n12026) );
  NANDN U4707 ( .A(x[2420]), .B(y[2420]), .Z(n2851) );
  NANDN U4708 ( .A(n12026), .B(n2851), .Z(n12030) );
  ANDN U4709 ( .B(x[2420]), .A(y[2420]), .Z(n12025) );
  NANDN U4710 ( .A(y[2417]), .B(x[2417]), .Z(n24976) );
  ANDN U4711 ( .B(x[2418]), .A(y[2418]), .Z(n16870) );
  ANDN U4712 ( .B(n24976), .A(n16870), .Z(n8949) );
  NANDN U4713 ( .A(y[2415]), .B(x[2415]), .Z(n2852) );
  ANDN U4714 ( .B(x[2416]), .A(y[2416]), .Z(n16862) );
  ANDN U4715 ( .B(n2852), .A(n16862), .Z(n24971) );
  ANDN U4716 ( .B(x[2414]), .A(y[2414]), .Z(n12031) );
  ANDN U4717 ( .B(x[2413]), .A(y[2413]), .Z(n12033) );
  NOR U4718 ( .A(n12031), .B(n12033), .Z(n24967) );
  ANDN U4719 ( .B(y[2411]), .A(x[2411]), .Z(n16852) );
  NANDN U4720 ( .A(y[2409]), .B(x[2409]), .Z(n24955) );
  NANDN U4721 ( .A(y[2407]), .B(x[2407]), .Z(n2854) );
  NANDN U4722 ( .A(y[2408]), .B(x[2408]), .Z(n2853) );
  NAND U4723 ( .A(n2854), .B(n2853), .Z(n24950) );
  NANDN U4724 ( .A(y[2406]), .B(x[2406]), .Z(n24946) );
  ANDN U4725 ( .B(x[2405]), .A(y[2405]), .Z(n16841) );
  NANDN U4726 ( .A(x[2404]), .B(y[2404]), .Z(n24939) );
  ANDN U4727 ( .B(x[2403]), .A(y[2403]), .Z(n24937) );
  NANDN U4728 ( .A(x[2399]), .B(y[2399]), .Z(n24927) );
  ANDN U4729 ( .B(y[2398]), .A(x[2398]), .Z(n16822) );
  ANDN U4730 ( .B(n24927), .A(n16822), .Z(n8916) );
  ANDN U4731 ( .B(x[2398]), .A(y[2398]), .Z(n24925) );
  NANDN U4732 ( .A(x[2392]), .B(y[2392]), .Z(n12039) );
  XNOR U4733 ( .A(y[2392]), .B(x[2392]), .Z(n8901) );
  XNOR U4734 ( .A(x[2391]), .B(y[2391]), .Z(n8898) );
  IV U4735 ( .A(y[2387]), .Z(n16798) );
  NAND U4736 ( .A(n16798), .B(x[2387]), .Z(n2856) );
  NANDN U4737 ( .A(y[2388]), .B(x[2388]), .Z(n2855) );
  NAND U4738 ( .A(n2856), .B(n2855), .Z(n24898) );
  IV U4739 ( .A(x[2384]), .Z(n16785) );
  NAND U4740 ( .A(n16785), .B(y[2384]), .Z(n2858) );
  NANDN U4741 ( .A(x[2385]), .B(y[2385]), .Z(n2857) );
  NAND U4742 ( .A(n2858), .B(n2857), .Z(n24891) );
  NANDN U4743 ( .A(y[2384]), .B(x[2384]), .Z(n2859) );
  ANDN U4744 ( .B(x[2383]), .A(y[2383]), .Z(n16779) );
  ANDN U4745 ( .B(n2859), .A(n16779), .Z(n24889) );
  NANDN U4746 ( .A(y[2379]), .B(x[2379]), .Z(n2861) );
  IV U4747 ( .A(y[2380]), .Z(n16770) );
  NAND U4748 ( .A(n16770), .B(x[2380]), .Z(n2860) );
  NAND U4749 ( .A(n2861), .B(n2860), .Z(n24881) );
  NANDN U4750 ( .A(x[2378]), .B(y[2378]), .Z(n16761) );
  NANDN U4751 ( .A(x[2379]), .B(y[2379]), .Z(n2862) );
  AND U4752 ( .A(n16761), .B(n2862), .Z(n24879) );
  ANDN U4753 ( .B(x[2378]), .A(y[2378]), .Z(n24875) );
  NANDN U4754 ( .A(y[2375]), .B(x[2375]), .Z(n24872) );
  ANDN U4755 ( .B(x[2376]), .A(y[2376]), .Z(n12044) );
  ANDN U4756 ( .B(n24872), .A(n12044), .Z(n8872) );
  NANDN U4757 ( .A(x[2371]), .B(y[2371]), .Z(n24861) );
  ANDN U4758 ( .B(y[2370]), .A(x[2370]), .Z(n12051) );
  ANDN U4759 ( .B(n24861), .A(n12051), .Z(n8864) );
  ANDN U4760 ( .B(x[2370]), .A(y[2370]), .Z(n24859) );
  NANDN U4761 ( .A(x[2368]), .B(y[2368]), .Z(n24853) );
  ANDN U4762 ( .B(x[2367]), .A(y[2367]), .Z(n24852) );
  IV U4763 ( .A(x[2365]), .Z(n12055) );
  NAND U4764 ( .A(n12055), .B(y[2365]), .Z(n12053) );
  NANDN U4765 ( .A(x[2363]), .B(y[2363]), .Z(n2863) );
  NANDN U4766 ( .A(x[2364]), .B(y[2364]), .Z(n12056) );
  AND U4767 ( .A(n2863), .B(n12056), .Z(n16728) );
  NANDN U4768 ( .A(y[2364]), .B(x[2364]), .Z(n8853) );
  NANDN U4769 ( .A(x[2362]), .B(y[2362]), .Z(n24840) );
  NANDN U4770 ( .A(x[2357]), .B(y[2357]), .Z(n2865) );
  NANDN U4771 ( .A(x[2356]), .B(y[2356]), .Z(n2864) );
  AND U4772 ( .A(n2865), .B(n2864), .Z(n24827) );
  NANDN U4773 ( .A(x[2355]), .B(y[2355]), .Z(n2867) );
  NANDN U4774 ( .A(x[2354]), .B(y[2354]), .Z(n2866) );
  NAND U4775 ( .A(n2867), .B(n2866), .Z(n12061) );
  NANDN U4776 ( .A(y[2354]), .B(x[2354]), .Z(n12060) );
  NANDN U4777 ( .A(y[2353]), .B(x[2353]), .Z(n2868) );
  NAND U4778 ( .A(n12060), .B(n2868), .Z(n2872) );
  ANDN U4779 ( .B(y[2352]), .A(x[2352]), .Z(n16706) );
  ANDN U4780 ( .B(y[2353]), .A(x[2353]), .Z(n12059) );
  OR U4781 ( .A(n16706), .B(n12059), .Z(n2869) );
  NANDN U4782 ( .A(n2872), .B(n2869), .Z(n2870) );
  NANDN U4783 ( .A(n12061), .B(n2870), .Z(n24824) );
  NANDN U4784 ( .A(y[2352]), .B(x[2352]), .Z(n2871) );
  NANDN U4785 ( .A(n2872), .B(n2871), .Z(n24822) );
  NANDN U4786 ( .A(x[2351]), .B(y[2351]), .Z(n24819) );
  ANDN U4787 ( .B(y[2350]), .A(x[2350]), .Z(n8837) );
  NANDN U4788 ( .A(y[2349]), .B(x[2349]), .Z(n16699) );
  ANDN U4789 ( .B(y[2347]), .A(x[2347]), .Z(n16696) );
  ANDN U4790 ( .B(y[2346]), .A(x[2346]), .Z(n12063) );
  NOR U4791 ( .A(n16696), .B(n12063), .Z(n24811) );
  NANDN U4792 ( .A(y[2345]), .B(x[2345]), .Z(n16688) );
  NANDN U4793 ( .A(y[2346]), .B(x[2346]), .Z(n16694) );
  NAND U4794 ( .A(n16688), .B(n16694), .Z(n24810) );
  ANDN U4795 ( .B(x[2343]), .A(y[2343]), .Z(n12067) );
  NANDN U4796 ( .A(y[2344]), .B(x[2344]), .Z(n24806) );
  NANDN U4797 ( .A(x[2343]), .B(y[2343]), .Z(n24803) );
  NANDN U4798 ( .A(x[2342]), .B(y[2342]), .Z(n16683) );
  XNOR U4799 ( .A(y[2342]), .B(x[2342]), .Z(n8834) );
  NANDN U4800 ( .A(y[2341]), .B(x[2341]), .Z(n24798) );
  NANDN U4801 ( .A(x[2337]), .B(y[2337]), .Z(n24787) );
  NANDN U4802 ( .A(y[2336]), .B(x[2336]), .Z(n2874) );
  NANDN U4803 ( .A(y[2337]), .B(x[2337]), .Z(n2873) );
  NAND U4804 ( .A(n2874), .B(n2873), .Z(n12074) );
  NANDN U4805 ( .A(y[2335]), .B(x[2335]), .Z(n12069) );
  NANDN U4806 ( .A(x[2336]), .B(y[2336]), .Z(n2875) );
  NANDN U4807 ( .A(n12069), .B(n2875), .Z(n8824) );
  NANDN U4808 ( .A(x[2334]), .B(y[2334]), .Z(n2877) );
  NANDN U4809 ( .A(x[2335]), .B(y[2335]), .Z(n2876) );
  NAND U4810 ( .A(n2876), .B(n2875), .Z(n12072) );
  ANDN U4811 ( .B(n2877), .A(n12072), .Z(n24783) );
  ANDN U4812 ( .B(x[2334]), .A(y[2334]), .Z(n12070) );
  NANDN U4813 ( .A(y[2333]), .B(x[2333]), .Z(n24782) );
  NANDN U4814 ( .A(y[2332]), .B(x[2332]), .Z(n2879) );
  NANDN U4815 ( .A(y[2331]), .B(x[2331]), .Z(n2878) );
  NAND U4816 ( .A(n2879), .B(n2878), .Z(n24777) );
  NANDN U4817 ( .A(y[2329]), .B(x[2329]), .Z(n2881) );
  NANDN U4818 ( .A(y[2330]), .B(x[2330]), .Z(n2880) );
  AND U4819 ( .A(n2881), .B(n2880), .Z(n24773) );
  NANDN U4820 ( .A(x[2328]), .B(y[2328]), .Z(n2882) );
  NANDN U4821 ( .A(x[2329]), .B(y[2329]), .Z(n24772) );
  NAND U4822 ( .A(n2882), .B(n24772), .Z(n16662) );
  NANDN U4823 ( .A(y[2327]), .B(x[2327]), .Z(n24764) );
  IV U4824 ( .A(y[2328]), .Z(n24767) );
  NAND U4825 ( .A(n24767), .B(x[2328]), .Z(n2883) );
  NAND U4826 ( .A(n24764), .B(n2883), .Z(n16661) );
  ANDN U4827 ( .B(y[2325]), .A(x[2325]), .Z(n12076) );
  NANDN U4828 ( .A(x[2324]), .B(y[2324]), .Z(n2884) );
  NANDN U4829 ( .A(n12076), .B(n2884), .Z(n8802) );
  NANDN U4830 ( .A(x[2323]), .B(y[2323]), .Z(n2885) );
  NANDN U4831 ( .A(n8802), .B(n2885), .Z(n24758) );
  ANDN U4832 ( .B(x[2321]), .A(y[2321]), .Z(n16650) );
  ANDN U4833 ( .B(x[2320]), .A(y[2320]), .Z(n16649) );
  NANDN U4834 ( .A(x[2318]), .B(y[2318]), .Z(n12081) );
  NANDN U4835 ( .A(x[2319]), .B(y[2319]), .Z(n16646) );
  NAND U4836 ( .A(n12081), .B(n16646), .Z(n24747) );
  NANDN U4837 ( .A(y[2317]), .B(x[2317]), .Z(n2886) );
  ANDN U4838 ( .B(x[2318]), .A(y[2318]), .Z(n12079) );
  ANDN U4839 ( .B(n2886), .A(n12079), .Z(n24744) );
  NANDN U4840 ( .A(x[2317]), .B(y[2317]), .Z(n12080) );
  ANDN U4841 ( .B(y[2314]), .A(x[2314]), .Z(n12083) );
  ANDN U4842 ( .B(y[2313]), .A(x[2313]), .Z(n12084) );
  NANDN U4843 ( .A(x[2312]), .B(y[2312]), .Z(n24730) );
  ANDN U4844 ( .B(y[2307]), .A(x[2307]), .Z(n12089) );
  ANDN U4845 ( .B(x[2307]), .A(y[2307]), .Z(n24721) );
  ANDN U4846 ( .B(x[2306]), .A(y[2306]), .Z(n24715) );
  NOR U4847 ( .A(n24721), .B(n24715), .Z(n16616) );
  ANDN U4848 ( .B(y[2306]), .A(x[2306]), .Z(n16611) );
  NOR U4849 ( .A(n12089), .B(n16611), .Z(n24716) );
  ANDN U4850 ( .B(y[2305]), .A(x[2305]), .Z(n16612) );
  ANDN U4851 ( .B(y[2304]), .A(x[2304]), .Z(n12091) );
  NOR U4852 ( .A(n16612), .B(n12091), .Z(n24710) );
  ANDN U4853 ( .B(y[2303]), .A(x[2303]), .Z(n12092) );
  ANDN U4854 ( .B(y[2302]), .A(x[2302]), .Z(n16601) );
  NOR U4855 ( .A(n12092), .B(n16601), .Z(n24706) );
  ANDN U4856 ( .B(y[2300]), .A(x[2300]), .Z(n16596) );
  NANDN U4857 ( .A(x[2301]), .B(y[2301]), .Z(n24702) );
  NANDN U4858 ( .A(y[2300]), .B(x[2300]), .Z(n24701) );
  NANDN U4859 ( .A(y[2299]), .B(x[2299]), .Z(n24697) );
  ANDN U4860 ( .B(y[2299]), .A(x[2299]), .Z(n16595) );
  NANDN U4861 ( .A(y[2297]), .B(x[2297]), .Z(n16588) );
  NANDN U4862 ( .A(y[2298]), .B(x[2298]), .Z(n12095) );
  NAND U4863 ( .A(n16588), .B(n12095), .Z(n24693) );
  NANDN U4864 ( .A(y[2296]), .B(x[2296]), .Z(n16589) );
  ANDN U4865 ( .B(x[2295]), .A(y[2295]), .Z(n12097) );
  ANDN U4866 ( .B(n16589), .A(n12097), .Z(n24688) );
  ANDN U4867 ( .B(y[2294]), .A(x[2294]), .Z(n12099) );
  ANDN U4868 ( .B(x[2293]), .A(y[2293]), .Z(n16578) );
  NANDN U4869 ( .A(y[2294]), .B(x[2294]), .Z(n24684) );
  NANDN U4870 ( .A(x[2292]), .B(y[2292]), .Z(n12100) );
  ANDN U4871 ( .B(y[2293]), .A(x[2293]), .Z(n12098) );
  ANDN U4872 ( .B(n12100), .A(n12098), .Z(n8768) );
  XNOR U4873 ( .A(y[2292]), .B(x[2292]), .Z(n8766) );
  NANDN U4874 ( .A(y[2291]), .B(x[2291]), .Z(n24676) );
  NANDN U4875 ( .A(y[2289]), .B(x[2289]), .Z(n2888) );
  NANDN U4876 ( .A(y[2290]), .B(x[2290]), .Z(n2887) );
  AND U4877 ( .A(n2888), .B(n2887), .Z(n24672) );
  NANDN U4878 ( .A(y[2288]), .B(x[2288]), .Z(n2890) );
  NANDN U4879 ( .A(y[2287]), .B(x[2287]), .Z(n2889) );
  AND U4880 ( .A(n2890), .B(n2889), .Z(n24668) );
  ANDN U4881 ( .B(y[2285]), .A(x[2285]), .Z(n8749) );
  NANDN U4882 ( .A(x[2284]), .B(y[2284]), .Z(n2891) );
  NANDN U4883 ( .A(n8749), .B(n2891), .Z(n24663) );
  NANDN U4884 ( .A(x[2282]), .B(y[2282]), .Z(n2895) );
  ANDN U4885 ( .B(x[2282]), .A(y[2282]), .Z(n2892) );
  NOR U4886 ( .A(n2892), .B(x[2281]), .Z(n2893) );
  NAND U4887 ( .A(n2893), .B(y[2281]), .Z(n2894) );
  NAND U4888 ( .A(n2895), .B(n2894), .Z(n16563) );
  NANDN U4889 ( .A(x[2283]), .B(y[2283]), .Z(n16567) );
  NANDN U4890 ( .A(n16563), .B(n16567), .Z(n24657) );
  XNOR U4891 ( .A(y[2270]), .B(x[2270]), .Z(n2896) );
  NANDN U4892 ( .A(y[2269]), .B(x[2269]), .Z(n16540) );
  NAND U4893 ( .A(n2896), .B(n16540), .Z(n24631) );
  NANDN U4894 ( .A(x[2266]), .B(y[2266]), .Z(n2897) );
  ANDN U4895 ( .B(y[2267]), .A(x[2267]), .Z(n12103) );
  ANDN U4896 ( .B(n2897), .A(n12103), .Z(n24624) );
  NANDN U4897 ( .A(y[2263]), .B(x[2263]), .Z(n24618) );
  NANDN U4898 ( .A(y[2262]), .B(x[2262]), .Z(n2899) );
  NANDN U4899 ( .A(y[2261]), .B(x[2261]), .Z(n2898) );
  AND U4900 ( .A(n2899), .B(n2898), .Z(n24614) );
  NANDN U4901 ( .A(y[2260]), .B(x[2260]), .Z(n2900) );
  ANDN U4902 ( .B(x[2259]), .A(y[2259]), .Z(n16520) );
  ANDN U4903 ( .B(n2900), .A(n16520), .Z(n24610) );
  NANDN U4904 ( .A(y[2249]), .B(x[2249]), .Z(n24591) );
  NANDN U4905 ( .A(x[2245]), .B(y[2245]), .Z(n24580) );
  ANDN U4906 ( .B(y[2244]), .A(x[2244]), .Z(n16478) );
  ANDN U4907 ( .B(n24580), .A(n16478), .Z(n8680) );
  NANDN U4908 ( .A(x[2242]), .B(y[2242]), .Z(n24573) );
  IV U4909 ( .A(x[2241]), .Z(n12112) );
  NAND U4910 ( .A(y[2241]), .B(n12112), .Z(n12110) );
  NANDN U4911 ( .A(x[2240]), .B(y[2240]), .Z(n16468) );
  NAND U4912 ( .A(n12110), .B(n16468), .Z(n24569) );
  NANDN U4913 ( .A(x[2239]), .B(y[2239]), .Z(n20251) );
  NANDN U4914 ( .A(x[2237]), .B(y[2237]), .Z(n24561) );
  NANDN U4915 ( .A(x[2238]), .B(y[2238]), .Z(n20252) );
  NAND U4916 ( .A(n24561), .B(n20252), .Z(n12116) );
  NANDN U4917 ( .A(x[2236]), .B(y[2236]), .Z(n24557) );
  NANDN U4918 ( .A(n12116), .B(n24557), .Z(n12119) );
  ANDN U4919 ( .B(x[2236]), .A(y[2236]), .Z(n12115) );
  NANDN U4920 ( .A(y[2235]), .B(x[2235]), .Z(n24554) );
  NANDN U4921 ( .A(x[2234]), .B(y[2234]), .Z(n16461) );
  NANDN U4922 ( .A(x[2235]), .B(y[2235]), .Z(n12120) );
  NAND U4923 ( .A(n16461), .B(n12120), .Z(n24552) );
  NANDN U4924 ( .A(x[2232]), .B(y[2232]), .Z(n2902) );
  NANDN U4925 ( .A(x[2233]), .B(y[2233]), .Z(n2901) );
  NAND U4926 ( .A(n2902), .B(n2901), .Z(n24549) );
  NANDN U4927 ( .A(x[2231]), .B(y[2231]), .Z(n24544) );
  IV U4928 ( .A(x[2227]), .Z(n20254) );
  NAND U4929 ( .A(y[2227]), .B(n20254), .Z(n24533) );
  NANDN U4930 ( .A(x[2228]), .B(y[2228]), .Z(n24537) );
  NAND U4931 ( .A(n24533), .B(n24537), .Z(n16444) );
  NANDN U4932 ( .A(y[2225]), .B(x[2225]), .Z(n24526) );
  NANDN U4933 ( .A(x[2220]), .B(y[2220]), .Z(n2903) );
  ANDN U4934 ( .B(y[2221]), .A(x[2221]), .Z(n16433) );
  ANDN U4935 ( .B(n2903), .A(n16433), .Z(n24514) );
  NANDN U4936 ( .A(y[2218]), .B(x[2218]), .Z(n20256) );
  NANDN U4937 ( .A(y[2217]), .B(x[2217]), .Z(n20255) );
  NAND U4938 ( .A(n20256), .B(n20255), .Z(n16427) );
  NANDN U4939 ( .A(x[2217]), .B(y[2217]), .Z(n2904) );
  NANDN U4940 ( .A(x[2216]), .B(y[2216]), .Z(n24505) );
  NAND U4941 ( .A(n2904), .B(n24505), .Z(n16424) );
  NANDN U4942 ( .A(x[2212]), .B(y[2212]), .Z(n2906) );
  NANDN U4943 ( .A(x[2213]), .B(y[2213]), .Z(n2905) );
  NAND U4944 ( .A(n2906), .B(n2905), .Z(n24496) );
  NANDN U4945 ( .A(y[2211]), .B(x[2211]), .Z(n12122) );
  IV U4946 ( .A(y[2212]), .Z(n12121) );
  NAND U4947 ( .A(n12121), .B(x[2212]), .Z(n2907) );
  NAND U4948 ( .A(n12122), .B(n2907), .Z(n8616) );
  ANDN U4949 ( .B(x[2210]), .A(y[2210]), .Z(n12124) );
  NANDN U4950 ( .A(x[2206]), .B(y[2206]), .Z(n2909) );
  NANDN U4951 ( .A(x[2207]), .B(y[2207]), .Z(n2908) );
  NAND U4952 ( .A(n2909), .B(n2908), .Z(n24485) );
  NANDN U4953 ( .A(x[2204]), .B(y[2204]), .Z(n2910) );
  NANDN U4954 ( .A(x[2205]), .B(y[2205]), .Z(n16411) );
  NAND U4955 ( .A(n2910), .B(n16411), .Z(n8599) );
  NANDN U4956 ( .A(x[2203]), .B(y[2203]), .Z(n2911) );
  NANDN U4957 ( .A(n8599), .B(n2911), .Z(n24480) );
  NANDN U4958 ( .A(y[2201]), .B(x[2201]), .Z(n24474) );
  NANDN U4959 ( .A(y[2200]), .B(x[2200]), .Z(n24468) );
  NAND U4960 ( .A(n24474), .B(n24468), .Z(n16403) );
  NANDN U4961 ( .A(x[2199]), .B(y[2199]), .Z(n2913) );
  NANDN U4962 ( .A(x[2198]), .B(y[2198]), .Z(n2912) );
  NAND U4963 ( .A(n2913), .B(n2912), .Z(n24466) );
  NANDN U4964 ( .A(y[2197]), .B(x[2197]), .Z(n2915) );
  NANDN U4965 ( .A(y[2198]), .B(x[2198]), .Z(n2914) );
  NAND U4966 ( .A(n2915), .B(n2914), .Z(n24465) );
  NANDN U4967 ( .A(x[2195]), .B(y[2195]), .Z(n2917) );
  NANDN U4968 ( .A(x[2196]), .B(y[2196]), .Z(n2916) );
  NAND U4969 ( .A(n2917), .B(n2916), .Z(n24459) );
  ANDN U4970 ( .B(x[2195]), .A(y[2195]), .Z(n12135) );
  ANDN U4971 ( .B(x[2194]), .A(y[2194]), .Z(n12134) );
  NANDN U4972 ( .A(y[2192]), .B(x[2192]), .Z(n16389) );
  NANDN U4973 ( .A(y[2191]), .B(x[2191]), .Z(n16381) );
  NAND U4974 ( .A(n16389), .B(n16381), .Z(n24449) );
  NANDN U4975 ( .A(y[2188]), .B(x[2188]), .Z(n24441) );
  NANDN U4976 ( .A(y[2187]), .B(x[2187]), .Z(n2919) );
  NANDN U4977 ( .A(y[2186]), .B(x[2186]), .Z(n2918) );
  NAND U4978 ( .A(n2919), .B(n2918), .Z(n24437) );
  NANDN U4979 ( .A(x[2186]), .B(y[2186]), .Z(n20258) );
  NANDN U4980 ( .A(x[2185]), .B(y[2185]), .Z(n20257) );
  NAND U4981 ( .A(n20258), .B(n20257), .Z(n16372) );
  NANDN U4982 ( .A(y[2185]), .B(x[2185]), .Z(n2920) );
  NANDN U4983 ( .A(y[2184]), .B(x[2184]), .Z(n24431) );
  NAND U4984 ( .A(n2920), .B(n24431), .Z(n16370) );
  IV U4985 ( .A(x[2181]), .Z(n12137) );
  ANDN U4986 ( .B(y[2180]), .A(x[2180]), .Z(n24420) );
  ANDN U4987 ( .B(x[2180]), .A(y[2180]), .Z(n12141) );
  IV U4988 ( .A(x[2176]), .Z(n16348) );
  NAND U4989 ( .A(n16348), .B(y[2176]), .Z(n2922) );
  NANDN U4990 ( .A(x[2177]), .B(y[2177]), .Z(n2921) );
  NAND U4991 ( .A(n2922), .B(n2921), .Z(n24413) );
  IV U4992 ( .A(y[2173]), .Z(n16335) );
  NAND U4993 ( .A(n16335), .B(x[2173]), .Z(n2924) );
  NANDN U4994 ( .A(y[2174]), .B(x[2174]), .Z(n2923) );
  NAND U4995 ( .A(n2924), .B(n2923), .Z(n24406) );
  NANDN U4996 ( .A(y[2171]), .B(x[2171]), .Z(n12143) );
  NANDN U4997 ( .A(y[2172]), .B(x[2172]), .Z(n2925) );
  NAND U4998 ( .A(n12143), .B(n2925), .Z(n24403) );
  NANDN U4999 ( .A(y[2169]), .B(x[2169]), .Z(n16322) );
  NANDN U5000 ( .A(y[2170]), .B(x[2170]), .Z(n12142) );
  NAND U5001 ( .A(n16322), .B(n12142), .Z(n24399) );
  ANDN U5002 ( .B(y[2168]), .A(x[2168]), .Z(n16319) );
  NANDN U5003 ( .A(x[2169]), .B(y[2169]), .Z(n24397) );
  NANDN U5004 ( .A(y[2168]), .B(x[2168]), .Z(n24394) );
  ANDN U5005 ( .B(x[2166]), .A(y[2166]), .Z(n12145) );
  NANDN U5006 ( .A(y[2165]), .B(x[2165]), .Z(n24386) );
  NANDN U5007 ( .A(x[2162]), .B(y[2162]), .Z(n2927) );
  NANDN U5008 ( .A(x[2163]), .B(y[2163]), .Z(n2926) );
  NAND U5009 ( .A(n2927), .B(n2926), .Z(n24381) );
  ANDN U5010 ( .B(x[2161]), .A(y[2161]), .Z(n16299) );
  XOR U5011 ( .A(x[2162]), .B(y[2162]), .Z(n16303) );
  NOR U5012 ( .A(n16299), .B(n16303), .Z(n24378) );
  NANDN U5013 ( .A(y[2159]), .B(x[2159]), .Z(n24370) );
  NANDN U5014 ( .A(y[2158]), .B(x[2158]), .Z(n24365) );
  NAND U5015 ( .A(n24370), .B(n24365), .Z(n16296) );
  NANDN U5016 ( .A(y[2157]), .B(x[2157]), .Z(n24366) );
  NANDN U5017 ( .A(x[2156]), .B(y[2156]), .Z(n12148) );
  NANDN U5018 ( .A(x[2157]), .B(y[2157]), .Z(n16293) );
  NAND U5019 ( .A(n12148), .B(n16293), .Z(n24363) );
  NANDN U5020 ( .A(y[2156]), .B(x[2156]), .Z(n12146) );
  NANDN U5021 ( .A(x[2149]), .B(y[2149]), .Z(n2929) );
  NANDN U5022 ( .A(x[2148]), .B(y[2148]), .Z(n2928) );
  AND U5023 ( .A(n2929), .B(n2928), .Z(n24346) );
  NANDN U5024 ( .A(x[2147]), .B(y[2147]), .Z(n2931) );
  NANDN U5025 ( .A(x[2146]), .B(y[2146]), .Z(n2930) );
  AND U5026 ( .A(n2931), .B(n2930), .Z(n24342) );
  NANDN U5027 ( .A(x[2145]), .B(y[2145]), .Z(n2933) );
  NANDN U5028 ( .A(x[2144]), .B(y[2144]), .Z(n2932) );
  AND U5029 ( .A(n2933), .B(n2932), .Z(n24338) );
  NANDN U5030 ( .A(x[2143]), .B(y[2143]), .Z(n24334) );
  NANDN U5031 ( .A(y[2140]), .B(x[2140]), .Z(n2935) );
  NANDN U5032 ( .A(y[2141]), .B(x[2141]), .Z(n2934) );
  NAND U5033 ( .A(n2935), .B(n2934), .Z(n12155) );
  NANDN U5034 ( .A(y[2139]), .B(x[2139]), .Z(n12150) );
  NANDN U5035 ( .A(x[2140]), .B(y[2140]), .Z(n2936) );
  NANDN U5036 ( .A(n12150), .B(n2936), .Z(n8483) );
  NANDN U5037 ( .A(x[2138]), .B(y[2138]), .Z(n2938) );
  NANDN U5038 ( .A(x[2139]), .B(y[2139]), .Z(n2937) );
  NAND U5039 ( .A(n2937), .B(n2936), .Z(n12153) );
  ANDN U5040 ( .B(n2938), .A(n12153), .Z(n24326) );
  NANDN U5041 ( .A(y[2137]), .B(x[2137]), .Z(n24325) );
  ANDN U5042 ( .B(x[2138]), .A(y[2138]), .Z(n12151) );
  ANDN U5043 ( .B(n24325), .A(n12151), .Z(n8480) );
  IV U5044 ( .A(y[2135]), .Z(n16252) );
  NAND U5045 ( .A(n16252), .B(x[2135]), .Z(n2939) );
  NANDN U5046 ( .A(y[2136]), .B(x[2136]), .Z(n16259) );
  AND U5047 ( .A(n2939), .B(n16259), .Z(n24320) );
  ANDN U5048 ( .B(x[2133]), .A(y[2133]), .Z(n12157) );
  NANDN U5049 ( .A(y[2131]), .B(x[2131]), .Z(n24308) );
  ANDN U5050 ( .B(x[2132]), .A(y[2132]), .Z(n12158) );
  ANDN U5051 ( .B(n24308), .A(n12158), .Z(n8470) );
  ANDN U5052 ( .B(y[2131]), .A(x[2131]), .Z(n16243) );
  NANDN U5053 ( .A(y[2129]), .B(x[2129]), .Z(n2940) );
  NANDN U5054 ( .A(y[2130]), .B(x[2130]), .Z(n12159) );
  NAND U5055 ( .A(n2940), .B(n12159), .Z(n24305) );
  ANDN U5056 ( .B(y[2126]), .A(x[2126]), .Z(n8454) );
  NANDN U5057 ( .A(y[2125]), .B(x[2125]), .Z(n16224) );
  OR U5058 ( .A(n8454), .B(n16224), .Z(n8461) );
  NANDN U5059 ( .A(x[2121]), .B(y[2121]), .Z(n2942) );
  NANDN U5060 ( .A(x[2120]), .B(y[2120]), .Z(n2941) );
  NAND U5061 ( .A(n2942), .B(n2941), .Z(n24287) );
  NANDN U5062 ( .A(x[2119]), .B(y[2119]), .Z(n2944) );
  NANDN U5063 ( .A(x[2118]), .B(y[2118]), .Z(n2943) );
  AND U5064 ( .A(n2944), .B(n2943), .Z(n24282) );
  NANDN U5065 ( .A(y[2117]), .B(x[2117]), .Z(n2945) );
  NANDN U5066 ( .A(y[2118]), .B(x[2118]), .Z(n24281) );
  NAND U5067 ( .A(n2945), .B(n24281), .Z(n16208) );
  NANDN U5068 ( .A(x[2116]), .B(y[2116]), .Z(n24273) );
  IV U5069 ( .A(x[2117]), .Z(n24276) );
  NAND U5070 ( .A(n24276), .B(y[2117]), .Z(n2946) );
  NAND U5071 ( .A(n24273), .B(n2946), .Z(n16204) );
  ANDN U5072 ( .B(y[2115]), .A(x[2115]), .Z(n16202) );
  ANDN U5073 ( .B(y[2114]), .A(x[2114]), .Z(n16196) );
  NOR U5074 ( .A(n16202), .B(n16196), .Z(n24269) );
  NANDN U5075 ( .A(x[2113]), .B(y[2113]), .Z(n24265) );
  ANDN U5076 ( .B(x[2111]), .A(y[2111]), .Z(n12161) );
  NANDN U5077 ( .A(x[2110]), .B(y[2110]), .Z(n24257) );
  NANDN U5078 ( .A(y[2109]), .B(x[2109]), .Z(n24255) );
  ANDN U5079 ( .B(x[2110]), .A(y[2110]), .Z(n12160) );
  ANDN U5080 ( .B(n24255), .A(n12160), .Z(n8428) );
  NANDN U5081 ( .A(y[2108]), .B(x[2108]), .Z(n2947) );
  ANDN U5082 ( .B(x[2107]), .A(y[2107]), .Z(n16182) );
  ANDN U5083 ( .B(n2947), .A(n16182), .Z(n24251) );
  NANDN U5084 ( .A(y[2106]), .B(x[2106]), .Z(n2949) );
  NANDN U5085 ( .A(y[2105]), .B(x[2105]), .Z(n2948) );
  NAND U5086 ( .A(n2949), .B(n2948), .Z(n24248) );
  XOR U5087 ( .A(x[2102]), .B(y[2102]), .Z(n16174) );
  NANDN U5088 ( .A(y[2101]), .B(x[2101]), .Z(n2950) );
  NANDN U5089 ( .A(n16174), .B(n2950), .Z(n24240) );
  NANDN U5090 ( .A(y[2100]), .B(x[2100]), .Z(n12162) );
  NANDN U5091 ( .A(x[2097]), .B(y[2097]), .Z(n20259) );
  NANDN U5092 ( .A(x[2091]), .B(y[2091]), .Z(n2952) );
  NANDN U5093 ( .A(x[2090]), .B(y[2090]), .Z(n2951) );
  NAND U5094 ( .A(n2952), .B(n2951), .Z(n16148) );
  NANDN U5095 ( .A(x[2088]), .B(y[2088]), .Z(n24214) );
  NANDN U5096 ( .A(y[2087]), .B(x[2087]), .Z(n2953) );
  NANDN U5097 ( .A(y[2088]), .B(x[2088]), .Z(n16143) );
  NAND U5098 ( .A(n2953), .B(n16143), .Z(n24211) );
  ANDN U5099 ( .B(y[2084]), .A(x[2084]), .Z(n12178) );
  NANDN U5100 ( .A(x[2085]), .B(y[2085]), .Z(n24205) );
  NANDN U5101 ( .A(y[2084]), .B(x[2084]), .Z(n24203) );
  NANDN U5102 ( .A(y[2083]), .B(x[2083]), .Z(n12179) );
  AND U5103 ( .A(n24203), .B(n12179), .Z(n8379) );
  XNOR U5104 ( .A(x[2083]), .B(y[2083]), .Z(n8377) );
  NANDN U5105 ( .A(x[2082]), .B(y[2082]), .Z(n24198) );
  NANDN U5106 ( .A(x[2080]), .B(y[2080]), .Z(n2954) );
  NANDN U5107 ( .A(x[2081]), .B(y[2081]), .Z(n16124) );
  AND U5108 ( .A(n2954), .B(n16124), .Z(n24193) );
  IV U5109 ( .A(y[2079]), .Z(n12181) );
  NAND U5110 ( .A(n12181), .B(x[2079]), .Z(n16120) );
  NANDN U5111 ( .A(y[2080]), .B(x[2080]), .Z(n16122) );
  NAND U5112 ( .A(n16120), .B(n16122), .Z(n24191) );
  ANDN U5113 ( .B(y[2078]), .A(x[2078]), .Z(n16115) );
  NANDN U5114 ( .A(x[2075]), .B(y[2075]), .Z(n8359) );
  NANDN U5115 ( .A(x[2074]), .B(y[2074]), .Z(n2955) );
  NAND U5116 ( .A(n8359), .B(n2955), .Z(n24181) );
  NANDN U5117 ( .A(y[2073]), .B(x[2073]), .Z(n24179) );
  ANDN U5118 ( .B(x[2069]), .A(y[2069]), .Z(n12183) );
  NANDN U5119 ( .A(x[2068]), .B(y[2068]), .Z(n24163) );
  ANDN U5120 ( .B(x[2068]), .A(y[2068]), .Z(n12182) );
  ANDN U5121 ( .B(x[2067]), .A(y[2067]), .Z(n24162) );
  IV U5122 ( .A(y[2065]), .Z(n16089) );
  NAND U5123 ( .A(n16089), .B(x[2065]), .Z(n2956) );
  NANDN U5124 ( .A(y[2066]), .B(x[2066]), .Z(n16094) );
  NAND U5125 ( .A(n2956), .B(n16094), .Z(n24158) );
  IV U5126 ( .A(x[2064]), .Z(n12184) );
  NAND U5127 ( .A(n12184), .B(y[2064]), .Z(n16086) );
  NANDN U5128 ( .A(x[2065]), .B(y[2065]), .Z(n2957) );
  AND U5129 ( .A(n16086), .B(n2957), .Z(n24155) );
  ANDN U5130 ( .B(y[2062]), .A(x[2062]), .Z(n12187) );
  NANDN U5131 ( .A(x[2063]), .B(y[2063]), .Z(n24151) );
  NANDN U5132 ( .A(x[2060]), .B(y[2060]), .Z(n24143) );
  ANDN U5133 ( .B(y[2061]), .A(x[2061]), .Z(n12186) );
  ANDN U5134 ( .B(n24143), .A(n12186), .Z(n8334) );
  NANDN U5135 ( .A(y[2060]), .B(x[2060]), .Z(n12188) );
  NANDN U5136 ( .A(x[2058]), .B(y[2058]), .Z(n2958) );
  IV U5137 ( .A(x[2059]), .Z(n12190) );
  NAND U5138 ( .A(n12190), .B(y[2059]), .Z(n12189) );
  NAND U5139 ( .A(n2958), .B(n12189), .Z(n24140) );
  NANDN U5140 ( .A(y[2058]), .B(x[2058]), .Z(n2959) );
  NANDN U5141 ( .A(y[2057]), .B(x[2057]), .Z(n16068) );
  NAND U5142 ( .A(n2959), .B(n16068), .Z(n24135) );
  NANDN U5143 ( .A(x[2054]), .B(y[2054]), .Z(n24129) );
  NANDN U5144 ( .A(y[2053]), .B(x[2053]), .Z(n24128) );
  NANDN U5145 ( .A(y[2050]), .B(x[2050]), .Z(n2961) );
  NANDN U5146 ( .A(y[2049]), .B(x[2049]), .Z(n2960) );
  NAND U5147 ( .A(n2961), .B(n2960), .Z(n24120) );
  NANDN U5148 ( .A(x[2049]), .B(y[2049]), .Z(n2963) );
  NANDN U5149 ( .A(x[2048]), .B(y[2048]), .Z(n2962) );
  AND U5150 ( .A(n2963), .B(n2962), .Z(n24117) );
  NANDN U5151 ( .A(x[2047]), .B(y[2047]), .Z(n2965) );
  NANDN U5152 ( .A(x[2046]), .B(y[2046]), .Z(n2964) );
  AND U5153 ( .A(n2965), .B(n2964), .Z(n24113) );
  NANDN U5154 ( .A(x[2043]), .B(y[2043]), .Z(n2967) );
  ANDN U5155 ( .B(y[2045]), .A(x[2045]), .Z(n16046) );
  NANDN U5156 ( .A(x[2044]), .B(y[2044]), .Z(n2966) );
  NANDN U5157 ( .A(n16046), .B(n2966), .Z(n8307) );
  ANDN U5158 ( .B(n2967), .A(n8307), .Z(n24109) );
  NANDN U5159 ( .A(x[2042]), .B(y[2042]), .Z(n8303) );
  ANDN U5160 ( .B(x[2041]), .A(y[2041]), .Z(n16035) );
  ANDN U5161 ( .B(x[2042]), .A(y[2042]), .Z(n16039) );
  ANDN U5162 ( .B(x[2040]), .A(y[2040]), .Z(n16036) );
  IV U5163 ( .A(y[2037]), .Z(n12194) );
  NAND U5164 ( .A(n12194), .B(x[2037]), .Z(n16026) );
  IV U5165 ( .A(y[2038]), .Z(n12193) );
  NAND U5166 ( .A(n12193), .B(x[2038]), .Z(n12192) );
  NAND U5167 ( .A(n16026), .B(n12192), .Z(n24099) );
  NANDN U5168 ( .A(x[2037]), .B(y[2037]), .Z(n2968) );
  ANDN U5169 ( .B(y[2036]), .A(x[2036]), .Z(n12195) );
  ANDN U5170 ( .B(n2968), .A(n12195), .Z(n24097) );
  ANDN U5171 ( .B(x[2035]), .A(y[2035]), .Z(n12197) );
  ANDN U5172 ( .B(x[2034]), .A(y[2034]), .Z(n12196) );
  IV U5173 ( .A(x[2030]), .Z(n16003) );
  NAND U5174 ( .A(n16003), .B(y[2030]), .Z(n2970) );
  NANDN U5175 ( .A(x[2031]), .B(y[2031]), .Z(n2969) );
  NAND U5176 ( .A(n2970), .B(n2969), .Z(n24082) );
  NANDN U5177 ( .A(y[2029]), .B(x[2029]), .Z(n15999) );
  NANDN U5178 ( .A(y[2030]), .B(x[2030]), .Z(n2971) );
  NAND U5179 ( .A(n15999), .B(n2971), .Z(n24079) );
  NANDN U5180 ( .A(y[2028]), .B(x[2028]), .Z(n24075) );
  ANDN U5181 ( .B(x[2027]), .A(y[2027]), .Z(n12200) );
  ANDN U5182 ( .B(n24075), .A(n12200), .Z(n8291) );
  ANDN U5183 ( .B(x[2020]), .A(y[2020]), .Z(n24055) );
  ANDN U5184 ( .B(y[2019]), .A(x[2019]), .Z(n12202) );
  NANDN U5185 ( .A(x[2018]), .B(y[2018]), .Z(n24050) );
  NANDN U5186 ( .A(y[2015]), .B(x[2015]), .Z(n8261) );
  XNOR U5187 ( .A(y[2015]), .B(x[2015]), .Z(n2973) );
  NANDN U5188 ( .A(x[2014]), .B(y[2014]), .Z(n2972) );
  NAND U5189 ( .A(n2973), .B(n2972), .Z(n2974) );
  NAND U5190 ( .A(n8261), .B(n2974), .Z(n2976) );
  NANDN U5191 ( .A(x[2016]), .B(y[2016]), .Z(n2975) );
  AND U5192 ( .A(n2976), .B(n2975), .Z(n2978) );
  NANDN U5193 ( .A(x[2017]), .B(y[2017]), .Z(n2977) );
  AND U5194 ( .A(n2978), .B(n2977), .Z(n24043) );
  NANDN U5195 ( .A(x[2010]), .B(y[2010]), .Z(n2980) );
  NANDN U5196 ( .A(x[2011]), .B(y[2011]), .Z(n2979) );
  AND U5197 ( .A(n2980), .B(n2979), .Z(n24029) );
  NANDN U5198 ( .A(x[2009]), .B(y[2009]), .Z(n2982) );
  NANDN U5199 ( .A(x[2008]), .B(y[2008]), .Z(n2981) );
  AND U5200 ( .A(n2982), .B(n2981), .Z(n24025) );
  NANDN U5201 ( .A(x[2007]), .B(y[2007]), .Z(n2984) );
  NANDN U5202 ( .A(x[2006]), .B(y[2006]), .Z(n2983) );
  AND U5203 ( .A(n2984), .B(n2983), .Z(n24021) );
  NANDN U5204 ( .A(x[2002]), .B(y[2002]), .Z(n2986) );
  NANDN U5205 ( .A(x[2003]), .B(y[2003]), .Z(n2985) );
  NAND U5206 ( .A(n2986), .B(n2985), .Z(n15954) );
  XOR U5207 ( .A(x[2002]), .B(y[2002]), .Z(n15953) );
  NANDN U5208 ( .A(y[2001]), .B(x[2001]), .Z(n2987) );
  NANDN U5209 ( .A(n15953), .B(n2987), .Z(n15950) );
  ANDN U5210 ( .B(y[2001]), .A(x[2001]), .Z(n15952) );
  NANDN U5211 ( .A(y[1999]), .B(x[1999]), .Z(n15945) );
  ANDN U5212 ( .B(x[2000]), .A(y[2000]), .Z(n15949) );
  ANDN U5213 ( .B(n15945), .A(n15949), .Z(n8236) );
  XNOR U5214 ( .A(x[1999]), .B(y[1999]), .Z(n8234) );
  NANDN U5215 ( .A(x[1998]), .B(y[1998]), .Z(n24005) );
  NANDN U5216 ( .A(x[1996]), .B(y[1996]), .Z(n12208) );
  NANDN U5217 ( .A(x[1997]), .B(y[1997]), .Z(n15942) );
  AND U5218 ( .A(n12208), .B(n15942), .Z(n24001) );
  NANDN U5219 ( .A(x[1994]), .B(y[1994]), .Z(n15935) );
  IV U5220 ( .A(x[1995]), .Z(n12209) );
  NAND U5221 ( .A(n12209), .B(y[1995]), .Z(n12207) );
  NAND U5222 ( .A(n15935), .B(n12207), .Z(n23998) );
  NANDN U5223 ( .A(y[1994]), .B(x[1994]), .Z(n2988) );
  NANDN U5224 ( .A(y[1993]), .B(x[1993]), .Z(n12210) );
  NAND U5225 ( .A(n2988), .B(n12210), .Z(n23996) );
  ANDN U5226 ( .B(y[1992]), .A(x[1992]), .Z(n12212) );
  ANDN U5227 ( .B(y[1991]), .A(x[1991]), .Z(n12211) );
  NANDN U5228 ( .A(y[1987]), .B(x[1987]), .Z(n2990) );
  NANDN U5229 ( .A(y[1988]), .B(x[1988]), .Z(n2989) );
  NAND U5230 ( .A(n2990), .B(n2989), .Z(n23978) );
  NANDN U5231 ( .A(y[1986]), .B(x[1986]), .Z(n23973) );
  ANDN U5232 ( .B(x[1985]), .A(y[1985]), .Z(n12214) );
  NANDN U5233 ( .A(y[1983]), .B(x[1983]), .Z(n23966) );
  ANDN U5234 ( .B(x[1984]), .A(y[1984]), .Z(n12213) );
  ANDN U5235 ( .B(n23966), .A(n12213), .Z(n8207) );
  NANDN U5236 ( .A(x[1982]), .B(y[1982]), .Z(n12217) );
  NANDN U5237 ( .A(x[1983]), .B(y[1983]), .Z(n15915) );
  NAND U5238 ( .A(n12217), .B(n15915), .Z(n23964) );
  NANDN U5239 ( .A(y[1979]), .B(x[1979]), .Z(n15902) );
  XNOR U5240 ( .A(y[1980]), .B(x[1980]), .Z(n2991) );
  NAND U5241 ( .A(n15902), .B(n2991), .Z(n23958) );
  NANDN U5242 ( .A(y[1978]), .B(x[1978]), .Z(n23954) );
  NANDN U5243 ( .A(y[1977]), .B(x[1977]), .Z(n2993) );
  NANDN U5244 ( .A(y[1976]), .B(x[1976]), .Z(n2992) );
  NAND U5245 ( .A(n2993), .B(n2992), .Z(n23950) );
  NANDN U5246 ( .A(y[1975]), .B(x[1975]), .Z(n23945) );
  IV U5247 ( .A(y[1974]), .Z(n20263) );
  NAND U5248 ( .A(n20263), .B(x[1974]), .Z(n23944) );
  AND U5249 ( .A(n23945), .B(n23944), .Z(n15896) );
  NANDN U5250 ( .A(x[1974]), .B(y[1974]), .Z(n2994) );
  NANDN U5251 ( .A(x[1973]), .B(y[1973]), .Z(n23937) );
  NAND U5252 ( .A(n2994), .B(n23937), .Z(n15895) );
  ANDN U5253 ( .B(x[1973]), .A(y[1973]), .Z(n23940) );
  ANDN U5254 ( .B(x[1972]), .A(y[1972]), .Z(n23936) );
  NOR U5255 ( .A(n23940), .B(n23936), .Z(n15892) );
  NANDN U5256 ( .A(y[1971]), .B(x[1971]), .Z(n12218) );
  AND U5257 ( .A(n15892), .B(n12218), .Z(n8187) );
  XNOR U5258 ( .A(x[1971]), .B(y[1971]), .Z(n8185) );
  NANDN U5259 ( .A(x[1970]), .B(y[1970]), .Z(n23929) );
  NANDN U5260 ( .A(x[1968]), .B(y[1968]), .Z(n2996) );
  NANDN U5261 ( .A(x[1969]), .B(y[1969]), .Z(n2995) );
  NAND U5262 ( .A(n2996), .B(n2995), .Z(n23925) );
  NANDN U5263 ( .A(x[1967]), .B(y[1967]), .Z(n2998) );
  NANDN U5264 ( .A(x[1966]), .B(y[1966]), .Z(n2997) );
  NAND U5265 ( .A(n2998), .B(n2997), .Z(n23922) );
  NANDN U5266 ( .A(x[1962]), .B(y[1962]), .Z(n3000) );
  NANDN U5267 ( .A(x[1963]), .B(y[1963]), .Z(n2999) );
  NAND U5268 ( .A(n3000), .B(n2999), .Z(n15874) );
  NANDN U5269 ( .A(y[1961]), .B(x[1961]), .Z(n3001) );
  XOR U5270 ( .A(x[1962]), .B(y[1962]), .Z(n15877) );
  ANDN U5271 ( .B(n3001), .A(n15877), .Z(n23910) );
  ANDN U5272 ( .B(y[1961]), .A(x[1961]), .Z(n15876) );
  NANDN U5273 ( .A(x[1960]), .B(y[1960]), .Z(n3002) );
  NANDN U5274 ( .A(n15876), .B(n3002), .Z(n3003) );
  NAND U5275 ( .A(n23910), .B(n3003), .Z(n3004) );
  NANDN U5276 ( .A(n15874), .B(n3004), .Z(n23913) );
  ANDN U5277 ( .B(x[1957]), .A(y[1957]), .Z(n12224) );
  NANDN U5278 ( .A(y[1951]), .B(x[1951]), .Z(n3005) );
  XNOR U5279 ( .A(x[1952]), .B(y[1952]), .Z(n12225) );
  AND U5280 ( .A(n3005), .B(n12225), .Z(n23890) );
  NANDN U5281 ( .A(y[1949]), .B(x[1949]), .Z(n15851) );
  ANDN U5282 ( .B(x[1950]), .A(y[1950]), .Z(n23886) );
  ANDN U5283 ( .B(n15851), .A(n23886), .Z(n23881) );
  NANDN U5284 ( .A(y[1947]), .B(x[1947]), .Z(n3007) );
  NANDN U5285 ( .A(y[1948]), .B(x[1948]), .Z(n3006) );
  NAND U5286 ( .A(n3007), .B(n3006), .Z(n23878) );
  NANDN U5287 ( .A(x[1947]), .B(y[1947]), .Z(n3009) );
  NANDN U5288 ( .A(x[1946]), .B(y[1946]), .Z(n3008) );
  AND U5289 ( .A(n3009), .B(n3008), .Z(n23875) );
  NANDN U5290 ( .A(x[1943]), .B(y[1943]), .Z(n3011) );
  NANDN U5291 ( .A(x[1942]), .B(y[1942]), .Z(n3010) );
  AND U5292 ( .A(n3011), .B(n3010), .Z(n23867) );
  NANDN U5293 ( .A(x[1939]), .B(y[1939]), .Z(n3013) );
  NANDN U5294 ( .A(x[1938]), .B(y[1938]), .Z(n3012) );
  AND U5295 ( .A(n3013), .B(n3012), .Z(n23859) );
  NANDN U5296 ( .A(x[1929]), .B(y[1929]), .Z(n23843) );
  ANDN U5297 ( .B(y[1930]), .A(x[1930]), .Z(n8101) );
  ANDN U5298 ( .B(n23843), .A(n8101), .Z(n15815) );
  NANDN U5299 ( .A(x[1928]), .B(y[1928]), .Z(n23839) );
  AND U5300 ( .A(n15815), .B(n23839), .Z(n8097) );
  IV U5301 ( .A(x[1932]), .Z(n15818) );
  NAND U5302 ( .A(n15818), .B(y[1932]), .Z(n15823) );
  NANDN U5303 ( .A(x[1933]), .B(y[1933]), .Z(n15828) );
  NAND U5304 ( .A(n15823), .B(n15828), .Z(n8104) );
  ANDN U5305 ( .B(y[1931]), .A(x[1931]), .Z(n15819) );
  NOR U5306 ( .A(n8104), .B(n15819), .Z(n8095) );
  NANDN U5307 ( .A(y[1926]), .B(x[1926]), .Z(n23833) );
  NANDN U5308 ( .A(x[1923]), .B(y[1923]), .Z(n23823) );
  IV U5309 ( .A(x[1924]), .Z(n20265) );
  NAND U5310 ( .A(y[1924]), .B(n20265), .Z(n23828) );
  NAND U5311 ( .A(n23823), .B(n23828), .Z(n15806) );
  ANDN U5312 ( .B(y[1922]), .A(x[1922]), .Z(n12230) );
  NANDN U5313 ( .A(y[1921]), .B(x[1921]), .Z(n23818) );
  ANDN U5314 ( .B(y[1919]), .A(x[1919]), .Z(n23809) );
  NANDN U5315 ( .A(x[1920]), .B(y[1920]), .Z(n23815) );
  NANDN U5316 ( .A(n23809), .B(n23815), .Z(n3014) );
  ANDN U5317 ( .B(x[1920]), .A(y[1920]), .Z(n3016) );
  ANDN U5318 ( .B(n3014), .A(n3016), .Z(n15801) );
  ANDN U5319 ( .B(y[1921]), .A(x[1921]), .Z(n12229) );
  NANDN U5320 ( .A(y[1919]), .B(x[1919]), .Z(n3015) );
  NANDN U5321 ( .A(n3016), .B(n3015), .Z(n23814) );
  NANDN U5322 ( .A(y[1916]), .B(x[1916]), .Z(n3018) );
  NANDN U5323 ( .A(y[1915]), .B(x[1915]), .Z(n3017) );
  NAND U5324 ( .A(n3018), .B(n3017), .Z(n12234) );
  NANDN U5325 ( .A(y[1913]), .B(x[1913]), .Z(n23800) );
  NANDN U5326 ( .A(y[1912]), .B(x[1912]), .Z(n3020) );
  NANDN U5327 ( .A(y[1911]), .B(x[1911]), .Z(n3019) );
  NAND U5328 ( .A(n3020), .B(n3019), .Z(n23796) );
  NANDN U5329 ( .A(y[1910]), .B(x[1910]), .Z(n3022) );
  NANDN U5330 ( .A(y[1909]), .B(x[1909]), .Z(n3021) );
  NAND U5331 ( .A(n3022), .B(n3021), .Z(n23792) );
  ANDN U5332 ( .B(x[1908]), .A(y[1908]), .Z(n23787) );
  ANDN U5333 ( .B(x[1903]), .A(y[1903]), .Z(n12236) );
  NANDN U5334 ( .A(x[1903]), .B(y[1903]), .Z(n23774) );
  NANDN U5335 ( .A(x[1902]), .B(y[1902]), .Z(n15771) );
  AND U5336 ( .A(n23774), .B(n15771), .Z(n8045) );
  XNOR U5337 ( .A(y[1902]), .B(x[1902]), .Z(n8043) );
  XNOR U5338 ( .A(x[1901]), .B(y[1901]), .Z(n8040) );
  ANDN U5339 ( .B(y[1900]), .A(x[1900]), .Z(n23766) );
  ANDN U5340 ( .B(x[1900]), .A(y[1900]), .Z(n12238) );
  NANDN U5341 ( .A(x[1897]), .B(y[1897]), .Z(n15761) );
  NANDN U5342 ( .A(y[1895]), .B(x[1895]), .Z(n15754) );
  IV U5343 ( .A(y[1896]), .Z(n12244) );
  NAND U5344 ( .A(n12244), .B(x[1896]), .Z(n12242) );
  NAND U5345 ( .A(n15754), .B(n12242), .Z(n23755) );
  NANDN U5346 ( .A(y[1894]), .B(x[1894]), .Z(n23751) );
  NANDN U5347 ( .A(y[1893]), .B(x[1893]), .Z(n23747) );
  NAND U5348 ( .A(n23751), .B(n23747), .Z(n8029) );
  NANDN U5349 ( .A(x[1890]), .B(y[1890]), .Z(n15734) );
  NANDN U5350 ( .A(x[1891]), .B(y[1891]), .Z(n3023) );
  NAND U5351 ( .A(n15734), .B(n3023), .Z(n23742) );
  NANDN U5352 ( .A(y[1888]), .B(x[1888]), .Z(n3025) );
  NANDN U5353 ( .A(y[1887]), .B(x[1887]), .Z(n3024) );
  AND U5354 ( .A(n3025), .B(n3024), .Z(n23735) );
  ANDN U5355 ( .B(x[1881]), .A(y[1881]), .Z(n15720) );
  NANDN U5356 ( .A(x[1881]), .B(y[1881]), .Z(n23725) );
  NANDN U5357 ( .A(x[1880]), .B(y[1880]), .Z(n12249) );
  AND U5358 ( .A(n23725), .B(n12249), .Z(n8001) );
  XNOR U5359 ( .A(y[1880]), .B(x[1880]), .Z(n7999) );
  NANDN U5360 ( .A(y[1879]), .B(x[1879]), .Z(n23719) );
  ANDN U5361 ( .B(y[1879]), .A(x[1879]), .Z(n12250) );
  NANDN U5362 ( .A(y[1878]), .B(x[1878]), .Z(n12251) );
  IV U5363 ( .A(x[1876]), .Z(n15709) );
  NAND U5364 ( .A(n15709), .B(y[1876]), .Z(n3026) );
  IV U5365 ( .A(x[1877]), .Z(n12253) );
  NAND U5366 ( .A(n12253), .B(y[1877]), .Z(n12252) );
  NAND U5367 ( .A(n3026), .B(n12252), .Z(n23714) );
  NANDN U5368 ( .A(x[1871]), .B(y[1871]), .Z(n15693) );
  NANDN U5369 ( .A(x[1870]), .B(y[1870]), .Z(n15687) );
  AND U5370 ( .A(n15693), .B(n15687), .Z(n23699) );
  NANDN U5371 ( .A(x[1869]), .B(y[1869]), .Z(n20268) );
  NANDN U5372 ( .A(x[1867]), .B(y[1867]), .Z(n3028) );
  NANDN U5373 ( .A(x[1866]), .B(y[1866]), .Z(n3027) );
  NAND U5374 ( .A(n3028), .B(n3027), .Z(n23688) );
  NANDN U5375 ( .A(y[1866]), .B(x[1866]), .Z(n3030) );
  NANDN U5376 ( .A(y[1865]), .B(x[1865]), .Z(n3029) );
  NAND U5377 ( .A(n3030), .B(n3029), .Z(n23685) );
  ANDN U5378 ( .B(x[1861]), .A(y[1861]), .Z(n15671) );
  NANDN U5379 ( .A(x[1861]), .B(y[1861]), .Z(n23679) );
  NANDN U5380 ( .A(x[1860]), .B(y[1860]), .Z(n12257) );
  AND U5381 ( .A(n23679), .B(n12257), .Z(n7965) );
  XNOR U5382 ( .A(y[1860]), .B(x[1860]), .Z(n7963) );
  XNOR U5383 ( .A(x[1859]), .B(y[1859]), .Z(n7960) );
  ANDN U5384 ( .B(x[1858]), .A(y[1858]), .Z(n12259) );
  NANDN U5385 ( .A(y[1857]), .B(x[1857]), .Z(n23670) );
  NANDN U5386 ( .A(y[1856]), .B(x[1856]), .Z(n3031) );
  NANDN U5387 ( .A(y[1855]), .B(x[1855]), .Z(n15660) );
  NAND U5388 ( .A(n3031), .B(n15660), .Z(n23666) );
  NANDN U5389 ( .A(x[1852]), .B(y[1852]), .Z(n3033) );
  NANDN U5390 ( .A(x[1853]), .B(y[1853]), .Z(n3032) );
  NAND U5391 ( .A(n3033), .B(n3032), .Z(n12264) );
  ANDN U5392 ( .B(y[1851]), .A(x[1851]), .Z(n12261) );
  NANDN U5393 ( .A(y[1849]), .B(x[1849]), .Z(n3034) );
  NANDN U5394 ( .A(y[1850]), .B(x[1850]), .Z(n12265) );
  NAND U5395 ( .A(n3034), .B(n12265), .Z(n23653) );
  NANDN U5396 ( .A(x[1845]), .B(y[1845]), .Z(n3035) );
  NANDN U5397 ( .A(x[1846]), .B(y[1846]), .Z(n7935) );
  NAND U5398 ( .A(n3035), .B(n7935), .Z(n15641) );
  NANDN U5399 ( .A(x[1844]), .B(y[1844]), .Z(n3036) );
  NANDN U5400 ( .A(n15641), .B(n3036), .Z(n23644) );
  ANDN U5401 ( .B(y[1841]), .A(x[1841]), .Z(n15633) );
  ANDN U5402 ( .B(y[1840]), .A(x[1840]), .Z(n15625) );
  NOR U5403 ( .A(n15633), .B(n15625), .Z(n23633) );
  NANDN U5404 ( .A(x[1839]), .B(y[1839]), .Z(n23627) );
  ANDN U5405 ( .B(x[1836]), .A(y[1836]), .Z(n12271) );
  ANDN U5406 ( .B(x[1831]), .A(y[1831]), .Z(n12273) );
  ANDN U5407 ( .B(x[1829]), .A(y[1829]), .Z(n23598) );
  ANDN U5408 ( .B(x[1830]), .A(y[1830]), .Z(n12272) );
  NANDN U5409 ( .A(x[1828]), .B(y[1828]), .Z(n12274) );
  NANDN U5410 ( .A(x[1829]), .B(y[1829]), .Z(n15610) );
  NAND U5411 ( .A(n12274), .B(n15610), .Z(n23597) );
  NANDN U5412 ( .A(x[1827]), .B(y[1827]), .Z(n23589) );
  ANDN U5413 ( .B(x[1823]), .A(y[1823]), .Z(n23577) );
  ANDN U5414 ( .B(y[1823]), .A(x[1823]), .Z(n12276) );
  NANDN U5415 ( .A(x[1818]), .B(y[1818]), .Z(n3038) );
  NANDN U5416 ( .A(x[1819]), .B(y[1819]), .Z(n3037) );
  AND U5417 ( .A(n3038), .B(n3037), .Z(n23566) );
  NANDN U5418 ( .A(y[1817]), .B(x[1817]), .Z(n15581) );
  NANDN U5419 ( .A(y[1818]), .B(x[1818]), .Z(n3039) );
  NAND U5420 ( .A(n15581), .B(n3039), .Z(n23565) );
  NANDN U5421 ( .A(y[1813]), .B(x[1813]), .Z(n15574) );
  IV U5422 ( .A(y[1814]), .Z(n12283) );
  NAND U5423 ( .A(n12283), .B(x[1814]), .Z(n12282) );
  NAND U5424 ( .A(n15574), .B(n12282), .Z(n23553) );
  NANDN U5425 ( .A(x[1812]), .B(y[1812]), .Z(n3041) );
  NANDN U5426 ( .A(x[1813]), .B(y[1813]), .Z(n3040) );
  NAND U5427 ( .A(n3041), .B(n3040), .Z(n23551) );
  NANDN U5428 ( .A(x[1811]), .B(y[1811]), .Z(n23546) );
  ANDN U5429 ( .B(y[1810]), .A(x[1810]), .Z(n12286) );
  ANDN U5430 ( .B(n23546), .A(n12286), .Z(n7883) );
  NANDN U5431 ( .A(y[1807]), .B(x[1807]), .Z(n3042) );
  ANDN U5432 ( .B(x[1808]), .A(y[1808]), .Z(n12287) );
  ANDN U5433 ( .B(n3042), .A(n12287), .Z(n23536) );
  NANDN U5434 ( .A(x[1806]), .B(y[1806]), .Z(n3044) );
  NANDN U5435 ( .A(x[1807]), .B(y[1807]), .Z(n3043) );
  NAND U5436 ( .A(n3044), .B(n3043), .Z(n23535) );
  NANDN U5437 ( .A(y[1806]), .B(x[1806]), .Z(n3045) );
  ANDN U5438 ( .B(x[1805]), .A(y[1805]), .Z(n12288) );
  ANDN U5439 ( .B(n3045), .A(n12288), .Z(n23532) );
  ANDN U5440 ( .B(y[1804]), .A(x[1804]), .Z(n12290) );
  ANDN U5441 ( .B(y[1805]), .A(x[1805]), .Z(n23530) );
  ANDN U5442 ( .B(x[1803]), .A(y[1803]), .Z(n15544) );
  ANDN U5443 ( .B(y[1799]), .A(x[1799]), .Z(n7859) );
  NANDN U5444 ( .A(x[1798]), .B(y[1798]), .Z(n3046) );
  NANDN U5445 ( .A(n7859), .B(n3046), .Z(n23515) );
  NANDN U5446 ( .A(x[1796]), .B(y[1796]), .Z(n3048) );
  NANDN U5447 ( .A(x[1797]), .B(y[1797]), .Z(n3047) );
  NAND U5448 ( .A(n3048), .B(n3047), .Z(n15535) );
  ANDN U5449 ( .B(y[1795]), .A(x[1795]), .Z(n15532) );
  NANDN U5450 ( .A(x[1791]), .B(y[1791]), .Z(n23496) );
  AND U5451 ( .A(n23496), .B(n12294), .Z(n7844) );
  XNOR U5452 ( .A(x[1790]), .B(y[1790]), .Z(n7842) );
  XNOR U5453 ( .A(x[1789]), .B(y[1789]), .Z(n7839) );
  NANDN U5454 ( .A(y[1787]), .B(x[1787]), .Z(n23486) );
  ANDN U5455 ( .B(x[1788]), .A(y[1788]), .Z(n12296) );
  ANDN U5456 ( .B(n23486), .A(n12296), .Z(n7836) );
  NANDN U5457 ( .A(x[1786]), .B(y[1786]), .Z(n3050) );
  NANDN U5458 ( .A(x[1787]), .B(y[1787]), .Z(n3049) );
  NAND U5459 ( .A(n3050), .B(n3049), .Z(n23485) );
  NANDN U5460 ( .A(y[1786]), .B(x[1786]), .Z(n3052) );
  NANDN U5461 ( .A(y[1785]), .B(x[1785]), .Z(n3051) );
  AND U5462 ( .A(n3052), .B(n3051), .Z(n23482) );
  NANDN U5463 ( .A(x[1783]), .B(y[1783]), .Z(n23476) );
  ANDN U5464 ( .B(y[1782]), .A(x[1782]), .Z(n12298) );
  ANDN U5465 ( .B(n23476), .A(n12298), .Z(n7828) );
  NANDN U5466 ( .A(x[1778]), .B(y[1778]), .Z(n3053) );
  NANDN U5467 ( .A(x[1779]), .B(y[1779]), .Z(n15524) );
  NAND U5468 ( .A(n3053), .B(n15524), .Z(n23464) );
  NANDN U5469 ( .A(y[1777]), .B(x[1777]), .Z(n15516) );
  IV U5470 ( .A(y[1778]), .Z(n15519) );
  NAND U5471 ( .A(n15519), .B(x[1778]), .Z(n3054) );
  NAND U5472 ( .A(n15516), .B(n3054), .Z(n23463) );
  NANDN U5473 ( .A(y[1775]), .B(x[1775]), .Z(n3056) );
  NANDN U5474 ( .A(y[1776]), .B(x[1776]), .Z(n3055) );
  NAND U5475 ( .A(n3056), .B(n3055), .Z(n12302) );
  ANDN U5476 ( .B(x[1774]), .A(y[1774]), .Z(n12299) );
  NANDN U5477 ( .A(y[1773]), .B(x[1773]), .Z(n23454) );
  NANDN U5478 ( .A(x[1771]), .B(y[1771]), .Z(n3058) );
  NANDN U5479 ( .A(x[1770]), .B(y[1770]), .Z(n3057) );
  NAND U5480 ( .A(n3058), .B(n3057), .Z(n23449) );
  NANDN U5481 ( .A(x[1762]), .B(y[1762]), .Z(n3060) );
  NANDN U5482 ( .A(x[1761]), .B(y[1761]), .Z(n3059) );
  NAND U5483 ( .A(n3060), .B(n3059), .Z(n23429) );
  ANDN U5484 ( .B(x[1761]), .A(y[1761]), .Z(n15490) );
  NANDN U5485 ( .A(x[1760]), .B(y[1760]), .Z(n23425) );
  ANDN U5486 ( .B(x[1760]), .A(y[1760]), .Z(n15489) );
  NANDN U5487 ( .A(x[1758]), .B(y[1758]), .Z(n3062) );
  NANDN U5488 ( .A(x[1759]), .B(y[1759]), .Z(n3061) );
  NAND U5489 ( .A(n3062), .B(n3061), .Z(n23421) );
  NANDN U5490 ( .A(y[1755]), .B(x[1755]), .Z(n3064) );
  NANDN U5491 ( .A(y[1756]), .B(x[1756]), .Z(n3063) );
  NAND U5492 ( .A(n3064), .B(n3063), .Z(n12308) );
  NANDN U5493 ( .A(x[1754]), .B(y[1754]), .Z(n3065) );
  ANDN U5494 ( .B(y[1755]), .A(x[1755]), .Z(n12306) );
  ANDN U5495 ( .B(n3065), .A(n12306), .Z(n23413) );
  ANDN U5496 ( .B(x[1754]), .A(y[1754]), .Z(n12305) );
  NANDN U5497 ( .A(x[1752]), .B(y[1752]), .Z(n12310) );
  NANDN U5498 ( .A(x[1753]), .B(y[1753]), .Z(n15481) );
  NAND U5499 ( .A(n12310), .B(n15481), .Z(n23409) );
  NANDN U5500 ( .A(x[1745]), .B(y[1745]), .Z(n3067) );
  NANDN U5501 ( .A(x[1744]), .B(y[1744]), .Z(n3066) );
  AND U5502 ( .A(n3067), .B(n3066), .Z(n23392) );
  NANDN U5503 ( .A(x[1742]), .B(y[1742]), .Z(n3069) );
  NANDN U5504 ( .A(x[1743]), .B(y[1743]), .Z(n3068) );
  NAND U5505 ( .A(n3069), .B(n3068), .Z(n23388) );
  NANDN U5506 ( .A(x[1738]), .B(y[1738]), .Z(n23380) );
  ANDN U5507 ( .B(y[1739]), .A(x[1739]), .Z(n15446) );
  ANDN U5508 ( .B(n23380), .A(n15446), .Z(n7739) );
  NANDN U5509 ( .A(x[1737]), .B(y[1737]), .Z(n3071) );
  NANDN U5510 ( .A(x[1736]), .B(y[1736]), .Z(n3070) );
  AND U5511 ( .A(n3071), .B(n3070), .Z(n23376) );
  NANDN U5512 ( .A(x[1735]), .B(y[1735]), .Z(n3073) );
  NANDN U5513 ( .A(x[1734]), .B(y[1734]), .Z(n3072) );
  AND U5514 ( .A(n3073), .B(n3072), .Z(n23372) );
  NANDN U5515 ( .A(x[1733]), .B(y[1733]), .Z(n3075) );
  NANDN U5516 ( .A(x[1732]), .B(y[1732]), .Z(n3074) );
  AND U5517 ( .A(n3075), .B(n3074), .Z(n23368) );
  NANDN U5518 ( .A(x[1722]), .B(y[1722]), .Z(n3077) );
  NANDN U5519 ( .A(x[1723]), .B(y[1723]), .Z(n3076) );
  NAND U5520 ( .A(n3077), .B(n3076), .Z(n23349) );
  ANDN U5521 ( .B(x[1719]), .A(y[1719]), .Z(n12312) );
  NANDN U5522 ( .A(x[1718]), .B(y[1718]), .Z(n23337) );
  NANDN U5523 ( .A(y[1713]), .B(x[1713]), .Z(n12315) );
  XNOR U5524 ( .A(x[1713]), .B(y[1713]), .Z(n7674) );
  XNOR U5525 ( .A(y[1712]), .B(x[1712]), .Z(n7671) );
  XNOR U5526 ( .A(y[1711]), .B(x[1711]), .Z(n7668) );
  ANDN U5527 ( .B(x[1710]), .A(y[1710]), .Z(n12320) );
  ANDN U5528 ( .B(y[1709]), .A(x[1709]), .Z(n23314) );
  NANDN U5529 ( .A(x[1710]), .B(y[1710]), .Z(n23320) );
  NANDN U5530 ( .A(n23314), .B(n23320), .Z(n15407) );
  NANDN U5531 ( .A(x[1708]), .B(y[1708]), .Z(n23315) );
  NANDN U5532 ( .A(y[1705]), .B(x[1705]), .Z(n3079) );
  NANDN U5533 ( .A(y[1706]), .B(x[1706]), .Z(n3078) );
  NAND U5534 ( .A(n3079), .B(n3078), .Z(n12324) );
  ANDN U5535 ( .B(x[1704]), .A(y[1704]), .Z(n12321) );
  NANDN U5536 ( .A(x[1702]), .B(y[1702]), .Z(n15398) );
  NANDN U5537 ( .A(x[1703]), .B(y[1703]), .Z(n12325) );
  NAND U5538 ( .A(n15398), .B(n12325), .Z(n23302) );
  NANDN U5539 ( .A(y[1697]), .B(x[1697]), .Z(n3080) );
  NANDN U5540 ( .A(y[1698]), .B(x[1698]), .Z(n12327) );
  AND U5541 ( .A(n3080), .B(n12327), .Z(n23292) );
  NANDN U5542 ( .A(x[1696]), .B(y[1696]), .Z(n15375) );
  NANDN U5543 ( .A(x[1697]), .B(y[1697]), .Z(n15382) );
  NAND U5544 ( .A(n15375), .B(n15382), .Z(n23290) );
  ANDN U5545 ( .B(y[1695]), .A(x[1695]), .Z(n15377) );
  ANDN U5546 ( .B(y[1693]), .A(x[1693]), .Z(n15367) );
  IV U5547 ( .A(n15367), .Z(n23283) );
  NANDN U5548 ( .A(y[1692]), .B(x[1692]), .Z(n23280) );
  NANDN U5549 ( .A(y[1691]), .B(x[1691]), .Z(n15362) );
  AND U5550 ( .A(n23280), .B(n15362), .Z(n7633) );
  XNOR U5551 ( .A(x[1691]), .B(y[1691]), .Z(n7631) );
  NANDN U5552 ( .A(x[1690]), .B(y[1690]), .Z(n23274) );
  NANDN U5553 ( .A(x[1688]), .B(y[1688]), .Z(n3081) );
  NANDN U5554 ( .A(x[1689]), .B(y[1689]), .Z(n12332) );
  NAND U5555 ( .A(n3081), .B(n12332), .Z(n23271) );
  NANDN U5556 ( .A(y[1687]), .B(x[1687]), .Z(n12334) );
  NANDN U5557 ( .A(y[1688]), .B(x[1688]), .Z(n3082) );
  NAND U5558 ( .A(n12334), .B(n3082), .Z(n23269) );
  NANDN U5559 ( .A(x[1687]), .B(y[1687]), .Z(n15352) );
  NANDN U5560 ( .A(y[1685]), .B(x[1685]), .Z(n15345) );
  IV U5561 ( .A(y[1686]), .Z(n12335) );
  NAND U5562 ( .A(n12335), .B(x[1686]), .Z(n12333) );
  NAND U5563 ( .A(n15345), .B(n12333), .Z(n23265) );
  NANDN U5564 ( .A(x[1685]), .B(y[1685]), .Z(n23262) );
  ANDN U5565 ( .B(y[1684]), .A(x[1684]), .Z(n12337) );
  ANDN U5566 ( .B(n23262), .A(n12337), .Z(n7622) );
  ANDN U5567 ( .B(x[1683]), .A(y[1683]), .Z(n23256) );
  ANDN U5568 ( .B(y[1683]), .A(x[1683]), .Z(n12336) );
  NANDN U5569 ( .A(x[1682]), .B(y[1682]), .Z(n23254) );
  NANDN U5570 ( .A(x[1678]), .B(y[1678]), .Z(n3083) );
  NANDN U5571 ( .A(x[1679]), .B(y[1679]), .Z(n12338) );
  AND U5572 ( .A(n3083), .B(n12338), .Z(n23246) );
  NANDN U5573 ( .A(y[1677]), .B(x[1677]), .Z(n15322) );
  NANDN U5574 ( .A(y[1678]), .B(x[1678]), .Z(n3084) );
  NAND U5575 ( .A(n15322), .B(n3084), .Z(n20272) );
  NANDN U5576 ( .A(y[1675]), .B(x[1675]), .Z(n23240) );
  ANDN U5577 ( .B(x[1676]), .A(y[1676]), .Z(n20270) );
  IV U5578 ( .A(n20270), .Z(n15321) );
  AND U5579 ( .A(n23240), .B(n15321), .Z(n7607) );
  ANDN U5580 ( .B(y[1672]), .A(x[1672]), .Z(n12344) );
  ANDN U5581 ( .B(x[1671]), .A(y[1671]), .Z(n12346) );
  NANDN U5582 ( .A(y[1672]), .B(x[1672]), .Z(n23233) );
  NANDN U5583 ( .A(x[1670]), .B(y[1670]), .Z(n12347) );
  ANDN U5584 ( .B(y[1671]), .A(x[1671]), .Z(n12343) );
  ANDN U5585 ( .B(n12347), .A(n12343), .Z(n7598) );
  XNOR U5586 ( .A(y[1670]), .B(x[1670]), .Z(n7596) );
  NANDN U5587 ( .A(y[1669]), .B(x[1669]), .Z(n23224) );
  ANDN U5588 ( .B(y[1669]), .A(x[1669]), .Z(n12348) );
  NANDN U5589 ( .A(y[1668]), .B(x[1668]), .Z(n12349) );
  NANDN U5590 ( .A(x[1666]), .B(y[1666]), .Z(n15294) );
  IV U5591 ( .A(x[1667]), .Z(n12351) );
  NAND U5592 ( .A(n12351), .B(y[1667]), .Z(n12350) );
  NAND U5593 ( .A(n15294), .B(n12350), .Z(n23219) );
  IV U5594 ( .A(y[1658]), .Z(n20274) );
  NAND U5595 ( .A(n20274), .B(x[1658]), .Z(n3085) );
  NANDN U5596 ( .A(y[1659]), .B(x[1659]), .Z(n23211) );
  NAND U5597 ( .A(n3085), .B(n23211), .Z(n15278) );
  NANDN U5598 ( .A(y[1656]), .B(x[1656]), .Z(n3087) );
  NANDN U5599 ( .A(y[1655]), .B(x[1655]), .Z(n3086) );
  AND U5600 ( .A(n3087), .B(n3086), .Z(n3088) );
  NANDN U5601 ( .A(y[1657]), .B(x[1657]), .Z(n7571) );
  NAND U5602 ( .A(n3088), .B(n7571), .Z(n23201) );
  NANDN U5603 ( .A(x[1655]), .B(y[1655]), .Z(n3090) );
  NANDN U5604 ( .A(x[1654]), .B(y[1654]), .Z(n3089) );
  NAND U5605 ( .A(n3090), .B(n3089), .Z(n23199) );
  ANDN U5606 ( .B(y[1652]), .A(x[1652]), .Z(n12353) );
  NANDN U5607 ( .A(x[1653]), .B(y[1653]), .Z(n23194) );
  NANDN U5608 ( .A(y[1652]), .B(x[1652]), .Z(n23192) );
  NANDN U5609 ( .A(y[1651]), .B(x[1651]), .Z(n15264) );
  AND U5610 ( .A(n23192), .B(n15264), .Z(n7562) );
  XNOR U5611 ( .A(x[1651]), .B(y[1651]), .Z(n7560) );
  NANDN U5612 ( .A(y[1649]), .B(x[1649]), .Z(n15260) );
  ANDN U5613 ( .B(x[1650]), .A(y[1650]), .Z(n15263) );
  ANDN U5614 ( .B(n15260), .A(n15263), .Z(n7557) );
  XNOR U5615 ( .A(x[1649]), .B(y[1649]), .Z(n7555) );
  NANDN U5616 ( .A(x[1648]), .B(y[1648]), .Z(n23182) );
  NANDN U5617 ( .A(y[1647]), .B(x[1647]), .Z(n23180) );
  ANDN U5618 ( .B(x[1648]), .A(y[1648]), .Z(n15259) );
  ANDN U5619 ( .B(n23180), .A(n15259), .Z(n7552) );
  NANDN U5620 ( .A(x[1642]), .B(y[1642]), .Z(n3092) );
  NANDN U5621 ( .A(x[1643]), .B(y[1643]), .Z(n3091) );
  NAND U5622 ( .A(n3092), .B(n3091), .Z(n12359) );
  IV U5623 ( .A(y[1639]), .Z(n15237) );
  NAND U5624 ( .A(n15237), .B(x[1639]), .Z(n3093) );
  NANDN U5625 ( .A(y[1640]), .B(x[1640]), .Z(n15244) );
  NAND U5626 ( .A(n3093), .B(n15244), .Z(n23164) );
  ANDN U5627 ( .B(x[1638]), .A(y[1638]), .Z(n23158) );
  NANDN U5628 ( .A(y[1636]), .B(x[1636]), .Z(n23153) );
  ANDN U5629 ( .B(x[1637]), .A(y[1637]), .Z(n23161) );
  ANDN U5630 ( .B(n23153), .A(n23161), .Z(n15232) );
  NANDN U5631 ( .A(x[1635]), .B(y[1635]), .Z(n3099) );
  XNOR U5632 ( .A(x[1635]), .B(y[1635]), .Z(n3095) );
  NANDN U5633 ( .A(y[1634]), .B(x[1634]), .Z(n3094) );
  NAND U5634 ( .A(n3095), .B(n3094), .Z(n3096) );
  NAND U5635 ( .A(n3099), .B(n3096), .Z(n23154) );
  NANDN U5636 ( .A(x[1634]), .B(y[1634]), .Z(n3098) );
  NANDN U5637 ( .A(x[1633]), .B(y[1633]), .Z(n3097) );
  AND U5638 ( .A(n3098), .B(n3097), .Z(n3100) );
  NAND U5639 ( .A(n3100), .B(n3099), .Z(n15228) );
  NANDN U5640 ( .A(y[1633]), .B(x[1633]), .Z(n7524) );
  ANDN U5641 ( .B(y[1632]), .A(x[1632]), .Z(n12361) );
  NAND U5642 ( .A(n7524), .B(n12361), .Z(n3101) );
  NANDN U5643 ( .A(n15228), .B(n3101), .Z(n23151) );
  NANDN U5644 ( .A(x[1631]), .B(y[1631]), .Z(n23146) );
  ANDN U5645 ( .B(x[1629]), .A(y[1629]), .Z(n12363) );
  NANDN U5646 ( .A(y[1627]), .B(x[1627]), .Z(n23136) );
  ANDN U5647 ( .B(x[1628]), .A(y[1628]), .Z(n12362) );
  ANDN U5648 ( .B(n23136), .A(n12362), .Z(n7514) );
  NANDN U5649 ( .A(y[1626]), .B(x[1626]), .Z(n20279) );
  IV U5650 ( .A(y[1624]), .Z(n23125) );
  NAND U5651 ( .A(n23125), .B(x[1624]), .Z(n3102) );
  NANDN U5652 ( .A(y[1625]), .B(x[1625]), .Z(n20278) );
  AND U5653 ( .A(n3102), .B(n20278), .Z(n15214) );
  ANDN U5654 ( .B(x[1623]), .A(y[1623]), .Z(n15209) );
  XNOR U5655 ( .A(x[1622]), .B(y[1622]), .Z(n7503) );
  XNOR U5656 ( .A(y[1621]), .B(x[1621]), .Z(n7500) );
  ANDN U5657 ( .B(x[1620]), .A(y[1620]), .Z(n12366) );
  NANDN U5658 ( .A(x[1620]), .B(y[1620]), .Z(n3104) );
  NANDN U5659 ( .A(x[1619]), .B(y[1619]), .Z(n3103) );
  NAND U5660 ( .A(n3104), .B(n3103), .Z(n23114) );
  ANDN U5661 ( .B(x[1615]), .A(y[1615]), .Z(n12369) );
  NANDN U5662 ( .A(x[1614]), .B(y[1614]), .Z(n23101) );
  IV U5663 ( .A(y[1611]), .Z(n15187) );
  NAND U5664 ( .A(n15187), .B(x[1611]), .Z(n3106) );
  NANDN U5665 ( .A(y[1612]), .B(x[1612]), .Z(n3105) );
  NAND U5666 ( .A(n3106), .B(n3105), .Z(n23096) );
  NANDN U5667 ( .A(x[1608]), .B(y[1608]), .Z(n15181) );
  XNOR U5668 ( .A(y[1608]), .B(x[1608]), .Z(n7471) );
  XNOR U5669 ( .A(x[1607]), .B(y[1607]), .Z(n7468) );
  NANDN U5670 ( .A(x[1600]), .B(y[1600]), .Z(n3108) );
  NANDN U5671 ( .A(x[1599]), .B(y[1599]), .Z(n3107) );
  AND U5672 ( .A(n3108), .B(n3107), .Z(n23069) );
  XNOR U5673 ( .A(y[1595]), .B(x[1595]), .Z(n7432) );
  ANDN U5674 ( .B(x[1594]), .A(y[1594]), .Z(n12378) );
  NANDN U5675 ( .A(y[1590]), .B(x[1590]), .Z(n3109) );
  ANDN U5676 ( .B(x[1591]), .A(y[1591]), .Z(n7422) );
  ANDN U5677 ( .B(n3109), .A(n7422), .Z(n23047) );
  ANDN U5678 ( .B(y[1589]), .A(x[1589]), .Z(n15154) );
  NANDN U5679 ( .A(x[1588]), .B(y[1588]), .Z(n3111) );
  NANDN U5680 ( .A(x[1587]), .B(y[1587]), .Z(n3110) );
  NAND U5681 ( .A(n3111), .B(n3110), .Z(n23042) );
  NANDN U5682 ( .A(y[1583]), .B(x[1583]), .Z(n12380) );
  XNOR U5683 ( .A(x[1583]), .B(y[1583]), .Z(n7404) );
  NANDN U5684 ( .A(x[1582]), .B(y[1582]), .Z(n23029) );
  ANDN U5685 ( .B(x[1581]), .A(y[1581]), .Z(n12383) );
  ANDN U5686 ( .B(y[1581]), .A(x[1581]), .Z(n12384) );
  ANDN U5687 ( .B(x[1579]), .A(y[1579]), .Z(n15138) );
  NANDN U5688 ( .A(y[1580]), .B(x[1580]), .Z(n12382) );
  NANDN U5689 ( .A(n15138), .B(n12382), .Z(n3112) );
  NANDN U5690 ( .A(n3116), .B(n3112), .Z(n3113) );
  NANDN U5691 ( .A(n12383), .B(n3113), .Z(n3114) );
  ANDN U5692 ( .B(x[1582]), .A(y[1582]), .Z(n12381) );
  NOR U5693 ( .A(n3114), .B(n12381), .Z(n7401) );
  NANDN U5694 ( .A(x[1579]), .B(y[1579]), .Z(n3115) );
  NANDN U5695 ( .A(n3116), .B(n3115), .Z(n23025) );
  NANDN U5696 ( .A(y[1577]), .B(x[1577]), .Z(n3118) );
  NANDN U5697 ( .A(y[1576]), .B(x[1576]), .Z(n3117) );
  AND U5698 ( .A(n3118), .B(n3117), .Z(n23019) );
  ANDN U5699 ( .B(y[1572]), .A(x[1572]), .Z(n7384) );
  ANDN U5700 ( .B(x[1571]), .A(y[1571]), .Z(n12386) );
  ANDN U5701 ( .B(x[1570]), .A(y[1570]), .Z(n12387) );
  NANDN U5702 ( .A(y[1569]), .B(x[1569]), .Z(n23007) );
  ANDN U5703 ( .B(y[1565]), .A(x[1565]), .Z(n12394) );
  NANDN U5704 ( .A(y[1565]), .B(x[1565]), .Z(n3120) );
  NANDN U5705 ( .A(y[1564]), .B(x[1564]), .Z(n3119) );
  AND U5706 ( .A(n3120), .B(n3119), .Z(n22995) );
  NANDN U5707 ( .A(y[1563]), .B(x[1563]), .Z(n3122) );
  NANDN U5708 ( .A(y[1562]), .B(x[1562]), .Z(n3121) );
  AND U5709 ( .A(n3122), .B(n3121), .Z(n22991) );
  NANDN U5710 ( .A(x[1560]), .B(y[1560]), .Z(n15115) );
  XNOR U5711 ( .A(y[1560]), .B(x[1560]), .Z(n7372) );
  XNOR U5712 ( .A(x[1559]), .B(y[1559]), .Z(n7369) );
  ANDN U5713 ( .B(y[1557]), .A(x[1557]), .Z(n12400) );
  ANDN U5714 ( .B(x[1556]), .A(y[1556]), .Z(n22976) );
  NANDN U5715 ( .A(x[1552]), .B(y[1552]), .Z(n3124) );
  NANDN U5716 ( .A(x[1551]), .B(y[1551]), .Z(n3123) );
  AND U5717 ( .A(n3124), .B(n3123), .Z(n22965) );
  NANDN U5718 ( .A(y[1547]), .B(x[1547]), .Z(n15095) );
  XNOR U5719 ( .A(x[1547]), .B(y[1547]), .Z(n7337) );
  XNOR U5720 ( .A(y[1546]), .B(x[1546]), .Z(n7334) );
  ANDN U5721 ( .B(y[1544]), .A(x[1544]), .Z(n12408) );
  ANDN U5722 ( .B(x[1544]), .A(y[1544]), .Z(n15091) );
  ANDN U5723 ( .B(y[1542]), .A(x[1542]), .Z(n12410) );
  ANDN U5724 ( .B(y[1543]), .A(x[1543]), .Z(n22947) );
  ANDN U5725 ( .B(x[1542]), .A(y[1542]), .Z(n15086) );
  ANDN U5726 ( .B(y[1541]), .A(x[1541]), .Z(n12409) );
  NANDN U5727 ( .A(y[1541]), .B(x[1541]), .Z(n3126) );
  NANDN U5728 ( .A(y[1540]), .B(x[1540]), .Z(n3125) );
  AND U5729 ( .A(n3126), .B(n3125), .Z(n22941) );
  NANDN U5730 ( .A(y[1539]), .B(x[1539]), .Z(n3128) );
  NANDN U5731 ( .A(y[1538]), .B(x[1538]), .Z(n3127) );
  AND U5732 ( .A(n3128), .B(n3127), .Z(n22937) );
  ANDN U5733 ( .B(x[1531]), .A(y[1531]), .Z(n12419) );
  NANDN U5734 ( .A(y[1530]), .B(x[1530]), .Z(n12418) );
  XNOR U5735 ( .A(x[1530]), .B(y[1530]), .Z(n7299) );
  NANDN U5736 ( .A(x[1528]), .B(y[1528]), .Z(n3130) );
  NANDN U5737 ( .A(x[1527]), .B(y[1527]), .Z(n3129) );
  AND U5738 ( .A(n3130), .B(n3129), .Z(n22915) );
  ANDN U5739 ( .B(x[1521]), .A(y[1521]), .Z(n7273) );
  NANDN U5740 ( .A(y[1520]), .B(x[1520]), .Z(n3131) );
  NANDN U5741 ( .A(n7273), .B(n3131), .Z(n22902) );
  NANDN U5742 ( .A(x[1519]), .B(y[1519]), .Z(n22899) );
  NANDN U5743 ( .A(x[1518]), .B(y[1518]), .Z(n12420) );
  AND U5744 ( .A(n22899), .B(n12420), .Z(n7270) );
  NANDN U5745 ( .A(x[1514]), .B(y[1514]), .Z(n3133) );
  NANDN U5746 ( .A(x[1513]), .B(y[1513]), .Z(n3132) );
  AND U5747 ( .A(n3133), .B(n3132), .Z(n22887) );
  NANDN U5748 ( .A(x[1508]), .B(y[1508]), .Z(n15037) );
  NANDN U5749 ( .A(y[1509]), .B(x[1509]), .Z(n3138) );
  NANDN U5750 ( .A(n15037), .B(n3138), .Z(n3136) );
  NANDN U5751 ( .A(x[1510]), .B(y[1510]), .Z(n3135) );
  NANDN U5752 ( .A(x[1509]), .B(y[1509]), .Z(n3134) );
  AND U5753 ( .A(n3135), .B(n3134), .Z(n15040) );
  NAND U5754 ( .A(n3136), .B(n15040), .Z(n22880) );
  ANDN U5755 ( .B(x[1507]), .A(y[1507]), .Z(n12424) );
  NANDN U5756 ( .A(y[1508]), .B(x[1508]), .Z(n3137) );
  NAND U5757 ( .A(n3138), .B(n3137), .Z(n20284) );
  ANDN U5758 ( .B(x[1506]), .A(y[1506]), .Z(n12425) );
  NANDN U5759 ( .A(x[1502]), .B(y[1502]), .Z(n3140) );
  NANDN U5760 ( .A(x[1501]), .B(y[1501]), .Z(n3139) );
  AND U5761 ( .A(n3140), .B(n3139), .Z(n22867) );
  XNOR U5762 ( .A(y[1499]), .B(x[1499]), .Z(n7220) );
  ANDN U5763 ( .B(y[1498]), .A(x[1498]), .Z(n22860) );
  ANDN U5764 ( .B(x[1498]), .A(y[1498]), .Z(n12431) );
  NANDN U5765 ( .A(y[1497]), .B(x[1497]), .Z(n22857) );
  NANDN U5766 ( .A(x[1490]), .B(y[1490]), .Z(n12433) );
  XNOR U5767 ( .A(y[1490]), .B(x[1490]), .Z(n7198) );
  XNOR U5768 ( .A(x[1489]), .B(y[1489]), .Z(n7195) );
  XNOR U5769 ( .A(x[1487]), .B(y[1487]), .Z(n7188) );
  ANDN U5770 ( .B(x[1486]), .A(y[1486]), .Z(n12440) );
  NANDN U5771 ( .A(y[1485]), .B(x[1485]), .Z(n22829) );
  NANDN U5772 ( .A(x[1483]), .B(y[1483]), .Z(n22823) );
  NANDN U5773 ( .A(y[1481]), .B(x[1481]), .Z(n3142) );
  NANDN U5774 ( .A(y[1480]), .B(x[1480]), .Z(n3141) );
  NAND U5775 ( .A(n3142), .B(n3141), .Z(n22818) );
  NANDN U5776 ( .A(y[1477]), .B(x[1477]), .Z(n12446) );
  XNOR U5777 ( .A(x[1477]), .B(y[1477]), .Z(n7165) );
  NANDN U5778 ( .A(y[1475]), .B(x[1475]), .Z(n12449) );
  ANDN U5779 ( .B(x[1476]), .A(y[1476]), .Z(n12447) );
  ANDN U5780 ( .B(n12449), .A(n12447), .Z(n7162) );
  XNOR U5781 ( .A(x[1475]), .B(y[1475]), .Z(n7160) );
  IV U5782 ( .A(x[1474]), .Z(n12450) );
  ANDN U5783 ( .B(y[1473]), .A(x[1473]), .Z(n12451) );
  ANDN U5784 ( .B(y[1472]), .A(x[1472]), .Z(n14979) );
  IV U5785 ( .A(x[1472]), .Z(n22797) );
  NOR U5786 ( .A(n22797), .B(y[1472]), .Z(n12453) );
  NANDN U5787 ( .A(x[1471]), .B(y[1471]), .Z(n22794) );
  NANDN U5788 ( .A(y[1469]), .B(x[1469]), .Z(n3144) );
  NANDN U5789 ( .A(y[1468]), .B(x[1468]), .Z(n3143) );
  NAND U5790 ( .A(n3144), .B(n3143), .Z(n22789) );
  NANDN U5791 ( .A(y[1467]), .B(x[1467]), .Z(n3146) );
  NANDN U5792 ( .A(y[1466]), .B(x[1466]), .Z(n3145) );
  NAND U5793 ( .A(n3146), .B(n3145), .Z(n22784) );
  ANDN U5794 ( .B(x[1463]), .A(y[1463]), .Z(n14966) );
  NANDN U5795 ( .A(y[1461]), .B(x[1461]), .Z(n22771) );
  ANDN U5796 ( .B(x[1462]), .A(y[1462]), .Z(n14965) );
  ANDN U5797 ( .B(n22771), .A(n14965), .Z(n7127) );
  ANDN U5798 ( .B(y[1461]), .A(x[1461]), .Z(n14962) );
  NANDN U5799 ( .A(x[1460]), .B(y[1460]), .Z(n14958) );
  NANDN U5800 ( .A(n14962), .B(n14958), .Z(n22770) );
  ANDN U5801 ( .B(x[1460]), .A(y[1460]), .Z(n12456) );
  NANDN U5802 ( .A(y[1459]), .B(x[1459]), .Z(n7119) );
  ANDN U5803 ( .B(y[1458]), .A(x[1458]), .Z(n14955) );
  NANDN U5804 ( .A(x[1459]), .B(y[1459]), .Z(n22766) );
  AND U5805 ( .A(n7119), .B(n3147), .Z(n7123) );
  ANDN U5806 ( .B(y[1457]), .A(x[1457]), .Z(n14954) );
  NANDN U5807 ( .A(y[1453]), .B(x[1453]), .Z(n12460) );
  XNOR U5808 ( .A(x[1453]), .B(y[1453]), .Z(n7106) );
  NANDN U5809 ( .A(y[1451]), .B(x[1451]), .Z(n12464) );
  ANDN U5810 ( .B(x[1452]), .A(y[1452]), .Z(n12459) );
  ANDN U5811 ( .B(n12464), .A(n12459), .Z(n7103) );
  XNOR U5812 ( .A(x[1451]), .B(y[1451]), .Z(n7101) );
  NANDN U5813 ( .A(x[1450]), .B(y[1450]), .Z(n22746) );
  ANDN U5814 ( .B(x[1450]), .A(y[1450]), .Z(n12463) );
  NANDN U5815 ( .A(x[1448]), .B(y[1448]), .Z(n14940) );
  NANDN U5816 ( .A(x[1449]), .B(y[1449]), .Z(n14944) );
  NAND U5817 ( .A(n14940), .B(n14944), .Z(n22742) );
  NANDN U5818 ( .A(y[1448]), .B(x[1448]), .Z(n22741) );
  NANDN U5819 ( .A(y[1446]), .B(x[1446]), .Z(n3149) );
  NANDN U5820 ( .A(y[1447]), .B(x[1447]), .Z(n3148) );
  NAND U5821 ( .A(n3149), .B(n3148), .Z(n22737) );
  NANDN U5822 ( .A(y[1445]), .B(x[1445]), .Z(n3151) );
  NANDN U5823 ( .A(y[1444]), .B(x[1444]), .Z(n3150) );
  NAND U5824 ( .A(n3151), .B(n3150), .Z(n22733) );
  NANDN U5825 ( .A(x[1442]), .B(y[1442]), .Z(n12467) );
  XNOR U5826 ( .A(y[1442]), .B(x[1442]), .Z(n7083) );
  NANDN U5827 ( .A(x[1440]), .B(y[1440]), .Z(n14929) );
  ANDN U5828 ( .B(y[1441]), .A(x[1441]), .Z(n12468) );
  ANDN U5829 ( .B(n14929), .A(n12468), .Z(n7080) );
  XNOR U5830 ( .A(y[1440]), .B(x[1440]), .Z(n7078) );
  XNOR U5831 ( .A(x[1439]), .B(y[1439]), .Z(n7075) );
  NANDN U5832 ( .A(x[1436]), .B(y[1436]), .Z(n14922) );
  NANDN U5833 ( .A(x[1437]), .B(y[1437]), .Z(n14926) );
  NAND U5834 ( .A(n14922), .B(n14926), .Z(n22715) );
  NANDN U5835 ( .A(x[1432]), .B(y[1432]), .Z(n3153) );
  NANDN U5836 ( .A(x[1431]), .B(y[1431]), .Z(n3152) );
  AND U5837 ( .A(n3153), .B(n3152), .Z(n22706) );
  NANDN U5838 ( .A(y[1429]), .B(x[1429]), .Z(n12475) );
  XNOR U5839 ( .A(x[1429]), .B(y[1429]), .Z(n7048) );
  XNOR U5840 ( .A(y[1428]), .B(x[1428]), .Z(n7045) );
  NANDN U5841 ( .A(y[1425]), .B(x[1425]), .Z(n22693) );
  ANDN U5842 ( .B(x[1426]), .A(y[1426]), .Z(n14912) );
  ANDN U5843 ( .B(n22693), .A(n14912), .Z(n7038) );
  ANDN U5844 ( .B(y[1423]), .A(x[1423]), .Z(n22687) );
  NANDN U5845 ( .A(y[1417]), .B(x[1417]), .Z(n14895) );
  XNOR U5846 ( .A(x[1417]), .B(y[1417]), .Z(n7016) );
  NANDN U5847 ( .A(y[1415]), .B(x[1415]), .Z(n12485) );
  ANDN U5848 ( .B(x[1416]), .A(y[1416]), .Z(n14896) );
  ANDN U5849 ( .B(n12485), .A(n14896), .Z(n7013) );
  XNOR U5850 ( .A(x[1415]), .B(y[1415]), .Z(n7011) );
  ANDN U5851 ( .B(x[1413]), .A(y[1413]), .Z(n14886) );
  IV U5852 ( .A(n14886), .Z(n14888) );
  ANDN U5853 ( .B(x[1414]), .A(y[1414]), .Z(n12486) );
  ANDN U5854 ( .B(n14888), .A(n12486), .Z(n7008) );
  NANDN U5855 ( .A(y[1407]), .B(x[1407]), .Z(n3155) );
  NANDN U5856 ( .A(y[1406]), .B(x[1406]), .Z(n3154) );
  NAND U5857 ( .A(n3155), .B(n3154), .Z(n22657) );
  NANDN U5858 ( .A(x[1404]), .B(y[1404]), .Z(n12490) );
  XNOR U5859 ( .A(y[1404]), .B(x[1404]), .Z(n6980) );
  NANDN U5860 ( .A(x[1402]), .B(y[1402]), .Z(n22646) );
  ANDN U5861 ( .B(y[1403]), .A(x[1403]), .Z(n12489) );
  ANDN U5862 ( .B(n22646), .A(n12489), .Z(n6977) );
  ANDN U5863 ( .B(x[1402]), .A(y[1402]), .Z(n12492) );
  NANDN U5864 ( .A(x[1400]), .B(y[1400]), .Z(n3156) );
  NANDN U5865 ( .A(x[1401]), .B(y[1401]), .Z(n14875) );
  NAND U5866 ( .A(n3156), .B(n14875), .Z(n22642) );
  IV U5867 ( .A(y[1400]), .Z(n14870) );
  NAND U5868 ( .A(n14870), .B(x[1400]), .Z(n3160) );
  ANDN U5869 ( .B(y[1399]), .A(x[1399]), .Z(n14867) );
  NANDN U5870 ( .A(y[1398]), .B(x[1398]), .Z(n3158) );
  NANDN U5871 ( .A(y[1399]), .B(x[1399]), .Z(n3157) );
  NAND U5872 ( .A(n3158), .B(n3157), .Z(n14865) );
  NANDN U5873 ( .A(n14867), .B(n14865), .Z(n3159) );
  NAND U5874 ( .A(n3160), .B(n3159), .Z(n22641) );
  NANDN U5875 ( .A(x[1394]), .B(y[1394]), .Z(n12495) );
  XNOR U5876 ( .A(y[1394]), .B(x[1394]), .Z(n6960) );
  NANDN U5877 ( .A(x[1392]), .B(y[1392]), .Z(n12499) );
  ANDN U5878 ( .B(y[1393]), .A(x[1393]), .Z(n12496) );
  ANDN U5879 ( .B(n12499), .A(n12496), .Z(n6957) );
  XNOR U5880 ( .A(y[1392]), .B(x[1392]), .Z(n6955) );
  NANDN U5881 ( .A(x[1390]), .B(y[1390]), .Z(n12501) );
  ANDN U5882 ( .B(y[1391]), .A(x[1391]), .Z(n12500) );
  ANDN U5883 ( .B(n12501), .A(n12500), .Z(n6952) );
  NANDN U5884 ( .A(y[1389]), .B(x[1389]), .Z(n6947) );
  NANDN U5885 ( .A(y[1388]), .B(x[1388]), .Z(n3161) );
  AND U5886 ( .A(n6947), .B(n3161), .Z(n3167) );
  NANDN U5887 ( .A(y[1386]), .B(x[1386]), .Z(n3162) );
  NANDN U5888 ( .A(x[1387]), .B(n3162), .Z(n3165) );
  XNOR U5889 ( .A(n3162), .B(x[1387]), .Z(n3163) );
  NAND U5890 ( .A(n3163), .B(y[1387]), .Z(n3164) );
  NAND U5891 ( .A(n3165), .B(n3164), .Z(n3166) );
  NAND U5892 ( .A(n3167), .B(n3166), .Z(n22621) );
  NANDN U5893 ( .A(x[1380]), .B(y[1380]), .Z(n12503) );
  XNOR U5894 ( .A(y[1380]), .B(x[1380]), .Z(n6923) );
  NANDN U5895 ( .A(x[1378]), .B(y[1378]), .Z(n12509) );
  ANDN U5896 ( .B(y[1379]), .A(x[1379]), .Z(n12504) );
  ANDN U5897 ( .B(n12509), .A(n12504), .Z(n6920) );
  XNOR U5898 ( .A(y[1378]), .B(x[1378]), .Z(n6918) );
  NANDN U5899 ( .A(x[1375]), .B(y[1375]), .Z(n6909) );
  XNOR U5900 ( .A(x[1375]), .B(y[1375]), .Z(n3169) );
  NANDN U5901 ( .A(y[1374]), .B(x[1374]), .Z(n3168) );
  NAND U5902 ( .A(n3169), .B(n3168), .Z(n3170) );
  NAND U5903 ( .A(n6909), .B(n3170), .Z(n3172) );
  NANDN U5904 ( .A(y[1376]), .B(x[1376]), .Z(n3171) );
  NAND U5905 ( .A(n3172), .B(n3171), .Z(n12511) );
  NANDN U5906 ( .A(x[1362]), .B(y[1362]), .Z(n3174) );
  NANDN U5907 ( .A(x[1361]), .B(y[1361]), .Z(n3173) );
  NAND U5908 ( .A(n3174), .B(n3173), .Z(n22575) );
  NANDN U5909 ( .A(y[1355]), .B(x[1355]), .Z(n12513) );
  XNOR U5910 ( .A(x[1355]), .B(y[1355]), .Z(n6858) );
  XNOR U5911 ( .A(y[1354]), .B(x[1354]), .Z(n6855) );
  ANDN U5912 ( .B(x[1353]), .A(y[1353]), .Z(n12519) );
  NANDN U5913 ( .A(y[1351]), .B(x[1351]), .Z(n3176) );
  ANDN U5914 ( .B(x[1352]), .A(y[1352]), .Z(n3175) );
  ANDN U5915 ( .B(n3176), .A(n3175), .Z(n3180) );
  XNOR U5916 ( .A(x[1351]), .B(y[1351]), .Z(n3178) );
  ANDN U5917 ( .B(x[1350]), .A(y[1350]), .Z(n3177) );
  NAND U5918 ( .A(n3178), .B(n3177), .Z(n3179) );
  NAND U5919 ( .A(n3180), .B(n3179), .Z(n12518) );
  NANDN U5920 ( .A(x[1350]), .B(y[1350]), .Z(n3182) );
  NANDN U5921 ( .A(x[1349]), .B(y[1349]), .Z(n3181) );
  AND U5922 ( .A(n3182), .B(n3181), .Z(n3184) );
  NANDN U5923 ( .A(x[1351]), .B(y[1351]), .Z(n3183) );
  NAND U5924 ( .A(n3184), .B(n3183), .Z(n12523) );
  NANDN U5925 ( .A(y[1345]), .B(x[1345]), .Z(n14800) );
  XNOR U5926 ( .A(x[1345]), .B(y[1345]), .Z(n6838) );
  NANDN U5927 ( .A(y[1343]), .B(x[1343]), .Z(n12528) );
  ANDN U5928 ( .B(x[1344]), .A(y[1344]), .Z(n14799) );
  ANDN U5929 ( .B(n12528), .A(n14799), .Z(n6835) );
  XNOR U5930 ( .A(x[1343]), .B(y[1343]), .Z(n6833) );
  NANDN U5931 ( .A(x[1342]), .B(y[1342]), .Z(n22538) );
  ANDN U5932 ( .B(x[1341]), .A(y[1341]), .Z(n22535) );
  NANDN U5933 ( .A(x[1341]), .B(y[1341]), .Z(n14793) );
  NANDN U5934 ( .A(x[1340]), .B(y[1340]), .Z(n3185) );
  NAND U5935 ( .A(n14793), .B(n3185), .Z(n22534) );
  IV U5936 ( .A(n22534), .Z(n12530) );
  ANDN U5937 ( .B(x[1340]), .A(y[1340]), .Z(n14792) );
  ANDN U5938 ( .B(x[1339]), .A(y[1339]), .Z(n6822) );
  NANDN U5939 ( .A(x[1339]), .B(y[1339]), .Z(n22530) );
  ANDN U5940 ( .B(y[1338]), .A(x[1338]), .Z(n14786) );
  ANDN U5941 ( .B(n22530), .A(n14786), .Z(n3186) );
  OR U5942 ( .A(n6822), .B(n3186), .Z(n6826) );
  ANDN U5943 ( .B(y[1337]), .A(x[1337]), .Z(n14787) );
  NANDN U5944 ( .A(y[1331]), .B(x[1331]), .Z(n12531) );
  XNOR U5945 ( .A(x[1331]), .B(y[1331]), .Z(n6803) );
  XNOR U5946 ( .A(y[1330]), .B(x[1330]), .Z(n6800) );
  ANDN U5947 ( .B(y[1329]), .A(x[1329]), .Z(n12534) );
  IV U5948 ( .A(y[1328]), .Z(n20288) );
  NANDN U5949 ( .A(y[1327]), .B(x[1327]), .Z(n6796) );
  ANDN U5950 ( .B(y[1327]), .A(x[1327]), .Z(n22504) );
  ANDN U5951 ( .B(y[1326]), .A(x[1326]), .Z(n14768) );
  ANDN U5952 ( .B(y[1325]), .A(x[1325]), .Z(n14767) );
  NANDN U5953 ( .A(y[1325]), .B(x[1325]), .Z(n3188) );
  NANDN U5954 ( .A(y[1324]), .B(x[1324]), .Z(n3187) );
  NAND U5955 ( .A(n3188), .B(n3187), .Z(n22499) );
  ANDN U5956 ( .B(x[1316]), .A(y[1316]), .Z(n22479) );
  NANDN U5957 ( .A(y[1315]), .B(x[1315]), .Z(n6789) );
  ANDN U5958 ( .B(y[1314]), .A(x[1314]), .Z(n12547) );
  NANDN U5959 ( .A(x[1315]), .B(y[1315]), .Z(n22476) );
  ANDN U5960 ( .B(y[1313]), .A(x[1313]), .Z(n12546) );
  NANDN U5961 ( .A(y[1311]), .B(x[1311]), .Z(n3190) );
  NANDN U5962 ( .A(y[1310]), .B(x[1310]), .Z(n3189) );
  AND U5963 ( .A(n3190), .B(n3189), .Z(n22466) );
  NANDN U5964 ( .A(x[1308]), .B(y[1308]), .Z(n14743) );
  XNOR U5965 ( .A(y[1308]), .B(x[1308]), .Z(n6780) );
  XNOR U5966 ( .A(x[1307]), .B(y[1307]), .Z(n6777) );
  ANDN U5967 ( .B(x[1305]), .A(y[1305]), .Z(n12553) );
  ANDN U5968 ( .B(y[1305]), .A(x[1305]), .Z(n12554) );
  NANDN U5969 ( .A(y[1304]), .B(x[1304]), .Z(n12552) );
  NANDN U5970 ( .A(x[1303]), .B(y[1303]), .Z(n12556) );
  NANDN U5971 ( .A(y[1303]), .B(x[1303]), .Z(n3192) );
  NANDN U5972 ( .A(y[1302]), .B(x[1302]), .Z(n3191) );
  AND U5973 ( .A(n3192), .B(n3191), .Z(n22450) );
  ANDN U5974 ( .B(y[1301]), .A(x[1301]), .Z(n14736) );
  NANDN U5975 ( .A(x[1298]), .B(y[1298]), .Z(n3194) );
  NANDN U5976 ( .A(x[1297]), .B(y[1297]), .Z(n3193) );
  AND U5977 ( .A(n3194), .B(n3193), .Z(n22440) );
  ANDN U5978 ( .B(x[1295]), .A(y[1295]), .Z(n12559) );
  ANDN U5979 ( .B(x[1294]), .A(y[1294]), .Z(n12558) );
  NANDN U5980 ( .A(y[1293]), .B(x[1293]), .Z(n22430) );
  NANDN U5981 ( .A(x[1291]), .B(y[1291]), .Z(n22424) );
  NANDN U5982 ( .A(y[1289]), .B(x[1289]), .Z(n3196) );
  NANDN U5983 ( .A(y[1288]), .B(x[1288]), .Z(n3195) );
  NAND U5984 ( .A(n3196), .B(n3195), .Z(n22419) );
  NANDN U5985 ( .A(y[1285]), .B(x[1285]), .Z(n12567) );
  XNOR U5986 ( .A(x[1285]), .B(y[1285]), .Z(n6726) );
  NANDN U5987 ( .A(y[1283]), .B(x[1283]), .Z(n12570) );
  ANDN U5988 ( .B(x[1284]), .A(y[1284]), .Z(n12566) );
  ANDN U5989 ( .B(n12570), .A(n12566), .Z(n6723) );
  XNOR U5990 ( .A(x[1283]), .B(y[1283]), .Z(n6721) );
  NANDN U5991 ( .A(x[1282]), .B(y[1282]), .Z(n22404) );
  ANDN U5992 ( .B(x[1282]), .A(y[1282]), .Z(n12571) );
  NANDN U5993 ( .A(y[1281]), .B(x[1281]), .Z(n12572) );
  ANDN U5994 ( .B(y[1281]), .A(x[1281]), .Z(n12574) );
  NANDN U5995 ( .A(x[1280]), .B(y[1280]), .Z(n3197) );
  NANDN U5996 ( .A(n12574), .B(n3197), .Z(n14706) );
  ANDN U5997 ( .B(x[1280]), .A(y[1280]), .Z(n12573) );
  NANDN U5998 ( .A(y[1279]), .B(x[1279]), .Z(n3199) );
  NANDN U5999 ( .A(y[1278]), .B(x[1278]), .Z(n3198) );
  NAND U6000 ( .A(n3199), .B(n3198), .Z(n22399) );
  ANDN U6001 ( .B(y[1277]), .A(x[1277]), .Z(n14702) );
  ANDN U6002 ( .B(x[1270]), .A(y[1270]), .Z(n12582) );
  ANDN U6003 ( .B(x[1267]), .A(y[1267]), .Z(n12584) );
  ANDN U6004 ( .B(y[1266]), .A(x[1266]), .Z(n14681) );
  NANDN U6005 ( .A(x[1267]), .B(y[1267]), .Z(n22372) );
  ANDN U6006 ( .B(x[1266]), .A(y[1266]), .Z(n12585) );
  ANDN U6007 ( .B(y[1265]), .A(x[1265]), .Z(n14680) );
  NANDN U6008 ( .A(y[1261]), .B(x[1261]), .Z(n12588) );
  XNOR U6009 ( .A(x[1261]), .B(y[1261]), .Z(n6666) );
  NANDN U6010 ( .A(y[1259]), .B(x[1259]), .Z(n12590) );
  ANDN U6011 ( .B(x[1260]), .A(y[1260]), .Z(n12589) );
  ANDN U6012 ( .B(n12590), .A(n12589), .Z(n6663) );
  XNOR U6013 ( .A(x[1259]), .B(y[1259]), .Z(n6661) );
  NANDN U6014 ( .A(y[1257]), .B(x[1257]), .Z(n22350) );
  ANDN U6015 ( .B(x[1258]), .A(y[1258]), .Z(n12591) );
  ANDN U6016 ( .B(n22350), .A(n12591), .Z(n6658) );
  NANDN U6017 ( .A(y[1255]), .B(x[1255]), .Z(n6650) );
  NANDN U6018 ( .A(x[1255]), .B(y[1255]), .Z(n22345) );
  NANDN U6019 ( .A(x[1254]), .B(y[1254]), .Z(n12592) );
  NAND U6020 ( .A(n22345), .B(n12592), .Z(n3200) );
  AND U6021 ( .A(n6650), .B(n3200), .Z(n6654) );
  ANDN U6022 ( .B(y[1253]), .A(x[1253]), .Z(n12593) );
  NANDN U6023 ( .A(y[1247]), .B(x[1247]), .Z(n12596) );
  XNOR U6024 ( .A(x[1247]), .B(y[1247]), .Z(n6631) );
  XNOR U6025 ( .A(y[1246]), .B(x[1246]), .Z(n6628) );
  ANDN U6026 ( .B(x[1245]), .A(y[1245]), .Z(n12601) );
  NANDN U6027 ( .A(x[1243]), .B(y[1243]), .Z(n6619) );
  XNOR U6028 ( .A(x[1243]), .B(y[1243]), .Z(n3202) );
  NANDN U6029 ( .A(y[1242]), .B(x[1242]), .Z(n3201) );
  NAND U6030 ( .A(n3202), .B(n3201), .Z(n3203) );
  NAND U6031 ( .A(n6619), .B(n3203), .Z(n3205) );
  NANDN U6032 ( .A(y[1244]), .B(x[1244]), .Z(n3204) );
  NAND U6033 ( .A(n3205), .B(n3204), .Z(n12602) );
  NANDN U6034 ( .A(y[1241]), .B(x[1241]), .Z(n3207) );
  NANDN U6035 ( .A(y[1240]), .B(x[1240]), .Z(n3206) );
  AND U6036 ( .A(n3207), .B(n3206), .Z(n22318) );
  NANDN U6037 ( .A(y[1237]), .B(x[1237]), .Z(n12605) );
  XNOR U6038 ( .A(x[1237]), .B(y[1237]), .Z(n6607) );
  NANDN U6039 ( .A(y[1235]), .B(x[1235]), .Z(n12607) );
  ANDN U6040 ( .B(x[1236]), .A(y[1236]), .Z(n12606) );
  ANDN U6041 ( .B(n12607), .A(n12606), .Z(n6604) );
  XNOR U6042 ( .A(x[1235]), .B(y[1235]), .Z(n6602) );
  NANDN U6043 ( .A(x[1234]), .B(y[1234]), .Z(n22304) );
  ANDN U6044 ( .B(x[1232]), .A(y[1232]), .Z(n14636) );
  NANDN U6045 ( .A(y[1230]), .B(x[1230]), .Z(n3208) );
  NANDN U6046 ( .A(y[1231]), .B(x[1231]), .Z(n6593) );
  AND U6047 ( .A(n3208), .B(n6593), .Z(n22294) );
  ANDN U6048 ( .B(y[1229]), .A(x[1229]), .Z(n12610) );
  NANDN U6049 ( .A(y[1229]), .B(x[1229]), .Z(n3210) );
  NANDN U6050 ( .A(y[1228]), .B(x[1228]), .Z(n3209) );
  NAND U6051 ( .A(n3210), .B(n3209), .Z(n22291) );
  ANDN U6052 ( .B(y[1224]), .A(x[1224]), .Z(n6583) );
  NANDN U6053 ( .A(y[1223]), .B(x[1223]), .Z(n14621) );
  NANDN U6054 ( .A(y[1225]), .B(x[1225]), .Z(n3212) );
  NANDN U6055 ( .A(y[1224]), .B(x[1224]), .Z(n3211) );
  NAND U6056 ( .A(n3212), .B(n3211), .Z(n14625) );
  ANDN U6057 ( .B(x[1221]), .A(y[1221]), .Z(n12615) );
  ANDN U6058 ( .B(y[1221]), .A(x[1221]), .Z(n12613) );
  NANDN U6059 ( .A(x[1220]), .B(y[1220]), .Z(n3213) );
  NANDN U6060 ( .A(n12613), .B(n3213), .Z(n14617) );
  ANDN U6061 ( .B(x[1220]), .A(y[1220]), .Z(n12612) );
  ANDN U6062 ( .B(y[1219]), .A(x[1219]), .Z(n14616) );
  ANDN U6063 ( .B(x[1211]), .A(y[1211]), .Z(n12617) );
  NANDN U6064 ( .A(x[1210]), .B(y[1210]), .Z(n22256) );
  ANDN U6065 ( .B(y[1209]), .A(x[1209]), .Z(n12618) );
  ANDN U6066 ( .B(y[1208]), .A(x[1208]), .Z(n14600) );
  NOR U6067 ( .A(n12618), .B(n14600), .Z(n22252) );
  ANDN U6068 ( .B(y[1206]), .A(x[1206]), .Z(n12619) );
  NANDN U6069 ( .A(x[1207]), .B(y[1207]), .Z(n22248) );
  NANDN U6070 ( .A(n12619), .B(n22248), .Z(n3214) );
  NANDN U6071 ( .A(y[1207]), .B(x[1207]), .Z(n3215) );
  NAND U6072 ( .A(n3214), .B(n3215), .Z(n6555) );
  NANDN U6073 ( .A(y[1206]), .B(x[1206]), .Z(n3216) );
  AND U6074 ( .A(n3216), .B(n3215), .Z(n22246) );
  ANDN U6075 ( .B(y[1205]), .A(x[1205]), .Z(n12620) );
  NANDN U6076 ( .A(y[1205]), .B(x[1205]), .Z(n3218) );
  NANDN U6077 ( .A(y[1204]), .B(x[1204]), .Z(n3217) );
  NAND U6078 ( .A(n3218), .B(n3217), .Z(n22243) );
  NANDN U6079 ( .A(y[1201]), .B(x[1201]), .Z(n3220) );
  NANDN U6080 ( .A(y[1200]), .B(x[1200]), .Z(n3219) );
  NAND U6081 ( .A(n3220), .B(n3219), .Z(n14591) );
  IV U6082 ( .A(n14591), .Z(n6538) );
  NANDN U6083 ( .A(x[1195]), .B(y[1195]), .Z(n22225) );
  NANDN U6084 ( .A(y[1189]), .B(x[1189]), .Z(n12623) );
  XNOR U6085 ( .A(y[1188]), .B(x[1188]), .Z(n6526) );
  ANDN U6086 ( .B(x[1187]), .A(y[1187]), .Z(n12626) );
  NANDN U6087 ( .A(y[1182]), .B(x[1182]), .Z(n3222) );
  NANDN U6088 ( .A(y[1183]), .B(x[1183]), .Z(n3221) );
  NAND U6089 ( .A(n3222), .B(n3221), .Z(n22195) );
  NANDN U6090 ( .A(x[1176]), .B(y[1176]), .Z(n14546) );
  XNOR U6091 ( .A(y[1176]), .B(x[1176]), .Z(n6498) );
  XNOR U6092 ( .A(x[1175]), .B(y[1175]), .Z(n6495) );
  ANDN U6093 ( .B(x[1174]), .A(y[1174]), .Z(n12631) );
  ANDN U6094 ( .B(y[1173]), .A(x[1173]), .Z(n12632) );
  NANDN U6095 ( .A(x[1172]), .B(y[1172]), .Z(n12634) );
  NANDN U6096 ( .A(n12632), .B(n12634), .Z(n3223) );
  ANDN U6097 ( .B(x[1173]), .A(y[1173]), .Z(n6485) );
  ANDN U6098 ( .B(n3223), .A(n6485), .Z(n22174) );
  NANDN U6099 ( .A(y[1169]), .B(x[1169]), .Z(n3225) );
  NANDN U6100 ( .A(y[1168]), .B(x[1168]), .Z(n3224) );
  NAND U6101 ( .A(n3225), .B(n3224), .Z(n22169) );
  NANDN U6102 ( .A(y[1167]), .B(x[1167]), .Z(n3227) );
  NANDN U6103 ( .A(y[1166]), .B(x[1166]), .Z(n3226) );
  NAND U6104 ( .A(n3227), .B(n3226), .Z(n22165) );
  ANDN U6105 ( .B(x[1161]), .A(y[1161]), .Z(n3231) );
  NANDN U6106 ( .A(x[1160]), .B(y[1160]), .Z(n3228) );
  NANDN U6107 ( .A(x[1161]), .B(y[1161]), .Z(n14523) );
  NAND U6108 ( .A(n3228), .B(n14523), .Z(n12636) );
  NANDN U6109 ( .A(n3231), .B(n12636), .Z(n3229) );
  NANDN U6110 ( .A(x[1162]), .B(y[1162]), .Z(n14527) );
  NAND U6111 ( .A(n3229), .B(n14527), .Z(n22155) );
  NANDN U6112 ( .A(y[1160]), .B(x[1160]), .Z(n3230) );
  NANDN U6113 ( .A(n3231), .B(n3230), .Z(n14522) );
  ANDN U6114 ( .B(y[1159]), .A(x[1159]), .Z(n12635) );
  NANDN U6115 ( .A(y[1158]), .B(x[1158]), .Z(n3233) );
  NANDN U6116 ( .A(y[1159]), .B(x[1159]), .Z(n3232) );
  NAND U6117 ( .A(n3233), .B(n3232), .Z(n14519) );
  NANDN U6118 ( .A(n12635), .B(n14519), .Z(n3234) );
  NANDN U6119 ( .A(n14522), .B(n3234), .Z(n22153) );
  NANDN U6120 ( .A(y[1157]), .B(x[1157]), .Z(n3236) );
  NANDN U6121 ( .A(y[1156]), .B(x[1156]), .Z(n3235) );
  NAND U6122 ( .A(n3236), .B(n3235), .Z(n22148) );
  NANDN U6123 ( .A(x[1152]), .B(y[1152]), .Z(n12637) );
  XNOR U6124 ( .A(y[1152]), .B(x[1152]), .Z(n6446) );
  NANDN U6125 ( .A(x[1150]), .B(y[1150]), .Z(n14503) );
  ANDN U6126 ( .B(y[1151]), .A(x[1151]), .Z(n12638) );
  ANDN U6127 ( .B(n14503), .A(n12638), .Z(n6443) );
  XNOR U6128 ( .A(y[1150]), .B(x[1150]), .Z(n6441) );
  NANDN U6129 ( .A(x[1148]), .B(y[1148]), .Z(n3238) );
  NANDN U6130 ( .A(x[1149]), .B(y[1149]), .Z(n3237) );
  NAND U6131 ( .A(n3238), .B(n3237), .Z(n14500) );
  NANDN U6132 ( .A(y[1147]), .B(x[1147]), .Z(n3240) );
  ANDN U6133 ( .B(x[1148]), .A(y[1148]), .Z(n3239) );
  ANDN U6134 ( .B(n3240), .A(n3239), .Z(n3244) );
  XNOR U6135 ( .A(x[1147]), .B(y[1147]), .Z(n3242) );
  ANDN U6136 ( .B(x[1146]), .A(y[1146]), .Z(n3241) );
  NAND U6137 ( .A(n3242), .B(n3241), .Z(n3243) );
  NAND U6138 ( .A(n3244), .B(n3243), .Z(n12639) );
  NANDN U6139 ( .A(x[1144]), .B(y[1144]), .Z(n3246) );
  NANDN U6140 ( .A(x[1143]), .B(y[1143]), .Z(n3245) );
  AND U6141 ( .A(n3246), .B(n3245), .Z(n22126) );
  ANDN U6142 ( .B(x[1139]), .A(y[1139]), .Z(n12641) );
  NANDN U6143 ( .A(x[1138]), .B(y[1138]), .Z(n22114) );
  ANDN U6144 ( .B(y[1137]), .A(x[1137]), .Z(n12642) );
  ANDN U6145 ( .B(y[1136]), .A(x[1136]), .Z(n12643) );
  NOR U6146 ( .A(n12642), .B(n12643), .Z(n22110) );
  NANDN U6147 ( .A(x[1135]), .B(y[1135]), .Z(n22106) );
  ANDN U6148 ( .B(y[1133]), .A(x[1133]), .Z(n14479) );
  NANDN U6149 ( .A(y[1133]), .B(x[1133]), .Z(n3248) );
  NANDN U6150 ( .A(y[1132]), .B(x[1132]), .Z(n3247) );
  NAND U6151 ( .A(n3248), .B(n3247), .Z(n22100) );
  NANDN U6152 ( .A(x[1128]), .B(y[1128]), .Z(n14471) );
  XNOR U6153 ( .A(y[1128]), .B(x[1128]), .Z(n6408) );
  XNOR U6154 ( .A(x[1127]), .B(y[1127]), .Z(n6405) );
  ANDN U6155 ( .B(x[1126]), .A(y[1126]), .Z(n12647) );
  ANDN U6156 ( .B(x[1123]), .A(y[1123]), .Z(n12651) );
  NANDN U6157 ( .A(y[1124]), .B(x[1124]), .Z(n22080) );
  NANDN U6158 ( .A(x[1123]), .B(y[1123]), .Z(n22078) );
  NANDN U6159 ( .A(y[1121]), .B(x[1121]), .Z(n3250) );
  NANDN U6160 ( .A(y[1120]), .B(x[1120]), .Z(n3249) );
  NAND U6161 ( .A(n3250), .B(n3249), .Z(n22072) );
  NANDN U6162 ( .A(x[1114]), .B(y[1114]), .Z(n3252) );
  NANDN U6163 ( .A(x[1113]), .B(y[1113]), .Z(n3251) );
  NAND U6164 ( .A(n3252), .B(n3251), .Z(n14454) );
  NANDN U6165 ( .A(y[1113]), .B(x[1113]), .Z(n3255) );
  ANDN U6166 ( .B(y[1112]), .A(x[1112]), .Z(n12655) );
  NAND U6167 ( .A(n3255), .B(n12655), .Z(n3253) );
  NANDN U6168 ( .A(n14454), .B(n3253), .Z(n22059) );
  NANDN U6169 ( .A(y[1112]), .B(x[1112]), .Z(n3254) );
  NAND U6170 ( .A(n3255), .B(n3254), .Z(n22057) );
  NANDN U6171 ( .A(x[1111]), .B(y[1111]), .Z(n22054) );
  NANDN U6172 ( .A(x[1110]), .B(y[1110]), .Z(n22050) );
  NAND U6173 ( .A(n22054), .B(n22050), .Z(n6369) );
  ANDN U6174 ( .B(x[1110]), .A(y[1110]), .Z(n12657) );
  NANDN U6175 ( .A(y[1107]), .B(x[1107]), .Z(n3257) );
  NANDN U6176 ( .A(y[1106]), .B(x[1106]), .Z(n3256) );
  AND U6177 ( .A(n3257), .B(n3256), .Z(n22042) );
  NANDN U6178 ( .A(y[1104]), .B(x[1104]), .Z(n3259) );
  NANDN U6179 ( .A(y[1105]), .B(x[1105]), .Z(n3258) );
  AND U6180 ( .A(n3259), .B(n3258), .Z(n12662) );
  NANDN U6181 ( .A(y[1103]), .B(x[1103]), .Z(n12658) );
  NANDN U6182 ( .A(x[1104]), .B(y[1104]), .Z(n6349) );
  NANDN U6183 ( .A(n12658), .B(n6349), .Z(n6354) );
  NANDN U6184 ( .A(y[1101]), .B(x[1101]), .Z(n22034) );
  ANDN U6185 ( .B(x[1102]), .A(y[1102]), .Z(n12659) );
  ANDN U6186 ( .B(n22034), .A(n12659), .Z(n6348) );
  NANDN U6187 ( .A(x[1099]), .B(y[1099]), .Z(n22028) );
  ANDN U6188 ( .B(y[1097]), .A(x[1097]), .Z(n14432) );
  NANDN U6189 ( .A(y[1097]), .B(x[1097]), .Z(n3261) );
  NANDN U6190 ( .A(y[1096]), .B(x[1096]), .Z(n3260) );
  AND U6191 ( .A(n3261), .B(n3260), .Z(n22022) );
  NANDN U6192 ( .A(y[1095]), .B(x[1095]), .Z(n3263) );
  NANDN U6193 ( .A(y[1094]), .B(x[1094]), .Z(n3262) );
  AND U6194 ( .A(n3263), .B(n3262), .Z(n22018) );
  ANDN U6195 ( .B(x[1089]), .A(y[1089]), .Z(n14415) );
  ANDN U6196 ( .B(y[1089]), .A(x[1089]), .Z(n14414) );
  NANDN U6197 ( .A(x[1088]), .B(y[1088]), .Z(n3264) );
  NANDN U6198 ( .A(n14414), .B(n3264), .Z(n12668) );
  ANDN U6199 ( .B(x[1088]), .A(y[1088]), .Z(n14413) );
  NANDN U6200 ( .A(x[1087]), .B(y[1087]), .Z(n12667) );
  ANDN U6201 ( .B(y[1085]), .A(x[1085]), .Z(n12670) );
  NANDN U6202 ( .A(x[1084]), .B(y[1084]), .Z(n3266) );
  NANDN U6203 ( .A(x[1083]), .B(y[1083]), .Z(n3265) );
  NAND U6204 ( .A(n3266), .B(n3265), .Z(n22000) );
  NANDN U6205 ( .A(y[1081]), .B(x[1081]), .Z(n12674) );
  XNOR U6206 ( .A(x[1081]), .B(y[1081]), .Z(n6299) );
  NANDN U6207 ( .A(y[1079]), .B(x[1079]), .Z(n14402) );
  ANDN U6208 ( .B(x[1080]), .A(y[1080]), .Z(n12673) );
  ANDN U6209 ( .B(n14402), .A(n12673), .Z(n6296) );
  XNOR U6210 ( .A(x[1079]), .B(y[1079]), .Z(n6294) );
  NANDN U6211 ( .A(x[1078]), .B(y[1078]), .Z(n21989) );
  NANDN U6212 ( .A(y[1075]), .B(x[1075]), .Z(n6284) );
  NANDN U6213 ( .A(y[1074]), .B(x[1074]), .Z(n3267) );
  NAND U6214 ( .A(n6284), .B(n3267), .Z(n21979) );
  ANDN U6215 ( .B(y[1073]), .A(x[1073]), .Z(n12679) );
  NANDN U6216 ( .A(x[1072]), .B(y[1072]), .Z(n3269) );
  NANDN U6217 ( .A(x[1071]), .B(y[1071]), .Z(n3268) );
  AND U6218 ( .A(n3269), .B(n3268), .Z(n21972) );
  NANDN U6219 ( .A(x[1070]), .B(y[1070]), .Z(n3271) );
  NANDN U6220 ( .A(x[1069]), .B(y[1069]), .Z(n3270) );
  AND U6221 ( .A(n3271), .B(n3270), .Z(n21968) );
  NANDN U6222 ( .A(x[1068]), .B(y[1068]), .Z(n3273) );
  NANDN U6223 ( .A(x[1067]), .B(y[1067]), .Z(n3272) );
  AND U6224 ( .A(n3273), .B(n3272), .Z(n21964) );
  NANDN U6225 ( .A(y[1065]), .B(x[1065]), .Z(n6262) );
  NANDN U6226 ( .A(y[1064]), .B(x[1064]), .Z(n3274) );
  AND U6227 ( .A(n6262), .B(n3274), .Z(n21959) );
  ANDN U6228 ( .B(x[1063]), .A(y[1063]), .Z(n12681) );
  ANDN U6229 ( .B(n21959), .A(n12681), .Z(n6261) );
  XNOR U6230 ( .A(x[1062]), .B(y[1062]), .Z(n6257) );
  ANDN U6231 ( .B(y[1061]), .A(x[1061]), .Z(n12683) );
  NANDN U6232 ( .A(y[1061]), .B(x[1061]), .Z(n3276) );
  NANDN U6233 ( .A(y[1060]), .B(x[1060]), .Z(n3275) );
  NAND U6234 ( .A(n3276), .B(n3275), .Z(n21951) );
  NANDN U6235 ( .A(y[1059]), .B(x[1059]), .Z(n3278) );
  NANDN U6236 ( .A(y[1058]), .B(x[1058]), .Z(n3277) );
  AND U6237 ( .A(n3278), .B(n3277), .Z(n21946) );
  NANDN U6238 ( .A(y[1056]), .B(x[1056]), .Z(n3280) );
  NANDN U6239 ( .A(y[1057]), .B(x[1057]), .Z(n3279) );
  AND U6240 ( .A(n3280), .B(n3279), .Z(n12688) );
  NANDN U6241 ( .A(y[1055]), .B(x[1055]), .Z(n12684) );
  NANDN U6242 ( .A(x[1056]), .B(y[1056]), .Z(n6240) );
  NANDN U6243 ( .A(n12684), .B(n6240), .Z(n6245) );
  NANDN U6244 ( .A(y[1053]), .B(x[1053]), .Z(n21938) );
  ANDN U6245 ( .B(x[1054]), .A(y[1054]), .Z(n12685) );
  ANDN U6246 ( .B(n21938), .A(n12685), .Z(n6239) );
  NANDN U6247 ( .A(x[1051]), .B(y[1051]), .Z(n21932) );
  ANDN U6248 ( .B(y[1049]), .A(x[1049]), .Z(n12696) );
  ANDN U6249 ( .B(y[1044]), .A(x[1044]), .Z(n6220) );
  NANDN U6250 ( .A(y[1043]), .B(x[1043]), .Z(n14353) );
  NANDN U6251 ( .A(y[1045]), .B(x[1045]), .Z(n3282) );
  NANDN U6252 ( .A(y[1044]), .B(x[1044]), .Z(n3281) );
  NAND U6253 ( .A(n3282), .B(n3281), .Z(n14357) );
  ANDN U6254 ( .B(x[1040]), .A(y[1040]), .Z(n21911) );
  NANDN U6255 ( .A(x[1039]), .B(y[1039]), .Z(n21908) );
  NANDN U6256 ( .A(y[1033]), .B(x[1033]), .Z(n12700) );
  XNOR U6257 ( .A(x[1033]), .B(y[1033]), .Z(n6205) );
  XNOR U6258 ( .A(y[1032]), .B(x[1032]), .Z(n6202) );
  ANDN U6259 ( .B(y[1029]), .A(x[1029]), .Z(n12704) );
  ANDN U6260 ( .B(y[1028]), .A(x[1028]), .Z(n14323) );
  NOR U6261 ( .A(n12704), .B(n14323), .Z(n21884) );
  NANDN U6262 ( .A(x[1027]), .B(y[1027]), .Z(n21880) );
  NANDN U6263 ( .A(y[1026]), .B(x[1026]), .Z(n12705) );
  XNOR U6264 ( .A(x[1026]), .B(y[1026]), .Z(n6188) );
  NANDN U6265 ( .A(x[1024]), .B(y[1024]), .Z(n21872) );
  NANDN U6266 ( .A(y[1021]), .B(x[1021]), .Z(n3283) );
  IV U6267 ( .A(y[1022]), .Z(n12709) );
  NAND U6268 ( .A(n12709), .B(x[1022]), .Z(n12708) );
  NAND U6269 ( .A(n3283), .B(n12708), .Z(n21867) );
  NANDN U6270 ( .A(x[1019]), .B(y[1019]), .Z(n3285) );
  NANDN U6271 ( .A(x[1018]), .B(y[1018]), .Z(n3284) );
  AND U6272 ( .A(n3285), .B(n3284), .Z(n21860) );
  NANDN U6273 ( .A(y[1017]), .B(x[1017]), .Z(n3287) );
  NANDN U6274 ( .A(y[1018]), .B(x[1018]), .Z(n3286) );
  NAND U6275 ( .A(n3287), .B(n3286), .Z(n14302) );
  NANDN U6276 ( .A(x[1012]), .B(y[1012]), .Z(n3289) );
  NANDN U6277 ( .A(x[1011]), .B(y[1011]), .Z(n3288) );
  AND U6278 ( .A(n3289), .B(n3288), .Z(n21844) );
  NANDN U6279 ( .A(x[1006]), .B(y[1006]), .Z(n3291) );
  NANDN U6280 ( .A(x[1007]), .B(y[1007]), .Z(n3290) );
  AND U6281 ( .A(n3291), .B(n3290), .Z(n21832) );
  NANDN U6282 ( .A(y[1003]), .B(x[1003]), .Z(n3292) );
  NANDN U6283 ( .A(y[1004]), .B(x[1004]), .Z(n20291) );
  NAND U6284 ( .A(n3292), .B(n20291), .Z(n6142) );
  NANDN U6285 ( .A(y[1002]), .B(x[1002]), .Z(n3293) );
  NANDN U6286 ( .A(n6142), .B(n3293), .Z(n21824) );
  NANDN U6287 ( .A(x[1000]), .B(y[1000]), .Z(n3295) );
  NANDN U6288 ( .A(x[999]), .B(y[999]), .Z(n3294) );
  AND U6289 ( .A(n3295), .B(n3294), .Z(n21816) );
  NANDN U6290 ( .A(x[994]), .B(y[994]), .Z(n3297) );
  NANDN U6291 ( .A(x[995]), .B(y[995]), .Z(n3296) );
  AND U6292 ( .A(n3297), .B(n3296), .Z(n21804) );
  NANDN U6293 ( .A(y[993]), .B(x[993]), .Z(n3299) );
  NANDN U6294 ( .A(y[994]), .B(x[994]), .Z(n3298) );
  NAND U6295 ( .A(n3299), .B(n3298), .Z(n12713) );
  ANDN U6296 ( .B(y[991]), .A(x[991]), .Z(n21801) );
  NANDN U6297 ( .A(x[990]), .B(y[990]), .Z(n21794) );
  NANDN U6298 ( .A(n21801), .B(n21794), .Z(n3300) );
  ANDN U6299 ( .B(x[991]), .A(y[991]), .Z(n6117) );
  ANDN U6300 ( .B(n3300), .A(n6117), .Z(n14269) );
  NANDN U6301 ( .A(y[989]), .B(x[989]), .Z(n3302) );
  NANDN U6302 ( .A(y[988]), .B(x[988]), .Z(n3301) );
  NAND U6303 ( .A(n3302), .B(n3301), .Z(n21791) );
  NANDN U6304 ( .A(y[985]), .B(x[985]), .Z(n3304) );
  NANDN U6305 ( .A(y[984]), .B(x[984]), .Z(n3303) );
  NAND U6306 ( .A(n3304), .B(n3303), .Z(n21782) );
  NANDN U6307 ( .A(y[980]), .B(x[980]), .Z(n3306) );
  NANDN U6308 ( .A(y[979]), .B(x[979]), .Z(n3305) );
  NAND U6309 ( .A(n3306), .B(n3305), .Z(n21770) );
  NANDN U6310 ( .A(y[975]), .B(x[975]), .Z(n3308) );
  NANDN U6311 ( .A(y[974]), .B(x[974]), .Z(n3307) );
  NAND U6312 ( .A(n3308), .B(n3307), .Z(n21758) );
  NANDN U6313 ( .A(y[973]), .B(x[973]), .Z(n3310) );
  NANDN U6314 ( .A(y[972]), .B(x[972]), .Z(n3309) );
  NAND U6315 ( .A(n3310), .B(n3309), .Z(n21755) );
  NANDN U6316 ( .A(y[971]), .B(x[971]), .Z(n21750) );
  NANDN U6317 ( .A(y[970]), .B(x[970]), .Z(n3312) );
  NANDN U6318 ( .A(y[969]), .B(x[969]), .Z(n3311) );
  NAND U6319 ( .A(n3312), .B(n3311), .Z(n21746) );
  NANDN U6320 ( .A(y[968]), .B(x[968]), .Z(n3314) );
  NANDN U6321 ( .A(y[967]), .B(x[967]), .Z(n3313) );
  NAND U6322 ( .A(n3314), .B(n3313), .Z(n21743) );
  NANDN U6323 ( .A(y[966]), .B(x[966]), .Z(n21738) );
  NANDN U6324 ( .A(y[964]), .B(x[964]), .Z(n3316) );
  NANDN U6325 ( .A(y[965]), .B(x[965]), .Z(n3315) );
  NAND U6326 ( .A(n3316), .B(n3315), .Z(n21734) );
  NANDN U6327 ( .A(y[963]), .B(x[963]), .Z(n3318) );
  NANDN U6328 ( .A(y[962]), .B(x[962]), .Z(n3317) );
  NAND U6329 ( .A(n3318), .B(n3317), .Z(n21731) );
  NANDN U6330 ( .A(x[960]), .B(y[960]), .Z(n3320) );
  NANDN U6331 ( .A(x[959]), .B(y[959]), .Z(n3319) );
  NAND U6332 ( .A(n3320), .B(n3319), .Z(n14231) );
  NANDN U6333 ( .A(x[958]), .B(y[958]), .Z(n14228) );
  NANDN U6334 ( .A(y[959]), .B(x[959]), .Z(n3323) );
  NANDN U6335 ( .A(n14228), .B(n3323), .Z(n3321) );
  NANDN U6336 ( .A(n14231), .B(n3321), .Z(n21725) );
  NANDN U6337 ( .A(y[958]), .B(x[958]), .Z(n3322) );
  NAND U6338 ( .A(n3323), .B(n3322), .Z(n21722) );
  NANDN U6339 ( .A(x[957]), .B(y[957]), .Z(n21720) );
  ANDN U6340 ( .B(y[956]), .A(x[956]), .Z(n21714) );
  ANDN U6341 ( .B(n21720), .A(n21714), .Z(n6047) );
  NANDN U6342 ( .A(x[954]), .B(y[954]), .Z(n21709) );
  NANDN U6343 ( .A(x[955]), .B(y[955]), .Z(n21715) );
  NAND U6344 ( .A(n21709), .B(n21715), .Z(n14223) );
  ANDN U6345 ( .B(y[953]), .A(x[953]), .Z(n21708) );
  NANDN U6346 ( .A(x[952]), .B(y[952]), .Z(n3325) );
  NANDN U6347 ( .A(x[951]), .B(y[951]), .Z(n3324) );
  AND U6348 ( .A(n3325), .B(n3324), .Z(n21704) );
  NANDN U6349 ( .A(x[946]), .B(y[946]), .Z(n3326) );
  ANDN U6350 ( .B(y[947]), .A(x[947]), .Z(n12716) );
  ANDN U6351 ( .B(n3326), .A(n12716), .Z(n21692) );
  NANDN U6352 ( .A(y[945]), .B(x[945]), .Z(n14204) );
  NANDN U6353 ( .A(y[946]), .B(x[946]), .Z(n3327) );
  NAND U6354 ( .A(n14204), .B(n3327), .Z(n21691) );
  ANDN U6355 ( .B(y[942]), .A(x[942]), .Z(n21680) );
  ANDN U6356 ( .B(y[943]), .A(x[943]), .Z(n20295) );
  NANDN U6357 ( .A(x[941]), .B(y[941]), .Z(n21681) );
  NANDN U6358 ( .A(x[940]), .B(y[940]), .Z(n3329) );
  NANDN U6359 ( .A(x[939]), .B(y[939]), .Z(n3328) );
  AND U6360 ( .A(n3329), .B(n3328), .Z(n21676) );
  NANDN U6361 ( .A(x[934]), .B(y[934]), .Z(n3331) );
  NANDN U6362 ( .A(x[935]), .B(y[935]), .Z(n3330) );
  AND U6363 ( .A(n3331), .B(n3330), .Z(n21664) );
  NANDN U6364 ( .A(x[933]), .B(y[933]), .Z(n21657) );
  NANDN U6365 ( .A(x[932]), .B(y[932]), .Z(n3332) );
  NAND U6366 ( .A(n21657), .B(n3332), .Z(n14185) );
  IV U6367 ( .A(y[931]), .Z(n21651) );
  NAND U6368 ( .A(n21651), .B(x[931]), .Z(n3334) );
  NANDN U6369 ( .A(y[932]), .B(x[932]), .Z(n3333) );
  NAND U6370 ( .A(n3334), .B(n3333), .Z(n14184) );
  NANDN U6371 ( .A(x[930]), .B(y[930]), .Z(n21645) );
  NANDN U6372 ( .A(x[931]), .B(y[931]), .Z(n3335) );
  NAND U6373 ( .A(n21645), .B(n3335), .Z(n14182) );
  NANDN U6374 ( .A(x[929]), .B(y[929]), .Z(n21647) );
  NANDN U6375 ( .A(x[924]), .B(y[924]), .Z(n21633) );
  NANDN U6376 ( .A(y[921]), .B(x[921]), .Z(n14162) );
  NANDN U6377 ( .A(y[922]), .B(x[922]), .Z(n3336) );
  NAND U6378 ( .A(n14162), .B(n3336), .Z(n21627) );
  NANDN U6379 ( .A(x[921]), .B(y[921]), .Z(n3338) );
  NANDN U6380 ( .A(x[920]), .B(y[920]), .Z(n3337) );
  NAND U6381 ( .A(n3338), .B(n3337), .Z(n21626) );
  NANDN U6382 ( .A(x[919]), .B(y[919]), .Z(n3340) );
  NANDN U6383 ( .A(x[918]), .B(y[918]), .Z(n3339) );
  AND U6384 ( .A(n3340), .B(n3339), .Z(n21621) );
  NANDN U6385 ( .A(x[914]), .B(y[914]), .Z(n3342) );
  NANDN U6386 ( .A(x[913]), .B(y[913]), .Z(n3341) );
  AND U6387 ( .A(n3342), .B(n3341), .Z(n21609) );
  IV U6388 ( .A(y[907]), .Z(n21587) );
  NAND U6389 ( .A(n21587), .B(x[907]), .Z(n3344) );
  NANDN U6390 ( .A(y[908]), .B(x[908]), .Z(n3343) );
  NAND U6391 ( .A(n3344), .B(n3343), .Z(n14143) );
  NANDN U6392 ( .A(x[906]), .B(y[906]), .Z(n21583) );
  NANDN U6393 ( .A(x[907]), .B(y[907]), .Z(n3345) );
  NAND U6394 ( .A(n21583), .B(n3345), .Z(n14141) );
  NANDN U6395 ( .A(x[904]), .B(y[904]), .Z(n3347) );
  NANDN U6396 ( .A(x[903]), .B(y[903]), .Z(n3346) );
  AND U6397 ( .A(n3347), .B(n3346), .Z(n21577) );
  NANDN U6398 ( .A(y[898]), .B(x[898]), .Z(n3349) );
  NANDN U6399 ( .A(y[897]), .B(x[897]), .Z(n3348) );
  NAND U6400 ( .A(n3349), .B(n3348), .Z(n21564) );
  NANDN U6401 ( .A(x[895]), .B(y[895]), .Z(n21557) );
  NANDN U6402 ( .A(x[894]), .B(y[894]), .Z(n21553) );
  NAND U6403 ( .A(n21557), .B(n21553), .Z(n14126) );
  NANDN U6404 ( .A(y[893]), .B(x[893]), .Z(n3351) );
  NANDN U6405 ( .A(y[892]), .B(x[892]), .Z(n3350) );
  NAND U6406 ( .A(n3351), .B(n3350), .Z(n21550) );
  NANDN U6407 ( .A(y[889]), .B(x[889]), .Z(n3353) );
  NANDN U6408 ( .A(y[888]), .B(x[888]), .Z(n3352) );
  NAND U6409 ( .A(n3353), .B(n3352), .Z(n21541) );
  NANDN U6410 ( .A(y[884]), .B(x[884]), .Z(n21530) );
  NANDN U6411 ( .A(y[879]), .B(x[879]), .Z(n3355) );
  NANDN U6412 ( .A(y[878]), .B(x[878]), .Z(n3354) );
  NAND U6413 ( .A(n3355), .B(n3354), .Z(n21514) );
  NANDN U6414 ( .A(y[877]), .B(x[877]), .Z(n3357) );
  NANDN U6415 ( .A(y[876]), .B(x[876]), .Z(n3356) );
  NAND U6416 ( .A(n3357), .B(n3356), .Z(n21510) );
  NANDN U6417 ( .A(y[875]), .B(x[875]), .Z(n21506) );
  NANDN U6418 ( .A(y[874]), .B(x[874]), .Z(n3359) );
  NANDN U6419 ( .A(y[873]), .B(x[873]), .Z(n3358) );
  NAND U6420 ( .A(n3359), .B(n3358), .Z(n21502) );
  NANDN U6421 ( .A(y[872]), .B(x[872]), .Z(n3361) );
  NANDN U6422 ( .A(y[871]), .B(x[871]), .Z(n3360) );
  NAND U6423 ( .A(n3361), .B(n3360), .Z(n21498) );
  NANDN U6424 ( .A(y[870]), .B(x[870]), .Z(n21494) );
  NANDN U6425 ( .A(y[868]), .B(x[868]), .Z(n3363) );
  NANDN U6426 ( .A(y[869]), .B(x[869]), .Z(n3362) );
  NAND U6427 ( .A(n3363), .B(n3362), .Z(n21490) );
  NANDN U6428 ( .A(y[867]), .B(x[867]), .Z(n3365) );
  NANDN U6429 ( .A(y[866]), .B(x[866]), .Z(n3364) );
  NAND U6430 ( .A(n3365), .B(n3364), .Z(n21486) );
  NANDN U6431 ( .A(x[866]), .B(y[866]), .Z(n3367) );
  NANDN U6432 ( .A(x[865]), .B(y[865]), .Z(n3366) );
  NAND U6433 ( .A(n3367), .B(n3366), .Z(n21484) );
  NANDN U6434 ( .A(y[865]), .B(x[865]), .Z(n3369) );
  NANDN U6435 ( .A(y[864]), .B(x[864]), .Z(n3368) );
  NAND U6436 ( .A(n3369), .B(n3368), .Z(n21482) );
  NANDN U6437 ( .A(x[862]), .B(y[862]), .Z(n14081) );
  NANDN U6438 ( .A(y[863]), .B(x[863]), .Z(n3374) );
  NANDN U6439 ( .A(n14081), .B(n3374), .Z(n3372) );
  NANDN U6440 ( .A(x[864]), .B(y[864]), .Z(n3371) );
  NANDN U6441 ( .A(x[863]), .B(y[863]), .Z(n3370) );
  AND U6442 ( .A(n3371), .B(n3370), .Z(n14084) );
  NAND U6443 ( .A(n3372), .B(n14084), .Z(n21480) );
  NANDN U6444 ( .A(y[862]), .B(x[862]), .Z(n3373) );
  NAND U6445 ( .A(n3374), .B(n3373), .Z(n21478) );
  ANDN U6446 ( .B(x[861]), .A(y[861]), .Z(n12719) );
  ANDN U6447 ( .B(x[860]), .A(y[860]), .Z(n12720) );
  ANDN U6448 ( .B(x[859]), .A(y[859]), .Z(n5847) );
  NANDN U6449 ( .A(y[858]), .B(x[858]), .Z(n3375) );
  NANDN U6450 ( .A(n5847), .B(n3375), .Z(n21467) );
  NANDN U6451 ( .A(x[854]), .B(y[854]), .Z(n3377) );
  NANDN U6452 ( .A(x[853]), .B(y[853]), .Z(n3376) );
  AND U6453 ( .A(n3377), .B(n3376), .Z(n21455) );
  NANDN U6454 ( .A(y[851]), .B(x[851]), .Z(n21450) );
  NANDN U6455 ( .A(x[850]), .B(y[850]), .Z(n3378) );
  NANDN U6456 ( .A(x[851]), .B(y[851]), .Z(n14067) );
  NAND U6457 ( .A(n3378), .B(n14067), .Z(n21448) );
  NANDN U6458 ( .A(y[850]), .B(x[850]), .Z(n3382) );
  ANDN U6459 ( .B(y[849]), .A(x[849]), .Z(n14059) );
  IV U6460 ( .A(n14059), .Z(n5826) );
  NANDN U6461 ( .A(y[849]), .B(x[849]), .Z(n3380) );
  NANDN U6462 ( .A(y[848]), .B(x[848]), .Z(n3379) );
  NAND U6463 ( .A(n3380), .B(n3379), .Z(n14058) );
  NAND U6464 ( .A(n5826), .B(n14058), .Z(n3381) );
  NAND U6465 ( .A(n3382), .B(n3381), .Z(n21446) );
  NANDN U6466 ( .A(y[847]), .B(x[847]), .Z(n3384) );
  NANDN U6467 ( .A(y[846]), .B(x[846]), .Z(n3383) );
  NAND U6468 ( .A(n3384), .B(n3383), .Z(n21442) );
  NANDN U6469 ( .A(y[843]), .B(x[843]), .Z(n3386) );
  NANDN U6470 ( .A(y[842]), .B(x[842]), .Z(n3385) );
  NAND U6471 ( .A(n3386), .B(n3385), .Z(n21434) );
  NANDN U6472 ( .A(x[840]), .B(y[840]), .Z(n14044) );
  NANDN U6473 ( .A(y[841]), .B(x[841]), .Z(n3391) );
  NANDN U6474 ( .A(n14044), .B(n3391), .Z(n3389) );
  NANDN U6475 ( .A(x[842]), .B(y[842]), .Z(n3388) );
  NANDN U6476 ( .A(x[841]), .B(y[841]), .Z(n3387) );
  AND U6477 ( .A(n3388), .B(n3387), .Z(n14048) );
  NAND U6478 ( .A(n3389), .B(n14048), .Z(n21432) );
  NANDN U6479 ( .A(y[840]), .B(x[840]), .Z(n3390) );
  NAND U6480 ( .A(n3391), .B(n3390), .Z(n21430) );
  NANDN U6481 ( .A(y[837]), .B(x[837]), .Z(n3393) );
  NANDN U6482 ( .A(y[836]), .B(x[836]), .Z(n3392) );
  NAND U6483 ( .A(n3393), .B(n3392), .Z(n21422) );
  NANDN U6484 ( .A(y[835]), .B(x[835]), .Z(n3395) );
  NANDN U6485 ( .A(y[834]), .B(x[834]), .Z(n3394) );
  NAND U6486 ( .A(n3395), .B(n3394), .Z(n21418) );
  NANDN U6487 ( .A(y[831]), .B(x[831]), .Z(n3397) );
  NANDN U6488 ( .A(y[830]), .B(x[830]), .Z(n3396) );
  NAND U6489 ( .A(n3397), .B(n3396), .Z(n21410) );
  NANDN U6490 ( .A(y[829]), .B(x[829]), .Z(n3399) );
  NANDN U6491 ( .A(y[828]), .B(x[828]), .Z(n3398) );
  NAND U6492 ( .A(n3399), .B(n3398), .Z(n21406) );
  NANDN U6493 ( .A(x[826]), .B(y[826]), .Z(n3401) );
  NANDN U6494 ( .A(x[825]), .B(y[825]), .Z(n3400) );
  AND U6495 ( .A(n3401), .B(n3400), .Z(n3402) );
  NANDN U6496 ( .A(x[827]), .B(y[827]), .Z(n5782) );
  NAND U6497 ( .A(n3402), .B(n5782), .Z(n12724) );
  NANDN U6498 ( .A(y[822]), .B(x[822]), .Z(n3404) );
  NANDN U6499 ( .A(y[823]), .B(x[823]), .Z(n3403) );
  NAND U6500 ( .A(n3404), .B(n3403), .Z(n21394) );
  NANDN U6501 ( .A(y[821]), .B(x[821]), .Z(n3406) );
  NANDN U6502 ( .A(y[820]), .B(x[820]), .Z(n3405) );
  NAND U6503 ( .A(n3406), .B(n3405), .Z(n21389) );
  NANDN U6504 ( .A(y[817]), .B(x[817]), .Z(n3408) );
  NANDN U6505 ( .A(y[816]), .B(x[816]), .Z(n3407) );
  NAND U6506 ( .A(n3408), .B(n3407), .Z(n21382) );
  NANDN U6507 ( .A(y[815]), .B(x[815]), .Z(n3414) );
  ANDN U6508 ( .B(x[813]), .A(y[813]), .Z(n3409) );
  OR U6509 ( .A(n3409), .B(x[814]), .Z(n3412) );
  XOR U6510 ( .A(x[814]), .B(n3409), .Z(n3410) );
  NAND U6511 ( .A(n3410), .B(y[814]), .Z(n3411) );
  NAND U6512 ( .A(n3412), .B(n3411), .Z(n3413) );
  NAND U6513 ( .A(n3414), .B(n3413), .Z(n21377) );
  NANDN U6514 ( .A(y[809]), .B(x[809]), .Z(n3416) );
  NANDN U6515 ( .A(y[808]), .B(x[808]), .Z(n3415) );
  NAND U6516 ( .A(n3416), .B(n3415), .Z(n21370) );
  NANDN U6517 ( .A(x[805]), .B(y[805]), .Z(n3418) );
  NANDN U6518 ( .A(x[806]), .B(y[806]), .Z(n3417) );
  NAND U6519 ( .A(n3418), .B(n3417), .Z(n12728) );
  ANDN U6520 ( .B(y[804]), .A(x[804]), .Z(n12725) );
  ANDN U6521 ( .B(x[803]), .A(y[803]), .Z(n12729) );
  NANDN U6522 ( .A(y[799]), .B(x[799]), .Z(n3420) );
  NANDN U6523 ( .A(y[798]), .B(x[798]), .Z(n3419) );
  AND U6524 ( .A(n3420), .B(n3419), .Z(n21353) );
  NANDN U6525 ( .A(y[793]), .B(x[793]), .Z(n3422) );
  NANDN U6526 ( .A(y[792]), .B(x[792]), .Z(n3421) );
  AND U6527 ( .A(n3422), .B(n3421), .Z(n21341) );
  NANDN U6528 ( .A(y[787]), .B(x[787]), .Z(n3424) );
  NANDN U6529 ( .A(y[786]), .B(x[786]), .Z(n3423) );
  AND U6530 ( .A(n3424), .B(n3423), .Z(n21329) );
  NANDN U6531 ( .A(y[781]), .B(x[781]), .Z(n3426) );
  NANDN U6532 ( .A(y[780]), .B(x[780]), .Z(n3425) );
  AND U6533 ( .A(n3426), .B(n3425), .Z(n21317) );
  ANDN U6534 ( .B(y[776]), .A(x[776]), .Z(n13983) );
  ANDN U6535 ( .B(y[775]), .A(x[775]), .Z(n13978) );
  NANDN U6536 ( .A(y[775]), .B(x[775]), .Z(n13980) );
  NANDN U6537 ( .A(y[774]), .B(x[774]), .Z(n3427) );
  NAND U6538 ( .A(n13980), .B(n3427), .Z(n21305) );
  NANDN U6539 ( .A(x[770]), .B(y[770]), .Z(n3429) );
  NANDN U6540 ( .A(x[769]), .B(y[769]), .Z(n3428) );
  AND U6541 ( .A(n3429), .B(n3428), .Z(n21295) );
  NANDN U6542 ( .A(y[767]), .B(x[767]), .Z(n12732) );
  NANDN U6543 ( .A(y[766]), .B(x[766]), .Z(n12731) );
  NAND U6544 ( .A(n12732), .B(n12731), .Z(n21289) );
  NANDN U6545 ( .A(x[764]), .B(y[764]), .Z(n3431) );
  NANDN U6546 ( .A(x[763]), .B(y[763]), .Z(n3430) );
  AND U6547 ( .A(n3431), .B(n3430), .Z(n21283) );
  NANDN U6548 ( .A(x[762]), .B(y[762]), .Z(n3433) );
  NANDN U6549 ( .A(x[761]), .B(y[761]), .Z(n3432) );
  AND U6550 ( .A(n3433), .B(n3432), .Z(n21279) );
  NANDN U6551 ( .A(x[756]), .B(y[756]), .Z(n3435) );
  NANDN U6552 ( .A(x[755]), .B(y[755]), .Z(n3434) );
  AND U6553 ( .A(n3435), .B(n3434), .Z(n21267) );
  NANDN U6554 ( .A(x[754]), .B(y[754]), .Z(n21263) );
  NANDN U6555 ( .A(x[753]), .B(y[753]), .Z(n3436) );
  NAND U6556 ( .A(n21263), .B(n3436), .Z(n5595) );
  NANDN U6557 ( .A(x[752]), .B(y[752]), .Z(n3437) );
  NANDN U6558 ( .A(n5595), .B(n3437), .Z(n21260) );
  ANDN U6559 ( .B(y[751]), .A(x[751]), .Z(n5590) );
  NANDN U6560 ( .A(y[750]), .B(x[750]), .Z(n13945) );
  ANDN U6561 ( .B(x[751]), .A(y[751]), .Z(n13948) );
  ANDN U6562 ( .B(n13945), .A(n13948), .Z(n3438) );
  NOR U6563 ( .A(n5590), .B(n3438), .Z(n21255) );
  NANDN U6564 ( .A(x[748]), .B(y[748]), .Z(n3440) );
  NANDN U6565 ( .A(x[747]), .B(y[747]), .Z(n3439) );
  AND U6566 ( .A(n3440), .B(n3439), .Z(n21249) );
  NANDN U6567 ( .A(x[742]), .B(y[742]), .Z(n3442) );
  NANDN U6568 ( .A(x[741]), .B(y[741]), .Z(n3441) );
  AND U6569 ( .A(n3442), .B(n3441), .Z(n3444) );
  NANDN U6570 ( .A(x[743]), .B(y[743]), .Z(n3443) );
  AND U6571 ( .A(n3444), .B(n3443), .Z(n21237) );
  NANDN U6572 ( .A(y[739]), .B(x[739]), .Z(n3446) );
  NANDN U6573 ( .A(y[738]), .B(x[738]), .Z(n3445) );
  AND U6574 ( .A(n3446), .B(n3445), .Z(n3452) );
  NANDN U6575 ( .A(y[736]), .B(x[736]), .Z(n3447) );
  NANDN U6576 ( .A(x[737]), .B(n3447), .Z(n3450) );
  XNOR U6577 ( .A(n3447), .B(x[737]), .Z(n3448) );
  NAND U6578 ( .A(n3448), .B(y[737]), .Z(n3449) );
  NAND U6579 ( .A(n3450), .B(n3449), .Z(n3451) );
  NAND U6580 ( .A(n3452), .B(n3451), .Z(n21232) );
  NANDN U6581 ( .A(y[735]), .B(x[735]), .Z(n3454) );
  NANDN U6582 ( .A(y[734]), .B(x[734]), .Z(n3453) );
  NAND U6583 ( .A(n3454), .B(n3453), .Z(n21228) );
  ANDN U6584 ( .B(y[733]), .A(x[733]), .Z(n12734) );
  NANDN U6585 ( .A(y[730]), .B(x[730]), .Z(n3456) );
  NANDN U6586 ( .A(y[731]), .B(x[731]), .Z(n3455) );
  NAND U6587 ( .A(n3456), .B(n3455), .Z(n21220) );
  NANDN U6588 ( .A(y[729]), .B(x[729]), .Z(n3458) );
  NANDN U6589 ( .A(y[728]), .B(x[728]), .Z(n3457) );
  NAND U6590 ( .A(n3458), .B(n3457), .Z(n21216) );
  NANDN U6591 ( .A(y[725]), .B(x[725]), .Z(n3460) );
  NANDN U6592 ( .A(y[724]), .B(x[724]), .Z(n3459) );
  NAND U6593 ( .A(n3460), .B(n3459), .Z(n21208) );
  NANDN U6594 ( .A(y[723]), .B(x[723]), .Z(n3462) );
  NANDN U6595 ( .A(y[722]), .B(x[722]), .Z(n3461) );
  NAND U6596 ( .A(n3462), .B(n3461), .Z(n21204) );
  NANDN U6597 ( .A(x[719]), .B(y[719]), .Z(n5517) );
  XNOR U6598 ( .A(x[719]), .B(y[719]), .Z(n3464) );
  NANDN U6599 ( .A(y[718]), .B(x[718]), .Z(n3463) );
  NAND U6600 ( .A(n3464), .B(n3463), .Z(n3465) );
  AND U6601 ( .A(n5517), .B(n3465), .Z(n21196) );
  NANDN U6602 ( .A(y[717]), .B(x[717]), .Z(n3467) );
  NANDN U6603 ( .A(y[716]), .B(x[716]), .Z(n3466) );
  NAND U6604 ( .A(n3467), .B(n3466), .Z(n21192) );
  NANDN U6605 ( .A(x[713]), .B(y[713]), .Z(n3469) );
  NANDN U6606 ( .A(x[714]), .B(y[714]), .Z(n3468) );
  NAND U6607 ( .A(n3469), .B(n3468), .Z(n13907) );
  NANDN U6608 ( .A(y[710]), .B(x[710]), .Z(n3471) );
  NANDN U6609 ( .A(y[711]), .B(x[711]), .Z(n3470) );
  NAND U6610 ( .A(n3471), .B(n3470), .Z(n21180) );
  NANDN U6611 ( .A(y[709]), .B(x[709]), .Z(n3473) );
  NANDN U6612 ( .A(y[708]), .B(x[708]), .Z(n3472) );
  NAND U6613 ( .A(n3473), .B(n3472), .Z(n21175) );
  NANDN U6614 ( .A(x[705]), .B(y[705]), .Z(n5487) );
  XNOR U6615 ( .A(x[705]), .B(y[705]), .Z(n3475) );
  NANDN U6616 ( .A(y[704]), .B(x[704]), .Z(n3474) );
  NAND U6617 ( .A(n3475), .B(n3474), .Z(n3476) );
  AND U6618 ( .A(n5487), .B(n3476), .Z(n21168) );
  NANDN U6619 ( .A(y[703]), .B(x[703]), .Z(n3478) );
  NANDN U6620 ( .A(y[702]), .B(x[702]), .Z(n3477) );
  NAND U6621 ( .A(n3478), .B(n3477), .Z(n21163) );
  NANDN U6622 ( .A(y[699]), .B(x[699]), .Z(n3480) );
  NANDN U6623 ( .A(y[698]), .B(x[698]), .Z(n3479) );
  NAND U6624 ( .A(n3480), .B(n3479), .Z(n21156) );
  NANDN U6625 ( .A(x[697]), .B(y[697]), .Z(n3482) );
  NANDN U6626 ( .A(x[698]), .B(y[698]), .Z(n3481) );
  NAND U6627 ( .A(n3482), .B(n3481), .Z(n12742) );
  ANDN U6628 ( .B(y[696]), .A(x[696]), .Z(n12739) );
  NANDN U6629 ( .A(y[692]), .B(x[692]), .Z(n3484) );
  NANDN U6630 ( .A(y[693]), .B(x[693]), .Z(n3483) );
  AND U6631 ( .A(n3484), .B(n3483), .Z(n21143) );
  NANDN U6632 ( .A(x[685]), .B(y[685]), .Z(n5442) );
  XNOR U6633 ( .A(x[685]), .B(y[685]), .Z(n3486) );
  NANDN U6634 ( .A(y[684]), .B(x[684]), .Z(n3485) );
  NAND U6635 ( .A(n3486), .B(n3485), .Z(n3487) );
  NAND U6636 ( .A(n5442), .B(n3487), .Z(n3489) );
  NANDN U6637 ( .A(y[686]), .B(x[686]), .Z(n3488) );
  AND U6638 ( .A(n3489), .B(n3488), .Z(n3491) );
  NANDN U6639 ( .A(y[687]), .B(x[687]), .Z(n3490) );
  AND U6640 ( .A(n3491), .B(n3490), .Z(n21131) );
  NANDN U6641 ( .A(y[679]), .B(x[679]), .Z(n3493) );
  NANDN U6642 ( .A(y[678]), .B(x[678]), .Z(n3492) );
  AND U6643 ( .A(n3493), .B(n3492), .Z(n21119) );
  NANDN U6644 ( .A(y[677]), .B(x[677]), .Z(n21112) );
  NANDN U6645 ( .A(y[676]), .B(x[676]), .Z(n3494) );
  NAND U6646 ( .A(n21112), .B(n3494), .Z(n13868) );
  IV U6647 ( .A(x[675]), .Z(n21106) );
  NAND U6648 ( .A(n21106), .B(y[675]), .Z(n3496) );
  NANDN U6649 ( .A(x[676]), .B(y[676]), .Z(n3495) );
  NAND U6650 ( .A(n3496), .B(n3495), .Z(n13866) );
  ANDN U6651 ( .B(x[674]), .A(y[674]), .Z(n21100) );
  NANDN U6652 ( .A(y[675]), .B(x[675]), .Z(n3497) );
  NANDN U6653 ( .A(n21100), .B(n3497), .Z(n13864) );
  NANDN U6654 ( .A(y[673]), .B(x[673]), .Z(n21101) );
  NANDN U6655 ( .A(x[672]), .B(y[672]), .Z(n13855) );
  NANDN U6656 ( .A(x[673]), .B(y[673]), .Z(n13861) );
  NAND U6657 ( .A(n13855), .B(n13861), .Z(n21098) );
  NANDN U6658 ( .A(y[670]), .B(x[670]), .Z(n3499) );
  NANDN U6659 ( .A(y[671]), .B(x[671]), .Z(n3498) );
  NAND U6660 ( .A(n3499), .B(n3498), .Z(n21092) );
  NANDN U6661 ( .A(y[665]), .B(x[665]), .Z(n3501) );
  NANDN U6662 ( .A(y[664]), .B(x[664]), .Z(n3500) );
  NAND U6663 ( .A(n3501), .B(n3500), .Z(n21080) );
  NANDN U6664 ( .A(x[663]), .B(y[663]), .Z(n3503) );
  NANDN U6665 ( .A(x[664]), .B(y[664]), .Z(n3502) );
  NAND U6666 ( .A(n3503), .B(n3502), .Z(n13846) );
  ANDN U6667 ( .B(y[662]), .A(x[662]), .Z(n13843) );
  NANDN U6668 ( .A(y[660]), .B(x[660]), .Z(n3505) );
  NANDN U6669 ( .A(y[661]), .B(x[661]), .Z(n3504) );
  NAND U6670 ( .A(n3505), .B(n3504), .Z(n21073) );
  NANDN U6671 ( .A(y[657]), .B(x[657]), .Z(n3507) );
  NANDN U6672 ( .A(y[656]), .B(x[656]), .Z(n3506) );
  NAND U6673 ( .A(n3507), .B(n3506), .Z(n21065) );
  NANDN U6674 ( .A(y[655]), .B(x[655]), .Z(n3509) );
  NANDN U6675 ( .A(y[654]), .B(x[654]), .Z(n3508) );
  NAND U6676 ( .A(n3509), .B(n3508), .Z(n21061) );
  NANDN U6677 ( .A(x[651]), .B(y[651]), .Z(n5368) );
  XNOR U6678 ( .A(x[651]), .B(y[651]), .Z(n3511) );
  NANDN U6679 ( .A(y[650]), .B(x[650]), .Z(n3510) );
  NAND U6680 ( .A(n3511), .B(n3510), .Z(n3512) );
  AND U6681 ( .A(n5368), .B(n3512), .Z(n21053) );
  NANDN U6682 ( .A(y[649]), .B(x[649]), .Z(n3514) );
  NANDN U6683 ( .A(y[648]), .B(x[648]), .Z(n3513) );
  NAND U6684 ( .A(n3514), .B(n3513), .Z(n21049) );
  NANDN U6685 ( .A(x[647]), .B(y[647]), .Z(n3516) );
  NANDN U6686 ( .A(x[648]), .B(y[648]), .Z(n3515) );
  NAND U6687 ( .A(n3516), .B(n3515), .Z(n12746) );
  NANDN U6688 ( .A(y[646]), .B(x[646]), .Z(n3517) );
  ANDN U6689 ( .B(x[647]), .A(y[647]), .Z(n12744) );
  ANDN U6690 ( .B(n3517), .A(n12744), .Z(n21044) );
  ANDN U6691 ( .B(y[646]), .A(x[646]), .Z(n12743) );
  NANDN U6692 ( .A(x[642]), .B(y[642]), .Z(n3519) );
  NANDN U6693 ( .A(x[641]), .B(y[641]), .Z(n3518) );
  NAND U6694 ( .A(n3519), .B(n3518), .Z(n21034) );
  NANDN U6695 ( .A(x[640]), .B(y[640]), .Z(n3521) );
  NANDN U6696 ( .A(x[639]), .B(y[639]), .Z(n3520) );
  NAND U6697 ( .A(n3521), .B(n3520), .Z(n21031) );
  NANDN U6698 ( .A(y[635]), .B(x[635]), .Z(n21020) );
  NANDN U6699 ( .A(y[634]), .B(x[634]), .Z(n21015) );
  NANDN U6700 ( .A(x[635]), .B(y[635]), .Z(n3524) );
  NANDN U6701 ( .A(n21015), .B(n3524), .Z(n3522) );
  NAND U6702 ( .A(n21020), .B(n3522), .Z(n13810) );
  NANDN U6703 ( .A(x[634]), .B(y[634]), .Z(n3523) );
  NAND U6704 ( .A(n3524), .B(n3523), .Z(n21019) );
  NANDN U6705 ( .A(y[633]), .B(x[633]), .Z(n13806) );
  IV U6706 ( .A(y[632]), .Z(n13801) );
  NAND U6707 ( .A(n13801), .B(x[632]), .Z(n3525) );
  AND U6708 ( .A(n13806), .B(n3525), .Z(n3526) );
  ANDN U6709 ( .B(y[633]), .A(x[633]), .Z(n5334) );
  NOR U6710 ( .A(n3526), .B(n5334), .Z(n21017) );
  NANDN U6711 ( .A(x[630]), .B(y[630]), .Z(n3528) );
  NANDN U6712 ( .A(x[629]), .B(y[629]), .Z(n3527) );
  NAND U6713 ( .A(n3528), .B(n3527), .Z(n21009) );
  NANDN U6714 ( .A(x[628]), .B(y[628]), .Z(n3530) );
  NANDN U6715 ( .A(x[627]), .B(y[627]), .Z(n3529) );
  NAND U6716 ( .A(n3530), .B(n3529), .Z(n21004) );
  NANDN U6717 ( .A(x[626]), .B(y[626]), .Z(n21000) );
  NANDN U6718 ( .A(x[624]), .B(y[624]), .Z(n3532) );
  NANDN U6719 ( .A(x[623]), .B(y[623]), .Z(n3531) );
  AND U6720 ( .A(n3532), .B(n3531), .Z(n3534) );
  IV U6721 ( .A(x[625]), .Z(n5315) );
  NAND U6722 ( .A(n5315), .B(y[625]), .Z(n3533) );
  NAND U6723 ( .A(n3534), .B(n3533), .Z(n20997) );
  NANDN U6724 ( .A(x[622]), .B(y[622]), .Z(n3536) );
  NANDN U6725 ( .A(x[621]), .B(y[621]), .Z(n3535) );
  NAND U6726 ( .A(n3536), .B(n3535), .Z(n20992) );
  NANDN U6727 ( .A(x[618]), .B(y[618]), .Z(n3538) );
  NANDN U6728 ( .A(x[617]), .B(y[617]), .Z(n3537) );
  NAND U6729 ( .A(n3538), .B(n3537), .Z(n20985) );
  NANDN U6730 ( .A(x[616]), .B(y[616]), .Z(n3540) );
  NANDN U6731 ( .A(x[615]), .B(y[615]), .Z(n3539) );
  NAND U6732 ( .A(n3540), .B(n3539), .Z(n20980) );
  NANDN U6733 ( .A(x[612]), .B(y[612]), .Z(n3542) );
  NANDN U6734 ( .A(x[611]), .B(y[611]), .Z(n3541) );
  NAND U6735 ( .A(n3542), .B(n3541), .Z(n20973) );
  NANDN U6736 ( .A(x[610]), .B(y[610]), .Z(n3544) );
  NANDN U6737 ( .A(x[609]), .B(y[609]), .Z(n3543) );
  NAND U6738 ( .A(n3544), .B(n3543), .Z(n20968) );
  NANDN U6739 ( .A(x[606]), .B(y[606]), .Z(n3546) );
  NANDN U6740 ( .A(x[605]), .B(y[605]), .Z(n3545) );
  NAND U6741 ( .A(n3546), .B(n3545), .Z(n20961) );
  NANDN U6742 ( .A(y[605]), .B(x[605]), .Z(n13768) );
  NANDN U6743 ( .A(y[604]), .B(x[604]), .Z(n3547) );
  NAND U6744 ( .A(n13768), .B(n3547), .Z(n20959) );
  NANDN U6745 ( .A(x[604]), .B(y[604]), .Z(n3549) );
  NANDN U6746 ( .A(x[603]), .B(y[603]), .Z(n3548) );
  NAND U6747 ( .A(n3549), .B(n3548), .Z(n20956) );
  NANDN U6748 ( .A(y[602]), .B(x[602]), .Z(n13761) );
  IV U6749 ( .A(y[603]), .Z(n12747) );
  NAND U6750 ( .A(n12747), .B(x[603]), .Z(n13766) );
  NAND U6751 ( .A(n13761), .B(n13766), .Z(n20955) );
  NANDN U6752 ( .A(x[600]), .B(y[600]), .Z(n3551) );
  NANDN U6753 ( .A(x[599]), .B(y[599]), .Z(n3550) );
  NAND U6754 ( .A(n3551), .B(n3550), .Z(n20949) );
  NANDN U6755 ( .A(x[598]), .B(y[598]), .Z(n3553) );
  NANDN U6756 ( .A(x[597]), .B(y[597]), .Z(n3552) );
  NAND U6757 ( .A(n3553), .B(n3552), .Z(n20944) );
  NANDN U6758 ( .A(x[594]), .B(y[594]), .Z(n3555) );
  NANDN U6759 ( .A(x[593]), .B(y[593]), .Z(n3554) );
  NAND U6760 ( .A(n3555), .B(n3554), .Z(n20937) );
  ANDN U6761 ( .B(x[591]), .A(y[591]), .Z(n13748) );
  ANDN U6762 ( .B(n13745), .A(n13748), .Z(n3556) );
  ANDN U6763 ( .B(y[591]), .A(x[591]), .Z(n5241) );
  NOR U6764 ( .A(n3556), .B(n5241), .Z(n20931) );
  NANDN U6765 ( .A(x[588]), .B(y[588]), .Z(n3558) );
  NANDN U6766 ( .A(x[587]), .B(y[587]), .Z(n3557) );
  NAND U6767 ( .A(n3558), .B(n3557), .Z(n20925) );
  NANDN U6768 ( .A(x[586]), .B(y[586]), .Z(n3560) );
  NANDN U6769 ( .A(x[585]), .B(y[585]), .Z(n3559) );
  NAND U6770 ( .A(n3560), .B(n3559), .Z(n20920) );
  NANDN U6771 ( .A(x[580]), .B(y[580]), .Z(n3562) );
  NANDN U6772 ( .A(x[579]), .B(y[579]), .Z(n3561) );
  AND U6773 ( .A(n3562), .B(n3561), .Z(n3564) );
  IV U6774 ( .A(x[581]), .Z(n5219) );
  NAND U6775 ( .A(n5219), .B(y[581]), .Z(n3563) );
  NAND U6776 ( .A(n3564), .B(n3563), .Z(n20908) );
  NANDN U6777 ( .A(x[572]), .B(y[572]), .Z(n3566) );
  NANDN U6778 ( .A(x[571]), .B(y[571]), .Z(n3565) );
  AND U6779 ( .A(n3566), .B(n3565), .Z(n20892) );
  NANDN U6780 ( .A(x[570]), .B(y[570]), .Z(n3568) );
  NANDN U6781 ( .A(x[569]), .B(y[569]), .Z(n3567) );
  NAND U6782 ( .A(n3568), .B(n3567), .Z(n12751) );
  NANDN U6783 ( .A(y[569]), .B(x[569]), .Z(n12748) );
  NANDN U6784 ( .A(y[568]), .B(x[568]), .Z(n3569) );
  NAND U6785 ( .A(n12748), .B(n3569), .Z(n20887) );
  NANDN U6786 ( .A(y[566]), .B(x[566]), .Z(n3570) );
  NANDN U6787 ( .A(y[567]), .B(x[567]), .Z(n20882) );
  AND U6788 ( .A(n3570), .B(n20882), .Z(n20879) );
  NANDN U6789 ( .A(x[565]), .B(y[565]), .Z(n20876) );
  NANDN U6790 ( .A(x[566]), .B(y[566]), .Z(n20881) );
  NAND U6791 ( .A(n20876), .B(n20881), .Z(n13718) );
  NANDN U6792 ( .A(y[564]), .B(x[564]), .Z(n3572) );
  NANDN U6793 ( .A(y[565]), .B(x[565]), .Z(n3571) );
  NAND U6794 ( .A(n3572), .B(n3571), .Z(n20875) );
  NANDN U6795 ( .A(y[563]), .B(x[563]), .Z(n3574) );
  NANDN U6796 ( .A(y[562]), .B(x[562]), .Z(n3573) );
  NAND U6797 ( .A(n3574), .B(n3573), .Z(n20871) );
  ANDN U6798 ( .B(y[559]), .A(x[559]), .Z(n3576) );
  NANDN U6799 ( .A(y[558]), .B(x[558]), .Z(n3575) );
  ANDN U6800 ( .B(x[559]), .A(y[559]), .Z(n13709) );
  ANDN U6801 ( .B(n3575), .A(n13709), .Z(n13705) );
  NOR U6802 ( .A(n3576), .B(n13705), .Z(n20863) );
  NANDN U6803 ( .A(x[557]), .B(y[557]), .Z(n13703) );
  NANDN U6804 ( .A(n13708), .B(n13703), .Z(n20861) );
  NANDN U6805 ( .A(y[557]), .B(x[557]), .Z(n3578) );
  NANDN U6806 ( .A(y[556]), .B(x[556]), .Z(n3577) );
  NAND U6807 ( .A(n3578), .B(n3577), .Z(n20859) );
  NANDN U6808 ( .A(y[553]), .B(x[553]), .Z(n3580) );
  NANDN U6809 ( .A(y[552]), .B(x[552]), .Z(n3579) );
  NAND U6810 ( .A(n3580), .B(n3579), .Z(n20851) );
  NANDN U6811 ( .A(y[551]), .B(x[551]), .Z(n3582) );
  NANDN U6812 ( .A(y[550]), .B(x[550]), .Z(n3581) );
  NAND U6813 ( .A(n3582), .B(n3581), .Z(n20847) );
  NANDN U6814 ( .A(x[547]), .B(y[547]), .Z(n5162) );
  XNOR U6815 ( .A(x[547]), .B(y[547]), .Z(n3584) );
  NANDN U6816 ( .A(y[546]), .B(x[546]), .Z(n3583) );
  NAND U6817 ( .A(n3584), .B(n3583), .Z(n3585) );
  AND U6818 ( .A(n5162), .B(n3585), .Z(n20839) );
  NANDN U6819 ( .A(y[545]), .B(x[545]), .Z(n3587) );
  NANDN U6820 ( .A(y[544]), .B(x[544]), .Z(n3586) );
  NAND U6821 ( .A(n3587), .B(n3586), .Z(n20835) );
  NANDN U6822 ( .A(y[541]), .B(x[541]), .Z(n3589) );
  NANDN U6823 ( .A(y[540]), .B(x[540]), .Z(n3588) );
  NAND U6824 ( .A(n3589), .B(n3588), .Z(n20827) );
  NANDN U6825 ( .A(y[539]), .B(x[539]), .Z(n3591) );
  NANDN U6826 ( .A(y[538]), .B(x[538]), .Z(n3590) );
  NAND U6827 ( .A(n3591), .B(n3590), .Z(n20823) );
  NANDN U6828 ( .A(y[535]), .B(x[535]), .Z(n3593) );
  NANDN U6829 ( .A(y[534]), .B(x[534]), .Z(n3592) );
  NAND U6830 ( .A(n3593), .B(n3592), .Z(n20815) );
  NANDN U6831 ( .A(y[533]), .B(x[533]), .Z(n3595) );
  NANDN U6832 ( .A(y[532]), .B(x[532]), .Z(n3594) );
  NAND U6833 ( .A(n3595), .B(n3594), .Z(n20811) );
  NANDN U6834 ( .A(x[531]), .B(y[531]), .Z(n3597) );
  NANDN U6835 ( .A(x[532]), .B(y[532]), .Z(n3596) );
  NAND U6836 ( .A(n3597), .B(n3596), .Z(n12755) );
  NANDN U6837 ( .A(y[530]), .B(x[530]), .Z(n3598) );
  ANDN U6838 ( .B(x[531]), .A(y[531]), .Z(n12753) );
  ANDN U6839 ( .B(n3598), .A(n12753), .Z(n20807) );
  NANDN U6840 ( .A(y[527]), .B(x[527]), .Z(n3600) );
  NANDN U6841 ( .A(y[526]), .B(x[526]), .Z(n3599) );
  NAND U6842 ( .A(n3600), .B(n3599), .Z(n20799) );
  NANDN U6843 ( .A(y[525]), .B(x[525]), .Z(n3602) );
  NANDN U6844 ( .A(y[524]), .B(x[524]), .Z(n3601) );
  NAND U6845 ( .A(n3602), .B(n3601), .Z(n20794) );
  NANDN U6846 ( .A(y[519]), .B(x[519]), .Z(n3604) );
  NANDN U6847 ( .A(y[518]), .B(x[518]), .Z(n3603) );
  NAND U6848 ( .A(n3604), .B(n3603), .Z(n20787) );
  NANDN U6849 ( .A(y[517]), .B(x[517]), .Z(n3606) );
  NANDN U6850 ( .A(y[516]), .B(x[516]), .Z(n3605) );
  NAND U6851 ( .A(n3606), .B(n3605), .Z(n20782) );
  NANDN U6852 ( .A(x[515]), .B(y[515]), .Z(n3608) );
  NANDN U6853 ( .A(x[516]), .B(y[516]), .Z(n3607) );
  NAND U6854 ( .A(n3608), .B(n3607), .Z(n12764) );
  NANDN U6855 ( .A(y[514]), .B(x[514]), .Z(n3609) );
  ANDN U6856 ( .B(x[515]), .A(y[515]), .Z(n12762) );
  ANDN U6857 ( .B(n3609), .A(n12762), .Z(n20778) );
  NANDN U6858 ( .A(x[511]), .B(y[511]), .Z(n5085) );
  XNOR U6859 ( .A(x[511]), .B(y[511]), .Z(n3611) );
  NANDN U6860 ( .A(y[510]), .B(x[510]), .Z(n3610) );
  NAND U6861 ( .A(n3611), .B(n3610), .Z(n3612) );
  AND U6862 ( .A(n5085), .B(n3612), .Z(n20770) );
  NANDN U6863 ( .A(y[509]), .B(x[509]), .Z(n3614) );
  NANDN U6864 ( .A(y[508]), .B(x[508]), .Z(n3613) );
  NAND U6865 ( .A(n3614), .B(n3613), .Z(n20767) );
  NANDN U6866 ( .A(y[505]), .B(x[505]), .Z(n3616) );
  NANDN U6867 ( .A(y[504]), .B(x[504]), .Z(n3615) );
  NAND U6868 ( .A(n3616), .B(n3615), .Z(n20758) );
  NANDN U6869 ( .A(y[503]), .B(x[503]), .Z(n3618) );
  NANDN U6870 ( .A(y[502]), .B(x[502]), .Z(n3617) );
  NAND U6871 ( .A(n3618), .B(n3617), .Z(n20755) );
  NANDN U6872 ( .A(y[499]), .B(x[499]), .Z(n3620) );
  NANDN U6873 ( .A(y[498]), .B(x[498]), .Z(n3619) );
  NAND U6874 ( .A(n3620), .B(n3619), .Z(n20746) );
  NANDN U6875 ( .A(y[497]), .B(x[497]), .Z(n3622) );
  NANDN U6876 ( .A(y[496]), .B(x[496]), .Z(n3621) );
  NAND U6877 ( .A(n3622), .B(n3621), .Z(n20743) );
  NANDN U6878 ( .A(y[493]), .B(x[493]), .Z(n3624) );
  NANDN U6879 ( .A(y[492]), .B(x[492]), .Z(n3623) );
  NAND U6880 ( .A(n3624), .B(n3623), .Z(n20734) );
  NANDN U6881 ( .A(y[491]), .B(x[491]), .Z(n3626) );
  NANDN U6882 ( .A(y[490]), .B(x[490]), .Z(n3625) );
  NAND U6883 ( .A(n3626), .B(n3625), .Z(n20731) );
  NANDN U6884 ( .A(y[487]), .B(x[487]), .Z(n3628) );
  NANDN U6885 ( .A(y[486]), .B(x[486]), .Z(n3627) );
  NAND U6886 ( .A(n3628), .B(n3627), .Z(n20722) );
  NANDN U6887 ( .A(y[485]), .B(x[485]), .Z(n3630) );
  NANDN U6888 ( .A(y[484]), .B(x[484]), .Z(n3629) );
  NAND U6889 ( .A(n3630), .B(n3629), .Z(n20719) );
  ANDN U6890 ( .B(y[484]), .A(x[484]), .Z(n13628) );
  ANDN U6891 ( .B(y[483]), .A(x[483]), .Z(n13623) );
  NANDN U6892 ( .A(y[483]), .B(x[483]), .Z(n13625) );
  NANDN U6893 ( .A(y[482]), .B(x[482]), .Z(n3631) );
  NAND U6894 ( .A(n13625), .B(n3631), .Z(n20715) );
  NANDN U6895 ( .A(x[481]), .B(y[481]), .Z(n20712) );
  NANDN U6896 ( .A(x[478]), .B(y[478]), .Z(n3633) );
  NANDN U6897 ( .A(x[477]), .B(y[477]), .Z(n3632) );
  AND U6898 ( .A(n3633), .B(n3632), .Z(n20704) );
  NANDN U6899 ( .A(x[472]), .B(y[472]), .Z(n3635) );
  NANDN U6900 ( .A(x[471]), .B(y[471]), .Z(n3634) );
  AND U6901 ( .A(n3635), .B(n3634), .Z(n20692) );
  NANDN U6902 ( .A(x[466]), .B(y[466]), .Z(n3637) );
  NANDN U6903 ( .A(x[465]), .B(y[465]), .Z(n3636) );
  AND U6904 ( .A(n3637), .B(n3636), .Z(n20680) );
  NANDN U6905 ( .A(x[460]), .B(y[460]), .Z(n3639) );
  NANDN U6906 ( .A(x[459]), .B(y[459]), .Z(n3638) );
  AND U6907 ( .A(n3639), .B(n3638), .Z(n20668) );
  NANDN U6908 ( .A(x[453]), .B(y[453]), .Z(n3641) );
  NANDN U6909 ( .A(x[454]), .B(y[454]), .Z(n3640) );
  NAND U6910 ( .A(n3641), .B(n3640), .Z(n3644) );
  NANDN U6911 ( .A(x[452]), .B(y[452]), .Z(n3643) );
  NANDN U6912 ( .A(x[451]), .B(y[451]), .Z(n3642) );
  AND U6913 ( .A(n3643), .B(n3642), .Z(n3645) );
  ANDN U6914 ( .B(n3645), .A(n3644), .Z(n20656) );
  NANDN U6915 ( .A(x[446]), .B(y[446]), .Z(n3647) );
  NANDN U6916 ( .A(x[445]), .B(y[445]), .Z(n3646) );
  AND U6917 ( .A(n3647), .B(n3646), .Z(n20644) );
  NANDN U6918 ( .A(x[440]), .B(y[440]), .Z(n3649) );
  NANDN U6919 ( .A(x[439]), .B(y[439]), .Z(n3648) );
  AND U6920 ( .A(n3649), .B(n3648), .Z(n3651) );
  NANDN U6921 ( .A(x[441]), .B(y[441]), .Z(n3650) );
  AND U6922 ( .A(n3651), .B(n3650), .Z(n20632) );
  NANDN U6923 ( .A(y[436]), .B(x[436]), .Z(n3652) );
  NANDN U6924 ( .A(y[437]), .B(x[437]), .Z(n20627) );
  NAND U6925 ( .A(n3652), .B(n20627), .Z(n13577) );
  NANDN U6926 ( .A(x[434]), .B(y[434]), .Z(n3654) );
  NANDN U6927 ( .A(x[433]), .B(y[433]), .Z(n3653) );
  AND U6928 ( .A(n3654), .B(n3653), .Z(n20615) );
  NANDN U6929 ( .A(x[428]), .B(y[428]), .Z(n20603) );
  ANDN U6930 ( .B(y[427]), .A(x[427]), .Z(n3656) );
  NANDN U6931 ( .A(y[426]), .B(x[426]), .Z(n20598) );
  ANDN U6932 ( .B(x[427]), .A(y[427]), .Z(n20601) );
  ANDN U6933 ( .B(n20598), .A(n20601), .Z(n3655) );
  NOR U6934 ( .A(n3656), .B(n3655), .Z(n13564) );
  NANDN U6935 ( .A(x[425]), .B(y[425]), .Z(n20595) );
  NANDN U6936 ( .A(n20600), .B(n20595), .Z(n13563) );
  NANDN U6937 ( .A(x[422]), .B(y[422]), .Z(n3658) );
  NANDN U6938 ( .A(x[421]), .B(y[421]), .Z(n3657) );
  AND U6939 ( .A(n3658), .B(n3657), .Z(n20587) );
  NANDN U6940 ( .A(x[416]), .B(y[416]), .Z(n3660) );
  NANDN U6941 ( .A(x[415]), .B(y[415]), .Z(n3659) );
  AND U6942 ( .A(n3660), .B(n3659), .Z(n20575) );
  NANDN U6943 ( .A(x[410]), .B(y[410]), .Z(n3662) );
  NANDN U6944 ( .A(x[409]), .B(y[409]), .Z(n3661) );
  AND U6945 ( .A(n3662), .B(n3661), .Z(n20563) );
  NANDN U6946 ( .A(x[404]), .B(y[404]), .Z(n3664) );
  NANDN U6947 ( .A(x[403]), .B(y[403]), .Z(n3663) );
  AND U6948 ( .A(n3664), .B(n3663), .Z(n20551) );
  NANDN U6949 ( .A(x[398]), .B(y[398]), .Z(n3666) );
  NANDN U6950 ( .A(x[397]), .B(y[397]), .Z(n3665) );
  AND U6951 ( .A(n3666), .B(n3665), .Z(n20539) );
  NANDN U6952 ( .A(x[392]), .B(y[392]), .Z(n3668) );
  NANDN U6953 ( .A(x[391]), .B(y[391]), .Z(n3667) );
  AND U6954 ( .A(n3668), .B(n3667), .Z(n20527) );
  NANDN U6955 ( .A(x[386]), .B(y[386]), .Z(n3670) );
  NANDN U6956 ( .A(x[385]), .B(y[385]), .Z(n3669) );
  AND U6957 ( .A(n3670), .B(n3669), .Z(n20515) );
  NANDN U6958 ( .A(x[380]), .B(y[380]), .Z(n3672) );
  NANDN U6959 ( .A(x[379]), .B(y[379]), .Z(n3671) );
  AND U6960 ( .A(n3672), .B(n3671), .Z(n3674) );
  NANDN U6961 ( .A(x[381]), .B(y[381]), .Z(n3673) );
  AND U6962 ( .A(n3674), .B(n3673), .Z(n20503) );
  ANDN U6963 ( .B(y[378]), .A(x[378]), .Z(n12771) );
  ANDN U6964 ( .B(y[377]), .A(x[377]), .Z(n12766) );
  NANDN U6965 ( .A(y[377]), .B(x[377]), .Z(n12768) );
  NANDN U6966 ( .A(y[376]), .B(x[376]), .Z(n3675) );
  NAND U6967 ( .A(n12768), .B(n3675), .Z(n20498) );
  NANDN U6968 ( .A(x[375]), .B(y[375]), .Z(n20495) );
  NANDN U6969 ( .A(x[372]), .B(y[372]), .Z(n3681) );
  ANDN U6970 ( .B(y[370]), .A(x[370]), .Z(n3676) );
  OR U6971 ( .A(n3676), .B(y[371]), .Z(n3679) );
  XOR U6972 ( .A(y[371]), .B(n3676), .Z(n3677) );
  NAND U6973 ( .A(n3677), .B(x[371]), .Z(n3678) );
  NAND U6974 ( .A(n3679), .B(n3678), .Z(n3680) );
  AND U6975 ( .A(n3681), .B(n3680), .Z(n20487) );
  NANDN U6976 ( .A(y[371]), .B(x[371]), .Z(n3683) );
  NANDN U6977 ( .A(y[370]), .B(x[370]), .Z(n3682) );
  AND U6978 ( .A(n3683), .B(n3682), .Z(n3689) );
  NANDN U6979 ( .A(y[368]), .B(x[368]), .Z(n3684) );
  NANDN U6980 ( .A(x[369]), .B(n3684), .Z(n3687) );
  XNOR U6981 ( .A(n3684), .B(x[369]), .Z(n3685) );
  NAND U6982 ( .A(n3685), .B(y[369]), .Z(n3686) );
  NAND U6983 ( .A(n3687), .B(n3686), .Z(n3688) );
  NAND U6984 ( .A(n3689), .B(n3688), .Z(n20486) );
  ANDN U6985 ( .B(y[365]), .A(x[365]), .Z(n4728) );
  ANDN U6986 ( .B(x[365]), .A(y[365]), .Z(n20477) );
  ANDN U6987 ( .B(n20474), .A(n20477), .Z(n3690) );
  NOR U6988 ( .A(n4728), .B(n3690), .Z(n13502) );
  NANDN U6989 ( .A(x[358]), .B(y[358]), .Z(n3692) );
  NANDN U6990 ( .A(x[357]), .B(y[357]), .Z(n3691) );
  AND U6991 ( .A(n3692), .B(n3691), .Z(n20459) );
  NANDN U6992 ( .A(x[354]), .B(y[354]), .Z(n3694) );
  NANDN U6993 ( .A(x[353]), .B(y[353]), .Z(n3693) );
  NAND U6994 ( .A(n3694), .B(n3693), .Z(n13489) );
  NANDN U6995 ( .A(x[351]), .B(y[351]), .Z(n20447) );
  ANDN U6996 ( .B(y[352]), .A(x[352]), .Z(n13486) );
  ANDN U6997 ( .B(n20447), .A(n13486), .Z(n4698) );
  NANDN U6998 ( .A(x[350]), .B(y[350]), .Z(n3696) );
  NANDN U6999 ( .A(x[349]), .B(y[349]), .Z(n3695) );
  AND U7000 ( .A(n3696), .B(n3695), .Z(n20443) );
  NANDN U7001 ( .A(x[344]), .B(y[344]), .Z(n3698) );
  NANDN U7002 ( .A(x[343]), .B(y[343]), .Z(n3697) );
  AND U7003 ( .A(n3698), .B(n3697), .Z(n20431) );
  NANDN U7004 ( .A(x[338]), .B(y[338]), .Z(n3700) );
  NANDN U7005 ( .A(x[337]), .B(y[337]), .Z(n3699) );
  AND U7006 ( .A(n3700), .B(n3699), .Z(n3702) );
  NANDN U7007 ( .A(x[339]), .B(y[339]), .Z(n3701) );
  AND U7008 ( .A(n3702), .B(n3701), .Z(n20419) );
  NANDN U7009 ( .A(x[332]), .B(y[332]), .Z(n20407) );
  NANDN U7010 ( .A(x[331]), .B(y[331]), .Z(n3705) );
  ANDN U7011 ( .B(x[330]), .A(y[330]), .Z(n20303) );
  NAND U7012 ( .A(n3705), .B(n20303), .Z(n3703) );
  NANDN U7013 ( .A(y[331]), .B(x[331]), .Z(n20405) );
  NAND U7014 ( .A(n3703), .B(n20405), .Z(n13463) );
  NANDN U7015 ( .A(x[330]), .B(y[330]), .Z(n3704) );
  NAND U7016 ( .A(n3705), .B(n3704), .Z(n20404) );
  NANDN U7017 ( .A(y[328]), .B(x[328]), .Z(n20306) );
  NANDN U7018 ( .A(y[329]), .B(x[329]), .Z(n20304) );
  AND U7019 ( .A(n20306), .B(n20304), .Z(n4638) );
  NANDN U7020 ( .A(y[326]), .B(x[326]), .Z(n20394) );
  NANDN U7021 ( .A(y[327]), .B(x[327]), .Z(n20305) );
  NAND U7022 ( .A(n20394), .B(n20305), .Z(n13456) );
  NANDN U7023 ( .A(y[325]), .B(x[325]), .Z(n3707) );
  NANDN U7024 ( .A(y[324]), .B(x[324]), .Z(n3706) );
  NAND U7025 ( .A(n3707), .B(n3706), .Z(n20390) );
  NANDN U7026 ( .A(y[317]), .B(x[317]), .Z(n3709) );
  NANDN U7027 ( .A(y[316]), .B(x[316]), .Z(n3708) );
  AND U7028 ( .A(n3709), .B(n3708), .Z(n20371) );
  NANDN U7029 ( .A(x[313]), .B(y[313]), .Z(n4598) );
  NANDN U7030 ( .A(y[313]), .B(x[313]), .Z(n20363) );
  NANDN U7031 ( .A(y[312]), .B(x[312]), .Z(n3710) );
  AND U7032 ( .A(n20363), .B(n3710), .Z(n3711) );
  ANDN U7033 ( .B(n4598), .A(n3711), .Z(n13439) );
  NANDN U7034 ( .A(x[310]), .B(y[310]), .Z(n3713) );
  NANDN U7035 ( .A(x[309]), .B(y[309]), .Z(n3712) );
  NAND U7036 ( .A(n3713), .B(n3712), .Z(n20353) );
  NANDN U7037 ( .A(x[306]), .B(y[306]), .Z(n3715) );
  NANDN U7038 ( .A(x[305]), .B(y[305]), .Z(n3714) );
  NAND U7039 ( .A(n3715), .B(n3714), .Z(n20346) );
  NANDN U7040 ( .A(x[304]), .B(y[304]), .Z(n3717) );
  NANDN U7041 ( .A(x[303]), .B(y[303]), .Z(n3716) );
  NAND U7042 ( .A(n3717), .B(n3716), .Z(n20341) );
  NANDN U7043 ( .A(x[300]), .B(y[300]), .Z(n3719) );
  NANDN U7044 ( .A(x[299]), .B(y[299]), .Z(n3718) );
  NAND U7045 ( .A(n3719), .B(n3718), .Z(n20334) );
  NANDN U7046 ( .A(x[298]), .B(y[298]), .Z(n3721) );
  NANDN U7047 ( .A(x[297]), .B(y[297]), .Z(n3720) );
  NAND U7048 ( .A(n3721), .B(n3720), .Z(n20329) );
  NANDN U7049 ( .A(x[294]), .B(y[294]), .Z(n3723) );
  NANDN U7050 ( .A(x[293]), .B(y[293]), .Z(n3722) );
  NAND U7051 ( .A(n3723), .B(n3722), .Z(n20322) );
  NANDN U7052 ( .A(x[292]), .B(y[292]), .Z(n3725) );
  NANDN U7053 ( .A(x[291]), .B(y[291]), .Z(n3724) );
  AND U7054 ( .A(n3725), .B(n3724), .Z(n3732) );
  NANDN U7055 ( .A(x[289]), .B(y[289]), .Z(n3727) );
  NANDN U7056 ( .A(x[290]), .B(y[290]), .Z(n3726) );
  AND U7057 ( .A(n3727), .B(n3726), .Z(n3730) );
  NANDN U7058 ( .A(y[291]), .B(x[291]), .Z(n3729) );
  NANDN U7059 ( .A(y[290]), .B(x[290]), .Z(n3728) );
  AND U7060 ( .A(n3729), .B(n3728), .Z(n3733) );
  NANDN U7061 ( .A(n3730), .B(n3733), .Z(n3731) );
  NAND U7062 ( .A(n3732), .B(n3731), .Z(n20317) );
  NANDN U7063 ( .A(y[289]), .B(x[289]), .Z(n3734) );
  NAND U7064 ( .A(n3734), .B(n3733), .Z(n20316) );
  NANDN U7065 ( .A(y[288]), .B(x[288]), .Z(n20311) );
  NANDN U7066 ( .A(n20316), .B(n20311), .Z(n13416) );
  NANDN U7067 ( .A(x[288]), .B(y[288]), .Z(n20313) );
  ANDN U7068 ( .B(y[287]), .A(x[287]), .Z(n4547) );
  NANDN U7069 ( .A(y[286]), .B(x[286]), .Z(n13410) );
  ANDN U7070 ( .B(x[287]), .A(y[287]), .Z(n13412) );
  ANDN U7071 ( .B(n13410), .A(n13412), .Z(n3735) );
  NOR U7072 ( .A(n4547), .B(n3735), .Z(n20309) );
  NANDN U7073 ( .A(y[284]), .B(x[284]), .Z(n3736) );
  NANDN U7074 ( .A(n3736), .B(x[285]), .Z(n3739) );
  IV U7075 ( .A(x[285]), .Z(n4542) );
  XOR U7076 ( .A(n3736), .B(n4542), .Z(n3737) );
  NANDN U7077 ( .A(y[285]), .B(n3737), .Z(n3738) );
  NAND U7078 ( .A(n3739), .B(n3738), .Z(n13408) );
  NANDN U7079 ( .A(y[282]), .B(x[282]), .Z(n3741) );
  NANDN U7080 ( .A(y[283]), .B(x[283]), .Z(n3740) );
  NAND U7081 ( .A(n3741), .B(n3740), .Z(n13404) );
  NANDN U7082 ( .A(x[282]), .B(y[282]), .Z(n3743) );
  NANDN U7083 ( .A(x[281]), .B(y[281]), .Z(n3742) );
  AND U7084 ( .A(n3743), .B(n3742), .Z(n13402) );
  NANDN U7085 ( .A(y[280]), .B(x[280]), .Z(n3745) );
  NANDN U7086 ( .A(y[281]), .B(x[281]), .Z(n3744) );
  NAND U7087 ( .A(n3745), .B(n3744), .Z(n13401) );
  NANDN U7088 ( .A(y[278]), .B(x[278]), .Z(n3747) );
  NANDN U7089 ( .A(y[279]), .B(x[279]), .Z(n3746) );
  NAND U7090 ( .A(n3747), .B(n3746), .Z(n13397) );
  NANDN U7091 ( .A(y[276]), .B(x[276]), .Z(n3749) );
  NANDN U7092 ( .A(y[277]), .B(x[277]), .Z(n3748) );
  NAND U7093 ( .A(n3749), .B(n3748), .Z(n13392) );
  NANDN U7094 ( .A(x[276]), .B(y[276]), .Z(n3751) );
  NANDN U7095 ( .A(x[275]), .B(y[275]), .Z(n3750) );
  AND U7096 ( .A(n3751), .B(n3750), .Z(n13390) );
  NANDN U7097 ( .A(y[274]), .B(x[274]), .Z(n3753) );
  NANDN U7098 ( .A(y[275]), .B(x[275]), .Z(n3752) );
  NAND U7099 ( .A(n3753), .B(n3752), .Z(n13389) );
  NANDN U7100 ( .A(y[272]), .B(x[272]), .Z(n3754) );
  NANDN U7101 ( .A(n3754), .B(x[273]), .Z(n3757) );
  IV U7102 ( .A(x[273]), .Z(n4521) );
  XOR U7103 ( .A(n3754), .B(n4521), .Z(n3755) );
  NANDN U7104 ( .A(y[273]), .B(n3755), .Z(n3756) );
  NAND U7105 ( .A(n3757), .B(n3756), .Z(n13385) );
  NANDN U7106 ( .A(x[269]), .B(y[269]), .Z(n13374) );
  NANDN U7107 ( .A(x[270]), .B(y[270]), .Z(n3758) );
  AND U7108 ( .A(n13374), .B(n3758), .Z(n4515) );
  NANDN U7109 ( .A(y[269]), .B(x[269]), .Z(n3760) );
  NANDN U7110 ( .A(y[268]), .B(x[268]), .Z(n3759) );
  NAND U7111 ( .A(n3760), .B(n3759), .Z(n13373) );
  NANDN U7112 ( .A(x[268]), .B(y[268]), .Z(n3762) );
  NANDN U7113 ( .A(x[267]), .B(y[267]), .Z(n3761) );
  AND U7114 ( .A(n3762), .B(n3761), .Z(n13370) );
  NANDN U7115 ( .A(y[266]), .B(x[266]), .Z(n3764) );
  NANDN U7116 ( .A(y[267]), .B(x[267]), .Z(n3763) );
  NAND U7117 ( .A(n3764), .B(n3763), .Z(n13368) );
  NANDN U7118 ( .A(y[264]), .B(x[264]), .Z(n3766) );
  ANDN U7119 ( .B(x[265]), .A(y[265]), .Z(n3765) );
  ANDN U7120 ( .B(n3766), .A(n3765), .Z(n3770) );
  XNOR U7121 ( .A(x[264]), .B(y[264]), .Z(n3768) );
  ANDN U7122 ( .B(x[263]), .A(y[263]), .Z(n3767) );
  NAND U7123 ( .A(n3768), .B(n3767), .Z(n3769) );
  NAND U7124 ( .A(n3770), .B(n3769), .Z(n13365) );
  NANDN U7125 ( .A(y[261]), .B(x[261]), .Z(n3772) );
  ANDN U7126 ( .B(x[262]), .A(y[262]), .Z(n3771) );
  ANDN U7127 ( .B(n3772), .A(n3771), .Z(n3776) );
  XNOR U7128 ( .A(x[261]), .B(y[261]), .Z(n3774) );
  ANDN U7129 ( .B(x[260]), .A(y[260]), .Z(n3773) );
  NAND U7130 ( .A(n3774), .B(n3773), .Z(n3775) );
  NAND U7131 ( .A(n3776), .B(n3775), .Z(n13361) );
  NANDN U7132 ( .A(x[260]), .B(y[260]), .Z(n3778) );
  NANDN U7133 ( .A(x[259]), .B(y[259]), .Z(n3777) );
  AND U7134 ( .A(n3778), .B(n3777), .Z(n3780) );
  NANDN U7135 ( .A(x[261]), .B(y[261]), .Z(n3779) );
  AND U7136 ( .A(n3780), .B(n3779), .Z(n13358) );
  NANDN U7137 ( .A(y[258]), .B(x[258]), .Z(n3782) );
  NANDN U7138 ( .A(y[259]), .B(x[259]), .Z(n3781) );
  NAND U7139 ( .A(n3782), .B(n3781), .Z(n13356) );
  NANDN U7140 ( .A(y[256]), .B(x[256]), .Z(n3784) );
  NANDN U7141 ( .A(y[257]), .B(x[257]), .Z(n3783) );
  NAND U7142 ( .A(n3784), .B(n3783), .Z(n13353) );
  NANDN U7143 ( .A(y[254]), .B(x[254]), .Z(n3786) );
  NANDN U7144 ( .A(y[255]), .B(x[255]), .Z(n3785) );
  NAND U7145 ( .A(n3786), .B(n3785), .Z(n13349) );
  NANDN U7146 ( .A(x[254]), .B(y[254]), .Z(n3788) );
  NANDN U7147 ( .A(x[253]), .B(y[253]), .Z(n3787) );
  AND U7148 ( .A(n3788), .B(n3787), .Z(n13346) );
  NANDN U7149 ( .A(y[252]), .B(x[252]), .Z(n3790) );
  NANDN U7150 ( .A(y[253]), .B(x[253]), .Z(n3789) );
  NAND U7151 ( .A(n3790), .B(n3789), .Z(n13344) );
  NANDN U7152 ( .A(y[250]), .B(x[250]), .Z(n3792) );
  NANDN U7153 ( .A(y[251]), .B(x[251]), .Z(n3791) );
  NAND U7154 ( .A(n3792), .B(n3791), .Z(n13341) );
  NANDN U7155 ( .A(y[248]), .B(x[248]), .Z(n3794) );
  NANDN U7156 ( .A(y[249]), .B(x[249]), .Z(n3793) );
  NAND U7157 ( .A(n3794), .B(n3793), .Z(n13337) );
  NANDN U7158 ( .A(y[247]), .B(x[247]), .Z(n3798) );
  XNOR U7159 ( .A(y[247]), .B(x[247]), .Z(n3796) );
  NANDN U7160 ( .A(x[246]), .B(y[246]), .Z(n3795) );
  NAND U7161 ( .A(n3796), .B(n3795), .Z(n3797) );
  NAND U7162 ( .A(n3798), .B(n3797), .Z(n3800) );
  NANDN U7163 ( .A(x[248]), .B(y[248]), .Z(n3799) );
  AND U7164 ( .A(n3800), .B(n3799), .Z(n13334) );
  ANDN U7165 ( .B(x[247]), .A(y[247]), .Z(n3806) );
  NANDN U7166 ( .A(y[244]), .B(x[244]), .Z(n3801) );
  NANDN U7167 ( .A(n3801), .B(x[245]), .Z(n3804) );
  IV U7168 ( .A(x[245]), .Z(n4475) );
  XOR U7169 ( .A(n3801), .B(n4475), .Z(n3802) );
  NANDN U7170 ( .A(y[245]), .B(n3802), .Z(n3803) );
  NAND U7171 ( .A(n3804), .B(n3803), .Z(n3805) );
  NOR U7172 ( .A(n3806), .B(n3805), .Z(n3808) );
  NANDN U7173 ( .A(y[246]), .B(x[246]), .Z(n3807) );
  NAND U7174 ( .A(n3808), .B(n3807), .Z(n13332) );
  NANDN U7175 ( .A(y[242]), .B(x[242]), .Z(n3810) );
  NANDN U7176 ( .A(y[243]), .B(x[243]), .Z(n3809) );
  NAND U7177 ( .A(n3810), .B(n3809), .Z(n13329) );
  NANDN U7178 ( .A(y[240]), .B(x[240]), .Z(n3812) );
  NANDN U7179 ( .A(y[241]), .B(x[241]), .Z(n3811) );
  NAND U7180 ( .A(n3812), .B(n3811), .Z(n13325) );
  NANDN U7181 ( .A(x[240]), .B(y[240]), .Z(n3814) );
  NANDN U7182 ( .A(x[239]), .B(y[239]), .Z(n3813) );
  AND U7183 ( .A(n3814), .B(n3813), .Z(n13322) );
  NANDN U7184 ( .A(y[238]), .B(x[238]), .Z(n3816) );
  NANDN U7185 ( .A(y[239]), .B(x[239]), .Z(n3815) );
  NAND U7186 ( .A(n3816), .B(n3815), .Z(n13320) );
  NANDN U7187 ( .A(y[236]), .B(x[236]), .Z(n3818) );
  NANDN U7188 ( .A(y[237]), .B(x[237]), .Z(n3817) );
  NAND U7189 ( .A(n3818), .B(n3817), .Z(n13317) );
  NANDN U7190 ( .A(y[234]), .B(x[234]), .Z(n3820) );
  NANDN U7191 ( .A(y[235]), .B(x[235]), .Z(n3819) );
  NAND U7192 ( .A(n3820), .B(n3819), .Z(n13313) );
  NANDN U7193 ( .A(x[234]), .B(y[234]), .Z(n3822) );
  NANDN U7194 ( .A(x[233]), .B(y[233]), .Z(n3821) );
  AND U7195 ( .A(n3822), .B(n3821), .Z(n13310) );
  NANDN U7196 ( .A(y[232]), .B(x[232]), .Z(n3824) );
  NANDN U7197 ( .A(y[233]), .B(x[233]), .Z(n3823) );
  NAND U7198 ( .A(n3824), .B(n3823), .Z(n13308) );
  NANDN U7199 ( .A(y[230]), .B(x[230]), .Z(n3826) );
  NANDN U7200 ( .A(y[231]), .B(x[231]), .Z(n3825) );
  NAND U7201 ( .A(n3826), .B(n3825), .Z(n13305) );
  NANDN U7202 ( .A(y[228]), .B(x[228]), .Z(n3828) );
  NANDN U7203 ( .A(y[229]), .B(x[229]), .Z(n3827) );
  NAND U7204 ( .A(n3828), .B(n3827), .Z(n13301) );
  NANDN U7205 ( .A(x[228]), .B(y[228]), .Z(n3830) );
  NANDN U7206 ( .A(x[227]), .B(y[227]), .Z(n3829) );
  AND U7207 ( .A(n3830), .B(n3829), .Z(n13298) );
  ANDN U7208 ( .B(x[225]), .A(y[225]), .Z(n13290) );
  NANDN U7209 ( .A(y[224]), .B(x[224]), .Z(n13283) );
  NANDN U7210 ( .A(x[224]), .B(y[224]), .Z(n13286) );
  NANDN U7211 ( .A(x[223]), .B(y[223]), .Z(n3836) );
  XNOR U7212 ( .A(x[223]), .B(y[223]), .Z(n3832) );
  NANDN U7213 ( .A(y[222]), .B(x[222]), .Z(n3831) );
  NAND U7214 ( .A(n3832), .B(n3831), .Z(n3833) );
  AND U7215 ( .A(n3836), .B(n3833), .Z(n13281) );
  NANDN U7216 ( .A(x[222]), .B(y[222]), .Z(n3835) );
  NANDN U7217 ( .A(x[221]), .B(y[221]), .Z(n3834) );
  AND U7218 ( .A(n3835), .B(n3834), .Z(n3837) );
  NAND U7219 ( .A(n3837), .B(n3836), .Z(n13280) );
  NANDN U7220 ( .A(y[221]), .B(x[221]), .Z(n3839) );
  NANDN U7221 ( .A(y[220]), .B(x[220]), .Z(n3838) );
  NAND U7222 ( .A(n3839), .B(n3838), .Z(n13278) );
  NANDN U7223 ( .A(x[219]), .B(y[219]), .Z(n3841) );
  NANDN U7224 ( .A(x[220]), .B(y[220]), .Z(n3840) );
  NAND U7225 ( .A(n3841), .B(n3840), .Z(n13276) );
  NANDN U7226 ( .A(x[217]), .B(y[217]), .Z(n3843) );
  NANDN U7227 ( .A(x[218]), .B(y[218]), .Z(n3842) );
  NAND U7228 ( .A(n3843), .B(n3842), .Z(n13272) );
  ANDN U7229 ( .B(x[217]), .A(y[217]), .Z(n13269) );
  NANDN U7230 ( .A(y[214]), .B(x[214]), .Z(n3845) );
  NANDN U7231 ( .A(y[215]), .B(x[215]), .Z(n3844) );
  NAND U7232 ( .A(n3845), .B(n3844), .Z(n13262) );
  NANDN U7233 ( .A(x[213]), .B(y[213]), .Z(n3847) );
  NANDN U7234 ( .A(x[214]), .B(y[214]), .Z(n3846) );
  NAND U7235 ( .A(n3847), .B(n3846), .Z(n13260) );
  NANDN U7236 ( .A(y[213]), .B(x[213]), .Z(n3849) );
  NANDN U7237 ( .A(y[212]), .B(x[212]), .Z(n3848) );
  NAND U7238 ( .A(n3849), .B(n3848), .Z(n13257) );
  NANDN U7239 ( .A(x[211]), .B(y[211]), .Z(n3851) );
  NANDN U7240 ( .A(x[212]), .B(y[212]), .Z(n3850) );
  NAND U7241 ( .A(n3851), .B(n3850), .Z(n13256) );
  NANDN U7242 ( .A(x[210]), .B(y[210]), .Z(n3853) );
  NANDN U7243 ( .A(x[209]), .B(y[209]), .Z(n3852) );
  AND U7244 ( .A(n3853), .B(n3852), .Z(n3863) );
  NANDN U7245 ( .A(y[208]), .B(x[208]), .Z(n3855) );
  NANDN U7246 ( .A(y[209]), .B(x[209]), .Z(n3854) );
  NAND U7247 ( .A(n3855), .B(n3854), .Z(n4429) );
  ANDN U7248 ( .B(y[206]), .A(x[206]), .Z(n3856) );
  OR U7249 ( .A(n3856), .B(y[207]), .Z(n3859) );
  XOR U7250 ( .A(y[207]), .B(n3856), .Z(n3857) );
  NAND U7251 ( .A(n3857), .B(x[207]), .Z(n3858) );
  NAND U7252 ( .A(n3859), .B(n3858), .Z(n3860) );
  ANDN U7253 ( .B(y[208]), .A(x[208]), .Z(n12775) );
  ANDN U7254 ( .B(n3860), .A(n12775), .Z(n3861) );
  OR U7255 ( .A(n4429), .B(n3861), .Z(n3862) );
  NAND U7256 ( .A(n3863), .B(n3862), .Z(n13252) );
  ANDN U7257 ( .B(x[207]), .A(y[207]), .Z(n12774) );
  NANDN U7258 ( .A(x[204]), .B(y[204]), .Z(n3865) );
  NANDN U7259 ( .A(x[203]), .B(y[203]), .Z(n3864) );
  AND U7260 ( .A(n3865), .B(n3864), .Z(n3867) );
  IV U7261 ( .A(x[205]), .Z(n4424) );
  NAND U7262 ( .A(n4424), .B(y[205]), .Z(n3866) );
  NAND U7263 ( .A(n3867), .B(n3866), .Z(n13248) );
  NANDN U7264 ( .A(y[203]), .B(x[203]), .Z(n3869) );
  NANDN U7265 ( .A(y[202]), .B(x[202]), .Z(n3868) );
  NAND U7266 ( .A(n3869), .B(n3868), .Z(n13246) );
  NANDN U7267 ( .A(x[201]), .B(y[201]), .Z(n3871) );
  NANDN U7268 ( .A(x[202]), .B(y[202]), .Z(n3870) );
  NAND U7269 ( .A(n3871), .B(n3870), .Z(n13244) );
  NANDN U7270 ( .A(y[201]), .B(x[201]), .Z(n3873) );
  NANDN U7271 ( .A(y[200]), .B(x[200]), .Z(n3872) );
  NAND U7272 ( .A(n3873), .B(n3872), .Z(n13241) );
  NANDN U7273 ( .A(x[199]), .B(y[199]), .Z(n3875) );
  ANDN U7274 ( .B(y[200]), .A(x[200]), .Z(n3874) );
  ANDN U7275 ( .B(n3875), .A(n3874), .Z(n3879) );
  XNOR U7276 ( .A(y[199]), .B(x[199]), .Z(n3877) );
  ANDN U7277 ( .B(y[198]), .A(x[198]), .Z(n3876) );
  NAND U7278 ( .A(n3877), .B(n3876), .Z(n3878) );
  NAND U7279 ( .A(n3879), .B(n3878), .Z(n13240) );
  NANDN U7280 ( .A(x[196]), .B(y[196]), .Z(n3881) );
  NANDN U7281 ( .A(x[195]), .B(y[195]), .Z(n3880) );
  AND U7282 ( .A(n3881), .B(n3880), .Z(n3883) );
  NANDN U7283 ( .A(x[197]), .B(y[197]), .Z(n3882) );
  NAND U7284 ( .A(n3883), .B(n3882), .Z(n13236) );
  NANDN U7285 ( .A(y[195]), .B(x[195]), .Z(n3885) );
  NANDN U7286 ( .A(y[194]), .B(x[194]), .Z(n3884) );
  NAND U7287 ( .A(n3885), .B(n3884), .Z(n13234) );
  NANDN U7288 ( .A(x[193]), .B(y[193]), .Z(n3887) );
  NANDN U7289 ( .A(x[194]), .B(y[194]), .Z(n3886) );
  NAND U7290 ( .A(n3887), .B(n3886), .Z(n13232) );
  NANDN U7291 ( .A(y[193]), .B(x[193]), .Z(n3889) );
  NANDN U7292 ( .A(y[192]), .B(x[192]), .Z(n3888) );
  NAND U7293 ( .A(n3889), .B(n3888), .Z(n13229) );
  NANDN U7294 ( .A(x[191]), .B(y[191]), .Z(n3891) );
  NANDN U7295 ( .A(x[192]), .B(y[192]), .Z(n3890) );
  NAND U7296 ( .A(n3891), .B(n3890), .Z(n13228) );
  NANDN U7297 ( .A(x[189]), .B(y[189]), .Z(n3893) );
  NANDN U7298 ( .A(x[190]), .B(y[190]), .Z(n3892) );
  NAND U7299 ( .A(n3893), .B(n3892), .Z(n13224) );
  NANDN U7300 ( .A(y[189]), .B(x[189]), .Z(n3895) );
  NANDN U7301 ( .A(y[188]), .B(x[188]), .Z(n3894) );
  NAND U7302 ( .A(n3895), .B(n3894), .Z(n13222) );
  NANDN U7303 ( .A(x[187]), .B(y[187]), .Z(n3897) );
  NANDN U7304 ( .A(x[188]), .B(y[188]), .Z(n3896) );
  NAND U7305 ( .A(n3897), .B(n3896), .Z(n13220) );
  ANDN U7306 ( .B(y[185]), .A(x[185]), .Z(n13211) );
  IV U7307 ( .A(x[186]), .Z(n13212) );
  AND U7308 ( .A(y[186]), .B(n13212), .Z(n4394) );
  NANDN U7309 ( .A(x[183]), .B(y[183]), .Z(n3899) );
  NANDN U7310 ( .A(x[184]), .B(y[184]), .Z(n3898) );
  NAND U7311 ( .A(n3899), .B(n3898), .Z(n13207) );
  NANDN U7312 ( .A(y[183]), .B(x[183]), .Z(n3901) );
  NANDN U7313 ( .A(y[182]), .B(x[182]), .Z(n3900) );
  AND U7314 ( .A(n3901), .B(n3900), .Z(n13204) );
  NANDN U7315 ( .A(x[181]), .B(y[181]), .Z(n3903) );
  NANDN U7316 ( .A(x[182]), .B(y[182]), .Z(n3902) );
  NAND U7317 ( .A(n3903), .B(n3902), .Z(n13202) );
  NANDN U7318 ( .A(x[179]), .B(y[179]), .Z(n3905) );
  NANDN U7319 ( .A(x[180]), .B(y[180]), .Z(n3904) );
  NAND U7320 ( .A(n3905), .B(n3904), .Z(n13199) );
  ANDN U7321 ( .B(y[178]), .A(x[178]), .Z(n13195) );
  NANDN U7322 ( .A(x[177]), .B(y[177]), .Z(n3913) );
  XNOR U7323 ( .A(x[177]), .B(y[177]), .Z(n3907) );
  NANDN U7324 ( .A(y[176]), .B(x[176]), .Z(n3906) );
  NAND U7325 ( .A(n3907), .B(n3906), .Z(n3908) );
  NAND U7326 ( .A(n3913), .B(n3908), .Z(n3910) );
  NANDN U7327 ( .A(y[178]), .B(x[178]), .Z(n3909) );
  AND U7328 ( .A(n3910), .B(n3909), .Z(n13192) );
  NANDN U7329 ( .A(x[176]), .B(y[176]), .Z(n3912) );
  NANDN U7330 ( .A(x[175]), .B(y[175]), .Z(n3911) );
  AND U7331 ( .A(n3912), .B(n3911), .Z(n3914) );
  NAND U7332 ( .A(n3914), .B(n3913), .Z(n13190) );
  NANDN U7333 ( .A(x[173]), .B(y[173]), .Z(n3916) );
  NANDN U7334 ( .A(x[174]), .B(y[174]), .Z(n3915) );
  NAND U7335 ( .A(n3916), .B(n3915), .Z(n13187) );
  NANDN U7336 ( .A(x[171]), .B(y[171]), .Z(n3918) );
  NANDN U7337 ( .A(x[172]), .B(y[172]), .Z(n3917) );
  NAND U7338 ( .A(n3918), .B(n3917), .Z(n13183) );
  NANDN U7339 ( .A(y[171]), .B(x[171]), .Z(n3920) );
  NANDN U7340 ( .A(y[170]), .B(x[170]), .Z(n3919) );
  AND U7341 ( .A(n3920), .B(n3919), .Z(n13180) );
  ANDN U7342 ( .B(y[170]), .A(x[170]), .Z(n13178) );
  NANDN U7343 ( .A(x[168]), .B(y[168]), .Z(n3922) );
  NANDN U7344 ( .A(x[167]), .B(y[167]), .Z(n3921) );
  AND U7345 ( .A(n3922), .B(n3921), .Z(n3923) );
  NANDN U7346 ( .A(x[169]), .B(y[169]), .Z(n4367) );
  NAND U7347 ( .A(n3923), .B(n4367), .Z(n13175) );
  NANDN U7348 ( .A(x[165]), .B(y[165]), .Z(n3925) );
  NANDN U7349 ( .A(x[166]), .B(y[166]), .Z(n3924) );
  NAND U7350 ( .A(n3925), .B(n3924), .Z(n13171) );
  NANDN U7351 ( .A(y[165]), .B(x[165]), .Z(n3927) );
  NANDN U7352 ( .A(y[164]), .B(x[164]), .Z(n3926) );
  AND U7353 ( .A(n3927), .B(n3926), .Z(n13168) );
  NANDN U7354 ( .A(x[163]), .B(y[163]), .Z(n3929) );
  NANDN U7355 ( .A(x[164]), .B(y[164]), .Z(n3928) );
  NAND U7356 ( .A(n3929), .B(n3928), .Z(n13166) );
  NANDN U7357 ( .A(x[161]), .B(y[161]), .Z(n3931) );
  NANDN U7358 ( .A(x[162]), .B(y[162]), .Z(n3930) );
  NAND U7359 ( .A(n3931), .B(n3930), .Z(n13163) );
  ANDN U7360 ( .B(y[159]), .A(x[159]), .Z(n13155) );
  ANDN U7361 ( .B(y[160]), .A(x[160]), .Z(n4348) );
  NANDN U7362 ( .A(x[157]), .B(y[157]), .Z(n3933) );
  NANDN U7363 ( .A(x[158]), .B(y[158]), .Z(n3932) );
  NAND U7364 ( .A(n3933), .B(n3932), .Z(n13151) );
  NANDN U7365 ( .A(y[157]), .B(x[157]), .Z(n3935) );
  NANDN U7366 ( .A(y[156]), .B(x[156]), .Z(n3934) );
  AND U7367 ( .A(n3935), .B(n3934), .Z(n13148) );
  NANDN U7368 ( .A(x[155]), .B(y[155]), .Z(n3937) );
  NANDN U7369 ( .A(x[156]), .B(y[156]), .Z(n3936) );
  NAND U7370 ( .A(n3937), .B(n3936), .Z(n13147) );
  NANDN U7371 ( .A(x[153]), .B(y[153]), .Z(n3939) );
  NANDN U7372 ( .A(x[154]), .B(y[154]), .Z(n3938) );
  NAND U7373 ( .A(n3939), .B(n3938), .Z(n13142) );
  NANDN U7374 ( .A(x[151]), .B(y[151]), .Z(n3941) );
  NANDN U7375 ( .A(x[152]), .B(y[152]), .Z(n3940) );
  NAND U7376 ( .A(n3941), .B(n3940), .Z(n13139) );
  NANDN U7377 ( .A(y[151]), .B(x[151]), .Z(n3943) );
  NANDN U7378 ( .A(y[150]), .B(x[150]), .Z(n3942) );
  AND U7379 ( .A(n3943), .B(n3942), .Z(n13136) );
  NANDN U7380 ( .A(x[149]), .B(y[149]), .Z(n3945) );
  NANDN U7381 ( .A(x[150]), .B(y[150]), .Z(n3944) );
  NAND U7382 ( .A(n3945), .B(n3944), .Z(n13135) );
  NANDN U7383 ( .A(x[147]), .B(y[147]), .Z(n3947) );
  NANDN U7384 ( .A(x[148]), .B(y[148]), .Z(n3946) );
  NAND U7385 ( .A(n3947), .B(n3946), .Z(n13130) );
  NANDN U7386 ( .A(x[145]), .B(y[145]), .Z(n3949) );
  NANDN U7387 ( .A(x[146]), .B(y[146]), .Z(n3948) );
  NAND U7388 ( .A(n3949), .B(n3948), .Z(n13127) );
  NANDN U7389 ( .A(y[145]), .B(x[145]), .Z(n3951) );
  NANDN U7390 ( .A(y[144]), .B(x[144]), .Z(n3950) );
  AND U7391 ( .A(n3951), .B(n3950), .Z(n13124) );
  NANDN U7392 ( .A(x[143]), .B(y[143]), .Z(n3953) );
  NANDN U7393 ( .A(x[144]), .B(y[144]), .Z(n3952) );
  NAND U7394 ( .A(n3953), .B(n3952), .Z(n13123) );
  NANDN U7395 ( .A(x[141]), .B(y[141]), .Z(n3955) );
  NANDN U7396 ( .A(x[142]), .B(y[142]), .Z(n3954) );
  NAND U7397 ( .A(n3955), .B(n3954), .Z(n13118) );
  NANDN U7398 ( .A(x[139]), .B(y[139]), .Z(n3957) );
  NANDN U7399 ( .A(x[140]), .B(y[140]), .Z(n3956) );
  NAND U7400 ( .A(n3957), .B(n3956), .Z(n13115) );
  NANDN U7401 ( .A(y[139]), .B(x[139]), .Z(n3959) );
  NANDN U7402 ( .A(y[138]), .B(x[138]), .Z(n3958) );
  AND U7403 ( .A(n3959), .B(n3958), .Z(n13112) );
  NANDN U7404 ( .A(x[137]), .B(y[137]), .Z(n3961) );
  NANDN U7405 ( .A(x[138]), .B(y[138]), .Z(n3960) );
  NAND U7406 ( .A(n3961), .B(n3960), .Z(n13111) );
  NANDN U7407 ( .A(x[135]), .B(y[135]), .Z(n3963) );
  NANDN U7408 ( .A(x[136]), .B(y[136]), .Z(n3962) );
  NAND U7409 ( .A(n3963), .B(n3962), .Z(n13106) );
  NANDN U7410 ( .A(x[133]), .B(y[133]), .Z(n3965) );
  NANDN U7411 ( .A(x[134]), .B(y[134]), .Z(n3964) );
  NAND U7412 ( .A(n3965), .B(n3964), .Z(n13103) );
  NANDN U7413 ( .A(y[133]), .B(x[133]), .Z(n3967) );
  NANDN U7414 ( .A(y[132]), .B(x[132]), .Z(n3966) );
  AND U7415 ( .A(n3967), .B(n3966), .Z(n13100) );
  NANDN U7416 ( .A(x[131]), .B(y[131]), .Z(n3969) );
  NANDN U7417 ( .A(x[132]), .B(y[132]), .Z(n3968) );
  NAND U7418 ( .A(n3969), .B(n3968), .Z(n13099) );
  NANDN U7419 ( .A(x[129]), .B(y[129]), .Z(n3971) );
  NANDN U7420 ( .A(x[130]), .B(y[130]), .Z(n3970) );
  NAND U7421 ( .A(n3971), .B(n3970), .Z(n13094) );
  NANDN U7422 ( .A(x[127]), .B(y[127]), .Z(n3973) );
  NANDN U7423 ( .A(x[128]), .B(y[128]), .Z(n3972) );
  NAND U7424 ( .A(n3973), .B(n3972), .Z(n13091) );
  NANDN U7425 ( .A(y[127]), .B(x[127]), .Z(n3975) );
  NANDN U7426 ( .A(y[126]), .B(x[126]), .Z(n3974) );
  AND U7427 ( .A(n3975), .B(n3974), .Z(n13088) );
  NANDN U7428 ( .A(x[125]), .B(y[125]), .Z(n3977) );
  NANDN U7429 ( .A(x[126]), .B(y[126]), .Z(n3976) );
  NAND U7430 ( .A(n3977), .B(n3976), .Z(n13087) );
  NANDN U7431 ( .A(x[123]), .B(y[123]), .Z(n3979) );
  NANDN U7432 ( .A(x[124]), .B(y[124]), .Z(n3978) );
  NAND U7433 ( .A(n3979), .B(n3978), .Z(n13082) );
  NANDN U7434 ( .A(x[121]), .B(y[121]), .Z(n3981) );
  NANDN U7435 ( .A(x[122]), .B(y[122]), .Z(n3980) );
  NAND U7436 ( .A(n3981), .B(n3980), .Z(n13079) );
  NANDN U7437 ( .A(y[121]), .B(x[121]), .Z(n3983) );
  NANDN U7438 ( .A(y[120]), .B(x[120]), .Z(n3982) );
  AND U7439 ( .A(n3983), .B(n3982), .Z(n13076) );
  NANDN U7440 ( .A(x[119]), .B(y[119]), .Z(n3985) );
  NANDN U7441 ( .A(x[120]), .B(y[120]), .Z(n3984) );
  NAND U7442 ( .A(n3985), .B(n3984), .Z(n13075) );
  NANDN U7443 ( .A(x[117]), .B(y[117]), .Z(n3987) );
  NANDN U7444 ( .A(x[118]), .B(y[118]), .Z(n3986) );
  NAND U7445 ( .A(n3987), .B(n3986), .Z(n13070) );
  NANDN U7446 ( .A(x[115]), .B(y[115]), .Z(n3989) );
  NANDN U7447 ( .A(x[116]), .B(y[116]), .Z(n3988) );
  NAND U7448 ( .A(n3989), .B(n3988), .Z(n13067) );
  NANDN U7449 ( .A(y[115]), .B(x[115]), .Z(n3991) );
  NANDN U7450 ( .A(y[114]), .B(x[114]), .Z(n3990) );
  AND U7451 ( .A(n3991), .B(n3990), .Z(n13064) );
  NANDN U7452 ( .A(x[113]), .B(y[113]), .Z(n3993) );
  NANDN U7453 ( .A(x[114]), .B(y[114]), .Z(n3992) );
  NAND U7454 ( .A(n3993), .B(n3992), .Z(n13063) );
  NANDN U7455 ( .A(x[111]), .B(y[111]), .Z(n3995) );
  NANDN U7456 ( .A(x[112]), .B(y[112]), .Z(n3994) );
  NAND U7457 ( .A(n3995), .B(n3994), .Z(n13058) );
  NANDN U7458 ( .A(x[109]), .B(y[109]), .Z(n3997) );
  NANDN U7459 ( .A(x[110]), .B(y[110]), .Z(n3996) );
  NAND U7460 ( .A(n3997), .B(n3996), .Z(n13055) );
  NANDN U7461 ( .A(y[109]), .B(x[109]), .Z(n3999) );
  NANDN U7462 ( .A(y[108]), .B(x[108]), .Z(n3998) );
  AND U7463 ( .A(n3999), .B(n3998), .Z(n13052) );
  NANDN U7464 ( .A(x[107]), .B(y[107]), .Z(n4001) );
  NANDN U7465 ( .A(x[108]), .B(y[108]), .Z(n4000) );
  NAND U7466 ( .A(n4001), .B(n4000), .Z(n13051) );
  NANDN U7467 ( .A(x[105]), .B(y[105]), .Z(n4003) );
  NANDN U7468 ( .A(x[106]), .B(y[106]), .Z(n4002) );
  NAND U7469 ( .A(n4003), .B(n4002), .Z(n13046) );
  NANDN U7470 ( .A(x[103]), .B(y[103]), .Z(n4005) );
  NANDN U7471 ( .A(x[104]), .B(y[104]), .Z(n4004) );
  NAND U7472 ( .A(n4005), .B(n4004), .Z(n13043) );
  NANDN U7473 ( .A(y[103]), .B(x[103]), .Z(n4007) );
  NANDN U7474 ( .A(y[102]), .B(x[102]), .Z(n4006) );
  AND U7475 ( .A(n4007), .B(n4006), .Z(n13040) );
  NANDN U7476 ( .A(x[101]), .B(y[101]), .Z(n4009) );
  NANDN U7477 ( .A(x[102]), .B(y[102]), .Z(n4008) );
  NAND U7478 ( .A(n4009), .B(n4008), .Z(n13039) );
  NANDN U7479 ( .A(x[99]), .B(y[99]), .Z(n4010) );
  NANDN U7480 ( .A(x[100]), .B(y[100]), .Z(n12778) );
  NAND U7481 ( .A(n4010), .B(n12778), .Z(n12781) );
  IV U7482 ( .A(x[96]), .Z(n13023) );
  NAND U7483 ( .A(n13023), .B(y[96]), .Z(n4256) );
  XOR U7484 ( .A(n13023), .B(y[96]), .Z(n4254) );
  ANDN U7485 ( .B(y[95]), .A(x[95]), .Z(n13022) );
  NANDN U7486 ( .A(y[95]), .B(x[95]), .Z(n4012) );
  NANDN U7487 ( .A(y[94]), .B(x[94]), .Z(n4011) );
  NAND U7488 ( .A(n4012), .B(n4011), .Z(n13020) );
  NANDN U7489 ( .A(x[94]), .B(y[94]), .Z(n4014) );
  NANDN U7490 ( .A(x[93]), .B(y[93]), .Z(n4013) );
  NAND U7491 ( .A(n4014), .B(n4013), .Z(n13018) );
  NANDN U7492 ( .A(y[92]), .B(x[92]), .Z(n4016) );
  NANDN U7493 ( .A(y[93]), .B(x[93]), .Z(n4015) );
  NAND U7494 ( .A(n4016), .B(n4015), .Z(n13016) );
  NANDN U7495 ( .A(y[90]), .B(x[90]), .Z(n4018) );
  NANDN U7496 ( .A(y[91]), .B(x[91]), .Z(n4017) );
  NAND U7497 ( .A(n4018), .B(n4017), .Z(n13012) );
  NANDN U7498 ( .A(x[90]), .B(y[90]), .Z(n4020) );
  NANDN U7499 ( .A(x[89]), .B(y[89]), .Z(n4019) );
  NAND U7500 ( .A(n4020), .B(n4019), .Z(n13009) );
  NANDN U7501 ( .A(y[88]), .B(x[88]), .Z(n4022) );
  NANDN U7502 ( .A(y[89]), .B(x[89]), .Z(n4021) );
  NAND U7503 ( .A(n4022), .B(n4021), .Z(n13008) );
  NANDN U7504 ( .A(x[88]), .B(y[88]), .Z(n4024) );
  NANDN U7505 ( .A(x[87]), .B(y[87]), .Z(n4023) );
  NAND U7506 ( .A(n4024), .B(n4023), .Z(n13006) );
  NANDN U7507 ( .A(y[86]), .B(x[86]), .Z(n4026) );
  NANDN U7508 ( .A(y[87]), .B(x[87]), .Z(n4025) );
  NAND U7509 ( .A(n4026), .B(n4025), .Z(n13004) );
  NANDN U7510 ( .A(y[84]), .B(x[84]), .Z(n4028) );
  NANDN U7511 ( .A(y[85]), .B(x[85]), .Z(n4027) );
  NAND U7512 ( .A(n4028), .B(n4027), .Z(n13000) );
  NANDN U7513 ( .A(x[84]), .B(y[84]), .Z(n4030) );
  NANDN U7514 ( .A(x[83]), .B(y[83]), .Z(n4029) );
  NAND U7515 ( .A(n4030), .B(n4029), .Z(n12997) );
  NANDN U7516 ( .A(y[82]), .B(x[82]), .Z(n4032) );
  NANDN U7517 ( .A(y[83]), .B(x[83]), .Z(n4031) );
  NAND U7518 ( .A(n4032), .B(n4031), .Z(n12996) );
  NANDN U7519 ( .A(x[82]), .B(y[82]), .Z(n4034) );
  NANDN U7520 ( .A(x[81]), .B(y[81]), .Z(n4033) );
  NAND U7521 ( .A(n4034), .B(n4033), .Z(n12994) );
  NANDN U7522 ( .A(y[80]), .B(x[80]), .Z(n4036) );
  NANDN U7523 ( .A(y[81]), .B(x[81]), .Z(n4035) );
  NAND U7524 ( .A(n4036), .B(n4035), .Z(n12992) );
  NANDN U7525 ( .A(y[78]), .B(x[78]), .Z(n4038) );
  NANDN U7526 ( .A(y[79]), .B(x[79]), .Z(n4037) );
  NAND U7527 ( .A(n4038), .B(n4037), .Z(n12988) );
  NANDN U7528 ( .A(x[78]), .B(y[78]), .Z(n4040) );
  NANDN U7529 ( .A(x[77]), .B(y[77]), .Z(n4039) );
  NAND U7530 ( .A(n4040), .B(n4039), .Z(n12985) );
  NANDN U7531 ( .A(y[76]), .B(x[76]), .Z(n4042) );
  NANDN U7532 ( .A(y[77]), .B(x[77]), .Z(n4041) );
  NAND U7533 ( .A(n4042), .B(n4041), .Z(n12984) );
  NANDN U7534 ( .A(x[76]), .B(y[76]), .Z(n4044) );
  NANDN U7535 ( .A(x[75]), .B(y[75]), .Z(n4043) );
  NAND U7536 ( .A(n4044), .B(n4043), .Z(n12982) );
  NANDN U7537 ( .A(y[74]), .B(x[74]), .Z(n4046) );
  NANDN U7538 ( .A(y[75]), .B(x[75]), .Z(n4045) );
  NAND U7539 ( .A(n4046), .B(n4045), .Z(n12980) );
  NANDN U7540 ( .A(y[72]), .B(x[72]), .Z(n4048) );
  NANDN U7541 ( .A(y[73]), .B(x[73]), .Z(n4047) );
  NAND U7542 ( .A(n4048), .B(n4047), .Z(n12976) );
  NANDN U7543 ( .A(x[72]), .B(y[72]), .Z(n4050) );
  NANDN U7544 ( .A(x[71]), .B(y[71]), .Z(n4049) );
  NAND U7545 ( .A(n4050), .B(n4049), .Z(n12973) );
  NANDN U7546 ( .A(y[70]), .B(x[70]), .Z(n4052) );
  NANDN U7547 ( .A(y[71]), .B(x[71]), .Z(n4051) );
  NAND U7548 ( .A(n4052), .B(n4051), .Z(n12972) );
  NANDN U7549 ( .A(x[70]), .B(y[70]), .Z(n4054) );
  NANDN U7550 ( .A(x[69]), .B(y[69]), .Z(n4053) );
  NAND U7551 ( .A(n4054), .B(n4053), .Z(n12970) );
  ANDN U7552 ( .B(y[67]), .A(x[67]), .Z(n12962) );
  NANDN U7553 ( .A(y[67]), .B(x[67]), .Z(n4056) );
  NANDN U7554 ( .A(y[66]), .B(x[66]), .Z(n4055) );
  NAND U7555 ( .A(n4056), .B(n4055), .Z(n12959) );
  NANDN U7556 ( .A(y[64]), .B(x[64]), .Z(n4058) );
  NANDN U7557 ( .A(y[65]), .B(x[65]), .Z(n4057) );
  NAND U7558 ( .A(n4058), .B(n4057), .Z(n12956) );
  NANDN U7559 ( .A(x[64]), .B(y[64]), .Z(n4060) );
  NANDN U7560 ( .A(x[63]), .B(y[63]), .Z(n4059) );
  NAND U7561 ( .A(n4060), .B(n4059), .Z(n12954) );
  NANDN U7562 ( .A(y[62]), .B(x[62]), .Z(n4062) );
  NANDN U7563 ( .A(y[63]), .B(x[63]), .Z(n4061) );
  NAND U7564 ( .A(n4062), .B(n4061), .Z(n12952) );
  NANDN U7565 ( .A(x[62]), .B(y[62]), .Z(n4064) );
  NANDN U7566 ( .A(x[61]), .B(y[61]), .Z(n4063) );
  NAND U7567 ( .A(n4064), .B(n4063), .Z(n12950) );
  NANDN U7568 ( .A(y[60]), .B(x[60]), .Z(n4066) );
  NANDN U7569 ( .A(y[61]), .B(x[61]), .Z(n4065) );
  NAND U7570 ( .A(n4066), .B(n4065), .Z(n12948) );
  NANDN U7571 ( .A(y[58]), .B(x[58]), .Z(n4068) );
  NANDN U7572 ( .A(y[59]), .B(x[59]), .Z(n4067) );
  NAND U7573 ( .A(n4068), .B(n4067), .Z(n12944) );
  ANDN U7574 ( .B(y[58]), .A(x[58]), .Z(n12942) );
  NANDN U7575 ( .A(y[55]), .B(x[55]), .Z(n4070) );
  NANDN U7576 ( .A(y[54]), .B(x[54]), .Z(n4069) );
  NAND U7577 ( .A(n4070), .B(n4069), .Z(n12929) );
  NANDN U7578 ( .A(x[54]), .B(y[54]), .Z(n4072) );
  NANDN U7579 ( .A(x[53]), .B(y[53]), .Z(n4071) );
  NAND U7580 ( .A(n4072), .B(n4071), .Z(n12927) );
  NANDN U7581 ( .A(y[52]), .B(x[52]), .Z(n4074) );
  NANDN U7582 ( .A(y[53]), .B(x[53]), .Z(n4073) );
  NAND U7583 ( .A(n4074), .B(n4073), .Z(n12925) );
  NANDN U7584 ( .A(x[52]), .B(y[52]), .Z(n4076) );
  NANDN U7585 ( .A(x[51]), .B(y[51]), .Z(n4075) );
  NAND U7586 ( .A(n4076), .B(n4075), .Z(n12923) );
  NANDN U7587 ( .A(y[50]), .B(x[50]), .Z(n4078) );
  NANDN U7588 ( .A(y[51]), .B(x[51]), .Z(n4077) );
  NAND U7589 ( .A(n4078), .B(n4077), .Z(n12921) );
  NANDN U7590 ( .A(y[48]), .B(x[48]), .Z(n4080) );
  NANDN U7591 ( .A(y[49]), .B(x[49]), .Z(n4079) );
  NAND U7592 ( .A(n4080), .B(n4079), .Z(n12917) );
  NANDN U7593 ( .A(x[48]), .B(y[48]), .Z(n4082) );
  NANDN U7594 ( .A(x[47]), .B(y[47]), .Z(n4081) );
  NAND U7595 ( .A(n4082), .B(n4081), .Z(n12915) );
  NANDN U7596 ( .A(y[46]), .B(x[46]), .Z(n4084) );
  NANDN U7597 ( .A(y[47]), .B(x[47]), .Z(n4083) );
  NAND U7598 ( .A(n4084), .B(n4083), .Z(n12913) );
  NANDN U7599 ( .A(x[46]), .B(y[46]), .Z(n4086) );
  NANDN U7600 ( .A(x[45]), .B(y[45]), .Z(n4085) );
  NAND U7601 ( .A(n4086), .B(n4085), .Z(n12911) );
  NANDN U7602 ( .A(y[44]), .B(x[44]), .Z(n4088) );
  NANDN U7603 ( .A(y[45]), .B(x[45]), .Z(n4087) );
  NAND U7604 ( .A(n4088), .B(n4087), .Z(n12909) );
  NANDN U7605 ( .A(y[42]), .B(x[42]), .Z(n4090) );
  NANDN U7606 ( .A(y[43]), .B(x[43]), .Z(n4089) );
  NAND U7607 ( .A(n4090), .B(n4089), .Z(n12905) );
  NANDN U7608 ( .A(x[42]), .B(y[42]), .Z(n4092) );
  NANDN U7609 ( .A(x[41]), .B(y[41]), .Z(n4091) );
  NAND U7610 ( .A(n4092), .B(n4091), .Z(n12903) );
  NANDN U7611 ( .A(y[40]), .B(x[40]), .Z(n4094) );
  NANDN U7612 ( .A(y[41]), .B(x[41]), .Z(n4093) );
  NAND U7613 ( .A(n4094), .B(n4093), .Z(n12901) );
  NANDN U7614 ( .A(x[40]), .B(y[40]), .Z(n4096) );
  NANDN U7615 ( .A(x[39]), .B(y[39]), .Z(n4095) );
  NAND U7616 ( .A(n4096), .B(n4095), .Z(n12899) );
  NANDN U7617 ( .A(y[38]), .B(x[38]), .Z(n4098) );
  NANDN U7618 ( .A(y[39]), .B(x[39]), .Z(n4097) );
  NAND U7619 ( .A(n4098), .B(n4097), .Z(n12897) );
  NANDN U7620 ( .A(y[36]), .B(x[36]), .Z(n4100) );
  NANDN U7621 ( .A(y[37]), .B(x[37]), .Z(n4099) );
  NAND U7622 ( .A(n4100), .B(n4099), .Z(n12893) );
  NANDN U7623 ( .A(x[36]), .B(y[36]), .Z(n4102) );
  NANDN U7624 ( .A(x[35]), .B(y[35]), .Z(n4101) );
  NAND U7625 ( .A(n4102), .B(n4101), .Z(n12891) );
  NANDN U7626 ( .A(y[34]), .B(x[34]), .Z(n4104) );
  NANDN U7627 ( .A(y[35]), .B(x[35]), .Z(n4103) );
  NAND U7628 ( .A(n4104), .B(n4103), .Z(n12889) );
  NANDN U7629 ( .A(x[34]), .B(y[34]), .Z(n4106) );
  NANDN U7630 ( .A(x[33]), .B(y[33]), .Z(n4105) );
  NAND U7631 ( .A(n4106), .B(n4105), .Z(n12887) );
  NANDN U7632 ( .A(y[32]), .B(x[32]), .Z(n4108) );
  NANDN U7633 ( .A(y[33]), .B(x[33]), .Z(n4107) );
  NAND U7634 ( .A(n4108), .B(n4107), .Z(n12885) );
  NANDN U7635 ( .A(y[30]), .B(x[30]), .Z(n4110) );
  NANDN U7636 ( .A(y[31]), .B(x[31]), .Z(n4109) );
  NAND U7637 ( .A(n4110), .B(n4109), .Z(n12881) );
  NANDN U7638 ( .A(x[30]), .B(y[30]), .Z(n4112) );
  NANDN U7639 ( .A(x[29]), .B(y[29]), .Z(n4111) );
  NAND U7640 ( .A(n4112), .B(n4111), .Z(n12879) );
  NANDN U7641 ( .A(y[28]), .B(x[28]), .Z(n4114) );
  NANDN U7642 ( .A(y[29]), .B(x[29]), .Z(n4113) );
  NAND U7643 ( .A(n4114), .B(n4113), .Z(n12877) );
  NANDN U7644 ( .A(x[28]), .B(y[28]), .Z(n4116) );
  NANDN U7645 ( .A(x[27]), .B(y[27]), .Z(n4115) );
  NAND U7646 ( .A(n4116), .B(n4115), .Z(n12875) );
  NANDN U7647 ( .A(y[26]), .B(x[26]), .Z(n4118) );
  NANDN U7648 ( .A(y[27]), .B(x[27]), .Z(n4117) );
  NAND U7649 ( .A(n4118), .B(n4117), .Z(n12873) );
  NANDN U7650 ( .A(y[24]), .B(x[24]), .Z(n4120) );
  NANDN U7651 ( .A(y[25]), .B(x[25]), .Z(n4119) );
  NAND U7652 ( .A(n4120), .B(n4119), .Z(n12869) );
  ANDN U7653 ( .B(y[24]), .A(x[24]), .Z(n12867) );
  NANDN U7654 ( .A(x[20]), .B(y[20]), .Z(n12786) );
  ANDN U7655 ( .B(y[19]), .A(x[19]), .Z(n12850) );
  ANDN U7656 ( .B(n12786), .A(n12850), .Z(n4159) );
  NANDN U7657 ( .A(y[19]), .B(x[19]), .Z(n4122) );
  NANDN U7658 ( .A(y[18]), .B(x[18]), .Z(n4121) );
  NAND U7659 ( .A(n4122), .B(n4121), .Z(n12847) );
  NANDN U7660 ( .A(x[16]), .B(y[16]), .Z(n12842) );
  NANDN U7661 ( .A(x[17]), .B(y[17]), .Z(n4123) );
  NANDN U7662 ( .A(x[18]), .B(y[18]), .Z(n4154) );
  NAND U7663 ( .A(n4123), .B(n4154), .Z(n12845) );
  ANDN U7664 ( .B(n12842), .A(n12845), .Z(n4153) );
  ANDN U7665 ( .B(x[16]), .A(y[16]), .Z(n12788) );
  NANDN U7666 ( .A(x[14]), .B(y[14]), .Z(n4125) );
  NANDN U7667 ( .A(x[15]), .B(y[15]), .Z(n4124) );
  NAND U7668 ( .A(n4125), .B(n4124), .Z(n12838) );
  ANDN U7669 ( .B(x[13]), .A(y[13]), .Z(n12832) );
  ANDN U7670 ( .B(y[13]), .A(x[13]), .Z(n12833) );
  NANDN U7671 ( .A(x[10]), .B(y[10]), .Z(n12821) );
  ANDN U7672 ( .B(y[11]), .A(x[11]), .Z(n12790) );
  ANDN U7673 ( .B(n12821), .A(n12790), .Z(n4142) );
  ANDN U7674 ( .B(x[9]), .A(y[9]), .Z(n12815) );
  ANDN U7675 ( .B(x[10]), .A(y[10]), .Z(n12826) );
  ANDN U7676 ( .B(y[8]), .A(x[8]), .Z(n12792) );
  ANDN U7677 ( .B(x[8]), .A(y[8]), .Z(n12818) );
  ANDN U7678 ( .B(y[6]), .A(x[6]), .Z(n12809) );
  NANDN U7679 ( .A(y[6]), .B(x[6]), .Z(n4127) );
  NANDN U7680 ( .A(y[5]), .B(x[5]), .Z(n4126) );
  NAND U7681 ( .A(n4127), .B(n4126), .Z(n12808) );
  NANDN U7682 ( .A(x[5]), .B(y[5]), .Z(n4129) );
  NANDN U7683 ( .A(x[4]), .B(y[4]), .Z(n4128) );
  NAND U7684 ( .A(n4129), .B(n4128), .Z(n12806) );
  NANDN U7685 ( .A(y[2]), .B(x[2]), .Z(n4131) );
  NANDN U7686 ( .A(y[1]), .B(x[1]), .Z(n4130) );
  NAND U7687 ( .A(n4131), .B(n4130), .Z(n12796) );
  NANDN U7688 ( .A(x[1]), .B(y[1]), .Z(n12793) );
  ANDN U7689 ( .B(y[2]), .A(x[2]), .Z(n12798) );
  NANDN U7690 ( .A(y[4]), .B(x[4]), .Z(n12800) );
  NANDN U7691 ( .A(n12808), .B(n4132), .Z(n4133) );
  ANDN U7692 ( .B(y[7]), .A(x[7]), .Z(n12791) );
  ANDN U7693 ( .B(n4133), .A(n12791), .Z(n4134) );
  NANDN U7694 ( .A(n12809), .B(n4134), .Z(n4135) );
  ANDN U7695 ( .B(x[7]), .A(y[7]), .Z(n12812) );
  ANDN U7696 ( .B(n4135), .A(n12812), .Z(n4136) );
  NANDN U7697 ( .A(n12818), .B(n4136), .Z(n4137) );
  ANDN U7698 ( .B(y[9]), .A(x[9]), .Z(n12819) );
  ANDN U7699 ( .B(n4137), .A(n12819), .Z(n4138) );
  NANDN U7700 ( .A(n12792), .B(n4138), .Z(n4139) );
  NANDN U7701 ( .A(n12826), .B(n4139), .Z(n4140) );
  OR U7702 ( .A(n12815), .B(n4140), .Z(n4141) );
  AND U7703 ( .A(n4142), .B(n4141), .Z(n4144) );
  NANDN U7704 ( .A(y[12]), .B(x[12]), .Z(n12829) );
  ANDN U7705 ( .B(x[11]), .A(y[11]), .Z(n12823) );
  ANDN U7706 ( .B(n12829), .A(n12823), .Z(n4143) );
  NANDN U7707 ( .A(n4144), .B(n4143), .Z(n4145) );
  ANDN U7708 ( .B(y[12]), .A(x[12]), .Z(n12789) );
  ANDN U7709 ( .B(n4145), .A(n12789), .Z(n4146) );
  NANDN U7710 ( .A(n12833), .B(n4146), .Z(n4147) );
  ANDN U7711 ( .B(x[14]), .A(y[14]), .Z(n12836) );
  ANDN U7712 ( .B(n4147), .A(n12836), .Z(n4148) );
  NANDN U7713 ( .A(n12832), .B(n4148), .Z(n4149) );
  NANDN U7714 ( .A(n12838), .B(n4149), .Z(n4150) );
  ANDN U7715 ( .B(x[15]), .A(y[15]), .Z(n12840) );
  ANDN U7716 ( .B(n4150), .A(n12840), .Z(n4151) );
  NANDN U7717 ( .A(n12788), .B(n4151), .Z(n4152) );
  NAND U7718 ( .A(n4153), .B(n4152), .Z(n4156) );
  ANDN U7719 ( .B(x[17]), .A(y[17]), .Z(n12787) );
  NAND U7720 ( .A(n4154), .B(n12787), .Z(n4155) );
  NAND U7721 ( .A(n4156), .B(n4155), .Z(n4157) );
  OR U7722 ( .A(n12847), .B(n4157), .Z(n4158) );
  AND U7723 ( .A(n4159), .B(n4158), .Z(n4161) );
  NANDN U7724 ( .A(y[21]), .B(x[21]), .Z(n12855) );
  ANDN U7725 ( .B(x[20]), .A(y[20]), .Z(n12852) );
  ANDN U7726 ( .B(n12855), .A(n12852), .Z(n4160) );
  NANDN U7727 ( .A(n4161), .B(n4160), .Z(n4162) );
  ANDN U7728 ( .B(y[21]), .A(x[21]), .Z(n12785) );
  ANDN U7729 ( .B(n4162), .A(n12785), .Z(n4163) );
  NAND U7730 ( .A(n4163), .B(n12861), .Z(n4166) );
  NANDN U7731 ( .A(y[23]), .B(x[23]), .Z(n12864) );
  IV U7732 ( .A(y[22]), .Z(n12857) );
  NAND U7733 ( .A(x[22]), .B(n12857), .Z(n4164) );
  AND U7734 ( .A(n12864), .B(n4164), .Z(n4165) );
  NAND U7735 ( .A(n4166), .B(n4165), .Z(n4167) );
  ANDN U7736 ( .B(y[23]), .A(x[23]), .Z(n12860) );
  ANDN U7737 ( .B(n4167), .A(n12860), .Z(n4168) );
  NANDN U7738 ( .A(n12867), .B(n4168), .Z(n4169) );
  NANDN U7739 ( .A(n12869), .B(n4169), .Z(n4172) );
  NANDN U7740 ( .A(x[26]), .B(y[26]), .Z(n4171) );
  NANDN U7741 ( .A(x[25]), .B(y[25]), .Z(n4170) );
  NAND U7742 ( .A(n4171), .B(n4170), .Z(n12870) );
  ANDN U7743 ( .B(n4172), .A(n12870), .Z(n4173) );
  OR U7744 ( .A(n12873), .B(n4173), .Z(n4174) );
  NANDN U7745 ( .A(n12875), .B(n4174), .Z(n4175) );
  NANDN U7746 ( .A(n12877), .B(n4175), .Z(n4176) );
  NANDN U7747 ( .A(n12879), .B(n4176), .Z(n4177) );
  NANDN U7748 ( .A(n12881), .B(n4177), .Z(n4180) );
  NANDN U7749 ( .A(x[32]), .B(y[32]), .Z(n4179) );
  NANDN U7750 ( .A(x[31]), .B(y[31]), .Z(n4178) );
  NAND U7751 ( .A(n4179), .B(n4178), .Z(n12882) );
  ANDN U7752 ( .B(n4180), .A(n12882), .Z(n4181) );
  OR U7753 ( .A(n12885), .B(n4181), .Z(n4182) );
  NANDN U7754 ( .A(n12887), .B(n4182), .Z(n4183) );
  NANDN U7755 ( .A(n12889), .B(n4183), .Z(n4184) );
  NANDN U7756 ( .A(n12891), .B(n4184), .Z(n4185) );
  NANDN U7757 ( .A(n12893), .B(n4185), .Z(n4188) );
  NANDN U7758 ( .A(x[38]), .B(y[38]), .Z(n4187) );
  NANDN U7759 ( .A(x[37]), .B(y[37]), .Z(n4186) );
  NAND U7760 ( .A(n4187), .B(n4186), .Z(n12894) );
  ANDN U7761 ( .B(n4188), .A(n12894), .Z(n4189) );
  OR U7762 ( .A(n12897), .B(n4189), .Z(n4190) );
  NANDN U7763 ( .A(n12899), .B(n4190), .Z(n4191) );
  NANDN U7764 ( .A(n12901), .B(n4191), .Z(n4192) );
  NANDN U7765 ( .A(n12903), .B(n4192), .Z(n4193) );
  NANDN U7766 ( .A(n12905), .B(n4193), .Z(n4196) );
  NANDN U7767 ( .A(x[44]), .B(y[44]), .Z(n4195) );
  NANDN U7768 ( .A(x[43]), .B(y[43]), .Z(n4194) );
  NAND U7769 ( .A(n4195), .B(n4194), .Z(n12906) );
  ANDN U7770 ( .B(n4196), .A(n12906), .Z(n4197) );
  OR U7771 ( .A(n12909), .B(n4197), .Z(n4198) );
  NANDN U7772 ( .A(n12911), .B(n4198), .Z(n4199) );
  NANDN U7773 ( .A(n12913), .B(n4199), .Z(n4200) );
  NANDN U7774 ( .A(n12915), .B(n4200), .Z(n4201) );
  NANDN U7775 ( .A(n12917), .B(n4201), .Z(n4204) );
  NANDN U7776 ( .A(x[50]), .B(y[50]), .Z(n4203) );
  NANDN U7777 ( .A(x[49]), .B(y[49]), .Z(n4202) );
  NAND U7778 ( .A(n4203), .B(n4202), .Z(n12918) );
  ANDN U7779 ( .B(n4204), .A(n12918), .Z(n4205) );
  OR U7780 ( .A(n12921), .B(n4205), .Z(n4206) );
  NANDN U7781 ( .A(n12923), .B(n4206), .Z(n4207) );
  NANDN U7782 ( .A(n12925), .B(n4207), .Z(n4208) );
  NANDN U7783 ( .A(n12927), .B(n4208), .Z(n4209) );
  NANDN U7784 ( .A(n12929), .B(n4209), .Z(n4210) );
  ANDN U7785 ( .B(y[55]), .A(x[55]), .Z(n12930) );
  ANDN U7786 ( .B(n4210), .A(n12930), .Z(n4211) );
  NAND U7787 ( .A(n4211), .B(n12936), .Z(n4214) );
  NANDN U7788 ( .A(y[57]), .B(x[57]), .Z(n12939) );
  IV U7789 ( .A(y[56]), .Z(n12932) );
  NAND U7790 ( .A(x[56]), .B(n12932), .Z(n4212) );
  AND U7791 ( .A(n12939), .B(n4212), .Z(n4213) );
  NAND U7792 ( .A(n4214), .B(n4213), .Z(n4215) );
  ANDN U7793 ( .B(y[57]), .A(x[57]), .Z(n12935) );
  ANDN U7794 ( .B(n4215), .A(n12935), .Z(n4216) );
  NANDN U7795 ( .A(n12942), .B(n4216), .Z(n4217) );
  NANDN U7796 ( .A(n12944), .B(n4217), .Z(n4220) );
  NANDN U7797 ( .A(x[60]), .B(y[60]), .Z(n4219) );
  NANDN U7798 ( .A(x[59]), .B(y[59]), .Z(n4218) );
  NAND U7799 ( .A(n4219), .B(n4218), .Z(n12945) );
  ANDN U7800 ( .B(n4220), .A(n12945), .Z(n4221) );
  OR U7801 ( .A(n12948), .B(n4221), .Z(n4222) );
  NANDN U7802 ( .A(n12950), .B(n4222), .Z(n4223) );
  NANDN U7803 ( .A(n12952), .B(n4223), .Z(n4224) );
  NANDN U7804 ( .A(n12954), .B(n4224), .Z(n4225) );
  NANDN U7805 ( .A(n12956), .B(n4225), .Z(n4228) );
  NANDN U7806 ( .A(x[66]), .B(y[66]), .Z(n4227) );
  NANDN U7807 ( .A(x[65]), .B(y[65]), .Z(n4226) );
  NAND U7808 ( .A(n4227), .B(n4226), .Z(n12957) );
  NANDN U7809 ( .A(y[69]), .B(x[69]), .Z(n12964) );
  NANDN U7810 ( .A(x[74]), .B(y[74]), .Z(n4230) );
  NANDN U7811 ( .A(x[73]), .B(y[73]), .Z(n4229) );
  NAND U7812 ( .A(n4230), .B(n4229), .Z(n12978) );
  NANDN U7813 ( .A(x[80]), .B(y[80]), .Z(n4232) );
  NANDN U7814 ( .A(x[79]), .B(y[79]), .Z(n4231) );
  NAND U7815 ( .A(n4232), .B(n4231), .Z(n12990) );
  OR U7816 ( .A(n12992), .B(n4233), .Z(n4234) );
  NANDN U7817 ( .A(n12994), .B(n4234), .Z(n4235) );
  NANDN U7818 ( .A(n12996), .B(n4235), .Z(n4236) );
  NANDN U7819 ( .A(n12997), .B(n4236), .Z(n4237) );
  NANDN U7820 ( .A(n13000), .B(n4237), .Z(n4240) );
  NANDN U7821 ( .A(x[86]), .B(y[86]), .Z(n4239) );
  NANDN U7822 ( .A(x[85]), .B(y[85]), .Z(n4238) );
  NAND U7823 ( .A(n4239), .B(n4238), .Z(n13002) );
  ANDN U7824 ( .B(n4240), .A(n13002), .Z(n4241) );
  OR U7825 ( .A(n13004), .B(n4241), .Z(n4242) );
  NANDN U7826 ( .A(n13006), .B(n4242), .Z(n4243) );
  NANDN U7827 ( .A(n13008), .B(n4243), .Z(n4244) );
  NANDN U7828 ( .A(n13009), .B(n4244), .Z(n4245) );
  NANDN U7829 ( .A(n13012), .B(n4245), .Z(n4248) );
  NANDN U7830 ( .A(x[92]), .B(y[92]), .Z(n4247) );
  NANDN U7831 ( .A(x[91]), .B(y[91]), .Z(n4246) );
  NAND U7832 ( .A(n4247), .B(n4246), .Z(n13014) );
  ANDN U7833 ( .B(n4248), .A(n13014), .Z(n4249) );
  OR U7834 ( .A(n13016), .B(n4249), .Z(n4250) );
  NANDN U7835 ( .A(n13018), .B(n4250), .Z(n4251) );
  NANDN U7836 ( .A(n13020), .B(n4251), .Z(n4252) );
  NANDN U7837 ( .A(n13022), .B(n4252), .Z(n4253) );
  NAND U7838 ( .A(n4254), .B(n4253), .Z(n4255) );
  AND U7839 ( .A(n4256), .B(n4255), .Z(n4257) );
  XNOR U7840 ( .A(n4257), .B(y[97]), .Z(n4258) );
  NANDN U7841 ( .A(x[97]), .B(n4258), .Z(n4259) );
  IV U7842 ( .A(x[98]), .Z(n12780) );
  NANDN U7843 ( .A(y[98]), .B(x[98]), .Z(n12784) );
  ANDN U7844 ( .B(x[99]), .A(y[99]), .Z(n12779) );
  NANDN U7845 ( .A(y[101]), .B(x[101]), .Z(n4261) );
  NANDN U7846 ( .A(y[100]), .B(x[100]), .Z(n4260) );
  AND U7847 ( .A(n4261), .B(n4260), .Z(n13036) );
  NANDN U7848 ( .A(y[105]), .B(x[105]), .Z(n4263) );
  NANDN U7849 ( .A(y[104]), .B(x[104]), .Z(n4262) );
  AND U7850 ( .A(n4263), .B(n4262), .Z(n13044) );
  NANDN U7851 ( .A(y[107]), .B(x[107]), .Z(n4265) );
  NANDN U7852 ( .A(y[106]), .B(x[106]), .Z(n4264) );
  AND U7853 ( .A(n4265), .B(n4264), .Z(n13048) );
  NANDN U7854 ( .A(y[111]), .B(x[111]), .Z(n4267) );
  NANDN U7855 ( .A(y[110]), .B(x[110]), .Z(n4266) );
  AND U7856 ( .A(n4267), .B(n4266), .Z(n13056) );
  NANDN U7857 ( .A(y[113]), .B(x[113]), .Z(n4269) );
  NANDN U7858 ( .A(y[112]), .B(x[112]), .Z(n4268) );
  AND U7859 ( .A(n4269), .B(n4268), .Z(n13060) );
  NAND U7860 ( .A(n4270), .B(n13060), .Z(n4271) );
  NANDN U7861 ( .A(n13063), .B(n4271), .Z(n4272) );
  AND U7862 ( .A(n13064), .B(n4272), .Z(n4273) );
  OR U7863 ( .A(n13067), .B(n4273), .Z(n4276) );
  NANDN U7864 ( .A(y[117]), .B(x[117]), .Z(n4275) );
  NANDN U7865 ( .A(y[116]), .B(x[116]), .Z(n4274) );
  AND U7866 ( .A(n4275), .B(n4274), .Z(n13068) );
  NAND U7867 ( .A(n4276), .B(n13068), .Z(n4277) );
  NANDN U7868 ( .A(n13070), .B(n4277), .Z(n4280) );
  NANDN U7869 ( .A(y[119]), .B(x[119]), .Z(n4279) );
  NANDN U7870 ( .A(y[118]), .B(x[118]), .Z(n4278) );
  AND U7871 ( .A(n4279), .B(n4278), .Z(n13072) );
  NAND U7872 ( .A(n4280), .B(n13072), .Z(n4281) );
  NANDN U7873 ( .A(n13075), .B(n4281), .Z(n4282) );
  AND U7874 ( .A(n13076), .B(n4282), .Z(n4283) );
  OR U7875 ( .A(n13079), .B(n4283), .Z(n4286) );
  NANDN U7876 ( .A(y[123]), .B(x[123]), .Z(n4285) );
  NANDN U7877 ( .A(y[122]), .B(x[122]), .Z(n4284) );
  AND U7878 ( .A(n4285), .B(n4284), .Z(n13080) );
  NAND U7879 ( .A(n4286), .B(n13080), .Z(n4287) );
  NANDN U7880 ( .A(n13082), .B(n4287), .Z(n4290) );
  NANDN U7881 ( .A(y[125]), .B(x[125]), .Z(n4289) );
  NANDN U7882 ( .A(y[124]), .B(x[124]), .Z(n4288) );
  AND U7883 ( .A(n4289), .B(n4288), .Z(n13084) );
  NAND U7884 ( .A(n4290), .B(n13084), .Z(n4291) );
  NANDN U7885 ( .A(n13087), .B(n4291), .Z(n4292) );
  AND U7886 ( .A(n13088), .B(n4292), .Z(n4293) );
  OR U7887 ( .A(n13091), .B(n4293), .Z(n4296) );
  NANDN U7888 ( .A(y[129]), .B(x[129]), .Z(n4295) );
  NANDN U7889 ( .A(y[128]), .B(x[128]), .Z(n4294) );
  AND U7890 ( .A(n4295), .B(n4294), .Z(n13092) );
  NAND U7891 ( .A(n4296), .B(n13092), .Z(n4297) );
  NANDN U7892 ( .A(n13094), .B(n4297), .Z(n4300) );
  NANDN U7893 ( .A(y[131]), .B(x[131]), .Z(n4299) );
  NANDN U7894 ( .A(y[130]), .B(x[130]), .Z(n4298) );
  AND U7895 ( .A(n4299), .B(n4298), .Z(n13096) );
  NAND U7896 ( .A(n4300), .B(n13096), .Z(n4301) );
  NANDN U7897 ( .A(n13099), .B(n4301), .Z(n4302) );
  AND U7898 ( .A(n13100), .B(n4302), .Z(n4303) );
  OR U7899 ( .A(n13103), .B(n4303), .Z(n4306) );
  NANDN U7900 ( .A(y[135]), .B(x[135]), .Z(n4305) );
  NANDN U7901 ( .A(y[134]), .B(x[134]), .Z(n4304) );
  AND U7902 ( .A(n4305), .B(n4304), .Z(n13104) );
  NAND U7903 ( .A(n4306), .B(n13104), .Z(n4307) );
  NANDN U7904 ( .A(n13106), .B(n4307), .Z(n4310) );
  NANDN U7905 ( .A(y[137]), .B(x[137]), .Z(n4309) );
  NANDN U7906 ( .A(y[136]), .B(x[136]), .Z(n4308) );
  AND U7907 ( .A(n4309), .B(n4308), .Z(n13108) );
  NAND U7908 ( .A(n4310), .B(n13108), .Z(n4311) );
  NANDN U7909 ( .A(n13111), .B(n4311), .Z(n4312) );
  AND U7910 ( .A(n13112), .B(n4312), .Z(n4313) );
  OR U7911 ( .A(n13115), .B(n4313), .Z(n4316) );
  NANDN U7912 ( .A(y[141]), .B(x[141]), .Z(n4315) );
  NANDN U7913 ( .A(y[140]), .B(x[140]), .Z(n4314) );
  AND U7914 ( .A(n4315), .B(n4314), .Z(n13116) );
  NAND U7915 ( .A(n4316), .B(n13116), .Z(n4317) );
  NANDN U7916 ( .A(n13118), .B(n4317), .Z(n4320) );
  NANDN U7917 ( .A(y[143]), .B(x[143]), .Z(n4319) );
  NANDN U7918 ( .A(y[142]), .B(x[142]), .Z(n4318) );
  AND U7919 ( .A(n4319), .B(n4318), .Z(n13120) );
  NAND U7920 ( .A(n4320), .B(n13120), .Z(n4321) );
  NANDN U7921 ( .A(n13123), .B(n4321), .Z(n4322) );
  AND U7922 ( .A(n13124), .B(n4322), .Z(n4323) );
  OR U7923 ( .A(n13127), .B(n4323), .Z(n4326) );
  NANDN U7924 ( .A(y[147]), .B(x[147]), .Z(n4325) );
  NANDN U7925 ( .A(y[146]), .B(x[146]), .Z(n4324) );
  AND U7926 ( .A(n4325), .B(n4324), .Z(n13128) );
  NAND U7927 ( .A(n4326), .B(n13128), .Z(n4327) );
  NANDN U7928 ( .A(n13130), .B(n4327), .Z(n4330) );
  NANDN U7929 ( .A(y[149]), .B(x[149]), .Z(n4329) );
  NANDN U7930 ( .A(y[148]), .B(x[148]), .Z(n4328) );
  AND U7931 ( .A(n4329), .B(n4328), .Z(n13132) );
  NAND U7932 ( .A(n4330), .B(n13132), .Z(n4331) );
  NANDN U7933 ( .A(n13135), .B(n4331), .Z(n4332) );
  AND U7934 ( .A(n13136), .B(n4332), .Z(n4333) );
  OR U7935 ( .A(n13139), .B(n4333), .Z(n4336) );
  NANDN U7936 ( .A(y[153]), .B(x[153]), .Z(n4335) );
  NANDN U7937 ( .A(y[152]), .B(x[152]), .Z(n4334) );
  AND U7938 ( .A(n4335), .B(n4334), .Z(n13140) );
  NAND U7939 ( .A(n4336), .B(n13140), .Z(n4337) );
  NANDN U7940 ( .A(n13142), .B(n4337), .Z(n4340) );
  NANDN U7941 ( .A(y[155]), .B(x[155]), .Z(n4339) );
  NANDN U7942 ( .A(y[154]), .B(x[154]), .Z(n4338) );
  AND U7943 ( .A(n4339), .B(n4338), .Z(n13144) );
  NAND U7944 ( .A(n4340), .B(n13144), .Z(n4341) );
  NANDN U7945 ( .A(n13147), .B(n4341), .Z(n4342) );
  AND U7946 ( .A(n13148), .B(n4342), .Z(n4343) );
  OR U7947 ( .A(n13151), .B(n4343), .Z(n4346) );
  NANDN U7948 ( .A(y[158]), .B(x[158]), .Z(n4345) );
  NANDN U7949 ( .A(y[159]), .B(x[159]), .Z(n4344) );
  AND U7950 ( .A(n4345), .B(n4344), .Z(n13152) );
  NAND U7951 ( .A(n4346), .B(n13152), .Z(n4347) );
  NANDN U7952 ( .A(n4348), .B(n4347), .Z(n4349) );
  OR U7953 ( .A(n13155), .B(n4349), .Z(n4352) );
  NANDN U7954 ( .A(y[161]), .B(x[161]), .Z(n13157) );
  NANDN U7955 ( .A(y[160]), .B(x[160]), .Z(n4350) );
  AND U7956 ( .A(n13157), .B(n4350), .Z(n4351) );
  NAND U7957 ( .A(n4352), .B(n4351), .Z(n4353) );
  NANDN U7958 ( .A(n13163), .B(n4353), .Z(n4356) );
  NANDN U7959 ( .A(y[163]), .B(x[163]), .Z(n4355) );
  NANDN U7960 ( .A(y[162]), .B(x[162]), .Z(n4354) );
  AND U7961 ( .A(n4355), .B(n4354), .Z(n13164) );
  NAND U7962 ( .A(n4356), .B(n13164), .Z(n4357) );
  NANDN U7963 ( .A(n13166), .B(n4357), .Z(n4358) );
  AND U7964 ( .A(n13168), .B(n4358), .Z(n4359) );
  OR U7965 ( .A(n13171), .B(n4359), .Z(n4362) );
  NANDN U7966 ( .A(y[167]), .B(x[167]), .Z(n4361) );
  NANDN U7967 ( .A(y[166]), .B(x[166]), .Z(n4360) );
  AND U7968 ( .A(n4361), .B(n4360), .Z(n13172) );
  NAND U7969 ( .A(n4362), .B(n13172), .Z(n4363) );
  NANDN U7970 ( .A(n13175), .B(n4363), .Z(n4368) );
  XNOR U7971 ( .A(x[169]), .B(y[169]), .Z(n4365) );
  NANDN U7972 ( .A(y[168]), .B(x[168]), .Z(n4364) );
  NAND U7973 ( .A(n4365), .B(n4364), .Z(n4366) );
  NAND U7974 ( .A(n4367), .B(n4366), .Z(n13176) );
  NAND U7975 ( .A(n4368), .B(n13176), .Z(n4369) );
  NANDN U7976 ( .A(n13178), .B(n4369), .Z(n4370) );
  AND U7977 ( .A(n13180), .B(n4370), .Z(n4371) );
  OR U7978 ( .A(n13183), .B(n4371), .Z(n4374) );
  NANDN U7979 ( .A(y[173]), .B(x[173]), .Z(n4373) );
  NANDN U7980 ( .A(y[172]), .B(x[172]), .Z(n4372) );
  AND U7981 ( .A(n4373), .B(n4372), .Z(n13184) );
  NAND U7982 ( .A(n4374), .B(n13184), .Z(n4375) );
  NANDN U7983 ( .A(n13187), .B(n4375), .Z(n4378) );
  NANDN U7984 ( .A(y[175]), .B(x[175]), .Z(n4377) );
  NANDN U7985 ( .A(y[174]), .B(x[174]), .Z(n4376) );
  AND U7986 ( .A(n4377), .B(n4376), .Z(n13188) );
  NAND U7987 ( .A(n4378), .B(n13188), .Z(n4379) );
  NANDN U7988 ( .A(n13190), .B(n4379), .Z(n4380) );
  AND U7989 ( .A(n13192), .B(n4380), .Z(n4381) );
  OR U7990 ( .A(n13195), .B(n4381), .Z(n4382) );
  NANDN U7991 ( .A(y[179]), .B(x[179]), .Z(n13196) );
  NAND U7992 ( .A(n4382), .B(n13196), .Z(n4383) );
  NANDN U7993 ( .A(n13199), .B(n4383), .Z(n4386) );
  NANDN U7994 ( .A(y[181]), .B(x[181]), .Z(n4385) );
  NANDN U7995 ( .A(y[180]), .B(x[180]), .Z(n4384) );
  AND U7996 ( .A(n4385), .B(n4384), .Z(n13200) );
  NAND U7997 ( .A(n4386), .B(n13200), .Z(n4387) );
  NANDN U7998 ( .A(n13202), .B(n4387), .Z(n4388) );
  AND U7999 ( .A(n13204), .B(n4388), .Z(n4389) );
  OR U8000 ( .A(n13207), .B(n4389), .Z(n4392) );
  NANDN U8001 ( .A(y[184]), .B(x[184]), .Z(n4391) );
  NANDN U8002 ( .A(y[185]), .B(x[185]), .Z(n4390) );
  AND U8003 ( .A(n4391), .B(n4390), .Z(n13208) );
  NAND U8004 ( .A(n4392), .B(n13208), .Z(n4393) );
  NANDN U8005 ( .A(n4394), .B(n4393), .Z(n4395) );
  OR U8006 ( .A(n13211), .B(n4395), .Z(n4398) );
  NANDN U8007 ( .A(y[186]), .B(x[186]), .Z(n4396) );
  ANDN U8008 ( .B(x[187]), .A(y[187]), .Z(n13217) );
  ANDN U8009 ( .B(n4396), .A(n13217), .Z(n4397) );
  NAND U8010 ( .A(n4398), .B(n4397), .Z(n4399) );
  NANDN U8011 ( .A(n13220), .B(n4399), .Z(n4400) );
  NANDN U8012 ( .A(n13222), .B(n4400), .Z(n4401) );
  NANDN U8013 ( .A(n13224), .B(n4401), .Z(n4404) );
  NANDN U8014 ( .A(y[191]), .B(x[191]), .Z(n4403) );
  NANDN U8015 ( .A(y[190]), .B(x[190]), .Z(n4402) );
  NAND U8016 ( .A(n4403), .B(n4402), .Z(n13226) );
  ANDN U8017 ( .B(n4404), .A(n13226), .Z(n4405) );
  OR U8018 ( .A(n13228), .B(n4405), .Z(n4406) );
  NANDN U8019 ( .A(n13229), .B(n4406), .Z(n4407) );
  NANDN U8020 ( .A(n13232), .B(n4407), .Z(n4408) );
  NANDN U8021 ( .A(n13234), .B(n4408), .Z(n4409) );
  NANDN U8022 ( .A(n13236), .B(n4409), .Z(n4418) );
  NANDN U8023 ( .A(y[199]), .B(x[199]), .Z(n4415) );
  ANDN U8024 ( .B(x[196]), .A(y[196]), .Z(n4410) );
  OR U8025 ( .A(n4410), .B(x[197]), .Z(n4413) );
  XOR U8026 ( .A(x[197]), .B(n4410), .Z(n4411) );
  NAND U8027 ( .A(n4411), .B(y[197]), .Z(n4412) );
  NAND U8028 ( .A(n4413), .B(n4412), .Z(n4414) );
  AND U8029 ( .A(n4415), .B(n4414), .Z(n4417) );
  NANDN U8030 ( .A(y[198]), .B(x[198]), .Z(n4416) );
  NAND U8031 ( .A(n4417), .B(n4416), .Z(n13238) );
  ANDN U8032 ( .B(n4418), .A(n13238), .Z(n4419) );
  OR U8033 ( .A(n13240), .B(n4419), .Z(n4420) );
  NANDN U8034 ( .A(n13241), .B(n4420), .Z(n4421) );
  NANDN U8035 ( .A(n13244), .B(n4421), .Z(n4422) );
  NANDN U8036 ( .A(n13246), .B(n4422), .Z(n4423) );
  NANDN U8037 ( .A(n13248), .B(n4423), .Z(n4433) );
  NANDN U8038 ( .A(y[204]), .B(x[204]), .Z(n4425) );
  NAND U8039 ( .A(n4424), .B(n4425), .Z(n4428) );
  XNOR U8040 ( .A(n4425), .B(x[205]), .Z(n4426) );
  NAND U8041 ( .A(n4426), .B(y[205]), .Z(n4427) );
  NAND U8042 ( .A(n4428), .B(n4427), .Z(n4430) );
  ANDN U8043 ( .B(n4430), .A(n4429), .Z(n4432) );
  NANDN U8044 ( .A(y[206]), .B(x[206]), .Z(n4431) );
  NAND U8045 ( .A(n4432), .B(n4431), .Z(n12776) );
  ANDN U8046 ( .B(n4433), .A(n12776), .Z(n4434) );
  NANDN U8047 ( .A(n12774), .B(n4434), .Z(n4435) );
  NANDN U8048 ( .A(n13252), .B(n4435), .Z(n4438) );
  NANDN U8049 ( .A(y[211]), .B(x[211]), .Z(n4437) );
  NANDN U8050 ( .A(y[210]), .B(x[210]), .Z(n4436) );
  NAND U8051 ( .A(n4437), .B(n4436), .Z(n13254) );
  ANDN U8052 ( .B(n4438), .A(n13254), .Z(n4439) );
  ANDN U8053 ( .B(y[215]), .A(x[215]), .Z(n13263) );
  NANDN U8054 ( .A(y[219]), .B(x[219]), .Z(n4441) );
  NANDN U8055 ( .A(y[218]), .B(x[218]), .Z(n4440) );
  NAND U8056 ( .A(n4441), .B(n4440), .Z(n13274) );
  ANDN U8057 ( .B(y[225]), .A(x[225]), .Z(n13285) );
  IV U8058 ( .A(x[226]), .Z(n13291) );
  NAND U8059 ( .A(n13291), .B(y[226]), .Z(n4442) );
  NAND U8060 ( .A(n4443), .B(n4442), .Z(n4446) );
  NANDN U8061 ( .A(y[226]), .B(x[226]), .Z(n4444) );
  ANDN U8062 ( .B(x[227]), .A(y[227]), .Z(n13296) );
  ANDN U8063 ( .B(n4444), .A(n13296), .Z(n4445) );
  NAND U8064 ( .A(n4446), .B(n4445), .Z(n4447) );
  AND U8065 ( .A(n13298), .B(n4447), .Z(n4448) );
  OR U8066 ( .A(n13301), .B(n4448), .Z(n4451) );
  NANDN U8067 ( .A(x[230]), .B(y[230]), .Z(n4450) );
  NANDN U8068 ( .A(x[229]), .B(y[229]), .Z(n4449) );
  AND U8069 ( .A(n4450), .B(n4449), .Z(n13302) );
  NAND U8070 ( .A(n4451), .B(n13302), .Z(n4452) );
  NANDN U8071 ( .A(n13305), .B(n4452), .Z(n4455) );
  NANDN U8072 ( .A(x[232]), .B(y[232]), .Z(n4454) );
  NANDN U8073 ( .A(x[231]), .B(y[231]), .Z(n4453) );
  AND U8074 ( .A(n4454), .B(n4453), .Z(n13306) );
  NAND U8075 ( .A(n4455), .B(n13306), .Z(n4456) );
  NANDN U8076 ( .A(n13308), .B(n4456), .Z(n4457) );
  AND U8077 ( .A(n13310), .B(n4457), .Z(n4458) );
  OR U8078 ( .A(n13313), .B(n4458), .Z(n4461) );
  NANDN U8079 ( .A(x[236]), .B(y[236]), .Z(n4460) );
  NANDN U8080 ( .A(x[235]), .B(y[235]), .Z(n4459) );
  AND U8081 ( .A(n4460), .B(n4459), .Z(n13314) );
  NAND U8082 ( .A(n4461), .B(n13314), .Z(n4462) );
  NANDN U8083 ( .A(n13317), .B(n4462), .Z(n4465) );
  NANDN U8084 ( .A(x[238]), .B(y[238]), .Z(n4464) );
  NANDN U8085 ( .A(x[237]), .B(y[237]), .Z(n4463) );
  AND U8086 ( .A(n4464), .B(n4463), .Z(n13318) );
  NAND U8087 ( .A(n4465), .B(n13318), .Z(n4466) );
  NANDN U8088 ( .A(n13320), .B(n4466), .Z(n4467) );
  AND U8089 ( .A(n13322), .B(n4467), .Z(n4468) );
  OR U8090 ( .A(n13325), .B(n4468), .Z(n4471) );
  NANDN U8091 ( .A(x[242]), .B(y[242]), .Z(n4470) );
  NANDN U8092 ( .A(x[241]), .B(y[241]), .Z(n4469) );
  AND U8093 ( .A(n4470), .B(n4469), .Z(n13326) );
  NAND U8094 ( .A(n4471), .B(n13326), .Z(n4472) );
  NANDN U8095 ( .A(n13329), .B(n4472), .Z(n4478) );
  NANDN U8096 ( .A(x[244]), .B(y[244]), .Z(n4474) );
  NANDN U8097 ( .A(x[243]), .B(y[243]), .Z(n4473) );
  AND U8098 ( .A(n4474), .B(n4473), .Z(n4477) );
  NAND U8099 ( .A(n4475), .B(y[245]), .Z(n4476) );
  AND U8100 ( .A(n4477), .B(n4476), .Z(n13330) );
  NAND U8101 ( .A(n4478), .B(n13330), .Z(n4479) );
  NANDN U8102 ( .A(n13332), .B(n4479), .Z(n4480) );
  AND U8103 ( .A(n13334), .B(n4480), .Z(n4481) );
  OR U8104 ( .A(n13337), .B(n4481), .Z(n4484) );
  NANDN U8105 ( .A(x[250]), .B(y[250]), .Z(n4483) );
  NANDN U8106 ( .A(x[249]), .B(y[249]), .Z(n4482) );
  AND U8107 ( .A(n4483), .B(n4482), .Z(n13338) );
  NAND U8108 ( .A(n4484), .B(n13338), .Z(n4485) );
  NANDN U8109 ( .A(n13341), .B(n4485), .Z(n4488) );
  NANDN U8110 ( .A(x[252]), .B(y[252]), .Z(n4487) );
  NANDN U8111 ( .A(x[251]), .B(y[251]), .Z(n4486) );
  AND U8112 ( .A(n4487), .B(n4486), .Z(n13342) );
  NAND U8113 ( .A(n4488), .B(n13342), .Z(n4489) );
  NANDN U8114 ( .A(n13344), .B(n4489), .Z(n4490) );
  AND U8115 ( .A(n13346), .B(n4490), .Z(n4491) );
  OR U8116 ( .A(n13349), .B(n4491), .Z(n4494) );
  NANDN U8117 ( .A(x[256]), .B(y[256]), .Z(n4493) );
  NANDN U8118 ( .A(x[255]), .B(y[255]), .Z(n4492) );
  AND U8119 ( .A(n4493), .B(n4492), .Z(n13350) );
  NAND U8120 ( .A(n4494), .B(n13350), .Z(n4495) );
  NANDN U8121 ( .A(n13353), .B(n4495), .Z(n4498) );
  NANDN U8122 ( .A(x[258]), .B(y[258]), .Z(n4497) );
  NANDN U8123 ( .A(x[257]), .B(y[257]), .Z(n4496) );
  AND U8124 ( .A(n4497), .B(n4496), .Z(n13354) );
  NAND U8125 ( .A(n4498), .B(n13354), .Z(n4499) );
  NANDN U8126 ( .A(n13356), .B(n4499), .Z(n4500) );
  AND U8127 ( .A(n13358), .B(n4500), .Z(n4501) );
  OR U8128 ( .A(n13361), .B(n4501), .Z(n4506) );
  NANDN U8129 ( .A(x[263]), .B(y[263]), .Z(n4503) );
  NANDN U8130 ( .A(x[262]), .B(y[262]), .Z(n4502) );
  AND U8131 ( .A(n4503), .B(n4502), .Z(n4505) );
  NANDN U8132 ( .A(x[264]), .B(y[264]), .Z(n4504) );
  AND U8133 ( .A(n4505), .B(n4504), .Z(n13362) );
  NAND U8134 ( .A(n4506), .B(n13362), .Z(n4507) );
  NANDN U8135 ( .A(n13365), .B(n4507), .Z(n4510) );
  NANDN U8136 ( .A(x[266]), .B(y[266]), .Z(n4509) );
  NANDN U8137 ( .A(x[265]), .B(y[265]), .Z(n4508) );
  AND U8138 ( .A(n4509), .B(n4508), .Z(n13366) );
  NAND U8139 ( .A(n4510), .B(n13366), .Z(n4511) );
  NANDN U8140 ( .A(n13368), .B(n4511), .Z(n4512) );
  AND U8141 ( .A(n13370), .B(n4512), .Z(n4513) );
  OR U8142 ( .A(n13373), .B(n4513), .Z(n4514) );
  AND U8143 ( .A(n4515), .B(n4514), .Z(n4518) );
  NANDN U8144 ( .A(y[270]), .B(x[270]), .Z(n4516) );
  ANDN U8145 ( .B(x[271]), .A(y[271]), .Z(n13380) );
  ANDN U8146 ( .B(n4516), .A(n13380), .Z(n4517) );
  NANDN U8147 ( .A(n4518), .B(n4517), .Z(n4524) );
  NANDN U8148 ( .A(x[272]), .B(y[272]), .Z(n4520) );
  NANDN U8149 ( .A(x[271]), .B(y[271]), .Z(n4519) );
  AND U8150 ( .A(n4520), .B(n4519), .Z(n4523) );
  NAND U8151 ( .A(n4521), .B(y[273]), .Z(n4522) );
  AND U8152 ( .A(n4523), .B(n4522), .Z(n13382) );
  NAND U8153 ( .A(n4524), .B(n13382), .Z(n4525) );
  NANDN U8154 ( .A(n13385), .B(n4525), .Z(n4526) );
  NANDN U8155 ( .A(x[274]), .B(y[274]), .Z(n13386) );
  NAND U8156 ( .A(n4526), .B(n13386), .Z(n4527) );
  NANDN U8157 ( .A(n13389), .B(n4527), .Z(n4528) );
  AND U8158 ( .A(n13390), .B(n4528), .Z(n4529) );
  OR U8159 ( .A(n13392), .B(n4529), .Z(n4532) );
  NANDN U8160 ( .A(x[278]), .B(y[278]), .Z(n4531) );
  NANDN U8161 ( .A(x[277]), .B(y[277]), .Z(n4530) );
  AND U8162 ( .A(n4531), .B(n4530), .Z(n13394) );
  NAND U8163 ( .A(n4532), .B(n13394), .Z(n4533) );
  NANDN U8164 ( .A(n13397), .B(n4533), .Z(n4536) );
  NANDN U8165 ( .A(x[280]), .B(y[280]), .Z(n4535) );
  NANDN U8166 ( .A(x[279]), .B(y[279]), .Z(n4534) );
  AND U8167 ( .A(n4535), .B(n4534), .Z(n13398) );
  NAND U8168 ( .A(n4536), .B(n13398), .Z(n4537) );
  NANDN U8169 ( .A(n13401), .B(n4537), .Z(n4538) );
  AND U8170 ( .A(n13402), .B(n4538), .Z(n4539) );
  OR U8171 ( .A(n13404), .B(n4539), .Z(n4545) );
  NANDN U8172 ( .A(x[284]), .B(y[284]), .Z(n4541) );
  NANDN U8173 ( .A(x[283]), .B(y[283]), .Z(n4540) );
  AND U8174 ( .A(n4541), .B(n4540), .Z(n4544) );
  NAND U8175 ( .A(n4542), .B(y[285]), .Z(n4543) );
  AND U8176 ( .A(n4544), .B(n4543), .Z(n13406) );
  NAND U8177 ( .A(n4545), .B(n13406), .Z(n4546) );
  NANDN U8178 ( .A(n13408), .B(n4546), .Z(n4548) );
  NAND U8179 ( .A(n4548), .B(n20307), .Z(n4549) );
  NANDN U8180 ( .A(n20309), .B(n4549), .Z(n4550) );
  AND U8181 ( .A(n20313), .B(n4550), .Z(n4551) );
  OR U8182 ( .A(n13416), .B(n4551), .Z(n4552) );
  NANDN U8183 ( .A(n20317), .B(n4552), .Z(n4555) );
  NANDN U8184 ( .A(y[292]), .B(x[292]), .Z(n4554) );
  NANDN U8185 ( .A(y[293]), .B(x[293]), .Z(n4553) );
  AND U8186 ( .A(n4554), .B(n4553), .Z(n20319) );
  NAND U8187 ( .A(n4555), .B(n20319), .Z(n4556) );
  NANDN U8188 ( .A(n20322), .B(n4556), .Z(n4559) );
  NANDN U8189 ( .A(y[294]), .B(x[294]), .Z(n4558) );
  NANDN U8190 ( .A(y[295]), .B(x[295]), .Z(n4557) );
  AND U8191 ( .A(n4558), .B(n4557), .Z(n20323) );
  NAND U8192 ( .A(n4559), .B(n20323), .Z(n4562) );
  NANDN U8193 ( .A(x[296]), .B(y[296]), .Z(n4561) );
  NANDN U8194 ( .A(x[295]), .B(y[295]), .Z(n4560) );
  NAND U8195 ( .A(n4561), .B(n4560), .Z(n20326) );
  ANDN U8196 ( .B(n4562), .A(n20326), .Z(n4565) );
  NANDN U8197 ( .A(y[296]), .B(x[296]), .Z(n4564) );
  NANDN U8198 ( .A(y[297]), .B(x[297]), .Z(n4563) );
  AND U8199 ( .A(n4564), .B(n4563), .Z(n20327) );
  NANDN U8200 ( .A(n4565), .B(n20327), .Z(n4566) );
  NANDN U8201 ( .A(n20329), .B(n4566), .Z(n4569) );
  NANDN U8202 ( .A(y[298]), .B(x[298]), .Z(n4568) );
  NANDN U8203 ( .A(y[299]), .B(x[299]), .Z(n4567) );
  AND U8204 ( .A(n4568), .B(n4567), .Z(n20331) );
  NAND U8205 ( .A(n4569), .B(n20331), .Z(n4570) );
  NANDN U8206 ( .A(n20334), .B(n4570), .Z(n4573) );
  NANDN U8207 ( .A(y[300]), .B(x[300]), .Z(n4572) );
  NANDN U8208 ( .A(y[301]), .B(x[301]), .Z(n4571) );
  AND U8209 ( .A(n4572), .B(n4571), .Z(n20335) );
  NAND U8210 ( .A(n4573), .B(n20335), .Z(n4576) );
  NANDN U8211 ( .A(x[302]), .B(y[302]), .Z(n4575) );
  NANDN U8212 ( .A(x[301]), .B(y[301]), .Z(n4574) );
  NAND U8213 ( .A(n4575), .B(n4574), .Z(n20338) );
  ANDN U8214 ( .B(n4576), .A(n20338), .Z(n4579) );
  NANDN U8215 ( .A(y[302]), .B(x[302]), .Z(n4578) );
  NANDN U8216 ( .A(y[303]), .B(x[303]), .Z(n4577) );
  AND U8217 ( .A(n4578), .B(n4577), .Z(n20339) );
  NANDN U8218 ( .A(n4579), .B(n20339), .Z(n4580) );
  NANDN U8219 ( .A(n20341), .B(n4580), .Z(n4583) );
  NANDN U8220 ( .A(y[304]), .B(x[304]), .Z(n4582) );
  NANDN U8221 ( .A(y[305]), .B(x[305]), .Z(n4581) );
  AND U8222 ( .A(n4582), .B(n4581), .Z(n20343) );
  NAND U8223 ( .A(n4583), .B(n20343), .Z(n4584) );
  NANDN U8224 ( .A(n20346), .B(n4584), .Z(n4587) );
  NANDN U8225 ( .A(y[306]), .B(x[306]), .Z(n4586) );
  NANDN U8226 ( .A(y[307]), .B(x[307]), .Z(n4585) );
  AND U8227 ( .A(n4586), .B(n4585), .Z(n20347) );
  NAND U8228 ( .A(n4587), .B(n20347), .Z(n4590) );
  NANDN U8229 ( .A(x[308]), .B(y[308]), .Z(n4589) );
  NANDN U8230 ( .A(x[307]), .B(y[307]), .Z(n4588) );
  NAND U8231 ( .A(n4589), .B(n4588), .Z(n20350) );
  ANDN U8232 ( .B(n4590), .A(n20350), .Z(n4593) );
  NANDN U8233 ( .A(y[308]), .B(x[308]), .Z(n4592) );
  NANDN U8234 ( .A(y[309]), .B(x[309]), .Z(n4591) );
  AND U8235 ( .A(n4592), .B(n4591), .Z(n20351) );
  NANDN U8236 ( .A(n4593), .B(n20351), .Z(n4594) );
  NANDN U8237 ( .A(n20353), .B(n4594), .Z(n4597) );
  NANDN U8238 ( .A(y[311]), .B(x[311]), .Z(n4596) );
  NANDN U8239 ( .A(y[310]), .B(x[310]), .Z(n4595) );
  AND U8240 ( .A(n4596), .B(n4595), .Z(n20355) );
  NAND U8241 ( .A(n4597), .B(n20355), .Z(n4600) );
  ANDN U8242 ( .B(y[311]), .A(x[311]), .Z(n20357) );
  NANDN U8243 ( .A(x[312]), .B(y[312]), .Z(n4599) );
  NAND U8244 ( .A(n4599), .B(n4598), .Z(n20362) );
  NOR U8245 ( .A(n20357), .B(n20362), .Z(n13437) );
  NAND U8246 ( .A(n4600), .B(n13437), .Z(n4601) );
  NANDN U8247 ( .A(n13439), .B(n4601), .Z(n4602) );
  NANDN U8248 ( .A(x[314]), .B(y[314]), .Z(n20365) );
  NAND U8249 ( .A(n4602), .B(n20365), .Z(n4605) );
  NANDN U8250 ( .A(y[315]), .B(x[315]), .Z(n4604) );
  NANDN U8251 ( .A(y[314]), .B(x[314]), .Z(n4603) );
  AND U8252 ( .A(n4604), .B(n4603), .Z(n20367) );
  NAND U8253 ( .A(n4605), .B(n20367), .Z(n4608) );
  NANDN U8254 ( .A(x[315]), .B(y[315]), .Z(n4607) );
  NANDN U8255 ( .A(x[316]), .B(y[316]), .Z(n4606) );
  AND U8256 ( .A(n4607), .B(n4606), .Z(n20370) );
  NAND U8257 ( .A(n4608), .B(n20370), .Z(n4609) );
  AND U8258 ( .A(n20371), .B(n4609), .Z(n4612) );
  NANDN U8259 ( .A(x[317]), .B(y[317]), .Z(n4611) );
  NANDN U8260 ( .A(x[318]), .B(y[318]), .Z(n4610) );
  AND U8261 ( .A(n4611), .B(n4610), .Z(n20373) );
  NANDN U8262 ( .A(n4612), .B(n20373), .Z(n4615) );
  NANDN U8263 ( .A(y[319]), .B(x[319]), .Z(n4614) );
  NANDN U8264 ( .A(y[318]), .B(x[318]), .Z(n4613) );
  AND U8265 ( .A(n4614), .B(n4613), .Z(n20375) );
  NAND U8266 ( .A(n4615), .B(n20375), .Z(n4618) );
  NANDN U8267 ( .A(x[319]), .B(y[319]), .Z(n4617) );
  NANDN U8268 ( .A(x[320]), .B(y[320]), .Z(n4616) );
  AND U8269 ( .A(n4617), .B(n4616), .Z(n20377) );
  NAND U8270 ( .A(n4618), .B(n20377), .Z(n4621) );
  NANDN U8271 ( .A(y[321]), .B(x[321]), .Z(n4620) );
  NANDN U8272 ( .A(y[320]), .B(x[320]), .Z(n4619) );
  AND U8273 ( .A(n4620), .B(n4619), .Z(n20379) );
  NAND U8274 ( .A(n4621), .B(n20379), .Z(n4622) );
  NANDN U8275 ( .A(x[321]), .B(y[321]), .Z(n20383) );
  NAND U8276 ( .A(n4622), .B(n20383), .Z(n4624) );
  NANDN U8277 ( .A(y[323]), .B(x[323]), .Z(n4627) );
  NANDN U8278 ( .A(y[322]), .B(x[322]), .Z(n4623) );
  NAND U8279 ( .A(n4627), .B(n4623), .Z(n20386) );
  ANDN U8280 ( .B(n4624), .A(n20386), .Z(n4629) );
  NANDN U8281 ( .A(x[324]), .B(y[324]), .Z(n4626) );
  NANDN U8282 ( .A(x[323]), .B(y[323]), .Z(n4625) );
  NAND U8283 ( .A(n4626), .B(n4625), .Z(n20387) );
  NANDN U8284 ( .A(x[322]), .B(y[322]), .Z(n20382) );
  NANDN U8285 ( .A(n20382), .B(n4627), .Z(n4628) );
  NANDN U8286 ( .A(n20387), .B(n4628), .Z(n13452) );
  OR U8287 ( .A(n4629), .B(n13452), .Z(n4630) );
  NANDN U8288 ( .A(n20390), .B(n4630), .Z(n4633) );
  NANDN U8289 ( .A(x[326]), .B(y[326]), .Z(n4632) );
  NANDN U8290 ( .A(x[325]), .B(y[325]), .Z(n4631) );
  AND U8291 ( .A(n4632), .B(n4631), .Z(n20391) );
  NAND U8292 ( .A(n4633), .B(n20391), .Z(n4634) );
  NANDN U8293 ( .A(n13456), .B(n4634), .Z(n4635) );
  ANDN U8294 ( .B(y[328]), .A(x[328]), .Z(n12773) );
  ANDN U8295 ( .B(n4635), .A(n12773), .Z(n4636) );
  NANDN U8296 ( .A(x[327]), .B(y[327]), .Z(n20395) );
  NAND U8297 ( .A(n4636), .B(n20395), .Z(n4637) );
  NAND U8298 ( .A(n4638), .B(n4637), .Z(n4639) );
  ANDN U8299 ( .B(y[329]), .A(x[329]), .Z(n12772) );
  ANDN U8300 ( .B(n4639), .A(n12772), .Z(n4640) );
  NANDN U8301 ( .A(n20404), .B(n4640), .Z(n4641) );
  NANDN U8302 ( .A(n13463), .B(n4641), .Z(n4642) );
  AND U8303 ( .A(n20407), .B(n4642), .Z(n4645) );
  NANDN U8304 ( .A(y[332]), .B(x[332]), .Z(n4644) );
  NANDN U8305 ( .A(y[333]), .B(x[333]), .Z(n4643) );
  AND U8306 ( .A(n4644), .B(n4643), .Z(n20409) );
  NANDN U8307 ( .A(n4645), .B(n20409), .Z(n4650) );
  NANDN U8308 ( .A(x[334]), .B(y[334]), .Z(n4647) );
  NANDN U8309 ( .A(x[333]), .B(y[333]), .Z(n4646) );
  AND U8310 ( .A(n4647), .B(n4646), .Z(n4649) );
  IV U8311 ( .A(x[335]), .Z(n4651) );
  NAND U8312 ( .A(n4651), .B(y[335]), .Z(n4648) );
  AND U8313 ( .A(n4649), .B(n4648), .Z(n20411) );
  NAND U8314 ( .A(n4650), .B(n20411), .Z(n4656) );
  NANDN U8315 ( .A(y[334]), .B(x[334]), .Z(n4652) );
  NANDN U8316 ( .A(n4652), .B(x[335]), .Z(n4655) );
  XOR U8317 ( .A(n4652), .B(n4651), .Z(n4653) );
  NANDN U8318 ( .A(y[335]), .B(n4653), .Z(n4654) );
  AND U8319 ( .A(n4655), .B(n4654), .Z(n20414) );
  NAND U8320 ( .A(n4656), .B(n20414), .Z(n4657) );
  NANDN U8321 ( .A(x[336]), .B(y[336]), .Z(n20415) );
  NAND U8322 ( .A(n4657), .B(n20415), .Z(n4660) );
  NANDN U8323 ( .A(y[336]), .B(x[336]), .Z(n4659) );
  NANDN U8324 ( .A(y[337]), .B(x[337]), .Z(n4658) );
  AND U8325 ( .A(n4659), .B(n4658), .Z(n20417) );
  NAND U8326 ( .A(n4660), .B(n20417), .Z(n4661) );
  AND U8327 ( .A(n20419), .B(n4661), .Z(n4666) );
  NANDN U8328 ( .A(y[338]), .B(x[338]), .Z(n4662) );
  NANDN U8329 ( .A(n4662), .B(x[339]), .Z(n4665) );
  XNOR U8330 ( .A(n4662), .B(x[339]), .Z(n4663) );
  NANDN U8331 ( .A(y[339]), .B(n4663), .Z(n4664) );
  AND U8332 ( .A(n4665), .B(n4664), .Z(n20421) );
  NANDN U8333 ( .A(n4666), .B(n20421), .Z(n4667) );
  NANDN U8334 ( .A(x[340]), .B(y[340]), .Z(n20423) );
  NAND U8335 ( .A(n4667), .B(n20423), .Z(n4670) );
  NANDN U8336 ( .A(y[340]), .B(x[340]), .Z(n4669) );
  NANDN U8337 ( .A(y[341]), .B(x[341]), .Z(n4668) );
  AND U8338 ( .A(n4669), .B(n4668), .Z(n20426) );
  NAND U8339 ( .A(n4670), .B(n20426), .Z(n4673) );
  NANDN U8340 ( .A(x[342]), .B(y[342]), .Z(n4672) );
  NANDN U8341 ( .A(x[341]), .B(y[341]), .Z(n4671) );
  AND U8342 ( .A(n4672), .B(n4671), .Z(n20427) );
  NAND U8343 ( .A(n4673), .B(n20427), .Z(n4676) );
  NANDN U8344 ( .A(y[342]), .B(x[342]), .Z(n4675) );
  NANDN U8345 ( .A(y[343]), .B(x[343]), .Z(n4674) );
  AND U8346 ( .A(n4675), .B(n4674), .Z(n20429) );
  NAND U8347 ( .A(n4676), .B(n20429), .Z(n4677) );
  AND U8348 ( .A(n20431), .B(n4677), .Z(n4680) );
  NANDN U8349 ( .A(y[344]), .B(x[344]), .Z(n4679) );
  NANDN U8350 ( .A(y[345]), .B(x[345]), .Z(n4678) );
  AND U8351 ( .A(n4679), .B(n4678), .Z(n20433) );
  NANDN U8352 ( .A(n4680), .B(n20433), .Z(n4683) );
  NANDN U8353 ( .A(x[346]), .B(y[346]), .Z(n4682) );
  NANDN U8354 ( .A(x[345]), .B(y[345]), .Z(n4681) );
  AND U8355 ( .A(n4682), .B(n4681), .Z(n20435) );
  NAND U8356 ( .A(n4683), .B(n20435), .Z(n4686) );
  NANDN U8357 ( .A(y[346]), .B(x[346]), .Z(n4685) );
  NANDN U8358 ( .A(y[347]), .B(x[347]), .Z(n4684) );
  AND U8359 ( .A(n4685), .B(n4684), .Z(n20438) );
  NAND U8360 ( .A(n4686), .B(n20438), .Z(n4689) );
  NANDN U8361 ( .A(x[348]), .B(y[348]), .Z(n4688) );
  NANDN U8362 ( .A(x[347]), .B(y[347]), .Z(n4687) );
  AND U8363 ( .A(n4688), .B(n4687), .Z(n20439) );
  NAND U8364 ( .A(n4689), .B(n20439), .Z(n4692) );
  NANDN U8365 ( .A(y[348]), .B(x[348]), .Z(n4691) );
  NANDN U8366 ( .A(y[349]), .B(x[349]), .Z(n4690) );
  AND U8367 ( .A(n4691), .B(n4690), .Z(n20441) );
  NAND U8368 ( .A(n4692), .B(n20441), .Z(n4693) );
  AND U8369 ( .A(n20443), .B(n4693), .Z(n4696) );
  NANDN U8370 ( .A(y[351]), .B(x[351]), .Z(n4695) );
  NANDN U8371 ( .A(y[350]), .B(x[350]), .Z(n4694) );
  AND U8372 ( .A(n4695), .B(n4694), .Z(n20445) );
  NANDN U8373 ( .A(n4696), .B(n20445), .Z(n4697) );
  AND U8374 ( .A(n4698), .B(n4697), .Z(n4700) );
  NANDN U8375 ( .A(y[352]), .B(x[352]), .Z(n4699) );
  ANDN U8376 ( .B(x[353]), .A(y[353]), .Z(n13487) );
  ANDN U8377 ( .B(n4699), .A(n13487), .Z(n20450) );
  NANDN U8378 ( .A(n4700), .B(n20450), .Z(n4701) );
  NANDN U8379 ( .A(n13489), .B(n4701), .Z(n4704) );
  NANDN U8380 ( .A(y[354]), .B(x[354]), .Z(n4703) );
  NANDN U8381 ( .A(y[355]), .B(x[355]), .Z(n4702) );
  AND U8382 ( .A(n4703), .B(n4702), .Z(n20453) );
  NAND U8383 ( .A(n4704), .B(n20453), .Z(n4707) );
  NANDN U8384 ( .A(x[356]), .B(y[356]), .Z(n4706) );
  NANDN U8385 ( .A(x[355]), .B(y[355]), .Z(n4705) );
  AND U8386 ( .A(n4706), .B(n4705), .Z(n20455) );
  NAND U8387 ( .A(n4707), .B(n20455), .Z(n4710) );
  NANDN U8388 ( .A(y[356]), .B(x[356]), .Z(n4709) );
  NANDN U8389 ( .A(y[357]), .B(x[357]), .Z(n4708) );
  AND U8390 ( .A(n4709), .B(n4708), .Z(n20457) );
  NAND U8391 ( .A(n4710), .B(n20457), .Z(n4711) );
  AND U8392 ( .A(n20459), .B(n4711), .Z(n4714) );
  NANDN U8393 ( .A(y[358]), .B(x[358]), .Z(n4713) );
  NANDN U8394 ( .A(y[359]), .B(x[359]), .Z(n4712) );
  AND U8395 ( .A(n4713), .B(n4712), .Z(n20462) );
  NANDN U8396 ( .A(n4714), .B(n20462), .Z(n4717) );
  NANDN U8397 ( .A(x[360]), .B(y[360]), .Z(n4716) );
  NANDN U8398 ( .A(x[359]), .B(y[359]), .Z(n4715) );
  AND U8399 ( .A(n4716), .B(n4715), .Z(n20463) );
  NAND U8400 ( .A(n4717), .B(n20463), .Z(n4720) );
  NANDN U8401 ( .A(y[360]), .B(x[360]), .Z(n4719) );
  NANDN U8402 ( .A(y[361]), .B(x[361]), .Z(n4718) );
  AND U8403 ( .A(n4719), .B(n4718), .Z(n20466) );
  NAND U8404 ( .A(n4720), .B(n20466), .Z(n4723) );
  NANDN U8405 ( .A(x[362]), .B(y[362]), .Z(n4722) );
  NANDN U8406 ( .A(x[361]), .B(y[361]), .Z(n4721) );
  AND U8407 ( .A(n4722), .B(n4721), .Z(n20467) );
  NAND U8408 ( .A(n4723), .B(n20467), .Z(n4726) );
  NANDN U8409 ( .A(y[363]), .B(x[363]), .Z(n4725) );
  NANDN U8410 ( .A(y[362]), .B(x[362]), .Z(n4724) );
  AND U8411 ( .A(n4725), .B(n4724), .Z(n20469) );
  NAND U8412 ( .A(n4726), .B(n20469), .Z(n4729) );
  NANDN U8413 ( .A(x[364]), .B(y[364]), .Z(n4727) );
  NANDN U8414 ( .A(n4728), .B(n4727), .Z(n20476) );
  NANDN U8415 ( .A(x[363]), .B(y[363]), .Z(n20471) );
  NANDN U8416 ( .A(n20476), .B(n20471), .Z(n13501) );
  ANDN U8417 ( .B(n4729), .A(n13501), .Z(n4730) );
  OR U8418 ( .A(n13502), .B(n4730), .Z(n4731) );
  NANDN U8419 ( .A(x[366]), .B(y[366]), .Z(n20479) );
  NAND U8420 ( .A(n4731), .B(n20479), .Z(n4734) );
  NANDN U8421 ( .A(y[366]), .B(x[366]), .Z(n4733) );
  NANDN U8422 ( .A(y[367]), .B(x[367]), .Z(n4732) );
  AND U8423 ( .A(n4733), .B(n4732), .Z(n20481) );
  NAND U8424 ( .A(n4734), .B(n20481), .Z(n4739) );
  NANDN U8425 ( .A(x[368]), .B(y[368]), .Z(n4736) );
  NANDN U8426 ( .A(x[367]), .B(y[367]), .Z(n4735) );
  AND U8427 ( .A(n4736), .B(n4735), .Z(n4738) );
  NANDN U8428 ( .A(x[369]), .B(y[369]), .Z(n4737) );
  AND U8429 ( .A(n4738), .B(n4737), .Z(n20483) );
  NAND U8430 ( .A(n4739), .B(n20483), .Z(n4740) );
  NANDN U8431 ( .A(n20486), .B(n4740), .Z(n4741) );
  AND U8432 ( .A(n20487), .B(n4741), .Z(n4744) );
  NANDN U8433 ( .A(y[372]), .B(x[372]), .Z(n4743) );
  NANDN U8434 ( .A(y[373]), .B(x[373]), .Z(n4742) );
  AND U8435 ( .A(n4743), .B(n4742), .Z(n20490) );
  NANDN U8436 ( .A(n4744), .B(n20490), .Z(n4747) );
  NANDN U8437 ( .A(x[374]), .B(y[374]), .Z(n4746) );
  NANDN U8438 ( .A(x[373]), .B(y[373]), .Z(n4745) );
  AND U8439 ( .A(n4746), .B(n4745), .Z(n20491) );
  NAND U8440 ( .A(n4747), .B(n20491), .Z(n4750) );
  NANDN U8441 ( .A(y[375]), .B(x[375]), .Z(n4749) );
  NANDN U8442 ( .A(y[374]), .B(x[374]), .Z(n4748) );
  AND U8443 ( .A(n4749), .B(n4748), .Z(n20493) );
  NAND U8444 ( .A(n4750), .B(n20493), .Z(n4751) );
  NAND U8445 ( .A(n20495), .B(n4751), .Z(n4753) );
  IV U8446 ( .A(x[376]), .Z(n12765) );
  AND U8447 ( .A(y[376]), .B(n12765), .Z(n4752) );
  OR U8448 ( .A(n4753), .B(n4752), .Z(n4754) );
  NANDN U8449 ( .A(n20498), .B(n4754), .Z(n4755) );
  NANDN U8450 ( .A(n12766), .B(n4755), .Z(n4756) );
  OR U8451 ( .A(n12771), .B(n4756), .Z(n4759) );
  NANDN U8452 ( .A(y[378]), .B(x[378]), .Z(n4758) );
  NANDN U8453 ( .A(y[379]), .B(x[379]), .Z(n4757) );
  AND U8454 ( .A(n4758), .B(n4757), .Z(n20502) );
  NAND U8455 ( .A(n4759), .B(n20502), .Z(n4760) );
  AND U8456 ( .A(n20503), .B(n4760), .Z(n4765) );
  NANDN U8457 ( .A(y[380]), .B(x[380]), .Z(n4761) );
  NANDN U8458 ( .A(n4761), .B(x[381]), .Z(n4764) );
  XNOR U8459 ( .A(n4761), .B(x[381]), .Z(n4762) );
  NANDN U8460 ( .A(y[381]), .B(n4762), .Z(n4763) );
  AND U8461 ( .A(n4764), .B(n4763), .Z(n20505) );
  NANDN U8462 ( .A(n4765), .B(n20505), .Z(n4766) );
  NANDN U8463 ( .A(x[382]), .B(y[382]), .Z(n20507) );
  NAND U8464 ( .A(n4766), .B(n20507), .Z(n4769) );
  NANDN U8465 ( .A(y[382]), .B(x[382]), .Z(n4768) );
  NANDN U8466 ( .A(y[383]), .B(x[383]), .Z(n4767) );
  AND U8467 ( .A(n4768), .B(n4767), .Z(n20509) );
  NAND U8468 ( .A(n4769), .B(n20509), .Z(n4772) );
  NANDN U8469 ( .A(x[384]), .B(y[384]), .Z(n4771) );
  NANDN U8470 ( .A(x[383]), .B(y[383]), .Z(n4770) );
  AND U8471 ( .A(n4771), .B(n4770), .Z(n20511) );
  NAND U8472 ( .A(n4772), .B(n20511), .Z(n4775) );
  NANDN U8473 ( .A(y[384]), .B(x[384]), .Z(n4774) );
  NANDN U8474 ( .A(y[385]), .B(x[385]), .Z(n4773) );
  AND U8475 ( .A(n4774), .B(n4773), .Z(n20514) );
  NAND U8476 ( .A(n4775), .B(n20514), .Z(n4776) );
  AND U8477 ( .A(n20515), .B(n4776), .Z(n4779) );
  NANDN U8478 ( .A(y[386]), .B(x[386]), .Z(n4778) );
  NANDN U8479 ( .A(y[387]), .B(x[387]), .Z(n4777) );
  AND U8480 ( .A(n4778), .B(n4777), .Z(n20517) );
  NANDN U8481 ( .A(n4779), .B(n20517), .Z(n4782) );
  NANDN U8482 ( .A(x[388]), .B(y[388]), .Z(n4781) );
  NANDN U8483 ( .A(x[387]), .B(y[387]), .Z(n4780) );
  AND U8484 ( .A(n4781), .B(n4780), .Z(n20519) );
  NAND U8485 ( .A(n4782), .B(n20519), .Z(n4785) );
  NANDN U8486 ( .A(y[388]), .B(x[388]), .Z(n4784) );
  NANDN U8487 ( .A(y[389]), .B(x[389]), .Z(n4783) );
  AND U8488 ( .A(n4784), .B(n4783), .Z(n20521) );
  NAND U8489 ( .A(n4785), .B(n20521), .Z(n4788) );
  NANDN U8490 ( .A(x[390]), .B(y[390]), .Z(n4787) );
  NANDN U8491 ( .A(x[389]), .B(y[389]), .Z(n4786) );
  AND U8492 ( .A(n4787), .B(n4786), .Z(n20523) );
  NAND U8493 ( .A(n4788), .B(n20523), .Z(n4791) );
  NANDN U8494 ( .A(y[390]), .B(x[390]), .Z(n4790) );
  NANDN U8495 ( .A(y[391]), .B(x[391]), .Z(n4789) );
  AND U8496 ( .A(n4790), .B(n4789), .Z(n20526) );
  NAND U8497 ( .A(n4791), .B(n20526), .Z(n4792) );
  AND U8498 ( .A(n20527), .B(n4792), .Z(n4795) );
  NANDN U8499 ( .A(y[392]), .B(x[392]), .Z(n4794) );
  NANDN U8500 ( .A(y[393]), .B(x[393]), .Z(n4793) );
  AND U8501 ( .A(n4794), .B(n4793), .Z(n20529) );
  NANDN U8502 ( .A(n4795), .B(n20529), .Z(n4800) );
  NANDN U8503 ( .A(x[394]), .B(y[394]), .Z(n4797) );
  NANDN U8504 ( .A(x[393]), .B(y[393]), .Z(n4796) );
  AND U8505 ( .A(n4797), .B(n4796), .Z(n4799) );
  IV U8506 ( .A(x[395]), .Z(n4801) );
  NAND U8507 ( .A(n4801), .B(y[395]), .Z(n4798) );
  AND U8508 ( .A(n4799), .B(n4798), .Z(n20531) );
  NAND U8509 ( .A(n4800), .B(n20531), .Z(n4806) );
  NANDN U8510 ( .A(y[394]), .B(x[394]), .Z(n4802) );
  NANDN U8511 ( .A(n4802), .B(x[395]), .Z(n4805) );
  XOR U8512 ( .A(n4802), .B(n4801), .Z(n4803) );
  NANDN U8513 ( .A(y[395]), .B(n4803), .Z(n4804) );
  AND U8514 ( .A(n4805), .B(n4804), .Z(n20533) );
  NAND U8515 ( .A(n4806), .B(n20533), .Z(n4807) );
  NANDN U8516 ( .A(x[396]), .B(y[396]), .Z(n20535) );
  NAND U8517 ( .A(n4807), .B(n20535), .Z(n4810) );
  NANDN U8518 ( .A(y[396]), .B(x[396]), .Z(n4809) );
  NANDN U8519 ( .A(y[397]), .B(x[397]), .Z(n4808) );
  AND U8520 ( .A(n4809), .B(n4808), .Z(n20538) );
  NAND U8521 ( .A(n4810), .B(n20538), .Z(n4811) );
  AND U8522 ( .A(n20539), .B(n4811), .Z(n4814) );
  NANDN U8523 ( .A(y[398]), .B(x[398]), .Z(n4813) );
  NANDN U8524 ( .A(y[399]), .B(x[399]), .Z(n4812) );
  AND U8525 ( .A(n4813), .B(n4812), .Z(n20541) );
  NANDN U8526 ( .A(n4814), .B(n20541), .Z(n4817) );
  NANDN U8527 ( .A(x[400]), .B(y[400]), .Z(n4816) );
  NANDN U8528 ( .A(x[399]), .B(y[399]), .Z(n4815) );
  AND U8529 ( .A(n4816), .B(n4815), .Z(n20543) );
  NAND U8530 ( .A(n4817), .B(n20543), .Z(n4820) );
  NANDN U8531 ( .A(y[400]), .B(x[400]), .Z(n4819) );
  NANDN U8532 ( .A(y[401]), .B(x[401]), .Z(n4818) );
  AND U8533 ( .A(n4819), .B(n4818), .Z(n20545) );
  NAND U8534 ( .A(n4820), .B(n20545), .Z(n4823) );
  NANDN U8535 ( .A(x[402]), .B(y[402]), .Z(n4822) );
  NANDN U8536 ( .A(x[401]), .B(y[401]), .Z(n4821) );
  AND U8537 ( .A(n4822), .B(n4821), .Z(n20547) );
  NAND U8538 ( .A(n4823), .B(n20547), .Z(n4826) );
  NANDN U8539 ( .A(y[402]), .B(x[402]), .Z(n4825) );
  NANDN U8540 ( .A(y[403]), .B(x[403]), .Z(n4824) );
  AND U8541 ( .A(n4825), .B(n4824), .Z(n20550) );
  NAND U8542 ( .A(n4826), .B(n20550), .Z(n4827) );
  AND U8543 ( .A(n20551), .B(n4827), .Z(n4830) );
  NANDN U8544 ( .A(y[404]), .B(x[404]), .Z(n4829) );
  NANDN U8545 ( .A(y[405]), .B(x[405]), .Z(n4828) );
  AND U8546 ( .A(n4829), .B(n4828), .Z(n20553) );
  NANDN U8547 ( .A(n4830), .B(n20553), .Z(n4833) );
  NANDN U8548 ( .A(x[406]), .B(y[406]), .Z(n4832) );
  NANDN U8549 ( .A(x[405]), .B(y[405]), .Z(n4831) );
  AND U8550 ( .A(n4832), .B(n4831), .Z(n20555) );
  NAND U8551 ( .A(n4833), .B(n20555), .Z(n4836) );
  NANDN U8552 ( .A(y[406]), .B(x[406]), .Z(n4835) );
  NANDN U8553 ( .A(y[407]), .B(x[407]), .Z(n4834) );
  AND U8554 ( .A(n4835), .B(n4834), .Z(n20557) );
  NAND U8555 ( .A(n4836), .B(n20557), .Z(n4839) );
  NANDN U8556 ( .A(x[408]), .B(y[408]), .Z(n4838) );
  NANDN U8557 ( .A(x[407]), .B(y[407]), .Z(n4837) );
  AND U8558 ( .A(n4838), .B(n4837), .Z(n20559) );
  NAND U8559 ( .A(n4839), .B(n20559), .Z(n4842) );
  NANDN U8560 ( .A(y[408]), .B(x[408]), .Z(n4841) );
  NANDN U8561 ( .A(y[409]), .B(x[409]), .Z(n4840) );
  AND U8562 ( .A(n4841), .B(n4840), .Z(n20562) );
  NAND U8563 ( .A(n4842), .B(n20562), .Z(n4843) );
  AND U8564 ( .A(n20563), .B(n4843), .Z(n4846) );
  NANDN U8565 ( .A(y[410]), .B(x[410]), .Z(n4845) );
  NANDN U8566 ( .A(y[411]), .B(x[411]), .Z(n4844) );
  AND U8567 ( .A(n4845), .B(n4844), .Z(n20565) );
  NANDN U8568 ( .A(n4846), .B(n20565), .Z(n4849) );
  NANDN U8569 ( .A(x[412]), .B(y[412]), .Z(n4848) );
  NANDN U8570 ( .A(x[411]), .B(y[411]), .Z(n4847) );
  AND U8571 ( .A(n4848), .B(n4847), .Z(n20567) );
  NAND U8572 ( .A(n4849), .B(n20567), .Z(n4852) );
  NANDN U8573 ( .A(y[412]), .B(x[412]), .Z(n4851) );
  NANDN U8574 ( .A(y[413]), .B(x[413]), .Z(n4850) );
  AND U8575 ( .A(n4851), .B(n4850), .Z(n20569) );
  NAND U8576 ( .A(n4852), .B(n20569), .Z(n4855) );
  NANDN U8577 ( .A(x[414]), .B(y[414]), .Z(n4854) );
  NANDN U8578 ( .A(x[413]), .B(y[413]), .Z(n4853) );
  AND U8579 ( .A(n4854), .B(n4853), .Z(n20571) );
  NAND U8580 ( .A(n4855), .B(n20571), .Z(n4858) );
  NANDN U8581 ( .A(y[414]), .B(x[414]), .Z(n4857) );
  NANDN U8582 ( .A(y[415]), .B(x[415]), .Z(n4856) );
  AND U8583 ( .A(n4857), .B(n4856), .Z(n20574) );
  NAND U8584 ( .A(n4858), .B(n20574), .Z(n4859) );
  AND U8585 ( .A(n20575), .B(n4859), .Z(n4862) );
  NANDN U8586 ( .A(y[416]), .B(x[416]), .Z(n4861) );
  NANDN U8587 ( .A(y[417]), .B(x[417]), .Z(n4860) );
  AND U8588 ( .A(n4861), .B(n4860), .Z(n20577) );
  NANDN U8589 ( .A(n4862), .B(n20577), .Z(n4865) );
  NANDN U8590 ( .A(x[418]), .B(y[418]), .Z(n4864) );
  NANDN U8591 ( .A(x[417]), .B(y[417]), .Z(n4863) );
  AND U8592 ( .A(n4864), .B(n4863), .Z(n20579) );
  NAND U8593 ( .A(n4865), .B(n20579), .Z(n4868) );
  NANDN U8594 ( .A(y[418]), .B(x[418]), .Z(n4867) );
  NANDN U8595 ( .A(y[419]), .B(x[419]), .Z(n4866) );
  AND U8596 ( .A(n4867), .B(n4866), .Z(n20581) );
  NAND U8597 ( .A(n4868), .B(n20581), .Z(n4871) );
  NANDN U8598 ( .A(x[420]), .B(y[420]), .Z(n4870) );
  NANDN U8599 ( .A(x[419]), .B(y[419]), .Z(n4869) );
  AND U8600 ( .A(n4870), .B(n4869), .Z(n20583) );
  NAND U8601 ( .A(n4871), .B(n20583), .Z(n4874) );
  NANDN U8602 ( .A(y[420]), .B(x[420]), .Z(n4873) );
  NANDN U8603 ( .A(y[421]), .B(x[421]), .Z(n4872) );
  AND U8604 ( .A(n4873), .B(n4872), .Z(n20586) );
  NAND U8605 ( .A(n4874), .B(n20586), .Z(n4875) );
  AND U8606 ( .A(n20587), .B(n4875), .Z(n4878) );
  NANDN U8607 ( .A(y[422]), .B(x[422]), .Z(n4877) );
  NANDN U8608 ( .A(y[423]), .B(x[423]), .Z(n4876) );
  AND U8609 ( .A(n4877), .B(n4876), .Z(n20590) );
  NANDN U8610 ( .A(n4878), .B(n20590), .Z(n4881) );
  NANDN U8611 ( .A(x[424]), .B(y[424]), .Z(n4880) );
  NANDN U8612 ( .A(x[423]), .B(y[423]), .Z(n4879) );
  AND U8613 ( .A(n4880), .B(n4879), .Z(n20591) );
  NAND U8614 ( .A(n4881), .B(n20591), .Z(n4884) );
  NANDN U8615 ( .A(y[425]), .B(x[425]), .Z(n4883) );
  NANDN U8616 ( .A(y[424]), .B(x[424]), .Z(n4882) );
  AND U8617 ( .A(n4883), .B(n4882), .Z(n20593) );
  NAND U8618 ( .A(n4884), .B(n20593), .Z(n4885) );
  NANDN U8619 ( .A(n13563), .B(n4885), .Z(n4886) );
  NANDN U8620 ( .A(n13564), .B(n4886), .Z(n4887) );
  AND U8621 ( .A(n20603), .B(n4887), .Z(n4890) );
  NANDN U8622 ( .A(y[428]), .B(x[428]), .Z(n4889) );
  NANDN U8623 ( .A(y[429]), .B(x[429]), .Z(n4888) );
  AND U8624 ( .A(n4889), .B(n4888), .Z(n20605) );
  NANDN U8625 ( .A(n4890), .B(n20605), .Z(n4893) );
  NANDN U8626 ( .A(x[430]), .B(y[430]), .Z(n4892) );
  NANDN U8627 ( .A(x[429]), .B(y[429]), .Z(n4891) );
  AND U8628 ( .A(n4892), .B(n4891), .Z(n20607) );
  NAND U8629 ( .A(n4893), .B(n20607), .Z(n4896) );
  NANDN U8630 ( .A(y[430]), .B(x[430]), .Z(n4895) );
  NANDN U8631 ( .A(y[431]), .B(x[431]), .Z(n4894) );
  AND U8632 ( .A(n4895), .B(n4894), .Z(n20609) );
  NAND U8633 ( .A(n4896), .B(n20609), .Z(n4899) );
  NANDN U8634 ( .A(x[432]), .B(y[432]), .Z(n4898) );
  NANDN U8635 ( .A(x[431]), .B(y[431]), .Z(n4897) );
  AND U8636 ( .A(n4898), .B(n4897), .Z(n20611) );
  NAND U8637 ( .A(n4899), .B(n20611), .Z(n4902) );
  NANDN U8638 ( .A(y[432]), .B(x[432]), .Z(n4901) );
  NANDN U8639 ( .A(y[433]), .B(x[433]), .Z(n4900) );
  AND U8640 ( .A(n4901), .B(n4900), .Z(n20614) );
  NAND U8641 ( .A(n4902), .B(n20614), .Z(n4903) );
  AND U8642 ( .A(n20615), .B(n4903), .Z(n4906) );
  NANDN U8643 ( .A(y[435]), .B(x[435]), .Z(n4905) );
  NANDN U8644 ( .A(y[434]), .B(x[434]), .Z(n4904) );
  AND U8645 ( .A(n4905), .B(n4904), .Z(n20617) );
  NANDN U8646 ( .A(n4906), .B(n20617), .Z(n4908) );
  NANDN U8647 ( .A(x[435]), .B(y[435]), .Z(n20619) );
  IV U8648 ( .A(x[436]), .Z(n20622) );
  NAND U8649 ( .A(n20622), .B(y[436]), .Z(n4907) );
  AND U8650 ( .A(n20619), .B(n4907), .Z(n13574) );
  NAND U8651 ( .A(n4908), .B(n13574), .Z(n4909) );
  NANDN U8652 ( .A(n13577), .B(n4909), .Z(n4912) );
  NANDN U8653 ( .A(x[438]), .B(y[438]), .Z(n4911) );
  NANDN U8654 ( .A(x[437]), .B(y[437]), .Z(n4910) );
  AND U8655 ( .A(n4911), .B(n4910), .Z(n20628) );
  NAND U8656 ( .A(n4912), .B(n20628), .Z(n4915) );
  NANDN U8657 ( .A(y[438]), .B(x[438]), .Z(n4914) );
  NANDN U8658 ( .A(y[439]), .B(x[439]), .Z(n4913) );
  AND U8659 ( .A(n4914), .B(n4913), .Z(n20630) );
  NAND U8660 ( .A(n4915), .B(n20630), .Z(n4916) );
  AND U8661 ( .A(n20632), .B(n4916), .Z(n4921) );
  NANDN U8662 ( .A(y[440]), .B(x[440]), .Z(n4917) );
  NANDN U8663 ( .A(n4917), .B(x[441]), .Z(n4920) );
  XNOR U8664 ( .A(n4917), .B(x[441]), .Z(n4918) );
  NANDN U8665 ( .A(y[441]), .B(n4918), .Z(n4919) );
  AND U8666 ( .A(n4920), .B(n4919), .Z(n20634) );
  NANDN U8667 ( .A(n4921), .B(n20634), .Z(n4922) );
  NANDN U8668 ( .A(x[442]), .B(y[442]), .Z(n20636) );
  NAND U8669 ( .A(n4922), .B(n20636), .Z(n4925) );
  NANDN U8670 ( .A(y[442]), .B(x[442]), .Z(n4924) );
  NANDN U8671 ( .A(y[443]), .B(x[443]), .Z(n4923) );
  AND U8672 ( .A(n4924), .B(n4923), .Z(n20639) );
  NAND U8673 ( .A(n4925), .B(n20639), .Z(n4928) );
  NANDN U8674 ( .A(x[444]), .B(y[444]), .Z(n4927) );
  NANDN U8675 ( .A(x[443]), .B(y[443]), .Z(n4926) );
  AND U8676 ( .A(n4927), .B(n4926), .Z(n20640) );
  NAND U8677 ( .A(n4928), .B(n20640), .Z(n4931) );
  NANDN U8678 ( .A(y[444]), .B(x[444]), .Z(n4930) );
  NANDN U8679 ( .A(y[445]), .B(x[445]), .Z(n4929) );
  AND U8680 ( .A(n4930), .B(n4929), .Z(n20642) );
  NAND U8681 ( .A(n4931), .B(n20642), .Z(n4932) );
  AND U8682 ( .A(n20644), .B(n4932), .Z(n4935) );
  NANDN U8683 ( .A(y[446]), .B(x[446]), .Z(n4934) );
  NANDN U8684 ( .A(y[447]), .B(x[447]), .Z(n4933) );
  AND U8685 ( .A(n4934), .B(n4933), .Z(n20646) );
  NANDN U8686 ( .A(n4935), .B(n20646), .Z(n4938) );
  NANDN U8687 ( .A(x[448]), .B(y[448]), .Z(n4937) );
  NANDN U8688 ( .A(x[447]), .B(y[447]), .Z(n4936) );
  AND U8689 ( .A(n4937), .B(n4936), .Z(n20648) );
  NAND U8690 ( .A(n4938), .B(n20648), .Z(n4941) );
  NANDN U8691 ( .A(y[448]), .B(x[448]), .Z(n4940) );
  NANDN U8692 ( .A(y[449]), .B(x[449]), .Z(n4939) );
  AND U8693 ( .A(n4940), .B(n4939), .Z(n20651) );
  NAND U8694 ( .A(n4941), .B(n20651), .Z(n4944) );
  NANDN U8695 ( .A(x[450]), .B(y[450]), .Z(n4943) );
  NANDN U8696 ( .A(x[449]), .B(y[449]), .Z(n4942) );
  AND U8697 ( .A(n4943), .B(n4942), .Z(n20652) );
  NAND U8698 ( .A(n4944), .B(n20652), .Z(n4947) );
  NANDN U8699 ( .A(y[450]), .B(x[450]), .Z(n4946) );
  NANDN U8700 ( .A(y[451]), .B(x[451]), .Z(n4945) );
  AND U8701 ( .A(n4946), .B(n4945), .Z(n20654) );
  NAND U8702 ( .A(n4947), .B(n20654), .Z(n4948) );
  AND U8703 ( .A(n20656), .B(n4948), .Z(n4949) );
  OR U8704 ( .A(n20659), .B(n4949), .Z(n4952) );
  NANDN U8705 ( .A(x[456]), .B(y[456]), .Z(n4951) );
  NANDN U8706 ( .A(x[455]), .B(y[455]), .Z(n4950) );
  AND U8707 ( .A(n4951), .B(n4950), .Z(n20660) );
  NAND U8708 ( .A(n4952), .B(n20660), .Z(n4955) );
  NANDN U8709 ( .A(y[456]), .B(x[456]), .Z(n4954) );
  NANDN U8710 ( .A(y[457]), .B(x[457]), .Z(n4953) );
  AND U8711 ( .A(n4954), .B(n4953), .Z(n20663) );
  NAND U8712 ( .A(n4955), .B(n20663), .Z(n4958) );
  NANDN U8713 ( .A(x[458]), .B(y[458]), .Z(n4957) );
  NANDN U8714 ( .A(x[457]), .B(y[457]), .Z(n4956) );
  AND U8715 ( .A(n4957), .B(n4956), .Z(n20664) );
  NAND U8716 ( .A(n4958), .B(n20664), .Z(n4961) );
  NANDN U8717 ( .A(y[458]), .B(x[458]), .Z(n4960) );
  NANDN U8718 ( .A(y[459]), .B(x[459]), .Z(n4959) );
  AND U8719 ( .A(n4960), .B(n4959), .Z(n20666) );
  NAND U8720 ( .A(n4961), .B(n20666), .Z(n4962) );
  AND U8721 ( .A(n20668), .B(n4962), .Z(n4965) );
  NANDN U8722 ( .A(y[460]), .B(x[460]), .Z(n4964) );
  NANDN U8723 ( .A(y[461]), .B(x[461]), .Z(n4963) );
  AND U8724 ( .A(n4964), .B(n4963), .Z(n20670) );
  NANDN U8725 ( .A(n4965), .B(n20670), .Z(n4968) );
  NANDN U8726 ( .A(x[462]), .B(y[462]), .Z(n4967) );
  NANDN U8727 ( .A(x[461]), .B(y[461]), .Z(n4966) );
  AND U8728 ( .A(n4967), .B(n4966), .Z(n20672) );
  NAND U8729 ( .A(n4968), .B(n20672), .Z(n4971) );
  NANDN U8730 ( .A(y[462]), .B(x[462]), .Z(n4970) );
  NANDN U8731 ( .A(y[463]), .B(x[463]), .Z(n4969) );
  AND U8732 ( .A(n4970), .B(n4969), .Z(n20675) );
  NAND U8733 ( .A(n4971), .B(n20675), .Z(n4974) );
  NANDN U8734 ( .A(x[464]), .B(y[464]), .Z(n4973) );
  NANDN U8735 ( .A(x[463]), .B(y[463]), .Z(n4972) );
  AND U8736 ( .A(n4973), .B(n4972), .Z(n20676) );
  NAND U8737 ( .A(n4974), .B(n20676), .Z(n4977) );
  NANDN U8738 ( .A(y[464]), .B(x[464]), .Z(n4976) );
  NANDN U8739 ( .A(y[465]), .B(x[465]), .Z(n4975) );
  AND U8740 ( .A(n4976), .B(n4975), .Z(n20678) );
  NAND U8741 ( .A(n4977), .B(n20678), .Z(n4978) );
  AND U8742 ( .A(n20680), .B(n4978), .Z(n4981) );
  NANDN U8743 ( .A(y[466]), .B(x[466]), .Z(n4980) );
  NANDN U8744 ( .A(y[467]), .B(x[467]), .Z(n4979) );
  AND U8745 ( .A(n4980), .B(n4979), .Z(n20682) );
  NANDN U8746 ( .A(n4981), .B(n20682), .Z(n4984) );
  NANDN U8747 ( .A(x[468]), .B(y[468]), .Z(n4983) );
  NANDN U8748 ( .A(x[467]), .B(y[467]), .Z(n4982) );
  AND U8749 ( .A(n4983), .B(n4982), .Z(n20684) );
  NAND U8750 ( .A(n4984), .B(n20684), .Z(n4987) );
  NANDN U8751 ( .A(y[468]), .B(x[468]), .Z(n4986) );
  NANDN U8752 ( .A(y[469]), .B(x[469]), .Z(n4985) );
  AND U8753 ( .A(n4986), .B(n4985), .Z(n20687) );
  NAND U8754 ( .A(n4987), .B(n20687), .Z(n4990) );
  NANDN U8755 ( .A(x[470]), .B(y[470]), .Z(n4989) );
  NANDN U8756 ( .A(x[469]), .B(y[469]), .Z(n4988) );
  AND U8757 ( .A(n4989), .B(n4988), .Z(n20688) );
  NAND U8758 ( .A(n4990), .B(n20688), .Z(n4993) );
  NANDN U8759 ( .A(y[470]), .B(x[470]), .Z(n4992) );
  NANDN U8760 ( .A(y[471]), .B(x[471]), .Z(n4991) );
  AND U8761 ( .A(n4992), .B(n4991), .Z(n20690) );
  NAND U8762 ( .A(n4993), .B(n20690), .Z(n4994) );
  AND U8763 ( .A(n20692), .B(n4994), .Z(n4997) );
  NANDN U8764 ( .A(y[472]), .B(x[472]), .Z(n4996) );
  NANDN U8765 ( .A(y[473]), .B(x[473]), .Z(n4995) );
  AND U8766 ( .A(n4996), .B(n4995), .Z(n20694) );
  NANDN U8767 ( .A(n4997), .B(n20694), .Z(n5000) );
  NANDN U8768 ( .A(x[474]), .B(y[474]), .Z(n4999) );
  NANDN U8769 ( .A(x[473]), .B(y[473]), .Z(n4998) );
  AND U8770 ( .A(n4999), .B(n4998), .Z(n20696) );
  NAND U8771 ( .A(n5000), .B(n20696), .Z(n5003) );
  NANDN U8772 ( .A(y[474]), .B(x[474]), .Z(n5002) );
  NANDN U8773 ( .A(y[475]), .B(x[475]), .Z(n5001) );
  AND U8774 ( .A(n5002), .B(n5001), .Z(n20699) );
  NAND U8775 ( .A(n5003), .B(n20699), .Z(n5006) );
  NANDN U8776 ( .A(x[476]), .B(y[476]), .Z(n5005) );
  NANDN U8777 ( .A(x[475]), .B(y[475]), .Z(n5004) );
  AND U8778 ( .A(n5005), .B(n5004), .Z(n20700) );
  NAND U8779 ( .A(n5006), .B(n20700), .Z(n5009) );
  NANDN U8780 ( .A(y[476]), .B(x[476]), .Z(n5008) );
  NANDN U8781 ( .A(y[477]), .B(x[477]), .Z(n5007) );
  AND U8782 ( .A(n5008), .B(n5007), .Z(n20702) );
  NAND U8783 ( .A(n5009), .B(n20702), .Z(n5010) );
  AND U8784 ( .A(n20704), .B(n5010), .Z(n5013) );
  NANDN U8785 ( .A(y[478]), .B(x[478]), .Z(n5012) );
  NANDN U8786 ( .A(y[479]), .B(x[479]), .Z(n5011) );
  AND U8787 ( .A(n5012), .B(n5011), .Z(n20706) );
  NANDN U8788 ( .A(n5013), .B(n20706), .Z(n5016) );
  NANDN U8789 ( .A(x[480]), .B(y[480]), .Z(n5015) );
  NANDN U8790 ( .A(x[479]), .B(y[479]), .Z(n5014) );
  AND U8791 ( .A(n5015), .B(n5014), .Z(n20708) );
  NAND U8792 ( .A(n5016), .B(n20708), .Z(n5019) );
  NANDN U8793 ( .A(y[481]), .B(x[481]), .Z(n5018) );
  NANDN U8794 ( .A(y[480]), .B(x[480]), .Z(n5017) );
  AND U8795 ( .A(n5018), .B(n5017), .Z(n20711) );
  NAND U8796 ( .A(n5019), .B(n20711), .Z(n5020) );
  NAND U8797 ( .A(n20712), .B(n5020), .Z(n5022) );
  IV U8798 ( .A(x[482]), .Z(n13622) );
  AND U8799 ( .A(y[482]), .B(n13622), .Z(n5021) );
  OR U8800 ( .A(n5022), .B(n5021), .Z(n5023) );
  NANDN U8801 ( .A(n20715), .B(n5023), .Z(n5024) );
  NANDN U8802 ( .A(n13623), .B(n5024), .Z(n5025) );
  OR U8803 ( .A(n13628), .B(n5025), .Z(n5026) );
  NANDN U8804 ( .A(n20719), .B(n5026), .Z(n5029) );
  NANDN U8805 ( .A(x[485]), .B(y[485]), .Z(n5028) );
  NANDN U8806 ( .A(x[486]), .B(y[486]), .Z(n5027) );
  AND U8807 ( .A(n5028), .B(n5027), .Z(n20720) );
  NAND U8808 ( .A(n5029), .B(n20720), .Z(n5030) );
  NANDN U8809 ( .A(n20722), .B(n5030), .Z(n5033) );
  NANDN U8810 ( .A(x[487]), .B(y[487]), .Z(n5032) );
  NANDN U8811 ( .A(x[488]), .B(y[488]), .Z(n5031) );
  AND U8812 ( .A(n5032), .B(n5031), .Z(n20724) );
  NAND U8813 ( .A(n5033), .B(n20724), .Z(n5036) );
  NANDN U8814 ( .A(y[489]), .B(x[489]), .Z(n5035) );
  NANDN U8815 ( .A(y[488]), .B(x[488]), .Z(n5034) );
  NAND U8816 ( .A(n5035), .B(n5034), .Z(n20727) );
  ANDN U8817 ( .B(n5036), .A(n20727), .Z(n5039) );
  NANDN U8818 ( .A(x[489]), .B(y[489]), .Z(n5038) );
  NANDN U8819 ( .A(x[490]), .B(y[490]), .Z(n5037) );
  AND U8820 ( .A(n5038), .B(n5037), .Z(n20728) );
  NANDN U8821 ( .A(n5039), .B(n20728), .Z(n5040) );
  NANDN U8822 ( .A(n20731), .B(n5040), .Z(n5043) );
  NANDN U8823 ( .A(x[491]), .B(y[491]), .Z(n5042) );
  NANDN U8824 ( .A(x[492]), .B(y[492]), .Z(n5041) );
  AND U8825 ( .A(n5042), .B(n5041), .Z(n20732) );
  NAND U8826 ( .A(n5043), .B(n20732), .Z(n5044) );
  NANDN U8827 ( .A(n20734), .B(n5044), .Z(n5047) );
  NANDN U8828 ( .A(x[493]), .B(y[493]), .Z(n5046) );
  NANDN U8829 ( .A(x[494]), .B(y[494]), .Z(n5045) );
  AND U8830 ( .A(n5046), .B(n5045), .Z(n20736) );
  NAND U8831 ( .A(n5047), .B(n20736), .Z(n5050) );
  NANDN U8832 ( .A(y[495]), .B(x[495]), .Z(n5049) );
  NANDN U8833 ( .A(y[494]), .B(x[494]), .Z(n5048) );
  NAND U8834 ( .A(n5049), .B(n5048), .Z(n20739) );
  ANDN U8835 ( .B(n5050), .A(n20739), .Z(n5053) );
  NANDN U8836 ( .A(x[495]), .B(y[495]), .Z(n5052) );
  NANDN U8837 ( .A(x[496]), .B(y[496]), .Z(n5051) );
  AND U8838 ( .A(n5052), .B(n5051), .Z(n20740) );
  NANDN U8839 ( .A(n5053), .B(n20740), .Z(n5054) );
  NANDN U8840 ( .A(n20743), .B(n5054), .Z(n5057) );
  NANDN U8841 ( .A(x[497]), .B(y[497]), .Z(n5056) );
  NANDN U8842 ( .A(x[498]), .B(y[498]), .Z(n5055) );
  AND U8843 ( .A(n5056), .B(n5055), .Z(n20744) );
  NAND U8844 ( .A(n5057), .B(n20744), .Z(n5058) );
  NANDN U8845 ( .A(n20746), .B(n5058), .Z(n5061) );
  NANDN U8846 ( .A(x[499]), .B(y[499]), .Z(n5060) );
  NANDN U8847 ( .A(x[500]), .B(y[500]), .Z(n5059) );
  AND U8848 ( .A(n5060), .B(n5059), .Z(n20748) );
  NAND U8849 ( .A(n5061), .B(n20748), .Z(n5064) );
  NANDN U8850 ( .A(y[501]), .B(x[501]), .Z(n5063) );
  NANDN U8851 ( .A(y[500]), .B(x[500]), .Z(n5062) );
  NAND U8852 ( .A(n5063), .B(n5062), .Z(n20751) );
  ANDN U8853 ( .B(n5064), .A(n20751), .Z(n5067) );
  NANDN U8854 ( .A(x[501]), .B(y[501]), .Z(n5066) );
  NANDN U8855 ( .A(x[502]), .B(y[502]), .Z(n5065) );
  AND U8856 ( .A(n5066), .B(n5065), .Z(n20752) );
  NANDN U8857 ( .A(n5067), .B(n20752), .Z(n5068) );
  NANDN U8858 ( .A(n20755), .B(n5068), .Z(n5071) );
  NANDN U8859 ( .A(x[503]), .B(y[503]), .Z(n5070) );
  NANDN U8860 ( .A(x[504]), .B(y[504]), .Z(n5069) );
  AND U8861 ( .A(n5070), .B(n5069), .Z(n20756) );
  NAND U8862 ( .A(n5071), .B(n20756), .Z(n5072) );
  NANDN U8863 ( .A(n20758), .B(n5072), .Z(n5075) );
  NANDN U8864 ( .A(x[505]), .B(y[505]), .Z(n5074) );
  NANDN U8865 ( .A(x[506]), .B(y[506]), .Z(n5073) );
  AND U8866 ( .A(n5074), .B(n5073), .Z(n20760) );
  NAND U8867 ( .A(n5075), .B(n20760), .Z(n5078) );
  NANDN U8868 ( .A(y[507]), .B(x[507]), .Z(n5077) );
  NANDN U8869 ( .A(y[506]), .B(x[506]), .Z(n5076) );
  NAND U8870 ( .A(n5077), .B(n5076), .Z(n20763) );
  ANDN U8871 ( .B(n5078), .A(n20763), .Z(n5081) );
  NANDN U8872 ( .A(x[507]), .B(y[507]), .Z(n5080) );
  NANDN U8873 ( .A(x[508]), .B(y[508]), .Z(n5079) );
  AND U8874 ( .A(n5080), .B(n5079), .Z(n20764) );
  NANDN U8875 ( .A(n5081), .B(n20764), .Z(n5082) );
  NANDN U8876 ( .A(n20767), .B(n5082), .Z(n5087) );
  NANDN U8877 ( .A(x[510]), .B(y[510]), .Z(n5084) );
  NANDN U8878 ( .A(x[509]), .B(y[509]), .Z(n5083) );
  AND U8879 ( .A(n5084), .B(n5083), .Z(n5086) );
  AND U8880 ( .A(n5086), .B(n5085), .Z(n20768) );
  NAND U8881 ( .A(n5087), .B(n20768), .Z(n5088) );
  NANDN U8882 ( .A(n20770), .B(n5088), .Z(n5089) );
  NANDN U8883 ( .A(x[512]), .B(y[512]), .Z(n20772) );
  NAND U8884 ( .A(n5089), .B(n20772), .Z(n5092) );
  NANDN U8885 ( .A(y[512]), .B(x[512]), .Z(n5091) );
  NANDN U8886 ( .A(y[513]), .B(x[513]), .Z(n5090) );
  NAND U8887 ( .A(n5091), .B(n5090), .Z(n20775) );
  ANDN U8888 ( .B(n5092), .A(n20775), .Z(n5094) );
  NANDN U8889 ( .A(x[513]), .B(y[513]), .Z(n20776) );
  ANDN U8890 ( .B(y[514]), .A(x[514]), .Z(n12761) );
  ANDN U8891 ( .B(n20776), .A(n12761), .Z(n5093) );
  NANDN U8892 ( .A(n5094), .B(n5093), .Z(n5095) );
  AND U8893 ( .A(n20778), .B(n5095), .Z(n5096) );
  OR U8894 ( .A(n12764), .B(n5096), .Z(n5097) );
  NANDN U8895 ( .A(n20782), .B(n5097), .Z(n5100) );
  NANDN U8896 ( .A(x[517]), .B(y[517]), .Z(n5099) );
  NANDN U8897 ( .A(x[518]), .B(y[518]), .Z(n5098) );
  AND U8898 ( .A(n5099), .B(n5098), .Z(n20784) );
  NAND U8899 ( .A(n5100), .B(n20784), .Z(n5101) );
  NANDN U8900 ( .A(n20787), .B(n5101), .Z(n5105) );
  ANDN U8901 ( .B(y[520]), .A(x[520]), .Z(n12757) );
  NANDN U8902 ( .A(x[522]), .B(y[522]), .Z(n5103) );
  NANDN U8903 ( .A(x[521]), .B(y[521]), .Z(n5102) );
  NAND U8904 ( .A(n5103), .B(n5102), .Z(n5110) );
  NANDN U8905 ( .A(x[519]), .B(y[519]), .Z(n5104) );
  NANDN U8906 ( .A(n5110), .B(n5104), .Z(n13666) );
  NOR U8907 ( .A(n12757), .B(n13666), .Z(n20788) );
  NAND U8908 ( .A(n5105), .B(n20788), .Z(n5112) );
  NANDN U8909 ( .A(y[523]), .B(x[523]), .Z(n5107) );
  NANDN U8910 ( .A(y[522]), .B(x[522]), .Z(n5106) );
  NAND U8911 ( .A(n5107), .B(n5106), .Z(n12756) );
  ANDN U8912 ( .B(x[521]), .A(y[521]), .Z(n12759) );
  NANDN U8913 ( .A(y[520]), .B(x[520]), .Z(n5108) );
  NANDN U8914 ( .A(n12759), .B(n5108), .Z(n5109) );
  NANDN U8915 ( .A(n5110), .B(n5109), .Z(n5111) );
  NANDN U8916 ( .A(n12756), .B(n5111), .Z(n20791) );
  ANDN U8917 ( .B(n5112), .A(n20791), .Z(n5115) );
  NANDN U8918 ( .A(x[523]), .B(y[523]), .Z(n5114) );
  NANDN U8919 ( .A(x[524]), .B(y[524]), .Z(n5113) );
  AND U8920 ( .A(n5114), .B(n5113), .Z(n20792) );
  NANDN U8921 ( .A(n5115), .B(n20792), .Z(n5116) );
  NANDN U8922 ( .A(n20794), .B(n5116), .Z(n5119) );
  NANDN U8923 ( .A(x[525]), .B(y[525]), .Z(n5118) );
  NANDN U8924 ( .A(x[526]), .B(y[526]), .Z(n5117) );
  AND U8925 ( .A(n5118), .B(n5117), .Z(n20796) );
  NAND U8926 ( .A(n5119), .B(n20796), .Z(n5120) );
  NANDN U8927 ( .A(n20799), .B(n5120), .Z(n5123) );
  NANDN U8928 ( .A(x[527]), .B(y[527]), .Z(n5122) );
  NANDN U8929 ( .A(x[528]), .B(y[528]), .Z(n5121) );
  AND U8930 ( .A(n5122), .B(n5121), .Z(n20800) );
  NAND U8931 ( .A(n5123), .B(n20800), .Z(n5126) );
  NANDN U8932 ( .A(y[528]), .B(x[528]), .Z(n5125) );
  NANDN U8933 ( .A(y[529]), .B(x[529]), .Z(n5124) );
  NAND U8934 ( .A(n5125), .B(n5124), .Z(n20803) );
  ANDN U8935 ( .B(n5126), .A(n20803), .Z(n5128) );
  NANDN U8936 ( .A(x[529]), .B(y[529]), .Z(n20804) );
  ANDN U8937 ( .B(y[530]), .A(x[530]), .Z(n12752) );
  ANDN U8938 ( .B(n20804), .A(n12752), .Z(n5127) );
  NANDN U8939 ( .A(n5128), .B(n5127), .Z(n5129) );
  AND U8940 ( .A(n20807), .B(n5129), .Z(n5130) );
  OR U8941 ( .A(n12755), .B(n5130), .Z(n5131) );
  NANDN U8942 ( .A(n20811), .B(n5131), .Z(n5134) );
  NANDN U8943 ( .A(x[533]), .B(y[533]), .Z(n5133) );
  NANDN U8944 ( .A(x[534]), .B(y[534]), .Z(n5132) );
  AND U8945 ( .A(n5133), .B(n5132), .Z(n20812) );
  NAND U8946 ( .A(n5134), .B(n20812), .Z(n5135) );
  NANDN U8947 ( .A(n20815), .B(n5135), .Z(n5138) );
  NANDN U8948 ( .A(x[535]), .B(y[535]), .Z(n5137) );
  NANDN U8949 ( .A(x[536]), .B(y[536]), .Z(n5136) );
  AND U8950 ( .A(n5137), .B(n5136), .Z(n20816) );
  NAND U8951 ( .A(n5138), .B(n20816), .Z(n5141) );
  NANDN U8952 ( .A(y[537]), .B(x[537]), .Z(n5140) );
  NANDN U8953 ( .A(y[536]), .B(x[536]), .Z(n5139) );
  NAND U8954 ( .A(n5140), .B(n5139), .Z(n20818) );
  ANDN U8955 ( .B(n5141), .A(n20818), .Z(n5144) );
  NANDN U8956 ( .A(x[537]), .B(y[537]), .Z(n5143) );
  NANDN U8957 ( .A(x[538]), .B(y[538]), .Z(n5142) );
  AND U8958 ( .A(n5143), .B(n5142), .Z(n20820) );
  NANDN U8959 ( .A(n5144), .B(n20820), .Z(n5145) );
  NANDN U8960 ( .A(n20823), .B(n5145), .Z(n5148) );
  NANDN U8961 ( .A(x[539]), .B(y[539]), .Z(n5147) );
  NANDN U8962 ( .A(x[540]), .B(y[540]), .Z(n5146) );
  AND U8963 ( .A(n5147), .B(n5146), .Z(n20824) );
  NAND U8964 ( .A(n5148), .B(n20824), .Z(n5149) );
  NANDN U8965 ( .A(n20827), .B(n5149), .Z(n5152) );
  NANDN U8966 ( .A(x[541]), .B(y[541]), .Z(n5151) );
  NANDN U8967 ( .A(x[542]), .B(y[542]), .Z(n5150) );
  AND U8968 ( .A(n5151), .B(n5150), .Z(n20828) );
  NAND U8969 ( .A(n5152), .B(n20828), .Z(n5155) );
  NANDN U8970 ( .A(y[543]), .B(x[543]), .Z(n5154) );
  NANDN U8971 ( .A(y[542]), .B(x[542]), .Z(n5153) );
  NAND U8972 ( .A(n5154), .B(n5153), .Z(n20830) );
  ANDN U8973 ( .B(n5155), .A(n20830), .Z(n5158) );
  NANDN U8974 ( .A(x[543]), .B(y[543]), .Z(n5157) );
  NANDN U8975 ( .A(x[544]), .B(y[544]), .Z(n5156) );
  AND U8976 ( .A(n5157), .B(n5156), .Z(n20832) );
  NANDN U8977 ( .A(n5158), .B(n20832), .Z(n5159) );
  NANDN U8978 ( .A(n20835), .B(n5159), .Z(n5164) );
  NANDN U8979 ( .A(x[546]), .B(y[546]), .Z(n5161) );
  NANDN U8980 ( .A(x[545]), .B(y[545]), .Z(n5160) );
  AND U8981 ( .A(n5161), .B(n5160), .Z(n5163) );
  AND U8982 ( .A(n5163), .B(n5162), .Z(n20836) );
  NAND U8983 ( .A(n5164), .B(n20836), .Z(n5165) );
  NANDN U8984 ( .A(n20839), .B(n5165), .Z(n5166) );
  NANDN U8985 ( .A(x[548]), .B(y[548]), .Z(n20840) );
  NAND U8986 ( .A(n5166), .B(n20840), .Z(n5169) );
  NANDN U8987 ( .A(y[549]), .B(x[549]), .Z(n5168) );
  NANDN U8988 ( .A(y[548]), .B(x[548]), .Z(n5167) );
  NAND U8989 ( .A(n5168), .B(n5167), .Z(n20842) );
  ANDN U8990 ( .B(n5169), .A(n20842), .Z(n5172) );
  NANDN U8991 ( .A(x[549]), .B(y[549]), .Z(n5171) );
  NANDN U8992 ( .A(x[550]), .B(y[550]), .Z(n5170) );
  AND U8993 ( .A(n5171), .B(n5170), .Z(n20844) );
  NANDN U8994 ( .A(n5172), .B(n20844), .Z(n5173) );
  NANDN U8995 ( .A(n20847), .B(n5173), .Z(n5176) );
  NANDN U8996 ( .A(x[551]), .B(y[551]), .Z(n5175) );
  NANDN U8997 ( .A(x[552]), .B(y[552]), .Z(n5174) );
  AND U8998 ( .A(n5175), .B(n5174), .Z(n20848) );
  NAND U8999 ( .A(n5176), .B(n20848), .Z(n5177) );
  NANDN U9000 ( .A(n20851), .B(n5177), .Z(n5180) );
  NANDN U9001 ( .A(x[553]), .B(y[553]), .Z(n5179) );
  NANDN U9002 ( .A(x[554]), .B(y[554]), .Z(n5178) );
  AND U9003 ( .A(n5179), .B(n5178), .Z(n20852) );
  NAND U9004 ( .A(n5180), .B(n20852), .Z(n5183) );
  NANDN U9005 ( .A(y[555]), .B(x[555]), .Z(n5182) );
  NANDN U9006 ( .A(y[554]), .B(x[554]), .Z(n5181) );
  NAND U9007 ( .A(n5182), .B(n5181), .Z(n20854) );
  ANDN U9008 ( .B(n5183), .A(n20854), .Z(n5186) );
  NANDN U9009 ( .A(x[555]), .B(y[555]), .Z(n5185) );
  NANDN U9010 ( .A(x[556]), .B(y[556]), .Z(n5184) );
  AND U9011 ( .A(n5185), .B(n5184), .Z(n20856) );
  NANDN U9012 ( .A(n5186), .B(n20856), .Z(n5187) );
  NANDN U9013 ( .A(n20859), .B(n5187), .Z(n5188) );
  NANDN U9014 ( .A(n20861), .B(n5188), .Z(n5189) );
  NANDN U9015 ( .A(n20863), .B(n5189), .Z(n5190) );
  NANDN U9016 ( .A(x[560]), .B(y[560]), .Z(n20864) );
  NAND U9017 ( .A(n5190), .B(n20864), .Z(n5193) );
  NANDN U9018 ( .A(y[561]), .B(x[561]), .Z(n5192) );
  NANDN U9019 ( .A(y[560]), .B(x[560]), .Z(n5191) );
  NAND U9020 ( .A(n5192), .B(n5191), .Z(n20866) );
  ANDN U9021 ( .B(n5193), .A(n20866), .Z(n5196) );
  NANDN U9022 ( .A(x[561]), .B(y[561]), .Z(n5195) );
  NANDN U9023 ( .A(x[562]), .B(y[562]), .Z(n5194) );
  AND U9024 ( .A(n5195), .B(n5194), .Z(n20868) );
  NANDN U9025 ( .A(n5196), .B(n20868), .Z(n5197) );
  NANDN U9026 ( .A(n20871), .B(n5197), .Z(n5200) );
  NANDN U9027 ( .A(x[563]), .B(y[563]), .Z(n5199) );
  NANDN U9028 ( .A(x[564]), .B(y[564]), .Z(n5198) );
  AND U9029 ( .A(n5199), .B(n5198), .Z(n20872) );
  NAND U9030 ( .A(n5200), .B(n20872), .Z(n5201) );
  NANDN U9031 ( .A(n20875), .B(n5201), .Z(n5202) );
  NANDN U9032 ( .A(x[567]), .B(y[567]), .Z(n20880) );
  ANDN U9033 ( .B(y[568]), .A(x[568]), .Z(n12749) );
  NANDN U9034 ( .A(y[570]), .B(x[570]), .Z(n5204) );
  NANDN U9035 ( .A(y[571]), .B(x[571]), .Z(n5203) );
  AND U9036 ( .A(n5204), .B(n5203), .Z(n20891) );
  NANDN U9037 ( .A(y[572]), .B(x[572]), .Z(n5206) );
  NANDN U9038 ( .A(y[573]), .B(x[573]), .Z(n5205) );
  AND U9039 ( .A(n5206), .B(n5205), .Z(n20894) );
  NANDN U9040 ( .A(x[574]), .B(y[574]), .Z(n5208) );
  NANDN U9041 ( .A(x[573]), .B(y[573]), .Z(n5207) );
  AND U9042 ( .A(n5208), .B(n5207), .Z(n20896) );
  NANDN U9043 ( .A(y[574]), .B(x[574]), .Z(n5210) );
  NANDN U9044 ( .A(y[575]), .B(x[575]), .Z(n5209) );
  AND U9045 ( .A(n5210), .B(n5209), .Z(n20898) );
  NANDN U9046 ( .A(x[576]), .B(y[576]), .Z(n5212) );
  NANDN U9047 ( .A(x[575]), .B(y[575]), .Z(n5211) );
  AND U9048 ( .A(n5212), .B(n5211), .Z(n20900) );
  NANDN U9049 ( .A(y[576]), .B(x[576]), .Z(n5214) );
  NANDN U9050 ( .A(y[577]), .B(x[577]), .Z(n5213) );
  AND U9051 ( .A(n5214), .B(n5213), .Z(n20903) );
  NANDN U9052 ( .A(x[578]), .B(y[578]), .Z(n5216) );
  NANDN U9053 ( .A(x[577]), .B(y[577]), .Z(n5215) );
  NAND U9054 ( .A(n5216), .B(n5215), .Z(n20905) );
  NANDN U9055 ( .A(y[578]), .B(x[578]), .Z(n5218) );
  NANDN U9056 ( .A(y[579]), .B(x[579]), .Z(n5217) );
  AND U9057 ( .A(n5218), .B(n5217), .Z(n20906) );
  NANDN U9058 ( .A(y[580]), .B(x[580]), .Z(n5220) );
  NANDN U9059 ( .A(n5220), .B(x[581]), .Z(n5223) );
  XOR U9060 ( .A(n5220), .B(n5219), .Z(n5221) );
  NANDN U9061 ( .A(y[581]), .B(n5221), .Z(n5222) );
  AND U9062 ( .A(n5223), .B(n5222), .Z(n20910) );
  NANDN U9063 ( .A(x[582]), .B(y[582]), .Z(n20912) );
  NANDN U9064 ( .A(y[582]), .B(x[582]), .Z(n5225) );
  NANDN U9065 ( .A(y[583]), .B(x[583]), .Z(n5224) );
  AND U9066 ( .A(n5225), .B(n5224), .Z(n20914) );
  NANDN U9067 ( .A(x[584]), .B(y[584]), .Z(n5227) );
  NANDN U9068 ( .A(x[583]), .B(y[583]), .Z(n5226) );
  NAND U9069 ( .A(n5227), .B(n5226), .Z(n20917) );
  ANDN U9070 ( .B(n5228), .A(n20917), .Z(n5231) );
  NANDN U9071 ( .A(y[584]), .B(x[584]), .Z(n5230) );
  NANDN U9072 ( .A(y[585]), .B(x[585]), .Z(n5229) );
  AND U9073 ( .A(n5230), .B(n5229), .Z(n20918) );
  NANDN U9074 ( .A(n5231), .B(n20918), .Z(n5232) );
  NANDN U9075 ( .A(n20920), .B(n5232), .Z(n5235) );
  NANDN U9076 ( .A(y[586]), .B(x[586]), .Z(n5234) );
  NANDN U9077 ( .A(y[587]), .B(x[587]), .Z(n5233) );
  AND U9078 ( .A(n5234), .B(n5233), .Z(n20922) );
  NAND U9079 ( .A(n5235), .B(n20922), .Z(n5236) );
  NANDN U9080 ( .A(n20925), .B(n5236), .Z(n5239) );
  NANDN U9081 ( .A(y[588]), .B(x[588]), .Z(n5238) );
  NANDN U9082 ( .A(y[589]), .B(x[589]), .Z(n5237) );
  AND U9083 ( .A(n5238), .B(n5237), .Z(n20926) );
  NAND U9084 ( .A(n5239), .B(n20926), .Z(n5242) );
  NANDN U9085 ( .A(x[590]), .B(y[590]), .Z(n5240) );
  NANDN U9086 ( .A(n5241), .B(n5240), .Z(n13747) );
  NANDN U9087 ( .A(x[589]), .B(y[589]), .Z(n13742) );
  NANDN U9088 ( .A(n13747), .B(n13742), .Z(n20929) );
  ANDN U9089 ( .B(n5242), .A(n20929), .Z(n5243) );
  OR U9090 ( .A(n20931), .B(n5243), .Z(n5244) );
  NANDN U9091 ( .A(x[592]), .B(y[592]), .Z(n20933) );
  NAND U9092 ( .A(n5244), .B(n20933), .Z(n5247) );
  NANDN U9093 ( .A(y[592]), .B(x[592]), .Z(n5246) );
  NANDN U9094 ( .A(y[593]), .B(x[593]), .Z(n5245) );
  AND U9095 ( .A(n5246), .B(n5245), .Z(n20934) );
  NAND U9096 ( .A(n5247), .B(n20934), .Z(n5248) );
  NANDN U9097 ( .A(n20937), .B(n5248), .Z(n5251) );
  NANDN U9098 ( .A(y[594]), .B(x[594]), .Z(n5250) );
  NANDN U9099 ( .A(y[595]), .B(x[595]), .Z(n5249) );
  AND U9100 ( .A(n5250), .B(n5249), .Z(n20938) );
  NAND U9101 ( .A(n5251), .B(n20938), .Z(n5254) );
  NANDN U9102 ( .A(x[596]), .B(y[596]), .Z(n5253) );
  NANDN U9103 ( .A(x[595]), .B(y[595]), .Z(n5252) );
  NAND U9104 ( .A(n5253), .B(n5252), .Z(n20941) );
  ANDN U9105 ( .B(n5254), .A(n20941), .Z(n5257) );
  NANDN U9106 ( .A(y[596]), .B(x[596]), .Z(n5256) );
  NANDN U9107 ( .A(y[597]), .B(x[597]), .Z(n5255) );
  AND U9108 ( .A(n5256), .B(n5255), .Z(n20942) );
  NANDN U9109 ( .A(n5257), .B(n20942), .Z(n5258) );
  NANDN U9110 ( .A(n20944), .B(n5258), .Z(n5261) );
  NANDN U9111 ( .A(y[598]), .B(x[598]), .Z(n5260) );
  NANDN U9112 ( .A(y[599]), .B(x[599]), .Z(n5259) );
  AND U9113 ( .A(n5260), .B(n5259), .Z(n20946) );
  NAND U9114 ( .A(n5261), .B(n20946), .Z(n5262) );
  NANDN U9115 ( .A(n20949), .B(n5262), .Z(n5265) );
  NANDN U9116 ( .A(y[600]), .B(x[600]), .Z(n5264) );
  NANDN U9117 ( .A(y[601]), .B(x[601]), .Z(n5263) );
  AND U9118 ( .A(n5264), .B(n5263), .Z(n20950) );
  NAND U9119 ( .A(n5265), .B(n20950), .Z(n5268) );
  NANDN U9120 ( .A(x[602]), .B(y[602]), .Z(n5267) );
  NANDN U9121 ( .A(x[601]), .B(y[601]), .Z(n5266) );
  NAND U9122 ( .A(n5267), .B(n5266), .Z(n20953) );
  ANDN U9123 ( .B(n5268), .A(n20953), .Z(n5269) );
  OR U9124 ( .A(n20955), .B(n5269), .Z(n5270) );
  NANDN U9125 ( .A(n20956), .B(n5270), .Z(n5271) );
  NANDN U9126 ( .A(n20959), .B(n5271), .Z(n5272) );
  NANDN U9127 ( .A(n20961), .B(n5272), .Z(n5275) );
  NANDN U9128 ( .A(y[606]), .B(x[606]), .Z(n5274) );
  NANDN U9129 ( .A(y[607]), .B(x[607]), .Z(n5273) );
  AND U9130 ( .A(n5274), .B(n5273), .Z(n20962) );
  NAND U9131 ( .A(n5275), .B(n20962), .Z(n5278) );
  NANDN U9132 ( .A(x[608]), .B(y[608]), .Z(n5277) );
  NANDN U9133 ( .A(x[607]), .B(y[607]), .Z(n5276) );
  NAND U9134 ( .A(n5277), .B(n5276), .Z(n20965) );
  ANDN U9135 ( .B(n5278), .A(n20965), .Z(n5281) );
  NANDN U9136 ( .A(y[608]), .B(x[608]), .Z(n5280) );
  NANDN U9137 ( .A(y[609]), .B(x[609]), .Z(n5279) );
  AND U9138 ( .A(n5280), .B(n5279), .Z(n20966) );
  NANDN U9139 ( .A(n5281), .B(n20966), .Z(n5282) );
  NANDN U9140 ( .A(n20968), .B(n5282), .Z(n5285) );
  NANDN U9141 ( .A(y[610]), .B(x[610]), .Z(n5284) );
  NANDN U9142 ( .A(y[611]), .B(x[611]), .Z(n5283) );
  AND U9143 ( .A(n5284), .B(n5283), .Z(n20970) );
  NAND U9144 ( .A(n5285), .B(n20970), .Z(n5286) );
  NANDN U9145 ( .A(n20973), .B(n5286), .Z(n5289) );
  NANDN U9146 ( .A(y[612]), .B(x[612]), .Z(n5288) );
  NANDN U9147 ( .A(y[613]), .B(x[613]), .Z(n5287) );
  AND U9148 ( .A(n5288), .B(n5287), .Z(n20974) );
  NAND U9149 ( .A(n5289), .B(n20974), .Z(n5292) );
  NANDN U9150 ( .A(x[614]), .B(y[614]), .Z(n5291) );
  NANDN U9151 ( .A(x[613]), .B(y[613]), .Z(n5290) );
  NAND U9152 ( .A(n5291), .B(n5290), .Z(n20977) );
  ANDN U9153 ( .B(n5292), .A(n20977), .Z(n5295) );
  NANDN U9154 ( .A(y[614]), .B(x[614]), .Z(n5294) );
  NANDN U9155 ( .A(y[615]), .B(x[615]), .Z(n5293) );
  AND U9156 ( .A(n5294), .B(n5293), .Z(n20978) );
  NANDN U9157 ( .A(n5295), .B(n20978), .Z(n5296) );
  NANDN U9158 ( .A(n20980), .B(n5296), .Z(n5299) );
  NANDN U9159 ( .A(y[616]), .B(x[616]), .Z(n5298) );
  NANDN U9160 ( .A(y[617]), .B(x[617]), .Z(n5297) );
  AND U9161 ( .A(n5298), .B(n5297), .Z(n20982) );
  NAND U9162 ( .A(n5299), .B(n20982), .Z(n5300) );
  NANDN U9163 ( .A(n20985), .B(n5300), .Z(n5303) );
  NANDN U9164 ( .A(y[618]), .B(x[618]), .Z(n5302) );
  NANDN U9165 ( .A(y[619]), .B(x[619]), .Z(n5301) );
  AND U9166 ( .A(n5302), .B(n5301), .Z(n20986) );
  NAND U9167 ( .A(n5303), .B(n20986), .Z(n5306) );
  NANDN U9168 ( .A(x[620]), .B(y[620]), .Z(n5305) );
  NANDN U9169 ( .A(x[619]), .B(y[619]), .Z(n5304) );
  NAND U9170 ( .A(n5305), .B(n5304), .Z(n20989) );
  ANDN U9171 ( .B(n5306), .A(n20989), .Z(n5309) );
  NANDN U9172 ( .A(y[620]), .B(x[620]), .Z(n5308) );
  NANDN U9173 ( .A(y[621]), .B(x[621]), .Z(n5307) );
  AND U9174 ( .A(n5308), .B(n5307), .Z(n20990) );
  NANDN U9175 ( .A(n5309), .B(n20990), .Z(n5310) );
  NANDN U9176 ( .A(n20992), .B(n5310), .Z(n5313) );
  NANDN U9177 ( .A(y[622]), .B(x[622]), .Z(n5312) );
  NANDN U9178 ( .A(y[623]), .B(x[623]), .Z(n5311) );
  AND U9179 ( .A(n5312), .B(n5311), .Z(n20994) );
  NAND U9180 ( .A(n5313), .B(n20994), .Z(n5314) );
  NANDN U9181 ( .A(n20997), .B(n5314), .Z(n5320) );
  NANDN U9182 ( .A(y[624]), .B(x[624]), .Z(n5316) );
  NANDN U9183 ( .A(n5316), .B(x[625]), .Z(n5319) );
  XOR U9184 ( .A(n5316), .B(n5315), .Z(n5317) );
  NANDN U9185 ( .A(y[625]), .B(n5317), .Z(n5318) );
  AND U9186 ( .A(n5319), .B(n5318), .Z(n20998) );
  NAND U9187 ( .A(n5320), .B(n20998), .Z(n5321) );
  AND U9188 ( .A(n21000), .B(n5321), .Z(n5324) );
  NANDN U9189 ( .A(y[626]), .B(x[626]), .Z(n5323) );
  NANDN U9190 ( .A(y[627]), .B(x[627]), .Z(n5322) );
  AND U9191 ( .A(n5323), .B(n5322), .Z(n21002) );
  NANDN U9192 ( .A(n5324), .B(n21002), .Z(n5325) );
  NANDN U9193 ( .A(n21004), .B(n5325), .Z(n5328) );
  NANDN U9194 ( .A(y[628]), .B(x[628]), .Z(n5327) );
  NANDN U9195 ( .A(y[629]), .B(x[629]), .Z(n5326) );
  AND U9196 ( .A(n5327), .B(n5326), .Z(n21006) );
  NAND U9197 ( .A(n5328), .B(n21006), .Z(n5329) );
  NANDN U9198 ( .A(n21009), .B(n5329), .Z(n5332) );
  NANDN U9199 ( .A(y[630]), .B(x[630]), .Z(n5331) );
  NANDN U9200 ( .A(y[631]), .B(x[631]), .Z(n5330) );
  AND U9201 ( .A(n5331), .B(n5330), .Z(n21010) );
  NAND U9202 ( .A(n5332), .B(n21010), .Z(n5335) );
  NANDN U9203 ( .A(x[632]), .B(y[632]), .Z(n5333) );
  NANDN U9204 ( .A(n5334), .B(n5333), .Z(n13805) );
  NANDN U9205 ( .A(x[631]), .B(y[631]), .Z(n13800) );
  NANDN U9206 ( .A(n13805), .B(n13800), .Z(n21013) );
  ANDN U9207 ( .B(n5335), .A(n21013), .Z(n5336) );
  OR U9208 ( .A(n21017), .B(n5336), .Z(n5337) );
  NANDN U9209 ( .A(n21019), .B(n5337), .Z(n5338) );
  NANDN U9210 ( .A(n13810), .B(n5338), .Z(n5339) );
  NANDN U9211 ( .A(x[636]), .B(y[636]), .Z(n21023) );
  NAND U9212 ( .A(n5339), .B(n21023), .Z(n5342) );
  NANDN U9213 ( .A(y[636]), .B(x[636]), .Z(n5341) );
  NANDN U9214 ( .A(y[637]), .B(x[637]), .Z(n5340) );
  AND U9215 ( .A(n5341), .B(n5340), .Z(n21024) );
  NAND U9216 ( .A(n5342), .B(n21024), .Z(n5345) );
  NANDN U9217 ( .A(x[638]), .B(y[638]), .Z(n5344) );
  NANDN U9218 ( .A(x[637]), .B(y[637]), .Z(n5343) );
  NAND U9219 ( .A(n5344), .B(n5343), .Z(n21027) );
  ANDN U9220 ( .B(n5345), .A(n21027), .Z(n5348) );
  NANDN U9221 ( .A(y[638]), .B(x[638]), .Z(n5347) );
  NANDN U9222 ( .A(y[639]), .B(x[639]), .Z(n5346) );
  AND U9223 ( .A(n5347), .B(n5346), .Z(n21028) );
  NANDN U9224 ( .A(n5348), .B(n21028), .Z(n5349) );
  NANDN U9225 ( .A(n21031), .B(n5349), .Z(n5352) );
  NANDN U9226 ( .A(y[640]), .B(x[640]), .Z(n5351) );
  NANDN U9227 ( .A(y[641]), .B(x[641]), .Z(n5350) );
  AND U9228 ( .A(n5351), .B(n5350), .Z(n21032) );
  NAND U9229 ( .A(n5352), .B(n21032), .Z(n5353) );
  NANDN U9230 ( .A(n21034), .B(n5353), .Z(n5356) );
  NANDN U9231 ( .A(y[643]), .B(x[643]), .Z(n5355) );
  NANDN U9232 ( .A(y[642]), .B(x[642]), .Z(n5354) );
  AND U9233 ( .A(n5355), .B(n5354), .Z(n21036) );
  NAND U9234 ( .A(n5356), .B(n21036), .Z(n5357) );
  ANDN U9235 ( .B(y[644]), .A(x[644]), .Z(n13821) );
  ANDN U9236 ( .B(n5357), .A(n13821), .Z(n5358) );
  NANDN U9237 ( .A(x[643]), .B(y[643]), .Z(n21039) );
  NAND U9238 ( .A(n5358), .B(n21039), .Z(n5360) );
  NANDN U9239 ( .A(y[644]), .B(x[644]), .Z(n5359) );
  ANDN U9240 ( .B(x[645]), .A(y[645]), .Z(n13822) );
  ANDN U9241 ( .B(n5359), .A(n13822), .Z(n21040) );
  NAND U9242 ( .A(n5360), .B(n21040), .Z(n5361) );
  ANDN U9243 ( .B(y[645]), .A(x[645]), .Z(n13824) );
  ANDN U9244 ( .B(n5361), .A(n13824), .Z(n5362) );
  NANDN U9245 ( .A(n12743), .B(n5362), .Z(n5363) );
  AND U9246 ( .A(n21044), .B(n5363), .Z(n5364) );
  OR U9247 ( .A(n12746), .B(n5364), .Z(n5365) );
  NANDN U9248 ( .A(n21049), .B(n5365), .Z(n5370) );
  NANDN U9249 ( .A(x[650]), .B(y[650]), .Z(n5367) );
  NANDN U9250 ( .A(x[649]), .B(y[649]), .Z(n5366) );
  AND U9251 ( .A(n5367), .B(n5366), .Z(n5369) );
  AND U9252 ( .A(n5369), .B(n5368), .Z(n21050) );
  NAND U9253 ( .A(n5370), .B(n21050), .Z(n5371) );
  NANDN U9254 ( .A(n21053), .B(n5371), .Z(n5372) );
  NANDN U9255 ( .A(x[652]), .B(y[652]), .Z(n21054) );
  NAND U9256 ( .A(n5372), .B(n21054), .Z(n5375) );
  NANDN U9257 ( .A(y[653]), .B(x[653]), .Z(n5374) );
  NANDN U9258 ( .A(y[652]), .B(x[652]), .Z(n5373) );
  NAND U9259 ( .A(n5374), .B(n5373), .Z(n21056) );
  ANDN U9260 ( .B(n5375), .A(n21056), .Z(n5378) );
  NANDN U9261 ( .A(x[653]), .B(y[653]), .Z(n5377) );
  NANDN U9262 ( .A(x[654]), .B(y[654]), .Z(n5376) );
  AND U9263 ( .A(n5377), .B(n5376), .Z(n21058) );
  NANDN U9264 ( .A(n5378), .B(n21058), .Z(n5379) );
  NANDN U9265 ( .A(n21061), .B(n5379), .Z(n5382) );
  NANDN U9266 ( .A(x[655]), .B(y[655]), .Z(n5381) );
  NANDN U9267 ( .A(x[656]), .B(y[656]), .Z(n5380) );
  AND U9268 ( .A(n5381), .B(n5380), .Z(n21062) );
  NAND U9269 ( .A(n5382), .B(n21062), .Z(n5383) );
  NANDN U9270 ( .A(n21065), .B(n5383), .Z(n5386) );
  NANDN U9271 ( .A(x[657]), .B(y[657]), .Z(n5385) );
  NANDN U9272 ( .A(x[658]), .B(y[658]), .Z(n5384) );
  AND U9273 ( .A(n5385), .B(n5384), .Z(n21066) );
  NAND U9274 ( .A(n5386), .B(n21066), .Z(n5389) );
  NANDN U9275 ( .A(y[659]), .B(x[659]), .Z(n5388) );
  NANDN U9276 ( .A(y[658]), .B(x[658]), .Z(n5387) );
  NAND U9277 ( .A(n5388), .B(n5387), .Z(n21068) );
  ANDN U9278 ( .B(n5389), .A(n21068), .Z(n5392) );
  NANDN U9279 ( .A(x[659]), .B(y[659]), .Z(n5391) );
  NANDN U9280 ( .A(x[660]), .B(y[660]), .Z(n5390) );
  AND U9281 ( .A(n5391), .B(n5390), .Z(n21070) );
  NANDN U9282 ( .A(n5392), .B(n21070), .Z(n5393) );
  NANDN U9283 ( .A(n21073), .B(n5393), .Z(n5394) );
  NANDN U9284 ( .A(x[661]), .B(y[661]), .Z(n21074) );
  NAND U9285 ( .A(n5394), .B(n21074), .Z(n5395) );
  OR U9286 ( .A(n13843), .B(n5395), .Z(n5397) );
  NANDN U9287 ( .A(y[662]), .B(x[662]), .Z(n5396) );
  ANDN U9288 ( .B(x[663]), .A(y[663]), .Z(n13844) );
  ANDN U9289 ( .B(n5396), .A(n13844), .Z(n21076) );
  NAND U9290 ( .A(n5397), .B(n21076), .Z(n5398) );
  NANDN U9291 ( .A(n13846), .B(n5398), .Z(n5399) );
  NANDN U9292 ( .A(n21080), .B(n5399), .Z(n5402) );
  NANDN U9293 ( .A(x[665]), .B(y[665]), .Z(n5401) );
  NANDN U9294 ( .A(x[666]), .B(y[666]), .Z(n5400) );
  AND U9295 ( .A(n5401), .B(n5400), .Z(n21082) );
  NAND U9296 ( .A(n5402), .B(n21082), .Z(n5405) );
  NANDN U9297 ( .A(y[667]), .B(x[667]), .Z(n5404) );
  NANDN U9298 ( .A(y[666]), .B(x[666]), .Z(n5403) );
  NAND U9299 ( .A(n5404), .B(n5403), .Z(n21085) );
  ANDN U9300 ( .B(n5405), .A(n21085), .Z(n5408) );
  NANDN U9301 ( .A(x[667]), .B(y[667]), .Z(n5407) );
  NANDN U9302 ( .A(x[668]), .B(y[668]), .Z(n5406) );
  AND U9303 ( .A(n5407), .B(n5406), .Z(n21086) );
  NANDN U9304 ( .A(n5408), .B(n21086), .Z(n5411) );
  NANDN U9305 ( .A(y[669]), .B(x[669]), .Z(n5410) );
  NANDN U9306 ( .A(y[668]), .B(x[668]), .Z(n5409) );
  NAND U9307 ( .A(n5410), .B(n5409), .Z(n21089) );
  ANDN U9308 ( .B(n5411), .A(n21089), .Z(n5414) );
  NANDN U9309 ( .A(x[669]), .B(y[669]), .Z(n5413) );
  NANDN U9310 ( .A(x[670]), .B(y[670]), .Z(n5412) );
  AND U9311 ( .A(n5413), .B(n5412), .Z(n21090) );
  NANDN U9312 ( .A(n5414), .B(n21090), .Z(n5415) );
  NANDN U9313 ( .A(n21092), .B(n5415), .Z(n5416) );
  NANDN U9314 ( .A(x[671]), .B(y[671]), .Z(n21094) );
  NAND U9315 ( .A(n5416), .B(n21094), .Z(n5417) );
  NANDN U9316 ( .A(y[672]), .B(x[672]), .Z(n21096) );
  NAND U9317 ( .A(n5417), .B(n21096), .Z(n5418) );
  NANDN U9318 ( .A(n21098), .B(n5418), .Z(n5419) );
  AND U9319 ( .A(n21101), .B(n5419), .Z(n5420) );
  NANDN U9320 ( .A(x[674]), .B(y[674]), .Z(n21104) );
  NANDN U9321 ( .A(n5420), .B(n21104), .Z(n5421) );
  NANDN U9322 ( .A(n13864), .B(n5421), .Z(n5422) );
  NANDN U9323 ( .A(n13866), .B(n5422), .Z(n5423) );
  NANDN U9324 ( .A(n13868), .B(n5423), .Z(n5426) );
  NANDN U9325 ( .A(x[677]), .B(y[677]), .Z(n5425) );
  NANDN U9326 ( .A(x[678]), .B(y[678]), .Z(n5424) );
  AND U9327 ( .A(n5425), .B(n5424), .Z(n21117) );
  NAND U9328 ( .A(n5426), .B(n21117), .Z(n5427) );
  AND U9329 ( .A(n21119), .B(n5427), .Z(n5430) );
  NANDN U9330 ( .A(x[679]), .B(y[679]), .Z(n5429) );
  NANDN U9331 ( .A(x[680]), .B(y[680]), .Z(n5428) );
  AND U9332 ( .A(n5429), .B(n5428), .Z(n21122) );
  NANDN U9333 ( .A(n5430), .B(n21122), .Z(n5433) );
  NANDN U9334 ( .A(y[681]), .B(x[681]), .Z(n5432) );
  NANDN U9335 ( .A(y[680]), .B(x[680]), .Z(n5431) );
  AND U9336 ( .A(n5432), .B(n5431), .Z(n21123) );
  NAND U9337 ( .A(n5433), .B(n21123), .Z(n5436) );
  NANDN U9338 ( .A(x[681]), .B(y[681]), .Z(n5435) );
  NANDN U9339 ( .A(x[682]), .B(y[682]), .Z(n5434) );
  AND U9340 ( .A(n5435), .B(n5434), .Z(n21125) );
  NAND U9341 ( .A(n5436), .B(n21125), .Z(n5439) );
  NANDN U9342 ( .A(y[683]), .B(x[683]), .Z(n5438) );
  NANDN U9343 ( .A(y[682]), .B(x[682]), .Z(n5437) );
  AND U9344 ( .A(n5438), .B(n5437), .Z(n21127) );
  NAND U9345 ( .A(n5439), .B(n21127), .Z(n5444) );
  NANDN U9346 ( .A(x[684]), .B(y[684]), .Z(n5441) );
  NANDN U9347 ( .A(x[683]), .B(y[683]), .Z(n5440) );
  AND U9348 ( .A(n5441), .B(n5440), .Z(n5443) );
  AND U9349 ( .A(n5443), .B(n5442), .Z(n21129) );
  NAND U9350 ( .A(n5444), .B(n21129), .Z(n5445) );
  AND U9351 ( .A(n21131), .B(n5445), .Z(n5452) );
  NANDN U9352 ( .A(x[687]), .B(y[687]), .Z(n5447) );
  ANDN U9353 ( .B(y[688]), .A(x[688]), .Z(n5446) );
  ANDN U9354 ( .B(n5447), .A(n5446), .Z(n5451) );
  XNOR U9355 ( .A(y[687]), .B(x[687]), .Z(n5449) );
  ANDN U9356 ( .B(y[686]), .A(x[686]), .Z(n5448) );
  NAND U9357 ( .A(n5449), .B(n5448), .Z(n5450) );
  AND U9358 ( .A(n5451), .B(n5450), .Z(n21134) );
  NANDN U9359 ( .A(n5452), .B(n21134), .Z(n5455) );
  NANDN U9360 ( .A(y[689]), .B(x[689]), .Z(n5454) );
  NANDN U9361 ( .A(y[688]), .B(x[688]), .Z(n5453) );
  AND U9362 ( .A(n5454), .B(n5453), .Z(n21135) );
  NAND U9363 ( .A(n5455), .B(n21135), .Z(n5458) );
  NANDN U9364 ( .A(x[689]), .B(y[689]), .Z(n5457) );
  NANDN U9365 ( .A(x[690]), .B(y[690]), .Z(n5456) );
  AND U9366 ( .A(n5457), .B(n5456), .Z(n21137) );
  NAND U9367 ( .A(n5458), .B(n21137), .Z(n5461) );
  NANDN U9368 ( .A(y[691]), .B(x[691]), .Z(n5460) );
  NANDN U9369 ( .A(y[690]), .B(x[690]), .Z(n5459) );
  AND U9370 ( .A(n5460), .B(n5459), .Z(n21139) );
  NAND U9371 ( .A(n5461), .B(n21139), .Z(n5464) );
  NANDN U9372 ( .A(x[691]), .B(y[691]), .Z(n5463) );
  NANDN U9373 ( .A(x[692]), .B(y[692]), .Z(n5462) );
  AND U9374 ( .A(n5463), .B(n5462), .Z(n21141) );
  NAND U9375 ( .A(n5464), .B(n21141), .Z(n5465) );
  AND U9376 ( .A(n21143), .B(n5465), .Z(n5466) );
  NANDN U9377 ( .A(x[694]), .B(y[694]), .Z(n20300) );
  ANDN U9378 ( .B(y[693]), .A(x[693]), .Z(n21145) );
  ANDN U9379 ( .B(n20300), .A(n21145), .Z(n13883) );
  NANDN U9380 ( .A(n5466), .B(n13883), .Z(n5468) );
  NANDN U9381 ( .A(y[694]), .B(x[694]), .Z(n5467) );
  NANDN U9382 ( .A(y[695]), .B(x[695]), .Z(n20302) );
  AND U9383 ( .A(n5467), .B(n20302), .Z(n21147) );
  NAND U9384 ( .A(n5468), .B(n21147), .Z(n5469) );
  NANDN U9385 ( .A(n12739), .B(n5469), .Z(n5470) );
  NANDN U9386 ( .A(x[695]), .B(y[695]), .Z(n20299) );
  NANDN U9387 ( .A(n5470), .B(n20299), .Z(n5472) );
  NANDN U9388 ( .A(y[696]), .B(x[696]), .Z(n5471) );
  ANDN U9389 ( .B(x[697]), .A(y[697]), .Z(n12740) );
  ANDN U9390 ( .B(n5471), .A(n12740), .Z(n21151) );
  NAND U9391 ( .A(n5472), .B(n21151), .Z(n5473) );
  NANDN U9392 ( .A(n12742), .B(n5473), .Z(n5474) );
  NANDN U9393 ( .A(n21156), .B(n5474), .Z(n5477) );
  NANDN U9394 ( .A(x[699]), .B(y[699]), .Z(n5476) );
  NANDN U9395 ( .A(x[700]), .B(y[700]), .Z(n5475) );
  AND U9396 ( .A(n5476), .B(n5475), .Z(n21157) );
  NAND U9397 ( .A(n5477), .B(n21157), .Z(n5480) );
  NANDN U9398 ( .A(y[701]), .B(x[701]), .Z(n5479) );
  NANDN U9399 ( .A(y[700]), .B(x[700]), .Z(n5478) );
  NAND U9400 ( .A(n5479), .B(n5478), .Z(n21160) );
  ANDN U9401 ( .B(n5480), .A(n21160), .Z(n5483) );
  NANDN U9402 ( .A(x[701]), .B(y[701]), .Z(n5482) );
  NANDN U9403 ( .A(x[702]), .B(y[702]), .Z(n5481) );
  AND U9404 ( .A(n5482), .B(n5481), .Z(n21161) );
  NANDN U9405 ( .A(n5483), .B(n21161), .Z(n5484) );
  NANDN U9406 ( .A(n21163), .B(n5484), .Z(n5489) );
  NANDN U9407 ( .A(x[704]), .B(y[704]), .Z(n5486) );
  NANDN U9408 ( .A(x[703]), .B(y[703]), .Z(n5485) );
  AND U9409 ( .A(n5486), .B(n5485), .Z(n5488) );
  AND U9410 ( .A(n5488), .B(n5487), .Z(n21165) );
  NAND U9411 ( .A(n5489), .B(n21165), .Z(n5490) );
  NANDN U9412 ( .A(n21168), .B(n5490), .Z(n5491) );
  NANDN U9413 ( .A(x[706]), .B(y[706]), .Z(n21169) );
  NAND U9414 ( .A(n5491), .B(n21169), .Z(n5494) );
  NANDN U9415 ( .A(y[707]), .B(x[707]), .Z(n5493) );
  NANDN U9416 ( .A(y[706]), .B(x[706]), .Z(n5492) );
  NAND U9417 ( .A(n5493), .B(n5492), .Z(n21172) );
  ANDN U9418 ( .B(n5494), .A(n21172), .Z(n5497) );
  NANDN U9419 ( .A(x[707]), .B(y[707]), .Z(n5496) );
  NANDN U9420 ( .A(x[708]), .B(y[708]), .Z(n5495) );
  AND U9421 ( .A(n5496), .B(n5495), .Z(n21173) );
  NANDN U9422 ( .A(n5497), .B(n21173), .Z(n5498) );
  NANDN U9423 ( .A(n21175), .B(n5498), .Z(n5501) );
  NANDN U9424 ( .A(x[709]), .B(y[709]), .Z(n5500) );
  NANDN U9425 ( .A(x[710]), .B(y[710]), .Z(n5499) );
  AND U9426 ( .A(n5500), .B(n5499), .Z(n21177) );
  NAND U9427 ( .A(n5501), .B(n21177), .Z(n5502) );
  NANDN U9428 ( .A(n21180), .B(n5502), .Z(n5503) );
  ANDN U9429 ( .B(y[712]), .A(x[712]), .Z(n13904) );
  ANDN U9430 ( .B(n5503), .A(n13904), .Z(n5504) );
  NANDN U9431 ( .A(x[711]), .B(y[711]), .Z(n21181) );
  NAND U9432 ( .A(n5504), .B(n21181), .Z(n5506) );
  NANDN U9433 ( .A(y[712]), .B(x[712]), .Z(n5505) );
  ANDN U9434 ( .B(x[713]), .A(y[713]), .Z(n13905) );
  ANDN U9435 ( .B(n5505), .A(n13905), .Z(n21183) );
  NAND U9436 ( .A(n5506), .B(n21183), .Z(n5507) );
  NANDN U9437 ( .A(n13907), .B(n5507), .Z(n5510) );
  NANDN U9438 ( .A(y[715]), .B(x[715]), .Z(n5509) );
  NANDN U9439 ( .A(y[714]), .B(x[714]), .Z(n5508) );
  NAND U9440 ( .A(n5509), .B(n5508), .Z(n21187) );
  ANDN U9441 ( .B(n5510), .A(n21187), .Z(n5513) );
  NANDN U9442 ( .A(x[715]), .B(y[715]), .Z(n5512) );
  NANDN U9443 ( .A(x[716]), .B(y[716]), .Z(n5511) );
  AND U9444 ( .A(n5512), .B(n5511), .Z(n21189) );
  NANDN U9445 ( .A(n5513), .B(n21189), .Z(n5514) );
  NANDN U9446 ( .A(n21192), .B(n5514), .Z(n5519) );
  NANDN U9447 ( .A(x[718]), .B(y[718]), .Z(n5516) );
  NANDN U9448 ( .A(x[717]), .B(y[717]), .Z(n5515) );
  AND U9449 ( .A(n5516), .B(n5515), .Z(n5518) );
  AND U9450 ( .A(n5518), .B(n5517), .Z(n21193) );
  NAND U9451 ( .A(n5519), .B(n21193), .Z(n5520) );
  NANDN U9452 ( .A(n21196), .B(n5520), .Z(n5521) );
  NANDN U9453 ( .A(x[720]), .B(y[720]), .Z(n21197) );
  NAND U9454 ( .A(n5521), .B(n21197), .Z(n5524) );
  NANDN U9455 ( .A(y[721]), .B(x[721]), .Z(n5523) );
  NANDN U9456 ( .A(y[720]), .B(x[720]), .Z(n5522) );
  NAND U9457 ( .A(n5523), .B(n5522), .Z(n21199) );
  ANDN U9458 ( .B(n5524), .A(n21199), .Z(n5527) );
  NANDN U9459 ( .A(x[721]), .B(y[721]), .Z(n5526) );
  NANDN U9460 ( .A(x[722]), .B(y[722]), .Z(n5525) );
  AND U9461 ( .A(n5526), .B(n5525), .Z(n21201) );
  NANDN U9462 ( .A(n5527), .B(n21201), .Z(n5528) );
  NANDN U9463 ( .A(n21204), .B(n5528), .Z(n5531) );
  NANDN U9464 ( .A(x[723]), .B(y[723]), .Z(n5530) );
  NANDN U9465 ( .A(x[724]), .B(y[724]), .Z(n5529) );
  AND U9466 ( .A(n5530), .B(n5529), .Z(n21205) );
  NAND U9467 ( .A(n5531), .B(n21205), .Z(n5532) );
  NANDN U9468 ( .A(n21208), .B(n5532), .Z(n5535) );
  NANDN U9469 ( .A(x[725]), .B(y[725]), .Z(n5534) );
  NANDN U9470 ( .A(x[726]), .B(y[726]), .Z(n5533) );
  AND U9471 ( .A(n5534), .B(n5533), .Z(n21209) );
  NAND U9472 ( .A(n5535), .B(n21209), .Z(n5538) );
  NANDN U9473 ( .A(y[727]), .B(x[727]), .Z(n5537) );
  NANDN U9474 ( .A(y[726]), .B(x[726]), .Z(n5536) );
  NAND U9475 ( .A(n5537), .B(n5536), .Z(n21211) );
  ANDN U9476 ( .B(n5538), .A(n21211), .Z(n5541) );
  NANDN U9477 ( .A(x[727]), .B(y[727]), .Z(n5540) );
  NANDN U9478 ( .A(x[728]), .B(y[728]), .Z(n5539) );
  AND U9479 ( .A(n5540), .B(n5539), .Z(n21213) );
  NANDN U9480 ( .A(n5541), .B(n21213), .Z(n5542) );
  NANDN U9481 ( .A(n21216), .B(n5542), .Z(n5545) );
  NANDN U9482 ( .A(x[729]), .B(y[729]), .Z(n5544) );
  NANDN U9483 ( .A(x[730]), .B(y[730]), .Z(n5543) );
  AND U9484 ( .A(n5544), .B(n5543), .Z(n21217) );
  NAND U9485 ( .A(n5545), .B(n21217), .Z(n5546) );
  NANDN U9486 ( .A(n21220), .B(n5546), .Z(n5547) );
  ANDN U9487 ( .B(y[732]), .A(x[732]), .Z(n12733) );
  ANDN U9488 ( .B(n5547), .A(n12733), .Z(n5548) );
  NANDN U9489 ( .A(x[731]), .B(y[731]), .Z(n21221) );
  NAND U9490 ( .A(n5548), .B(n21221), .Z(n5550) );
  NANDN U9491 ( .A(y[732]), .B(x[732]), .Z(n5549) );
  NANDN U9492 ( .A(y[733]), .B(x[733]), .Z(n12735) );
  AND U9493 ( .A(n5549), .B(n12735), .Z(n21224) );
  NAND U9494 ( .A(n5550), .B(n21224), .Z(n5551) );
  ANDN U9495 ( .B(y[734]), .A(x[734]), .Z(n12738) );
  ANDN U9496 ( .B(n5551), .A(n12738), .Z(n5552) );
  NANDN U9497 ( .A(n12734), .B(n5552), .Z(n5553) );
  NANDN U9498 ( .A(n21228), .B(n5553), .Z(n5558) );
  NANDN U9499 ( .A(x[736]), .B(y[736]), .Z(n5555) );
  NANDN U9500 ( .A(x[735]), .B(y[735]), .Z(n5554) );
  AND U9501 ( .A(n5555), .B(n5554), .Z(n5557) );
  NANDN U9502 ( .A(x[737]), .B(y[737]), .Z(n5556) );
  AND U9503 ( .A(n5557), .B(n5556), .Z(n21229) );
  NAND U9504 ( .A(n5558), .B(n21229), .Z(n5559) );
  NANDN U9505 ( .A(n21232), .B(n5559), .Z(n5566) );
  NANDN U9506 ( .A(x[740]), .B(y[740]), .Z(n5565) );
  ANDN U9507 ( .B(y[738]), .A(x[738]), .Z(n5560) );
  OR U9508 ( .A(n5560), .B(y[739]), .Z(n5563) );
  XOR U9509 ( .A(y[739]), .B(n5560), .Z(n5561) );
  NAND U9510 ( .A(n5561), .B(x[739]), .Z(n5562) );
  NAND U9511 ( .A(n5563), .B(n5562), .Z(n5564) );
  AND U9512 ( .A(n5565), .B(n5564), .Z(n21233) );
  NAND U9513 ( .A(n5566), .B(n21233), .Z(n5569) );
  NANDN U9514 ( .A(y[740]), .B(x[740]), .Z(n5568) );
  NANDN U9515 ( .A(y[741]), .B(x[741]), .Z(n5567) );
  AND U9516 ( .A(n5568), .B(n5567), .Z(n21236) );
  NAND U9517 ( .A(n5569), .B(n21236), .Z(n5570) );
  AND U9518 ( .A(n21237), .B(n5570), .Z(n5575) );
  NANDN U9519 ( .A(y[742]), .B(x[742]), .Z(n5571) );
  NANDN U9520 ( .A(n5571), .B(x[743]), .Z(n5574) );
  XNOR U9521 ( .A(n5571), .B(x[743]), .Z(n5572) );
  NANDN U9522 ( .A(y[743]), .B(n5572), .Z(n5573) );
  AND U9523 ( .A(n5574), .B(n5573), .Z(n21239) );
  NANDN U9524 ( .A(n5575), .B(n21239), .Z(n5576) );
  NANDN U9525 ( .A(x[744]), .B(y[744]), .Z(n21241) );
  NAND U9526 ( .A(n5576), .B(n21241), .Z(n5579) );
  NANDN U9527 ( .A(y[744]), .B(x[744]), .Z(n5578) );
  NANDN U9528 ( .A(y[745]), .B(x[745]), .Z(n5577) );
  AND U9529 ( .A(n5578), .B(n5577), .Z(n21243) );
  NAND U9530 ( .A(n5579), .B(n21243), .Z(n5582) );
  NANDN U9531 ( .A(x[746]), .B(y[746]), .Z(n5581) );
  NANDN U9532 ( .A(x[745]), .B(y[745]), .Z(n5580) );
  AND U9533 ( .A(n5581), .B(n5580), .Z(n21245) );
  NAND U9534 ( .A(n5582), .B(n21245), .Z(n5585) );
  NANDN U9535 ( .A(y[746]), .B(x[746]), .Z(n5584) );
  NANDN U9536 ( .A(y[747]), .B(x[747]), .Z(n5583) );
  AND U9537 ( .A(n5584), .B(n5583), .Z(n21248) );
  NAND U9538 ( .A(n5585), .B(n21248), .Z(n5586) );
  AND U9539 ( .A(n21249), .B(n5586), .Z(n5589) );
  NANDN U9540 ( .A(y[748]), .B(x[748]), .Z(n5588) );
  NANDN U9541 ( .A(y[749]), .B(x[749]), .Z(n5587) );
  AND U9542 ( .A(n5588), .B(n5587), .Z(n21251) );
  NANDN U9543 ( .A(n5589), .B(n21251), .Z(n5591) );
  ANDN U9544 ( .B(y[749]), .A(x[749]), .Z(n13943) );
  ANDN U9545 ( .B(n13946), .A(n13943), .Z(n21253) );
  NAND U9546 ( .A(n5591), .B(n21253), .Z(n5592) );
  NANDN U9547 ( .A(n21255), .B(n5592), .Z(n5593) );
  NANDN U9548 ( .A(n21260), .B(n5593), .Z(n5599) );
  NANDN U9549 ( .A(y[753]), .B(x[753]), .Z(n21264) );
  NANDN U9550 ( .A(y[752]), .B(x[752]), .Z(n21257) );
  NAND U9551 ( .A(n21264), .B(n21257), .Z(n5594) );
  NANDN U9552 ( .A(n5595), .B(n5594), .Z(n5598) );
  NANDN U9553 ( .A(y[754]), .B(x[754]), .Z(n5597) );
  NANDN U9554 ( .A(y[755]), .B(x[755]), .Z(n5596) );
  NAND U9555 ( .A(n5597), .B(n5596), .Z(n21261) );
  ANDN U9556 ( .B(n5598), .A(n21261), .Z(n13951) );
  NAND U9557 ( .A(n5599), .B(n13951), .Z(n5600) );
  AND U9558 ( .A(n21267), .B(n5600), .Z(n5603) );
  NANDN U9559 ( .A(y[756]), .B(x[756]), .Z(n5602) );
  NANDN U9560 ( .A(y[757]), .B(x[757]), .Z(n5601) );
  AND U9561 ( .A(n5602), .B(n5601), .Z(n21269) );
  NANDN U9562 ( .A(n5603), .B(n21269), .Z(n5606) );
  NANDN U9563 ( .A(x[758]), .B(y[758]), .Z(n5605) );
  NANDN U9564 ( .A(x[757]), .B(y[757]), .Z(n5604) );
  AND U9565 ( .A(n5605), .B(n5604), .Z(n21271) );
  NAND U9566 ( .A(n5606), .B(n21271), .Z(n5609) );
  NANDN U9567 ( .A(y[758]), .B(x[758]), .Z(n5608) );
  NANDN U9568 ( .A(y[759]), .B(x[759]), .Z(n5607) );
  AND U9569 ( .A(n5608), .B(n5607), .Z(n21273) );
  NAND U9570 ( .A(n5609), .B(n21273), .Z(n5612) );
  NANDN U9571 ( .A(x[760]), .B(y[760]), .Z(n5611) );
  NANDN U9572 ( .A(x[759]), .B(y[759]), .Z(n5610) );
  AND U9573 ( .A(n5611), .B(n5610), .Z(n21275) );
  NAND U9574 ( .A(n5612), .B(n21275), .Z(n5615) );
  NANDN U9575 ( .A(y[760]), .B(x[760]), .Z(n5614) );
  NANDN U9576 ( .A(y[761]), .B(x[761]), .Z(n5613) );
  AND U9577 ( .A(n5614), .B(n5613), .Z(n21278) );
  NAND U9578 ( .A(n5615), .B(n21278), .Z(n5616) );
  AND U9579 ( .A(n21279), .B(n5616), .Z(n5619) );
  NANDN U9580 ( .A(y[762]), .B(x[762]), .Z(n5618) );
  NANDN U9581 ( .A(y[763]), .B(x[763]), .Z(n5617) );
  AND U9582 ( .A(n5618), .B(n5617), .Z(n21281) );
  NANDN U9583 ( .A(n5619), .B(n21281), .Z(n5620) );
  AND U9584 ( .A(n21283), .B(n5620), .Z(n5623) );
  NANDN U9585 ( .A(y[764]), .B(x[764]), .Z(n5622) );
  NANDN U9586 ( .A(y[765]), .B(x[765]), .Z(n5621) );
  AND U9587 ( .A(n5622), .B(n5621), .Z(n21285) );
  NANDN U9588 ( .A(n5623), .B(n21285), .Z(n5625) );
  NANDN U9589 ( .A(x[766]), .B(y[766]), .Z(n5624) );
  ANDN U9590 ( .B(y[765]), .A(x[765]), .Z(n13963) );
  ANDN U9591 ( .B(n5624), .A(n13963), .Z(n21287) );
  NAND U9592 ( .A(n5625), .B(n21287), .Z(n5626) );
  NANDN U9593 ( .A(n21289), .B(n5626), .Z(n5629) );
  NANDN U9594 ( .A(x[768]), .B(y[768]), .Z(n5628) );
  NANDN U9595 ( .A(x[767]), .B(y[767]), .Z(n5627) );
  AND U9596 ( .A(n5628), .B(n5627), .Z(n21291) );
  NAND U9597 ( .A(n5629), .B(n21291), .Z(n5632) );
  NANDN U9598 ( .A(y[768]), .B(x[768]), .Z(n5631) );
  NANDN U9599 ( .A(y[769]), .B(x[769]), .Z(n5630) );
  AND U9600 ( .A(n5631), .B(n5630), .Z(n21293) );
  NAND U9601 ( .A(n5632), .B(n21293), .Z(n5633) );
  AND U9602 ( .A(n21295), .B(n5633), .Z(n5636) );
  NANDN U9603 ( .A(y[770]), .B(x[770]), .Z(n5635) );
  NANDN U9604 ( .A(y[771]), .B(x[771]), .Z(n5634) );
  AND U9605 ( .A(n5635), .B(n5634), .Z(n21297) );
  NANDN U9606 ( .A(n5636), .B(n21297), .Z(n5639) );
  NANDN U9607 ( .A(x[772]), .B(y[772]), .Z(n5638) );
  NANDN U9608 ( .A(x[771]), .B(y[771]), .Z(n5637) );
  AND U9609 ( .A(n5638), .B(n5637), .Z(n21299) );
  NAND U9610 ( .A(n5639), .B(n21299), .Z(n5642) );
  NANDN U9611 ( .A(y[773]), .B(x[773]), .Z(n5641) );
  NANDN U9612 ( .A(y[772]), .B(x[772]), .Z(n5640) );
  AND U9613 ( .A(n5641), .B(n5640), .Z(n21302) );
  NAND U9614 ( .A(n5642), .B(n21302), .Z(n5643) );
  NANDN U9615 ( .A(x[773]), .B(y[773]), .Z(n21303) );
  NAND U9616 ( .A(n5643), .B(n21303), .Z(n5645) );
  IV U9617 ( .A(x[774]), .Z(n13977) );
  AND U9618 ( .A(y[774]), .B(n13977), .Z(n5644) );
  OR U9619 ( .A(n5645), .B(n5644), .Z(n5646) );
  NANDN U9620 ( .A(n21305), .B(n5646), .Z(n5647) );
  NANDN U9621 ( .A(n13978), .B(n5647), .Z(n5648) );
  OR U9622 ( .A(n13983), .B(n5648), .Z(n5651) );
  NANDN U9623 ( .A(y[777]), .B(x[777]), .Z(n5650) );
  NANDN U9624 ( .A(y[776]), .B(x[776]), .Z(n5649) );
  AND U9625 ( .A(n5650), .B(n5649), .Z(n21309) );
  NAND U9626 ( .A(n5651), .B(n21309), .Z(n5654) );
  NANDN U9627 ( .A(x[777]), .B(y[777]), .Z(n5653) );
  NANDN U9628 ( .A(x[778]), .B(y[778]), .Z(n5652) );
  AND U9629 ( .A(n5653), .B(n5652), .Z(n21312) );
  NAND U9630 ( .A(n5654), .B(n21312), .Z(n5657) );
  NANDN U9631 ( .A(y[779]), .B(x[779]), .Z(n5656) );
  NANDN U9632 ( .A(y[778]), .B(x[778]), .Z(n5655) );
  AND U9633 ( .A(n5656), .B(n5655), .Z(n21313) );
  NAND U9634 ( .A(n5657), .B(n21313), .Z(n5660) );
  NANDN U9635 ( .A(x[779]), .B(y[779]), .Z(n5659) );
  NANDN U9636 ( .A(x[780]), .B(y[780]), .Z(n5658) );
  AND U9637 ( .A(n5659), .B(n5658), .Z(n21315) );
  NAND U9638 ( .A(n5660), .B(n21315), .Z(n5661) );
  AND U9639 ( .A(n21317), .B(n5661), .Z(n5664) );
  NANDN U9640 ( .A(x[781]), .B(y[781]), .Z(n5663) );
  NANDN U9641 ( .A(x[782]), .B(y[782]), .Z(n5662) );
  AND U9642 ( .A(n5663), .B(n5662), .Z(n21319) );
  NANDN U9643 ( .A(n5664), .B(n21319), .Z(n5667) );
  NANDN U9644 ( .A(y[783]), .B(x[783]), .Z(n5666) );
  NANDN U9645 ( .A(y[782]), .B(x[782]), .Z(n5665) );
  AND U9646 ( .A(n5666), .B(n5665), .Z(n21321) );
  NAND U9647 ( .A(n5667), .B(n21321), .Z(n5670) );
  NANDN U9648 ( .A(x[783]), .B(y[783]), .Z(n5669) );
  NANDN U9649 ( .A(x[784]), .B(y[784]), .Z(n5668) );
  AND U9650 ( .A(n5669), .B(n5668), .Z(n21324) );
  NAND U9651 ( .A(n5670), .B(n21324), .Z(n5673) );
  NANDN U9652 ( .A(y[785]), .B(x[785]), .Z(n5672) );
  NANDN U9653 ( .A(y[784]), .B(x[784]), .Z(n5671) );
  AND U9654 ( .A(n5672), .B(n5671), .Z(n21325) );
  NAND U9655 ( .A(n5673), .B(n21325), .Z(n5676) );
  NANDN U9656 ( .A(x[785]), .B(y[785]), .Z(n5675) );
  NANDN U9657 ( .A(x[786]), .B(y[786]), .Z(n5674) );
  AND U9658 ( .A(n5675), .B(n5674), .Z(n21327) );
  NAND U9659 ( .A(n5676), .B(n21327), .Z(n5677) );
  AND U9660 ( .A(n21329), .B(n5677), .Z(n5681) );
  NANDN U9661 ( .A(x[788]), .B(y[788]), .Z(n5679) );
  NANDN U9662 ( .A(x[787]), .B(y[787]), .Z(n5678) );
  AND U9663 ( .A(n5679), .B(n5678), .Z(n5680) );
  NANDN U9664 ( .A(x[789]), .B(y[789]), .Z(n5685) );
  AND U9665 ( .A(n5680), .B(n5685), .Z(n21331) );
  NANDN U9666 ( .A(n5681), .B(n21331), .Z(n5686) );
  XNOR U9667 ( .A(x[789]), .B(y[789]), .Z(n5683) );
  NANDN U9668 ( .A(y[788]), .B(x[788]), .Z(n5682) );
  NAND U9669 ( .A(n5683), .B(n5682), .Z(n5684) );
  NAND U9670 ( .A(n5685), .B(n5684), .Z(n21333) );
  NAND U9671 ( .A(n5686), .B(n21333), .Z(n5687) );
  NANDN U9672 ( .A(x[790]), .B(y[790]), .Z(n21336) );
  NAND U9673 ( .A(n5687), .B(n21336), .Z(n5690) );
  NANDN U9674 ( .A(y[791]), .B(x[791]), .Z(n5689) );
  NANDN U9675 ( .A(y[790]), .B(x[790]), .Z(n5688) );
  AND U9676 ( .A(n5689), .B(n5688), .Z(n21337) );
  NAND U9677 ( .A(n5690), .B(n21337), .Z(n5693) );
  NANDN U9678 ( .A(x[791]), .B(y[791]), .Z(n5692) );
  NANDN U9679 ( .A(x[792]), .B(y[792]), .Z(n5691) );
  AND U9680 ( .A(n5692), .B(n5691), .Z(n21339) );
  NAND U9681 ( .A(n5693), .B(n21339), .Z(n5694) );
  AND U9682 ( .A(n21341), .B(n5694), .Z(n5697) );
  NANDN U9683 ( .A(x[793]), .B(y[793]), .Z(n5696) );
  NANDN U9684 ( .A(x[794]), .B(y[794]), .Z(n5695) );
  AND U9685 ( .A(n5696), .B(n5695), .Z(n21343) );
  NANDN U9686 ( .A(n5697), .B(n21343), .Z(n5700) );
  NANDN U9687 ( .A(y[795]), .B(x[795]), .Z(n5699) );
  NANDN U9688 ( .A(y[794]), .B(x[794]), .Z(n5698) );
  AND U9689 ( .A(n5699), .B(n5698), .Z(n21345) );
  NAND U9690 ( .A(n5700), .B(n21345), .Z(n5703) );
  NANDN U9691 ( .A(x[795]), .B(y[795]), .Z(n5702) );
  NANDN U9692 ( .A(x[796]), .B(y[796]), .Z(n5701) );
  AND U9693 ( .A(n5702), .B(n5701), .Z(n21348) );
  NAND U9694 ( .A(n5703), .B(n21348), .Z(n5706) );
  NANDN U9695 ( .A(y[797]), .B(x[797]), .Z(n5705) );
  NANDN U9696 ( .A(y[796]), .B(x[796]), .Z(n5704) );
  AND U9697 ( .A(n5705), .B(n5704), .Z(n21349) );
  NAND U9698 ( .A(n5706), .B(n21349), .Z(n5709) );
  NANDN U9699 ( .A(x[797]), .B(y[797]), .Z(n5708) );
  NANDN U9700 ( .A(x[798]), .B(y[798]), .Z(n5707) );
  AND U9701 ( .A(n5708), .B(n5707), .Z(n21351) );
  NAND U9702 ( .A(n5709), .B(n21351), .Z(n5710) );
  AND U9703 ( .A(n21353), .B(n5710), .Z(n5715) );
  NANDN U9704 ( .A(x[800]), .B(y[800]), .Z(n5712) );
  NANDN U9705 ( .A(x[799]), .B(y[799]), .Z(n5711) );
  AND U9706 ( .A(n5712), .B(n5711), .Z(n5714) );
  NANDN U9707 ( .A(x[801]), .B(y[801]), .Z(n5713) );
  AND U9708 ( .A(n5714), .B(n5713), .Z(n21355) );
  NANDN U9709 ( .A(n5715), .B(n21355), .Z(n5722) );
  NANDN U9710 ( .A(y[802]), .B(x[802]), .Z(n5721) );
  ANDN U9711 ( .B(x[800]), .A(y[800]), .Z(n5716) );
  OR U9712 ( .A(n5716), .B(x[801]), .Z(n5719) );
  XOR U9713 ( .A(x[801]), .B(n5716), .Z(n5717) );
  NAND U9714 ( .A(n5717), .B(y[801]), .Z(n5718) );
  NAND U9715 ( .A(n5719), .B(n5718), .Z(n5720) );
  AND U9716 ( .A(n5721), .B(n5720), .Z(n21357) );
  NAND U9717 ( .A(n5722), .B(n21357), .Z(n5725) );
  NANDN U9718 ( .A(x[802]), .B(y[802]), .Z(n5724) );
  NANDN U9719 ( .A(x[803]), .B(y[803]), .Z(n5723) );
  AND U9720 ( .A(n5724), .B(n5723), .Z(n21360) );
  NAND U9721 ( .A(n5725), .B(n21360), .Z(n5726) );
  NANDN U9722 ( .A(n12729), .B(n5726), .Z(n5727) );
  NANDN U9723 ( .A(n12725), .B(n5727), .Z(n5729) );
  ANDN U9724 ( .B(x[805]), .A(y[805]), .Z(n12726) );
  NANDN U9725 ( .A(y[804]), .B(x[804]), .Z(n5728) );
  NANDN U9726 ( .A(n12726), .B(n5728), .Z(n12730) );
  ANDN U9727 ( .B(n5729), .A(n12730), .Z(n5730) );
  OR U9728 ( .A(n12728), .B(n5730), .Z(n5733) );
  NANDN U9729 ( .A(y[807]), .B(x[807]), .Z(n5732) );
  NANDN U9730 ( .A(y[806]), .B(x[806]), .Z(n5731) );
  AND U9731 ( .A(n5732), .B(n5731), .Z(n21365) );
  NAND U9732 ( .A(n5733), .B(n21365), .Z(n5736) );
  NANDN U9733 ( .A(x[807]), .B(y[807]), .Z(n5735) );
  NANDN U9734 ( .A(x[808]), .B(y[808]), .Z(n5734) );
  AND U9735 ( .A(n5735), .B(n5734), .Z(n21367) );
  NAND U9736 ( .A(n5736), .B(n21367), .Z(n5737) );
  NANDN U9737 ( .A(n21370), .B(n5737), .Z(n5742) );
  NANDN U9738 ( .A(x[810]), .B(y[810]), .Z(n5739) );
  NANDN U9739 ( .A(x[809]), .B(y[809]), .Z(n5738) );
  AND U9740 ( .A(n5739), .B(n5738), .Z(n5741) );
  NANDN U9741 ( .A(x[811]), .B(y[811]), .Z(n5740) );
  AND U9742 ( .A(n5741), .B(n5740), .Z(n21371) );
  NAND U9743 ( .A(n5742), .B(n21371), .Z(n5749) );
  NANDN U9744 ( .A(y[812]), .B(x[812]), .Z(n5748) );
  ANDN U9745 ( .B(x[810]), .A(y[810]), .Z(n5743) );
  OR U9746 ( .A(n5743), .B(x[811]), .Z(n5746) );
  XOR U9747 ( .A(x[811]), .B(n5743), .Z(n5744) );
  NAND U9748 ( .A(n5744), .B(y[811]), .Z(n5745) );
  NAND U9749 ( .A(n5746), .B(n5745), .Z(n5747) );
  NAND U9750 ( .A(n5748), .B(n5747), .Z(n21374) );
  ANDN U9751 ( .B(n5749), .A(n21374), .Z(n5754) );
  NANDN U9752 ( .A(x[813]), .B(y[813]), .Z(n5751) );
  NANDN U9753 ( .A(x[812]), .B(y[812]), .Z(n5750) );
  AND U9754 ( .A(n5751), .B(n5750), .Z(n5753) );
  NANDN U9755 ( .A(x[814]), .B(y[814]), .Z(n5752) );
  AND U9756 ( .A(n5753), .B(n5752), .Z(n21375) );
  NANDN U9757 ( .A(n5754), .B(n21375), .Z(n5755) );
  NANDN U9758 ( .A(n21377), .B(n5755), .Z(n5758) );
  NANDN U9759 ( .A(x[815]), .B(y[815]), .Z(n5757) );
  NANDN U9760 ( .A(x[816]), .B(y[816]), .Z(n5756) );
  AND U9761 ( .A(n5757), .B(n5756), .Z(n21379) );
  NAND U9762 ( .A(n5758), .B(n21379), .Z(n5759) );
  NANDN U9763 ( .A(n21382), .B(n5759), .Z(n5762) );
  NANDN U9764 ( .A(x[817]), .B(y[817]), .Z(n5761) );
  NANDN U9765 ( .A(x[818]), .B(y[818]), .Z(n5760) );
  AND U9766 ( .A(n5761), .B(n5760), .Z(n21383) );
  NAND U9767 ( .A(n5762), .B(n21383), .Z(n5765) );
  NANDN U9768 ( .A(y[819]), .B(x[819]), .Z(n5764) );
  NANDN U9769 ( .A(y[818]), .B(x[818]), .Z(n5763) );
  NAND U9770 ( .A(n5764), .B(n5763), .Z(n21386) );
  ANDN U9771 ( .B(n5765), .A(n21386), .Z(n5768) );
  NANDN U9772 ( .A(x[819]), .B(y[819]), .Z(n5767) );
  NANDN U9773 ( .A(x[820]), .B(y[820]), .Z(n5766) );
  AND U9774 ( .A(n5767), .B(n5766), .Z(n21387) );
  NANDN U9775 ( .A(n5768), .B(n21387), .Z(n5769) );
  NANDN U9776 ( .A(n21389), .B(n5769), .Z(n5772) );
  NANDN U9777 ( .A(x[821]), .B(y[821]), .Z(n5771) );
  NANDN U9778 ( .A(x[822]), .B(y[822]), .Z(n5770) );
  AND U9779 ( .A(n5771), .B(n5770), .Z(n21391) );
  NAND U9780 ( .A(n5772), .B(n21391), .Z(n5773) );
  NANDN U9781 ( .A(n21394), .B(n5773), .Z(n5774) );
  ANDN U9782 ( .B(y[824]), .A(x[824]), .Z(n12721) );
  ANDN U9783 ( .B(n5774), .A(n12721), .Z(n5775) );
  NANDN U9784 ( .A(x[823]), .B(y[823]), .Z(n21395) );
  NAND U9785 ( .A(n5775), .B(n21395), .Z(n5777) );
  NANDN U9786 ( .A(y[824]), .B(x[824]), .Z(n5776) );
  ANDN U9787 ( .B(x[825]), .A(y[825]), .Z(n12722) );
  ANDN U9788 ( .B(n5776), .A(n12722), .Z(n21397) );
  NAND U9789 ( .A(n5777), .B(n21397), .Z(n5778) );
  NANDN U9790 ( .A(n12724), .B(n5778), .Z(n5783) );
  XNOR U9791 ( .A(x[827]), .B(y[827]), .Z(n5780) );
  NANDN U9792 ( .A(y[826]), .B(x[826]), .Z(n5779) );
  NAND U9793 ( .A(n5780), .B(n5779), .Z(n5781) );
  AND U9794 ( .A(n5782), .B(n5781), .Z(n21401) );
  ANDN U9795 ( .B(n5783), .A(n21401), .Z(n5784) );
  NANDN U9796 ( .A(x[828]), .B(y[828]), .Z(n21403) );
  NANDN U9797 ( .A(n5784), .B(n21403), .Z(n5785) );
  NANDN U9798 ( .A(n21406), .B(n5785), .Z(n5788) );
  NANDN U9799 ( .A(x[829]), .B(y[829]), .Z(n5787) );
  NANDN U9800 ( .A(x[830]), .B(y[830]), .Z(n5786) );
  AND U9801 ( .A(n5787), .B(n5786), .Z(n21407) );
  NAND U9802 ( .A(n5788), .B(n21407), .Z(n5789) );
  NANDN U9803 ( .A(n21410), .B(n5789), .Z(n5792) );
  NANDN U9804 ( .A(x[831]), .B(y[831]), .Z(n5791) );
  NANDN U9805 ( .A(x[832]), .B(y[832]), .Z(n5790) );
  AND U9806 ( .A(n5791), .B(n5790), .Z(n21411) );
  NAND U9807 ( .A(n5792), .B(n21411), .Z(n5795) );
  NANDN U9808 ( .A(y[833]), .B(x[833]), .Z(n5794) );
  NANDN U9809 ( .A(y[832]), .B(x[832]), .Z(n5793) );
  NAND U9810 ( .A(n5794), .B(n5793), .Z(n21413) );
  ANDN U9811 ( .B(n5795), .A(n21413), .Z(n5798) );
  NANDN U9812 ( .A(x[833]), .B(y[833]), .Z(n5797) );
  NANDN U9813 ( .A(x[834]), .B(y[834]), .Z(n5796) );
  AND U9814 ( .A(n5797), .B(n5796), .Z(n21415) );
  NANDN U9815 ( .A(n5798), .B(n21415), .Z(n5799) );
  NANDN U9816 ( .A(n21418), .B(n5799), .Z(n5802) );
  NANDN U9817 ( .A(x[835]), .B(y[835]), .Z(n5801) );
  NANDN U9818 ( .A(x[836]), .B(y[836]), .Z(n5800) );
  AND U9819 ( .A(n5801), .B(n5800), .Z(n21419) );
  NAND U9820 ( .A(n5802), .B(n21419), .Z(n5803) );
  NANDN U9821 ( .A(n21422), .B(n5803), .Z(n5806) );
  NANDN U9822 ( .A(x[837]), .B(y[837]), .Z(n5805) );
  NANDN U9823 ( .A(x[838]), .B(y[838]), .Z(n5804) );
  AND U9824 ( .A(n5805), .B(n5804), .Z(n21423) );
  NAND U9825 ( .A(n5806), .B(n21423), .Z(n5809) );
  NANDN U9826 ( .A(y[838]), .B(x[838]), .Z(n5808) );
  NANDN U9827 ( .A(y[839]), .B(x[839]), .Z(n5807) );
  NAND U9828 ( .A(n5808), .B(n5807), .Z(n21425) );
  ANDN U9829 ( .B(n5809), .A(n21425), .Z(n5810) );
  NANDN U9830 ( .A(x[839]), .B(y[839]), .Z(n21427) );
  NANDN U9831 ( .A(n5810), .B(n21427), .Z(n5811) );
  NANDN U9832 ( .A(n21430), .B(n5811), .Z(n5812) );
  NANDN U9833 ( .A(n21432), .B(n5812), .Z(n5813) );
  NANDN U9834 ( .A(n21434), .B(n5813), .Z(n5816) );
  NANDN U9835 ( .A(x[843]), .B(y[843]), .Z(n5815) );
  NANDN U9836 ( .A(x[844]), .B(y[844]), .Z(n5814) );
  AND U9837 ( .A(n5815), .B(n5814), .Z(n21435) );
  NAND U9838 ( .A(n5816), .B(n21435), .Z(n5819) );
  NANDN U9839 ( .A(y[845]), .B(x[845]), .Z(n5818) );
  NANDN U9840 ( .A(y[844]), .B(x[844]), .Z(n5817) );
  NAND U9841 ( .A(n5818), .B(n5817), .Z(n21437) );
  ANDN U9842 ( .B(n5819), .A(n21437), .Z(n5822) );
  NANDN U9843 ( .A(x[845]), .B(y[845]), .Z(n5821) );
  NANDN U9844 ( .A(x[846]), .B(y[846]), .Z(n5820) );
  AND U9845 ( .A(n5821), .B(n5820), .Z(n21439) );
  NANDN U9846 ( .A(n5822), .B(n21439), .Z(n5823) );
  NANDN U9847 ( .A(n21442), .B(n5823), .Z(n5827) );
  NANDN U9848 ( .A(x[848]), .B(y[848]), .Z(n5825) );
  NANDN U9849 ( .A(x[847]), .B(y[847]), .Z(n5824) );
  NAND U9850 ( .A(n5825), .B(n5824), .Z(n14056) );
  ANDN U9851 ( .B(n5826), .A(n14056), .Z(n21443) );
  NAND U9852 ( .A(n5827), .B(n21443), .Z(n5828) );
  NANDN U9853 ( .A(n21446), .B(n5828), .Z(n5829) );
  NANDN U9854 ( .A(n21448), .B(n5829), .Z(n5830) );
  AND U9855 ( .A(n21450), .B(n5830), .Z(n5831) );
  NANDN U9856 ( .A(x[852]), .B(y[852]), .Z(n21451) );
  NANDN U9857 ( .A(n5831), .B(n21451), .Z(n5834) );
  NANDN U9858 ( .A(y[852]), .B(x[852]), .Z(n5833) );
  NANDN U9859 ( .A(y[853]), .B(x[853]), .Z(n5832) );
  AND U9860 ( .A(n5833), .B(n5832), .Z(n21453) );
  NAND U9861 ( .A(n5834), .B(n21453), .Z(n5835) );
  AND U9862 ( .A(n21455), .B(n5835), .Z(n5838) );
  NANDN U9863 ( .A(y[854]), .B(x[854]), .Z(n5837) );
  NANDN U9864 ( .A(y[855]), .B(x[855]), .Z(n5836) );
  AND U9865 ( .A(n5837), .B(n5836), .Z(n21457) );
  NANDN U9866 ( .A(n5838), .B(n21457), .Z(n5841) );
  NANDN U9867 ( .A(x[856]), .B(y[856]), .Z(n5840) );
  NANDN U9868 ( .A(x[855]), .B(y[855]), .Z(n5839) );
  AND U9869 ( .A(n5840), .B(n5839), .Z(n21459) );
  NAND U9870 ( .A(n5841), .B(n21459), .Z(n5844) );
  NANDN U9871 ( .A(y[856]), .B(x[856]), .Z(n5843) );
  NANDN U9872 ( .A(y[857]), .B(x[857]), .Z(n5842) );
  AND U9873 ( .A(n5843), .B(n5842), .Z(n21462) );
  NAND U9874 ( .A(n5844), .B(n21462), .Z(n5845) );
  NANDN U9875 ( .A(x[857]), .B(y[857]), .Z(n21464) );
  NAND U9876 ( .A(n5845), .B(n21464), .Z(n5846) );
  NANDN U9877 ( .A(n21467), .B(n5846), .Z(n5849) );
  NANDN U9878 ( .A(x[858]), .B(y[858]), .Z(n21463) );
  OR U9879 ( .A(n5847), .B(n21463), .Z(n5848) );
  NANDN U9880 ( .A(x[859]), .B(y[859]), .Z(n21470) );
  NAND U9881 ( .A(n5848), .B(n21470), .Z(n14078) );
  ANDN U9882 ( .B(n5849), .A(n14078), .Z(n5850) );
  OR U9883 ( .A(n12720), .B(n5850), .Z(n5852) );
  NANDN U9884 ( .A(x[861]), .B(y[861]), .Z(n21476) );
  NANDN U9885 ( .A(x[860]), .B(y[860]), .Z(n21471) );
  AND U9886 ( .A(n21476), .B(n21471), .Z(n5851) );
  NAND U9887 ( .A(n5852), .B(n5851), .Z(n5853) );
  NANDN U9888 ( .A(n12719), .B(n5853), .Z(n5854) );
  OR U9889 ( .A(n21478), .B(n5854), .Z(n5855) );
  NANDN U9890 ( .A(n21480), .B(n5855), .Z(n5856) );
  NANDN U9891 ( .A(n21482), .B(n5856), .Z(n5857) );
  NANDN U9892 ( .A(n21484), .B(n5857), .Z(n5858) );
  NANDN U9893 ( .A(n21486), .B(n5858), .Z(n5861) );
  NANDN U9894 ( .A(x[867]), .B(y[867]), .Z(n5860) );
  NANDN U9895 ( .A(x[868]), .B(y[868]), .Z(n5859) );
  AND U9896 ( .A(n5860), .B(n5859), .Z(n21487) );
  NAND U9897 ( .A(n5861), .B(n21487), .Z(n5862) );
  NANDN U9898 ( .A(n21490), .B(n5862), .Z(n5863) );
  NANDN U9899 ( .A(x[869]), .B(y[869]), .Z(n21491) );
  NAND U9900 ( .A(n5863), .B(n21491), .Z(n5864) );
  AND U9901 ( .A(n21494), .B(n5864), .Z(n5867) );
  NANDN U9902 ( .A(x[870]), .B(y[870]), .Z(n5866) );
  NANDN U9903 ( .A(x[871]), .B(y[871]), .Z(n5865) );
  AND U9904 ( .A(n5866), .B(n5865), .Z(n21495) );
  NANDN U9905 ( .A(n5867), .B(n21495), .Z(n5868) );
  NANDN U9906 ( .A(n21498), .B(n5868), .Z(n5871) );
  NANDN U9907 ( .A(x[872]), .B(y[872]), .Z(n5870) );
  NANDN U9908 ( .A(x[873]), .B(y[873]), .Z(n5869) );
  AND U9909 ( .A(n5870), .B(n5869), .Z(n21499) );
  NAND U9910 ( .A(n5871), .B(n21499), .Z(n5872) );
  NANDN U9911 ( .A(n21502), .B(n5872), .Z(n5875) );
  NANDN U9912 ( .A(x[875]), .B(y[875]), .Z(n5874) );
  NANDN U9913 ( .A(x[874]), .B(y[874]), .Z(n5873) );
  AND U9914 ( .A(n5874), .B(n5873), .Z(n21503) );
  NAND U9915 ( .A(n5875), .B(n21503), .Z(n5876) );
  AND U9916 ( .A(n21506), .B(n5876), .Z(n5877) );
  NANDN U9917 ( .A(x[876]), .B(y[876]), .Z(n21507) );
  NANDN U9918 ( .A(n5877), .B(n21507), .Z(n5878) );
  NANDN U9919 ( .A(n21510), .B(n5878), .Z(n5881) );
  NANDN U9920 ( .A(x[877]), .B(y[877]), .Z(n5880) );
  NANDN U9921 ( .A(x[878]), .B(y[878]), .Z(n5879) );
  AND U9922 ( .A(n5880), .B(n5879), .Z(n21511) );
  NAND U9923 ( .A(n5881), .B(n21511), .Z(n5882) );
  NANDN U9924 ( .A(n21514), .B(n5882), .Z(n5885) );
  NANDN U9925 ( .A(x[879]), .B(y[879]), .Z(n5884) );
  NANDN U9926 ( .A(x[880]), .B(y[880]), .Z(n5883) );
  AND U9927 ( .A(n5884), .B(n5883), .Z(n21515) );
  NAND U9928 ( .A(n5885), .B(n21515), .Z(n5888) );
  NANDN U9929 ( .A(y[881]), .B(x[881]), .Z(n5887) );
  NANDN U9930 ( .A(y[880]), .B(x[880]), .Z(n5886) );
  NAND U9931 ( .A(n5887), .B(n5886), .Z(n21517) );
  ANDN U9932 ( .B(n5888), .A(n21517), .Z(n5889) );
  NANDN U9933 ( .A(x[881]), .B(y[881]), .Z(n21520) );
  NANDN U9934 ( .A(n5889), .B(n21520), .Z(n5890) );
  NANDN U9935 ( .A(y[882]), .B(x[882]), .Z(n21523) );
  NAND U9936 ( .A(n5890), .B(n21523), .Z(n5892) );
  NANDN U9937 ( .A(x[883]), .B(y[883]), .Z(n5891) );
  ANDN U9938 ( .B(y[882]), .A(x[882]), .Z(n21519) );
  ANDN U9939 ( .B(n5891), .A(n21519), .Z(n14107) );
  NAND U9940 ( .A(n5892), .B(n14107), .Z(n5893) );
  NANDN U9941 ( .A(n14110), .B(n5893), .Z(n5896) );
  NANDN U9942 ( .A(x[884]), .B(y[884]), .Z(n5895) );
  NANDN U9943 ( .A(x[885]), .B(y[885]), .Z(n5894) );
  AND U9944 ( .A(n5895), .B(n5894), .Z(n21531) );
  NAND U9945 ( .A(n5896), .B(n21531), .Z(n5899) );
  NANDN U9946 ( .A(y[886]), .B(x[886]), .Z(n5898) );
  NANDN U9947 ( .A(y[885]), .B(x[885]), .Z(n5897) );
  NAND U9948 ( .A(n5898), .B(n5897), .Z(n21534) );
  ANDN U9949 ( .B(n5899), .A(n21534), .Z(n5900) );
  ANDN U9950 ( .B(y[887]), .A(x[887]), .Z(n12718) );
  ANDN U9951 ( .B(y[886]), .A(x[886]), .Z(n14113) );
  NOR U9952 ( .A(n12718), .B(n14113), .Z(n21535) );
  NANDN U9953 ( .A(n5900), .B(n21535), .Z(n5901) );
  NANDN U9954 ( .A(y[887]), .B(x[887]), .Z(n21537) );
  NAND U9955 ( .A(n5901), .B(n21537), .Z(n5902) );
  NANDN U9956 ( .A(x[888]), .B(y[888]), .Z(n21539) );
  NAND U9957 ( .A(n5902), .B(n21539), .Z(n5903) );
  NANDN U9958 ( .A(n21541), .B(n5903), .Z(n5906) );
  NANDN U9959 ( .A(x[889]), .B(y[889]), .Z(n5905) );
  NANDN U9960 ( .A(x[890]), .B(y[890]), .Z(n5904) );
  AND U9961 ( .A(n5905), .B(n5904), .Z(n21543) );
  NAND U9962 ( .A(n5906), .B(n21543), .Z(n5909) );
  NANDN U9963 ( .A(y[891]), .B(x[891]), .Z(n5908) );
  NANDN U9964 ( .A(y[890]), .B(x[890]), .Z(n5907) );
  NAND U9965 ( .A(n5908), .B(n5907), .Z(n21546) );
  ANDN U9966 ( .B(n5909), .A(n21546), .Z(n5912) );
  NANDN U9967 ( .A(x[891]), .B(y[891]), .Z(n5911) );
  NANDN U9968 ( .A(x[892]), .B(y[892]), .Z(n5910) );
  AND U9969 ( .A(n5911), .B(n5910), .Z(n21547) );
  NANDN U9970 ( .A(n5912), .B(n21547), .Z(n5913) );
  NANDN U9971 ( .A(n21550), .B(n5913), .Z(n5914) );
  NANDN U9972 ( .A(x[893]), .B(y[893]), .Z(n21552) );
  NAND U9973 ( .A(n5914), .B(n21552), .Z(n5915) );
  NANDN U9974 ( .A(y[894]), .B(x[894]), .Z(n21555) );
  NAND U9975 ( .A(n5915), .B(n21555), .Z(n5916) );
  NANDN U9976 ( .A(n14126), .B(n5916), .Z(n5919) );
  NANDN U9977 ( .A(y[896]), .B(x[896]), .Z(n5918) );
  NANDN U9978 ( .A(y[895]), .B(x[895]), .Z(n5917) );
  NAND U9979 ( .A(n5918), .B(n5917), .Z(n21559) );
  ANDN U9980 ( .B(n5919), .A(n21559), .Z(n5922) );
  NANDN U9981 ( .A(x[896]), .B(y[896]), .Z(n5921) );
  NANDN U9982 ( .A(x[897]), .B(y[897]), .Z(n5920) );
  AND U9983 ( .A(n5921), .B(n5920), .Z(n21561) );
  NANDN U9984 ( .A(n5922), .B(n21561), .Z(n5923) );
  NANDN U9985 ( .A(n21564), .B(n5923), .Z(n5926) );
  NANDN U9986 ( .A(x[899]), .B(y[899]), .Z(n5925) );
  NANDN U9987 ( .A(x[898]), .B(y[898]), .Z(n5924) );
  AND U9988 ( .A(n5925), .B(n5924), .Z(n21565) );
  NAND U9989 ( .A(n5926), .B(n21565), .Z(n5927) );
  NANDN U9990 ( .A(y[899]), .B(x[899]), .Z(n21567) );
  NAND U9991 ( .A(n5927), .B(n21567), .Z(n5928) );
  NANDN U9992 ( .A(x[900]), .B(y[900]), .Z(n21569) );
  NAND U9993 ( .A(n5928), .B(n21569), .Z(n5931) );
  NANDN U9994 ( .A(y[900]), .B(x[900]), .Z(n5930) );
  NANDN U9995 ( .A(y[901]), .B(x[901]), .Z(n5929) );
  AND U9996 ( .A(n5930), .B(n5929), .Z(n21572) );
  NAND U9997 ( .A(n5931), .B(n21572), .Z(n5934) );
  NANDN U9998 ( .A(x[902]), .B(y[902]), .Z(n5933) );
  NANDN U9999 ( .A(x[901]), .B(y[901]), .Z(n5932) );
  AND U10000 ( .A(n5933), .B(n5932), .Z(n21573) );
  NAND U10001 ( .A(n5934), .B(n21573), .Z(n5937) );
  NANDN U10002 ( .A(y[902]), .B(x[902]), .Z(n5936) );
  NANDN U10003 ( .A(y[903]), .B(x[903]), .Z(n5935) );
  AND U10004 ( .A(n5936), .B(n5935), .Z(n21575) );
  NAND U10005 ( .A(n5937), .B(n21575), .Z(n5938) );
  AND U10006 ( .A(n21577), .B(n5938), .Z(n5941) );
  NANDN U10007 ( .A(y[904]), .B(x[904]), .Z(n5940) );
  NANDN U10008 ( .A(y[905]), .B(x[905]), .Z(n5939) );
  AND U10009 ( .A(n5940), .B(n5939), .Z(n21579) );
  NANDN U10010 ( .A(n5941), .B(n21579), .Z(n5942) );
  NANDN U10011 ( .A(x[905]), .B(y[905]), .Z(n21582) );
  NAND U10012 ( .A(n5942), .B(n21582), .Z(n5943) );
  NANDN U10013 ( .A(y[906]), .B(x[906]), .Z(n21585) );
  NAND U10014 ( .A(n5943), .B(n21585), .Z(n5944) );
  NANDN U10015 ( .A(n14141), .B(n5944), .Z(n5945) );
  NANDN U10016 ( .A(n14143), .B(n5945), .Z(n5947) );
  NANDN U10017 ( .A(x[909]), .B(y[909]), .Z(n21593) );
  IV U10018 ( .A(x[908]), .Z(n21595) );
  NAND U10019 ( .A(n21595), .B(y[908]), .Z(n5946) );
  NAND U10020 ( .A(n21593), .B(n5946), .Z(n14144) );
  ANDN U10021 ( .B(n5947), .A(n14144), .Z(n5950) );
  NANDN U10022 ( .A(y[909]), .B(x[909]), .Z(n5949) );
  NANDN U10023 ( .A(y[910]), .B(x[910]), .Z(n5948) );
  AND U10024 ( .A(n5949), .B(n5948), .Z(n21599) );
  NANDN U10025 ( .A(n5950), .B(n21599), .Z(n5953) );
  NANDN U10026 ( .A(x[910]), .B(y[910]), .Z(n5952) );
  NANDN U10027 ( .A(x[911]), .B(y[911]), .Z(n5951) );
  AND U10028 ( .A(n5952), .B(n5951), .Z(n21601) );
  NAND U10029 ( .A(n5953), .B(n21601), .Z(n5954) );
  NANDN U10030 ( .A(y[911]), .B(x[911]), .Z(n21604) );
  NAND U10031 ( .A(n5954), .B(n21604), .Z(n5955) );
  NANDN U10032 ( .A(x[912]), .B(y[912]), .Z(n21605) );
  NAND U10033 ( .A(n5955), .B(n21605), .Z(n5958) );
  NANDN U10034 ( .A(y[912]), .B(x[912]), .Z(n5957) );
  NANDN U10035 ( .A(y[913]), .B(x[913]), .Z(n5956) );
  AND U10036 ( .A(n5957), .B(n5956), .Z(n21607) );
  NAND U10037 ( .A(n5958), .B(n21607), .Z(n5959) );
  AND U10038 ( .A(n21609), .B(n5959), .Z(n5962) );
  NANDN U10039 ( .A(y[914]), .B(x[914]), .Z(n5961) );
  NANDN U10040 ( .A(y[915]), .B(x[915]), .Z(n5960) );
  AND U10041 ( .A(n5961), .B(n5960), .Z(n21611) );
  NANDN U10042 ( .A(n5962), .B(n21611), .Z(n5965) );
  NANDN U10043 ( .A(x[916]), .B(y[916]), .Z(n5964) );
  NANDN U10044 ( .A(x[915]), .B(y[915]), .Z(n5963) );
  AND U10045 ( .A(n5964), .B(n5963), .Z(n21613) );
  NAND U10046 ( .A(n5965), .B(n21613), .Z(n5968) );
  NANDN U10047 ( .A(y[917]), .B(x[917]), .Z(n5967) );
  NANDN U10048 ( .A(y[916]), .B(x[916]), .Z(n5966) );
  AND U10049 ( .A(n5967), .B(n5966), .Z(n21616) );
  NAND U10050 ( .A(n5968), .B(n21616), .Z(n5969) );
  NANDN U10051 ( .A(x[917]), .B(y[917]), .Z(n21617) );
  NAND U10052 ( .A(n5969), .B(n21617), .Z(n5970) );
  NANDN U10053 ( .A(y[918]), .B(x[918]), .Z(n21619) );
  NAND U10054 ( .A(n5970), .B(n21619), .Z(n5971) );
  AND U10055 ( .A(n21621), .B(n5971), .Z(n5972) );
  NANDN U10056 ( .A(y[919]), .B(x[919]), .Z(n14158) );
  ANDN U10057 ( .B(x[920]), .A(y[920]), .Z(n14164) );
  NANDN U10058 ( .A(n5972), .B(n21623), .Z(n5973) );
  NANDN U10059 ( .A(n21626), .B(n5973), .Z(n5974) );
  NANDN U10060 ( .A(n21627), .B(n5974), .Z(n5975) );
  ANDN U10061 ( .B(y[923]), .A(x[923]), .Z(n12717) );
  NAND U10062 ( .A(n5975), .B(n21629), .Z(n5976) );
  NANDN U10063 ( .A(y[923]), .B(x[923]), .Z(n21631) );
  NAND U10064 ( .A(n5976), .B(n21631), .Z(n5977) );
  AND U10065 ( .A(n21633), .B(n5977), .Z(n5980) );
  NANDN U10066 ( .A(y[924]), .B(x[924]), .Z(n5979) );
  NANDN U10067 ( .A(y[925]), .B(x[925]), .Z(n5978) );
  AND U10068 ( .A(n5979), .B(n5978), .Z(n21635) );
  NANDN U10069 ( .A(n5980), .B(n21635), .Z(n5983) );
  NANDN U10070 ( .A(x[926]), .B(y[926]), .Z(n5982) );
  NANDN U10071 ( .A(x[925]), .B(y[925]), .Z(n5981) );
  AND U10072 ( .A(n5982), .B(n5981), .Z(n21637) );
  NAND U10073 ( .A(n5983), .B(n21637), .Z(n5986) );
  NANDN U10074 ( .A(y[926]), .B(x[926]), .Z(n5985) );
  NANDN U10075 ( .A(y[927]), .B(x[927]), .Z(n5984) );
  AND U10076 ( .A(n5985), .B(n5984), .Z(n21640) );
  NAND U10077 ( .A(n5986), .B(n21640), .Z(n5989) );
  NANDN U10078 ( .A(x[928]), .B(y[928]), .Z(n5988) );
  NANDN U10079 ( .A(x[927]), .B(y[927]), .Z(n5987) );
  AND U10080 ( .A(n5988), .B(n5987), .Z(n21641) );
  NAND U10081 ( .A(n5989), .B(n21641), .Z(n5992) );
  NANDN U10082 ( .A(y[928]), .B(x[928]), .Z(n5991) );
  NANDN U10083 ( .A(y[929]), .B(x[929]), .Z(n5990) );
  AND U10084 ( .A(n5991), .B(n5990), .Z(n21643) );
  NAND U10085 ( .A(n5992), .B(n21643), .Z(n5993) );
  AND U10086 ( .A(n21647), .B(n5993), .Z(n5994) );
  NANDN U10087 ( .A(y[930]), .B(x[930]), .Z(n21649) );
  NANDN U10088 ( .A(n5994), .B(n21649), .Z(n5995) );
  NANDN U10089 ( .A(n14182), .B(n5995), .Z(n5996) );
  NANDN U10090 ( .A(n14184), .B(n5996), .Z(n5997) );
  NANDN U10091 ( .A(n14185), .B(n5997), .Z(n6000) );
  NANDN U10092 ( .A(y[933]), .B(x[933]), .Z(n5999) );
  NANDN U10093 ( .A(y[934]), .B(x[934]), .Z(n5998) );
  AND U10094 ( .A(n5999), .B(n5998), .Z(n21662) );
  NAND U10095 ( .A(n6000), .B(n21662), .Z(n6001) );
  AND U10096 ( .A(n21664), .B(n6001), .Z(n6002) );
  NANDN U10097 ( .A(y[935]), .B(x[935]), .Z(n21667) );
  NANDN U10098 ( .A(n6002), .B(n21667), .Z(n6003) );
  NANDN U10099 ( .A(x[936]), .B(y[936]), .Z(n21668) );
  NAND U10100 ( .A(n6003), .B(n21668), .Z(n6006) );
  NANDN U10101 ( .A(y[936]), .B(x[936]), .Z(n6005) );
  NANDN U10102 ( .A(y[937]), .B(x[937]), .Z(n6004) );
  AND U10103 ( .A(n6005), .B(n6004), .Z(n21670) );
  NAND U10104 ( .A(n6006), .B(n21670), .Z(n6009) );
  NANDN U10105 ( .A(x[938]), .B(y[938]), .Z(n6008) );
  NANDN U10106 ( .A(x[937]), .B(y[937]), .Z(n6007) );
  AND U10107 ( .A(n6008), .B(n6007), .Z(n21672) );
  NAND U10108 ( .A(n6009), .B(n21672), .Z(n6012) );
  NANDN U10109 ( .A(y[938]), .B(x[938]), .Z(n6011) );
  NANDN U10110 ( .A(y[939]), .B(x[939]), .Z(n6010) );
  AND U10111 ( .A(n6011), .B(n6010), .Z(n21674) );
  NAND U10112 ( .A(n6012), .B(n21674), .Z(n6013) );
  AND U10113 ( .A(n21676), .B(n6013), .Z(n6016) );
  NANDN U10114 ( .A(y[940]), .B(x[940]), .Z(n6015) );
  NANDN U10115 ( .A(y[941]), .B(x[941]), .Z(n6014) );
  AND U10116 ( .A(n6015), .B(n6014), .Z(n21679) );
  NANDN U10117 ( .A(n6016), .B(n21679), .Z(n6017) );
  AND U10118 ( .A(n21681), .B(n6017), .Z(n6018) );
  NANDN U10119 ( .A(y[942]), .B(x[942]), .Z(n20297) );
  NANDN U10120 ( .A(n6018), .B(n20297), .Z(n6019) );
  NANDN U10121 ( .A(n14198), .B(n6019), .Z(n6020) );
  NANDN U10122 ( .A(y[943]), .B(x[943]), .Z(n14200) );
  ANDN U10123 ( .B(x[944]), .A(y[944]), .Z(n20296) );
  ANDN U10124 ( .B(n14200), .A(n20296), .Z(n20298) );
  NAND U10125 ( .A(n6020), .B(n20298), .Z(n6023) );
  NANDN U10126 ( .A(x[945]), .B(y[945]), .Z(n6022) );
  NANDN U10127 ( .A(x[944]), .B(y[944]), .Z(n6021) );
  AND U10128 ( .A(n6022), .B(n6021), .Z(n21688) );
  NAND U10129 ( .A(n6023), .B(n21688), .Z(n6024) );
  NANDN U10130 ( .A(n21691), .B(n6024), .Z(n6025) );
  AND U10131 ( .A(n21692), .B(n6025), .Z(n6026) );
  NANDN U10132 ( .A(y[947]), .B(x[947]), .Z(n21695) );
  NANDN U10133 ( .A(n6026), .B(n21695), .Z(n6027) );
  NANDN U10134 ( .A(x[948]), .B(y[948]), .Z(n21696) );
  NAND U10135 ( .A(n6027), .B(n21696), .Z(n6030) );
  NANDN U10136 ( .A(y[948]), .B(x[948]), .Z(n6029) );
  NANDN U10137 ( .A(y[949]), .B(x[949]), .Z(n6028) );
  AND U10138 ( .A(n6029), .B(n6028), .Z(n21698) );
  NAND U10139 ( .A(n6030), .B(n21698), .Z(n6033) );
  NANDN U10140 ( .A(x[950]), .B(y[950]), .Z(n6032) );
  NANDN U10141 ( .A(x[949]), .B(y[949]), .Z(n6031) );
  AND U10142 ( .A(n6032), .B(n6031), .Z(n21700) );
  NAND U10143 ( .A(n6033), .B(n21700), .Z(n6036) );
  NANDN U10144 ( .A(y[950]), .B(x[950]), .Z(n6035) );
  NANDN U10145 ( .A(y[951]), .B(x[951]), .Z(n6034) );
  AND U10146 ( .A(n6035), .B(n6034), .Z(n21702) );
  NAND U10147 ( .A(n6036), .B(n21702), .Z(n6037) );
  AND U10148 ( .A(n21704), .B(n6037), .Z(n6040) );
  NANDN U10149 ( .A(y[952]), .B(x[952]), .Z(n6039) );
  NANDN U10150 ( .A(y[953]), .B(x[953]), .Z(n6038) );
  AND U10151 ( .A(n6039), .B(n6038), .Z(n21707) );
  NANDN U10152 ( .A(n6040), .B(n21707), .Z(n6041) );
  NANDN U10153 ( .A(n21708), .B(n6041), .Z(n6042) );
  NANDN U10154 ( .A(y[954]), .B(x[954]), .Z(n20293) );
  NAND U10155 ( .A(n6042), .B(n20293), .Z(n6043) );
  NANDN U10156 ( .A(n14223), .B(n6043), .Z(n6044) );
  ANDN U10157 ( .B(x[956]), .A(y[956]), .Z(n12715) );
  ANDN U10158 ( .B(n6044), .A(n12715), .Z(n6045) );
  NANDN U10159 ( .A(y[955]), .B(x[955]), .Z(n20294) );
  NAND U10160 ( .A(n6045), .B(n20294), .Z(n6046) );
  NAND U10161 ( .A(n6047), .B(n6046), .Z(n6048) );
  ANDN U10162 ( .B(x[957]), .A(y[957]), .Z(n12714) );
  ANDN U10163 ( .B(n6048), .A(n12714), .Z(n6049) );
  NANDN U10164 ( .A(n21722), .B(n6049), .Z(n6050) );
  NANDN U10165 ( .A(n21725), .B(n6050), .Z(n6053) );
  NANDN U10166 ( .A(y[961]), .B(x[961]), .Z(n6052) );
  NANDN U10167 ( .A(y[960]), .B(x[960]), .Z(n6051) );
  NAND U10168 ( .A(n6052), .B(n6051), .Z(n21727) );
  ANDN U10169 ( .B(n6053), .A(n21727), .Z(n6056) );
  NANDN U10170 ( .A(x[961]), .B(y[961]), .Z(n6055) );
  NANDN U10171 ( .A(x[962]), .B(y[962]), .Z(n6054) );
  AND U10172 ( .A(n6055), .B(n6054), .Z(n21728) );
  NANDN U10173 ( .A(n6056), .B(n21728), .Z(n6057) );
  NANDN U10174 ( .A(n21731), .B(n6057), .Z(n6060) );
  NANDN U10175 ( .A(x[963]), .B(y[963]), .Z(n6059) );
  NANDN U10176 ( .A(x[964]), .B(y[964]), .Z(n6058) );
  AND U10177 ( .A(n6059), .B(n6058), .Z(n21732) );
  NAND U10178 ( .A(n6060), .B(n21732), .Z(n6061) );
  NANDN U10179 ( .A(n21734), .B(n6061), .Z(n6062) );
  NANDN U10180 ( .A(x[965]), .B(y[965]), .Z(n21736) );
  NAND U10181 ( .A(n6062), .B(n21736), .Z(n6063) );
  AND U10182 ( .A(n21738), .B(n6063), .Z(n6066) );
  NANDN U10183 ( .A(x[966]), .B(y[966]), .Z(n6065) );
  NANDN U10184 ( .A(x[967]), .B(y[967]), .Z(n6064) );
  AND U10185 ( .A(n6065), .B(n6064), .Z(n21740) );
  NANDN U10186 ( .A(n6066), .B(n21740), .Z(n6067) );
  NANDN U10187 ( .A(n21743), .B(n6067), .Z(n6070) );
  NANDN U10188 ( .A(x[968]), .B(y[968]), .Z(n6069) );
  NANDN U10189 ( .A(x[969]), .B(y[969]), .Z(n6068) );
  AND U10190 ( .A(n6069), .B(n6068), .Z(n21744) );
  NAND U10191 ( .A(n6070), .B(n21744), .Z(n6071) );
  NANDN U10192 ( .A(n21746), .B(n6071), .Z(n6074) );
  NANDN U10193 ( .A(x[971]), .B(y[971]), .Z(n6073) );
  NANDN U10194 ( .A(x[970]), .B(y[970]), .Z(n6072) );
  AND U10195 ( .A(n6073), .B(n6072), .Z(n21748) );
  NAND U10196 ( .A(n6074), .B(n21748), .Z(n6075) );
  AND U10197 ( .A(n21750), .B(n6075), .Z(n6076) );
  NANDN U10198 ( .A(x[972]), .B(y[972]), .Z(n21752) );
  NANDN U10199 ( .A(n6076), .B(n21752), .Z(n6077) );
  NANDN U10200 ( .A(n21755), .B(n6077), .Z(n6080) );
  NANDN U10201 ( .A(x[973]), .B(y[973]), .Z(n6079) );
  NANDN U10202 ( .A(x[974]), .B(y[974]), .Z(n6078) );
  AND U10203 ( .A(n6079), .B(n6078), .Z(n21756) );
  NAND U10204 ( .A(n6080), .B(n21756), .Z(n6081) );
  NANDN U10205 ( .A(n21758), .B(n6081), .Z(n6084) );
  NANDN U10206 ( .A(x[975]), .B(y[975]), .Z(n6083) );
  NANDN U10207 ( .A(x[976]), .B(y[976]), .Z(n6082) );
  AND U10208 ( .A(n6083), .B(n6082), .Z(n21760) );
  NAND U10209 ( .A(n6084), .B(n21760), .Z(n6087) );
  NANDN U10210 ( .A(y[976]), .B(x[976]), .Z(n6086) );
  NANDN U10211 ( .A(y[977]), .B(x[977]), .Z(n6085) );
  NAND U10212 ( .A(n6086), .B(n6085), .Z(n21763) );
  ANDN U10213 ( .B(n6087), .A(n21763), .Z(n6088) );
  NANDN U10214 ( .A(x[977]), .B(y[977]), .Z(n21764) );
  NANDN U10215 ( .A(n6088), .B(n21764), .Z(n6089) );
  NANDN U10216 ( .A(y[978]), .B(x[978]), .Z(n21766) );
  NAND U10217 ( .A(n6089), .B(n21766), .Z(n6092) );
  NANDN U10218 ( .A(x[978]), .B(y[978]), .Z(n6091) );
  NANDN U10219 ( .A(x[979]), .B(y[979]), .Z(n6090) );
  AND U10220 ( .A(n6091), .B(n6090), .Z(n21768) );
  NAND U10221 ( .A(n6092), .B(n21768), .Z(n6093) );
  NANDN U10222 ( .A(n21770), .B(n6093), .Z(n6096) );
  NANDN U10223 ( .A(x[980]), .B(y[980]), .Z(n6095) );
  NANDN U10224 ( .A(x[981]), .B(y[981]), .Z(n6094) );
  AND U10225 ( .A(n6095), .B(n6094), .Z(n21772) );
  NAND U10226 ( .A(n6096), .B(n21772), .Z(n6099) );
  NANDN U10227 ( .A(y[982]), .B(x[982]), .Z(n6098) );
  NANDN U10228 ( .A(y[981]), .B(x[981]), .Z(n6097) );
  NAND U10229 ( .A(n6098), .B(n6097), .Z(n21775) );
  ANDN U10230 ( .B(n6099), .A(n21775), .Z(n6102) );
  NANDN U10231 ( .A(x[983]), .B(y[983]), .Z(n6101) );
  NANDN U10232 ( .A(x[982]), .B(y[982]), .Z(n6100) );
  AND U10233 ( .A(n6101), .B(n6100), .Z(n21776) );
  NANDN U10234 ( .A(n6102), .B(n21776), .Z(n6103) );
  NANDN U10235 ( .A(y[983]), .B(x[983]), .Z(n21778) );
  NAND U10236 ( .A(n6103), .B(n21778), .Z(n6104) );
  NANDN U10237 ( .A(x[984]), .B(y[984]), .Z(n21780) );
  NAND U10238 ( .A(n6104), .B(n21780), .Z(n6105) );
  NANDN U10239 ( .A(n21782), .B(n6105), .Z(n6108) );
  NANDN U10240 ( .A(x[985]), .B(y[985]), .Z(n6107) );
  NANDN U10241 ( .A(x[986]), .B(y[986]), .Z(n6106) );
  AND U10242 ( .A(n6107), .B(n6106), .Z(n21784) );
  NAND U10243 ( .A(n6108), .B(n21784), .Z(n6111) );
  NANDN U10244 ( .A(y[987]), .B(x[987]), .Z(n6110) );
  NANDN U10245 ( .A(y[986]), .B(x[986]), .Z(n6109) );
  NAND U10246 ( .A(n6110), .B(n6109), .Z(n21787) );
  ANDN U10247 ( .B(n6111), .A(n21787), .Z(n6114) );
  NANDN U10248 ( .A(x[987]), .B(y[987]), .Z(n6113) );
  NANDN U10249 ( .A(x[988]), .B(y[988]), .Z(n6112) );
  AND U10250 ( .A(n6113), .B(n6112), .Z(n21788) );
  NANDN U10251 ( .A(n6114), .B(n21788), .Z(n6115) );
  NANDN U10252 ( .A(n21791), .B(n6115), .Z(n6116) );
  NANDN U10253 ( .A(x[989]), .B(y[989]), .Z(n21793) );
  NAND U10254 ( .A(n6116), .B(n21793), .Z(n6118) );
  NAND U10255 ( .A(n6118), .B(n21796), .Z(n6119) );
  NANDN U10256 ( .A(n14269), .B(n6119), .Z(n6120) );
  ANDN U10257 ( .B(x[992]), .A(y[992]), .Z(n12710) );
  ANDN U10258 ( .B(n6120), .A(n12710), .Z(n6122) );
  NANDN U10259 ( .A(x[992]), .B(y[992]), .Z(n6121) );
  ANDN U10260 ( .B(y[993]), .A(x[993]), .Z(n12711) );
  ANDN U10261 ( .B(n6121), .A(n12711), .Z(n21799) );
  NANDN U10262 ( .A(n6122), .B(n21799), .Z(n6123) );
  NANDN U10263 ( .A(n12713), .B(n6123), .Z(n6124) );
  AND U10264 ( .A(n21804), .B(n6124), .Z(n6125) );
  NANDN U10265 ( .A(y[995]), .B(x[995]), .Z(n21807) );
  NANDN U10266 ( .A(n6125), .B(n21807), .Z(n6126) );
  NANDN U10267 ( .A(x[996]), .B(y[996]), .Z(n21808) );
  NAND U10268 ( .A(n6126), .B(n21808), .Z(n6129) );
  NANDN U10269 ( .A(y[996]), .B(x[996]), .Z(n6128) );
  NANDN U10270 ( .A(y[997]), .B(x[997]), .Z(n6127) );
  AND U10271 ( .A(n6128), .B(n6127), .Z(n21810) );
  NAND U10272 ( .A(n6129), .B(n21810), .Z(n6132) );
  NANDN U10273 ( .A(x[998]), .B(y[998]), .Z(n6131) );
  NANDN U10274 ( .A(x[997]), .B(y[997]), .Z(n6130) );
  AND U10275 ( .A(n6131), .B(n6130), .Z(n21812) );
  NAND U10276 ( .A(n6132), .B(n21812), .Z(n6135) );
  NANDN U10277 ( .A(y[998]), .B(x[998]), .Z(n6134) );
  NANDN U10278 ( .A(y[999]), .B(x[999]), .Z(n6133) );
  AND U10279 ( .A(n6134), .B(n6133), .Z(n21814) );
  NAND U10280 ( .A(n6135), .B(n21814), .Z(n6136) );
  AND U10281 ( .A(n21816), .B(n6136), .Z(n6139) );
  NANDN U10282 ( .A(y[1000]), .B(x[1000]), .Z(n6138) );
  NANDN U10283 ( .A(y[1001]), .B(x[1001]), .Z(n6137) );
  AND U10284 ( .A(n6138), .B(n6137), .Z(n21819) );
  NANDN U10285 ( .A(n6139), .B(n21819), .Z(n6140) );
  NANDN U10286 ( .A(x[1001]), .B(y[1001]), .Z(n21821) );
  NAND U10287 ( .A(n6140), .B(n21821), .Z(n6141) );
  NANDN U10288 ( .A(n21824), .B(n6141), .Z(n6145) );
  ANDN U10289 ( .B(y[1003]), .A(x[1003]), .Z(n20292) );
  NANDN U10290 ( .A(x[1002]), .B(y[1002]), .Z(n21820) );
  NANDN U10291 ( .A(x[1005]), .B(y[1005]), .Z(n6144) );
  NANDN U10292 ( .A(x[1004]), .B(y[1004]), .Z(n6143) );
  AND U10293 ( .A(n6144), .B(n6143), .Z(n21828) );
  NAND U10294 ( .A(n6145), .B(n14282), .Z(n6148) );
  NANDN U10295 ( .A(y[1005]), .B(x[1005]), .Z(n6147) );
  NANDN U10296 ( .A(y[1006]), .B(x[1006]), .Z(n6146) );
  AND U10297 ( .A(n6147), .B(n6146), .Z(n21830) );
  NAND U10298 ( .A(n6148), .B(n21830), .Z(n6149) );
  AND U10299 ( .A(n21832), .B(n6149), .Z(n6150) );
  NANDN U10300 ( .A(y[1007]), .B(x[1007]), .Z(n21835) );
  NANDN U10301 ( .A(n6150), .B(n21835), .Z(n6151) );
  NANDN U10302 ( .A(x[1008]), .B(y[1008]), .Z(n21836) );
  NAND U10303 ( .A(n6151), .B(n21836), .Z(n6154) );
  NANDN U10304 ( .A(y[1008]), .B(x[1008]), .Z(n6153) );
  NANDN U10305 ( .A(y[1009]), .B(x[1009]), .Z(n6152) );
  AND U10306 ( .A(n6153), .B(n6152), .Z(n21838) );
  NAND U10307 ( .A(n6154), .B(n21838), .Z(n6157) );
  NANDN U10308 ( .A(x[1010]), .B(y[1010]), .Z(n6156) );
  NANDN U10309 ( .A(x[1009]), .B(y[1009]), .Z(n6155) );
  AND U10310 ( .A(n6156), .B(n6155), .Z(n21840) );
  NAND U10311 ( .A(n6157), .B(n21840), .Z(n6160) );
  NANDN U10312 ( .A(y[1010]), .B(x[1010]), .Z(n6159) );
  NANDN U10313 ( .A(y[1011]), .B(x[1011]), .Z(n6158) );
  AND U10314 ( .A(n6159), .B(n6158), .Z(n21842) );
  NAND U10315 ( .A(n6160), .B(n21842), .Z(n6161) );
  AND U10316 ( .A(n21844), .B(n6161), .Z(n6164) );
  NANDN U10317 ( .A(y[1012]), .B(x[1012]), .Z(n6163) );
  NANDN U10318 ( .A(y[1013]), .B(x[1013]), .Z(n6162) );
  AND U10319 ( .A(n6163), .B(n6162), .Z(n21847) );
  NANDN U10320 ( .A(n6164), .B(n21847), .Z(n6165) );
  NANDN U10321 ( .A(x[1013]), .B(y[1013]), .Z(n21849) );
  NAND U10322 ( .A(n6165), .B(n21849), .Z(n6166) );
  NANDN U10323 ( .A(y[1014]), .B(x[1014]), .Z(n20289) );
  NAND U10324 ( .A(n6166), .B(n20289), .Z(n6167) );
  NANDN U10325 ( .A(x[1014]), .B(y[1014]), .Z(n21848) );
  NANDN U10326 ( .A(x[1015]), .B(y[1015]), .Z(n21855) );
  AND U10327 ( .A(n21848), .B(n21855), .Z(n14295) );
  NAND U10328 ( .A(n6167), .B(n14295), .Z(n6168) );
  ANDN U10329 ( .B(x[1016]), .A(y[1016]), .Z(n14299) );
  ANDN U10330 ( .B(n6168), .A(n14299), .Z(n6169) );
  NANDN U10331 ( .A(y[1015]), .B(x[1015]), .Z(n20290) );
  NAND U10332 ( .A(n6169), .B(n20290), .Z(n6171) );
  NANDN U10333 ( .A(x[1016]), .B(y[1016]), .Z(n6170) );
  ANDN U10334 ( .B(y[1017]), .A(x[1017]), .Z(n14300) );
  ANDN U10335 ( .B(n6170), .A(n14300), .Z(n21856) );
  NAND U10336 ( .A(n6171), .B(n21856), .Z(n6172) );
  NANDN U10337 ( .A(n14302), .B(n6172), .Z(n6173) );
  AND U10338 ( .A(n21860), .B(n6173), .Z(n6176) );
  NANDN U10339 ( .A(y[1019]), .B(x[1019]), .Z(n6175) );
  NANDN U10340 ( .A(y[1020]), .B(x[1020]), .Z(n6174) );
  AND U10341 ( .A(n6175), .B(n6174), .Z(n21862) );
  NANDN U10342 ( .A(n6176), .B(n21862), .Z(n6178) );
  NANDN U10343 ( .A(x[1021]), .B(y[1021]), .Z(n6177) );
  ANDN U10344 ( .B(y[1020]), .A(x[1020]), .Z(n14307) );
  ANDN U10345 ( .B(n6177), .A(n14307), .Z(n21864) );
  NAND U10346 ( .A(n6178), .B(n21864), .Z(n6179) );
  NANDN U10347 ( .A(n21867), .B(n6179), .Z(n6180) );
  ANDN U10348 ( .B(y[1023]), .A(x[1023]), .Z(n12707) );
  NAND U10349 ( .A(n6180), .B(n21868), .Z(n6181) );
  NANDN U10350 ( .A(y[1023]), .B(x[1023]), .Z(n21871) );
  NAND U10351 ( .A(n6181), .B(n21871), .Z(n6182) );
  AND U10352 ( .A(n21872), .B(n6182), .Z(n6185) );
  NANDN U10353 ( .A(y[1024]), .B(x[1024]), .Z(n6184) );
  NANDN U10354 ( .A(y[1025]), .B(x[1025]), .Z(n6183) );
  AND U10355 ( .A(n6184), .B(n6183), .Z(n21874) );
  NANDN U10356 ( .A(n6185), .B(n21874), .Z(n6186) );
  ANDN U10357 ( .B(y[1025]), .A(x[1025]), .Z(n14319) );
  ANDN U10358 ( .B(n6186), .A(n14319), .Z(n6187) );
  NAND U10359 ( .A(n6188), .B(n6187), .Z(n6189) );
  NAND U10360 ( .A(n12705), .B(n6189), .Z(n6190) );
  AND U10361 ( .A(n21880), .B(n6190), .Z(n6192) );
  NANDN U10362 ( .A(y[1028]), .B(x[1028]), .Z(n21883) );
  ANDN U10363 ( .B(x[1027]), .A(y[1027]), .Z(n12706) );
  ANDN U10364 ( .B(n21883), .A(n12706), .Z(n6191) );
  NANDN U10365 ( .A(n6192), .B(n6191), .Z(n6193) );
  AND U10366 ( .A(n21884), .B(n6193), .Z(n6195) );
  NANDN U10367 ( .A(y[1029]), .B(x[1029]), .Z(n21886) );
  ANDN U10368 ( .B(x[1030]), .A(y[1030]), .Z(n12703) );
  ANDN U10369 ( .B(n21886), .A(n12703), .Z(n6194) );
  NANDN U10370 ( .A(n6195), .B(n6194), .Z(n6196) );
  NANDN U10371 ( .A(x[1030]), .B(y[1030]), .Z(n21888) );
  NAND U10372 ( .A(n6196), .B(n21888), .Z(n6197) );
  NANDN U10373 ( .A(n6197), .B(x[1031]), .Z(n6200) );
  XNOR U10374 ( .A(n6197), .B(x[1031]), .Z(n6198) );
  NANDN U10375 ( .A(y[1031]), .B(n6198), .Z(n6199) );
  NAND U10376 ( .A(n6200), .B(n6199), .Z(n6201) );
  NAND U10377 ( .A(n6202), .B(n6201), .Z(n6203) );
  NAND U10378 ( .A(n12701), .B(n6203), .Z(n6204) );
  NAND U10379 ( .A(n6205), .B(n6204), .Z(n6206) );
  NAND U10380 ( .A(n12700), .B(n6206), .Z(n6207) );
  ANDN U10381 ( .B(y[1034]), .A(x[1034]), .Z(n14336) );
  ANDN U10382 ( .B(n6207), .A(n14336), .Z(n6210) );
  NANDN U10383 ( .A(y[1034]), .B(x[1034]), .Z(n6209) );
  NANDN U10384 ( .A(y[1035]), .B(x[1035]), .Z(n6208) );
  AND U10385 ( .A(n6209), .B(n6208), .Z(n21898) );
  NANDN U10386 ( .A(n6210), .B(n21898), .Z(n6213) );
  NANDN U10387 ( .A(x[1036]), .B(y[1036]), .Z(n6212) );
  NANDN U10388 ( .A(x[1035]), .B(y[1035]), .Z(n6211) );
  AND U10389 ( .A(n6212), .B(n6211), .Z(n21900) );
  NAND U10390 ( .A(n6213), .B(n21900), .Z(n6216) );
  NANDN U10391 ( .A(y[1036]), .B(x[1036]), .Z(n6215) );
  NANDN U10392 ( .A(y[1037]), .B(x[1037]), .Z(n6214) );
  AND U10393 ( .A(n6215), .B(n6214), .Z(n21902) );
  NAND U10394 ( .A(n6216), .B(n21902), .Z(n6217) );
  ANDN U10395 ( .B(y[1037]), .A(x[1037]), .Z(n14342) );
  ANDN U10396 ( .B(n6217), .A(n14342), .Z(n6218) );
  IV U10397 ( .A(x[1038]), .Z(n14341) );
  ANDN U10398 ( .B(x[1039]), .A(y[1039]), .Z(n12699) );
  ANDN U10399 ( .B(y[1041]), .A(x[1041]), .Z(n12697) );
  ANDN U10400 ( .B(y[1040]), .A(x[1040]), .Z(n14346) );
  NOR U10401 ( .A(n12697), .B(n14346), .Z(n21912) );
  ANDN U10402 ( .B(x[1042]), .A(y[1042]), .Z(n14354) );
  NANDN U10403 ( .A(y[1041]), .B(x[1041]), .Z(n21914) );
  NANDN U10404 ( .A(x[1042]), .B(y[1042]), .Z(n6221) );
  NANDN U10405 ( .A(x[1043]), .B(y[1043]), .Z(n6219) );
  NANDN U10406 ( .A(n6220), .B(n6219), .Z(n14356) );
  ANDN U10407 ( .B(n6221), .A(n14356), .Z(n21916) );
  NANDN U10408 ( .A(x[1045]), .B(y[1045]), .Z(n6223) );
  NANDN U10409 ( .A(x[1046]), .B(y[1046]), .Z(n6222) );
  AND U10410 ( .A(n6223), .B(n6222), .Z(n21920) );
  NANDN U10411 ( .A(y[1047]), .B(x[1047]), .Z(n6225) );
  NANDN U10412 ( .A(y[1046]), .B(x[1046]), .Z(n6224) );
  NAND U10413 ( .A(n6225), .B(n6224), .Z(n21923) );
  NANDN U10414 ( .A(x[1047]), .B(y[1047]), .Z(n6227) );
  NANDN U10415 ( .A(x[1048]), .B(y[1048]), .Z(n6226) );
  AND U10416 ( .A(n6227), .B(n6226), .Z(n21924) );
  NANDN U10417 ( .A(y[1049]), .B(x[1049]), .Z(n6229) );
  NANDN U10418 ( .A(y[1048]), .B(x[1048]), .Z(n6228) );
  NAND U10419 ( .A(n6229), .B(n6228), .Z(n21927) );
  IV U10420 ( .A(x[1050]), .Z(n12694) );
  NANDN U10421 ( .A(n6231), .B(n12694), .Z(n6230) );
  AND U10422 ( .A(n21932), .B(n6230), .Z(n6234) );
  XOR U10423 ( .A(x[1050]), .B(n6231), .Z(n6232) );
  NAND U10424 ( .A(n6232), .B(y[1050]), .Z(n6233) );
  NAND U10425 ( .A(n6234), .B(n6233), .Z(n6235) );
  ANDN U10426 ( .B(x[1051]), .A(y[1051]), .Z(n12693) );
  ANDN U10427 ( .B(n6235), .A(n12693), .Z(n6236) );
  NANDN U10428 ( .A(y[1052]), .B(x[1052]), .Z(n21934) );
  NAND U10429 ( .A(n6236), .B(n21934), .Z(n6237) );
  ANDN U10430 ( .B(y[1053]), .A(x[1053]), .Z(n12690) );
  ANDN U10431 ( .B(y[1052]), .A(x[1052]), .Z(n12691) );
  NOR U10432 ( .A(n12690), .B(n12691), .Z(n21937) );
  NAND U10433 ( .A(n6237), .B(n21937), .Z(n6238) );
  NAND U10434 ( .A(n6239), .B(n6238), .Z(n6243) );
  NANDN U10435 ( .A(x[1055]), .B(y[1055]), .Z(n6241) );
  NAND U10436 ( .A(n6241), .B(n6240), .Z(n12687) );
  NANDN U10437 ( .A(x[1054]), .B(y[1054]), .Z(n6242) );
  NANDN U10438 ( .A(n12687), .B(n6242), .Z(n21941) );
  ANDN U10439 ( .B(n6243), .A(n21941), .Z(n6244) );
  ANDN U10440 ( .B(n6245), .A(n6244), .Z(n6246) );
  AND U10441 ( .A(n12688), .B(n6246), .Z(n6249) );
  NANDN U10442 ( .A(x[1057]), .B(y[1057]), .Z(n6248) );
  NANDN U10443 ( .A(x[1058]), .B(y[1058]), .Z(n6247) );
  AND U10444 ( .A(n6248), .B(n6247), .Z(n21944) );
  NANDN U10445 ( .A(n6249), .B(n21944), .Z(n6250) );
  AND U10446 ( .A(n21946), .B(n6250), .Z(n6253) );
  NANDN U10447 ( .A(x[1059]), .B(y[1059]), .Z(n6252) );
  NANDN U10448 ( .A(x[1060]), .B(y[1060]), .Z(n6251) );
  AND U10449 ( .A(n6252), .B(n6251), .Z(n21949) );
  NANDN U10450 ( .A(n6253), .B(n21949), .Z(n6254) );
  NANDN U10451 ( .A(n21951), .B(n6254), .Z(n6255) );
  NANDN U10452 ( .A(n12683), .B(n6255), .Z(n6256) );
  NAND U10453 ( .A(n6257), .B(n6256), .Z(n6258) );
  NAND U10454 ( .A(n12682), .B(n6258), .Z(n6259) );
  NANDN U10455 ( .A(x[1063]), .B(y[1063]), .Z(n21956) );
  NANDN U10456 ( .A(n6259), .B(n21956), .Z(n6260) );
  AND U10457 ( .A(n6261), .B(n6260), .Z(n6266) );
  NANDN U10458 ( .A(x[1064]), .B(y[1064]), .Z(n14380) );
  NANDN U10459 ( .A(n14380), .B(n6262), .Z(n6265) );
  NANDN U10460 ( .A(x[1066]), .B(y[1066]), .Z(n6264) );
  NANDN U10461 ( .A(x[1065]), .B(y[1065]), .Z(n6263) );
  AND U10462 ( .A(n6264), .B(n6263), .Z(n14383) );
  NAND U10463 ( .A(n6265), .B(n14383), .Z(n21961) );
  OR U10464 ( .A(n6266), .B(n21961), .Z(n6269) );
  NANDN U10465 ( .A(y[1066]), .B(x[1066]), .Z(n6268) );
  NANDN U10466 ( .A(y[1067]), .B(x[1067]), .Z(n6267) );
  AND U10467 ( .A(n6268), .B(n6267), .Z(n21962) );
  NAND U10468 ( .A(n6269), .B(n21962), .Z(n6270) );
  AND U10469 ( .A(n21964), .B(n6270), .Z(n6273) );
  NANDN U10470 ( .A(y[1068]), .B(x[1068]), .Z(n6272) );
  NANDN U10471 ( .A(y[1069]), .B(x[1069]), .Z(n6271) );
  AND U10472 ( .A(n6272), .B(n6271), .Z(n21966) );
  NANDN U10473 ( .A(n6273), .B(n21966), .Z(n6274) );
  AND U10474 ( .A(n21968), .B(n6274), .Z(n6277) );
  NANDN U10475 ( .A(y[1070]), .B(x[1070]), .Z(n6276) );
  NANDN U10476 ( .A(y[1071]), .B(x[1071]), .Z(n6275) );
  AND U10477 ( .A(n6276), .B(n6275), .Z(n21971) );
  NANDN U10478 ( .A(n6277), .B(n21971), .Z(n6278) );
  AND U10479 ( .A(n21972), .B(n6278), .Z(n6281) );
  NANDN U10480 ( .A(y[1072]), .B(x[1072]), .Z(n6280) );
  NANDN U10481 ( .A(y[1073]), .B(x[1073]), .Z(n6279) );
  AND U10482 ( .A(n6280), .B(n6279), .Z(n21974) );
  NANDN U10483 ( .A(n6281), .B(n21974), .Z(n6282) );
  NANDN U10484 ( .A(n12679), .B(n6282), .Z(n6283) );
  NANDN U10485 ( .A(n21979), .B(n6283), .Z(n6287) );
  ANDN U10486 ( .B(y[1074]), .A(x[1074]), .Z(n12678) );
  NANDN U10487 ( .A(x[1075]), .B(y[1075]), .Z(n21980) );
  NANDN U10488 ( .A(n12678), .B(n21980), .Z(n6285) );
  NAND U10489 ( .A(n6285), .B(n6284), .Z(n6286) );
  AND U10490 ( .A(n6287), .B(n6286), .Z(n6288) );
  NANDN U10491 ( .A(y[1076]), .B(x[1076]), .Z(n21982) );
  NANDN U10492 ( .A(n6288), .B(n21982), .Z(n6289) );
  ANDN U10493 ( .B(y[1077]), .A(x[1077]), .Z(n12677) );
  NANDN U10494 ( .A(x[1076]), .B(y[1076]), .Z(n14394) );
  NANDN U10495 ( .A(n12677), .B(n14394), .Z(n21985) );
  ANDN U10496 ( .B(n6289), .A(n21985), .Z(n6291) );
  NANDN U10497 ( .A(y[1077]), .B(x[1077]), .Z(n21986) );
  ANDN U10498 ( .B(x[1078]), .A(y[1078]), .Z(n14401) );
  ANDN U10499 ( .B(n21986), .A(n14401), .Z(n6290) );
  NANDN U10500 ( .A(n6291), .B(n6290), .Z(n6292) );
  AND U10501 ( .A(n21989), .B(n6292), .Z(n6293) );
  NAND U10502 ( .A(n6294), .B(n6293), .Z(n6295) );
  NAND U10503 ( .A(n6296), .B(n6295), .Z(n6297) );
  ANDN U10504 ( .B(y[1080]), .A(x[1080]), .Z(n12676) );
  ANDN U10505 ( .B(n6297), .A(n12676), .Z(n6298) );
  NAND U10506 ( .A(n6299), .B(n6298), .Z(n6300) );
  NAND U10507 ( .A(n12674), .B(n6300), .Z(n6301) );
  ANDN U10508 ( .B(y[1082]), .A(x[1082]), .Z(n12672) );
  ANDN U10509 ( .B(n6301), .A(n12672), .Z(n6304) );
  NANDN U10510 ( .A(y[1082]), .B(x[1082]), .Z(n6303) );
  NANDN U10511 ( .A(y[1083]), .B(x[1083]), .Z(n6302) );
  AND U10512 ( .A(n6303), .B(n6302), .Z(n21998) );
  NANDN U10513 ( .A(n6304), .B(n21998), .Z(n6305) );
  NANDN U10514 ( .A(n22000), .B(n6305), .Z(n6308) );
  NANDN U10515 ( .A(y[1084]), .B(x[1084]), .Z(n6307) );
  NANDN U10516 ( .A(y[1085]), .B(x[1085]), .Z(n6306) );
  AND U10517 ( .A(n6307), .B(n6306), .Z(n22002) );
  NAND U10518 ( .A(n6308), .B(n22002), .Z(n6309) );
  NANDN U10519 ( .A(n12670), .B(n6309), .Z(n6312) );
  NANDN U10520 ( .A(y[1087]), .B(x[1087]), .Z(n6311) );
  NANDN U10521 ( .A(y[1086]), .B(x[1086]), .Z(n6310) );
  NAND U10522 ( .A(n6311), .B(n6310), .Z(n22007) );
  ANDN U10523 ( .B(n6312), .A(n22007), .Z(n6313) );
  ANDN U10524 ( .B(n12667), .A(n6313), .Z(n6316) );
  XNOR U10525 ( .A(y[1087]), .B(x[1087]), .Z(n6314) );
  ANDN U10526 ( .B(y[1086]), .A(x[1086]), .Z(n12669) );
  NAND U10527 ( .A(n6314), .B(n12669), .Z(n6315) );
  NAND U10528 ( .A(n6316), .B(n6315), .Z(n6317) );
  NANDN U10529 ( .A(n14413), .B(n6317), .Z(n6318) );
  NANDN U10530 ( .A(n12668), .B(n6318), .Z(n6319) );
  ANDN U10531 ( .B(x[1090]), .A(y[1090]), .Z(n14420) );
  ANDN U10532 ( .B(n6319), .A(n14420), .Z(n6320) );
  NANDN U10533 ( .A(n14415), .B(n6320), .Z(n6323) );
  NANDN U10534 ( .A(x[1090]), .B(y[1090]), .Z(n6322) );
  NANDN U10535 ( .A(x[1091]), .B(y[1091]), .Z(n6321) );
  NANDN U10536 ( .A(x[1092]), .B(y[1092]), .Z(n6324) );
  NAND U10537 ( .A(n6321), .B(n6324), .Z(n14422) );
  ANDN U10538 ( .B(n6322), .A(n14422), .Z(n22013) );
  NAND U10539 ( .A(n6323), .B(n22013), .Z(n6326) );
  ANDN U10540 ( .B(x[1091]), .A(y[1091]), .Z(n14419) );
  NAND U10541 ( .A(n6324), .B(n14419), .Z(n6325) );
  NAND U10542 ( .A(n6326), .B(n6325), .Z(n6329) );
  NANDN U10543 ( .A(y[1093]), .B(x[1093]), .Z(n6328) );
  NANDN U10544 ( .A(y[1092]), .B(x[1092]), .Z(n6327) );
  NAND U10545 ( .A(n6328), .B(n6327), .Z(n14423) );
  OR U10546 ( .A(n6329), .B(n14423), .Z(n6332) );
  NANDN U10547 ( .A(x[1093]), .B(y[1093]), .Z(n6331) );
  NANDN U10548 ( .A(x[1094]), .B(y[1094]), .Z(n6330) );
  AND U10549 ( .A(n6331), .B(n6330), .Z(n22016) );
  NAND U10550 ( .A(n6332), .B(n22016), .Z(n6333) );
  AND U10551 ( .A(n22018), .B(n6333), .Z(n6336) );
  NANDN U10552 ( .A(x[1095]), .B(y[1095]), .Z(n6335) );
  NANDN U10553 ( .A(x[1096]), .B(y[1096]), .Z(n6334) );
  AND U10554 ( .A(n6335), .B(n6334), .Z(n22020) );
  NANDN U10555 ( .A(n6336), .B(n22020), .Z(n6337) );
  AND U10556 ( .A(n22022), .B(n6337), .Z(n6338) );
  NOR U10557 ( .A(n14432), .B(n6338), .Z(n6340) );
  IV U10558 ( .A(x[1098]), .Z(n14430) );
  NANDN U10559 ( .A(n6340), .B(n14430), .Z(n6339) );
  AND U10560 ( .A(n22028), .B(n6339), .Z(n6343) );
  XOR U10561 ( .A(x[1098]), .B(n6340), .Z(n6341) );
  NAND U10562 ( .A(n6341), .B(y[1098]), .Z(n6342) );
  NAND U10563 ( .A(n6343), .B(n6342), .Z(n6344) );
  ANDN U10564 ( .B(x[1099]), .A(y[1099]), .Z(n12666) );
  ANDN U10565 ( .B(n6344), .A(n12666), .Z(n6345) );
  NANDN U10566 ( .A(y[1100]), .B(x[1100]), .Z(n22030) );
  NAND U10567 ( .A(n6345), .B(n22030), .Z(n6346) );
  ANDN U10568 ( .B(y[1101]), .A(x[1101]), .Z(n14441) );
  ANDN U10569 ( .B(y[1100]), .A(x[1100]), .Z(n12664) );
  NOR U10570 ( .A(n14441), .B(n12664), .Z(n22032) );
  NAND U10571 ( .A(n6346), .B(n22032), .Z(n6347) );
  NAND U10572 ( .A(n6348), .B(n6347), .Z(n6352) );
  NANDN U10573 ( .A(x[1103]), .B(y[1103]), .Z(n6350) );
  NAND U10574 ( .A(n6350), .B(n6349), .Z(n12661) );
  NANDN U10575 ( .A(x[1102]), .B(y[1102]), .Z(n6351) );
  NANDN U10576 ( .A(n12661), .B(n6351), .Z(n22036) );
  ANDN U10577 ( .B(n6352), .A(n22036), .Z(n6353) );
  ANDN U10578 ( .B(n6354), .A(n6353), .Z(n6355) );
  AND U10579 ( .A(n12662), .B(n6355), .Z(n6358) );
  NANDN U10580 ( .A(x[1105]), .B(y[1105]), .Z(n6357) );
  NANDN U10581 ( .A(x[1106]), .B(y[1106]), .Z(n6356) );
  AND U10582 ( .A(n6357), .B(n6356), .Z(n22040) );
  NANDN U10583 ( .A(n6358), .B(n22040), .Z(n6359) );
  AND U10584 ( .A(n22042), .B(n6359), .Z(n6362) );
  NANDN U10585 ( .A(x[1107]), .B(y[1107]), .Z(n6361) );
  NANDN U10586 ( .A(x[1108]), .B(y[1108]), .Z(n6360) );
  AND U10587 ( .A(n6361), .B(n6360), .Z(n22044) );
  NANDN U10588 ( .A(n6362), .B(n22044), .Z(n6365) );
  NANDN U10589 ( .A(y[1109]), .B(x[1109]), .Z(n6364) );
  NANDN U10590 ( .A(y[1108]), .B(x[1108]), .Z(n6363) );
  AND U10591 ( .A(n6364), .B(n6363), .Z(n22046) );
  NAND U10592 ( .A(n6365), .B(n22046), .Z(n6366) );
  NANDN U10593 ( .A(x[1109]), .B(y[1109]), .Z(n22049) );
  NAND U10594 ( .A(n6366), .B(n22049), .Z(n6367) );
  NANDN U10595 ( .A(n12657), .B(n6367), .Z(n6368) );
  NANDN U10596 ( .A(n6369), .B(n6368), .Z(n6370) );
  ANDN U10597 ( .B(x[1111]), .A(y[1111]), .Z(n12656) );
  ANDN U10598 ( .B(n6370), .A(n12656), .Z(n6371) );
  NANDN U10599 ( .A(n22057), .B(n6371), .Z(n6372) );
  NANDN U10600 ( .A(n22059), .B(n6372), .Z(n6375) );
  NANDN U10601 ( .A(y[1115]), .B(x[1115]), .Z(n6374) );
  NANDN U10602 ( .A(y[1114]), .B(x[1114]), .Z(n6373) );
  NAND U10603 ( .A(n6374), .B(n6373), .Z(n22060) );
  ANDN U10604 ( .B(n6375), .A(n22060), .Z(n6378) );
  NANDN U10605 ( .A(x[1115]), .B(y[1115]), .Z(n6377) );
  NANDN U10606 ( .A(x[1116]), .B(y[1116]), .Z(n6376) );
  AND U10607 ( .A(n6377), .B(n6376), .Z(n22062) );
  NANDN U10608 ( .A(n6378), .B(n22062), .Z(n6381) );
  NANDN U10609 ( .A(y[1117]), .B(x[1117]), .Z(n6380) );
  NANDN U10610 ( .A(y[1116]), .B(x[1116]), .Z(n6379) );
  NAND U10611 ( .A(n6380), .B(n6379), .Z(n22065) );
  ANDN U10612 ( .B(n6381), .A(n22065), .Z(n6384) );
  NANDN U10613 ( .A(x[1117]), .B(y[1117]), .Z(n6383) );
  NANDN U10614 ( .A(x[1118]), .B(y[1118]), .Z(n6382) );
  AND U10615 ( .A(n6383), .B(n6382), .Z(n22066) );
  NANDN U10616 ( .A(n6384), .B(n22066), .Z(n6387) );
  NANDN U10617 ( .A(y[1119]), .B(x[1119]), .Z(n6386) );
  NANDN U10618 ( .A(y[1118]), .B(x[1118]), .Z(n6385) );
  NAND U10619 ( .A(n6386), .B(n6385), .Z(n22069) );
  ANDN U10620 ( .B(n6387), .A(n22069), .Z(n6390) );
  NANDN U10621 ( .A(x[1119]), .B(y[1119]), .Z(n6389) );
  NANDN U10622 ( .A(x[1120]), .B(y[1120]), .Z(n6388) );
  AND U10623 ( .A(n6389), .B(n6388), .Z(n22070) );
  NANDN U10624 ( .A(n6390), .B(n22070), .Z(n6391) );
  NANDN U10625 ( .A(n22072), .B(n6391), .Z(n6392) );
  ANDN U10626 ( .B(y[1121]), .A(x[1121]), .Z(n12653) );
  ANDN U10627 ( .B(n6392), .A(n12653), .Z(n6394) );
  IV U10628 ( .A(x[1122]), .Z(n12652) );
  NANDN U10629 ( .A(n6394), .B(n12652), .Z(n6393) );
  AND U10630 ( .A(n22078), .B(n6393), .Z(n6397) );
  XOR U10631 ( .A(x[1122]), .B(n6394), .Z(n6395) );
  NAND U10632 ( .A(n6395), .B(y[1122]), .Z(n6396) );
  NAND U10633 ( .A(n6397), .B(n6396), .Z(n6398) );
  AND U10634 ( .A(n22080), .B(n6398), .Z(n6399) );
  NANDN U10635 ( .A(n12651), .B(n6399), .Z(n6400) );
  ANDN U10636 ( .B(y[1125]), .A(x[1125]), .Z(n12648) );
  ANDN U10637 ( .B(y[1124]), .A(x[1124]), .Z(n12649) );
  NOR U10638 ( .A(n12648), .B(n12649), .Z(n22082) );
  NAND U10639 ( .A(n6400), .B(n22082), .Z(n6401) );
  ANDN U10640 ( .B(x[1125]), .A(y[1125]), .Z(n22084) );
  ANDN U10641 ( .B(n6401), .A(n22084), .Z(n6402) );
  NANDN U10642 ( .A(n12647), .B(n6402), .Z(n6403) );
  NANDN U10643 ( .A(x[1126]), .B(y[1126]), .Z(n22086) );
  NAND U10644 ( .A(n6403), .B(n22086), .Z(n6404) );
  NAND U10645 ( .A(n6405), .B(n6404), .Z(n6406) );
  NAND U10646 ( .A(n14472), .B(n6406), .Z(n6407) );
  NAND U10647 ( .A(n6408), .B(n6407), .Z(n6409) );
  NAND U10648 ( .A(n14471), .B(n6409), .Z(n6410) );
  ANDN U10649 ( .B(x[1129]), .A(y[1129]), .Z(n12645) );
  NANDN U10650 ( .A(x[1129]), .B(y[1129]), .Z(n6412) );
  NANDN U10651 ( .A(x[1130]), .B(y[1130]), .Z(n6411) );
  AND U10652 ( .A(n6412), .B(n6411), .Z(n22094) );
  NANDN U10653 ( .A(y[1131]), .B(x[1131]), .Z(n6414) );
  NANDN U10654 ( .A(y[1130]), .B(x[1130]), .Z(n6413) );
  NAND U10655 ( .A(n6414), .B(n6413), .Z(n22096) );
  NANDN U10656 ( .A(x[1131]), .B(y[1131]), .Z(n6416) );
  NANDN U10657 ( .A(x[1132]), .B(y[1132]), .Z(n6415) );
  AND U10658 ( .A(n6416), .B(n6415), .Z(n22098) );
  NANDN U10659 ( .A(y[1136]), .B(x[1136]), .Z(n22108) );
  ANDN U10660 ( .B(x[1135]), .A(y[1135]), .Z(n14482) );
  NANDN U10661 ( .A(y[1137]), .B(x[1137]), .Z(n22113) );
  ANDN U10662 ( .B(x[1138]), .A(y[1138]), .Z(n12640) );
  NANDN U10663 ( .A(x[1140]), .B(y[1140]), .Z(n6418) );
  NANDN U10664 ( .A(x[1139]), .B(y[1139]), .Z(n6417) );
  AND U10665 ( .A(n6418), .B(n6417), .Z(n22118) );
  NANDN U10666 ( .A(y[1140]), .B(x[1140]), .Z(n6420) );
  NANDN U10667 ( .A(y[1141]), .B(x[1141]), .Z(n6419) );
  AND U10668 ( .A(n6420), .B(n6419), .Z(n22120) );
  NAND U10669 ( .A(n6421), .B(n22120), .Z(n6424) );
  NANDN U10670 ( .A(x[1142]), .B(y[1142]), .Z(n6423) );
  NANDN U10671 ( .A(x[1141]), .B(y[1141]), .Z(n6422) );
  AND U10672 ( .A(n6423), .B(n6422), .Z(n22122) );
  NAND U10673 ( .A(n6424), .B(n22122), .Z(n6427) );
  NANDN U10674 ( .A(y[1142]), .B(x[1142]), .Z(n6426) );
  NANDN U10675 ( .A(y[1143]), .B(x[1143]), .Z(n6425) );
  AND U10676 ( .A(n6426), .B(n6425), .Z(n22125) );
  NAND U10677 ( .A(n6427), .B(n22125), .Z(n6428) );
  AND U10678 ( .A(n22126), .B(n6428), .Z(n6431) );
  NANDN U10679 ( .A(y[1144]), .B(x[1144]), .Z(n6430) );
  NANDN U10680 ( .A(y[1145]), .B(x[1145]), .Z(n6429) );
  AND U10681 ( .A(n6430), .B(n6429), .Z(n22128) );
  NANDN U10682 ( .A(n6431), .B(n22128), .Z(n6436) );
  NANDN U10683 ( .A(x[1146]), .B(y[1146]), .Z(n6433) );
  NANDN U10684 ( .A(x[1145]), .B(y[1145]), .Z(n6432) );
  AND U10685 ( .A(n6433), .B(n6432), .Z(n6435) );
  NANDN U10686 ( .A(x[1147]), .B(y[1147]), .Z(n6434) );
  AND U10687 ( .A(n6435), .B(n6434), .Z(n22130) );
  NAND U10688 ( .A(n6436), .B(n22130), .Z(n6437) );
  NANDN U10689 ( .A(n12639), .B(n6437), .Z(n6438) );
  NANDN U10690 ( .A(n14500), .B(n6438), .Z(n6439) );
  ANDN U10691 ( .B(x[1149]), .A(y[1149]), .Z(n14501) );
  ANDN U10692 ( .B(n6439), .A(n14501), .Z(n6440) );
  NAND U10693 ( .A(n6441), .B(n6440), .Z(n6442) );
  NAND U10694 ( .A(n6443), .B(n6442), .Z(n6444) );
  ANDN U10695 ( .B(x[1151]), .A(y[1151]), .Z(n14506) );
  ANDN U10696 ( .B(n6444), .A(n14506), .Z(n6445) );
  NAND U10697 ( .A(n6446), .B(n6445), .Z(n6447) );
  NAND U10698 ( .A(n12637), .B(n6447), .Z(n6448) );
  ANDN U10699 ( .B(x[1153]), .A(y[1153]), .Z(n14510) );
  ANDN U10700 ( .B(n6448), .A(n14510), .Z(n6451) );
  NANDN U10701 ( .A(x[1153]), .B(y[1153]), .Z(n6450) );
  NANDN U10702 ( .A(x[1154]), .B(y[1154]), .Z(n6449) );
  AND U10703 ( .A(n6450), .B(n6449), .Z(n22142) );
  NANDN U10704 ( .A(n6451), .B(n22142), .Z(n6454) );
  NANDN U10705 ( .A(y[1155]), .B(x[1155]), .Z(n6453) );
  NANDN U10706 ( .A(y[1154]), .B(x[1154]), .Z(n6452) );
  NAND U10707 ( .A(n6453), .B(n6452), .Z(n22145) );
  ANDN U10708 ( .B(n6454), .A(n22145), .Z(n6457) );
  NANDN U10709 ( .A(x[1155]), .B(y[1155]), .Z(n6456) );
  NANDN U10710 ( .A(x[1156]), .B(y[1156]), .Z(n6455) );
  AND U10711 ( .A(n6456), .B(n6455), .Z(n22146) );
  NANDN U10712 ( .A(n6457), .B(n22146), .Z(n6458) );
  NANDN U10713 ( .A(n22148), .B(n6458), .Z(n6461) );
  NANDN U10714 ( .A(x[1158]), .B(y[1158]), .Z(n6460) );
  NANDN U10715 ( .A(x[1157]), .B(y[1157]), .Z(n6459) );
  NAND U10716 ( .A(n6460), .B(n6459), .Z(n14516) );
  NOR U10717 ( .A(n12635), .B(n14516), .Z(n22150) );
  NAND U10718 ( .A(n6461), .B(n22150), .Z(n6462) );
  NANDN U10719 ( .A(n22153), .B(n6462), .Z(n6463) );
  NANDN U10720 ( .A(n22155), .B(n6463), .Z(n6466) );
  NANDN U10721 ( .A(y[1163]), .B(x[1163]), .Z(n6465) );
  NANDN U10722 ( .A(y[1162]), .B(x[1162]), .Z(n6464) );
  NAND U10723 ( .A(n6465), .B(n6464), .Z(n22157) );
  ANDN U10724 ( .B(n6466), .A(n22157), .Z(n6469) );
  NANDN U10725 ( .A(x[1163]), .B(y[1163]), .Z(n6468) );
  NANDN U10726 ( .A(x[1164]), .B(y[1164]), .Z(n6467) );
  AND U10727 ( .A(n6468), .B(n6467), .Z(n22158) );
  NANDN U10728 ( .A(n6469), .B(n22158), .Z(n6472) );
  NANDN U10729 ( .A(y[1165]), .B(x[1165]), .Z(n6471) );
  NANDN U10730 ( .A(y[1164]), .B(x[1164]), .Z(n6470) );
  NAND U10731 ( .A(n6471), .B(n6470), .Z(n22160) );
  ANDN U10732 ( .B(n6472), .A(n22160), .Z(n6475) );
  NANDN U10733 ( .A(x[1165]), .B(y[1165]), .Z(n6474) );
  NANDN U10734 ( .A(x[1166]), .B(y[1166]), .Z(n6473) );
  AND U10735 ( .A(n6474), .B(n6473), .Z(n22162) );
  NANDN U10736 ( .A(n6475), .B(n22162), .Z(n6476) );
  NANDN U10737 ( .A(n22165), .B(n6476), .Z(n6479) );
  NANDN U10738 ( .A(x[1167]), .B(y[1167]), .Z(n6478) );
  NANDN U10739 ( .A(x[1168]), .B(y[1168]), .Z(n6477) );
  AND U10740 ( .A(n6478), .B(n6477), .Z(n22166) );
  NAND U10741 ( .A(n6479), .B(n22166), .Z(n6480) );
  NANDN U10742 ( .A(n22169), .B(n6480), .Z(n6483) );
  ANDN U10743 ( .B(y[1171]), .A(x[1171]), .Z(n6486) );
  NANDN U10744 ( .A(x[1170]), .B(y[1170]), .Z(n6482) );
  NANDN U10745 ( .A(x[1169]), .B(y[1169]), .Z(n6481) );
  NAND U10746 ( .A(n6482), .B(n6481), .Z(n14536) );
  NOR U10747 ( .A(n6486), .B(n14536), .Z(n22170) );
  NAND U10748 ( .A(n6483), .B(n22170), .Z(n6490) );
  NANDN U10749 ( .A(y[1172]), .B(x[1172]), .Z(n6484) );
  NANDN U10750 ( .A(n6485), .B(n6484), .Z(n14542) );
  IV U10751 ( .A(n6486), .Z(n12633) );
  NANDN U10752 ( .A(y[1170]), .B(x[1170]), .Z(n6488) );
  NANDN U10753 ( .A(y[1171]), .B(x[1171]), .Z(n6487) );
  NAND U10754 ( .A(n6488), .B(n6487), .Z(n14538) );
  NAND U10755 ( .A(n12633), .B(n14538), .Z(n6489) );
  NANDN U10756 ( .A(n14542), .B(n6489), .Z(n22172) );
  ANDN U10757 ( .B(n6490), .A(n22172), .Z(n6491) );
  OR U10758 ( .A(n22174), .B(n6491), .Z(n6492) );
  NANDN U10759 ( .A(n12631), .B(n6492), .Z(n6493) );
  NANDN U10760 ( .A(x[1174]), .B(y[1174]), .Z(n22175) );
  NAND U10761 ( .A(n6493), .B(n22175), .Z(n6494) );
  NAND U10762 ( .A(n6495), .B(n6494), .Z(n6496) );
  NAND U10763 ( .A(n14547), .B(n6496), .Z(n6497) );
  NAND U10764 ( .A(n6498), .B(n6497), .Z(n6499) );
  NAND U10765 ( .A(n14546), .B(n6499), .Z(n6500) );
  ANDN U10766 ( .B(x[1177]), .A(y[1177]), .Z(n12629) );
  ANDN U10767 ( .B(n6500), .A(n12629), .Z(n6503) );
  NANDN U10768 ( .A(x[1177]), .B(y[1177]), .Z(n6502) );
  NANDN U10769 ( .A(x[1178]), .B(y[1178]), .Z(n6501) );
  AND U10770 ( .A(n6502), .B(n6501), .Z(n22184) );
  NANDN U10771 ( .A(n6503), .B(n22184), .Z(n6506) );
  NANDN U10772 ( .A(y[1179]), .B(x[1179]), .Z(n6505) );
  NANDN U10773 ( .A(y[1178]), .B(x[1178]), .Z(n6504) );
  NAND U10774 ( .A(n6505), .B(n6504), .Z(n22187) );
  ANDN U10775 ( .B(n6506), .A(n22187), .Z(n6509) );
  NANDN U10776 ( .A(x[1179]), .B(y[1179]), .Z(n6508) );
  NANDN U10777 ( .A(x[1180]), .B(y[1180]), .Z(n6507) );
  AND U10778 ( .A(n6508), .B(n6507), .Z(n22188) );
  NANDN U10779 ( .A(n6509), .B(n22188), .Z(n6512) );
  NANDN U10780 ( .A(y[1181]), .B(x[1181]), .Z(n6511) );
  NANDN U10781 ( .A(y[1180]), .B(x[1180]), .Z(n6510) );
  NAND U10782 ( .A(n6511), .B(n6510), .Z(n22190) );
  ANDN U10783 ( .B(n6512), .A(n22190), .Z(n6515) );
  NANDN U10784 ( .A(x[1181]), .B(y[1181]), .Z(n6514) );
  NANDN U10785 ( .A(x[1182]), .B(y[1182]), .Z(n6513) );
  AND U10786 ( .A(n6514), .B(n6513), .Z(n22192) );
  NANDN U10787 ( .A(n6515), .B(n22192), .Z(n6516) );
  NANDN U10788 ( .A(n22195), .B(n6516), .Z(n6517) );
  NANDN U10789 ( .A(x[1183]), .B(y[1183]), .Z(n22196) );
  NAND U10790 ( .A(n6517), .B(n22196), .Z(n6518) );
  NANDN U10791 ( .A(y[1184]), .B(x[1184]), .Z(n22198) );
  NAND U10792 ( .A(n6518), .B(n22198), .Z(n6519) );
  ANDN U10793 ( .B(y[1185]), .A(x[1185]), .Z(n12627) );
  ANDN U10794 ( .B(y[1184]), .A(x[1184]), .Z(n14556) );
  NOR U10795 ( .A(n12627), .B(n14556), .Z(n22200) );
  NAND U10796 ( .A(n6519), .B(n22200), .Z(n6520) );
  ANDN U10797 ( .B(x[1186]), .A(y[1186]), .Z(n12625) );
  ANDN U10798 ( .B(n6520), .A(n12625), .Z(n6521) );
  NANDN U10799 ( .A(y[1185]), .B(x[1185]), .Z(n22203) );
  NAND U10800 ( .A(n6521), .B(n22203), .Z(n6522) );
  ANDN U10801 ( .B(y[1187]), .A(x[1187]), .Z(n14564) );
  ANDN U10802 ( .B(n6522), .A(n14564), .Z(n6523) );
  NANDN U10803 ( .A(x[1186]), .B(y[1186]), .Z(n22204) );
  NAND U10804 ( .A(n6523), .B(n22204), .Z(n6524) );
  NANDN U10805 ( .A(n12626), .B(n6524), .Z(n6525) );
  NAND U10806 ( .A(n6526), .B(n6525), .Z(n6527) );
  NAND U10807 ( .A(n12624), .B(n6527), .Z(n6528) );
  ANDN U10808 ( .B(y[1190]), .A(x[1190]), .Z(n14569) );
  NANDN U10809 ( .A(y[1190]), .B(x[1190]), .Z(n6530) );
  NANDN U10810 ( .A(y[1191]), .B(x[1191]), .Z(n6529) );
  AND U10811 ( .A(n6530), .B(n6529), .Z(n22214) );
  NANDN U10812 ( .A(x[1192]), .B(y[1192]), .Z(n6532) );
  NANDN U10813 ( .A(x[1191]), .B(y[1191]), .Z(n6531) );
  NAND U10814 ( .A(n6532), .B(n6531), .Z(n22217) );
  NANDN U10815 ( .A(y[1192]), .B(x[1192]), .Z(n6534) );
  NANDN U10816 ( .A(y[1193]), .B(x[1193]), .Z(n6533) );
  AND U10817 ( .A(n6534), .B(n6533), .Z(n22218) );
  NANDN U10818 ( .A(x[1193]), .B(y[1193]), .Z(n12621) );
  IV U10819 ( .A(y[1194]), .Z(n14575) );
  NANDN U10820 ( .A(y[1196]), .B(x[1196]), .Z(n22226) );
  ANDN U10821 ( .B(x[1195]), .A(y[1195]), .Z(n14576) );
  NANDN U10822 ( .A(x[1196]), .B(y[1196]), .Z(n14580) );
  NANDN U10823 ( .A(x[1197]), .B(y[1197]), .Z(n14585) );
  NAND U10824 ( .A(n14580), .B(n14585), .Z(n22229) );
  NANDN U10825 ( .A(y[1197]), .B(x[1197]), .Z(n22230) );
  ANDN U10826 ( .B(x[1198]), .A(y[1198]), .Z(n14588) );
  NANDN U10827 ( .A(x[1200]), .B(y[1200]), .Z(n6539) );
  NANDN U10828 ( .A(x[1199]), .B(y[1199]), .Z(n6535) );
  NAND U10829 ( .A(n6539), .B(n6535), .Z(n14590) );
  NANDN U10830 ( .A(x[1198]), .B(y[1198]), .Z(n6536) );
  NANDN U10831 ( .A(n14590), .B(n6536), .Z(n22232) );
  ANDN U10832 ( .B(n6538), .A(n6537), .Z(n6541) );
  NANDN U10833 ( .A(y[1199]), .B(x[1199]), .Z(n14587) );
  NANDN U10834 ( .A(n14587), .B(n6539), .Z(n6540) );
  AND U10835 ( .A(n6541), .B(n6540), .Z(n6544) );
  NANDN U10836 ( .A(x[1201]), .B(y[1201]), .Z(n6543) );
  NANDN U10837 ( .A(x[1202]), .B(y[1202]), .Z(n6542) );
  AND U10838 ( .A(n6543), .B(n6542), .Z(n22236) );
  NANDN U10839 ( .A(n6544), .B(n22236), .Z(n6547) );
  NANDN U10840 ( .A(y[1203]), .B(x[1203]), .Z(n6546) );
  NANDN U10841 ( .A(y[1202]), .B(x[1202]), .Z(n6545) );
  AND U10842 ( .A(n6546), .B(n6545), .Z(n22239) );
  NAND U10843 ( .A(n6547), .B(n22239), .Z(n6550) );
  NANDN U10844 ( .A(x[1203]), .B(y[1203]), .Z(n6549) );
  NANDN U10845 ( .A(x[1204]), .B(y[1204]), .Z(n6548) );
  AND U10846 ( .A(n6549), .B(n6548), .Z(n22240) );
  NAND U10847 ( .A(n6550), .B(n22240), .Z(n6551) );
  NANDN U10848 ( .A(n22243), .B(n6551), .Z(n6552) );
  NANDN U10849 ( .A(n12620), .B(n6552), .Z(n6553) );
  AND U10850 ( .A(n22246), .B(n6553), .Z(n6554) );
  ANDN U10851 ( .B(n6555), .A(n6554), .Z(n6556) );
  NANDN U10852 ( .A(y[1208]), .B(x[1208]), .Z(n22251) );
  NANDN U10853 ( .A(n6556), .B(n22251), .Z(n6557) );
  AND U10854 ( .A(n22252), .B(n6557), .Z(n6559) );
  NANDN U10855 ( .A(y[1209]), .B(x[1209]), .Z(n22255) );
  ANDN U10856 ( .B(x[1210]), .A(y[1210]), .Z(n12616) );
  ANDN U10857 ( .B(n22255), .A(n12616), .Z(n6558) );
  NANDN U10858 ( .A(n6559), .B(n6558), .Z(n6560) );
  AND U10859 ( .A(n22256), .B(n6560), .Z(n6561) );
  OR U10860 ( .A(n12617), .B(n6561), .Z(n6564) );
  NANDN U10861 ( .A(x[1212]), .B(y[1212]), .Z(n6563) );
  NANDN U10862 ( .A(x[1211]), .B(y[1211]), .Z(n6562) );
  NAND U10863 ( .A(n6563), .B(n6562), .Z(n22260) );
  ANDN U10864 ( .B(n6564), .A(n22260), .Z(n6567) );
  NANDN U10865 ( .A(y[1212]), .B(x[1212]), .Z(n6566) );
  NANDN U10866 ( .A(y[1213]), .B(x[1213]), .Z(n6565) );
  AND U10867 ( .A(n6566), .B(n6565), .Z(n22262) );
  NANDN U10868 ( .A(n6567), .B(n22262), .Z(n6570) );
  NANDN U10869 ( .A(x[1214]), .B(y[1214]), .Z(n6569) );
  NANDN U10870 ( .A(x[1213]), .B(y[1213]), .Z(n6568) );
  NAND U10871 ( .A(n6569), .B(n6568), .Z(n22265) );
  ANDN U10872 ( .B(n6570), .A(n22265), .Z(n6573) );
  NANDN U10873 ( .A(y[1214]), .B(x[1214]), .Z(n6572) );
  NANDN U10874 ( .A(y[1215]), .B(x[1215]), .Z(n6571) );
  AND U10875 ( .A(n6572), .B(n6571), .Z(n22266) );
  NANDN U10876 ( .A(x[1216]), .B(y[1216]), .Z(n6575) );
  NANDN U10877 ( .A(x[1215]), .B(y[1215]), .Z(n6574) );
  AND U10878 ( .A(n6575), .B(n6574), .Z(n22268) );
  NANDN U10879 ( .A(y[1216]), .B(x[1216]), .Z(n6577) );
  NANDN U10880 ( .A(y[1217]), .B(x[1217]), .Z(n6576) );
  AND U10881 ( .A(n6577), .B(n6576), .Z(n22271) );
  NANDN U10882 ( .A(x[1217]), .B(y[1217]), .Z(n6579) );
  NANDN U10883 ( .A(x[1218]), .B(y[1218]), .Z(n6578) );
  AND U10884 ( .A(n6579), .B(n6578), .Z(n22272) );
  NANDN U10885 ( .A(y[1219]), .B(x[1219]), .Z(n6581) );
  NANDN U10886 ( .A(y[1218]), .B(x[1218]), .Z(n6580) );
  NAND U10887 ( .A(n6581), .B(n6580), .Z(n22275) );
  ANDN U10888 ( .B(x[1222]), .A(y[1222]), .Z(n14622) );
  NANDN U10889 ( .A(x[1222]), .B(y[1222]), .Z(n6584) );
  NANDN U10890 ( .A(x[1223]), .B(y[1223]), .Z(n6582) );
  NANDN U10891 ( .A(n6583), .B(n6582), .Z(n14624) );
  ANDN U10892 ( .B(n6584), .A(n14624), .Z(n22280) );
  NANDN U10893 ( .A(x[1225]), .B(y[1225]), .Z(n6586) );
  NANDN U10894 ( .A(x[1226]), .B(y[1226]), .Z(n6585) );
  AND U10895 ( .A(n6586), .B(n6585), .Z(n22284) );
  NANDN U10896 ( .A(y[1227]), .B(x[1227]), .Z(n6588) );
  NANDN U10897 ( .A(y[1226]), .B(x[1226]), .Z(n6587) );
  NAND U10898 ( .A(n6588), .B(n6587), .Z(n22286) );
  NANDN U10899 ( .A(x[1227]), .B(y[1227]), .Z(n6590) );
  NANDN U10900 ( .A(x[1228]), .B(y[1228]), .Z(n6589) );
  AND U10901 ( .A(n6590), .B(n6589), .Z(n22288) );
  AND U10902 ( .A(n22294), .B(n6591), .Z(n6595) );
  ANDN U10903 ( .B(y[1230]), .A(x[1230]), .Z(n12611) );
  NANDN U10904 ( .A(x[1231]), .B(y[1231]), .Z(n22296) );
  NANDN U10905 ( .A(n12611), .B(n22296), .Z(n6592) );
  AND U10906 ( .A(n6593), .B(n6592), .Z(n6594) );
  OR U10907 ( .A(n6595), .B(n6594), .Z(n6596) );
  NANDN U10908 ( .A(n14636), .B(n6596), .Z(n6597) );
  NANDN U10909 ( .A(x[1232]), .B(y[1232]), .Z(n12609) );
  NANDN U10910 ( .A(x[1233]), .B(y[1233]), .Z(n14640) );
  NAND U10911 ( .A(n12609), .B(n14640), .Z(n22300) );
  ANDN U10912 ( .B(n6597), .A(n22300), .Z(n6599) );
  ANDN U10913 ( .B(x[1233]), .A(y[1233]), .Z(n14637) );
  IV U10914 ( .A(n14637), .Z(n22301) );
  ANDN U10915 ( .B(x[1234]), .A(y[1234]), .Z(n12608) );
  ANDN U10916 ( .B(n22301), .A(n12608), .Z(n6598) );
  NANDN U10917 ( .A(n6599), .B(n6598), .Z(n6600) );
  AND U10918 ( .A(n22304), .B(n6600), .Z(n6601) );
  NAND U10919 ( .A(n6602), .B(n6601), .Z(n6603) );
  NAND U10920 ( .A(n6604), .B(n6603), .Z(n6605) );
  ANDN U10921 ( .B(y[1236]), .A(x[1236]), .Z(n14644) );
  ANDN U10922 ( .B(n6605), .A(n14644), .Z(n6606) );
  NAND U10923 ( .A(n6607), .B(n6606), .Z(n6608) );
  NAND U10924 ( .A(n12605), .B(n6608), .Z(n6609) );
  ANDN U10925 ( .B(y[1238]), .A(x[1238]), .Z(n12604) );
  ANDN U10926 ( .B(n6609), .A(n12604), .Z(n6612) );
  NANDN U10927 ( .A(y[1238]), .B(x[1238]), .Z(n6611) );
  NANDN U10928 ( .A(y[1239]), .B(x[1239]), .Z(n6610) );
  AND U10929 ( .A(n6611), .B(n6610), .Z(n22314) );
  NANDN U10930 ( .A(n6612), .B(n22314), .Z(n6615) );
  NANDN U10931 ( .A(x[1240]), .B(y[1240]), .Z(n6614) );
  NANDN U10932 ( .A(x[1239]), .B(y[1239]), .Z(n6613) );
  NAND U10933 ( .A(n6614), .B(n6613), .Z(n22317) );
  ANDN U10934 ( .B(n6615), .A(n22317), .Z(n6616) );
  ANDN U10935 ( .B(n22318), .A(n6616), .Z(n6621) );
  NANDN U10936 ( .A(x[1242]), .B(y[1242]), .Z(n6618) );
  NANDN U10937 ( .A(x[1241]), .B(y[1241]), .Z(n6617) );
  AND U10938 ( .A(n6618), .B(n6617), .Z(n6620) );
  AND U10939 ( .A(n6620), .B(n6619), .Z(n22321) );
  NANDN U10940 ( .A(n6621), .B(n22321), .Z(n6622) );
  NANDN U10941 ( .A(n12602), .B(n6622), .Z(n6625) );
  NANDN U10942 ( .A(x[1245]), .B(y[1245]), .Z(n6624) );
  NANDN U10943 ( .A(x[1244]), .B(y[1244]), .Z(n6623) );
  AND U10944 ( .A(n6624), .B(n6623), .Z(n12598) );
  NAND U10945 ( .A(n6625), .B(n12598), .Z(n6626) );
  NANDN U10946 ( .A(n12601), .B(n6626), .Z(n6627) );
  NAND U10947 ( .A(n6628), .B(n6627), .Z(n6629) );
  NAND U10948 ( .A(n12597), .B(n6629), .Z(n6630) );
  NAND U10949 ( .A(n6631), .B(n6630), .Z(n6632) );
  NAND U10950 ( .A(n12596), .B(n6632), .Z(n6633) );
  ANDN U10951 ( .B(y[1248]), .A(x[1248]), .Z(n12595) );
  ANDN U10952 ( .B(n6633), .A(n12595), .Z(n6636) );
  NANDN U10953 ( .A(y[1248]), .B(x[1248]), .Z(n6635) );
  NANDN U10954 ( .A(y[1249]), .B(x[1249]), .Z(n6634) );
  AND U10955 ( .A(n6635), .B(n6634), .Z(n22330) );
  NANDN U10956 ( .A(n6636), .B(n22330), .Z(n6639) );
  NANDN U10957 ( .A(x[1250]), .B(y[1250]), .Z(n6638) );
  NANDN U10958 ( .A(x[1249]), .B(y[1249]), .Z(n6637) );
  NAND U10959 ( .A(n6638), .B(n6637), .Z(n22332) );
  ANDN U10960 ( .B(n6639), .A(n22332), .Z(n6642) );
  NANDN U10961 ( .A(y[1250]), .B(x[1250]), .Z(n6641) );
  NANDN U10962 ( .A(y[1251]), .B(x[1251]), .Z(n6640) );
  AND U10963 ( .A(n6641), .B(n6640), .Z(n22334) );
  NANDN U10964 ( .A(n6642), .B(n22334), .Z(n6645) );
  NANDN U10965 ( .A(x[1252]), .B(y[1252]), .Z(n6644) );
  NANDN U10966 ( .A(x[1251]), .B(y[1251]), .Z(n6643) );
  NAND U10967 ( .A(n6644), .B(n6643), .Z(n22337) );
  ANDN U10968 ( .B(n6645), .A(n22337), .Z(n6648) );
  NANDN U10969 ( .A(y[1252]), .B(x[1252]), .Z(n6647) );
  NANDN U10970 ( .A(y[1253]), .B(x[1253]), .Z(n6646) );
  AND U10971 ( .A(n6647), .B(n6646), .Z(n22338) );
  NANDN U10972 ( .A(n6648), .B(n22338), .Z(n6649) );
  NANDN U10973 ( .A(n12593), .B(n6649), .Z(n6652) );
  NANDN U10974 ( .A(y[1254]), .B(x[1254]), .Z(n6651) );
  AND U10975 ( .A(n6651), .B(n6650), .Z(n22342) );
  NAND U10976 ( .A(n6652), .B(n22342), .Z(n6653) );
  NANDN U10977 ( .A(n6654), .B(n6653), .Z(n6655) );
  NANDN U10978 ( .A(y[1256]), .B(x[1256]), .Z(n22346) );
  NAND U10979 ( .A(n6655), .B(n22346), .Z(n6656) );
  NANDN U10980 ( .A(x[1256]), .B(y[1256]), .Z(n14663) );
  ANDN U10981 ( .B(y[1257]), .A(x[1257]), .Z(n14668) );
  ANDN U10982 ( .B(n14663), .A(n14668), .Z(n22348) );
  NAND U10983 ( .A(n6656), .B(n22348), .Z(n6657) );
  NAND U10984 ( .A(n6658), .B(n6657), .Z(n6659) );
  ANDN U10985 ( .B(y[1258]), .A(x[1258]), .Z(n22352) );
  ANDN U10986 ( .B(n6659), .A(n22352), .Z(n6660) );
  NAND U10987 ( .A(n6661), .B(n6660), .Z(n6662) );
  NAND U10988 ( .A(n6663), .B(n6662), .Z(n6664) );
  ANDN U10989 ( .B(y[1260]), .A(x[1260]), .Z(n14673) );
  ANDN U10990 ( .B(n6664), .A(n14673), .Z(n6665) );
  NAND U10991 ( .A(n6666), .B(n6665), .Z(n6667) );
  NAND U10992 ( .A(n12588), .B(n6667), .Z(n6668) );
  ANDN U10993 ( .B(y[1262]), .A(x[1262]), .Z(n12587) );
  ANDN U10994 ( .B(n6668), .A(n12587), .Z(n6671) );
  NANDN U10995 ( .A(y[1262]), .B(x[1262]), .Z(n6670) );
  NANDN U10996 ( .A(y[1263]), .B(x[1263]), .Z(n6669) );
  AND U10997 ( .A(n6670), .B(n6669), .Z(n22362) );
  NANDN U10998 ( .A(n6671), .B(n22362), .Z(n6674) );
  NANDN U10999 ( .A(x[1264]), .B(y[1264]), .Z(n6673) );
  NANDN U11000 ( .A(x[1263]), .B(y[1263]), .Z(n6672) );
  NAND U11001 ( .A(n6673), .B(n6672), .Z(n22364) );
  ANDN U11002 ( .B(n6674), .A(n22364), .Z(n6677) );
  NANDN U11003 ( .A(y[1264]), .B(x[1264]), .Z(n6676) );
  NANDN U11004 ( .A(y[1265]), .B(x[1265]), .Z(n6675) );
  AND U11005 ( .A(n6676), .B(n6675), .Z(n22366) );
  NANDN U11006 ( .A(n6677), .B(n22366), .Z(n6678) );
  NANDN U11007 ( .A(n14680), .B(n6678), .Z(n6679) );
  NANDN U11008 ( .A(n12585), .B(n6679), .Z(n6680) );
  AND U11009 ( .A(n22372), .B(n6680), .Z(n6681) );
  NANDN U11010 ( .A(n14681), .B(n6681), .Z(n6682) );
  NANDN U11011 ( .A(n12584), .B(n6682), .Z(n6683) );
  NANDN U11012 ( .A(y[1268]), .B(x[1268]), .Z(n22374) );
  NANDN U11013 ( .A(n6683), .B(n22374), .Z(n6684) );
  ANDN U11014 ( .B(y[1269]), .A(x[1269]), .Z(n12583) );
  ANDN U11015 ( .B(y[1268]), .A(x[1268]), .Z(n14684) );
  NOR U11016 ( .A(n12583), .B(n14684), .Z(n22376) );
  NAND U11017 ( .A(n6684), .B(n22376), .Z(n6685) );
  ANDN U11018 ( .B(x[1269]), .A(y[1269]), .Z(n22378) );
  ANDN U11019 ( .B(n6685), .A(n22378), .Z(n6686) );
  NANDN U11020 ( .A(n12582), .B(n6686), .Z(n6687) );
  NANDN U11021 ( .A(x[1270]), .B(y[1270]), .Z(n22380) );
  AND U11022 ( .A(n6687), .B(n22380), .Z(n6689) );
  IV U11023 ( .A(x[1271]), .Z(n14692) );
  NANDN U11024 ( .A(n6689), .B(n14692), .Z(n6688) );
  ANDN U11025 ( .B(y[1272]), .A(x[1272]), .Z(n14694) );
  ANDN U11026 ( .B(n6688), .A(n14694), .Z(n6692) );
  XOR U11027 ( .A(x[1271]), .B(n6689), .Z(n6690) );
  NAND U11028 ( .A(n6690), .B(y[1271]), .Z(n6691) );
  NAND U11029 ( .A(n6692), .B(n6691), .Z(n6693) );
  ANDN U11030 ( .B(x[1272]), .A(y[1272]), .Z(n12580) );
  ANDN U11031 ( .B(n6693), .A(n12580), .Z(n6694) );
  IV U11032 ( .A(y[1273]), .Z(n12578) );
  NANDN U11033 ( .A(n6694), .B(n12578), .Z(n6697) );
  XOR U11034 ( .A(y[1273]), .B(n6694), .Z(n6695) );
  NAND U11035 ( .A(n6695), .B(x[1273]), .Z(n6696) );
  NAND U11036 ( .A(n6697), .B(n6696), .Z(n6698) );
  ANDN U11037 ( .B(y[1274]), .A(x[1274]), .Z(n12577) );
  ANDN U11038 ( .B(n6698), .A(n12577), .Z(n6701) );
  NANDN U11039 ( .A(y[1274]), .B(x[1274]), .Z(n6700) );
  NANDN U11040 ( .A(y[1275]), .B(x[1275]), .Z(n6699) );
  AND U11041 ( .A(n6700), .B(n6699), .Z(n22390) );
  NANDN U11042 ( .A(n6701), .B(n22390), .Z(n6704) );
  NANDN U11043 ( .A(x[1276]), .B(y[1276]), .Z(n6703) );
  NANDN U11044 ( .A(x[1275]), .B(y[1275]), .Z(n6702) );
  NAND U11045 ( .A(n6703), .B(n6702), .Z(n22392) );
  ANDN U11046 ( .B(n6704), .A(n22392), .Z(n6707) );
  NANDN U11047 ( .A(y[1276]), .B(x[1276]), .Z(n6706) );
  NANDN U11048 ( .A(y[1277]), .B(x[1277]), .Z(n6705) );
  AND U11049 ( .A(n6706), .B(n6705), .Z(n22394) );
  NANDN U11050 ( .A(n6707), .B(n22394), .Z(n6708) );
  NANDN U11051 ( .A(n14702), .B(n6708), .Z(n6709) );
  NANDN U11052 ( .A(n22399), .B(n6709), .Z(n6714) );
  NANDN U11053 ( .A(x[1278]), .B(y[1278]), .Z(n14701) );
  NANDN U11054 ( .A(y[1279]), .B(n14701), .Z(n6712) );
  XNOR U11055 ( .A(y[1279]), .B(n14701), .Z(n6710) );
  NAND U11056 ( .A(n6710), .B(x[1279]), .Z(n6711) );
  NAND U11057 ( .A(n6712), .B(n6711), .Z(n6713) );
  AND U11058 ( .A(n6714), .B(n6713), .Z(n6715) );
  OR U11059 ( .A(n12573), .B(n6715), .Z(n6716) );
  NANDN U11060 ( .A(n14706), .B(n6716), .Z(n6717) );
  AND U11061 ( .A(n12572), .B(n6717), .Z(n6718) );
  NANDN U11062 ( .A(n12571), .B(n6718), .Z(n6719) );
  AND U11063 ( .A(n22404), .B(n6719), .Z(n6720) );
  NAND U11064 ( .A(n6721), .B(n6720), .Z(n6722) );
  NAND U11065 ( .A(n6723), .B(n6722), .Z(n6724) );
  ANDN U11066 ( .B(y[1284]), .A(x[1284]), .Z(n12569) );
  ANDN U11067 ( .B(n6724), .A(n12569), .Z(n6725) );
  NAND U11068 ( .A(n6726), .B(n6725), .Z(n6727) );
  NAND U11069 ( .A(n12567), .B(n6727), .Z(n6728) );
  ANDN U11070 ( .B(y[1286]), .A(x[1286]), .Z(n14714) );
  ANDN U11071 ( .B(n6728), .A(n14714), .Z(n6731) );
  NANDN U11072 ( .A(y[1286]), .B(x[1286]), .Z(n6730) );
  NANDN U11073 ( .A(y[1287]), .B(x[1287]), .Z(n6729) );
  AND U11074 ( .A(n6730), .B(n6729), .Z(n22414) );
  NANDN U11075 ( .A(n6731), .B(n22414), .Z(n6734) );
  NANDN U11076 ( .A(x[1288]), .B(y[1288]), .Z(n6733) );
  NANDN U11077 ( .A(x[1287]), .B(y[1287]), .Z(n6732) );
  NAND U11078 ( .A(n6733), .B(n6732), .Z(n22417) );
  ANDN U11079 ( .B(n6734), .A(n22417), .Z(n6735) );
  OR U11080 ( .A(n22419), .B(n6735), .Z(n6736) );
  ANDN U11081 ( .B(y[1289]), .A(x[1289]), .Z(n12565) );
  ANDN U11082 ( .B(n6736), .A(n12565), .Z(n6738) );
  IV U11083 ( .A(x[1290]), .Z(n12563) );
  NANDN U11084 ( .A(n6738), .B(n12563), .Z(n6737) );
  AND U11085 ( .A(n22424), .B(n6737), .Z(n6741) );
  XOR U11086 ( .A(x[1290]), .B(n6738), .Z(n6739) );
  NAND U11087 ( .A(n6739), .B(y[1290]), .Z(n6740) );
  NAND U11088 ( .A(n6741), .B(n6740), .Z(n6742) );
  ANDN U11089 ( .B(x[1291]), .A(y[1291]), .Z(n12562) );
  ANDN U11090 ( .B(n6742), .A(n12562), .Z(n6743) );
  NANDN U11091 ( .A(y[1292]), .B(x[1292]), .Z(n22426) );
  NAND U11092 ( .A(n6743), .B(n22426), .Z(n6744) );
  ANDN U11093 ( .B(y[1293]), .A(x[1293]), .Z(n12560) );
  ANDN U11094 ( .B(y[1292]), .A(x[1292]), .Z(n14721) );
  NOR U11095 ( .A(n12560), .B(n14721), .Z(n22428) );
  NAND U11096 ( .A(n6744), .B(n22428), .Z(n6745) );
  AND U11097 ( .A(n22430), .B(n6745), .Z(n6746) );
  NANDN U11098 ( .A(n12558), .B(n6746), .Z(n6747) );
  NANDN U11099 ( .A(x[1294]), .B(y[1294]), .Z(n22432) );
  NAND U11100 ( .A(n6747), .B(n22432), .Z(n6748) );
  NANDN U11101 ( .A(n12559), .B(n6748), .Z(n6751) );
  NANDN U11102 ( .A(x[1296]), .B(y[1296]), .Z(n6750) );
  NANDN U11103 ( .A(x[1295]), .B(y[1295]), .Z(n6749) );
  AND U11104 ( .A(n6750), .B(n6749), .Z(n22436) );
  NAND U11105 ( .A(n6751), .B(n22436), .Z(n6754) );
  NANDN U11106 ( .A(y[1296]), .B(x[1296]), .Z(n6753) );
  NANDN U11107 ( .A(y[1297]), .B(x[1297]), .Z(n6752) );
  AND U11108 ( .A(n6753), .B(n6752), .Z(n22439) );
  NAND U11109 ( .A(n6754), .B(n22439), .Z(n6755) );
  AND U11110 ( .A(n22440), .B(n6755), .Z(n6758) );
  NANDN U11111 ( .A(y[1298]), .B(x[1298]), .Z(n6757) );
  NANDN U11112 ( .A(y[1299]), .B(x[1299]), .Z(n6756) );
  AND U11113 ( .A(n6757), .B(n6756), .Z(n22443) );
  NANDN U11114 ( .A(n6758), .B(n22443), .Z(n6761) );
  NANDN U11115 ( .A(x[1300]), .B(y[1300]), .Z(n6760) );
  NANDN U11116 ( .A(x[1299]), .B(y[1299]), .Z(n6759) );
  AND U11117 ( .A(n6760), .B(n6759), .Z(n22444) );
  NAND U11118 ( .A(n6761), .B(n22444), .Z(n6764) );
  NANDN U11119 ( .A(y[1300]), .B(x[1300]), .Z(n6763) );
  NANDN U11120 ( .A(y[1301]), .B(x[1301]), .Z(n6762) );
  AND U11121 ( .A(n6763), .B(n6762), .Z(n22446) );
  NAND U11122 ( .A(n6764), .B(n22446), .Z(n6765) );
  NANDN U11123 ( .A(n14736), .B(n6765), .Z(n6766) );
  AND U11124 ( .A(n22450), .B(n6766), .Z(n6767) );
  ANDN U11125 ( .B(n12556), .A(n6767), .Z(n6770) );
  XNOR U11126 ( .A(y[1303]), .B(x[1303]), .Z(n6768) );
  ANDN U11127 ( .B(y[1302]), .A(x[1302]), .Z(n14735) );
  NAND U11128 ( .A(n6768), .B(n14735), .Z(n6769) );
  NAND U11129 ( .A(n6770), .B(n6769), .Z(n6771) );
  NAND U11130 ( .A(n12552), .B(n6771), .Z(n6772) );
  NANDN U11131 ( .A(n12557), .B(n6772), .Z(n6773) );
  ANDN U11132 ( .B(x[1306]), .A(y[1306]), .Z(n12551) );
  ANDN U11133 ( .B(n6773), .A(n12551), .Z(n6774) );
  NANDN U11134 ( .A(n12553), .B(n6774), .Z(n6775) );
  NANDN U11135 ( .A(x[1306]), .B(y[1306]), .Z(n22456) );
  NAND U11136 ( .A(n6775), .B(n22456), .Z(n6776) );
  NAND U11137 ( .A(n6777), .B(n6776), .Z(n6778) );
  NAND U11138 ( .A(n14744), .B(n6778), .Z(n6779) );
  NAND U11139 ( .A(n6780), .B(n6779), .Z(n6781) );
  NAND U11140 ( .A(n14743), .B(n6781), .Z(n6782) );
  ANDN U11141 ( .B(x[1309]), .A(y[1309]), .Z(n12548) );
  NANDN U11142 ( .A(x[1309]), .B(y[1309]), .Z(n6784) );
  NANDN U11143 ( .A(x[1310]), .B(y[1310]), .Z(n6783) );
  AND U11144 ( .A(n6784), .B(n6783), .Z(n22465) );
  NANDN U11145 ( .A(x[1311]), .B(y[1311]), .Z(n6786) );
  NANDN U11146 ( .A(x[1312]), .B(y[1312]), .Z(n6785) );
  AND U11147 ( .A(n6786), .B(n6785), .Z(n22468) );
  NANDN U11148 ( .A(y[1313]), .B(x[1313]), .Z(n6788) );
  NANDN U11149 ( .A(y[1312]), .B(x[1312]), .Z(n6787) );
  AND U11150 ( .A(n6788), .B(n6787), .Z(n22470) );
  NANDN U11151 ( .A(y[1314]), .B(x[1314]), .Z(n6790) );
  AND U11152 ( .A(n6790), .B(n6789), .Z(n22475) );
  NANDN U11153 ( .A(x[1317]), .B(y[1317]), .Z(n14758) );
  ANDN U11154 ( .B(y[1316]), .A(x[1316]), .Z(n12545) );
  ANDN U11155 ( .B(n14758), .A(n12545), .Z(n22480) );
  ANDN U11156 ( .B(x[1318]), .A(y[1318]), .Z(n12543) );
  NANDN U11157 ( .A(y[1317]), .B(x[1317]), .Z(n22482) );
  NANDN U11158 ( .A(x[1318]), .B(y[1318]), .Z(n22484) );
  IV U11159 ( .A(y[1319]), .Z(n12542) );
  ANDN U11160 ( .B(y[1322]), .A(x[1322]), .Z(n12537) );
  NANDN U11161 ( .A(y[1323]), .B(x[1323]), .Z(n6793) );
  NANDN U11162 ( .A(y[1322]), .B(x[1322]), .Z(n6792) );
  NAND U11163 ( .A(n6793), .B(n6792), .Z(n22494) );
  NANDN U11164 ( .A(x[1323]), .B(y[1323]), .Z(n6795) );
  NANDN U11165 ( .A(x[1324]), .B(y[1324]), .Z(n6794) );
  AND U11166 ( .A(n6795), .B(n6794), .Z(n22496) );
  NANDN U11167 ( .A(y[1326]), .B(x[1326]), .Z(n6797) );
  AND U11168 ( .A(n6797), .B(n6796), .Z(n22502) );
  ANDN U11169 ( .B(y[1328]), .A(x[1328]), .Z(n12535) );
  NANDN U11170 ( .A(y[1329]), .B(x[1329]), .Z(n20287) );
  NAND U11171 ( .A(n6798), .B(n20287), .Z(n6799) );
  NAND U11172 ( .A(n6800), .B(n6799), .Z(n6801) );
  NAND U11173 ( .A(n12532), .B(n6801), .Z(n6802) );
  NAND U11174 ( .A(n6803), .B(n6802), .Z(n6804) );
  NAND U11175 ( .A(n12531), .B(n6804), .Z(n6805) );
  ANDN U11176 ( .B(y[1332]), .A(x[1332]), .Z(n14779) );
  ANDN U11177 ( .B(n6805), .A(n14779), .Z(n6808) );
  NANDN U11178 ( .A(y[1332]), .B(x[1332]), .Z(n6807) );
  NANDN U11179 ( .A(y[1333]), .B(x[1333]), .Z(n6806) );
  AND U11180 ( .A(n6807), .B(n6806), .Z(n22516) );
  NANDN U11181 ( .A(n6808), .B(n22516), .Z(n6811) );
  NANDN U11182 ( .A(x[1334]), .B(y[1334]), .Z(n6810) );
  NANDN U11183 ( .A(x[1333]), .B(y[1333]), .Z(n6809) );
  NAND U11184 ( .A(n6810), .B(n6809), .Z(n22518) );
  ANDN U11185 ( .B(n6811), .A(n22518), .Z(n6814) );
  NANDN U11186 ( .A(y[1334]), .B(x[1334]), .Z(n6813) );
  NANDN U11187 ( .A(y[1335]), .B(x[1335]), .Z(n6812) );
  AND U11188 ( .A(n6813), .B(n6812), .Z(n22520) );
  NANDN U11189 ( .A(n6814), .B(n22520), .Z(n6817) );
  NANDN U11190 ( .A(x[1336]), .B(y[1336]), .Z(n6816) );
  NANDN U11191 ( .A(x[1335]), .B(y[1335]), .Z(n6815) );
  NAND U11192 ( .A(n6816), .B(n6815), .Z(n22522) );
  ANDN U11193 ( .B(n6817), .A(n22522), .Z(n6820) );
  NANDN U11194 ( .A(y[1336]), .B(x[1336]), .Z(n6819) );
  NANDN U11195 ( .A(y[1337]), .B(x[1337]), .Z(n6818) );
  AND U11196 ( .A(n6819), .B(n6818), .Z(n22524) );
  NANDN U11197 ( .A(n6820), .B(n22524), .Z(n6821) );
  NANDN U11198 ( .A(n14787), .B(n6821), .Z(n6824) );
  NANDN U11199 ( .A(y[1338]), .B(x[1338]), .Z(n6823) );
  ANDN U11200 ( .B(n6823), .A(n6822), .Z(n22528) );
  NAND U11201 ( .A(n6824), .B(n22528), .Z(n6825) );
  NAND U11202 ( .A(n6826), .B(n6825), .Z(n6827) );
  NANDN U11203 ( .A(n14792), .B(n6827), .Z(n6828) );
  NAND U11204 ( .A(n12530), .B(n6828), .Z(n6829) );
  ANDN U11205 ( .B(x[1342]), .A(y[1342]), .Z(n12529) );
  ANDN U11206 ( .B(n6829), .A(n12529), .Z(n6830) );
  NANDN U11207 ( .A(n22535), .B(n6830), .Z(n6831) );
  AND U11208 ( .A(n22538), .B(n6831), .Z(n6832) );
  NAND U11209 ( .A(n6833), .B(n6832), .Z(n6834) );
  NAND U11210 ( .A(n6835), .B(n6834), .Z(n6836) );
  ANDN U11211 ( .B(y[1344]), .A(x[1344]), .Z(n12527) );
  ANDN U11212 ( .B(n6836), .A(n12527), .Z(n6837) );
  NAND U11213 ( .A(n6838), .B(n6837), .Z(n6839) );
  NAND U11214 ( .A(n14800), .B(n6839), .Z(n6840) );
  ANDN U11215 ( .B(y[1346]), .A(x[1346]), .Z(n12525) );
  ANDN U11216 ( .B(n6840), .A(n12525), .Z(n6843) );
  NANDN U11217 ( .A(y[1347]), .B(x[1347]), .Z(n6842) );
  NANDN U11218 ( .A(y[1346]), .B(x[1346]), .Z(n6841) );
  AND U11219 ( .A(n6842), .B(n6841), .Z(n22548) );
  NANDN U11220 ( .A(n6843), .B(n22548), .Z(n6844) );
  ANDN U11221 ( .B(y[1348]), .A(x[1348]), .Z(n12520) );
  ANDN U11222 ( .B(n6844), .A(n12520), .Z(n6845) );
  NANDN U11223 ( .A(x[1347]), .B(y[1347]), .Z(n22551) );
  NAND U11224 ( .A(n6845), .B(n22551), .Z(n6847) );
  NANDN U11225 ( .A(y[1348]), .B(x[1348]), .Z(n6846) );
  ANDN U11226 ( .B(x[1349]), .A(y[1349]), .Z(n12521) );
  ANDN U11227 ( .B(n6846), .A(n12521), .Z(n22552) );
  NAND U11228 ( .A(n6847), .B(n22552), .Z(n6848) );
  NANDN U11229 ( .A(n12523), .B(n6848), .Z(n6849) );
  NANDN U11230 ( .A(n12518), .B(n6849), .Z(n6852) );
  NANDN U11231 ( .A(x[1352]), .B(y[1352]), .Z(n6851) );
  NANDN U11232 ( .A(x[1353]), .B(y[1353]), .Z(n6850) );
  NAND U11233 ( .A(n6851), .B(n6850), .Z(n12515) );
  ANDN U11234 ( .B(n6852), .A(n12515), .Z(n6853) );
  OR U11235 ( .A(n12519), .B(n6853), .Z(n6854) );
  NAND U11236 ( .A(n6855), .B(n6854), .Z(n6856) );
  NAND U11237 ( .A(n12514), .B(n6856), .Z(n6857) );
  NAND U11238 ( .A(n6858), .B(n6857), .Z(n6859) );
  NAND U11239 ( .A(n12513), .B(n6859), .Z(n6860) );
  ANDN U11240 ( .B(y[1356]), .A(x[1356]), .Z(n14811) );
  ANDN U11241 ( .B(n6860), .A(n14811), .Z(n6863) );
  NANDN U11242 ( .A(y[1356]), .B(x[1356]), .Z(n6862) );
  NANDN U11243 ( .A(y[1357]), .B(x[1357]), .Z(n6861) );
  AND U11244 ( .A(n6862), .B(n6861), .Z(n22564) );
  NANDN U11245 ( .A(n6863), .B(n22564), .Z(n6866) );
  NANDN U11246 ( .A(x[1358]), .B(y[1358]), .Z(n6865) );
  NANDN U11247 ( .A(x[1357]), .B(y[1357]), .Z(n6864) );
  NAND U11248 ( .A(n6865), .B(n6864), .Z(n22566) );
  ANDN U11249 ( .B(n6866), .A(n22566), .Z(n6869) );
  NANDN U11250 ( .A(y[1358]), .B(x[1358]), .Z(n6868) );
  NANDN U11251 ( .A(y[1359]), .B(x[1359]), .Z(n6867) );
  AND U11252 ( .A(n6868), .B(n6867), .Z(n22568) );
  NANDN U11253 ( .A(n6869), .B(n22568), .Z(n6872) );
  NANDN U11254 ( .A(x[1360]), .B(y[1360]), .Z(n6871) );
  NANDN U11255 ( .A(x[1359]), .B(y[1359]), .Z(n6870) );
  NAND U11256 ( .A(n6871), .B(n6870), .Z(n22570) );
  ANDN U11257 ( .B(n6872), .A(n22570), .Z(n6875) );
  NANDN U11258 ( .A(y[1360]), .B(x[1360]), .Z(n6874) );
  NANDN U11259 ( .A(y[1361]), .B(x[1361]), .Z(n6873) );
  AND U11260 ( .A(n6874), .B(n6873), .Z(n22572) );
  NANDN U11261 ( .A(n6875), .B(n22572), .Z(n6876) );
  NANDN U11262 ( .A(n22575), .B(n6876), .Z(n6879) );
  NANDN U11263 ( .A(y[1363]), .B(x[1363]), .Z(n6878) );
  NANDN U11264 ( .A(y[1362]), .B(x[1362]), .Z(n6877) );
  AND U11265 ( .A(n6878), .B(n6877), .Z(n22576) );
  NAND U11266 ( .A(n6879), .B(n22576), .Z(n6880) );
  NANDN U11267 ( .A(x[1363]), .B(y[1363]), .Z(n22578) );
  NAND U11268 ( .A(n6880), .B(n22578), .Z(n6881) );
  NANDN U11269 ( .A(y[1364]), .B(x[1364]), .Z(n22580) );
  NAND U11270 ( .A(n6881), .B(n22580), .Z(n6882) );
  ANDN U11271 ( .B(y[1365]), .A(x[1365]), .Z(n14826) );
  ANDN U11272 ( .B(y[1364]), .A(x[1364]), .Z(n12512) );
  NOR U11273 ( .A(n14826), .B(n12512), .Z(n22583) );
  NAND U11274 ( .A(n6882), .B(n22583), .Z(n6883) );
  ANDN U11275 ( .B(x[1366]), .A(y[1366]), .Z(n14828) );
  ANDN U11276 ( .B(n6883), .A(n14828), .Z(n6884) );
  NANDN U11277 ( .A(y[1365]), .B(x[1365]), .Z(n22584) );
  NAND U11278 ( .A(n6884), .B(n22584), .Z(n6887) );
  NANDN U11279 ( .A(x[1366]), .B(y[1366]), .Z(n6886) );
  NANDN U11280 ( .A(x[1368]), .B(y[1368]), .Z(n6892) );
  NANDN U11281 ( .A(x[1367]), .B(y[1367]), .Z(n6885) );
  NAND U11282 ( .A(n6892), .B(n6885), .Z(n14830) );
  ANDN U11283 ( .B(n6886), .A(n14830), .Z(n22586) );
  NAND U11284 ( .A(n6887), .B(n22586), .Z(n6891) );
  NANDN U11285 ( .A(y[1369]), .B(x[1369]), .Z(n6889) );
  NANDN U11286 ( .A(y[1368]), .B(x[1368]), .Z(n6888) );
  NAND U11287 ( .A(n6889), .B(n6888), .Z(n14831) );
  IV U11288 ( .A(n14831), .Z(n6890) );
  AND U11289 ( .A(n6891), .B(n6890), .Z(n6894) );
  NANDN U11290 ( .A(y[1367]), .B(x[1367]), .Z(n14827) );
  NANDN U11291 ( .A(n14827), .B(n6892), .Z(n6893) );
  AND U11292 ( .A(n6894), .B(n6893), .Z(n6897) );
  NANDN U11293 ( .A(x[1369]), .B(y[1369]), .Z(n6896) );
  NANDN U11294 ( .A(x[1370]), .B(y[1370]), .Z(n6895) );
  AND U11295 ( .A(n6896), .B(n6895), .Z(n22590) );
  NANDN U11296 ( .A(n6897), .B(n22590), .Z(n6900) );
  NANDN U11297 ( .A(y[1371]), .B(x[1371]), .Z(n6899) );
  NANDN U11298 ( .A(y[1370]), .B(x[1370]), .Z(n6898) );
  NAND U11299 ( .A(n6899), .B(n6898), .Z(n22593) );
  ANDN U11300 ( .B(n6900), .A(n22593), .Z(n6903) );
  NANDN U11301 ( .A(x[1371]), .B(y[1371]), .Z(n6902) );
  NANDN U11302 ( .A(x[1372]), .B(y[1372]), .Z(n6901) );
  AND U11303 ( .A(n6902), .B(n6901), .Z(n22594) );
  NANDN U11304 ( .A(n6903), .B(n22594), .Z(n6906) );
  NANDN U11305 ( .A(y[1373]), .B(x[1373]), .Z(n6905) );
  NANDN U11306 ( .A(y[1372]), .B(x[1372]), .Z(n6904) );
  NAND U11307 ( .A(n6905), .B(n6904), .Z(n22597) );
  ANDN U11308 ( .B(n6906), .A(n22597), .Z(n6911) );
  NANDN U11309 ( .A(x[1374]), .B(y[1374]), .Z(n6908) );
  NANDN U11310 ( .A(x[1373]), .B(y[1373]), .Z(n6907) );
  AND U11311 ( .A(n6908), .B(n6907), .Z(n6910) );
  AND U11312 ( .A(n6910), .B(n6909), .Z(n22598) );
  NANDN U11313 ( .A(n6911), .B(n22598), .Z(n6912) );
  NANDN U11314 ( .A(n12511), .B(n6912), .Z(n6915) );
  NANDN U11315 ( .A(x[1377]), .B(y[1377]), .Z(n6914) );
  NANDN U11316 ( .A(x[1376]), .B(y[1376]), .Z(n6913) );
  AND U11317 ( .A(n6914), .B(n6913), .Z(n12507) );
  NAND U11318 ( .A(n6915), .B(n12507), .Z(n6916) );
  ANDN U11319 ( .B(x[1377]), .A(y[1377]), .Z(n12510) );
  ANDN U11320 ( .B(n6916), .A(n12510), .Z(n6917) );
  NAND U11321 ( .A(n6918), .B(n6917), .Z(n6919) );
  NAND U11322 ( .A(n6920), .B(n6919), .Z(n6921) );
  ANDN U11323 ( .B(x[1379]), .A(y[1379]), .Z(n12506) );
  ANDN U11324 ( .B(n6921), .A(n12506), .Z(n6922) );
  NAND U11325 ( .A(n6923), .B(n6922), .Z(n6924) );
  NAND U11326 ( .A(n12503), .B(n6924), .Z(n6925) );
  ANDN U11327 ( .B(x[1381]), .A(y[1381]), .Z(n14844) );
  ANDN U11328 ( .B(n6925), .A(n14844), .Z(n6928) );
  NANDN U11329 ( .A(x[1381]), .B(y[1381]), .Z(n6927) );
  NANDN U11330 ( .A(x[1382]), .B(y[1382]), .Z(n6926) );
  AND U11331 ( .A(n6927), .B(n6926), .Z(n22610) );
  NANDN U11332 ( .A(n6928), .B(n22610), .Z(n6931) );
  NANDN U11333 ( .A(y[1383]), .B(x[1383]), .Z(n6930) );
  NANDN U11334 ( .A(y[1382]), .B(x[1382]), .Z(n6929) );
  NAND U11335 ( .A(n6930), .B(n6929), .Z(n22613) );
  ANDN U11336 ( .B(n6931), .A(n22613), .Z(n6934) );
  NANDN U11337 ( .A(x[1383]), .B(y[1383]), .Z(n6933) );
  NANDN U11338 ( .A(x[1384]), .B(y[1384]), .Z(n6932) );
  AND U11339 ( .A(n6933), .B(n6932), .Z(n22614) );
  NANDN U11340 ( .A(n6934), .B(n22614), .Z(n6937) );
  NANDN U11341 ( .A(y[1385]), .B(x[1385]), .Z(n6936) );
  NANDN U11342 ( .A(y[1384]), .B(x[1384]), .Z(n6935) );
  AND U11343 ( .A(n6936), .B(n6935), .Z(n22616) );
  NAND U11344 ( .A(n6937), .B(n22616), .Z(n6942) );
  NANDN U11345 ( .A(x[1386]), .B(y[1386]), .Z(n6939) );
  NANDN U11346 ( .A(x[1385]), .B(y[1385]), .Z(n6938) );
  AND U11347 ( .A(n6939), .B(n6938), .Z(n6941) );
  NANDN U11348 ( .A(x[1387]), .B(y[1387]), .Z(n6940) );
  AND U11349 ( .A(n6941), .B(n6940), .Z(n22619) );
  NAND U11350 ( .A(n6942), .B(n22619), .Z(n6943) );
  NANDN U11351 ( .A(n22621), .B(n6943), .Z(n6948) );
  XNOR U11352 ( .A(y[1389]), .B(x[1389]), .Z(n6945) );
  NANDN U11353 ( .A(x[1388]), .B(y[1388]), .Z(n6944) );
  NAND U11354 ( .A(n6945), .B(n6944), .Z(n6946) );
  AND U11355 ( .A(n6947), .B(n6946), .Z(n12502) );
  ANDN U11356 ( .B(n6948), .A(n12502), .Z(n6950) );
  XNOR U11357 ( .A(y[1390]), .B(x[1390]), .Z(n6949) );
  NANDN U11358 ( .A(n6950), .B(n6949), .Z(n6951) );
  NAND U11359 ( .A(n6952), .B(n6951), .Z(n6953) );
  ANDN U11360 ( .B(x[1391]), .A(y[1391]), .Z(n14854) );
  ANDN U11361 ( .B(n6953), .A(n14854), .Z(n6954) );
  NAND U11362 ( .A(n6955), .B(n6954), .Z(n6956) );
  NAND U11363 ( .A(n6957), .B(n6956), .Z(n6958) );
  ANDN U11364 ( .B(x[1393]), .A(y[1393]), .Z(n12498) );
  ANDN U11365 ( .B(n6958), .A(n12498), .Z(n6959) );
  NAND U11366 ( .A(n6960), .B(n6959), .Z(n6961) );
  NAND U11367 ( .A(n12495), .B(n6961), .Z(n6962) );
  ANDN U11368 ( .B(x[1395]), .A(y[1395]), .Z(n12494) );
  ANDN U11369 ( .B(n6962), .A(n12494), .Z(n6965) );
  NANDN U11370 ( .A(x[1395]), .B(y[1395]), .Z(n6964) );
  NANDN U11371 ( .A(x[1396]), .B(y[1396]), .Z(n6963) );
  AND U11372 ( .A(n6964), .B(n6963), .Z(n22634) );
  NANDN U11373 ( .A(n6965), .B(n22634), .Z(n6968) );
  NANDN U11374 ( .A(y[1397]), .B(x[1397]), .Z(n6967) );
  NANDN U11375 ( .A(y[1396]), .B(x[1396]), .Z(n6966) );
  AND U11376 ( .A(n6967), .B(n6966), .Z(n22636) );
  NAND U11377 ( .A(n6968), .B(n22636), .Z(n6971) );
  NANDN U11378 ( .A(x[1398]), .B(y[1398]), .Z(n6970) );
  NANDN U11379 ( .A(x[1397]), .B(y[1397]), .Z(n6969) );
  NAND U11380 ( .A(n6970), .B(n6969), .Z(n14863) );
  NOR U11381 ( .A(n14867), .B(n14863), .Z(n22638) );
  NAND U11382 ( .A(n6971), .B(n22638), .Z(n6972) );
  NANDN U11383 ( .A(n22641), .B(n6972), .Z(n6973) );
  NANDN U11384 ( .A(n22642), .B(n6973), .Z(n6974) );
  NANDN U11385 ( .A(y[1401]), .B(x[1401]), .Z(n22644) );
  NAND U11386 ( .A(n6974), .B(n22644), .Z(n6975) );
  OR U11387 ( .A(n12492), .B(n6975), .Z(n6976) );
  NAND U11388 ( .A(n6977), .B(n6976), .Z(n6978) );
  ANDN U11389 ( .B(x[1403]), .A(y[1403]), .Z(n12491) );
  ANDN U11390 ( .B(n6978), .A(n12491), .Z(n6979) );
  NAND U11391 ( .A(n6980), .B(n6979), .Z(n6981) );
  NAND U11392 ( .A(n12490), .B(n6981), .Z(n6982) );
  ANDN U11393 ( .B(x[1405]), .A(y[1405]), .Z(n12488) );
  ANDN U11394 ( .B(n6982), .A(n12488), .Z(n6985) );
  NANDN U11395 ( .A(x[1405]), .B(y[1405]), .Z(n6984) );
  NANDN U11396 ( .A(x[1406]), .B(y[1406]), .Z(n6983) );
  AND U11397 ( .A(n6984), .B(n6983), .Z(n22654) );
  NANDN U11398 ( .A(n6985), .B(n22654), .Z(n6986) );
  NANDN U11399 ( .A(n22657), .B(n6986), .Z(n6989) );
  NANDN U11400 ( .A(x[1407]), .B(y[1407]), .Z(n6988) );
  NANDN U11401 ( .A(x[1408]), .B(y[1408]), .Z(n6987) );
  AND U11402 ( .A(n6988), .B(n6987), .Z(n22658) );
  NAND U11403 ( .A(n6989), .B(n22658), .Z(n6992) );
  NANDN U11404 ( .A(y[1409]), .B(x[1409]), .Z(n6991) );
  NANDN U11405 ( .A(y[1408]), .B(x[1408]), .Z(n6990) );
  NAND U11406 ( .A(n6991), .B(n6990), .Z(n22661) );
  ANDN U11407 ( .B(n6992), .A(n22661), .Z(n6996) );
  NANDN U11408 ( .A(x[1410]), .B(y[1410]), .Z(n6994) );
  NANDN U11409 ( .A(x[1409]), .B(y[1409]), .Z(n6993) );
  AND U11410 ( .A(n6994), .B(n6993), .Z(n6995) );
  NANDN U11411 ( .A(x[1411]), .B(y[1411]), .Z(n7000) );
  AND U11412 ( .A(n6995), .B(n7000), .Z(n22662) );
  NANDN U11413 ( .A(n6996), .B(n22662), .Z(n7003) );
  XNOR U11414 ( .A(x[1411]), .B(y[1411]), .Z(n6998) );
  NANDN U11415 ( .A(y[1410]), .B(x[1410]), .Z(n6997) );
  NAND U11416 ( .A(n6998), .B(n6997), .Z(n6999) );
  NAND U11417 ( .A(n7000), .B(n6999), .Z(n7002) );
  NANDN U11418 ( .A(y[1412]), .B(x[1412]), .Z(n7001) );
  NAND U11419 ( .A(n7002), .B(n7001), .Z(n14885) );
  ANDN U11420 ( .B(n7003), .A(n14885), .Z(n7006) );
  NANDN U11421 ( .A(x[1413]), .B(y[1413]), .Z(n7005) );
  NANDN U11422 ( .A(x[1412]), .B(y[1412]), .Z(n7004) );
  AND U11423 ( .A(n7005), .B(n7004), .Z(n14889) );
  NANDN U11424 ( .A(n7006), .B(n14889), .Z(n7007) );
  NAND U11425 ( .A(n7008), .B(n7007), .Z(n7009) );
  ANDN U11426 ( .B(y[1414]), .A(x[1414]), .Z(n14890) );
  ANDN U11427 ( .B(n7009), .A(n14890), .Z(n7010) );
  NAND U11428 ( .A(n7011), .B(n7010), .Z(n7012) );
  NAND U11429 ( .A(n7013), .B(n7012), .Z(n7014) );
  ANDN U11430 ( .B(y[1416]), .A(x[1416]), .Z(n12484) );
  ANDN U11431 ( .B(n7014), .A(n12484), .Z(n7015) );
  NAND U11432 ( .A(n7016), .B(n7015), .Z(n7017) );
  NAND U11433 ( .A(n14895), .B(n7017), .Z(n7018) );
  ANDN U11434 ( .B(y[1418]), .A(x[1418]), .Z(n12482) );
  ANDN U11435 ( .B(n7018), .A(n12482), .Z(n7021) );
  NANDN U11436 ( .A(y[1418]), .B(x[1418]), .Z(n7020) );
  NANDN U11437 ( .A(y[1419]), .B(x[1419]), .Z(n7019) );
  AND U11438 ( .A(n7020), .B(n7019), .Z(n22677) );
  NANDN U11439 ( .A(n7021), .B(n22677), .Z(n7024) );
  NANDN U11440 ( .A(x[1420]), .B(y[1420]), .Z(n7023) );
  NANDN U11441 ( .A(x[1419]), .B(y[1419]), .Z(n7022) );
  AND U11442 ( .A(n7023), .B(n7022), .Z(n22678) );
  NAND U11443 ( .A(n7024), .B(n22678), .Z(n7027) );
  NANDN U11444 ( .A(y[1420]), .B(x[1420]), .Z(n7026) );
  NANDN U11445 ( .A(y[1421]), .B(x[1421]), .Z(n7025) );
  AND U11446 ( .A(n7026), .B(n7025), .Z(n22680) );
  NAND U11447 ( .A(n7027), .B(n22680), .Z(n7030) );
  NANDN U11448 ( .A(x[1421]), .B(y[1421]), .Z(n7029) );
  NANDN U11449 ( .A(x[1422]), .B(y[1422]), .Z(n7028) );
  AND U11450 ( .A(n7029), .B(n7028), .Z(n22682) );
  NAND U11451 ( .A(n7030), .B(n22682), .Z(n7033) );
  NANDN U11452 ( .A(y[1422]), .B(x[1422]), .Z(n7032) );
  NANDN U11453 ( .A(y[1423]), .B(x[1423]), .Z(n7031) );
  NAND U11454 ( .A(n7032), .B(n7031), .Z(n22685) );
  ANDN U11455 ( .B(n7033), .A(n22685), .Z(n7034) );
  OR U11456 ( .A(n22687), .B(n7034), .Z(n7035) );
  NANDN U11457 ( .A(y[1424]), .B(x[1424]), .Z(n22688) );
  NAND U11458 ( .A(n7035), .B(n22688), .Z(n7036) );
  NANDN U11459 ( .A(x[1425]), .B(y[1425]), .Z(n12479) );
  ANDN U11460 ( .B(y[1424]), .A(x[1424]), .Z(n12480) );
  ANDN U11461 ( .B(n12479), .A(n12480), .Z(n22690) );
  NAND U11462 ( .A(n7036), .B(n22690), .Z(n7037) );
  NAND U11463 ( .A(n7038), .B(n7037), .Z(n7039) );
  NANDN U11464 ( .A(x[1426]), .B(y[1426]), .Z(n22694) );
  NAND U11465 ( .A(n7039), .B(n22694), .Z(n7040) );
  NANDN U11466 ( .A(n7040), .B(x[1427]), .Z(n7043) );
  IV U11467 ( .A(y[1427]), .Z(n14910) );
  XNOR U11468 ( .A(n7040), .B(x[1427]), .Z(n7041) );
  NAND U11469 ( .A(n14910), .B(n7041), .Z(n7042) );
  NAND U11470 ( .A(n7043), .B(n7042), .Z(n7044) );
  NAND U11471 ( .A(n7045), .B(n7044), .Z(n7046) );
  NAND U11472 ( .A(n12476), .B(n7046), .Z(n7047) );
  NAND U11473 ( .A(n7048), .B(n7047), .Z(n7049) );
  NAND U11474 ( .A(n12475), .B(n7049), .Z(n7050) );
  ANDN U11475 ( .B(y[1430]), .A(x[1430]), .Z(n12474) );
  ANDN U11476 ( .B(n7050), .A(n12474), .Z(n7053) );
  NANDN U11477 ( .A(y[1430]), .B(x[1430]), .Z(n7052) );
  NANDN U11478 ( .A(y[1431]), .B(x[1431]), .Z(n7051) );
  AND U11479 ( .A(n7052), .B(n7051), .Z(n22705) );
  NANDN U11480 ( .A(n7053), .B(n22705), .Z(n7054) );
  AND U11481 ( .A(n22706), .B(n7054), .Z(n7057) );
  NANDN U11482 ( .A(y[1432]), .B(x[1432]), .Z(n7056) );
  NANDN U11483 ( .A(y[1433]), .B(x[1433]), .Z(n7055) );
  AND U11484 ( .A(n7056), .B(n7055), .Z(n22708) );
  NANDN U11485 ( .A(n7057), .B(n22708), .Z(n7062) );
  NANDN U11486 ( .A(x[1434]), .B(y[1434]), .Z(n7059) );
  NANDN U11487 ( .A(x[1433]), .B(y[1433]), .Z(n7058) );
  AND U11488 ( .A(n7059), .B(n7058), .Z(n7061) );
  NANDN U11489 ( .A(x[1435]), .B(y[1435]), .Z(n7060) );
  AND U11490 ( .A(n7061), .B(n7060), .Z(n22710) );
  NAND U11491 ( .A(n7062), .B(n22710), .Z(n7069) );
  NANDN U11492 ( .A(y[1435]), .B(x[1435]), .Z(n7064) );
  ANDN U11493 ( .B(x[1436]), .A(y[1436]), .Z(n7063) );
  ANDN U11494 ( .B(n7064), .A(n7063), .Z(n7068) );
  XNOR U11495 ( .A(x[1435]), .B(y[1435]), .Z(n7066) );
  ANDN U11496 ( .B(x[1434]), .A(y[1434]), .Z(n7065) );
  NAND U11497 ( .A(n7066), .B(n7065), .Z(n7067) );
  AND U11498 ( .A(n7068), .B(n7067), .Z(n22712) );
  NAND U11499 ( .A(n7069), .B(n22712), .Z(n7070) );
  NANDN U11500 ( .A(n22715), .B(n7070), .Z(n7071) );
  ANDN U11501 ( .B(x[1438]), .A(y[1438]), .Z(n12472) );
  ANDN U11502 ( .B(n7071), .A(n12472), .Z(n7072) );
  NANDN U11503 ( .A(y[1437]), .B(x[1437]), .Z(n22716) );
  NAND U11504 ( .A(n7072), .B(n22716), .Z(n7073) );
  NANDN U11505 ( .A(x[1438]), .B(y[1438]), .Z(n22718) );
  NAND U11506 ( .A(n7073), .B(n22718), .Z(n7074) );
  NAND U11507 ( .A(n7075), .B(n7074), .Z(n7076) );
  NAND U11508 ( .A(n14930), .B(n7076), .Z(n7077) );
  NAND U11509 ( .A(n7078), .B(n7077), .Z(n7079) );
  NAND U11510 ( .A(n7080), .B(n7079), .Z(n7081) );
  ANDN U11511 ( .B(x[1441]), .A(y[1441]), .Z(n12470) );
  ANDN U11512 ( .B(n7081), .A(n12470), .Z(n7082) );
  NAND U11513 ( .A(n7083), .B(n7082), .Z(n7084) );
  NAND U11514 ( .A(n12467), .B(n7084), .Z(n7085) );
  ANDN U11515 ( .B(x[1443]), .A(y[1443]), .Z(n12466) );
  ANDN U11516 ( .B(n7085), .A(n12466), .Z(n7088) );
  NANDN U11517 ( .A(x[1443]), .B(y[1443]), .Z(n7087) );
  NANDN U11518 ( .A(x[1444]), .B(y[1444]), .Z(n7086) );
  AND U11519 ( .A(n7087), .B(n7086), .Z(n22730) );
  NANDN U11520 ( .A(n7088), .B(n22730), .Z(n7089) );
  NANDN U11521 ( .A(n22733), .B(n7089), .Z(n7092) );
  NANDN U11522 ( .A(x[1445]), .B(y[1445]), .Z(n7091) );
  NANDN U11523 ( .A(x[1446]), .B(y[1446]), .Z(n7090) );
  AND U11524 ( .A(n7091), .B(n7090), .Z(n22734) );
  NAND U11525 ( .A(n7092), .B(n22734), .Z(n7093) );
  NANDN U11526 ( .A(n22737), .B(n7093), .Z(n7094) );
  NANDN U11527 ( .A(x[1447]), .B(y[1447]), .Z(n22738) );
  NAND U11528 ( .A(n7094), .B(n22738), .Z(n7095) );
  AND U11529 ( .A(n22741), .B(n7095), .Z(n7096) );
  OR U11530 ( .A(n22742), .B(n7096), .Z(n7097) );
  ANDN U11531 ( .B(x[1449]), .A(y[1449]), .Z(n22744) );
  ANDN U11532 ( .B(n7097), .A(n22744), .Z(n7098) );
  NANDN U11533 ( .A(n12463), .B(n7098), .Z(n7099) );
  AND U11534 ( .A(n22746), .B(n7099), .Z(n7100) );
  NAND U11535 ( .A(n7101), .B(n7100), .Z(n7102) );
  NAND U11536 ( .A(n7103), .B(n7102), .Z(n7104) );
  ANDN U11537 ( .B(y[1452]), .A(x[1452]), .Z(n12462) );
  ANDN U11538 ( .B(n7104), .A(n12462), .Z(n7105) );
  NAND U11539 ( .A(n7106), .B(n7105), .Z(n7107) );
  NAND U11540 ( .A(n12460), .B(n7107), .Z(n7108) );
  ANDN U11541 ( .B(y[1454]), .A(x[1454]), .Z(n12458) );
  ANDN U11542 ( .B(n7108), .A(n12458), .Z(n7111) );
  NANDN U11543 ( .A(y[1454]), .B(x[1454]), .Z(n7110) );
  NANDN U11544 ( .A(y[1455]), .B(x[1455]), .Z(n7109) );
  AND U11545 ( .A(n7110), .B(n7109), .Z(n22756) );
  NANDN U11546 ( .A(n7111), .B(n22756), .Z(n7114) );
  NANDN U11547 ( .A(x[1456]), .B(y[1456]), .Z(n7113) );
  NANDN U11548 ( .A(x[1455]), .B(y[1455]), .Z(n7112) );
  NAND U11549 ( .A(n7113), .B(n7112), .Z(n22759) );
  ANDN U11550 ( .B(n7114), .A(n22759), .Z(n7117) );
  NANDN U11551 ( .A(y[1456]), .B(x[1456]), .Z(n7116) );
  NANDN U11552 ( .A(y[1457]), .B(x[1457]), .Z(n7115) );
  AND U11553 ( .A(n7116), .B(n7115), .Z(n22760) );
  NANDN U11554 ( .A(n7117), .B(n22760), .Z(n7118) );
  NANDN U11555 ( .A(n14954), .B(n7118), .Z(n7121) );
  NANDN U11556 ( .A(y[1458]), .B(x[1458]), .Z(n7120) );
  AND U11557 ( .A(n7120), .B(n7119), .Z(n22764) );
  NAND U11558 ( .A(n7121), .B(n22764), .Z(n7122) );
  NANDN U11559 ( .A(n7123), .B(n7122), .Z(n7124) );
  NANDN U11560 ( .A(n12456), .B(n7124), .Z(n7125) );
  NANDN U11561 ( .A(n22770), .B(n7125), .Z(n7126) );
  NAND U11562 ( .A(n7127), .B(n7126), .Z(n7128) );
  ANDN U11563 ( .B(y[1462]), .A(x[1462]), .Z(n22775) );
  ANDN U11564 ( .B(n7128), .A(n22775), .Z(n7129) );
  OR U11565 ( .A(n14966), .B(n7129), .Z(n7132) );
  NANDN U11566 ( .A(x[1464]), .B(y[1464]), .Z(n7131) );
  NANDN U11567 ( .A(x[1463]), .B(y[1463]), .Z(n7130) );
  AND U11568 ( .A(n7131), .B(n7130), .Z(n22778) );
  NAND U11569 ( .A(n7132), .B(n22778), .Z(n7135) );
  NANDN U11570 ( .A(y[1464]), .B(x[1464]), .Z(n7134) );
  NANDN U11571 ( .A(y[1465]), .B(x[1465]), .Z(n7133) );
  AND U11572 ( .A(n7134), .B(n7133), .Z(n22781) );
  NAND U11573 ( .A(n7135), .B(n22781), .Z(n7138) );
  NANDN U11574 ( .A(x[1466]), .B(y[1466]), .Z(n7137) );
  NANDN U11575 ( .A(x[1465]), .B(y[1465]), .Z(n7136) );
  AND U11576 ( .A(n7137), .B(n7136), .Z(n22782) );
  NAND U11577 ( .A(n7138), .B(n22782), .Z(n7139) );
  NANDN U11578 ( .A(n22784), .B(n7139), .Z(n7142) );
  NANDN U11579 ( .A(x[1467]), .B(y[1467]), .Z(n7141) );
  NANDN U11580 ( .A(x[1468]), .B(y[1468]), .Z(n7140) );
  AND U11581 ( .A(n7141), .B(n7140), .Z(n22786) );
  NAND U11582 ( .A(n7142), .B(n22786), .Z(n7143) );
  NANDN U11583 ( .A(n22789), .B(n7143), .Z(n7144) );
  ANDN U11584 ( .B(y[1469]), .A(x[1469]), .Z(n14975) );
  ANDN U11585 ( .B(n7144), .A(n14975), .Z(n7146) );
  IV U11586 ( .A(x[1470]), .Z(n14974) );
  NANDN U11587 ( .A(n7146), .B(n14974), .Z(n7145) );
  AND U11588 ( .A(n22794), .B(n7145), .Z(n7149) );
  XOR U11589 ( .A(x[1470]), .B(n7146), .Z(n7147) );
  NAND U11590 ( .A(n7147), .B(y[1470]), .Z(n7148) );
  NAND U11591 ( .A(n7149), .B(n7148), .Z(n7150) );
  ANDN U11592 ( .B(x[1471]), .A(y[1471]), .Z(n12455) );
  ANDN U11593 ( .B(n7150), .A(n12455), .Z(n7151) );
  NANDN U11594 ( .A(n12453), .B(n7151), .Z(n7152) );
  NANDN U11595 ( .A(n14979), .B(n7152), .Z(n7153) );
  OR U11596 ( .A(n12451), .B(n7153), .Z(n7154) );
  NANDN U11597 ( .A(y[1473]), .B(x[1473]), .Z(n22802) );
  NAND U11598 ( .A(n7154), .B(n22802), .Z(n7156) );
  XNOR U11599 ( .A(y[1474]), .B(n7156), .Z(n7155) );
  NAND U11600 ( .A(n12450), .B(n7155), .Z(n7158) );
  NANDN U11601 ( .A(n7156), .B(y[1474]), .Z(n7157) );
  AND U11602 ( .A(n7158), .B(n7157), .Z(n7159) );
  NAND U11603 ( .A(n7160), .B(n7159), .Z(n7161) );
  NAND U11604 ( .A(n7162), .B(n7161), .Z(n7163) );
  ANDN U11605 ( .B(y[1476]), .A(x[1476]), .Z(n14986) );
  ANDN U11606 ( .B(n7163), .A(n14986), .Z(n7164) );
  NAND U11607 ( .A(n7165), .B(n7164), .Z(n7166) );
  NAND U11608 ( .A(n12446), .B(n7166), .Z(n7167) );
  ANDN U11609 ( .B(y[1478]), .A(x[1478]), .Z(n12445) );
  ANDN U11610 ( .B(n7167), .A(n12445), .Z(n7170) );
  NANDN U11611 ( .A(y[1478]), .B(x[1478]), .Z(n7169) );
  NANDN U11612 ( .A(y[1479]), .B(x[1479]), .Z(n7168) );
  AND U11613 ( .A(n7169), .B(n7168), .Z(n22813) );
  NANDN U11614 ( .A(n7170), .B(n22813), .Z(n7173) );
  NANDN U11615 ( .A(x[1480]), .B(y[1480]), .Z(n7172) );
  NANDN U11616 ( .A(x[1479]), .B(y[1479]), .Z(n7171) );
  NAND U11617 ( .A(n7172), .B(n7171), .Z(n22816) );
  ANDN U11618 ( .B(n7173), .A(n22816), .Z(n7174) );
  OR U11619 ( .A(n22818), .B(n7174), .Z(n7175) );
  ANDN U11620 ( .B(y[1481]), .A(x[1481]), .Z(n14995) );
  ANDN U11621 ( .B(n7175), .A(n14995), .Z(n7177) );
  IV U11622 ( .A(x[1482]), .Z(n14994) );
  NANDN U11623 ( .A(n7177), .B(n14994), .Z(n7176) );
  AND U11624 ( .A(n22823), .B(n7176), .Z(n7180) );
  XOR U11625 ( .A(x[1482]), .B(n7177), .Z(n7178) );
  NAND U11626 ( .A(n7178), .B(y[1482]), .Z(n7179) );
  NAND U11627 ( .A(n7180), .B(n7179), .Z(n7181) );
  ANDN U11628 ( .B(x[1483]), .A(y[1483]), .Z(n12443) );
  ANDN U11629 ( .B(n7181), .A(n12443), .Z(n7182) );
  NANDN U11630 ( .A(y[1484]), .B(x[1484]), .Z(n22825) );
  NAND U11631 ( .A(n7182), .B(n22825), .Z(n7183) );
  ANDN U11632 ( .B(y[1485]), .A(x[1485]), .Z(n15003) );
  ANDN U11633 ( .B(y[1484]), .A(x[1484]), .Z(n12441) );
  NOR U11634 ( .A(n15003), .B(n12441), .Z(n22827) );
  NAND U11635 ( .A(n7183), .B(n22827), .Z(n7184) );
  AND U11636 ( .A(n22829), .B(n7184), .Z(n7185) );
  NANDN U11637 ( .A(n12440), .B(n7185), .Z(n7186) );
  NANDN U11638 ( .A(x[1486]), .B(y[1486]), .Z(n22831) );
  NAND U11639 ( .A(n7186), .B(n22831), .Z(n7187) );
  NAND U11640 ( .A(n7188), .B(n7187), .Z(n7189) );
  AND U11641 ( .A(n12438), .B(n7189), .Z(n7190) );
  NANDN U11642 ( .A(n7190), .B(y[1488]), .Z(n7193) );
  XNOR U11643 ( .A(n7190), .B(y[1488]), .Z(n7191) );
  NANDN U11644 ( .A(x[1488]), .B(n7191), .Z(n7192) );
  NAND U11645 ( .A(n7193), .B(n7192), .Z(n7194) );
  NAND U11646 ( .A(n7195), .B(n7194), .Z(n7196) );
  NAND U11647 ( .A(n12434), .B(n7196), .Z(n7197) );
  NAND U11648 ( .A(n7198), .B(n7197), .Z(n7199) );
  NAND U11649 ( .A(n12433), .B(n7199), .Z(n7200) );
  ANDN U11650 ( .B(x[1491]), .A(y[1491]), .Z(n15011) );
  ANDN U11651 ( .B(n7200), .A(n15011), .Z(n7203) );
  NANDN U11652 ( .A(x[1491]), .B(y[1491]), .Z(n7202) );
  NANDN U11653 ( .A(x[1492]), .B(y[1492]), .Z(n7201) );
  AND U11654 ( .A(n7202), .B(n7201), .Z(n22843) );
  NANDN U11655 ( .A(n7203), .B(n22843), .Z(n7206) );
  NANDN U11656 ( .A(y[1493]), .B(x[1493]), .Z(n7205) );
  NANDN U11657 ( .A(y[1492]), .B(x[1492]), .Z(n7204) );
  NAND U11658 ( .A(n7205), .B(n7204), .Z(n22845) );
  ANDN U11659 ( .B(n7206), .A(n22845), .Z(n7209) );
  NANDN U11660 ( .A(x[1493]), .B(y[1493]), .Z(n7208) );
  NANDN U11661 ( .A(x[1494]), .B(y[1494]), .Z(n7207) );
  AND U11662 ( .A(n7208), .B(n7207), .Z(n22847) );
  NANDN U11663 ( .A(n7209), .B(n22847), .Z(n7212) );
  NANDN U11664 ( .A(y[1495]), .B(x[1495]), .Z(n7211) );
  NANDN U11665 ( .A(y[1494]), .B(x[1494]), .Z(n7210) );
  NAND U11666 ( .A(n7211), .B(n7210), .Z(n22849) );
  ANDN U11667 ( .B(n7212), .A(n22849), .Z(n7213) );
  NANDN U11668 ( .A(x[1495]), .B(y[1495]), .Z(n22852) );
  NANDN U11669 ( .A(n7213), .B(n22852), .Z(n7214) );
  NANDN U11670 ( .A(y[1496]), .B(x[1496]), .Z(n22853) );
  NAND U11671 ( .A(n7214), .B(n22853), .Z(n7215) );
  ANDN U11672 ( .B(y[1497]), .A(x[1497]), .Z(n15022) );
  ANDN U11673 ( .B(y[1496]), .A(x[1496]), .Z(n15017) );
  NOR U11674 ( .A(n15022), .B(n15017), .Z(n22855) );
  NAND U11675 ( .A(n7215), .B(n22855), .Z(n7216) );
  AND U11676 ( .A(n22857), .B(n7216), .Z(n7217) );
  NANDN U11677 ( .A(n12431), .B(n7217), .Z(n7218) );
  NANDN U11678 ( .A(n22860), .B(n7218), .Z(n7219) );
  NAND U11679 ( .A(n7220), .B(n7219), .Z(n7221) );
  NANDN U11680 ( .A(x[1499]), .B(y[1499]), .Z(n12430) );
  NAND U11681 ( .A(n7221), .B(n12430), .Z(n7223) );
  IV U11682 ( .A(y[1500]), .Z(n12426) );
  NANDN U11683 ( .A(n7223), .B(n12426), .Z(n7222) );
  ANDN U11684 ( .B(x[1501]), .A(y[1501]), .Z(n12428) );
  ANDN U11685 ( .B(n7222), .A(n12428), .Z(n7226) );
  XOR U11686 ( .A(n7223), .B(y[1500]), .Z(n7224) );
  NAND U11687 ( .A(x[1500]), .B(n7224), .Z(n7225) );
  NAND U11688 ( .A(n7226), .B(n7225), .Z(n7227) );
  AND U11689 ( .A(n22867), .B(n7227), .Z(n7230) );
  NANDN U11690 ( .A(y[1502]), .B(x[1502]), .Z(n7229) );
  NANDN U11691 ( .A(y[1503]), .B(x[1503]), .Z(n7228) );
  AND U11692 ( .A(n7229), .B(n7228), .Z(n22870) );
  NANDN U11693 ( .A(n7230), .B(n22870), .Z(n7235) );
  NANDN U11694 ( .A(x[1504]), .B(y[1504]), .Z(n7232) );
  NANDN U11695 ( .A(x[1503]), .B(y[1503]), .Z(n7231) );
  AND U11696 ( .A(n7232), .B(n7231), .Z(n7234) );
  IV U11697 ( .A(x[1505]), .Z(n7236) );
  NAND U11698 ( .A(n7236), .B(y[1505]), .Z(n7233) );
  AND U11699 ( .A(n7234), .B(n7233), .Z(n22871) );
  NAND U11700 ( .A(n7235), .B(n22871), .Z(n7241) );
  NANDN U11701 ( .A(y[1504]), .B(x[1504]), .Z(n7237) );
  NANDN U11702 ( .A(n7237), .B(x[1505]), .Z(n7240) );
  XOR U11703 ( .A(n7237), .B(n7236), .Z(n7238) );
  NANDN U11704 ( .A(y[1505]), .B(n7238), .Z(n7239) );
  AND U11705 ( .A(n7240), .B(n7239), .Z(n22873) );
  NAND U11706 ( .A(n7241), .B(n22873), .Z(n7242) );
  OR U11707 ( .A(n12425), .B(n7242), .Z(n7243) );
  ANDN U11708 ( .B(y[1507]), .A(x[1507]), .Z(n20283) );
  ANDN U11709 ( .B(y[1506]), .A(x[1506]), .Z(n15033) );
  NOR U11710 ( .A(n20283), .B(n15033), .Z(n22875) );
  NAND U11711 ( .A(n7243), .B(n22875), .Z(n7244) );
  NANDN U11712 ( .A(n20284), .B(n7244), .Z(n7245) );
  OR U11713 ( .A(n12424), .B(n7245), .Z(n7246) );
  NANDN U11714 ( .A(n22880), .B(n7246), .Z(n7247) );
  ANDN U11715 ( .B(x[1510]), .A(y[1510]), .Z(n15044) );
  ANDN U11716 ( .B(n7247), .A(n15044), .Z(n7248) );
  IV U11717 ( .A(y[1511]), .Z(n15042) );
  NANDN U11718 ( .A(n7248), .B(n15042), .Z(n7251) );
  XOR U11719 ( .A(y[1511]), .B(n7248), .Z(n7249) );
  NAND U11720 ( .A(n7249), .B(x[1511]), .Z(n7250) );
  NAND U11721 ( .A(n7251), .B(n7250), .Z(n7252) );
  ANDN U11722 ( .B(y[1512]), .A(x[1512]), .Z(n12423) );
  ANDN U11723 ( .B(n7252), .A(n12423), .Z(n7255) );
  NANDN U11724 ( .A(y[1512]), .B(x[1512]), .Z(n7254) );
  NANDN U11725 ( .A(y[1513]), .B(x[1513]), .Z(n7253) );
  AND U11726 ( .A(n7254), .B(n7253), .Z(n22886) );
  NANDN U11727 ( .A(n7255), .B(n22886), .Z(n7256) );
  AND U11728 ( .A(n22887), .B(n7256), .Z(n7259) );
  NANDN U11729 ( .A(y[1514]), .B(x[1514]), .Z(n7258) );
  NANDN U11730 ( .A(y[1515]), .B(x[1515]), .Z(n7257) );
  AND U11731 ( .A(n7258), .B(n7257), .Z(n22890) );
  NANDN U11732 ( .A(n7259), .B(n22890), .Z(n7262) );
  NANDN U11733 ( .A(x[1516]), .B(y[1516]), .Z(n7261) );
  NANDN U11734 ( .A(x[1515]), .B(y[1515]), .Z(n7260) );
  AND U11735 ( .A(n7261), .B(n7260), .Z(n22891) );
  NAND U11736 ( .A(n7262), .B(n22891), .Z(n7265) );
  NANDN U11737 ( .A(y[1516]), .B(x[1516]), .Z(n7264) );
  NANDN U11738 ( .A(y[1517]), .B(x[1517]), .Z(n7263) );
  AND U11739 ( .A(n7264), .B(n7263), .Z(n22894) );
  NAND U11740 ( .A(n7265), .B(n22894), .Z(n7266) );
  ANDN U11741 ( .B(y[1517]), .A(x[1517]), .Z(n12421) );
  ANDN U11742 ( .B(n7266), .A(n12421), .Z(n7268) );
  XNOR U11743 ( .A(y[1518]), .B(x[1518]), .Z(n7267) );
  NANDN U11744 ( .A(n7268), .B(n7267), .Z(n7269) );
  NAND U11745 ( .A(n7270), .B(n7269), .Z(n7271) );
  ANDN U11746 ( .B(x[1519]), .A(y[1519]), .Z(n15054) );
  ANDN U11747 ( .B(n7271), .A(n15054), .Z(n7272) );
  NANDN U11748 ( .A(n22902), .B(n7272), .Z(n7277) );
  ANDN U11749 ( .B(y[1520]), .A(x[1520]), .Z(n15056) );
  NANDN U11750 ( .A(n7273), .B(n15056), .Z(n7276) );
  NANDN U11751 ( .A(x[1522]), .B(y[1522]), .Z(n7275) );
  NANDN U11752 ( .A(x[1521]), .B(y[1521]), .Z(n7274) );
  AND U11753 ( .A(n7275), .B(n7274), .Z(n15060) );
  NAND U11754 ( .A(n7276), .B(n15060), .Z(n22904) );
  ANDN U11755 ( .B(n7277), .A(n22904), .Z(n7280) );
  NANDN U11756 ( .A(y[1522]), .B(x[1522]), .Z(n7279) );
  NANDN U11757 ( .A(y[1523]), .B(x[1523]), .Z(n7278) );
  AND U11758 ( .A(n7279), .B(n7278), .Z(n22906) );
  NANDN U11759 ( .A(n7280), .B(n22906), .Z(n7283) );
  NANDN U11760 ( .A(x[1524]), .B(y[1524]), .Z(n7282) );
  NANDN U11761 ( .A(x[1523]), .B(y[1523]), .Z(n7281) );
  AND U11762 ( .A(n7282), .B(n7281), .Z(n22907) );
  NAND U11763 ( .A(n7283), .B(n22907), .Z(n7286) );
  NANDN U11764 ( .A(y[1524]), .B(x[1524]), .Z(n7285) );
  NANDN U11765 ( .A(y[1525]), .B(x[1525]), .Z(n7284) );
  AND U11766 ( .A(n7285), .B(n7284), .Z(n22910) );
  NAND U11767 ( .A(n7286), .B(n22910), .Z(n7289) );
  NANDN U11768 ( .A(x[1526]), .B(y[1526]), .Z(n7288) );
  NANDN U11769 ( .A(x[1525]), .B(y[1525]), .Z(n7287) );
  AND U11770 ( .A(n7288), .B(n7287), .Z(n22911) );
  NAND U11771 ( .A(n7289), .B(n22911), .Z(n7292) );
  NANDN U11772 ( .A(y[1526]), .B(x[1526]), .Z(n7291) );
  NANDN U11773 ( .A(y[1527]), .B(x[1527]), .Z(n7290) );
  AND U11774 ( .A(n7291), .B(n7290), .Z(n22914) );
  NAND U11775 ( .A(n7292), .B(n22914), .Z(n7293) );
  AND U11776 ( .A(n22915), .B(n7293), .Z(n7296) );
  NANDN U11777 ( .A(y[1528]), .B(x[1528]), .Z(n7295) );
  NANDN U11778 ( .A(y[1529]), .B(x[1529]), .Z(n7294) );
  AND U11779 ( .A(n7295), .B(n7294), .Z(n22917) );
  NANDN U11780 ( .A(n7296), .B(n22917), .Z(n7297) );
  ANDN U11781 ( .B(y[1529]), .A(x[1529]), .Z(n15069) );
  ANDN U11782 ( .B(n7297), .A(n15069), .Z(n7298) );
  NAND U11783 ( .A(n7299), .B(n7298), .Z(n7300) );
  NAND U11784 ( .A(n12418), .B(n7300), .Z(n7301) );
  NANDN U11785 ( .A(x[1531]), .B(y[1531]), .Z(n22923) );
  NAND U11786 ( .A(n7301), .B(n22923), .Z(n7302) );
  ANDN U11787 ( .B(x[1532]), .A(y[1532]), .Z(n22926) );
  ANDN U11788 ( .B(n7302), .A(n22926), .Z(n7303) );
  NANDN U11789 ( .A(n12419), .B(n7303), .Z(n7304) );
  NANDN U11790 ( .A(x[1533]), .B(y[1533]), .Z(n15078) );
  ANDN U11791 ( .B(y[1532]), .A(x[1532]), .Z(n12417) );
  ANDN U11792 ( .B(n15078), .A(n12417), .Z(n22927) );
  NAND U11793 ( .A(n7304), .B(n22927), .Z(n7305) );
  ANDN U11794 ( .B(x[1534]), .A(y[1534]), .Z(n12412) );
  ANDN U11795 ( .B(n7305), .A(n12412), .Z(n7306) );
  NANDN U11796 ( .A(y[1533]), .B(x[1533]), .Z(n22930) );
  NAND U11797 ( .A(n7306), .B(n22930), .Z(n7309) );
  NANDN U11798 ( .A(x[1534]), .B(y[1534]), .Z(n7308) );
  NANDN U11799 ( .A(x[1536]), .B(y[1536]), .Z(n7313) );
  NANDN U11800 ( .A(x[1535]), .B(y[1535]), .Z(n7307) );
  NAND U11801 ( .A(n7313), .B(n7307), .Z(n12414) );
  ANDN U11802 ( .B(n7308), .A(n12414), .Z(n22932) );
  NAND U11803 ( .A(n7309), .B(n22932), .Z(n7312) );
  NANDN U11804 ( .A(y[1537]), .B(x[1537]), .Z(n7311) );
  NANDN U11805 ( .A(y[1536]), .B(x[1536]), .Z(n7310) );
  NAND U11806 ( .A(n7311), .B(n7310), .Z(n12415) );
  ANDN U11807 ( .B(n7312), .A(n12415), .Z(n7315) );
  ANDN U11808 ( .B(x[1535]), .A(y[1535]), .Z(n12411) );
  NAND U11809 ( .A(n7313), .B(n12411), .Z(n7314) );
  AND U11810 ( .A(n7315), .B(n7314), .Z(n7318) );
  NANDN U11811 ( .A(x[1537]), .B(y[1537]), .Z(n7317) );
  NANDN U11812 ( .A(x[1538]), .B(y[1538]), .Z(n7316) );
  AND U11813 ( .A(n7317), .B(n7316), .Z(n22936) );
  NANDN U11814 ( .A(n7318), .B(n22936), .Z(n7319) );
  AND U11815 ( .A(n22937), .B(n7319), .Z(n7322) );
  NANDN U11816 ( .A(x[1539]), .B(y[1539]), .Z(n7321) );
  NANDN U11817 ( .A(x[1540]), .B(y[1540]), .Z(n7320) );
  AND U11818 ( .A(n7321), .B(n7320), .Z(n22939) );
  NANDN U11819 ( .A(n7322), .B(n22939), .Z(n7323) );
  AND U11820 ( .A(n22941), .B(n7323), .Z(n7324) );
  OR U11821 ( .A(n12409), .B(n7324), .Z(n7325) );
  NANDN U11822 ( .A(n15086), .B(n7325), .Z(n7326) );
  NANDN U11823 ( .A(n22947), .B(n7326), .Z(n7327) );
  OR U11824 ( .A(n12410), .B(n7327), .Z(n7328) );
  ANDN U11825 ( .B(x[1543]), .A(y[1543]), .Z(n15087) );
  ANDN U11826 ( .B(n7328), .A(n15087), .Z(n7329) );
  NANDN U11827 ( .A(n15091), .B(n7329), .Z(n7330) );
  ANDN U11828 ( .B(y[1545]), .A(x[1545]), .Z(n12407) );
  ANDN U11829 ( .B(n7330), .A(n12407), .Z(n7331) );
  NANDN U11830 ( .A(n12408), .B(n7331), .Z(n7332) );
  NANDN U11831 ( .A(y[1545]), .B(x[1545]), .Z(n20281) );
  NAND U11832 ( .A(n7332), .B(n20281), .Z(n7333) );
  NAND U11833 ( .A(n7334), .B(n7333), .Z(n7335) );
  NAND U11834 ( .A(n15096), .B(n7335), .Z(n7336) );
  NAND U11835 ( .A(n7337), .B(n7336), .Z(n7338) );
  NAND U11836 ( .A(n15095), .B(n7338), .Z(n7339) );
  ANDN U11837 ( .B(y[1548]), .A(x[1548]), .Z(n12405) );
  ANDN U11838 ( .B(n7339), .A(n12405), .Z(n7342) );
  NANDN U11839 ( .A(y[1548]), .B(x[1548]), .Z(n7341) );
  NANDN U11840 ( .A(y[1549]), .B(x[1549]), .Z(n7340) );
  AND U11841 ( .A(n7341), .B(n7340), .Z(n22959) );
  NANDN U11842 ( .A(n7342), .B(n22959), .Z(n7345) );
  NANDN U11843 ( .A(x[1550]), .B(y[1550]), .Z(n7344) );
  NANDN U11844 ( .A(x[1549]), .B(y[1549]), .Z(n7343) );
  NAND U11845 ( .A(n7344), .B(n7343), .Z(n22961) );
  ANDN U11846 ( .B(n7345), .A(n22961), .Z(n7348) );
  NANDN U11847 ( .A(y[1550]), .B(x[1550]), .Z(n7347) );
  NANDN U11848 ( .A(y[1551]), .B(x[1551]), .Z(n7346) );
  AND U11849 ( .A(n7347), .B(n7346), .Z(n22963) );
  NANDN U11850 ( .A(n7348), .B(n22963), .Z(n7349) );
  AND U11851 ( .A(n22965), .B(n7349), .Z(n7352) );
  NANDN U11852 ( .A(y[1553]), .B(x[1553]), .Z(n7351) );
  NANDN U11853 ( .A(y[1552]), .B(x[1552]), .Z(n7350) );
  AND U11854 ( .A(n7351), .B(n7350), .Z(n22967) );
  NANDN U11855 ( .A(n7352), .B(n22967), .Z(n7353) );
  ANDN U11856 ( .B(y[1553]), .A(x[1553]), .Z(n15105) );
  ANDN U11857 ( .B(n7353), .A(n15105), .Z(n7355) );
  IV U11858 ( .A(x[1554]), .Z(n15104) );
  NANDN U11859 ( .A(n7355), .B(n15104), .Z(n7354) );
  ANDN U11860 ( .B(y[1555]), .A(x[1555]), .Z(n22974) );
  ANDN U11861 ( .B(n7354), .A(n22974), .Z(n7358) );
  XOR U11862 ( .A(x[1554]), .B(n7355), .Z(n7356) );
  NAND U11863 ( .A(n7356), .B(y[1554]), .Z(n7357) );
  NAND U11864 ( .A(n7358), .B(n7357), .Z(n7359) );
  ANDN U11865 ( .B(x[1555]), .A(y[1555]), .Z(n12403) );
  ANDN U11866 ( .B(n7359), .A(n12403), .Z(n7360) );
  NANDN U11867 ( .A(n22976), .B(n7360), .Z(n7361) );
  NANDN U11868 ( .A(x[1556]), .B(y[1556]), .Z(n22977) );
  NAND U11869 ( .A(n7361), .B(n22977), .Z(n7362) );
  OR U11870 ( .A(n12400), .B(n7362), .Z(n7363) );
  NANDN U11871 ( .A(y[1557]), .B(x[1557]), .Z(n22980) );
  NAND U11872 ( .A(n7363), .B(n22980), .Z(n7364) );
  NANDN U11873 ( .A(n7364), .B(y[1558]), .Z(n7367) );
  IV U11874 ( .A(x[1558]), .Z(n12399) );
  XNOR U11875 ( .A(n7364), .B(y[1558]), .Z(n7365) );
  NAND U11876 ( .A(n12399), .B(n7365), .Z(n7366) );
  NAND U11877 ( .A(n7367), .B(n7366), .Z(n7368) );
  NAND U11878 ( .A(n7369), .B(n7368), .Z(n7370) );
  NAND U11879 ( .A(n15116), .B(n7370), .Z(n7371) );
  NAND U11880 ( .A(n7372), .B(n7371), .Z(n7373) );
  NAND U11881 ( .A(n15115), .B(n7373), .Z(n7374) );
  ANDN U11882 ( .B(x[1561]), .A(y[1561]), .Z(n12396) );
  ANDN U11883 ( .B(n7374), .A(n12396), .Z(n7377) );
  NANDN U11884 ( .A(x[1561]), .B(y[1561]), .Z(n7376) );
  NANDN U11885 ( .A(x[1562]), .B(y[1562]), .Z(n7375) );
  AND U11886 ( .A(n7376), .B(n7375), .Z(n22989) );
  NANDN U11887 ( .A(n7377), .B(n22989), .Z(n7378) );
  NANDN U11888 ( .A(x[1563]), .B(y[1563]), .Z(n7380) );
  NANDN U11889 ( .A(x[1564]), .B(y[1564]), .Z(n7379) );
  AND U11890 ( .A(n7380), .B(n7379), .Z(n22993) );
  NANDN U11891 ( .A(y[1566]), .B(x[1566]), .Z(n7381) );
  ANDN U11892 ( .B(x[1567]), .A(y[1567]), .Z(n7382) );
  ANDN U11893 ( .B(n7381), .A(n7382), .Z(n22999) );
  NANDN U11894 ( .A(x[1567]), .B(y[1567]), .Z(n23001) );
  NANDN U11895 ( .A(x[1566]), .B(y[1566]), .Z(n12393) );
  NANDN U11896 ( .A(y[1568]), .B(x[1568]), .Z(n23003) );
  NANDN U11897 ( .A(x[1569]), .B(y[1569]), .Z(n15130) );
  NANDN U11898 ( .A(x[1568]), .B(y[1568]), .Z(n12392) );
  NAND U11899 ( .A(n15130), .B(n12392), .Z(n23006) );
  NANDN U11900 ( .A(x[1570]), .B(y[1570]), .Z(n7385) );
  NANDN U11901 ( .A(x[1571]), .B(y[1571]), .Z(n7383) );
  NANDN U11902 ( .A(n7384), .B(n7383), .Z(n12389) );
  ANDN U11903 ( .B(n7385), .A(n12389), .Z(n23010) );
  NANDN U11904 ( .A(y[1573]), .B(x[1573]), .Z(n7387) );
  NANDN U11905 ( .A(y[1572]), .B(x[1572]), .Z(n7386) );
  NAND U11906 ( .A(n7387), .B(n7386), .Z(n12390) );
  NANDN U11907 ( .A(x[1573]), .B(y[1573]), .Z(n7389) );
  NANDN U11908 ( .A(x[1574]), .B(y[1574]), .Z(n7388) );
  AND U11909 ( .A(n7389), .B(n7388), .Z(n23014) );
  NANDN U11910 ( .A(y[1575]), .B(x[1575]), .Z(n7391) );
  NANDN U11911 ( .A(y[1574]), .B(x[1574]), .Z(n7390) );
  AND U11912 ( .A(n7391), .B(n7390), .Z(n23015) );
  NANDN U11913 ( .A(x[1575]), .B(y[1575]), .Z(n7393) );
  NANDN U11914 ( .A(x[1576]), .B(y[1576]), .Z(n7392) );
  AND U11915 ( .A(n7393), .B(n7392), .Z(n23018) );
  AND U11916 ( .A(n23019), .B(n7394), .Z(n7397) );
  NANDN U11917 ( .A(x[1577]), .B(y[1577]), .Z(n7396) );
  NANDN U11918 ( .A(x[1578]), .B(y[1578]), .Z(n7395) );
  AND U11919 ( .A(n7396), .B(n7395), .Z(n23022) );
  NANDN U11920 ( .A(n7397), .B(n23022), .Z(n7398) );
  ANDN U11921 ( .B(x[1578]), .A(y[1578]), .Z(n15139) );
  ANDN U11922 ( .B(n7398), .A(n15139), .Z(n7399) );
  OR U11923 ( .A(n23025), .B(n7399), .Z(n7400) );
  NAND U11924 ( .A(n7401), .B(n7400), .Z(n7402) );
  AND U11925 ( .A(n23029), .B(n7402), .Z(n7403) );
  NAND U11926 ( .A(n7404), .B(n7403), .Z(n7405) );
  NAND U11927 ( .A(n12380), .B(n7405), .Z(n7406) );
  ANDN U11928 ( .B(y[1584]), .A(x[1584]), .Z(n15146) );
  ANDN U11929 ( .B(n7406), .A(n15146), .Z(n7409) );
  NANDN U11930 ( .A(y[1584]), .B(x[1584]), .Z(n7408) );
  NANDN U11931 ( .A(y[1585]), .B(x[1585]), .Z(n7407) );
  AND U11932 ( .A(n7408), .B(n7407), .Z(n23035) );
  NANDN U11933 ( .A(n7409), .B(n23035), .Z(n7412) );
  NANDN U11934 ( .A(x[1586]), .B(y[1586]), .Z(n7411) );
  NANDN U11935 ( .A(x[1585]), .B(y[1585]), .Z(n7410) );
  NAND U11936 ( .A(n7411), .B(n7410), .Z(n23037) );
  ANDN U11937 ( .B(n7412), .A(n23037), .Z(n7415) );
  NANDN U11938 ( .A(y[1586]), .B(x[1586]), .Z(n7414) );
  NANDN U11939 ( .A(y[1587]), .B(x[1587]), .Z(n7413) );
  AND U11940 ( .A(n7414), .B(n7413), .Z(n23039) );
  NANDN U11941 ( .A(n7415), .B(n23039), .Z(n7416) );
  NANDN U11942 ( .A(n23042), .B(n7416), .Z(n7419) );
  NANDN U11943 ( .A(y[1588]), .B(x[1588]), .Z(n7418) );
  NANDN U11944 ( .A(y[1589]), .B(x[1589]), .Z(n7417) );
  AND U11945 ( .A(n7418), .B(n7417), .Z(n23043) );
  NAND U11946 ( .A(n7419), .B(n23043), .Z(n7420) );
  NANDN U11947 ( .A(n15154), .B(n7420), .Z(n7421) );
  AND U11948 ( .A(n23047), .B(n7421), .Z(n7425) );
  NANDN U11949 ( .A(x[1591]), .B(y[1591]), .Z(n23049) );
  NANDN U11950 ( .A(x[1590]), .B(y[1590]), .Z(n15153) );
  NAND U11951 ( .A(n23049), .B(n15153), .Z(n7423) );
  ANDN U11952 ( .B(n7423), .A(n7422), .Z(n7424) );
  OR U11953 ( .A(n7425), .B(n7424), .Z(n7426) );
  NANDN U11954 ( .A(y[1592]), .B(x[1592]), .Z(n23051) );
  NAND U11955 ( .A(n7426), .B(n23051), .Z(n7427) );
  ANDN U11956 ( .B(y[1593]), .A(x[1593]), .Z(n12379) );
  ANDN U11957 ( .B(y[1592]), .A(x[1592]), .Z(n15157) );
  NOR U11958 ( .A(n12379), .B(n15157), .Z(n23053) );
  NAND U11959 ( .A(n7427), .B(n23053), .Z(n7428) );
  ANDN U11960 ( .B(x[1593]), .A(y[1593]), .Z(n23055) );
  ANDN U11961 ( .B(n7428), .A(n23055), .Z(n7429) );
  NANDN U11962 ( .A(n12378), .B(n7429), .Z(n7430) );
  NANDN U11963 ( .A(x[1594]), .B(y[1594]), .Z(n23057) );
  NAND U11964 ( .A(n7430), .B(n23057), .Z(n7431) );
  NAND U11965 ( .A(n7432), .B(n7431), .Z(n7433) );
  NANDN U11966 ( .A(x[1595]), .B(y[1595]), .Z(n12376) );
  NAND U11967 ( .A(n7433), .B(n12376), .Z(n7435) );
  IV U11968 ( .A(y[1596]), .Z(n15166) );
  NANDN U11969 ( .A(n7435), .B(n15166), .Z(n7434) );
  ANDN U11970 ( .B(x[1597]), .A(y[1597]), .Z(n15168) );
  ANDN U11971 ( .B(n7434), .A(n15168), .Z(n7438) );
  XOR U11972 ( .A(n7435), .B(y[1596]), .Z(n7436) );
  NAND U11973 ( .A(n7436), .B(x[1596]), .Z(n7437) );
  NAND U11974 ( .A(n7438), .B(n7437), .Z(n7441) );
  NANDN U11975 ( .A(x[1598]), .B(y[1598]), .Z(n7440) );
  NANDN U11976 ( .A(x[1597]), .B(y[1597]), .Z(n7439) );
  AND U11977 ( .A(n7440), .B(n7439), .Z(n23065) );
  NAND U11978 ( .A(n7441), .B(n23065), .Z(n7444) );
  NANDN U11979 ( .A(y[1598]), .B(x[1598]), .Z(n7443) );
  NANDN U11980 ( .A(y[1599]), .B(x[1599]), .Z(n7442) );
  AND U11981 ( .A(n7443), .B(n7442), .Z(n23067) );
  NAND U11982 ( .A(n7444), .B(n23067), .Z(n7445) );
  AND U11983 ( .A(n23069), .B(n7445), .Z(n7448) );
  NANDN U11984 ( .A(y[1600]), .B(x[1600]), .Z(n7447) );
  NANDN U11985 ( .A(y[1601]), .B(x[1601]), .Z(n7446) );
  AND U11986 ( .A(n7447), .B(n7446), .Z(n23071) );
  NANDN U11987 ( .A(n7448), .B(n23071), .Z(n7453) );
  NANDN U11988 ( .A(x[1602]), .B(y[1602]), .Z(n7450) );
  NANDN U11989 ( .A(x[1601]), .B(y[1601]), .Z(n7449) );
  AND U11990 ( .A(n7450), .B(n7449), .Z(n7452) );
  NANDN U11991 ( .A(x[1603]), .B(y[1603]), .Z(n7451) );
  AND U11992 ( .A(n7452), .B(n7451), .Z(n23073) );
  NAND U11993 ( .A(n7453), .B(n23073), .Z(n7460) );
  NANDN U11994 ( .A(y[1603]), .B(x[1603]), .Z(n7455) );
  ANDN U11995 ( .B(x[1604]), .A(y[1604]), .Z(n7454) );
  ANDN U11996 ( .B(n7455), .A(n7454), .Z(n7459) );
  XNOR U11997 ( .A(x[1603]), .B(y[1603]), .Z(n7457) );
  ANDN U11998 ( .B(x[1602]), .A(y[1602]), .Z(n7456) );
  NAND U11999 ( .A(n7457), .B(n7456), .Z(n7458) );
  AND U12000 ( .A(n7459), .B(n7458), .Z(n23076) );
  NAND U12001 ( .A(n7460), .B(n23076), .Z(n7463) );
  NANDN U12002 ( .A(x[1604]), .B(y[1604]), .Z(n7462) );
  NANDN U12003 ( .A(x[1605]), .B(y[1605]), .Z(n7461) );
  AND U12004 ( .A(n7462), .B(n7461), .Z(n23077) );
  NAND U12005 ( .A(n7463), .B(n23077), .Z(n7464) );
  ANDN U12006 ( .B(x[1606]), .A(y[1606]), .Z(n12374) );
  ANDN U12007 ( .B(n7464), .A(n12374), .Z(n7465) );
  NANDN U12008 ( .A(y[1605]), .B(x[1605]), .Z(n23079) );
  NAND U12009 ( .A(n7465), .B(n23079), .Z(n7466) );
  NANDN U12010 ( .A(x[1606]), .B(y[1606]), .Z(n23081) );
  NAND U12011 ( .A(n7466), .B(n23081), .Z(n7467) );
  NAND U12012 ( .A(n7468), .B(n7467), .Z(n7469) );
  NAND U12013 ( .A(n15180), .B(n7469), .Z(n7470) );
  NAND U12014 ( .A(n7471), .B(n7470), .Z(n7472) );
  NAND U12015 ( .A(n15181), .B(n7472), .Z(n7473) );
  ANDN U12016 ( .B(x[1609]), .A(y[1609]), .Z(n12372) );
  ANDN U12017 ( .B(n7473), .A(n12372), .Z(n7474) );
  NANDN U12018 ( .A(x[1609]), .B(y[1609]), .Z(n23089) );
  NANDN U12019 ( .A(n7474), .B(n23089), .Z(n7475) );
  NANDN U12020 ( .A(y[1610]), .B(x[1610]), .Z(n23091) );
  NAND U12021 ( .A(n7475), .B(n23091), .Z(n7477) );
  NANDN U12022 ( .A(x[1611]), .B(y[1611]), .Z(n7476) );
  ANDN U12023 ( .B(y[1610]), .A(x[1610]), .Z(n12370) );
  ANDN U12024 ( .B(n7476), .A(n12370), .Z(n23093) );
  NAND U12025 ( .A(n7477), .B(n23093), .Z(n7478) );
  NANDN U12026 ( .A(n23096), .B(n7478), .Z(n7480) );
  IV U12027 ( .A(x[1612]), .Z(n15193) );
  NAND U12028 ( .A(n15193), .B(y[1612]), .Z(n7479) );
  NANDN U12029 ( .A(x[1613]), .B(y[1613]), .Z(n15198) );
  NAND U12030 ( .A(n7479), .B(n15198), .Z(n23097) );
  ANDN U12031 ( .B(n7480), .A(n23097), .Z(n7482) );
  NANDN U12032 ( .A(y[1613]), .B(x[1613]), .Z(n23099) );
  ANDN U12033 ( .B(x[1614]), .A(y[1614]), .Z(n12368) );
  ANDN U12034 ( .B(n23099), .A(n12368), .Z(n7481) );
  NANDN U12035 ( .A(n7482), .B(n7481), .Z(n7483) );
  AND U12036 ( .A(n23101), .B(n7483), .Z(n7484) );
  OR U12037 ( .A(n12369), .B(n7484), .Z(n7487) );
  NANDN U12038 ( .A(x[1616]), .B(y[1616]), .Z(n7486) );
  NANDN U12039 ( .A(x[1615]), .B(y[1615]), .Z(n7485) );
  NAND U12040 ( .A(n7486), .B(n7485), .Z(n23106) );
  ANDN U12041 ( .B(n7487), .A(n23106), .Z(n7490) );
  NANDN U12042 ( .A(y[1616]), .B(x[1616]), .Z(n7489) );
  NANDN U12043 ( .A(y[1617]), .B(x[1617]), .Z(n7488) );
  AND U12044 ( .A(n7489), .B(n7488), .Z(n23107) );
  NANDN U12045 ( .A(n7490), .B(n23107), .Z(n7493) );
  NANDN U12046 ( .A(x[1618]), .B(y[1618]), .Z(n7492) );
  NANDN U12047 ( .A(x[1617]), .B(y[1617]), .Z(n7491) );
  NAND U12048 ( .A(n7492), .B(n7491), .Z(n23109) );
  ANDN U12049 ( .B(n7493), .A(n23109), .Z(n7496) );
  NANDN U12050 ( .A(y[1618]), .B(x[1618]), .Z(n7495) );
  NANDN U12051 ( .A(y[1619]), .B(x[1619]), .Z(n7494) );
  AND U12052 ( .A(n7495), .B(n7494), .Z(n23111) );
  NANDN U12053 ( .A(n7496), .B(n23111), .Z(n7497) );
  NANDN U12054 ( .A(n23114), .B(n7497), .Z(n7498) );
  NANDN U12055 ( .A(n12366), .B(n7498), .Z(n7499) );
  NAND U12056 ( .A(n7500), .B(n7499), .Z(n7501) );
  NAND U12057 ( .A(n12367), .B(n7501), .Z(n7502) );
  NAND U12058 ( .A(n7503), .B(n7502), .Z(n7504) );
  NANDN U12059 ( .A(y[1622]), .B(x[1622]), .Z(n15210) );
  AND U12060 ( .A(n7504), .B(n15210), .Z(n7505) );
  NANDN U12061 ( .A(n15209), .B(n7505), .Z(n7507) );
  NANDN U12062 ( .A(x[1624]), .B(y[1624]), .Z(n7506) );
  ANDN U12063 ( .B(y[1623]), .A(x[1623]), .Z(n23122) );
  ANDN U12064 ( .B(n7506), .A(n23122), .Z(n15212) );
  NAND U12065 ( .A(n7507), .B(n15212), .Z(n7508) );
  AND U12066 ( .A(n15214), .B(n7508), .Z(n7510) );
  NANDN U12067 ( .A(x[1625]), .B(y[1625]), .Z(n7509) );
  ANDN U12068 ( .B(y[1626]), .A(x[1626]), .Z(n23135) );
  ANDN U12069 ( .B(n7509), .A(n23135), .Z(n15217) );
  NANDN U12070 ( .A(n7510), .B(n15217), .Z(n7511) );
  AND U12071 ( .A(n20279), .B(n7511), .Z(n7512) );
  XNOR U12072 ( .A(y[1627]), .B(x[1627]), .Z(n23133) );
  NANDN U12073 ( .A(n7512), .B(n23133), .Z(n7513) );
  AND U12074 ( .A(n7514), .B(n7513), .Z(n7515) );
  NANDN U12075 ( .A(x[1628]), .B(y[1628]), .Z(n23138) );
  NANDN U12076 ( .A(n7515), .B(n23138), .Z(n7516) );
  NANDN U12077 ( .A(n12363), .B(n7516), .Z(n7519) );
  NANDN U12078 ( .A(x[1629]), .B(y[1629]), .Z(n7518) );
  NANDN U12079 ( .A(x[1630]), .B(y[1630]), .Z(n7517) );
  AND U12080 ( .A(n7518), .B(n7517), .Z(n23143) );
  NAND U12081 ( .A(n7519), .B(n23143), .Z(n7522) );
  NANDN U12082 ( .A(y[1631]), .B(x[1631]), .Z(n7521) );
  NANDN U12083 ( .A(y[1630]), .B(x[1630]), .Z(n7520) );
  AND U12084 ( .A(n7521), .B(n7520), .Z(n23144) );
  NAND U12085 ( .A(n7522), .B(n23144), .Z(n7523) );
  AND U12086 ( .A(n23146), .B(n7523), .Z(n7526) );
  NANDN U12087 ( .A(y[1632]), .B(x[1632]), .Z(n7525) );
  AND U12088 ( .A(n7525), .B(n7524), .Z(n23148) );
  NANDN U12089 ( .A(n7526), .B(n23148), .Z(n7527) );
  NANDN U12090 ( .A(n23151), .B(n7527), .Z(n7528) );
  AND U12091 ( .A(n23154), .B(n7528), .Z(n7529) );
  NANDN U12092 ( .A(x[1636]), .B(y[1636]), .Z(n20277) );
  NANDN U12093 ( .A(n7529), .B(n20277), .Z(n7530) );
  AND U12094 ( .A(n15232), .B(n7530), .Z(n7531) );
  NANDN U12095 ( .A(x[1637]), .B(y[1637]), .Z(n20276) );
  NANDN U12096 ( .A(n7531), .B(n20276), .Z(n7532) );
  NANDN U12097 ( .A(n23158), .B(n7532), .Z(n7534) );
  NANDN U12098 ( .A(x[1639]), .B(y[1639]), .Z(n7533) );
  ANDN U12099 ( .B(y[1638]), .A(x[1638]), .Z(n12360) );
  ANDN U12100 ( .B(n7533), .A(n12360), .Z(n23162) );
  NAND U12101 ( .A(n7534), .B(n23162), .Z(n7535) );
  NANDN U12102 ( .A(n23164), .B(n7535), .Z(n7536) );
  ANDN U12103 ( .B(y[1641]), .A(x[1641]), .Z(n12356) );
  ANDN U12104 ( .B(n7536), .A(n12356), .Z(n7537) );
  NANDN U12105 ( .A(x[1640]), .B(y[1640]), .Z(n23166) );
  NAND U12106 ( .A(n7537), .B(n23166), .Z(n7539) );
  NANDN U12107 ( .A(y[1641]), .B(x[1641]), .Z(n7538) );
  ANDN U12108 ( .B(x[1642]), .A(y[1642]), .Z(n12357) );
  ANDN U12109 ( .B(n7538), .A(n12357), .Z(n23169) );
  NAND U12110 ( .A(n7539), .B(n23169), .Z(n7540) );
  NANDN U12111 ( .A(n12359), .B(n7540), .Z(n7543) );
  NANDN U12112 ( .A(y[1644]), .B(x[1644]), .Z(n7542) );
  NANDN U12113 ( .A(y[1643]), .B(x[1643]), .Z(n7541) );
  NAND U12114 ( .A(n7542), .B(n7541), .Z(n23173) );
  ANDN U12115 ( .B(n7543), .A(n23173), .Z(n7546) );
  NANDN U12116 ( .A(x[1644]), .B(y[1644]), .Z(n7545) );
  NANDN U12117 ( .A(x[1645]), .B(y[1645]), .Z(n7544) );
  AND U12118 ( .A(n7545), .B(n7544), .Z(n23174) );
  NANDN U12119 ( .A(n7546), .B(n23174), .Z(n7548) );
  NANDN U12120 ( .A(y[1646]), .B(x[1646]), .Z(n7547) );
  ANDN U12121 ( .B(x[1645]), .A(y[1645]), .Z(n15250) );
  ANDN U12122 ( .B(n7547), .A(n15250), .Z(n23176) );
  NAND U12123 ( .A(n7548), .B(n23176), .Z(n7550) );
  NANDN U12124 ( .A(x[1646]), .B(y[1646]), .Z(n7549) );
  ANDN U12125 ( .B(y[1647]), .A(x[1647]), .Z(n15256) );
  ANDN U12126 ( .B(n7549), .A(n15256), .Z(n23179) );
  NAND U12127 ( .A(n7550), .B(n23179), .Z(n7551) );
  NAND U12128 ( .A(n7552), .B(n7551), .Z(n7553) );
  AND U12129 ( .A(n23182), .B(n7553), .Z(n7554) );
  NAND U12130 ( .A(n7555), .B(n7554), .Z(n7556) );
  NAND U12131 ( .A(n7557), .B(n7556), .Z(n7558) );
  ANDN U12132 ( .B(y[1650]), .A(x[1650]), .Z(n12355) );
  ANDN U12133 ( .B(n7558), .A(n12355), .Z(n7559) );
  NAND U12134 ( .A(n7560), .B(n7559), .Z(n7561) );
  NAND U12135 ( .A(n7562), .B(n7561), .Z(n7563) );
  AND U12136 ( .A(n23194), .B(n7563), .Z(n7564) );
  NANDN U12137 ( .A(n12353), .B(n7564), .Z(n7565) );
  ANDN U12138 ( .B(x[1653]), .A(y[1653]), .Z(n15267) );
  ANDN U12139 ( .B(x[1654]), .A(y[1654]), .Z(n15271) );
  NOR U12140 ( .A(n15267), .B(n15271), .Z(n23196) );
  NAND U12141 ( .A(n7565), .B(n23196), .Z(n7566) );
  NANDN U12142 ( .A(n23199), .B(n7566), .Z(n7567) );
  NANDN U12143 ( .A(n23201), .B(n7567), .Z(n7572) );
  IV U12144 ( .A(x[1658]), .Z(n20275) );
  NAND U12145 ( .A(y[1658]), .B(n20275), .Z(n23207) );
  XNOR U12146 ( .A(y[1657]), .B(x[1657]), .Z(n7569) );
  NANDN U12147 ( .A(x[1656]), .B(y[1656]), .Z(n7568) );
  NAND U12148 ( .A(n7569), .B(n7568), .Z(n7570) );
  NAND U12149 ( .A(n7571), .B(n7570), .Z(n23202) );
  AND U12150 ( .A(n23207), .B(n23202), .Z(n15275) );
  NAND U12151 ( .A(n7572), .B(n15275), .Z(n7573) );
  NANDN U12152 ( .A(n15278), .B(n7573), .Z(n7574) );
  NANDN U12153 ( .A(x[1659]), .B(y[1659]), .Z(n23208) );
  NAND U12154 ( .A(n7574), .B(n23208), .Z(n7577) );
  NANDN U12155 ( .A(y[1661]), .B(x[1661]), .Z(n7575) );
  NANDN U12156 ( .A(y[1662]), .B(x[1662]), .Z(n15283) );
  NAND U12157 ( .A(n7575), .B(n15283), .Z(n7579) );
  NANDN U12158 ( .A(y[1660]), .B(x[1660]), .Z(n7576) );
  NANDN U12159 ( .A(n7579), .B(n7576), .Z(n23213) );
  ANDN U12160 ( .B(n7577), .A(n23213), .Z(n7582) );
  NANDN U12161 ( .A(x[1665]), .B(y[1665]), .Z(n7578) );
  ANDN U12162 ( .B(y[1664]), .A(x[1664]), .Z(n15292) );
  ANDN U12163 ( .B(n7578), .A(n15292), .Z(n7586) );
  ANDN U12164 ( .B(y[1661]), .A(x[1661]), .Z(n15284) );
  NANDN U12165 ( .A(x[1660]), .B(y[1660]), .Z(n15280) );
  NANDN U12166 ( .A(x[1663]), .B(y[1663]), .Z(n7581) );
  NANDN U12167 ( .A(x[1662]), .B(y[1662]), .Z(n7580) );
  AND U12168 ( .A(n7581), .B(n7580), .Z(n15287) );
  NANDN U12169 ( .A(n7582), .B(n23214), .Z(n7589) );
  NANDN U12170 ( .A(y[1665]), .B(x[1665]), .Z(n7583) );
  ANDN U12171 ( .B(x[1666]), .A(y[1666]), .Z(n15299) );
  ANDN U12172 ( .B(n7583), .A(n15299), .Z(n7588) );
  NANDN U12173 ( .A(y[1663]), .B(x[1663]), .Z(n7585) );
  NANDN U12174 ( .A(y[1664]), .B(x[1664]), .Z(n7584) );
  NAND U12175 ( .A(n7585), .B(n7584), .Z(n15289) );
  NAND U12176 ( .A(n15289), .B(n7586), .Z(n7587) );
  NAND U12177 ( .A(n7588), .B(n7587), .Z(n23216) );
  ANDN U12178 ( .B(n7589), .A(n23216), .Z(n7590) );
  OR U12179 ( .A(n23219), .B(n7590), .Z(n7591) );
  NANDN U12180 ( .A(n23221), .B(n7591), .Z(n7592) );
  NANDN U12181 ( .A(x[1668]), .B(y[1668]), .Z(n23222) );
  NAND U12182 ( .A(n7592), .B(n23222), .Z(n7593) );
  OR U12183 ( .A(n12348), .B(n7593), .Z(n7594) );
  AND U12184 ( .A(n23224), .B(n7594), .Z(n7595) );
  NAND U12185 ( .A(n7596), .B(n7595), .Z(n7597) );
  NAND U12186 ( .A(n7598), .B(n7597), .Z(n7599) );
  AND U12187 ( .A(n23233), .B(n7599), .Z(n7600) );
  NANDN U12188 ( .A(n12346), .B(n7600), .Z(n7601) );
  NANDN U12189 ( .A(x[1673]), .B(y[1673]), .Z(n23234) );
  NAND U12190 ( .A(n7601), .B(n23234), .Z(n7602) );
  OR U12191 ( .A(n12344), .B(n7602), .Z(n7603) );
  NANDN U12192 ( .A(y[1673]), .B(x[1673]), .Z(n15311) );
  NANDN U12193 ( .A(y[1674]), .B(x[1674]), .Z(n12342) );
  NAND U12194 ( .A(n15311), .B(n12342), .Z(n23237) );
  ANDN U12195 ( .B(n7603), .A(n23237), .Z(n7605) );
  NANDN U12196 ( .A(x[1674]), .B(y[1674]), .Z(n7604) );
  ANDN U12197 ( .B(y[1675]), .A(x[1675]), .Z(n12341) );
  ANDN U12198 ( .B(n7604), .A(n12341), .Z(n23238) );
  NANDN U12199 ( .A(n7605), .B(n23238), .Z(n7606) );
  NAND U12200 ( .A(n7607), .B(n7606), .Z(n7608) );
  ANDN U12201 ( .B(y[1677]), .A(x[1677]), .Z(n20271) );
  ANDN U12202 ( .B(y[1676]), .A(x[1676]), .Z(n12340) );
  NOR U12203 ( .A(n20271), .B(n12340), .Z(n23242) );
  NAND U12204 ( .A(n7608), .B(n23242), .Z(n7609) );
  NANDN U12205 ( .A(n20272), .B(n7609), .Z(n7610) );
  AND U12206 ( .A(n23246), .B(n7610), .Z(n7612) );
  NANDN U12207 ( .A(y[1679]), .B(x[1679]), .Z(n7611) );
  ANDN U12208 ( .B(x[1680]), .A(y[1680]), .Z(n15334) );
  ANDN U12209 ( .B(n7611), .A(n15334), .Z(n23248) );
  NANDN U12210 ( .A(n7612), .B(n23248), .Z(n7614) );
  NANDN U12211 ( .A(x[1680]), .B(y[1680]), .Z(n12339) );
  NANDN U12212 ( .A(x[1681]), .B(y[1681]), .Z(n7613) );
  AND U12213 ( .A(n12339), .B(n7613), .Z(n23250) );
  NAND U12214 ( .A(n7614), .B(n23250), .Z(n7616) );
  NANDN U12215 ( .A(y[1681]), .B(x[1681]), .Z(n7615) );
  ANDN U12216 ( .B(x[1682]), .A(y[1682]), .Z(n15340) );
  ANDN U12217 ( .B(n7615), .A(n15340), .Z(n23252) );
  NAND U12218 ( .A(n7616), .B(n23252), .Z(n7617) );
  AND U12219 ( .A(n23254), .B(n7617), .Z(n7618) );
  NANDN U12220 ( .A(n12336), .B(n7618), .Z(n7619) );
  NANDN U12221 ( .A(y[1684]), .B(x[1684]), .Z(n23261) );
  NAND U12222 ( .A(n7619), .B(n23261), .Z(n7620) );
  OR U12223 ( .A(n23256), .B(n7620), .Z(n7621) );
  AND U12224 ( .A(n7622), .B(n7621), .Z(n7623) );
  OR U12225 ( .A(n23265), .B(n7623), .Z(n7624) );
  NANDN U12226 ( .A(n23266), .B(n7624), .Z(n7625) );
  NANDN U12227 ( .A(n23269), .B(n7625), .Z(n7626) );
  NANDN U12228 ( .A(n23271), .B(n7626), .Z(n7627) );
  ANDN U12229 ( .B(x[1690]), .A(y[1690]), .Z(n15361) );
  ANDN U12230 ( .B(n7627), .A(n15361), .Z(n7628) );
  NANDN U12231 ( .A(y[1689]), .B(x[1689]), .Z(n23272) );
  NAND U12232 ( .A(n7628), .B(n23272), .Z(n7629) );
  AND U12233 ( .A(n23274), .B(n7629), .Z(n7630) );
  NAND U12234 ( .A(n7631), .B(n7630), .Z(n7632) );
  NAND U12235 ( .A(n7633), .B(n7632), .Z(n7634) );
  ANDN U12236 ( .B(y[1692]), .A(x[1692]), .Z(n12331) );
  ANDN U12237 ( .B(n7634), .A(n12331), .Z(n7635) );
  NAND U12238 ( .A(n23283), .B(n7635), .Z(n7637) );
  NANDN U12239 ( .A(y[1694]), .B(x[1694]), .Z(n7636) );
  ANDN U12240 ( .B(x[1693]), .A(y[1693]), .Z(n12329) );
  ANDN U12241 ( .B(n7636), .A(n12329), .Z(n23284) );
  NAND U12242 ( .A(n7637), .B(n23284), .Z(n7638) );
  NANDN U12243 ( .A(n23287), .B(n7638), .Z(n7641) );
  NANDN U12244 ( .A(y[1696]), .B(x[1696]), .Z(n7640) );
  NANDN U12245 ( .A(y[1695]), .B(x[1695]), .Z(n7639) );
  AND U12246 ( .A(n7640), .B(n7639), .Z(n23288) );
  NAND U12247 ( .A(n7641), .B(n23288), .Z(n7642) );
  NANDN U12248 ( .A(n23290), .B(n7642), .Z(n7643) );
  AND U12249 ( .A(n23292), .B(n7643), .Z(n7645) );
  NANDN U12250 ( .A(x[1698]), .B(y[1698]), .Z(n7644) );
  ANDN U12251 ( .B(y[1699]), .A(x[1699]), .Z(n15388) );
  ANDN U12252 ( .B(n7644), .A(n15388), .Z(n23294) );
  NANDN U12253 ( .A(n7645), .B(n23294), .Z(n7646) );
  NANDN U12254 ( .A(y[1699]), .B(x[1699]), .Z(n12328) );
  IV U12255 ( .A(y[1700]), .Z(n12326) );
  NAND U12256 ( .A(n12326), .B(x[1700]), .Z(n15393) );
  AND U12257 ( .A(n12328), .B(n15393), .Z(n23296) );
  NAND U12258 ( .A(n7646), .B(n23296), .Z(n7647) );
  ANDN U12259 ( .B(y[1701]), .A(x[1701]), .Z(n15394) );
  NAND U12260 ( .A(n7647), .B(n23299), .Z(n7650) );
  NANDN U12261 ( .A(y[1702]), .B(x[1702]), .Z(n7649) );
  NANDN U12262 ( .A(y[1701]), .B(x[1701]), .Z(n7648) );
  AND U12263 ( .A(n7649), .B(n7648), .Z(n23300) );
  NAND U12264 ( .A(n7650), .B(n23300), .Z(n7651) );
  NANDN U12265 ( .A(n23302), .B(n7651), .Z(n7652) );
  NANDN U12266 ( .A(y[1703]), .B(x[1703]), .Z(n23304) );
  NAND U12267 ( .A(n7652), .B(n23304), .Z(n7653) );
  OR U12268 ( .A(n12321), .B(n7653), .Z(n7655) );
  NANDN U12269 ( .A(x[1704]), .B(y[1704]), .Z(n7654) );
  ANDN U12270 ( .B(y[1705]), .A(x[1705]), .Z(n12322) );
  ANDN U12271 ( .B(n7654), .A(n12322), .Z(n23306) );
  NAND U12272 ( .A(n7655), .B(n23306), .Z(n7656) );
  NANDN U12273 ( .A(n12324), .B(n7656), .Z(n7659) );
  NANDN U12274 ( .A(x[1707]), .B(y[1707]), .Z(n7658) );
  NANDN U12275 ( .A(x[1706]), .B(y[1706]), .Z(n7657) );
  AND U12276 ( .A(n7658), .B(n7657), .Z(n23310) );
  NAND U12277 ( .A(n7659), .B(n23310), .Z(n7662) );
  NANDN U12278 ( .A(y[1707]), .B(x[1707]), .Z(n7661) );
  NANDN U12279 ( .A(y[1708]), .B(x[1708]), .Z(n7660) );
  AND U12280 ( .A(n7661), .B(n7660), .Z(n23313) );
  NAND U12281 ( .A(n7662), .B(n23313), .Z(n7663) );
  AND U12282 ( .A(n23315), .B(n7663), .Z(n7664) );
  NANDN U12283 ( .A(y[1709]), .B(x[1709]), .Z(n23318) );
  NANDN U12284 ( .A(n7664), .B(n23318), .Z(n7665) );
  NANDN U12285 ( .A(n15407), .B(n7665), .Z(n7666) );
  NANDN U12286 ( .A(n12320), .B(n7666), .Z(n7667) );
  NAND U12287 ( .A(n7668), .B(n7667), .Z(n7669) );
  NAND U12288 ( .A(n12319), .B(n7669), .Z(n7670) );
  NAND U12289 ( .A(n7671), .B(n7670), .Z(n7672) );
  NAND U12290 ( .A(n12316), .B(n7672), .Z(n7673) );
  NAND U12291 ( .A(n7674), .B(n7673), .Z(n7675) );
  NAND U12292 ( .A(n12315), .B(n7675), .Z(n7678) );
  NANDN U12293 ( .A(x[1715]), .B(y[1715]), .Z(n7677) );
  NANDN U12294 ( .A(x[1714]), .B(y[1714]), .Z(n7676) );
  NAND U12295 ( .A(n7677), .B(n7676), .Z(n12314) );
  ANDN U12296 ( .B(n7678), .A(n12314), .Z(n7685) );
  NANDN U12297 ( .A(y[1715]), .B(x[1715]), .Z(n7680) );
  ANDN U12298 ( .B(x[1716]), .A(y[1716]), .Z(n7679) );
  ANDN U12299 ( .B(n7680), .A(n7679), .Z(n7684) );
  XNOR U12300 ( .A(x[1715]), .B(y[1715]), .Z(n7682) );
  ANDN U12301 ( .B(x[1714]), .A(y[1714]), .Z(n7681) );
  NAND U12302 ( .A(n7682), .B(n7681), .Z(n7683) );
  AND U12303 ( .A(n7684), .B(n7683), .Z(n23330) );
  NANDN U12304 ( .A(n7685), .B(n23330), .Z(n7688) );
  NANDN U12305 ( .A(x[1716]), .B(y[1716]), .Z(n7687) );
  NANDN U12306 ( .A(x[1717]), .B(y[1717]), .Z(n7686) );
  NAND U12307 ( .A(n7687), .B(n7686), .Z(n23333) );
  ANDN U12308 ( .B(n7688), .A(n23333), .Z(n7690) );
  NANDN U12309 ( .A(y[1717]), .B(x[1717]), .Z(n23334) );
  ANDN U12310 ( .B(x[1718]), .A(y[1718]), .Z(n12311) );
  ANDN U12311 ( .B(n23334), .A(n12311), .Z(n7689) );
  NANDN U12312 ( .A(n7690), .B(n7689), .Z(n7691) );
  AND U12313 ( .A(n23337), .B(n7691), .Z(n7692) );
  OR U12314 ( .A(n12312), .B(n7692), .Z(n7695) );
  NANDN U12315 ( .A(x[1720]), .B(y[1720]), .Z(n7694) );
  NANDN U12316 ( .A(x[1719]), .B(y[1719]), .Z(n7693) );
  NAND U12317 ( .A(n7694), .B(n7693), .Z(n23340) );
  ANDN U12318 ( .B(n7695), .A(n23340), .Z(n7696) );
  NANDN U12319 ( .A(y[1720]), .B(x[1720]), .Z(n23342) );
  NANDN U12320 ( .A(n7696), .B(n23342), .Z(n7697) );
  NANDN U12321 ( .A(x[1721]), .B(y[1721]), .Z(n23344) );
  NAND U12322 ( .A(n7697), .B(n23344), .Z(n7698) );
  ANDN U12323 ( .B(x[1721]), .A(y[1721]), .Z(n15419) );
  XOR U12324 ( .A(x[1722]), .B(y[1722]), .Z(n15424) );
  NOR U12325 ( .A(n15419), .B(n15424), .Z(n23346) );
  NAND U12326 ( .A(n7698), .B(n23346), .Z(n7699) );
  NANDN U12327 ( .A(n23349), .B(n7699), .Z(n7702) );
  NANDN U12328 ( .A(y[1723]), .B(x[1723]), .Z(n7701) );
  NANDN U12329 ( .A(y[1724]), .B(x[1724]), .Z(n7700) );
  AND U12330 ( .A(n7701), .B(n7700), .Z(n23350) );
  NAND U12331 ( .A(n7702), .B(n23350), .Z(n7705) );
  NANDN U12332 ( .A(x[1725]), .B(y[1725]), .Z(n7704) );
  NANDN U12333 ( .A(x[1724]), .B(y[1724]), .Z(n7703) );
  NAND U12334 ( .A(n7704), .B(n7703), .Z(n23352) );
  ANDN U12335 ( .B(n7705), .A(n23352), .Z(n7708) );
  NANDN U12336 ( .A(y[1725]), .B(x[1725]), .Z(n7707) );
  NANDN U12337 ( .A(y[1726]), .B(x[1726]), .Z(n7706) );
  AND U12338 ( .A(n7707), .B(n7706), .Z(n23354) );
  NANDN U12339 ( .A(n7708), .B(n23354), .Z(n7711) );
  NANDN U12340 ( .A(x[1727]), .B(y[1727]), .Z(n7710) );
  NANDN U12341 ( .A(x[1726]), .B(y[1726]), .Z(n7709) );
  NAND U12342 ( .A(n7710), .B(n7709), .Z(n23356) );
  ANDN U12343 ( .B(n7711), .A(n23356), .Z(n7714) );
  NANDN U12344 ( .A(y[1727]), .B(x[1727]), .Z(n7713) );
  NANDN U12345 ( .A(y[1728]), .B(x[1728]), .Z(n7712) );
  AND U12346 ( .A(n7713), .B(n7712), .Z(n23358) );
  NANDN U12347 ( .A(n7714), .B(n23358), .Z(n7717) );
  NANDN U12348 ( .A(x[1729]), .B(y[1729]), .Z(n7716) );
  NANDN U12349 ( .A(x[1728]), .B(y[1728]), .Z(n7715) );
  AND U12350 ( .A(n7716), .B(n7715), .Z(n23360) );
  NAND U12351 ( .A(n7717), .B(n23360), .Z(n7719) );
  NANDN U12352 ( .A(y[1730]), .B(x[1730]), .Z(n7718) );
  ANDN U12353 ( .B(x[1729]), .A(y[1729]), .Z(n15432) );
  ANDN U12354 ( .B(n7718), .A(n15432), .Z(n23363) );
  NAND U12355 ( .A(n7719), .B(n23363), .Z(n7722) );
  NANDN U12356 ( .A(x[1730]), .B(y[1730]), .Z(n7721) );
  ANDN U12357 ( .B(y[1731]), .A(x[1731]), .Z(n7720) );
  ANDN U12358 ( .B(n7721), .A(n7720), .Z(n23364) );
  NAND U12359 ( .A(n7722), .B(n23364), .Z(n7725) );
  NANDN U12360 ( .A(y[1731]), .B(x[1731]), .Z(n7724) );
  NANDN U12361 ( .A(y[1732]), .B(x[1732]), .Z(n7723) );
  AND U12362 ( .A(n7724), .B(n7723), .Z(n23366) );
  NAND U12363 ( .A(n7725), .B(n23366), .Z(n7726) );
  AND U12364 ( .A(n23368), .B(n7726), .Z(n7729) );
  NANDN U12365 ( .A(y[1733]), .B(x[1733]), .Z(n7728) );
  NANDN U12366 ( .A(y[1734]), .B(x[1734]), .Z(n7727) );
  AND U12367 ( .A(n7728), .B(n7727), .Z(n23370) );
  NANDN U12368 ( .A(n7729), .B(n23370), .Z(n7730) );
  AND U12369 ( .A(n23372), .B(n7730), .Z(n7733) );
  NANDN U12370 ( .A(y[1735]), .B(x[1735]), .Z(n7732) );
  NANDN U12371 ( .A(y[1736]), .B(x[1736]), .Z(n7731) );
  AND U12372 ( .A(n7732), .B(n7731), .Z(n23375) );
  NANDN U12373 ( .A(n7733), .B(n23375), .Z(n7734) );
  AND U12374 ( .A(n23376), .B(n7734), .Z(n7737) );
  NANDN U12375 ( .A(y[1738]), .B(x[1738]), .Z(n7736) );
  NANDN U12376 ( .A(y[1737]), .B(x[1737]), .Z(n7735) );
  AND U12377 ( .A(n7736), .B(n7735), .Z(n23379) );
  NANDN U12378 ( .A(n7737), .B(n23379), .Z(n7738) );
  AND U12379 ( .A(n7739), .B(n7738), .Z(n7741) );
  NANDN U12380 ( .A(y[1739]), .B(x[1739]), .Z(n7740) );
  ANDN U12381 ( .B(x[1740]), .A(y[1740]), .Z(n15447) );
  ANDN U12382 ( .B(n7740), .A(n15447), .Z(n23382) );
  NANDN U12383 ( .A(n7741), .B(n23382), .Z(n7744) );
  NANDN U12384 ( .A(x[1741]), .B(y[1741]), .Z(n7743) );
  NANDN U12385 ( .A(x[1740]), .B(y[1740]), .Z(n7742) );
  NAND U12386 ( .A(n7743), .B(n7742), .Z(n15449) );
  ANDN U12387 ( .B(n7744), .A(n15449), .Z(n7747) );
  XNOR U12388 ( .A(x[1742]), .B(y[1742]), .Z(n7746) );
  NANDN U12389 ( .A(y[1741]), .B(x[1741]), .Z(n7745) );
  AND U12390 ( .A(n7746), .B(n7745), .Z(n23386) );
  NANDN U12391 ( .A(n7747), .B(n23386), .Z(n7748) );
  NANDN U12392 ( .A(n23388), .B(n7748), .Z(n7751) );
  NANDN U12393 ( .A(y[1743]), .B(x[1743]), .Z(n7750) );
  NANDN U12394 ( .A(y[1744]), .B(x[1744]), .Z(n7749) );
  AND U12395 ( .A(n7750), .B(n7749), .Z(n23390) );
  NAND U12396 ( .A(n7751), .B(n23390), .Z(n7752) );
  AND U12397 ( .A(n23392), .B(n7752), .Z(n7754) );
  IV U12398 ( .A(y[1746]), .Z(n15458) );
  NAND U12399 ( .A(n15458), .B(x[1746]), .Z(n7753) );
  ANDN U12400 ( .B(x[1745]), .A(y[1745]), .Z(n15456) );
  ANDN U12401 ( .B(n7753), .A(n15456), .Z(n23395) );
  NANDN U12402 ( .A(n7754), .B(n23395), .Z(n7756) );
  NANDN U12403 ( .A(x[1746]), .B(y[1746]), .Z(n7755) );
  ANDN U12404 ( .B(y[1747]), .A(x[1747]), .Z(n15462) );
  ANDN U12405 ( .B(n7755), .A(n15462), .Z(n23396) );
  NAND U12406 ( .A(n7756), .B(n23396), .Z(n7759) );
  NANDN U12407 ( .A(y[1747]), .B(x[1747]), .Z(n7758) );
  NANDN U12408 ( .A(y[1748]), .B(x[1748]), .Z(n7757) );
  AND U12409 ( .A(n7758), .B(n7757), .Z(n23398) );
  NAND U12410 ( .A(n7759), .B(n23398), .Z(n7762) );
  NANDN U12411 ( .A(x[1749]), .B(y[1749]), .Z(n7761) );
  NANDN U12412 ( .A(x[1748]), .B(y[1748]), .Z(n7760) );
  AND U12413 ( .A(n7761), .B(n7760), .Z(n23400) );
  NAND U12414 ( .A(n7762), .B(n23400), .Z(n7764) );
  NANDN U12415 ( .A(y[1750]), .B(x[1750]), .Z(n7763) );
  ANDN U12416 ( .B(x[1749]), .A(y[1749]), .Z(n15466) );
  ANDN U12417 ( .B(n7763), .A(n15466), .Z(n23402) );
  NAND U12418 ( .A(n7764), .B(n23402), .Z(n7766) );
  IV U12419 ( .A(x[1750]), .Z(n15470) );
  NAND U12420 ( .A(n15470), .B(y[1750]), .Z(n7765) );
  NANDN U12421 ( .A(x[1751]), .B(y[1751]), .Z(n12309) );
  NAND U12422 ( .A(n7765), .B(n12309), .Z(n23405) );
  ANDN U12423 ( .B(n7766), .A(n23405), .Z(n7768) );
  NANDN U12424 ( .A(y[1751]), .B(x[1751]), .Z(n7767) );
  ANDN U12425 ( .B(x[1752]), .A(y[1752]), .Z(n15477) );
  ANDN U12426 ( .B(n7767), .A(n15477), .Z(n23406) );
  NANDN U12427 ( .A(n7768), .B(n23406), .Z(n7769) );
  NANDN U12428 ( .A(n23409), .B(n7769), .Z(n7770) );
  NANDN U12429 ( .A(y[1753]), .B(x[1753]), .Z(n23410) );
  NAND U12430 ( .A(n7770), .B(n23410), .Z(n7771) );
  OR U12431 ( .A(n12305), .B(n7771), .Z(n7772) );
  AND U12432 ( .A(n23413), .B(n7772), .Z(n7773) );
  OR U12433 ( .A(n12308), .B(n7773), .Z(n7776) );
  NANDN U12434 ( .A(x[1757]), .B(y[1757]), .Z(n7775) );
  NANDN U12435 ( .A(x[1756]), .B(y[1756]), .Z(n7774) );
  NAND U12436 ( .A(n7775), .B(n7774), .Z(n23417) );
  ANDN U12437 ( .B(n7776), .A(n23417), .Z(n7779) );
  NANDN U12438 ( .A(y[1757]), .B(x[1757]), .Z(n7778) );
  NANDN U12439 ( .A(y[1758]), .B(x[1758]), .Z(n7777) );
  AND U12440 ( .A(n7778), .B(n7777), .Z(n23418) );
  NANDN U12441 ( .A(n7779), .B(n23418), .Z(n7780) );
  NANDN U12442 ( .A(n23421), .B(n7780), .Z(n7781) );
  NANDN U12443 ( .A(y[1759]), .B(x[1759]), .Z(n23422) );
  NAND U12444 ( .A(n7781), .B(n23422), .Z(n7782) );
  OR U12445 ( .A(n15489), .B(n7782), .Z(n7783) );
  AND U12446 ( .A(n23425), .B(n7783), .Z(n7784) );
  OR U12447 ( .A(n15490), .B(n7784), .Z(n7785) );
  NANDN U12448 ( .A(n23429), .B(n7785), .Z(n7786) );
  NANDN U12449 ( .A(y[1762]), .B(x[1762]), .Z(n23430) );
  NAND U12450 ( .A(n7786), .B(n23430), .Z(n7787) );
  NANDN U12451 ( .A(x[1763]), .B(y[1763]), .Z(n23432) );
  NAND U12452 ( .A(n7787), .B(n23432), .Z(n7788) );
  XNOR U12453 ( .A(x[1764]), .B(y[1764]), .Z(n15496) );
  ANDN U12454 ( .B(x[1763]), .A(y[1763]), .Z(n15493) );
  ANDN U12455 ( .B(n15496), .A(n15493), .Z(n23434) );
  NAND U12456 ( .A(n7788), .B(n23434), .Z(n7789) );
  ANDN U12457 ( .B(y[1765]), .A(x[1765]), .Z(n12303) );
  IV U12458 ( .A(y[1764]), .Z(n15500) );
  ANDN U12459 ( .B(n7789), .A(n23436), .Z(n7791) );
  NANDN U12460 ( .A(y[1765]), .B(x[1765]), .Z(n7790) );
  ANDN U12461 ( .B(x[1766]), .A(y[1766]), .Z(n12304) );
  ANDN U12462 ( .B(n7790), .A(n12304), .Z(n23438) );
  NANDN U12463 ( .A(n7791), .B(n23438), .Z(n7794) );
  NANDN U12464 ( .A(x[1767]), .B(y[1767]), .Z(n7793) );
  NANDN U12465 ( .A(x[1766]), .B(y[1766]), .Z(n7792) );
  NAND U12466 ( .A(n7793), .B(n7792), .Z(n23440) );
  ANDN U12467 ( .B(n7794), .A(n23440), .Z(n7797) );
  NANDN U12468 ( .A(y[1767]), .B(x[1767]), .Z(n7796) );
  NANDN U12469 ( .A(y[1768]), .B(x[1768]), .Z(n7795) );
  AND U12470 ( .A(n7796), .B(n7795), .Z(n23442) );
  NANDN U12471 ( .A(n7797), .B(n23442), .Z(n7800) );
  NANDN U12472 ( .A(x[1769]), .B(y[1769]), .Z(n7799) );
  NANDN U12473 ( .A(x[1768]), .B(y[1768]), .Z(n7798) );
  NAND U12474 ( .A(n7799), .B(n7798), .Z(n23445) );
  ANDN U12475 ( .B(n7800), .A(n23445), .Z(n7803) );
  NANDN U12476 ( .A(y[1769]), .B(x[1769]), .Z(n7802) );
  NANDN U12477 ( .A(y[1770]), .B(x[1770]), .Z(n7801) );
  AND U12478 ( .A(n7802), .B(n7801), .Z(n23446) );
  NANDN U12479 ( .A(n7803), .B(n23446), .Z(n7804) );
  NANDN U12480 ( .A(n23449), .B(n7804), .Z(n7807) );
  NANDN U12481 ( .A(y[1771]), .B(x[1771]), .Z(n7806) );
  NANDN U12482 ( .A(y[1772]), .B(x[1772]), .Z(n7805) );
  AND U12483 ( .A(n7806), .B(n7805), .Z(n23450) );
  NAND U12484 ( .A(n7807), .B(n23450), .Z(n7810) );
  NANDN U12485 ( .A(x[1773]), .B(y[1773]), .Z(n7809) );
  NANDN U12486 ( .A(x[1772]), .B(y[1772]), .Z(n7808) );
  AND U12487 ( .A(n7809), .B(n7808), .Z(n23453) );
  NAND U12488 ( .A(n7810), .B(n23453), .Z(n7811) );
  AND U12489 ( .A(n23454), .B(n7811), .Z(n7812) );
  NANDN U12490 ( .A(n12299), .B(n7812), .Z(n7814) );
  NANDN U12491 ( .A(x[1774]), .B(y[1774]), .Z(n7813) );
  ANDN U12492 ( .B(y[1775]), .A(x[1775]), .Z(n12300) );
  ANDN U12493 ( .B(n7813), .A(n12300), .Z(n23456) );
  NAND U12494 ( .A(n7814), .B(n23456), .Z(n7815) );
  NANDN U12495 ( .A(n12302), .B(n7815), .Z(n7818) );
  NANDN U12496 ( .A(x[1777]), .B(y[1777]), .Z(n7817) );
  NANDN U12497 ( .A(x[1776]), .B(y[1776]), .Z(n7816) );
  NAND U12498 ( .A(n7817), .B(n7816), .Z(n23461) );
  ANDN U12499 ( .B(n7818), .A(n23461), .Z(n7819) );
  OR U12500 ( .A(n23463), .B(n7819), .Z(n7820) );
  NANDN U12501 ( .A(n23464), .B(n7820), .Z(n7823) );
  NANDN U12502 ( .A(y[1780]), .B(x[1780]), .Z(n7822) );
  NANDN U12503 ( .A(y[1779]), .B(x[1779]), .Z(n7821) );
  AND U12504 ( .A(n7822), .B(n7821), .Z(n23466) );
  NAND U12505 ( .A(n7823), .B(n23466), .Z(n7824) );
  ANDN U12506 ( .B(y[1781]), .A(x[1781]), .Z(n12297) );
  ANDN U12507 ( .B(n7824), .A(n12297), .Z(n7825) );
  NANDN U12508 ( .A(x[1780]), .B(y[1780]), .Z(n23468) );
  NAND U12509 ( .A(n7825), .B(n23468), .Z(n7826) );
  NANDN U12510 ( .A(y[1781]), .B(x[1781]), .Z(n15525) );
  ANDN U12511 ( .B(x[1782]), .A(y[1782]), .Z(n23473) );
  ANDN U12512 ( .B(n15525), .A(n23473), .Z(n23470) );
  NAND U12513 ( .A(n7826), .B(n23470), .Z(n7827) );
  NAND U12514 ( .A(n7828), .B(n7827), .Z(n7829) );
  NANDN U12515 ( .A(y[1784]), .B(x[1784]), .Z(n15527) );
  NANDN U12516 ( .A(y[1783]), .B(x[1783]), .Z(n15526) );
  NAND U12517 ( .A(n15527), .B(n15526), .Z(n23479) );
  ANDN U12518 ( .B(n7829), .A(n23479), .Z(n7832) );
  NANDN U12519 ( .A(x[1784]), .B(y[1784]), .Z(n7831) );
  NANDN U12520 ( .A(x[1785]), .B(y[1785]), .Z(n7830) );
  AND U12521 ( .A(n7831), .B(n7830), .Z(n23480) );
  NANDN U12522 ( .A(n7832), .B(n23480), .Z(n7833) );
  AND U12523 ( .A(n23482), .B(n7833), .Z(n7834) );
  OR U12524 ( .A(n23485), .B(n7834), .Z(n7835) );
  NAND U12525 ( .A(n7836), .B(n7835), .Z(n7837) );
  NANDN U12526 ( .A(x[1788]), .B(y[1788]), .Z(n23489) );
  NAND U12527 ( .A(n7837), .B(n23489), .Z(n7838) );
  NAND U12528 ( .A(n7839), .B(n7838), .Z(n7840) );
  NAND U12529 ( .A(n12293), .B(n7840), .Z(n7841) );
  NAND U12530 ( .A(n7842), .B(n7841), .Z(n7843) );
  AND U12531 ( .A(n7844), .B(n7843), .Z(n7845) );
  ANDN U12532 ( .B(x[1791]), .A(y[1791]), .Z(n12292) );
  NOR U12533 ( .A(n7845), .B(n12292), .Z(n7847) );
  XNOR U12534 ( .A(x[1792]), .B(y[1792]), .Z(n7846) );
  NAND U12535 ( .A(n7847), .B(n7846), .Z(n7848) );
  NANDN U12536 ( .A(n23500), .B(n7848), .Z(n7851) );
  NANDN U12537 ( .A(y[1793]), .B(x[1793]), .Z(n7850) );
  NANDN U12538 ( .A(y[1794]), .B(x[1794]), .Z(n7849) );
  AND U12539 ( .A(n7850), .B(n7849), .Z(n23502) );
  NAND U12540 ( .A(n7851), .B(n23502), .Z(n7852) );
  NANDN U12541 ( .A(x[1794]), .B(y[1794]), .Z(n23504) );
  NAND U12542 ( .A(n7852), .B(n23504), .Z(n7853) );
  OR U12543 ( .A(n15532), .B(n7853), .Z(n7855) );
  NANDN U12544 ( .A(y[1795]), .B(x[1795]), .Z(n7854) );
  ANDN U12545 ( .B(x[1796]), .A(y[1796]), .Z(n15533) );
  ANDN U12546 ( .B(n7854), .A(n15533), .Z(n23506) );
  NAND U12547 ( .A(n7855), .B(n23506), .Z(n7856) );
  NANDN U12548 ( .A(n15535), .B(n7856), .Z(n7857) );
  NANDN U12549 ( .A(y[1797]), .B(x[1797]), .Z(n23511) );
  NAND U12550 ( .A(n7857), .B(n23511), .Z(n7858) );
  NANDN U12551 ( .A(n23515), .B(n7858), .Z(n7863) );
  NANDN U12552 ( .A(y[1798]), .B(x[1798]), .Z(n23512) );
  OR U12553 ( .A(n7859), .B(n23512), .Z(n7862) );
  NANDN U12554 ( .A(y[1800]), .B(x[1800]), .Z(n7861) );
  NANDN U12555 ( .A(y[1799]), .B(x[1799]), .Z(n7860) );
  AND U12556 ( .A(n7861), .B(n7860), .Z(n23516) );
  NAND U12557 ( .A(n7862), .B(n23516), .Z(n15540) );
  ANDN U12558 ( .B(n7863), .A(n15540), .Z(n7866) );
  NANDN U12559 ( .A(x[1801]), .B(y[1801]), .Z(n7865) );
  NANDN U12560 ( .A(x[1800]), .B(y[1800]), .Z(n7864) );
  AND U12561 ( .A(n7865), .B(n7864), .Z(n23519) );
  NANDN U12562 ( .A(n7866), .B(n23519), .Z(n7867) );
  ANDN U12563 ( .B(x[1802]), .A(y[1802]), .Z(n15545) );
  ANDN U12564 ( .B(n7867), .A(n15545), .Z(n7868) );
  NANDN U12565 ( .A(y[1801]), .B(x[1801]), .Z(n23520) );
  NAND U12566 ( .A(n7868), .B(n23520), .Z(n7869) );
  ANDN U12567 ( .B(y[1803]), .A(x[1803]), .Z(n12289) );
  ANDN U12568 ( .B(n7869), .A(n12289), .Z(n7870) );
  NANDN U12569 ( .A(x[1802]), .B(y[1802]), .Z(n23522) );
  NAND U12570 ( .A(n7870), .B(n23522), .Z(n7871) );
  NANDN U12571 ( .A(y[1804]), .B(x[1804]), .Z(n23528) );
  AND U12572 ( .A(n7871), .B(n23528), .Z(n7872) );
  NANDN U12573 ( .A(n15544), .B(n7872), .Z(n7873) );
  NANDN U12574 ( .A(n23530), .B(n7873), .Z(n7874) );
  OR U12575 ( .A(n12290), .B(n7874), .Z(n7875) );
  AND U12576 ( .A(n23532), .B(n7875), .Z(n7876) );
  OR U12577 ( .A(n23535), .B(n7876), .Z(n7877) );
  AND U12578 ( .A(n23536), .B(n7877), .Z(n7879) );
  NANDN U12579 ( .A(x[1808]), .B(y[1808]), .Z(n23538) );
  ANDN U12580 ( .B(y[1809]), .A(x[1809]), .Z(n12285) );
  ANDN U12581 ( .B(n23538), .A(n12285), .Z(n7878) );
  NANDN U12582 ( .A(n7879), .B(n7878), .Z(n7880) );
  NANDN U12583 ( .A(y[1810]), .B(x[1810]), .Z(n23544) );
  NAND U12584 ( .A(n7880), .B(n23544), .Z(n7881) );
  NANDN U12585 ( .A(y[1809]), .B(x[1809]), .Z(n23540) );
  NANDN U12586 ( .A(n7881), .B(n23540), .Z(n7882) );
  AND U12587 ( .A(n7883), .B(n7882), .Z(n7885) );
  IV U12588 ( .A(y[1812]), .Z(n15568) );
  NAND U12589 ( .A(n15568), .B(x[1812]), .Z(n7884) );
  ANDN U12590 ( .B(x[1811]), .A(y[1811]), .Z(n12284) );
  ANDN U12591 ( .B(n7884), .A(n12284), .Z(n23548) );
  NANDN U12592 ( .A(n7885), .B(n23548), .Z(n7886) );
  NANDN U12593 ( .A(n23551), .B(n7886), .Z(n7887) );
  NANDN U12594 ( .A(n23553), .B(n7887), .Z(n7888) );
  ANDN U12595 ( .B(y[1815]), .A(x[1815]), .Z(n12281) );
  NAND U12596 ( .A(n7888), .B(n23554), .Z(n7889) );
  ANDN U12597 ( .B(x[1815]), .A(y[1815]), .Z(n23556) );
  ANDN U12598 ( .B(n7889), .A(n23556), .Z(n7890) );
  IV U12599 ( .A(y[1816]), .Z(n12280) );
  NANDN U12600 ( .A(n7890), .B(n12280), .Z(n7893) );
  XOR U12601 ( .A(y[1816]), .B(n7890), .Z(n7891) );
  NAND U12602 ( .A(n7891), .B(x[1816]), .Z(n7892) );
  NAND U12603 ( .A(n7893), .B(n7892), .Z(n7894) );
  ANDN U12604 ( .B(y[1817]), .A(x[1817]), .Z(n23560) );
  ANDN U12605 ( .B(n7894), .A(n23560), .Z(n7895) );
  OR U12606 ( .A(n23565), .B(n7895), .Z(n7896) );
  AND U12607 ( .A(n23566), .B(n7896), .Z(n7898) );
  NANDN U12608 ( .A(y[1819]), .B(x[1819]), .Z(n7897) );
  ANDN U12609 ( .B(x[1820]), .A(y[1820]), .Z(n12277) );
  ANDN U12610 ( .B(n7897), .A(n12277), .Z(n23569) );
  NANDN U12611 ( .A(n7898), .B(n23569), .Z(n7900) );
  NANDN U12612 ( .A(x[1820]), .B(y[1820]), .Z(n7899) );
  ANDN U12613 ( .B(y[1821]), .A(x[1821]), .Z(n12278) );
  ANDN U12614 ( .B(n7899), .A(n12278), .Z(n23570) );
  NAND U12615 ( .A(n7900), .B(n23570), .Z(n7903) );
  NANDN U12616 ( .A(y[1822]), .B(x[1822]), .Z(n7902) );
  NANDN U12617 ( .A(y[1821]), .B(x[1821]), .Z(n7901) );
  AND U12618 ( .A(n7902), .B(n7901), .Z(n23573) );
  NAND U12619 ( .A(n7903), .B(n23573), .Z(n7904) );
  NANDN U12620 ( .A(x[1822]), .B(y[1822]), .Z(n23574) );
  AND U12621 ( .A(n7904), .B(n23574), .Z(n7905) );
  NANDN U12622 ( .A(n12276), .B(n7905), .Z(n7906) );
  NANDN U12623 ( .A(n23577), .B(n7906), .Z(n7908) );
  NANDN U12624 ( .A(y[1824]), .B(n7908), .Z(n7907) );
  ANDN U12625 ( .B(x[1825]), .A(y[1825]), .Z(n23587) );
  ANDN U12626 ( .B(n7907), .A(n23587), .Z(n7911) );
  XNOR U12627 ( .A(n7908), .B(y[1824]), .Z(n7909) );
  NAND U12628 ( .A(x[1824]), .B(n7909), .Z(n7910) );
  NAND U12629 ( .A(n7911), .B(n7910), .Z(n7912) );
  NANDN U12630 ( .A(x[1825]), .B(y[1825]), .Z(n23582) );
  NANDN U12631 ( .A(x[1826]), .B(y[1826]), .Z(n23590) );
  AND U12632 ( .A(n23582), .B(n23590), .Z(n15601) );
  NAND U12633 ( .A(n7912), .B(n15601), .Z(n7913) );
  ANDN U12634 ( .B(x[1827]), .A(y[1827]), .Z(n23593) );
  ANDN U12635 ( .B(x[1826]), .A(y[1826]), .Z(n23584) );
  NOR U12636 ( .A(n23593), .B(n23584), .Z(n15603) );
  NAND U12637 ( .A(n7913), .B(n15603), .Z(n7914) );
  AND U12638 ( .A(n23589), .B(n7914), .Z(n7915) );
  NANDN U12639 ( .A(y[1828]), .B(x[1828]), .Z(n23594) );
  NANDN U12640 ( .A(n7915), .B(n23594), .Z(n7916) );
  NANDN U12641 ( .A(n23597), .B(n7916), .Z(n7917) );
  NANDN U12642 ( .A(n12272), .B(n7917), .Z(n7918) );
  OR U12643 ( .A(n23598), .B(n7918), .Z(n7919) );
  NANDN U12644 ( .A(x[1830]), .B(y[1830]), .Z(n23600) );
  NAND U12645 ( .A(n7919), .B(n23600), .Z(n7920) );
  NANDN U12646 ( .A(n12273), .B(n7920), .Z(n7923) );
  NANDN U12647 ( .A(x[1832]), .B(y[1832]), .Z(n7922) );
  NANDN U12648 ( .A(x[1831]), .B(y[1831]), .Z(n7921) );
  AND U12649 ( .A(n7922), .B(n7921), .Z(n23604) );
  NAND U12650 ( .A(n7923), .B(n23604), .Z(n7925) );
  NANDN U12651 ( .A(y[1833]), .B(x[1833]), .Z(n7924) );
  ANDN U12652 ( .B(x[1832]), .A(y[1832]), .Z(n23607) );
  ANDN U12653 ( .B(n7924), .A(n23607), .Z(n15614) );
  NAND U12654 ( .A(n7925), .B(n15614), .Z(n7927) );
  NANDN U12655 ( .A(x[1834]), .B(y[1834]), .Z(n23616) );
  IV U12656 ( .A(x[1833]), .Z(n23610) );
  NAND U12657 ( .A(n23610), .B(y[1833]), .Z(n7926) );
  NAND U12658 ( .A(n23616), .B(n7926), .Z(n15617) );
  ANDN U12659 ( .B(n7927), .A(n15617), .Z(n7929) );
  NANDN U12660 ( .A(y[1834]), .B(x[1834]), .Z(n7928) );
  ANDN U12661 ( .B(x[1835]), .A(y[1835]), .Z(n23617) );
  ANDN U12662 ( .B(n7928), .A(n23617), .Z(n15618) );
  NANDN U12663 ( .A(n7929), .B(n15618), .Z(n7932) );
  NANDN U12664 ( .A(x[1836]), .B(y[1836]), .Z(n7931) );
  NANDN U12665 ( .A(x[1835]), .B(y[1835]), .Z(n7930) );
  AND U12666 ( .A(n7931), .B(n7930), .Z(n23619) );
  NAND U12667 ( .A(n7932), .B(n23619), .Z(n7933) );
  NANDN U12668 ( .A(n12271), .B(n7933), .Z(n7934) );
  NANDN U12669 ( .A(y[1838]), .B(x[1838]), .Z(n23625) );
  ANDN U12670 ( .B(y[1838]), .A(x[1838]), .Z(n12268) );
  NANDN U12671 ( .A(y[1839]), .B(x[1839]), .Z(n23630) );
  ANDN U12672 ( .B(x[1841]), .A(y[1841]), .Z(n23635) );
  ANDN U12673 ( .B(x[1840]), .A(y[1840]), .Z(n23632) );
  NOR U12674 ( .A(n23635), .B(n23632), .Z(n15629) );
  NANDN U12675 ( .A(y[1842]), .B(x[1842]), .Z(n23637) );
  ANDN U12676 ( .B(y[1843]), .A(x[1843]), .Z(n12267) );
  ANDN U12677 ( .B(y[1842]), .A(x[1842]), .Z(n15630) );
  NOR U12678 ( .A(n12267), .B(n15630), .Z(n23639) );
  ANDN U12679 ( .B(x[1844]), .A(y[1844]), .Z(n15639) );
  NANDN U12680 ( .A(y[1843]), .B(x[1843]), .Z(n23641) );
  NANDN U12681 ( .A(y[1845]), .B(x[1845]), .Z(n15638) );
  NANDN U12682 ( .A(y[1847]), .B(x[1847]), .Z(n7937) );
  NANDN U12683 ( .A(y[1846]), .B(x[1846]), .Z(n7936) );
  NAND U12684 ( .A(n7937), .B(n7936), .Z(n15642) );
  NANDN U12685 ( .A(x[1847]), .B(y[1847]), .Z(n23647) );
  NAND U12686 ( .A(n7938), .B(n23647), .Z(n7939) );
  ANDN U12687 ( .B(x[1848]), .A(y[1848]), .Z(n23650) );
  ANDN U12688 ( .B(n7939), .A(n23650), .Z(n7941) );
  IV U12689 ( .A(x[1849]), .Z(n15650) );
  NAND U12690 ( .A(n15650), .B(y[1849]), .Z(n7940) );
  ANDN U12691 ( .B(y[1848]), .A(x[1848]), .Z(n12266) );
  ANDN U12692 ( .B(n7940), .A(n12266), .Z(n23651) );
  NANDN U12693 ( .A(n7941), .B(n23651), .Z(n7942) );
  NANDN U12694 ( .A(n23653), .B(n7942), .Z(n7943) );
  NANDN U12695 ( .A(x[1850]), .B(y[1850]), .Z(n23655) );
  NAND U12696 ( .A(n7943), .B(n23655), .Z(n7944) );
  OR U12697 ( .A(n12261), .B(n7944), .Z(n7946) );
  NANDN U12698 ( .A(y[1851]), .B(x[1851]), .Z(n7945) );
  ANDN U12699 ( .B(x[1852]), .A(y[1852]), .Z(n12262) );
  ANDN U12700 ( .B(n7945), .A(n12262), .Z(n23658) );
  NAND U12701 ( .A(n7946), .B(n23658), .Z(n7947) );
  NANDN U12702 ( .A(n12264), .B(n7947), .Z(n7950) );
  NANDN U12703 ( .A(y[1854]), .B(x[1854]), .Z(n7949) );
  NANDN U12704 ( .A(y[1853]), .B(x[1853]), .Z(n7948) );
  NAND U12705 ( .A(n7949), .B(n7948), .Z(n23662) );
  ANDN U12706 ( .B(n7950), .A(n23662), .Z(n7953) );
  NANDN U12707 ( .A(x[1854]), .B(y[1854]), .Z(n7952) );
  NANDN U12708 ( .A(x[1855]), .B(y[1855]), .Z(n7951) );
  AND U12709 ( .A(n7952), .B(n7951), .Z(n23663) );
  NANDN U12710 ( .A(n7953), .B(n23663), .Z(n7954) );
  NANDN U12711 ( .A(n23666), .B(n7954), .Z(n7955) );
  ANDN U12712 ( .B(y[1857]), .A(x[1857]), .Z(n12260) );
  NAND U12713 ( .A(n7955), .B(n23667), .Z(n7956) );
  AND U12714 ( .A(n23670), .B(n7956), .Z(n7957) );
  NANDN U12715 ( .A(n12259), .B(n7957), .Z(n7958) );
  NANDN U12716 ( .A(x[1858]), .B(y[1858]), .Z(n23671) );
  NAND U12717 ( .A(n7958), .B(n23671), .Z(n7959) );
  NAND U12718 ( .A(n7960), .B(n7959), .Z(n7961) );
  NAND U12719 ( .A(n12256), .B(n7961), .Z(n7962) );
  NAND U12720 ( .A(n7963), .B(n7962), .Z(n7964) );
  NAND U12721 ( .A(n7965), .B(n7964), .Z(n7968) );
  NANDN U12722 ( .A(y[1864]), .B(x[1864]), .Z(n12254) );
  NANDN U12723 ( .A(y[1863]), .B(x[1863]), .Z(n7966) );
  NAND U12724 ( .A(n12254), .B(n7966), .Z(n7971) );
  NANDN U12725 ( .A(y[1862]), .B(x[1862]), .Z(n7967) );
  NANDN U12726 ( .A(n7971), .B(n7967), .Z(n23681) );
  ANDN U12727 ( .B(n7968), .A(n23681), .Z(n7969) );
  NANDN U12728 ( .A(n15671), .B(n7969), .Z(n7975) );
  NANDN U12729 ( .A(x[1863]), .B(y[1863]), .Z(n12255) );
  NANDN U12730 ( .A(x[1862]), .B(y[1862]), .Z(n15673) );
  NAND U12731 ( .A(n12255), .B(n15673), .Z(n7970) );
  NANDN U12732 ( .A(n7971), .B(n7970), .Z(n7974) );
  NANDN U12733 ( .A(x[1864]), .B(y[1864]), .Z(n7973) );
  NANDN U12734 ( .A(x[1865]), .B(y[1865]), .Z(n7972) );
  NAND U12735 ( .A(n7973), .B(n7972), .Z(n15677) );
  ANDN U12736 ( .B(n7974), .A(n15677), .Z(n23683) );
  NAND U12737 ( .A(n7975), .B(n23683), .Z(n7976) );
  NANDN U12738 ( .A(n23685), .B(n7976), .Z(n7977) );
  NANDN U12739 ( .A(n23688), .B(n7977), .Z(n7978) );
  NANDN U12740 ( .A(y[1867]), .B(x[1867]), .Z(n23690) );
  NAND U12741 ( .A(n7978), .B(n23690), .Z(n7979) );
  NANDN U12742 ( .A(x[1868]), .B(y[1868]), .Z(n20269) );
  NAND U12743 ( .A(n7979), .B(n20269), .Z(n7980) );
  ANDN U12744 ( .B(x[1869]), .A(y[1869]), .Z(n23695) );
  ANDN U12745 ( .B(x[1868]), .A(y[1868]), .Z(n23692) );
  NOR U12746 ( .A(n23695), .B(n23692), .Z(n15685) );
  NAND U12747 ( .A(n7980), .B(n15685), .Z(n7981) );
  AND U12748 ( .A(n20268), .B(n7981), .Z(n7982) );
  NANDN U12749 ( .A(y[1870]), .B(x[1870]), .Z(n23697) );
  NANDN U12750 ( .A(n7982), .B(n23697), .Z(n7983) );
  AND U12751 ( .A(n23699), .B(n7983), .Z(n7984) );
  NANDN U12752 ( .A(y[1872]), .B(x[1872]), .Z(n20267) );
  NANDN U12753 ( .A(y[1871]), .B(x[1871]), .Z(n23701) );
  AND U12754 ( .A(n20267), .B(n23701), .Z(n15690) );
  NANDN U12755 ( .A(n7984), .B(n15690), .Z(n7985) );
  NANDN U12756 ( .A(x[1873]), .B(y[1873]), .Z(n20266) );
  ANDN U12757 ( .B(y[1872]), .A(x[1872]), .Z(n15697) );
  ANDN U12758 ( .B(n20266), .A(n15697), .Z(n23703) );
  NAND U12759 ( .A(n7985), .B(n23703), .Z(n7987) );
  NANDN U12760 ( .A(y[1873]), .B(x[1873]), .Z(n7986) );
  NANDN U12761 ( .A(y[1874]), .B(x[1874]), .Z(n15703) );
  NAND U12762 ( .A(n7986), .B(n15703), .Z(n23705) );
  ANDN U12763 ( .B(n7987), .A(n23705), .Z(n7990) );
  NANDN U12764 ( .A(x[1874]), .B(y[1874]), .Z(n7989) );
  NANDN U12765 ( .A(x[1875]), .B(y[1875]), .Z(n7988) );
  AND U12766 ( .A(n7989), .B(n7988), .Z(n23709) );
  NANDN U12767 ( .A(n7990), .B(n23709), .Z(n7992) );
  NANDN U12768 ( .A(y[1876]), .B(x[1876]), .Z(n7991) );
  NANDN U12769 ( .A(y[1875]), .B(x[1875]), .Z(n15706) );
  NAND U12770 ( .A(n7991), .B(n15706), .Z(n23712) );
  ANDN U12771 ( .B(n7992), .A(n23712), .Z(n7993) );
  OR U12772 ( .A(n23714), .B(n7993), .Z(n7994) );
  NANDN U12773 ( .A(n23715), .B(n7994), .Z(n7995) );
  NANDN U12774 ( .A(x[1878]), .B(y[1878]), .Z(n23717) );
  NAND U12775 ( .A(n7995), .B(n23717), .Z(n7996) );
  OR U12776 ( .A(n12250), .B(n7996), .Z(n7997) );
  AND U12777 ( .A(n23719), .B(n7997), .Z(n7998) );
  NAND U12778 ( .A(n7999), .B(n7998), .Z(n8000) );
  NAND U12779 ( .A(n8001), .B(n8000), .Z(n8004) );
  ANDN U12780 ( .B(x[1884]), .A(y[1884]), .Z(n12246) );
  NANDN U12781 ( .A(y[1883]), .B(x[1883]), .Z(n8002) );
  NANDN U12782 ( .A(n12246), .B(n8002), .Z(n8007) );
  NANDN U12783 ( .A(y[1882]), .B(x[1882]), .Z(n8003) );
  NANDN U12784 ( .A(n8007), .B(n8003), .Z(n23728) );
  ANDN U12785 ( .B(n8004), .A(n23728), .Z(n8005) );
  NANDN U12786 ( .A(n15720), .B(n8005), .Z(n8011) );
  ANDN U12787 ( .B(y[1883]), .A(x[1883]), .Z(n12245) );
  NANDN U12788 ( .A(x[1882]), .B(y[1882]), .Z(n15722) );
  NANDN U12789 ( .A(n12245), .B(n15722), .Z(n8006) );
  NANDN U12790 ( .A(n8007), .B(n8006), .Z(n8010) );
  NANDN U12791 ( .A(x[1884]), .B(y[1884]), .Z(n8009) );
  NANDN U12792 ( .A(x[1885]), .B(y[1885]), .Z(n8008) );
  NAND U12793 ( .A(n8009), .B(n8008), .Z(n12248) );
  ANDN U12794 ( .B(n8010), .A(n12248), .Z(n23729) );
  NAND U12795 ( .A(n8011), .B(n23729), .Z(n8014) );
  NANDN U12796 ( .A(y[1886]), .B(x[1886]), .Z(n8013) );
  NANDN U12797 ( .A(y[1885]), .B(x[1885]), .Z(n8012) );
  AND U12798 ( .A(n8013), .B(n8012), .Z(n23731) );
  NAND U12799 ( .A(n8014), .B(n23731), .Z(n8017) );
  NANDN U12800 ( .A(x[1886]), .B(y[1886]), .Z(n8016) );
  NANDN U12801 ( .A(x[1887]), .B(y[1887]), .Z(n8015) );
  AND U12802 ( .A(n8016), .B(n8015), .Z(n23734) );
  NAND U12803 ( .A(n8017), .B(n23734), .Z(n8018) );
  AND U12804 ( .A(n23735), .B(n8018), .Z(n8020) );
  IV U12805 ( .A(x[1889]), .Z(n15736) );
  NAND U12806 ( .A(n15736), .B(y[1889]), .Z(n8019) );
  ANDN U12807 ( .B(y[1888]), .A(x[1888]), .Z(n15732) );
  ANDN U12808 ( .B(n8019), .A(n15732), .Z(n23737) );
  NANDN U12809 ( .A(n8020), .B(n23737), .Z(n8022) );
  NANDN U12810 ( .A(y[1889]), .B(x[1889]), .Z(n8021) );
  ANDN U12811 ( .B(x[1890]), .A(y[1890]), .Z(n15741) );
  ANDN U12812 ( .B(n8021), .A(n15741), .Z(n23739) );
  NAND U12813 ( .A(n8022), .B(n23739), .Z(n8023) );
  NANDN U12814 ( .A(n23742), .B(n8023), .Z(n8025) );
  NANDN U12815 ( .A(y[1891]), .B(x[1891]), .Z(n8024) );
  ANDN U12816 ( .B(x[1892]), .A(y[1892]), .Z(n15747) );
  ANDN U12817 ( .B(n8024), .A(n15747), .Z(n23743) );
  NAND U12818 ( .A(n8025), .B(n23743), .Z(n8026) );
  ANDN U12819 ( .B(y[1893]), .A(x[1893]), .Z(n15750) );
  ANDN U12820 ( .B(n8026), .A(n15750), .Z(n8027) );
  NANDN U12821 ( .A(x[1892]), .B(y[1892]), .Z(n23746) );
  NAND U12822 ( .A(n8027), .B(n23746), .Z(n8028) );
  NANDN U12823 ( .A(n8029), .B(n8028), .Z(n8030) );
  ANDN U12824 ( .B(y[1894]), .A(x[1894]), .Z(n15751) );
  ANDN U12825 ( .B(n8030), .A(n15751), .Z(n8031) );
  NANDN U12826 ( .A(x[1895]), .B(y[1895]), .Z(n23754) );
  NAND U12827 ( .A(n8031), .B(n23754), .Z(n8032) );
  NANDN U12828 ( .A(n23755), .B(n8032), .Z(n8033) );
  NANDN U12829 ( .A(n23757), .B(n8033), .Z(n8034) );
  NANDN U12830 ( .A(y[1897]), .B(x[1897]), .Z(n12243) );
  IV U12831 ( .A(y[1898]), .Z(n12241) );
  NAND U12832 ( .A(n12241), .B(x[1898]), .Z(n12240) );
  AND U12833 ( .A(n12243), .B(n12240), .Z(n23759) );
  NAND U12834 ( .A(n8034), .B(n23759), .Z(n8035) );
  ANDN U12835 ( .B(y[1899]), .A(x[1899]), .Z(n12239) );
  NAND U12836 ( .A(n8035), .B(n23761), .Z(n8036) );
  NANDN U12837 ( .A(y[1899]), .B(x[1899]), .Z(n23763) );
  AND U12838 ( .A(n8036), .B(n23763), .Z(n8037) );
  NANDN U12839 ( .A(n12238), .B(n8037), .Z(n8038) );
  NANDN U12840 ( .A(n23766), .B(n8038), .Z(n8039) );
  NAND U12841 ( .A(n8040), .B(n8039), .Z(n8041) );
  NAND U12842 ( .A(n15770), .B(n8041), .Z(n8042) );
  NAND U12843 ( .A(n8043), .B(n8042), .Z(n8044) );
  NAND U12844 ( .A(n8045), .B(n8044), .Z(n8046) );
  NANDN U12845 ( .A(y[1904]), .B(x[1904]), .Z(n23775) );
  AND U12846 ( .A(n8046), .B(n23775), .Z(n8047) );
  NANDN U12847 ( .A(n12236), .B(n8047), .Z(n8048) );
  ANDN U12848 ( .B(y[1904]), .A(x[1904]), .Z(n15774) );
  ANDN U12849 ( .B(y[1905]), .A(x[1905]), .Z(n15778) );
  NOR U12850 ( .A(n15774), .B(n15778), .Z(n23777) );
  NAND U12851 ( .A(n8048), .B(n23777), .Z(n8051) );
  NANDN U12852 ( .A(y[1906]), .B(x[1906]), .Z(n8050) );
  NANDN U12853 ( .A(y[1905]), .B(x[1905]), .Z(n8049) );
  AND U12854 ( .A(n8050), .B(n8049), .Z(n23779) );
  NAND U12855 ( .A(n8051), .B(n23779), .Z(n8053) );
  NANDN U12856 ( .A(x[1907]), .B(y[1907]), .Z(n8052) );
  NANDN U12857 ( .A(x[1906]), .B(y[1906]), .Z(n23782) );
  NAND U12858 ( .A(n8052), .B(n23782), .Z(n15781) );
  ANDN U12859 ( .B(n8053), .A(n15781), .Z(n8054) );
  ANDN U12860 ( .B(n15783), .A(n8054), .Z(n8057) );
  NANDN U12861 ( .A(x[1908]), .B(y[1908]), .Z(n8056) );
  NANDN U12862 ( .A(x[1909]), .B(y[1909]), .Z(n8055) );
  AND U12863 ( .A(n8056), .B(n8055), .Z(n23789) );
  NANDN U12864 ( .A(n8057), .B(n23789), .Z(n8058) );
  NANDN U12865 ( .A(n23792), .B(n8058), .Z(n8061) );
  NANDN U12866 ( .A(x[1910]), .B(y[1910]), .Z(n8060) );
  NANDN U12867 ( .A(x[1911]), .B(y[1911]), .Z(n8059) );
  AND U12868 ( .A(n8060), .B(n8059), .Z(n23793) );
  NAND U12869 ( .A(n8061), .B(n23793), .Z(n8062) );
  NANDN U12870 ( .A(n23796), .B(n8062), .Z(n8063) );
  ANDN U12871 ( .B(y[1913]), .A(x[1913]), .Z(n15794) );
  ANDN U12872 ( .B(y[1912]), .A(x[1912]), .Z(n15790) );
  NOR U12873 ( .A(n15794), .B(n15790), .Z(n23797) );
  NAND U12874 ( .A(n8063), .B(n23797), .Z(n8064) );
  AND U12875 ( .A(n23800), .B(n8064), .Z(n8065) );
  ANDN U12876 ( .B(x[1914]), .A(y[1914]), .Z(n12231) );
  ANDN U12877 ( .B(n8065), .A(n12231), .Z(n8067) );
  NANDN U12878 ( .A(x[1914]), .B(y[1914]), .Z(n8066) );
  ANDN U12879 ( .B(y[1915]), .A(x[1915]), .Z(n12232) );
  ANDN U12880 ( .B(n8066), .A(n12232), .Z(n23801) );
  NANDN U12881 ( .A(n8067), .B(n23801), .Z(n8068) );
  NANDN U12882 ( .A(n12234), .B(n8068), .Z(n8071) );
  NANDN U12883 ( .A(x[1916]), .B(y[1916]), .Z(n8070) );
  NANDN U12884 ( .A(x[1917]), .B(y[1917]), .Z(n8069) );
  AND U12885 ( .A(n8070), .B(n8069), .Z(n23805) );
  NAND U12886 ( .A(n8071), .B(n23805), .Z(n8074) );
  NANDN U12887 ( .A(y[1918]), .B(x[1918]), .Z(n8073) );
  NANDN U12888 ( .A(y[1917]), .B(x[1917]), .Z(n8072) );
  NAND U12889 ( .A(n8073), .B(n8072), .Z(n23808) );
  ANDN U12890 ( .B(n8074), .A(n23808), .Z(n8075) );
  NANDN U12891 ( .A(x[1918]), .B(y[1918]), .Z(n23811) );
  NANDN U12892 ( .A(n8075), .B(n23811), .Z(n8076) );
  NANDN U12893 ( .A(n23814), .B(n8076), .Z(n8077) );
  NANDN U12894 ( .A(n12229), .B(n8077), .Z(n8078) );
  OR U12895 ( .A(n15801), .B(n8078), .Z(n8079) );
  AND U12896 ( .A(n23818), .B(n8079), .Z(n8080) );
  OR U12897 ( .A(n12230), .B(n8080), .Z(n8083) );
  NANDN U12898 ( .A(y[1922]), .B(x[1922]), .Z(n8082) );
  NANDN U12899 ( .A(y[1923]), .B(x[1923]), .Z(n8081) );
  NAND U12900 ( .A(n8082), .B(n8081), .Z(n23822) );
  ANDN U12901 ( .B(n8083), .A(n23822), .Z(n8084) );
  OR U12902 ( .A(n15806), .B(n8084), .Z(n8086) );
  IV U12903 ( .A(y[1924]), .Z(n20264) );
  NAND U12904 ( .A(n20264), .B(x[1924]), .Z(n8085) );
  NANDN U12905 ( .A(y[1925]), .B(x[1925]), .Z(n23832) );
  NAND U12906 ( .A(n8085), .B(n23832), .Z(n15808) );
  ANDN U12907 ( .B(n8086), .A(n15808), .Z(n8087) );
  NANDN U12908 ( .A(x[1925]), .B(y[1925]), .Z(n23829) );
  NANDN U12909 ( .A(n8087), .B(n23829), .Z(n8088) );
  AND U12910 ( .A(n23833), .B(n8088), .Z(n8091) );
  NANDN U12911 ( .A(x[1927]), .B(y[1927]), .Z(n8090) );
  NANDN U12912 ( .A(x[1926]), .B(y[1926]), .Z(n8089) );
  AND U12913 ( .A(n8090), .B(n8089), .Z(n23835) );
  NANDN U12914 ( .A(n8091), .B(n23835), .Z(n8092) );
  ANDN U12915 ( .B(x[1928]), .A(y[1928]), .Z(n12228) );
  ANDN U12916 ( .B(n8092), .A(n12228), .Z(n8093) );
  NANDN U12917 ( .A(y[1927]), .B(x[1927]), .Z(n23838) );
  NAND U12918 ( .A(n8093), .B(n23838), .Z(n8094) );
  AND U12919 ( .A(n8095), .B(n8094), .Z(n8096) );
  AND U12920 ( .A(n8097), .B(n8096), .Z(n8110) );
  XNOR U12921 ( .A(x[1932]), .B(y[1932]), .Z(n8099) );
  NANDN U12922 ( .A(y[1931]), .B(x[1931]), .Z(n8098) );
  NAND U12923 ( .A(n8099), .B(n8098), .Z(n8103) );
  NANDN U12924 ( .A(y[1930]), .B(x[1930]), .Z(n8100) );
  NANDN U12925 ( .A(n8103), .B(n8100), .Z(n23846) );
  NANDN U12926 ( .A(y[1929]), .B(x[1929]), .Z(n12227) );
  NANDN U12927 ( .A(n23846), .B(n12227), .Z(n8106) );
  OR U12928 ( .A(n15819), .B(n8101), .Z(n8102) );
  NANDN U12929 ( .A(n8103), .B(n8102), .Z(n8105) );
  ANDN U12930 ( .B(n8105), .A(n8104), .Z(n23847) );
  NAND U12931 ( .A(n8106), .B(n23847), .Z(n8108) );
  NANDN U12932 ( .A(y[1934]), .B(x[1934]), .Z(n8107) );
  ANDN U12933 ( .B(x[1933]), .A(y[1933]), .Z(n15825) );
  ANDN U12934 ( .B(n8107), .A(n15825), .Z(n23850) );
  NAND U12935 ( .A(n8108), .B(n23850), .Z(n8109) );
  OR U12936 ( .A(n8110), .B(n8109), .Z(n8112) );
  NANDN U12937 ( .A(x[1935]), .B(y[1935]), .Z(n15830) );
  IV U12938 ( .A(x[1934]), .Z(n15831) );
  NAND U12939 ( .A(n15831), .B(y[1934]), .Z(n8111) );
  NAND U12940 ( .A(n15830), .B(n8111), .Z(n23852) );
  ANDN U12941 ( .B(n8112), .A(n23852), .Z(n8115) );
  NANDN U12942 ( .A(y[1935]), .B(x[1935]), .Z(n8114) );
  NANDN U12943 ( .A(y[1936]), .B(x[1936]), .Z(n8113) );
  AND U12944 ( .A(n8114), .B(n8113), .Z(n23854) );
  NANDN U12945 ( .A(n8115), .B(n23854), .Z(n8118) );
  NANDN U12946 ( .A(x[1937]), .B(y[1937]), .Z(n8117) );
  NANDN U12947 ( .A(x[1936]), .B(y[1936]), .Z(n8116) );
  AND U12948 ( .A(n8117), .B(n8116), .Z(n23855) );
  NAND U12949 ( .A(n8118), .B(n23855), .Z(n8121) );
  NANDN U12950 ( .A(y[1937]), .B(x[1937]), .Z(n8120) );
  NANDN U12951 ( .A(y[1938]), .B(x[1938]), .Z(n8119) );
  AND U12952 ( .A(n8120), .B(n8119), .Z(n23857) );
  NAND U12953 ( .A(n8121), .B(n23857), .Z(n8122) );
  AND U12954 ( .A(n23859), .B(n8122), .Z(n8125) );
  NANDN U12955 ( .A(y[1939]), .B(x[1939]), .Z(n8124) );
  NANDN U12956 ( .A(y[1940]), .B(x[1940]), .Z(n8123) );
  AND U12957 ( .A(n8124), .B(n8123), .Z(n23861) );
  NANDN U12958 ( .A(n8125), .B(n23861), .Z(n8128) );
  NANDN U12959 ( .A(x[1941]), .B(y[1941]), .Z(n8127) );
  NANDN U12960 ( .A(x[1940]), .B(y[1940]), .Z(n8126) );
  AND U12961 ( .A(n8127), .B(n8126), .Z(n23863) );
  NAND U12962 ( .A(n8128), .B(n23863), .Z(n8131) );
  NANDN U12963 ( .A(y[1941]), .B(x[1941]), .Z(n8130) );
  NANDN U12964 ( .A(y[1942]), .B(x[1942]), .Z(n8129) );
  AND U12965 ( .A(n8130), .B(n8129), .Z(n23866) );
  NAND U12966 ( .A(n8131), .B(n23866), .Z(n8132) );
  AND U12967 ( .A(n23867), .B(n8132), .Z(n8135) );
  NANDN U12968 ( .A(y[1943]), .B(x[1943]), .Z(n8134) );
  NANDN U12969 ( .A(y[1944]), .B(x[1944]), .Z(n8133) );
  AND U12970 ( .A(n8134), .B(n8133), .Z(n23870) );
  NANDN U12971 ( .A(n8135), .B(n23870), .Z(n8138) );
  NANDN U12972 ( .A(x[1945]), .B(y[1945]), .Z(n8137) );
  NANDN U12973 ( .A(x[1944]), .B(y[1944]), .Z(n8136) );
  AND U12974 ( .A(n8137), .B(n8136), .Z(n23871) );
  NAND U12975 ( .A(n8138), .B(n23871), .Z(n8141) );
  NANDN U12976 ( .A(y[1945]), .B(x[1945]), .Z(n8140) );
  NANDN U12977 ( .A(y[1946]), .B(x[1946]), .Z(n8139) );
  AND U12978 ( .A(n8140), .B(n8139), .Z(n23874) );
  NAND U12979 ( .A(n8141), .B(n23874), .Z(n8142) );
  AND U12980 ( .A(n23875), .B(n8142), .Z(n8143) );
  OR U12981 ( .A(n23878), .B(n8143), .Z(n8144) );
  NANDN U12982 ( .A(x[1948]), .B(y[1948]), .Z(n23879) );
  ANDN U12983 ( .B(y[1949]), .A(x[1949]), .Z(n23885) );
  ANDN U12984 ( .B(n23879), .A(n23885), .Z(n15849) );
  NAND U12985 ( .A(n8144), .B(n15849), .Z(n8145) );
  AND U12986 ( .A(n23881), .B(n8145), .Z(n8146) );
  NANDN U12987 ( .A(x[1951]), .B(y[1951]), .Z(n12226) );
  NANDN U12988 ( .A(x[1950]), .B(y[1950]), .Z(n15853) );
  AND U12989 ( .A(n12226), .B(n15853), .Z(n23883) );
  NANDN U12990 ( .A(n8146), .B(n23883), .Z(n8147) );
  AND U12991 ( .A(n23890), .B(n8147), .Z(n8150) );
  NANDN U12992 ( .A(x[1952]), .B(y[1952]), .Z(n8149) );
  NANDN U12993 ( .A(x[1953]), .B(y[1953]), .Z(n8148) );
  AND U12994 ( .A(n8149), .B(n8148), .Z(n23891) );
  NANDN U12995 ( .A(n8150), .B(n23891), .Z(n8153) );
  NANDN U12996 ( .A(y[1954]), .B(x[1954]), .Z(n8152) );
  NANDN U12997 ( .A(y[1953]), .B(x[1953]), .Z(n8151) );
  NAND U12998 ( .A(n8152), .B(n8151), .Z(n23894) );
  ANDN U12999 ( .B(n8153), .A(n23894), .Z(n8156) );
  NANDN U13000 ( .A(x[1955]), .B(y[1955]), .Z(n8155) );
  NANDN U13001 ( .A(x[1954]), .B(y[1954]), .Z(n8154) );
  AND U13002 ( .A(n8155), .B(n8154), .Z(n23895) );
  NANDN U13003 ( .A(n8156), .B(n23895), .Z(n8157) );
  ANDN U13004 ( .B(x[1956]), .A(y[1956]), .Z(n12221) );
  ANDN U13005 ( .B(n8157), .A(n12221), .Z(n8158) );
  NANDN U13006 ( .A(y[1955]), .B(x[1955]), .Z(n23897) );
  NAND U13007 ( .A(n8158), .B(n23897), .Z(n8160) );
  NANDN U13008 ( .A(x[1956]), .B(y[1956]), .Z(n8159) );
  ANDN U13009 ( .B(y[1957]), .A(x[1957]), .Z(n12222) );
  ANDN U13010 ( .B(n8159), .A(n12222), .Z(n23899) );
  NAND U13011 ( .A(n8160), .B(n23899), .Z(n8161) );
  NANDN U13012 ( .A(n12224), .B(n8161), .Z(n8162) );
  ANDN U13013 ( .B(y[1959]), .A(x[1959]), .Z(n15869) );
  NANDN U13014 ( .A(x[1958]), .B(y[1958]), .Z(n15866) );
  NANDN U13015 ( .A(n15869), .B(n15866), .Z(n23906) );
  ANDN U13016 ( .B(n8162), .A(n23906), .Z(n8164) );
  NANDN U13017 ( .A(y[1959]), .B(x[1959]), .Z(n23911) );
  NANDN U13018 ( .A(y[1958]), .B(x[1958]), .Z(n23901) );
  AND U13019 ( .A(n23911), .B(n23901), .Z(n15867) );
  OR U13020 ( .A(n15869), .B(n15867), .Z(n8163) );
  NANDN U13021 ( .A(n8164), .B(n8163), .Z(n8165) );
  IV U13022 ( .A(y[1960]), .Z(n12220) );
  NANDN U13023 ( .A(n8165), .B(n15872), .Z(n8166) );
  NANDN U13024 ( .A(n23913), .B(n8166), .Z(n8169) );
  NANDN U13025 ( .A(y[1963]), .B(x[1963]), .Z(n8168) );
  NANDN U13026 ( .A(y[1964]), .B(x[1964]), .Z(n8167) );
  AND U13027 ( .A(n8168), .B(n8167), .Z(n23915) );
  NAND U13028 ( .A(n8169), .B(n23915), .Z(n8172) );
  NANDN U13029 ( .A(x[1965]), .B(y[1965]), .Z(n8171) );
  NANDN U13030 ( .A(x[1964]), .B(y[1964]), .Z(n8170) );
  NAND U13031 ( .A(n8171), .B(n8170), .Z(n23918) );
  ANDN U13032 ( .B(n8172), .A(n23918), .Z(n8175) );
  NANDN U13033 ( .A(y[1965]), .B(x[1965]), .Z(n8174) );
  NANDN U13034 ( .A(y[1966]), .B(x[1966]), .Z(n8173) );
  AND U13035 ( .A(n8174), .B(n8173), .Z(n23919) );
  NANDN U13036 ( .A(n8175), .B(n23919), .Z(n8176) );
  NANDN U13037 ( .A(n23922), .B(n8176), .Z(n8179) );
  NANDN U13038 ( .A(y[1967]), .B(x[1967]), .Z(n8178) );
  NANDN U13039 ( .A(y[1968]), .B(x[1968]), .Z(n8177) );
  AND U13040 ( .A(n8178), .B(n8177), .Z(n23923) );
  NAND U13041 ( .A(n8179), .B(n23923), .Z(n8180) );
  NANDN U13042 ( .A(n23925), .B(n8180), .Z(n8181) );
  ANDN U13043 ( .B(x[1970]), .A(y[1970]), .Z(n12219) );
  ANDN U13044 ( .B(n8181), .A(n12219), .Z(n8182) );
  NANDN U13045 ( .A(y[1969]), .B(x[1969]), .Z(n23927) );
  NAND U13046 ( .A(n8182), .B(n23927), .Z(n8183) );
  AND U13047 ( .A(n23929), .B(n8183), .Z(n8184) );
  NAND U13048 ( .A(n8185), .B(n8184), .Z(n8186) );
  NAND U13049 ( .A(n8187), .B(n8186), .Z(n8189) );
  NANDN U13050 ( .A(x[1972]), .B(y[1972]), .Z(n15889) );
  OR U13051 ( .A(n23940), .B(n15889), .Z(n8188) );
  AND U13052 ( .A(n8189), .B(n8188), .Z(n8190) );
  NANDN U13053 ( .A(n15895), .B(n8190), .Z(n8191) );
  AND U13054 ( .A(n15896), .B(n8191), .Z(n8194) );
  NANDN U13055 ( .A(x[1975]), .B(y[1975]), .Z(n8193) );
  NANDN U13056 ( .A(x[1976]), .B(y[1976]), .Z(n8192) );
  AND U13057 ( .A(n8193), .B(n8192), .Z(n23948) );
  NANDN U13058 ( .A(n8194), .B(n23948), .Z(n8195) );
  NANDN U13059 ( .A(n23950), .B(n8195), .Z(n8198) );
  NANDN U13060 ( .A(x[1978]), .B(y[1978]), .Z(n8197) );
  NANDN U13061 ( .A(x[1977]), .B(y[1977]), .Z(n8196) );
  AND U13062 ( .A(n8197), .B(n8196), .Z(n23951) );
  NAND U13063 ( .A(n8198), .B(n23951), .Z(n8199) );
  AND U13064 ( .A(n23954), .B(n8199), .Z(n8200) );
  NANDN U13065 ( .A(x[1979]), .B(y[1979]), .Z(n23955) );
  NANDN U13066 ( .A(n8200), .B(n23955), .Z(n8201) );
  NANDN U13067 ( .A(n23958), .B(n8201), .Z(n8202) );
  NANDN U13068 ( .A(x[1981]), .B(y[1981]), .Z(n12216) );
  ANDN U13069 ( .B(y[1980]), .A(x[1980]), .Z(n15904) );
  ANDN U13070 ( .B(n12216), .A(n15904), .Z(n23959) );
  NAND U13071 ( .A(n8202), .B(n23959), .Z(n8204) );
  NANDN U13072 ( .A(y[1981]), .B(x[1981]), .Z(n8203) );
  NANDN U13073 ( .A(y[1982]), .B(x[1982]), .Z(n12215) );
  NAND U13074 ( .A(n8203), .B(n12215), .Z(n23962) );
  ANDN U13075 ( .B(n8204), .A(n23962), .Z(n8205) );
  OR U13076 ( .A(n23964), .B(n8205), .Z(n8206) );
  AND U13077 ( .A(n8207), .B(n8206), .Z(n8208) );
  NANDN U13078 ( .A(x[1984]), .B(y[1984]), .Z(n23967) );
  NANDN U13079 ( .A(n8208), .B(n23967), .Z(n8209) );
  NANDN U13080 ( .A(n12214), .B(n8209), .Z(n8212) );
  NANDN U13081 ( .A(x[1986]), .B(y[1986]), .Z(n8211) );
  NANDN U13082 ( .A(x[1985]), .B(y[1985]), .Z(n8210) );
  AND U13083 ( .A(n8211), .B(n8210), .Z(n23971) );
  NAND U13084 ( .A(n8212), .B(n23971), .Z(n8213) );
  AND U13085 ( .A(n23973), .B(n8213), .Z(n8214) );
  XNOR U13086 ( .A(y[1987]), .B(x[1987]), .Z(n23976) );
  NANDN U13087 ( .A(n8214), .B(n23976), .Z(n8215) );
  NANDN U13088 ( .A(n23978), .B(n8215), .Z(n8218) );
  NANDN U13089 ( .A(x[1988]), .B(y[1988]), .Z(n8217) );
  NANDN U13090 ( .A(x[1989]), .B(y[1989]), .Z(n8216) );
  AND U13091 ( .A(n8217), .B(n8216), .Z(n23980) );
  NAND U13092 ( .A(n8218), .B(n23980), .Z(n8219) );
  NANDN U13093 ( .A(y[1989]), .B(x[1989]), .Z(n23982) );
  NAND U13094 ( .A(n8219), .B(n23982), .Z(n8220) );
  NANDN U13095 ( .A(x[1990]), .B(y[1990]), .Z(n23985) );
  NAND U13096 ( .A(n8220), .B(n23985), .Z(n8221) );
  ANDN U13097 ( .B(x[1990]), .A(y[1990]), .Z(n23981) );
  NANDN U13098 ( .A(y[1991]), .B(x[1991]), .Z(n23987) );
  NANDN U13099 ( .A(n23981), .B(n23987), .Z(n15927) );
  ANDN U13100 ( .B(n8221), .A(n15927), .Z(n8222) );
  OR U13101 ( .A(n12211), .B(n8222), .Z(n8223) );
  NANDN U13102 ( .A(y[1992]), .B(x[1992]), .Z(n23992) );
  NAND U13103 ( .A(n8223), .B(n23992), .Z(n8224) );
  NANDN U13104 ( .A(x[1993]), .B(y[1993]), .Z(n23993) );
  NAND U13105 ( .A(n8224), .B(n23993), .Z(n8225) );
  OR U13106 ( .A(n12212), .B(n8225), .Z(n8226) );
  NANDN U13107 ( .A(n23996), .B(n8226), .Z(n8227) );
  NANDN U13108 ( .A(n23998), .B(n8227), .Z(n8228) );
  ANDN U13109 ( .B(x[1996]), .A(y[1996]), .Z(n12206) );
  NAND U13110 ( .A(n8228), .B(n23999), .Z(n8229) );
  AND U13111 ( .A(n24001), .B(n8229), .Z(n8231) );
  NANDN U13112 ( .A(y[1997]), .B(x[1997]), .Z(n24004) );
  ANDN U13113 ( .B(x[1998]), .A(y[1998]), .Z(n15946) );
  ANDN U13114 ( .B(n24004), .A(n15946), .Z(n8230) );
  NANDN U13115 ( .A(n8231), .B(n8230), .Z(n8232) );
  AND U13116 ( .A(n24005), .B(n8232), .Z(n8233) );
  NAND U13117 ( .A(n8234), .B(n8233), .Z(n8235) );
  NAND U13118 ( .A(n8236), .B(n8235), .Z(n8237) );
  ANDN U13119 ( .B(y[2000]), .A(x[2000]), .Z(n12205) );
  ANDN U13120 ( .B(n8237), .A(n12205), .Z(n8238) );
  NANDN U13121 ( .A(n15952), .B(n8238), .Z(n8239) );
  NANDN U13122 ( .A(n15950), .B(n8239), .Z(n8240) );
  NANDN U13123 ( .A(n15954), .B(n8240), .Z(n8242) );
  IV U13124 ( .A(y[2004]), .Z(n15960) );
  NAND U13125 ( .A(n15960), .B(x[2004]), .Z(n8241) );
  NANDN U13126 ( .A(y[2003]), .B(x[2003]), .Z(n15958) );
  NAND U13127 ( .A(n8241), .B(n15958), .Z(n24015) );
  ANDN U13128 ( .B(n8242), .A(n24015), .Z(n8244) );
  NANDN U13129 ( .A(x[2004]), .B(y[2004]), .Z(n8243) );
  NANDN U13130 ( .A(x[2005]), .B(y[2005]), .Z(n15965) );
  NAND U13131 ( .A(n8243), .B(n15965), .Z(n24018) );
  OR U13132 ( .A(n8244), .B(n24018), .Z(n8247) );
  NANDN U13133 ( .A(y[2005]), .B(x[2005]), .Z(n8246) );
  NANDN U13134 ( .A(y[2006]), .B(x[2006]), .Z(n8245) );
  AND U13135 ( .A(n8246), .B(n8245), .Z(n24020) );
  NAND U13136 ( .A(n8247), .B(n24020), .Z(n8248) );
  AND U13137 ( .A(n24021), .B(n8248), .Z(n8251) );
  NANDN U13138 ( .A(y[2007]), .B(x[2007]), .Z(n8250) );
  NANDN U13139 ( .A(y[2008]), .B(x[2008]), .Z(n8249) );
  AND U13140 ( .A(n8250), .B(n8249), .Z(n24023) );
  NANDN U13141 ( .A(n8251), .B(n24023), .Z(n8252) );
  AND U13142 ( .A(n24025), .B(n8252), .Z(n8255) );
  NANDN U13143 ( .A(y[2009]), .B(x[2009]), .Z(n8254) );
  NANDN U13144 ( .A(y[2010]), .B(x[2010]), .Z(n8253) );
  AND U13145 ( .A(n8254), .B(n8253), .Z(n24027) );
  NANDN U13146 ( .A(n8255), .B(n24027), .Z(n8256) );
  AND U13147 ( .A(n24029), .B(n8256), .Z(n8258) );
  NANDN U13148 ( .A(y[2012]), .B(x[2012]), .Z(n8257) );
  ANDN U13149 ( .B(x[2011]), .A(y[2011]), .Z(n24031) );
  ANDN U13150 ( .B(n8257), .A(n24031), .Z(n15972) );
  NANDN U13151 ( .A(n8258), .B(n15972), .Z(n8259) );
  NANDN U13152 ( .A(x[2013]), .B(y[2013]), .Z(n24039) );
  NANDN U13153 ( .A(x[2012]), .B(y[2012]), .Z(n24036) );
  AND U13154 ( .A(n24039), .B(n24036), .Z(n15974) );
  NAND U13155 ( .A(n8259), .B(n15974), .Z(n8262) );
  ANDN U13156 ( .B(x[2013]), .A(y[2013]), .Z(n24037) );
  NANDN U13157 ( .A(y[2014]), .B(x[2014]), .Z(n8260) );
  NAND U13158 ( .A(n8261), .B(n8260), .Z(n24041) );
  NOR U13159 ( .A(n24037), .B(n24041), .Z(n15977) );
  NAND U13160 ( .A(n8262), .B(n15977), .Z(n8263) );
  AND U13161 ( .A(n24043), .B(n8263), .Z(n8268) );
  NANDN U13162 ( .A(y[2016]), .B(x[2016]), .Z(n8264) );
  NANDN U13163 ( .A(n8264), .B(x[2017]), .Z(n8267) );
  XNOR U13164 ( .A(n8264), .B(x[2017]), .Z(n8265) );
  NANDN U13165 ( .A(y[2017]), .B(n8265), .Z(n8266) );
  AND U13166 ( .A(n8267), .B(n8266), .Z(n24046) );
  NANDN U13167 ( .A(n8268), .B(n24046), .Z(n8269) );
  AND U13168 ( .A(n24050), .B(n8269), .Z(n8271) );
  NANDN U13169 ( .A(y[2018]), .B(x[2018]), .Z(n8270) );
  ANDN U13170 ( .B(x[2019]), .A(y[2019]), .Z(n24051) );
  ANDN U13171 ( .B(n8270), .A(n24051), .Z(n15981) );
  NANDN U13172 ( .A(n8271), .B(n15981), .Z(n8272) );
  NANDN U13173 ( .A(n12202), .B(n8272), .Z(n8273) );
  NANDN U13174 ( .A(n24055), .B(n8273), .Z(n8274) );
  ANDN U13175 ( .B(y[2020]), .A(x[2020]), .Z(n12203) );
  ANDN U13176 ( .B(n8274), .A(n12203), .Z(n8275) );
  NANDN U13177 ( .A(x[2021]), .B(y[2021]), .Z(n24058) );
  NAND U13178 ( .A(n8275), .B(n24058), .Z(n8276) );
  XNOR U13179 ( .A(x[2022]), .B(y[2022]), .Z(n15988) );
  ANDN U13180 ( .B(x[2021]), .A(y[2021]), .Z(n12201) );
  ANDN U13181 ( .B(n15988), .A(n12201), .Z(n24059) );
  NAND U13182 ( .A(n8276), .B(n24059), .Z(n8279) );
  NANDN U13183 ( .A(x[2022]), .B(y[2022]), .Z(n8278) );
  NANDN U13184 ( .A(x[2023]), .B(y[2023]), .Z(n8277) );
  NAND U13185 ( .A(n8278), .B(n8277), .Z(n24062) );
  ANDN U13186 ( .B(n8279), .A(n24062), .Z(n8282) );
  NANDN U13187 ( .A(y[2023]), .B(x[2023]), .Z(n8281) );
  NANDN U13188 ( .A(y[2024]), .B(x[2024]), .Z(n8280) );
  AND U13189 ( .A(n8281), .B(n8280), .Z(n24063) );
  NANDN U13190 ( .A(n8282), .B(n24063), .Z(n8285) );
  NANDN U13191 ( .A(x[2024]), .B(y[2024]), .Z(n8284) );
  NANDN U13192 ( .A(x[2025]), .B(y[2025]), .Z(n8283) );
  NAND U13193 ( .A(n8284), .B(n8283), .Z(n24066) );
  ANDN U13194 ( .B(n8285), .A(n24066), .Z(n8287) );
  NANDN U13195 ( .A(y[2025]), .B(x[2025]), .Z(n24067) );
  ANDN U13196 ( .B(x[2026]), .A(y[2026]), .Z(n12199) );
  ANDN U13197 ( .B(n24067), .A(n12199), .Z(n8286) );
  NANDN U13198 ( .A(n8287), .B(n8286), .Z(n8288) );
  NANDN U13199 ( .A(x[2027]), .B(y[2027]), .Z(n24074) );
  NAND U13200 ( .A(n8288), .B(n24074), .Z(n8289) );
  NANDN U13201 ( .A(x[2026]), .B(y[2026]), .Z(n24070) );
  NANDN U13202 ( .A(n8289), .B(n24070), .Z(n8290) );
  AND U13203 ( .A(n8291), .B(n8290), .Z(n8292) );
  ANDN U13204 ( .B(y[2029]), .A(x[2029]), .Z(n16002) );
  ANDN U13205 ( .B(y[2028]), .A(x[2028]), .Z(n15995) );
  NOR U13206 ( .A(n16002), .B(n15995), .Z(n24077) );
  NANDN U13207 ( .A(n8292), .B(n24077), .Z(n8293) );
  NANDN U13208 ( .A(n24079), .B(n8293), .Z(n8294) );
  NANDN U13209 ( .A(n24082), .B(n8294), .Z(n8296) );
  NANDN U13210 ( .A(y[2031]), .B(x[2031]), .Z(n8295) );
  ANDN U13211 ( .B(x[2032]), .A(y[2032]), .Z(n12198) );
  ANDN U13212 ( .B(n8295), .A(n12198), .Z(n24083) );
  NAND U13213 ( .A(n8296), .B(n24083), .Z(n8297) );
  ANDN U13214 ( .B(y[2033]), .A(x[2033]), .Z(n16016) );
  ANDN U13215 ( .B(y[2032]), .A(x[2032]), .Z(n16012) );
  NOR U13216 ( .A(n16016), .B(n16012), .Z(n24085) );
  NAND U13217 ( .A(n8297), .B(n24085), .Z(n8298) );
  ANDN U13218 ( .B(x[2033]), .A(y[2033]), .Z(n24087) );
  ANDN U13219 ( .B(n8298), .A(n24087), .Z(n8299) );
  NANDN U13220 ( .A(n12196), .B(n8299), .Z(n8301) );
  NANDN U13221 ( .A(x[2035]), .B(y[2035]), .Z(n24093) );
  NANDN U13222 ( .A(x[2034]), .B(y[2034]), .Z(n24089) );
  AND U13223 ( .A(n24093), .B(n24089), .Z(n8300) );
  NAND U13224 ( .A(n8301), .B(n8300), .Z(n8302) );
  NANDN U13225 ( .A(y[2036]), .B(x[2036]), .Z(n24095) );
  ANDN U13226 ( .B(y[2039]), .A(x[2039]), .Z(n12191) );
  NANDN U13227 ( .A(y[2039]), .B(x[2039]), .Z(n24103) );
  NANDN U13228 ( .A(x[2040]), .B(y[2040]), .Z(n8305) );
  NANDN U13229 ( .A(x[2041]), .B(y[2041]), .Z(n8304) );
  NAND U13230 ( .A(n8304), .B(n8303), .Z(n16038) );
  ANDN U13231 ( .B(n8305), .A(n16038), .Z(n24105) );
  ANDN U13232 ( .B(x[2044]), .A(y[2044]), .Z(n16045) );
  NANDN U13233 ( .A(y[2043]), .B(x[2043]), .Z(n16033) );
  NANDN U13234 ( .A(n16045), .B(n16033), .Z(n8306) );
  NANDN U13235 ( .A(n8307), .B(n8306), .Z(n8310) );
  NANDN U13236 ( .A(y[2045]), .B(x[2045]), .Z(n8309) );
  NANDN U13237 ( .A(y[2046]), .B(x[2046]), .Z(n8308) );
  NAND U13238 ( .A(n8309), .B(n8308), .Z(n16044) );
  ANDN U13239 ( .B(n8310), .A(n16044), .Z(n24112) );
  NANDN U13240 ( .A(y[2047]), .B(x[2047]), .Z(n8312) );
  NANDN U13241 ( .A(y[2048]), .B(x[2048]), .Z(n8311) );
  AND U13242 ( .A(n8312), .B(n8311), .Z(n24115) );
  NANDN U13243 ( .A(x[2050]), .B(y[2050]), .Z(n8314) );
  NANDN U13244 ( .A(x[2051]), .B(y[2051]), .Z(n8313) );
  AND U13245 ( .A(n8314), .B(n8313), .Z(n24121) );
  NANDN U13246 ( .A(y[2052]), .B(x[2052]), .Z(n8316) );
  NANDN U13247 ( .A(y[2051]), .B(x[2051]), .Z(n8315) );
  NAND U13248 ( .A(n8316), .B(n8315), .Z(n24123) );
  NANDN U13249 ( .A(x[2053]), .B(y[2053]), .Z(n8318) );
  NANDN U13250 ( .A(x[2052]), .B(y[2052]), .Z(n8317) );
  AND U13251 ( .A(n8318), .B(n8317), .Z(n24125) );
  NANDN U13252 ( .A(n8319), .B(n24125), .Z(n8320) );
  AND U13253 ( .A(n24128), .B(n8320), .Z(n8321) );
  ANDN U13254 ( .B(x[2054]), .A(y[2054]), .Z(n16059) );
  ANDN U13255 ( .B(n8321), .A(n16059), .Z(n8322) );
  ANDN U13256 ( .B(n24129), .A(n8322), .Z(n8323) );
  IV U13257 ( .A(x[2055]), .Z(n16061) );
  NANDN U13258 ( .A(n8323), .B(n16061), .Z(n8326) );
  XOR U13259 ( .A(x[2055]), .B(n8323), .Z(n8324) );
  NAND U13260 ( .A(n8324), .B(y[2055]), .Z(n8325) );
  NAND U13261 ( .A(n8326), .B(n8325), .Z(n8327) );
  ANDN U13262 ( .B(x[2056]), .A(y[2056]), .Z(n16066) );
  ANDN U13263 ( .B(n8327), .A(n16066), .Z(n8329) );
  NANDN U13264 ( .A(x[2056]), .B(y[2056]), .Z(n8328) );
  ANDN U13265 ( .B(y[2057]), .A(x[2057]), .Z(n16065) );
  ANDN U13266 ( .B(n8328), .A(n16065), .Z(n16062) );
  NANDN U13267 ( .A(n8329), .B(n16062), .Z(n8330) );
  NANDN U13268 ( .A(n24135), .B(n8330), .Z(n8331) );
  NANDN U13269 ( .A(n24140), .B(n8331), .Z(n8332) );
  NANDN U13270 ( .A(n24141), .B(n8332), .Z(n8333) );
  AND U13271 ( .A(n8334), .B(n8333), .Z(n8336) );
  NANDN U13272 ( .A(y[2062]), .B(x[2062]), .Z(n24149) );
  NANDN U13273 ( .A(y[2061]), .B(x[2061]), .Z(n24145) );
  AND U13274 ( .A(n24149), .B(n24145), .Z(n8335) );
  NANDN U13275 ( .A(n8336), .B(n8335), .Z(n8337) );
  AND U13276 ( .A(n24151), .B(n8337), .Z(n8338) );
  NANDN U13277 ( .A(n12187), .B(n8338), .Z(n8339) );
  ANDN U13278 ( .B(x[2063]), .A(y[2063]), .Z(n12185) );
  NAND U13279 ( .A(n8339), .B(n24154), .Z(n8340) );
  AND U13280 ( .A(n24155), .B(n8340), .Z(n8341) );
  OR U13281 ( .A(n24158), .B(n8341), .Z(n8343) );
  NANDN U13282 ( .A(x[2066]), .B(y[2066]), .Z(n8342) );
  ANDN U13283 ( .B(y[2067]), .A(x[2067]), .Z(n16096) );
  ANDN U13284 ( .B(n8342), .A(n16096), .Z(n24159) );
  NAND U13285 ( .A(n8343), .B(n24159), .Z(n8344) );
  NANDN U13286 ( .A(n24162), .B(n8344), .Z(n8345) );
  OR U13287 ( .A(n12182), .B(n8345), .Z(n8346) );
  AND U13288 ( .A(n24163), .B(n8346), .Z(n8347) );
  OR U13289 ( .A(n12183), .B(n8347), .Z(n8350) );
  NANDN U13290 ( .A(x[2069]), .B(y[2069]), .Z(n8349) );
  NANDN U13291 ( .A(x[2070]), .B(y[2070]), .Z(n8348) );
  NAND U13292 ( .A(n8349), .B(n8348), .Z(n24168) );
  ANDN U13293 ( .B(n8350), .A(n24168), .Z(n8351) );
  NANDN U13294 ( .A(y[2070]), .B(x[2070]), .Z(n24169) );
  NANDN U13295 ( .A(n8351), .B(n24169), .Z(n8352) );
  NANDN U13296 ( .A(x[2071]), .B(y[2071]), .Z(n24172) );
  NAND U13297 ( .A(n8352), .B(n24172), .Z(n8353) );
  NANDN U13298 ( .A(y[2071]), .B(x[2071]), .Z(n16103) );
  XOR U13299 ( .A(x[2072]), .B(y[2072]), .Z(n16106) );
  ANDN U13300 ( .B(n16103), .A(n16106), .Z(n24173) );
  NAND U13301 ( .A(n8353), .B(n24173), .Z(n8356) );
  NANDN U13302 ( .A(x[2072]), .B(y[2072]), .Z(n8355) );
  NANDN U13303 ( .A(x[2073]), .B(y[2073]), .Z(n8354) );
  NAND U13304 ( .A(n8355), .B(n8354), .Z(n24176) );
  ANDN U13305 ( .B(n8356), .A(n24176), .Z(n8357) );
  ANDN U13306 ( .B(n24179), .A(n8357), .Z(n8358) );
  OR U13307 ( .A(n24181), .B(n8358), .Z(n8363) );
  NANDN U13308 ( .A(y[2074]), .B(x[2074]), .Z(n24177) );
  NANDN U13309 ( .A(n24177), .B(n8359), .Z(n8362) );
  NANDN U13310 ( .A(y[2076]), .B(x[2076]), .Z(n8361) );
  NANDN U13311 ( .A(y[2075]), .B(x[2075]), .Z(n8360) );
  AND U13312 ( .A(n8361), .B(n8360), .Z(n24183) );
  AND U13313 ( .A(n8362), .B(n24183), .Z(n16111) );
  NAND U13314 ( .A(n8363), .B(n16111), .Z(n8366) );
  NANDN U13315 ( .A(x[2076]), .B(y[2076]), .Z(n8365) );
  NANDN U13316 ( .A(x[2077]), .B(y[2077]), .Z(n8364) );
  AND U13317 ( .A(n8365), .B(n8364), .Z(n24185) );
  NAND U13318 ( .A(n8366), .B(n24185), .Z(n8369) );
  NANDN U13319 ( .A(y[2077]), .B(x[2077]), .Z(n8368) );
  NANDN U13320 ( .A(y[2078]), .B(x[2078]), .Z(n8367) );
  AND U13321 ( .A(n8368), .B(n8367), .Z(n24187) );
  NAND U13322 ( .A(n8369), .B(n24187), .Z(n8370) );
  AND U13323 ( .A(n24189), .B(n8370), .Z(n8371) );
  OR U13324 ( .A(n24191), .B(n8371), .Z(n8372) );
  AND U13325 ( .A(n24193), .B(n8372), .Z(n8374) );
  NANDN U13326 ( .A(y[2081]), .B(x[2081]), .Z(n24195) );
  ANDN U13327 ( .B(x[2082]), .A(y[2082]), .Z(n12180) );
  ANDN U13328 ( .B(n24195), .A(n12180), .Z(n8373) );
  NANDN U13329 ( .A(n8374), .B(n8373), .Z(n8375) );
  AND U13330 ( .A(n24198), .B(n8375), .Z(n8376) );
  NAND U13331 ( .A(n8377), .B(n8376), .Z(n8378) );
  NAND U13332 ( .A(n8379), .B(n8378), .Z(n8380) );
  AND U13333 ( .A(n24205), .B(n8380), .Z(n8381) );
  NANDN U13334 ( .A(n12178), .B(n8381), .Z(n8383) );
  XNOR U13335 ( .A(y[2086]), .B(x[2086]), .Z(n8382) );
  ANDN U13336 ( .B(x[2085]), .A(y[2085]), .Z(n16132) );
  ANDN U13337 ( .B(n8382), .A(n16132), .Z(n24207) );
  NAND U13338 ( .A(n8383), .B(n24207), .Z(n8384) );
  NANDN U13339 ( .A(x[2087]), .B(y[2087]), .Z(n12176) );
  NANDN U13340 ( .A(x[2086]), .B(y[2086]), .Z(n16134) );
  NAND U13341 ( .A(n12176), .B(n16134), .Z(n24209) );
  ANDN U13342 ( .B(n8384), .A(n24209), .Z(n8385) );
  OR U13343 ( .A(n24211), .B(n8385), .Z(n8386) );
  AND U13344 ( .A(n24214), .B(n8386), .Z(n8387) );
  ANDN U13345 ( .B(y[2089]), .A(x[2089]), .Z(n16145) );
  ANDN U13346 ( .B(n8387), .A(n16145), .Z(n8389) );
  NANDN U13347 ( .A(y[2089]), .B(x[2089]), .Z(n8388) );
  ANDN U13348 ( .B(x[2090]), .A(y[2090]), .Z(n16146) );
  ANDN U13349 ( .B(n8388), .A(n16146), .Z(n24215) );
  NANDN U13350 ( .A(n8389), .B(n24215), .Z(n8390) );
  NANDN U13351 ( .A(n16148), .B(n8390), .Z(n8391) );
  NANDN U13352 ( .A(y[2091]), .B(x[2091]), .Z(n16150) );
  ANDN U13353 ( .B(x[2092]), .A(y[2092]), .Z(n12172) );
  ANDN U13354 ( .B(n16150), .A(n12172), .Z(n24219) );
  NAND U13355 ( .A(n8391), .B(n24219), .Z(n8394) );
  NANDN U13356 ( .A(x[2093]), .B(y[2093]), .Z(n8393) );
  NANDN U13357 ( .A(x[2092]), .B(y[2092]), .Z(n8392) );
  NAND U13358 ( .A(n8393), .B(n8392), .Z(n24222) );
  ANDN U13359 ( .B(n8394), .A(n24222), .Z(n8396) );
  NANDN U13360 ( .A(y[2093]), .B(x[2093]), .Z(n8395) );
  ANDN U13361 ( .B(x[2094]), .A(y[2094]), .Z(n12169) );
  ANDN U13362 ( .B(n8395), .A(n12169), .Z(n24223) );
  NANDN U13363 ( .A(n8396), .B(n24223), .Z(n8398) );
  NANDN U13364 ( .A(x[2094]), .B(y[2094]), .Z(n8397) );
  ANDN U13365 ( .B(y[2095]), .A(x[2095]), .Z(n12170) );
  ANDN U13366 ( .B(n8397), .A(n12170), .Z(n24225) );
  NAND U13367 ( .A(n8398), .B(n24225), .Z(n8399) );
  ANDN U13368 ( .B(x[2095]), .A(y[2095]), .Z(n20261) );
  ANDN U13369 ( .B(n8399), .A(n20261), .Z(n8400) );
  OR U13370 ( .A(n8400), .B(y[2096]), .Z(n8403) );
  XOR U13371 ( .A(y[2096]), .B(n8400), .Z(n8401) );
  NAND U13372 ( .A(x[2096]), .B(n8401), .Z(n8402) );
  NAND U13373 ( .A(n8403), .B(n8402), .Z(n8404) );
  AND U13374 ( .A(n20259), .B(n8404), .Z(n8406) );
  IV U13375 ( .A(y[2098]), .Z(n12166) );
  NAND U13376 ( .A(n12166), .B(x[2098]), .Z(n8405) );
  ANDN U13377 ( .B(x[2097]), .A(y[2097]), .Z(n12168) );
  ANDN U13378 ( .B(n8405), .A(n12168), .Z(n24232) );
  NANDN U13379 ( .A(n8406), .B(n24232), .Z(n8407) );
  IV U13380 ( .A(x[2098]), .Z(n12167) );
  NAND U13381 ( .A(y[2098]), .B(n12167), .Z(n16165) );
  IV U13382 ( .A(x[2099]), .Z(n12165) );
  NAND U13383 ( .A(n12165), .B(y[2099]), .Z(n12163) );
  AND U13384 ( .A(n16165), .B(n12163), .Z(n24233) );
  NAND U13385 ( .A(n8407), .B(n24233), .Z(n8408) );
  NANDN U13386 ( .A(n24236), .B(n8408), .Z(n8409) );
  NANDN U13387 ( .A(x[2100]), .B(y[2100]), .Z(n12164) );
  ANDN U13388 ( .B(y[2101]), .A(x[2101]), .Z(n16173) );
  NAND U13389 ( .A(n8409), .B(n24237), .Z(n8410) );
  NANDN U13390 ( .A(n24240), .B(n8410), .Z(n8413) );
  NANDN U13391 ( .A(x[2102]), .B(y[2102]), .Z(n8412) );
  NANDN U13392 ( .A(x[2103]), .B(y[2103]), .Z(n8411) );
  AND U13393 ( .A(n8412), .B(n8411), .Z(n24241) );
  NAND U13394 ( .A(n8413), .B(n24241), .Z(n8416) );
  NANDN U13395 ( .A(y[2104]), .B(x[2104]), .Z(n8415) );
  NANDN U13396 ( .A(y[2103]), .B(x[2103]), .Z(n8414) );
  NAND U13397 ( .A(n8415), .B(n8414), .Z(n24243) );
  ANDN U13398 ( .B(n8416), .A(n24243), .Z(n8419) );
  NANDN U13399 ( .A(x[2104]), .B(y[2104]), .Z(n8418) );
  NANDN U13400 ( .A(x[2105]), .B(y[2105]), .Z(n8417) );
  AND U13401 ( .A(n8418), .B(n8417), .Z(n24245) );
  NANDN U13402 ( .A(n8419), .B(n24245), .Z(n8420) );
  NANDN U13403 ( .A(n24248), .B(n8420), .Z(n8423) );
  NANDN U13404 ( .A(x[2106]), .B(y[2106]), .Z(n8422) );
  NANDN U13405 ( .A(x[2107]), .B(y[2107]), .Z(n8421) );
  AND U13406 ( .A(n8422), .B(n8421), .Z(n24249) );
  NAND U13407 ( .A(n8423), .B(n24249), .Z(n8424) );
  AND U13408 ( .A(n24251), .B(n8424), .Z(n8426) );
  NANDN U13409 ( .A(x[2108]), .B(y[2108]), .Z(n8425) );
  NANDN U13410 ( .A(x[2109]), .B(y[2109]), .Z(n16188) );
  NAND U13411 ( .A(n8425), .B(n16188), .Z(n24253) );
  OR U13412 ( .A(n8426), .B(n24253), .Z(n8427) );
  NAND U13413 ( .A(n8428), .B(n8427), .Z(n8429) );
  AND U13414 ( .A(n24257), .B(n8429), .Z(n8430) );
  OR U13415 ( .A(n12161), .B(n8430), .Z(n8433) );
  NANDN U13416 ( .A(x[2111]), .B(y[2111]), .Z(n8432) );
  NANDN U13417 ( .A(x[2112]), .B(y[2112]), .Z(n8431) );
  AND U13418 ( .A(n8432), .B(n8431), .Z(n24261) );
  NAND U13419 ( .A(n8433), .B(n24261), .Z(n8434) );
  NANDN U13420 ( .A(y[2112]), .B(x[2112]), .Z(n24264) );
  NAND U13421 ( .A(n8434), .B(n24264), .Z(n8435) );
  AND U13422 ( .A(n24265), .B(n8435), .Z(n8436) );
  NANDN U13423 ( .A(y[2113]), .B(x[2113]), .Z(n16194) );
  NANDN U13424 ( .A(y[2114]), .B(x[2114]), .Z(n16199) );
  NAND U13425 ( .A(n16194), .B(n16199), .Z(n24267) );
  OR U13426 ( .A(n8436), .B(n24267), .Z(n8437) );
  AND U13427 ( .A(n24269), .B(n8437), .Z(n8439) );
  NANDN U13428 ( .A(y[2115]), .B(x[2115]), .Z(n8438) );
  ANDN U13429 ( .B(x[2116]), .A(y[2116]), .Z(n16203) );
  ANDN U13430 ( .B(n8438), .A(n16203), .Z(n24271) );
  NANDN U13431 ( .A(n8439), .B(n24271), .Z(n8440) );
  NANDN U13432 ( .A(n16204), .B(n8440), .Z(n8441) );
  NANDN U13433 ( .A(n16208), .B(n8441), .Z(n8442) );
  AND U13434 ( .A(n24282), .B(n8442), .Z(n8445) );
  NANDN U13435 ( .A(y[2119]), .B(x[2119]), .Z(n8444) );
  NANDN U13436 ( .A(y[2120]), .B(x[2120]), .Z(n8443) );
  AND U13437 ( .A(n8444), .B(n8443), .Z(n24285) );
  NANDN U13438 ( .A(n8445), .B(n24285), .Z(n8446) );
  NANDN U13439 ( .A(n24287), .B(n8446), .Z(n8448) );
  NANDN U13440 ( .A(y[2122]), .B(x[2122]), .Z(n8447) );
  ANDN U13441 ( .B(x[2121]), .A(y[2121]), .Z(n16214) );
  ANDN U13442 ( .B(n8447), .A(n16214), .Z(n24288) );
  NAND U13443 ( .A(n8448), .B(n24288), .Z(n8450) );
  IV U13444 ( .A(x[2122]), .Z(n16217) );
  NAND U13445 ( .A(n16217), .B(y[2122]), .Z(n8449) );
  NANDN U13446 ( .A(x[2123]), .B(y[2123]), .Z(n16222) );
  NAND U13447 ( .A(n8449), .B(n16222), .Z(n24290) );
  ANDN U13448 ( .B(n8450), .A(n24290), .Z(n8452) );
  NANDN U13449 ( .A(y[2124]), .B(x[2124]), .Z(n16225) );
  NANDN U13450 ( .A(y[2123]), .B(x[2123]), .Z(n24292) );
  AND U13451 ( .A(n16225), .B(n24292), .Z(n8451) );
  NANDN U13452 ( .A(n8452), .B(n8451), .Z(n8456) );
  NANDN U13453 ( .A(x[2124]), .B(y[2124]), .Z(n8455) );
  NANDN U13454 ( .A(x[2125]), .B(y[2125]), .Z(n8453) );
  NANDN U13455 ( .A(n8454), .B(n8453), .Z(n16227) );
  ANDN U13456 ( .B(n8455), .A(n16227), .Z(n24294) );
  NAND U13457 ( .A(n8456), .B(n24294), .Z(n8459) );
  NANDN U13458 ( .A(y[2127]), .B(x[2127]), .Z(n8458) );
  NANDN U13459 ( .A(y[2126]), .B(x[2126]), .Z(n8457) );
  NAND U13460 ( .A(n8458), .B(n8457), .Z(n16228) );
  ANDN U13461 ( .B(n8459), .A(n16228), .Z(n8460) );
  NAND U13462 ( .A(n8461), .B(n8460), .Z(n8462) );
  NANDN U13463 ( .A(x[2127]), .B(y[2127]), .Z(n24298) );
  NAND U13464 ( .A(n8462), .B(n24298), .Z(n8463) );
  ANDN U13465 ( .B(x[2128]), .A(y[2128]), .Z(n16234) );
  IV U13466 ( .A(n16234), .Z(n24300) );
  AND U13467 ( .A(n8463), .B(n24300), .Z(n8465) );
  NANDN U13468 ( .A(x[2129]), .B(y[2129]), .Z(n8464) );
  ANDN U13469 ( .B(y[2128]), .A(x[2128]), .Z(n16231) );
  ANDN U13470 ( .B(n8464), .A(n16231), .Z(n24302) );
  NANDN U13471 ( .A(n8465), .B(n24302), .Z(n8466) );
  NANDN U13472 ( .A(n24305), .B(n8466), .Z(n8467) );
  NANDN U13473 ( .A(x[2130]), .B(y[2130]), .Z(n24306) );
  NAND U13474 ( .A(n8467), .B(n24306), .Z(n8468) );
  OR U13475 ( .A(n16243), .B(n8468), .Z(n8469) );
  AND U13476 ( .A(n8470), .B(n8469), .Z(n8472) );
  NANDN U13477 ( .A(x[2133]), .B(y[2133]), .Z(n24314) );
  ANDN U13478 ( .B(y[2132]), .A(x[2132]), .Z(n16244) );
  ANDN U13479 ( .B(n24314), .A(n16244), .Z(n8471) );
  NANDN U13480 ( .A(n8472), .B(n8471), .Z(n8473) );
  ANDN U13481 ( .B(x[2134]), .A(y[2134]), .Z(n16249) );
  IV U13482 ( .A(n16249), .Z(n24317) );
  AND U13483 ( .A(n8473), .B(n24317), .Z(n8474) );
  NANDN U13484 ( .A(n12157), .B(n8474), .Z(n8476) );
  NANDN U13485 ( .A(x[2135]), .B(y[2135]), .Z(n8475) );
  ANDN U13486 ( .B(y[2134]), .A(x[2134]), .Z(n12156) );
  ANDN U13487 ( .B(n8475), .A(n12156), .Z(n24318) );
  NAND U13488 ( .A(n8476), .B(n24318), .Z(n8477) );
  AND U13489 ( .A(n24320), .B(n8477), .Z(n8478) );
  NANDN U13490 ( .A(x[2136]), .B(y[2136]), .Z(n16257) );
  NANDN U13491 ( .A(x[2137]), .B(y[2137]), .Z(n16262) );
  NAND U13492 ( .A(n16257), .B(n16262), .Z(n24322) );
  OR U13493 ( .A(n8478), .B(n24322), .Z(n8479) );
  NAND U13494 ( .A(n8480), .B(n8479), .Z(n8481) );
  AND U13495 ( .A(n24326), .B(n8481), .Z(n8482) );
  ANDN U13496 ( .B(n8483), .A(n8482), .Z(n8484) );
  NANDN U13497 ( .A(n12155), .B(n8484), .Z(n8487) );
  NANDN U13498 ( .A(x[2141]), .B(y[2141]), .Z(n8486) );
  NANDN U13499 ( .A(x[2142]), .B(y[2142]), .Z(n8485) );
  AND U13500 ( .A(n8486), .B(n8485), .Z(n24330) );
  NAND U13501 ( .A(n8487), .B(n24330), .Z(n8488) );
  NANDN U13502 ( .A(y[2142]), .B(x[2142]), .Z(n24333) );
  NAND U13503 ( .A(n8488), .B(n24333), .Z(n8489) );
  AND U13504 ( .A(n24334), .B(n8489), .Z(n8490) );
  ANDN U13505 ( .B(x[2143]), .A(y[2143]), .Z(n16266) );
  ANDN U13506 ( .B(x[2144]), .A(y[2144]), .Z(n16270) );
  NOR U13507 ( .A(n16266), .B(n16270), .Z(n24336) );
  NANDN U13508 ( .A(n8490), .B(n24336), .Z(n8491) );
  AND U13509 ( .A(n24338), .B(n8491), .Z(n8494) );
  NANDN U13510 ( .A(y[2145]), .B(x[2145]), .Z(n8493) );
  NANDN U13511 ( .A(y[2146]), .B(x[2146]), .Z(n8492) );
  AND U13512 ( .A(n8493), .B(n8492), .Z(n24341) );
  NANDN U13513 ( .A(n8494), .B(n24341), .Z(n8495) );
  AND U13514 ( .A(n24342), .B(n8495), .Z(n8498) );
  NANDN U13515 ( .A(y[2147]), .B(x[2147]), .Z(n8497) );
  NANDN U13516 ( .A(y[2148]), .B(x[2148]), .Z(n8496) );
  AND U13517 ( .A(n8497), .B(n8496), .Z(n24344) );
  NANDN U13518 ( .A(n8498), .B(n24344), .Z(n8499) );
  AND U13519 ( .A(n24346), .B(n8499), .Z(n8502) );
  NANDN U13520 ( .A(y[2149]), .B(x[2149]), .Z(n8501) );
  NANDN U13521 ( .A(y[2150]), .B(x[2150]), .Z(n8500) );
  AND U13522 ( .A(n8501), .B(n8500), .Z(n24348) );
  NANDN U13523 ( .A(n8502), .B(n24348), .Z(n8505) );
  NANDN U13524 ( .A(x[2151]), .B(y[2151]), .Z(n8504) );
  NANDN U13525 ( .A(x[2150]), .B(y[2150]), .Z(n8503) );
  NAND U13526 ( .A(n8504), .B(n8503), .Z(n24351) );
  ANDN U13527 ( .B(n8505), .A(n24351), .Z(n8508) );
  NANDN U13528 ( .A(y[2151]), .B(x[2151]), .Z(n8507) );
  NANDN U13529 ( .A(y[2152]), .B(x[2152]), .Z(n8506) );
  AND U13530 ( .A(n8507), .B(n8506), .Z(n24352) );
  NANDN U13531 ( .A(n8508), .B(n24352), .Z(n8509) );
  NANDN U13532 ( .A(x[2152]), .B(y[2152]), .Z(n24355) );
  NAND U13533 ( .A(n8509), .B(n24355), .Z(n8511) );
  NANDN U13534 ( .A(y[2154]), .B(x[2154]), .Z(n8513) );
  NANDN U13535 ( .A(y[2153]), .B(x[2153]), .Z(n8510) );
  NAND U13536 ( .A(n8513), .B(n8510), .Z(n16283) );
  IV U13537 ( .A(n16283), .Z(n24357) );
  AND U13538 ( .A(n8511), .B(n24357), .Z(n8514) );
  IV U13539 ( .A(x[2155]), .Z(n12149) );
  NAND U13540 ( .A(n12149), .B(y[2155]), .Z(n12147) );
  NANDN U13541 ( .A(x[2153]), .B(y[2153]), .Z(n8512) );
  ANDN U13542 ( .B(y[2154]), .A(x[2154]), .Z(n16284) );
  ANDN U13543 ( .B(n8512), .A(n16284), .Z(n16280) );
  OR U13544 ( .A(n8514), .B(n24359), .Z(n8515) );
  NANDN U13545 ( .A(n24361), .B(n8515), .Z(n8516) );
  NANDN U13546 ( .A(n24363), .B(n8516), .Z(n8517) );
  AND U13547 ( .A(n24366), .B(n8517), .Z(n8518) );
  NANDN U13548 ( .A(x[2158]), .B(y[2158]), .Z(n24368) );
  NANDN U13549 ( .A(n8518), .B(n24368), .Z(n8519) );
  NANDN U13550 ( .A(n16296), .B(n8519), .Z(n8522) );
  NANDN U13551 ( .A(x[2160]), .B(y[2160]), .Z(n8521) );
  NANDN U13552 ( .A(x[2159]), .B(y[2159]), .Z(n8520) );
  AND U13553 ( .A(n8521), .B(n8520), .Z(n24372) );
  NAND U13554 ( .A(n8522), .B(n24372), .Z(n8523) );
  NANDN U13555 ( .A(y[2160]), .B(x[2160]), .Z(n24374) );
  NAND U13556 ( .A(n8523), .B(n24374), .Z(n8524) );
  NANDN U13557 ( .A(x[2161]), .B(y[2161]), .Z(n24377) );
  NAND U13558 ( .A(n8524), .B(n24377), .Z(n8525) );
  AND U13559 ( .A(n24378), .B(n8525), .Z(n8526) );
  OR U13560 ( .A(n24381), .B(n8526), .Z(n8528) );
  NANDN U13561 ( .A(y[2164]), .B(x[2164]), .Z(n8527) );
  ANDN U13562 ( .B(x[2163]), .A(y[2163]), .Z(n16306) );
  ANDN U13563 ( .B(n8527), .A(n16306), .Z(n24382) );
  NAND U13564 ( .A(n8528), .B(n24382), .Z(n8529) );
  NANDN U13565 ( .A(x[2164]), .B(y[2164]), .Z(n16311) );
  ANDN U13566 ( .B(y[2165]), .A(x[2165]), .Z(n16313) );
  ANDN U13567 ( .B(n16311), .A(n16313), .Z(n24384) );
  NAND U13568 ( .A(n8529), .B(n24384), .Z(n8530) );
  AND U13569 ( .A(n24386), .B(n8530), .Z(n8531) );
  NANDN U13570 ( .A(n12145), .B(n8531), .Z(n8532) );
  NANDN U13571 ( .A(x[2166]), .B(y[2166]), .Z(n24388) );
  AND U13572 ( .A(n8532), .B(n24388), .Z(n8533) );
  IV U13573 ( .A(x[2167]), .Z(n16317) );
  NANDN U13574 ( .A(n8533), .B(n16317), .Z(n8536) );
  XOR U13575 ( .A(x[2167]), .B(n8533), .Z(n8534) );
  NAND U13576 ( .A(n8534), .B(y[2167]), .Z(n8535) );
  NAND U13577 ( .A(n8536), .B(n8535), .Z(n8537) );
  NAND U13578 ( .A(n24394), .B(n8537), .Z(n8538) );
  AND U13579 ( .A(n24397), .B(n8538), .Z(n8539) );
  NANDN U13580 ( .A(n16319), .B(n8539), .Z(n8540) );
  NANDN U13581 ( .A(n24399), .B(n8540), .Z(n8542) );
  NANDN U13582 ( .A(x[2170]), .B(y[2170]), .Z(n8541) );
  NANDN U13583 ( .A(x[2171]), .B(y[2171]), .Z(n16329) );
  NAND U13584 ( .A(n8541), .B(n16329), .Z(n24401) );
  ANDN U13585 ( .B(n8542), .A(n24401), .Z(n8543) );
  OR U13586 ( .A(n24403), .B(n8543), .Z(n8544) );
  NAND U13587 ( .A(n8544), .B(n24404), .Z(n8545) );
  NANDN U13588 ( .A(n24406), .B(n8545), .Z(n8547) );
  NANDN U13589 ( .A(x[2174]), .B(y[2174]), .Z(n8546) );
  ANDN U13590 ( .B(y[2175]), .A(x[2175]), .Z(n16347) );
  ANDN U13591 ( .B(n8546), .A(n16347), .Z(n24408) );
  NAND U13592 ( .A(n8547), .B(n24408), .Z(n8549) );
  NANDN U13593 ( .A(y[2176]), .B(x[2176]), .Z(n8548) );
  NANDN U13594 ( .A(y[2175]), .B(x[2175]), .Z(n16345) );
  NAND U13595 ( .A(n8548), .B(n16345), .Z(n24411) );
  ANDN U13596 ( .B(n8549), .A(n24411), .Z(n8550) );
  OR U13597 ( .A(n24413), .B(n8550), .Z(n8552) );
  NANDN U13598 ( .A(y[2177]), .B(x[2177]), .Z(n8551) );
  NANDN U13599 ( .A(y[2178]), .B(x[2178]), .Z(n16360) );
  AND U13600 ( .A(n8551), .B(n16360), .Z(n24414) );
  NAND U13601 ( .A(n8552), .B(n24414), .Z(n8553) );
  ANDN U13602 ( .B(y[2179]), .A(x[2179]), .Z(n16363) );
  ANDN U13603 ( .B(y[2178]), .A(x[2178]), .Z(n16357) );
  NOR U13604 ( .A(n16363), .B(n16357), .Z(n24417) );
  NAND U13605 ( .A(n8553), .B(n24417), .Z(n8554) );
  NANDN U13606 ( .A(y[2179]), .B(x[2179]), .Z(n24418) );
  AND U13607 ( .A(n8554), .B(n24418), .Z(n8555) );
  NANDN U13608 ( .A(n12141), .B(n8555), .Z(n8556) );
  NANDN U13609 ( .A(n24420), .B(n8556), .Z(n8558) );
  NAND U13610 ( .A(n12137), .B(n8558), .Z(n8557) );
  ANDN U13611 ( .B(y[2182]), .A(x[2182]), .Z(n12139) );
  ANDN U13612 ( .B(n8557), .A(n12139), .Z(n8561) );
  XNOR U13613 ( .A(n8558), .B(x[2181]), .Z(n8559) );
  NAND U13614 ( .A(y[2181]), .B(n8559), .Z(n8560) );
  NAND U13615 ( .A(n8561), .B(n8560), .Z(n8564) );
  NANDN U13616 ( .A(y[2183]), .B(x[2183]), .Z(n8563) );
  NANDN U13617 ( .A(y[2182]), .B(x[2182]), .Z(n8562) );
  NAND U13618 ( .A(n8563), .B(n8562), .Z(n24426) );
  ANDN U13619 ( .B(n8564), .A(n24426), .Z(n8567) );
  NANDN U13620 ( .A(x[2183]), .B(y[2183]), .Z(n8566) );
  NANDN U13621 ( .A(x[2184]), .B(y[2184]), .Z(n8565) );
  AND U13622 ( .A(n8566), .B(n8565), .Z(n24428) );
  NANDN U13623 ( .A(n8567), .B(n24428), .Z(n8568) );
  NANDN U13624 ( .A(n16370), .B(n8568), .Z(n8569) );
  NANDN U13625 ( .A(n16372), .B(n8569), .Z(n8570) );
  NANDN U13626 ( .A(n24437), .B(n8570), .Z(n8573) );
  NANDN U13627 ( .A(x[2188]), .B(y[2188]), .Z(n8572) );
  NANDN U13628 ( .A(x[2187]), .B(y[2187]), .Z(n8571) );
  AND U13629 ( .A(n8572), .B(n8571), .Z(n24438) );
  NAND U13630 ( .A(n8573), .B(n24438), .Z(n8574) );
  AND U13631 ( .A(n24441), .B(n8574), .Z(n8575) );
  NANDN U13632 ( .A(x[2189]), .B(y[2189]), .Z(n24442) );
  NANDN U13633 ( .A(n8575), .B(n24442), .Z(n8577) );
  XNOR U13634 ( .A(y[2190]), .B(x[2190]), .Z(n8576) );
  NANDN U13635 ( .A(y[2189]), .B(x[2189]), .Z(n16376) );
  NAND U13636 ( .A(n8576), .B(n16376), .Z(n24444) );
  ANDN U13637 ( .B(n8577), .A(n24444), .Z(n8578) );
  ANDN U13638 ( .B(y[2190]), .A(x[2190]), .Z(n12136) );
  ANDN U13639 ( .B(y[2191]), .A(x[2191]), .Z(n16384) );
  NOR U13640 ( .A(n12136), .B(n16384), .Z(n24446) );
  NANDN U13641 ( .A(n8578), .B(n24446), .Z(n8579) );
  NANDN U13642 ( .A(n24449), .B(n8579), .Z(n8580) );
  ANDN U13643 ( .B(y[2193]), .A(x[2193]), .Z(n16392) );
  ANDN U13644 ( .B(y[2192]), .A(x[2192]), .Z(n16385) );
  NOR U13645 ( .A(n16392), .B(n16385), .Z(n24450) );
  NAND U13646 ( .A(n8580), .B(n24450), .Z(n8581) );
  NANDN U13647 ( .A(y[2193]), .B(x[2193]), .Z(n24452) );
  AND U13648 ( .A(n8581), .B(n24452), .Z(n8582) );
  NANDN U13649 ( .A(n12134), .B(n8582), .Z(n8583) );
  NANDN U13650 ( .A(x[2194]), .B(y[2194]), .Z(n24454) );
  NAND U13651 ( .A(n8583), .B(n24454), .Z(n8584) );
  NANDN U13652 ( .A(n12135), .B(n8584), .Z(n8585) );
  NANDN U13653 ( .A(n24459), .B(n8585), .Z(n8586) );
  NANDN U13654 ( .A(y[2196]), .B(x[2196]), .Z(n24460) );
  NAND U13655 ( .A(n8586), .B(n24460), .Z(n8587) );
  XOR U13656 ( .A(y[2197]), .B(x[2197]), .Z(n24462) );
  ANDN U13657 ( .B(n8587), .A(n24462), .Z(n8588) );
  OR U13658 ( .A(n24465), .B(n8588), .Z(n8589) );
  NANDN U13659 ( .A(n24466), .B(n8589), .Z(n8590) );
  NANDN U13660 ( .A(y[2199]), .B(x[2199]), .Z(n24469) );
  NAND U13661 ( .A(n8590), .B(n24469), .Z(n8591) );
  NANDN U13662 ( .A(x[2200]), .B(y[2200]), .Z(n24473) );
  NAND U13663 ( .A(n8591), .B(n24473), .Z(n8592) );
  NANDN U13664 ( .A(n16403), .B(n8592), .Z(n8595) );
  NANDN U13665 ( .A(x[2202]), .B(y[2202]), .Z(n8594) );
  NANDN U13666 ( .A(x[2201]), .B(y[2201]), .Z(n8593) );
  NAND U13667 ( .A(n8594), .B(n8593), .Z(n24476) );
  ANDN U13668 ( .B(n8595), .A(n24476), .Z(n8596) );
  NANDN U13669 ( .A(y[2202]), .B(x[2202]), .Z(n24478) );
  NANDN U13670 ( .A(n8596), .B(n24478), .Z(n8597) );
  NANDN U13671 ( .A(n24480), .B(n8597), .Z(n8603) );
  ANDN U13672 ( .B(x[2204]), .A(y[2204]), .Z(n16410) );
  NANDN U13673 ( .A(y[2203]), .B(x[2203]), .Z(n12133) );
  NANDN U13674 ( .A(n16410), .B(n12133), .Z(n8598) );
  NANDN U13675 ( .A(n8599), .B(n8598), .Z(n8602) );
  NANDN U13676 ( .A(y[2205]), .B(x[2205]), .Z(n8601) );
  NANDN U13677 ( .A(y[2206]), .B(x[2206]), .Z(n8600) );
  NAND U13678 ( .A(n8601), .B(n8600), .Z(n16409) );
  ANDN U13679 ( .B(n8602), .A(n16409), .Z(n24482) );
  NAND U13680 ( .A(n8603), .B(n24482), .Z(n8604) );
  NANDN U13681 ( .A(n24485), .B(n8604), .Z(n8605) );
  ANDN U13682 ( .B(x[2208]), .A(y[2208]), .Z(n12132) );
  ANDN U13683 ( .B(n8605), .A(n12132), .Z(n8606) );
  NANDN U13684 ( .A(y[2207]), .B(x[2207]), .Z(n24486) );
  NAND U13685 ( .A(n8606), .B(n24486), .Z(n8607) );
  ANDN U13686 ( .B(y[2208]), .A(x[2208]), .Z(n24488) );
  ANDN U13687 ( .B(n8607), .A(n24488), .Z(n8608) );
  IV U13688 ( .A(x[2209]), .Z(n12128) );
  NANDN U13689 ( .A(n8608), .B(n12128), .Z(n8611) );
  XOR U13690 ( .A(x[2209]), .B(n8608), .Z(n8609) );
  NAND U13691 ( .A(y[2209]), .B(n8609), .Z(n8610) );
  NAND U13692 ( .A(n8611), .B(n8610), .Z(n8612) );
  NANDN U13693 ( .A(n12124), .B(n8612), .Z(n8614) );
  ANDN U13694 ( .B(y[2211]), .A(x[2211]), .Z(n12125) );
  NANDN U13695 ( .A(x[2210]), .B(y[2210]), .Z(n8613) );
  NANDN U13696 ( .A(n12125), .B(n8613), .Z(n12130) );
  ANDN U13697 ( .B(n8614), .A(n12130), .Z(n8615) );
  OR U13698 ( .A(n8616), .B(n8615), .Z(n8617) );
  NANDN U13699 ( .A(n24496), .B(n8617), .Z(n8620) );
  NANDN U13700 ( .A(y[2213]), .B(x[2213]), .Z(n8619) );
  NANDN U13701 ( .A(y[2214]), .B(x[2214]), .Z(n8618) );
  AND U13702 ( .A(n8619), .B(n8618), .Z(n24498) );
  NAND U13703 ( .A(n8620), .B(n24498), .Z(n8623) );
  NANDN U13704 ( .A(x[2215]), .B(y[2215]), .Z(n8622) );
  NANDN U13705 ( .A(x[2214]), .B(y[2214]), .Z(n8621) );
  NAND U13706 ( .A(n8622), .B(n8621), .Z(n24500) );
  ANDN U13707 ( .B(n8623), .A(n24500), .Z(n8626) );
  NANDN U13708 ( .A(y[2216]), .B(x[2216]), .Z(n8625) );
  NANDN U13709 ( .A(y[2215]), .B(x[2215]), .Z(n8624) );
  AND U13710 ( .A(n8625), .B(n8624), .Z(n24502) );
  NANDN U13711 ( .A(n8626), .B(n24502), .Z(n8627) );
  NANDN U13712 ( .A(n16424), .B(n8627), .Z(n8628) );
  NANDN U13713 ( .A(n16427), .B(n8628), .Z(n8631) );
  NANDN U13714 ( .A(x[2219]), .B(y[2219]), .Z(n8630) );
  NANDN U13715 ( .A(x[2218]), .B(y[2218]), .Z(n8629) );
  NAND U13716 ( .A(n8630), .B(n8629), .Z(n24510) );
  ANDN U13717 ( .B(n8631), .A(n24510), .Z(n8632) );
  NANDN U13718 ( .A(y[2219]), .B(x[2219]), .Z(n16429) );
  ANDN U13719 ( .B(x[2220]), .A(y[2220]), .Z(n16432) );
  ANDN U13720 ( .B(n16429), .A(n16432), .Z(n24512) );
  NANDN U13721 ( .A(n8632), .B(n24512), .Z(n8633) );
  AND U13722 ( .A(n24514), .B(n8633), .Z(n8636) );
  NANDN U13723 ( .A(y[2222]), .B(x[2222]), .Z(n8635) );
  NANDN U13724 ( .A(y[2221]), .B(x[2221]), .Z(n8634) );
  AND U13725 ( .A(n8635), .B(n8634), .Z(n24516) );
  NANDN U13726 ( .A(n8636), .B(n24516), .Z(n8639) );
  NANDN U13727 ( .A(x[2222]), .B(y[2222]), .Z(n8638) );
  NANDN U13728 ( .A(x[2223]), .B(y[2223]), .Z(n8637) );
  AND U13729 ( .A(n8638), .B(n8637), .Z(n24518) );
  NAND U13730 ( .A(n8639), .B(n24518), .Z(n8642) );
  NANDN U13731 ( .A(y[2224]), .B(x[2224]), .Z(n8641) );
  NANDN U13732 ( .A(y[2223]), .B(x[2223]), .Z(n8640) );
  NAND U13733 ( .A(n8641), .B(n8640), .Z(n24521) );
  ANDN U13734 ( .B(n8642), .A(n24521), .Z(n8645) );
  NANDN U13735 ( .A(x[2224]), .B(y[2224]), .Z(n8644) );
  NANDN U13736 ( .A(x[2225]), .B(y[2225]), .Z(n8643) );
  AND U13737 ( .A(n8644), .B(n8643), .Z(n24522) );
  NANDN U13738 ( .A(n8645), .B(n24522), .Z(n8646) );
  AND U13739 ( .A(n24526), .B(n8646), .Z(n8647) );
  NANDN U13740 ( .A(x[2226]), .B(y[2226]), .Z(n24528) );
  NANDN U13741 ( .A(n8647), .B(n24528), .Z(n8649) );
  IV U13742 ( .A(y[2227]), .Z(n20253) );
  NAND U13743 ( .A(n20253), .B(x[2227]), .Z(n8648) );
  NANDN U13744 ( .A(y[2226]), .B(x[2226]), .Z(n24524) );
  NAND U13745 ( .A(n8648), .B(n24524), .Z(n16442) );
  ANDN U13746 ( .B(n8649), .A(n16442), .Z(n8650) );
  OR U13747 ( .A(n16444), .B(n8650), .Z(n8652) );
  NANDN U13748 ( .A(y[2228]), .B(x[2228]), .Z(n8651) );
  NANDN U13749 ( .A(y[2229]), .B(x[2229]), .Z(n24539) );
  NAND U13750 ( .A(n8651), .B(n24539), .Z(n16446) );
  ANDN U13751 ( .B(n8652), .A(n16446), .Z(n8655) );
  NANDN U13752 ( .A(x[2230]), .B(y[2230]), .Z(n8654) );
  NANDN U13753 ( .A(x[2229]), .B(y[2229]), .Z(n8653) );
  AND U13754 ( .A(n8654), .B(n8653), .Z(n24540) );
  NANDN U13755 ( .A(n8655), .B(n24540), .Z(n8656) );
  NANDN U13756 ( .A(y[2230]), .B(x[2230]), .Z(n24542) );
  NAND U13757 ( .A(n8656), .B(n24542), .Z(n8657) );
  AND U13758 ( .A(n24544), .B(n8657), .Z(n8658) );
  ANDN U13759 ( .B(x[2231]), .A(y[2231]), .Z(n16449) );
  XOR U13760 ( .A(x[2232]), .B(y[2232]), .Z(n16453) );
  NOR U13761 ( .A(n16449), .B(n16453), .Z(n24547) );
  NANDN U13762 ( .A(n8658), .B(n24547), .Z(n8659) );
  NANDN U13763 ( .A(n24549), .B(n8659), .Z(n8661) );
  NANDN U13764 ( .A(y[2234]), .B(x[2234]), .Z(n8660) );
  ANDN U13765 ( .B(x[2233]), .A(y[2233]), .Z(n16456) );
  ANDN U13766 ( .B(n8660), .A(n16456), .Z(n24550) );
  NAND U13767 ( .A(n8661), .B(n24550), .Z(n8662) );
  NANDN U13768 ( .A(n24552), .B(n8662), .Z(n8663) );
  AND U13769 ( .A(n24554), .B(n8663), .Z(n8664) );
  NANDN U13770 ( .A(n12115), .B(n8664), .Z(n8665) );
  NANDN U13771 ( .A(n12119), .B(n8665), .Z(n8668) );
  NANDN U13772 ( .A(y[2238]), .B(x[2238]), .Z(n24562) );
  ANDN U13773 ( .B(x[2237]), .A(y[2237]), .Z(n12114) );
  NAND U13774 ( .A(n20252), .B(n12114), .Z(n8666) );
  AND U13775 ( .A(n24562), .B(n8666), .Z(n8667) );
  NAND U13776 ( .A(n8668), .B(n8667), .Z(n8669) );
  AND U13777 ( .A(n20251), .B(n8669), .Z(n8671) );
  XNOR U13778 ( .A(y[2240]), .B(x[2240]), .Z(n8670) );
  ANDN U13779 ( .B(x[2239]), .A(y[2239]), .Z(n12113) );
  ANDN U13780 ( .B(n8670), .A(n12113), .Z(n24566) );
  NANDN U13781 ( .A(n8671), .B(n24566), .Z(n8672) );
  NANDN U13782 ( .A(n24569), .B(n8672), .Z(n8674) );
  IV U13783 ( .A(y[2241]), .Z(n12111) );
  NAND U13784 ( .A(n12111), .B(x[2241]), .Z(n8673) );
  ANDN U13785 ( .B(x[2242]), .A(y[2242]), .Z(n12109) );
  ANDN U13786 ( .B(n8673), .A(n12109), .Z(n24570) );
  NAND U13787 ( .A(n8674), .B(n24570), .Z(n8675) );
  AND U13788 ( .A(n24573), .B(n8675), .Z(n8676) );
  XNOR U13789 ( .A(x[2243]), .B(y[2243]), .Z(n24574) );
  NANDN U13790 ( .A(n8676), .B(n24574), .Z(n8677) );
  ANDN U13791 ( .B(y[2243]), .A(x[2243]), .Z(n16479) );
  ANDN U13792 ( .B(n8677), .A(n16479), .Z(n8678) );
  NANDN U13793 ( .A(y[2244]), .B(x[2244]), .Z(n24579) );
  NANDN U13794 ( .A(n8678), .B(n24579), .Z(n8679) );
  AND U13795 ( .A(n8680), .B(n8679), .Z(n8681) );
  NANDN U13796 ( .A(y[2245]), .B(x[2245]), .Z(n16481) );
  ANDN U13797 ( .B(x[2246]), .A(y[2246]), .Z(n16487) );
  ANDN U13798 ( .B(n16481), .A(n16487), .Z(n24582) );
  NANDN U13799 ( .A(n8681), .B(n24582), .Z(n8683) );
  NANDN U13800 ( .A(x[2246]), .B(y[2246]), .Z(n12108) );
  NANDN U13801 ( .A(x[2247]), .B(y[2247]), .Z(n8682) );
  AND U13802 ( .A(n12108), .B(n8682), .Z(n24584) );
  NAND U13803 ( .A(n8683), .B(n24584), .Z(n8684) );
  NANDN U13804 ( .A(n24586), .B(n8684), .Z(n8686) );
  IV U13805 ( .A(x[2248]), .Z(n16492) );
  NAND U13806 ( .A(n16492), .B(y[2248]), .Z(n8685) );
  ANDN U13807 ( .B(y[2249]), .A(x[2249]), .Z(n12107) );
  ANDN U13808 ( .B(n8685), .A(n12107), .Z(n24588) );
  NAND U13809 ( .A(n8686), .B(n24588), .Z(n8687) );
  ANDN U13810 ( .B(x[2250]), .A(y[2250]), .Z(n16501) );
  ANDN U13811 ( .B(n8687), .A(n16501), .Z(n8688) );
  NANDN U13812 ( .A(x[2250]), .B(y[2250]), .Z(n8691) );
  NANDN U13813 ( .A(x[2252]), .B(y[2252]), .Z(n8690) );
  NANDN U13814 ( .A(x[2251]), .B(y[2251]), .Z(n8689) );
  NAND U13815 ( .A(n8690), .B(n8689), .Z(n16503) );
  ANDN U13816 ( .B(n8691), .A(n16503), .Z(n24592) );
  NANDN U13817 ( .A(y[2251]), .B(x[2251]), .Z(n16500) );
  XNOR U13818 ( .A(x[2252]), .B(n16500), .Z(n8692) );
  NAND U13819 ( .A(n8692), .B(y[2252]), .Z(n8693) );
  NANDN U13820 ( .A(x[2253]), .B(y[2253]), .Z(n24596) );
  NANDN U13821 ( .A(y[2254]), .B(x[2254]), .Z(n16513) );
  NANDN U13822 ( .A(y[2253]), .B(x[2253]), .Z(n16506) );
  NAND U13823 ( .A(n16513), .B(n16506), .Z(n24598) );
  NANDN U13824 ( .A(x[2254]), .B(y[2254]), .Z(n8694) );
  ANDN U13825 ( .B(y[2255]), .A(x[2255]), .Z(n16514) );
  ANDN U13826 ( .B(n8694), .A(n16514), .Z(n24600) );
  NANDN U13827 ( .A(y[2256]), .B(x[2256]), .Z(n8696) );
  NANDN U13828 ( .A(y[2255]), .B(x[2255]), .Z(n8695) );
  NAND U13829 ( .A(n8696), .B(n8695), .Z(n24603) );
  NANDN U13830 ( .A(x[2256]), .B(y[2256]), .Z(n8698) );
  NANDN U13831 ( .A(x[2257]), .B(y[2257]), .Z(n8697) );
  AND U13832 ( .A(n8698), .B(n8697), .Z(n24604) );
  NANDN U13833 ( .A(y[2258]), .B(x[2258]), .Z(n8700) );
  NANDN U13834 ( .A(y[2257]), .B(x[2257]), .Z(n8699) );
  NAND U13835 ( .A(n8700), .B(n8699), .Z(n24606) );
  NANDN U13836 ( .A(x[2258]), .B(y[2258]), .Z(n8702) );
  NANDN U13837 ( .A(x[2259]), .B(y[2259]), .Z(n8701) );
  AND U13838 ( .A(n8702), .B(n8701), .Z(n24608) );
  NANDN U13839 ( .A(x[2261]), .B(y[2261]), .Z(n12106) );
  NANDN U13840 ( .A(x[2260]), .B(y[2260]), .Z(n12105) );
  NAND U13841 ( .A(n12106), .B(n12105), .Z(n24612) );
  NANDN U13842 ( .A(x[2263]), .B(y[2263]), .Z(n8704) );
  NANDN U13843 ( .A(x[2262]), .B(y[2262]), .Z(n8703) );
  AND U13844 ( .A(n8704), .B(n8703), .Z(n24616) );
  ANDN U13845 ( .B(x[2264]), .A(y[2264]), .Z(n16530) );
  NANDN U13846 ( .A(x[2264]), .B(y[2264]), .Z(n8705) );
  NANDN U13847 ( .A(x[2265]), .B(y[2265]), .Z(n16531) );
  AND U13848 ( .A(n8705), .B(n16531), .Z(n24621) );
  ANDN U13849 ( .B(x[2266]), .A(y[2266]), .Z(n12102) );
  ANDN U13850 ( .B(x[2265]), .A(y[2265]), .Z(n16532) );
  NOR U13851 ( .A(n12102), .B(n16532), .Z(n20249) );
  NAND U13852 ( .A(n8706), .B(n20249), .Z(n8707) );
  AND U13853 ( .A(n24624), .B(n8707), .Z(n8710) );
  NANDN U13854 ( .A(y[2267]), .B(x[2267]), .Z(n8709) );
  NANDN U13855 ( .A(y[2268]), .B(x[2268]), .Z(n8708) );
  AND U13856 ( .A(n8709), .B(n8708), .Z(n24626) );
  NANDN U13857 ( .A(n8710), .B(n24626), .Z(n8713) );
  NANDN U13858 ( .A(x[2269]), .B(y[2269]), .Z(n8712) );
  NANDN U13859 ( .A(x[2268]), .B(y[2268]), .Z(n8711) );
  NAND U13860 ( .A(n8712), .B(n8711), .Z(n24628) );
  ANDN U13861 ( .B(n8713), .A(n24628), .Z(n8714) );
  OR U13862 ( .A(n24631), .B(n8714), .Z(n8716) );
  NANDN U13863 ( .A(x[2270]), .B(y[2270]), .Z(n16543) );
  NANDN U13864 ( .A(x[2271]), .B(y[2271]), .Z(n8715) );
  NAND U13865 ( .A(n16543), .B(n8715), .Z(n24633) );
  ANDN U13866 ( .B(n8716), .A(n24633), .Z(n8718) );
  NANDN U13867 ( .A(y[2271]), .B(x[2271]), .Z(n8717) );
  ANDN U13868 ( .B(x[2272]), .A(y[2272]), .Z(n16549) );
  ANDN U13869 ( .B(n8717), .A(n16549), .Z(n24634) );
  NANDN U13870 ( .A(n8718), .B(n24634), .Z(n8721) );
  NANDN U13871 ( .A(x[2273]), .B(y[2273]), .Z(n8720) );
  NANDN U13872 ( .A(x[2272]), .B(y[2272]), .Z(n8719) );
  NAND U13873 ( .A(n8720), .B(n8719), .Z(n24636) );
  ANDN U13874 ( .B(n8721), .A(n24636), .Z(n8724) );
  NANDN U13875 ( .A(y[2273]), .B(x[2273]), .Z(n8723) );
  NANDN U13876 ( .A(y[2274]), .B(x[2274]), .Z(n8722) );
  AND U13877 ( .A(n8723), .B(n8722), .Z(n24638) );
  NANDN U13878 ( .A(n8724), .B(n24638), .Z(n8727) );
  NANDN U13879 ( .A(x[2275]), .B(y[2275]), .Z(n8726) );
  NANDN U13880 ( .A(x[2274]), .B(y[2274]), .Z(n8725) );
  NAND U13881 ( .A(n8726), .B(n8725), .Z(n24641) );
  ANDN U13882 ( .B(n8727), .A(n24641), .Z(n8730) );
  NANDN U13883 ( .A(y[2275]), .B(x[2275]), .Z(n8729) );
  NANDN U13884 ( .A(y[2276]), .B(x[2276]), .Z(n8728) );
  AND U13885 ( .A(n8729), .B(n8728), .Z(n24642) );
  NANDN U13886 ( .A(n8730), .B(n24642), .Z(n8733) );
  NANDN U13887 ( .A(x[2276]), .B(y[2276]), .Z(n8732) );
  NANDN U13888 ( .A(x[2277]), .B(y[2277]), .Z(n8731) );
  NAND U13889 ( .A(n8732), .B(n8731), .Z(n24645) );
  ANDN U13890 ( .B(n8733), .A(n24645), .Z(n8735) );
  NANDN U13891 ( .A(y[2277]), .B(x[2277]), .Z(n24646) );
  ANDN U13892 ( .B(x[2278]), .A(y[2278]), .Z(n16558) );
  ANDN U13893 ( .B(n24646), .A(n16558), .Z(n8734) );
  NANDN U13894 ( .A(n8735), .B(n8734), .Z(n8736) );
  NANDN U13895 ( .A(x[2278]), .B(y[2278]), .Z(n24649) );
  NAND U13896 ( .A(n8736), .B(n24649), .Z(n8737) );
  ANDN U13897 ( .B(x[2279]), .A(y[2279]), .Z(n16559) );
  ANDN U13898 ( .B(n8737), .A(n16559), .Z(n8740) );
  NANDN U13899 ( .A(x[2280]), .B(y[2280]), .Z(n8739) );
  NANDN U13900 ( .A(x[2279]), .B(y[2279]), .Z(n8738) );
  NAND U13901 ( .A(n8739), .B(n8738), .Z(n24652) );
  NOR U13902 ( .A(n8740), .B(n24652), .Z(n8745) );
  XNOR U13903 ( .A(x[2282]), .B(y[2282]), .Z(n8744) );
  NANDN U13904 ( .A(y[2280]), .B(x[2280]), .Z(n8742) );
  NANDN U13905 ( .A(y[2281]), .B(x[2281]), .Z(n8741) );
  NAND U13906 ( .A(n8742), .B(n8741), .Z(n8743) );
  ANDN U13907 ( .B(n8744), .A(n8743), .Z(n24654) );
  NANDN U13908 ( .A(n8745), .B(n24654), .Z(n8746) );
  NANDN U13909 ( .A(n24657), .B(n8746), .Z(n8747) );
  NANDN U13910 ( .A(y[2283]), .B(x[2283]), .Z(n24660) );
  NAND U13911 ( .A(n8747), .B(n24660), .Z(n8748) );
  NANDN U13912 ( .A(n24663), .B(n8748), .Z(n8753) );
  NANDN U13913 ( .A(y[2284]), .B(x[2284]), .Z(n24658) );
  OR U13914 ( .A(n8749), .B(n24658), .Z(n8752) );
  NANDN U13915 ( .A(y[2286]), .B(x[2286]), .Z(n8751) );
  NANDN U13916 ( .A(y[2285]), .B(x[2285]), .Z(n8750) );
  AND U13917 ( .A(n8751), .B(n8750), .Z(n24664) );
  NAND U13918 ( .A(n8752), .B(n24664), .Z(n16569) );
  ANDN U13919 ( .B(n8753), .A(n16569), .Z(n8756) );
  NANDN U13920 ( .A(x[2286]), .B(y[2286]), .Z(n8755) );
  NANDN U13921 ( .A(x[2287]), .B(y[2287]), .Z(n8754) );
  AND U13922 ( .A(n8755), .B(n8754), .Z(n24667) );
  NANDN U13923 ( .A(n8756), .B(n24667), .Z(n8757) );
  AND U13924 ( .A(n24668), .B(n8757), .Z(n8760) );
  NANDN U13925 ( .A(x[2288]), .B(y[2288]), .Z(n8759) );
  NANDN U13926 ( .A(x[2289]), .B(y[2289]), .Z(n8758) );
  AND U13927 ( .A(n8759), .B(n8758), .Z(n24670) );
  NANDN U13928 ( .A(n8760), .B(n24670), .Z(n8761) );
  AND U13929 ( .A(n24672), .B(n8761), .Z(n8763) );
  NANDN U13930 ( .A(x[2290]), .B(y[2290]), .Z(n24675) );
  ANDN U13931 ( .B(y[2291]), .A(x[2291]), .Z(n12101) );
  ANDN U13932 ( .B(n24675), .A(n12101), .Z(n8762) );
  NANDN U13933 ( .A(n8763), .B(n8762), .Z(n8764) );
  AND U13934 ( .A(n24676), .B(n8764), .Z(n8765) );
  NAND U13935 ( .A(n8766), .B(n8765), .Z(n8767) );
  NAND U13936 ( .A(n8768), .B(n8767), .Z(n8769) );
  AND U13937 ( .A(n24684), .B(n8769), .Z(n8770) );
  NANDN U13938 ( .A(n16578), .B(n8770), .Z(n8771) );
  NANDN U13939 ( .A(x[2295]), .B(y[2295]), .Z(n24686) );
  NAND U13940 ( .A(n8771), .B(n24686), .Z(n8772) );
  OR U13941 ( .A(n12099), .B(n8772), .Z(n8773) );
  AND U13942 ( .A(n24688), .B(n8773), .Z(n8774) );
  NANDN U13943 ( .A(x[2296]), .B(y[2296]), .Z(n16584) );
  ANDN U13944 ( .B(y[2297]), .A(x[2297]), .Z(n12096) );
  ANDN U13945 ( .B(n16584), .A(n12096), .Z(n24691) );
  NANDN U13946 ( .A(n8774), .B(n24691), .Z(n8775) );
  NANDN U13947 ( .A(n24693), .B(n8775), .Z(n8776) );
  NANDN U13948 ( .A(x[2298]), .B(y[2298]), .Z(n24694) );
  NANDN U13949 ( .A(y[2301]), .B(x[2301]), .Z(n16598) );
  ANDN U13950 ( .B(x[2302]), .A(y[2302]), .Z(n12094) );
  ANDN U13951 ( .B(n16598), .A(n12094), .Z(n24705) );
  NANDN U13952 ( .A(y[2304]), .B(x[2304]), .Z(n16609) );
  ANDN U13953 ( .B(x[2303]), .A(y[2303]), .Z(n12093) );
  ANDN U13954 ( .B(n16609), .A(n12093), .Z(n24708) );
  NANDN U13955 ( .A(y[2305]), .B(x[2305]), .Z(n24713) );
  NANDN U13956 ( .A(y[2308]), .B(x[2308]), .Z(n24719) );
  NANDN U13957 ( .A(x[2309]), .B(y[2309]), .Z(n8777) );
  ANDN U13958 ( .B(y[2308]), .A(x[2308]), .Z(n12090) );
  ANDN U13959 ( .B(n8777), .A(n12090), .Z(n24722) );
  IV U13960 ( .A(y[2309]), .Z(n12088) );
  NAND U13961 ( .A(n12088), .B(x[2309]), .Z(n16623) );
  NANDN U13962 ( .A(y[2310]), .B(x[2310]), .Z(n8778) );
  NAND U13963 ( .A(n16623), .B(n8778), .Z(n24724) );
  NANDN U13964 ( .A(x[2310]), .B(y[2310]), .Z(n8779) );
  ANDN U13965 ( .B(y[2311]), .A(x[2311]), .Z(n12085) );
  ANDN U13966 ( .B(n8779), .A(n12085), .Z(n24726) );
  NANDN U13967 ( .A(y[2311]), .B(x[2311]), .Z(n8780) );
  XOR U13968 ( .A(x[2312]), .B(y[2312]), .Z(n12086) );
  ANDN U13969 ( .B(n8780), .A(n12086), .Z(n24729) );
  AND U13970 ( .A(n24730), .B(n8781), .Z(n8782) );
  XNOR U13971 ( .A(x[2313]), .B(y[2313]), .Z(n24733) );
  NANDN U13972 ( .A(n8782), .B(n24733), .Z(n8783) );
  NANDN U13973 ( .A(n12084), .B(n8783), .Z(n8784) );
  NANDN U13974 ( .A(y[2314]), .B(x[2314]), .Z(n24736) );
  NAND U13975 ( .A(n8784), .B(n24736), .Z(n8785) );
  ANDN U13976 ( .B(y[2315]), .A(x[2315]), .Z(n24738) );
  ANDN U13977 ( .B(n8785), .A(n24738), .Z(n8786) );
  NANDN U13978 ( .A(n12083), .B(n8786), .Z(n8788) );
  NANDN U13979 ( .A(y[2316]), .B(x[2316]), .Z(n8787) );
  ANDN U13980 ( .B(x[2315]), .A(y[2315]), .Z(n12082) );
  ANDN U13981 ( .B(n8787), .A(n12082), .Z(n24740) );
  NAND U13982 ( .A(n8788), .B(n24740), .Z(n8789) );
  NANDN U13983 ( .A(n24743), .B(n8789), .Z(n8790) );
  AND U13984 ( .A(n24744), .B(n8790), .Z(n8791) );
  OR U13985 ( .A(n24747), .B(n8791), .Z(n8792) );
  ANDN U13986 ( .B(x[2319]), .A(y[2319]), .Z(n24749) );
  ANDN U13987 ( .B(n8792), .A(n24749), .Z(n8793) );
  NANDN U13988 ( .A(n16649), .B(n8793), .Z(n8794) );
  NANDN U13989 ( .A(x[2320]), .B(y[2320]), .Z(n24750) );
  NAND U13990 ( .A(n8794), .B(n24750), .Z(n8795) );
  NANDN U13991 ( .A(n16650), .B(n8795), .Z(n8798) );
  NANDN U13992 ( .A(x[2321]), .B(y[2321]), .Z(n8797) );
  NANDN U13993 ( .A(x[2322]), .B(y[2322]), .Z(n8796) );
  NAND U13994 ( .A(n8797), .B(n8796), .Z(n24755) );
  ANDN U13995 ( .B(n8798), .A(n24755), .Z(n8799) );
  NANDN U13996 ( .A(y[2322]), .B(x[2322]), .Z(n24756) );
  NANDN U13997 ( .A(n8799), .B(n24756), .Z(n8800) );
  NANDN U13998 ( .A(n24758), .B(n8800), .Z(n8806) );
  ANDN U13999 ( .B(x[2324]), .A(y[2324]), .Z(n12075) );
  NANDN U14000 ( .A(y[2323]), .B(x[2323]), .Z(n16653) );
  NANDN U14001 ( .A(n12075), .B(n16653), .Z(n8801) );
  NANDN U14002 ( .A(n8802), .B(n8801), .Z(n8805) );
  NANDN U14003 ( .A(y[2325]), .B(x[2325]), .Z(n8804) );
  NANDN U14004 ( .A(y[2326]), .B(x[2326]), .Z(n8803) );
  NAND U14005 ( .A(n8804), .B(n8803), .Z(n12077) );
  ANDN U14006 ( .B(n8805), .A(n12077), .Z(n24760) );
  NAND U14007 ( .A(n8806), .B(n24760), .Z(n8809) );
  NANDN U14008 ( .A(x[2326]), .B(y[2326]), .Z(n8808) );
  NANDN U14009 ( .A(x[2327]), .B(y[2327]), .Z(n8807) );
  NAND U14010 ( .A(n8808), .B(n8807), .Z(n24763) );
  ANDN U14011 ( .B(n8809), .A(n24763), .Z(n8810) );
  OR U14012 ( .A(n16661), .B(n8810), .Z(n8811) );
  NANDN U14013 ( .A(n16662), .B(n8811), .Z(n8812) );
  AND U14014 ( .A(n24773), .B(n8812), .Z(n8815) );
  NANDN U14015 ( .A(x[2330]), .B(y[2330]), .Z(n8814) );
  NANDN U14016 ( .A(x[2331]), .B(y[2331]), .Z(n8813) );
  AND U14017 ( .A(n8814), .B(n8813), .Z(n24775) );
  NANDN U14018 ( .A(n8815), .B(n24775), .Z(n8816) );
  NANDN U14019 ( .A(n24777), .B(n8816), .Z(n8819) );
  NANDN U14020 ( .A(x[2333]), .B(y[2333]), .Z(n8818) );
  NANDN U14021 ( .A(x[2332]), .B(y[2332]), .Z(n8817) );
  AND U14022 ( .A(n8818), .B(n8817), .Z(n24779) );
  NAND U14023 ( .A(n8819), .B(n24779), .Z(n8820) );
  AND U14024 ( .A(n24782), .B(n8820), .Z(n8821) );
  NANDN U14025 ( .A(n12070), .B(n8821), .Z(n8822) );
  AND U14026 ( .A(n24783), .B(n8822), .Z(n8823) );
  ANDN U14027 ( .B(n8824), .A(n8823), .Z(n8825) );
  NANDN U14028 ( .A(n12074), .B(n8825), .Z(n8826) );
  AND U14029 ( .A(n24787), .B(n8826), .Z(n8827) );
  NANDN U14030 ( .A(y[2338]), .B(x[2338]), .Z(n24790) );
  NANDN U14031 ( .A(n8827), .B(n24790), .Z(n8828) );
  ANDN U14032 ( .B(y[2339]), .A(x[2339]), .Z(n12068) );
  ANDN U14033 ( .B(y[2338]), .A(x[2338]), .Z(n16671) );
  NOR U14034 ( .A(n12068), .B(n16671), .Z(n24791) );
  NAND U14035 ( .A(n8828), .B(n24791), .Z(n8829) );
  NANDN U14036 ( .A(y[2339]), .B(x[2339]), .Z(n16675) );
  NANDN U14037 ( .A(y[2340]), .B(x[2340]), .Z(n16680) );
  NAND U14038 ( .A(n16675), .B(n16680), .Z(n24794) );
  ANDN U14039 ( .B(n8829), .A(n24794), .Z(n8831) );
  NANDN U14040 ( .A(x[2340]), .B(y[2340]), .Z(n24795) );
  ANDN U14041 ( .B(y[2341]), .A(x[2341]), .Z(n16682) );
  ANDN U14042 ( .B(n24795), .A(n16682), .Z(n8830) );
  NANDN U14043 ( .A(n8831), .B(n8830), .Z(n8832) );
  AND U14044 ( .A(n24798), .B(n8832), .Z(n8833) );
  NAND U14045 ( .A(n8834), .B(n8833), .Z(n8835) );
  ANDN U14046 ( .B(y[2345]), .A(x[2345]), .Z(n12064) );
  ANDN U14047 ( .B(y[2344]), .A(x[2344]), .Z(n12065) );
  NOR U14048 ( .A(n12064), .B(n12065), .Z(n24807) );
  NANDN U14049 ( .A(y[2347]), .B(x[2347]), .Z(n24813) );
  ANDN U14050 ( .B(x[2348]), .A(y[2348]), .Z(n16700) );
  NANDN U14051 ( .A(x[2348]), .B(y[2348]), .Z(n8838) );
  NANDN U14052 ( .A(x[2349]), .B(y[2349]), .Z(n8836) );
  NANDN U14053 ( .A(n8837), .B(n8836), .Z(n16702) );
  ANDN U14054 ( .B(n8838), .A(n16702), .Z(n24815) );
  NANDN U14055 ( .A(y[2351]), .B(x[2351]), .Z(n8840) );
  NANDN U14056 ( .A(y[2350]), .B(x[2350]), .Z(n8839) );
  NAND U14057 ( .A(n8840), .B(n8839), .Z(n16703) );
  NANDN U14058 ( .A(y[2355]), .B(x[2355]), .Z(n8842) );
  NANDN U14059 ( .A(y[2356]), .B(x[2356]), .Z(n8841) );
  AND U14060 ( .A(n8842), .B(n8841), .Z(n24826) );
  NANDN U14061 ( .A(y[2357]), .B(x[2357]), .Z(n8844) );
  NANDN U14062 ( .A(y[2358]), .B(x[2358]), .Z(n8843) );
  AND U14063 ( .A(n8844), .B(n8843), .Z(n24829) );
  NANDN U14064 ( .A(x[2359]), .B(y[2359]), .Z(n8846) );
  NANDN U14065 ( .A(x[2358]), .B(y[2358]), .Z(n8845) );
  AND U14066 ( .A(n8846), .B(n8845), .Z(n24831) );
  NAND U14067 ( .A(n8847), .B(n24831), .Z(n8848) );
  ANDN U14068 ( .B(x[2359]), .A(y[2359]), .Z(n16716) );
  NAND U14069 ( .A(n8848), .B(n24833), .Z(n8849) );
  NANDN U14070 ( .A(x[2361]), .B(y[2361]), .Z(n16724) );
  IV U14071 ( .A(x[2360]), .Z(n12058) );
  NAND U14072 ( .A(n12058), .B(y[2360]), .Z(n16721) );
  NAND U14073 ( .A(n16724), .B(n16721), .Z(n24835) );
  ANDN U14074 ( .B(n8849), .A(n24835), .Z(n8850) );
  ANDN U14075 ( .B(x[2361]), .A(y[2361]), .Z(n16722) );
  ANDN U14076 ( .B(x[2362]), .A(y[2362]), .Z(n16726) );
  NOR U14077 ( .A(n16722), .B(n16726), .Z(n24837) );
  NANDN U14078 ( .A(n8850), .B(n24837), .Z(n8851) );
  AND U14079 ( .A(n24840), .B(n8851), .Z(n8854) );
  NANDN U14080 ( .A(y[2363]), .B(x[2363]), .Z(n8852) );
  NAND U14081 ( .A(n8853), .B(n8852), .Z(n12057) );
  IV U14082 ( .A(n12057), .Z(n24841) );
  NANDN U14083 ( .A(n8854), .B(n24841), .Z(n8855) );
  NANDN U14084 ( .A(n24844), .B(n8855), .Z(n8856) );
  ANDN U14085 ( .B(x[2366]), .A(y[2366]), .Z(n12052) );
  NAND U14086 ( .A(n8856), .B(n24845), .Z(n8857) );
  NANDN U14087 ( .A(x[2366]), .B(y[2366]), .Z(n12054) );
  NANDN U14088 ( .A(x[2367]), .B(y[2367]), .Z(n16739) );
  AND U14089 ( .A(n12054), .B(n16739), .Z(n24847) );
  NAND U14090 ( .A(n8857), .B(n24847), .Z(n8858) );
  NANDN U14091 ( .A(n24852), .B(n8858), .Z(n8859) );
  AND U14092 ( .A(n24853), .B(n8859), .Z(n8860) );
  ANDN U14093 ( .B(x[2368]), .A(y[2368]), .Z(n24849) );
  ANDN U14094 ( .B(x[2369]), .A(y[2369]), .Z(n24855) );
  NOR U14095 ( .A(n24849), .B(n24855), .Z(n16743) );
  NANDN U14096 ( .A(n8860), .B(n16743), .Z(n8861) );
  ANDN U14097 ( .B(y[2369]), .A(x[2369]), .Z(n12050) );
  ANDN U14098 ( .B(n8861), .A(n12050), .Z(n8862) );
  OR U14099 ( .A(n24859), .B(n8862), .Z(n8863) );
  AND U14100 ( .A(n8864), .B(n8863), .Z(n8865) );
  ANDN U14101 ( .B(x[2371]), .A(y[2371]), .Z(n16745) );
  XOR U14102 ( .A(x[2372]), .B(y[2372]), .Z(n16749) );
  NOR U14103 ( .A(n16745), .B(n16749), .Z(n24864) );
  NANDN U14104 ( .A(n8865), .B(n24864), .Z(n8868) );
  NANDN U14105 ( .A(x[2372]), .B(y[2372]), .Z(n8867) );
  NANDN U14106 ( .A(x[2373]), .B(y[2373]), .Z(n8866) );
  AND U14107 ( .A(n8867), .B(n8866), .Z(n24865) );
  NAND U14108 ( .A(n8868), .B(n24865), .Z(n8869) );
  ANDN U14109 ( .B(x[2374]), .A(y[2374]), .Z(n12049) );
  ANDN U14110 ( .B(x[2373]), .A(y[2373]), .Z(n16753) );
  NOR U14111 ( .A(n12049), .B(n16753), .Z(n24867) );
  NAND U14112 ( .A(n8869), .B(n24867), .Z(n8870) );
  NANDN U14113 ( .A(x[2374]), .B(y[2374]), .Z(n16754) );
  ANDN U14114 ( .B(y[2375]), .A(x[2375]), .Z(n12048) );
  ANDN U14115 ( .B(n16754), .A(n12048), .Z(n24869) );
  NAND U14116 ( .A(n8870), .B(n24869), .Z(n8871) );
  AND U14117 ( .A(n8872), .B(n8871), .Z(n8874) );
  NANDN U14118 ( .A(x[2376]), .B(y[2376]), .Z(n8873) );
  ANDN U14119 ( .B(y[2377]), .A(x[2377]), .Z(n12045) );
  ANDN U14120 ( .B(n8873), .A(n12045), .Z(n24873) );
  NANDN U14121 ( .A(n8874), .B(n24873), .Z(n8875) );
  ANDN U14122 ( .B(x[2377]), .A(y[2377]), .Z(n12047) );
  ANDN U14123 ( .B(n8875), .A(n12047), .Z(n8876) );
  NANDN U14124 ( .A(n24875), .B(n8876), .Z(n8877) );
  AND U14125 ( .A(n24879), .B(n8877), .Z(n8878) );
  OR U14126 ( .A(n24881), .B(n8878), .Z(n8881) );
  NANDN U14127 ( .A(x[2380]), .B(y[2380]), .Z(n8880) );
  NANDN U14128 ( .A(x[2381]), .B(y[2381]), .Z(n8879) );
  AND U14129 ( .A(n8880), .B(n8879), .Z(n24883) );
  NAND U14130 ( .A(n8881), .B(n24883), .Z(n8883) );
  NANDN U14131 ( .A(y[2381]), .B(x[2381]), .Z(n8882) );
  ANDN U14132 ( .B(x[2382]), .A(y[2382]), .Z(n16780) );
  ANDN U14133 ( .B(n8882), .A(n16780), .Z(n24885) );
  NAND U14134 ( .A(n8883), .B(n24885), .Z(n8884) );
  ANDN U14135 ( .B(y[2383]), .A(x[2383]), .Z(n16784) );
  ANDN U14136 ( .B(y[2382]), .A(x[2382]), .Z(n16777) );
  NOR U14137 ( .A(n16784), .B(n16777), .Z(n24887) );
  NAND U14138 ( .A(n8884), .B(n24887), .Z(n8885) );
  AND U14139 ( .A(n24889), .B(n8885), .Z(n8886) );
  OR U14140 ( .A(n24891), .B(n8886), .Z(n8888) );
  NANDN U14141 ( .A(y[2385]), .B(x[2385]), .Z(n8887) );
  ANDN U14142 ( .B(x[2386]), .A(y[2386]), .Z(n16797) );
  ANDN U14143 ( .B(n8887), .A(n16797), .Z(n24893) );
  NAND U14144 ( .A(n8888), .B(n24893), .Z(n8890) );
  NANDN U14145 ( .A(x[2387]), .B(y[2387]), .Z(n8889) );
  ANDN U14146 ( .B(y[2386]), .A(x[2386]), .Z(n16795) );
  ANDN U14147 ( .B(n8889), .A(n16795), .Z(n24895) );
  NAND U14148 ( .A(n8890), .B(n24895), .Z(n8891) );
  NANDN U14149 ( .A(n24898), .B(n8891), .Z(n8893) );
  IV U14150 ( .A(x[2388]), .Z(n16804) );
  NAND U14151 ( .A(n16804), .B(y[2388]), .Z(n8892) );
  NANDN U14152 ( .A(x[2389]), .B(y[2389]), .Z(n12043) );
  NAND U14153 ( .A(n8892), .B(n12043), .Z(n24900) );
  ANDN U14154 ( .B(n8893), .A(n24900), .Z(n8895) );
  NANDN U14155 ( .A(y[2389]), .B(x[2389]), .Z(n24901) );
  ANDN U14156 ( .B(x[2390]), .A(y[2390]), .Z(n12042) );
  ANDN U14157 ( .B(n24901), .A(n12042), .Z(n8894) );
  NANDN U14158 ( .A(n8895), .B(n8894), .Z(n8896) );
  NANDN U14159 ( .A(x[2390]), .B(y[2390]), .Z(n24903) );
  NAND U14160 ( .A(n8896), .B(n24903), .Z(n8897) );
  NAND U14161 ( .A(n8898), .B(n8897), .Z(n8899) );
  NAND U14162 ( .A(n12040), .B(n8899), .Z(n8900) );
  NAND U14163 ( .A(n8901), .B(n8900), .Z(n8902) );
  NAND U14164 ( .A(n12039), .B(n8902), .Z(n8903) );
  ANDN U14165 ( .B(x[2393]), .A(y[2393]), .Z(n16814) );
  ANDN U14166 ( .B(n8903), .A(n16814), .Z(n8904) );
  NANDN U14167 ( .A(x[2393]), .B(y[2393]), .Z(n24911) );
  ANDN U14168 ( .B(y[2394]), .A(x[2394]), .Z(n24915) );
  ANDN U14169 ( .B(n24911), .A(n24915), .Z(n16816) );
  NANDN U14170 ( .A(n8904), .B(n16816), .Z(n8906) );
  NANDN U14171 ( .A(y[2394]), .B(x[2394]), .Z(n8905) );
  ANDN U14172 ( .B(x[2395]), .A(y[2395]), .Z(n24916) );
  ANDN U14173 ( .B(n8905), .A(n24916), .Z(n24914) );
  NAND U14174 ( .A(n8906), .B(n24914), .Z(n8909) );
  NANDN U14175 ( .A(x[2396]), .B(y[2396]), .Z(n8908) );
  NANDN U14176 ( .A(x[2395]), .B(y[2395]), .Z(n8907) );
  NAND U14177 ( .A(n8908), .B(n8907), .Z(n24917) );
  ANDN U14178 ( .B(n8909), .A(n24917), .Z(n8912) );
  NANDN U14179 ( .A(y[2396]), .B(x[2396]), .Z(n8911) );
  NANDN U14180 ( .A(y[2397]), .B(x[2397]), .Z(n8910) );
  AND U14181 ( .A(n8911), .B(n8910), .Z(n24921) );
  NANDN U14182 ( .A(n8912), .B(n24921), .Z(n8913) );
  ANDN U14183 ( .B(y[2397]), .A(x[2397]), .Z(n16821) );
  ANDN U14184 ( .B(n8913), .A(n16821), .Z(n8914) );
  OR U14185 ( .A(n24925), .B(n8914), .Z(n8915) );
  AND U14186 ( .A(n8916), .B(n8915), .Z(n8918) );
  XNOR U14187 ( .A(y[2400]), .B(x[2400]), .Z(n8917) );
  ANDN U14188 ( .B(x[2399]), .A(y[2399]), .Z(n12038) );
  ANDN U14189 ( .B(n8917), .A(n12038), .Z(n24929) );
  NANDN U14190 ( .A(n8918), .B(n24929), .Z(n8919) );
  IV U14191 ( .A(x[2401]), .Z(n12037) );
  NAND U14192 ( .A(n12037), .B(y[2401]), .Z(n12035) );
  ANDN U14193 ( .B(y[2400]), .A(x[2400]), .Z(n16828) );
  ANDN U14194 ( .B(n12035), .A(n16828), .Z(n24931) );
  NAND U14195 ( .A(n8919), .B(n24931), .Z(n8920) );
  ANDN U14196 ( .B(x[2402]), .A(y[2402]), .Z(n12034) );
  NAND U14197 ( .A(n8920), .B(n24934), .Z(n8921) );
  NANDN U14198 ( .A(x[2402]), .B(y[2402]), .Z(n12036) );
  NANDN U14199 ( .A(x[2403]), .B(y[2403]), .Z(n16837) );
  AND U14200 ( .A(n12036), .B(n16837), .Z(n24935) );
  NAND U14201 ( .A(n8921), .B(n24935), .Z(n8922) );
  ANDN U14202 ( .B(x[2404]), .A(y[2404]), .Z(n16840) );
  ANDN U14203 ( .B(n8922), .A(n16840), .Z(n8923) );
  NANDN U14204 ( .A(n24937), .B(n8923), .Z(n8924) );
  AND U14205 ( .A(n24939), .B(n8924), .Z(n8925) );
  OR U14206 ( .A(n16841), .B(n8925), .Z(n8928) );
  NANDN U14207 ( .A(x[2405]), .B(y[2405]), .Z(n8927) );
  NANDN U14208 ( .A(x[2406]), .B(y[2406]), .Z(n8926) );
  AND U14209 ( .A(n8927), .B(n8926), .Z(n24943) );
  NAND U14210 ( .A(n8928), .B(n24943), .Z(n8929) );
  AND U14211 ( .A(n24946), .B(n8929), .Z(n8930) );
  XNOR U14212 ( .A(y[2407]), .B(x[2407]), .Z(n24947) );
  NANDN U14213 ( .A(n8930), .B(n24947), .Z(n8931) );
  NANDN U14214 ( .A(n24950), .B(n8931), .Z(n8934) );
  NANDN U14215 ( .A(x[2408]), .B(y[2408]), .Z(n8933) );
  NANDN U14216 ( .A(x[2409]), .B(y[2409]), .Z(n8932) );
  AND U14217 ( .A(n8933), .B(n8932), .Z(n24951) );
  NAND U14218 ( .A(n8934), .B(n24951), .Z(n8935) );
  AND U14219 ( .A(n24955), .B(n8935), .Z(n8936) );
  NANDN U14220 ( .A(x[2410]), .B(y[2410]), .Z(n24957) );
  NANDN U14221 ( .A(n8936), .B(n24957), .Z(n8937) );
  NANDN U14222 ( .A(y[2411]), .B(x[2411]), .Z(n24959) );
  ANDN U14223 ( .B(x[2410]), .A(y[2410]), .Z(n24953) );
  ANDN U14224 ( .B(n24959), .A(n24953), .Z(n16850) );
  NAND U14225 ( .A(n8937), .B(n16850), .Z(n8938) );
  NANDN U14226 ( .A(n16852), .B(n8938), .Z(n8939) );
  NANDN U14227 ( .A(y[2412]), .B(x[2412]), .Z(n24963) );
  NAND U14228 ( .A(n8939), .B(n24963), .Z(n8940) );
  ANDN U14229 ( .B(y[2412]), .A(x[2412]), .Z(n16853) );
  ANDN U14230 ( .B(n8940), .A(n16853), .Z(n8941) );
  NANDN U14231 ( .A(x[2413]), .B(y[2413]), .Z(n24966) );
  NAND U14232 ( .A(n8941), .B(n24966), .Z(n8942) );
  AND U14233 ( .A(n24967), .B(n8942), .Z(n8943) );
  ANDN U14234 ( .B(y[2415]), .A(x[2415]), .Z(n16861) );
  ANDN U14235 ( .B(y[2414]), .A(x[2414]), .Z(n12032) );
  NOR U14236 ( .A(n16861), .B(n12032), .Z(n24970) );
  NANDN U14237 ( .A(n8943), .B(n24970), .Z(n8944) );
  AND U14238 ( .A(n24971), .B(n8944), .Z(n8947) );
  NANDN U14239 ( .A(x[2416]), .B(y[2416]), .Z(n8946) );
  NANDN U14240 ( .A(x[2417]), .B(y[2417]), .Z(n8945) );
  AND U14241 ( .A(n8946), .B(n8945), .Z(n24973) );
  NANDN U14242 ( .A(n8947), .B(n24973), .Z(n8948) );
  NAND U14243 ( .A(n8949), .B(n8948), .Z(n8950) );
  NANDN U14244 ( .A(x[2418]), .B(y[2418]), .Z(n24977) );
  NAND U14245 ( .A(n8950), .B(n24977), .Z(n8951) );
  NANDN U14246 ( .A(n8951), .B(x[2419]), .Z(n8954) );
  IV U14247 ( .A(y[2419]), .Z(n16868) );
  XNOR U14248 ( .A(n8951), .B(x[2419]), .Z(n8952) );
  NAND U14249 ( .A(n16868), .B(n8952), .Z(n8953) );
  NAND U14250 ( .A(n8954), .B(n8953), .Z(n8955) );
  OR U14251 ( .A(n12025), .B(n8955), .Z(n8956) );
  NANDN U14252 ( .A(n12030), .B(n8956), .Z(n8959) );
  NANDN U14253 ( .A(y[2421]), .B(x[2421]), .Z(n8958) );
  NANDN U14254 ( .A(y[2422]), .B(x[2422]), .Z(n8957) );
  NAND U14255 ( .A(n8958), .B(n8957), .Z(n12028) );
  ANDN U14256 ( .B(n8959), .A(n12028), .Z(n8962) );
  NANDN U14257 ( .A(x[2422]), .B(y[2422]), .Z(n8961) );
  NANDN U14258 ( .A(x[2423]), .B(y[2423]), .Z(n8960) );
  AND U14259 ( .A(n8961), .B(n8960), .Z(n24985) );
  NANDN U14260 ( .A(n8962), .B(n24985), .Z(n8963) );
  NANDN U14261 ( .A(n24987), .B(n8963), .Z(n8966) );
  NANDN U14262 ( .A(x[2425]), .B(y[2425]), .Z(n8965) );
  NANDN U14263 ( .A(x[2424]), .B(y[2424]), .Z(n8964) );
  AND U14264 ( .A(n8965), .B(n8964), .Z(n24989) );
  NAND U14265 ( .A(n8966), .B(n24989), .Z(n8967) );
  AND U14266 ( .A(n16877), .B(n8967), .Z(n8968) );
  OR U14267 ( .A(n16879), .B(n8968), .Z(n8969) );
  AND U14268 ( .A(n8970), .B(n8969), .Z(n8972) );
  NANDN U14269 ( .A(x[2429]), .B(y[2429]), .Z(n8971) );
  ANDN U14270 ( .B(y[2428]), .A(x[2428]), .Z(n16883) );
  ANDN U14271 ( .B(n8971), .A(n16883), .Z(n25003) );
  NANDN U14272 ( .A(n8972), .B(n25003), .Z(n8974) );
  NANDN U14273 ( .A(y[2429]), .B(x[2429]), .Z(n8973) );
  ANDN U14274 ( .B(x[2430]), .A(y[2430]), .Z(n16891) );
  ANDN U14275 ( .B(n8973), .A(n16891), .Z(n25005) );
  NAND U14276 ( .A(n8974), .B(n25005), .Z(n8976) );
  NANDN U14277 ( .A(x[2430]), .B(y[2430]), .Z(n8975) );
  ANDN U14278 ( .B(y[2431]), .A(x[2431]), .Z(n16892) );
  ANDN U14279 ( .B(n8975), .A(n16892), .Z(n25008) );
  NAND U14280 ( .A(n8976), .B(n25008), .Z(n8977) );
  NANDN U14281 ( .A(n16893), .B(n8977), .Z(n8978) );
  AND U14282 ( .A(n8979), .B(n8978), .Z(n8980) );
  NANDN U14283 ( .A(y[2433]), .B(x[2433]), .Z(n25015) );
  NANDN U14284 ( .A(n8980), .B(n25015), .Z(n8981) );
  ANDN U14285 ( .B(y[2434]), .A(x[2434]), .Z(n16900) );
  ANDN U14286 ( .B(n8981), .A(n16900), .Z(n8984) );
  NANDN U14287 ( .A(y[2434]), .B(x[2434]), .Z(n8983) );
  NANDN U14288 ( .A(y[2435]), .B(x[2435]), .Z(n8982) );
  AND U14289 ( .A(n8983), .B(n8982), .Z(n25019) );
  NANDN U14290 ( .A(n8984), .B(n25019), .Z(n8987) );
  NANDN U14291 ( .A(x[2436]), .B(y[2436]), .Z(n8986) );
  NANDN U14292 ( .A(x[2435]), .B(y[2435]), .Z(n8985) );
  NAND U14293 ( .A(n8986), .B(n8985), .Z(n25021) );
  ANDN U14294 ( .B(n8987), .A(n25021), .Z(n8990) );
  NANDN U14295 ( .A(y[2436]), .B(x[2436]), .Z(n8989) );
  NANDN U14296 ( .A(y[2437]), .B(x[2437]), .Z(n8988) );
  AND U14297 ( .A(n8989), .B(n8988), .Z(n25023) );
  NANDN U14298 ( .A(n8990), .B(n25023), .Z(n8991) );
  AND U14299 ( .A(n16905), .B(n8991), .Z(n8992) );
  NANDN U14300 ( .A(y[2439]), .B(x[2439]), .Z(n20248) );
  NANDN U14301 ( .A(y[2438]), .B(x[2438]), .Z(n20247) );
  NAND U14302 ( .A(n20248), .B(n20247), .Z(n16908) );
  OR U14303 ( .A(n8992), .B(n16908), .Z(n8993) );
  NANDN U14304 ( .A(n12023), .B(n8993), .Z(n8994) );
  NANDN U14305 ( .A(y[2440]), .B(x[2440]), .Z(n25033) );
  NAND U14306 ( .A(n8994), .B(n25033), .Z(n8995) );
  ANDN U14307 ( .B(y[2440]), .A(x[2440]), .Z(n12024) );
  ANDN U14308 ( .B(n8995), .A(n12024), .Z(n8996) );
  NANDN U14309 ( .A(x[2441]), .B(y[2441]), .Z(n25036) );
  NAND U14310 ( .A(n8996), .B(n25036), .Z(n8997) );
  ANDN U14311 ( .B(x[2441]), .A(y[2441]), .Z(n12022) );
  XOR U14312 ( .A(x[2442]), .B(y[2442]), .Z(n16914) );
  NOR U14313 ( .A(n12022), .B(n16914), .Z(n25037) );
  NAND U14314 ( .A(n8997), .B(n25037), .Z(n8998) );
  NANDN U14315 ( .A(n25040), .B(n8998), .Z(n8999) );
  AND U14316 ( .A(n25041), .B(n8999), .Z(n9001) );
  NANDN U14317 ( .A(x[2444]), .B(y[2444]), .Z(n9000) );
  ANDN U14318 ( .B(y[2445]), .A(x[2445]), .Z(n12021) );
  ANDN U14319 ( .B(n9000), .A(n12021), .Z(n25043) );
  NANDN U14320 ( .A(n9001), .B(n25043), .Z(n9002) );
  AND U14321 ( .A(n25045), .B(n9002), .Z(n9003) );
  NANDN U14322 ( .A(n12017), .B(n9003), .Z(n9005) );
  NANDN U14323 ( .A(x[2446]), .B(y[2446]), .Z(n9004) );
  ANDN U14324 ( .B(y[2447]), .A(x[2447]), .Z(n12018) );
  ANDN U14325 ( .B(n9004), .A(n12018), .Z(n25047) );
  NAND U14326 ( .A(n9005), .B(n25047), .Z(n9006) );
  NANDN U14327 ( .A(n25052), .B(n9006), .Z(n9007) );
  OR U14328 ( .A(n12020), .B(n9007), .Z(n9008) );
  AND U14329 ( .A(n25053), .B(n9008), .Z(n9009) );
  OR U14330 ( .A(n25055), .B(n9009), .Z(n9010) );
  ANDN U14331 ( .B(y[2451]), .A(x[2451]), .Z(n16937) );
  NAND U14332 ( .A(n9010), .B(n25057), .Z(n9011) );
  NANDN U14333 ( .A(n25060), .B(n9011), .Z(n9012) );
  AND U14334 ( .A(n25061), .B(n9012), .Z(n9013) );
  XNOR U14335 ( .A(y[2453]), .B(x[2453]), .Z(n25064) );
  NANDN U14336 ( .A(n9013), .B(n25064), .Z(n9014) );
  ANDN U14337 ( .B(y[2453]), .A(x[2453]), .Z(n16944) );
  ANDN U14338 ( .B(n9014), .A(n16944), .Z(n9015) );
  OR U14339 ( .A(n25067), .B(n9015), .Z(n9016) );
  AND U14340 ( .A(n9017), .B(n9016), .Z(n9019) );
  NANDN U14341 ( .A(y[2456]), .B(x[2456]), .Z(n9018) );
  ANDN U14342 ( .B(x[2455]), .A(y[2455]), .Z(n12013) );
  ANDN U14343 ( .B(n9018), .A(n12013), .Z(n25071) );
  NANDN U14344 ( .A(n9019), .B(n25071), .Z(n9020) );
  IV U14345 ( .A(x[2457]), .Z(n12012) );
  NAND U14346 ( .A(n12012), .B(y[2457]), .Z(n12011) );
  NAND U14347 ( .A(n9020), .B(n25073), .Z(n9021) );
  ANDN U14348 ( .B(x[2458]), .A(y[2458]), .Z(n12010) );
  NAND U14349 ( .A(n9021), .B(n25076), .Z(n9022) );
  NANDN U14350 ( .A(x[2458]), .B(y[2458]), .Z(n25077) );
  AND U14351 ( .A(n9022), .B(n25077), .Z(n9023) );
  NANDN U14352 ( .A(n12009), .B(n9023), .Z(n9024) );
  NANDN U14353 ( .A(n25080), .B(n9024), .Z(n9025) );
  NAND U14354 ( .A(n16960), .B(n9025), .Z(n9028) );
  XNOR U14355 ( .A(n9025), .B(y[2460]), .Z(n9026) );
  NAND U14356 ( .A(n9026), .B(x[2460]), .Z(n9027) );
  NAND U14357 ( .A(n9028), .B(n9027), .Z(n9029) );
  AND U14358 ( .A(n25085), .B(n9029), .Z(n9033) );
  NANDN U14359 ( .A(y[2462]), .B(x[2462]), .Z(n25087) );
  NANDN U14360 ( .A(y[2461]), .B(x[2461]), .Z(n16961) );
  NAND U14361 ( .A(n25087), .B(n16961), .Z(n9031) );
  ANDN U14362 ( .B(n9031), .A(n9030), .Z(n9032) );
  OR U14363 ( .A(n9033), .B(n9032), .Z(n9034) );
  NANDN U14364 ( .A(x[2463]), .B(y[2463]), .Z(n25089) );
  NAND U14365 ( .A(n9034), .B(n25089), .Z(n9035) );
  ANDN U14366 ( .B(x[2464]), .A(y[2464]), .Z(n12007) );
  ANDN U14367 ( .B(x[2463]), .A(y[2463]), .Z(n16965) );
  NOR U14368 ( .A(n12007), .B(n16965), .Z(n25092) );
  NAND U14369 ( .A(n9035), .B(n25092), .Z(n9036) );
  AND U14370 ( .A(n25093), .B(n9036), .Z(n9038) );
  NANDN U14371 ( .A(y[2465]), .B(x[2465]), .Z(n9037) );
  ANDN U14372 ( .B(x[2466]), .A(y[2466]), .Z(n16974) );
  ANDN U14373 ( .B(n9037), .A(n16974), .Z(n25096) );
  NANDN U14374 ( .A(n9038), .B(n25096), .Z(n9041) );
  NANDN U14375 ( .A(x[2467]), .B(y[2467]), .Z(n9040) );
  NANDN U14376 ( .A(x[2466]), .B(y[2466]), .Z(n9039) );
  AND U14377 ( .A(n9040), .B(n9039), .Z(n25097) );
  NAND U14378 ( .A(n9041), .B(n25097), .Z(n9044) );
  NANDN U14379 ( .A(y[2467]), .B(x[2467]), .Z(n9043) );
  NANDN U14380 ( .A(y[2468]), .B(x[2468]), .Z(n9042) );
  AND U14381 ( .A(n9043), .B(n9042), .Z(n25099) );
  NAND U14382 ( .A(n9044), .B(n25099), .Z(n9045) );
  AND U14383 ( .A(n25101), .B(n9045), .Z(n9048) );
  NANDN U14384 ( .A(y[2469]), .B(x[2469]), .Z(n9047) );
  NANDN U14385 ( .A(y[2470]), .B(x[2470]), .Z(n9046) );
  AND U14386 ( .A(n9047), .B(n9046), .Z(n25104) );
  NANDN U14387 ( .A(n9048), .B(n25104), .Z(n9051) );
  NANDN U14388 ( .A(x[2471]), .B(y[2471]), .Z(n9050) );
  NANDN U14389 ( .A(x[2470]), .B(y[2470]), .Z(n9049) );
  AND U14390 ( .A(n9050), .B(n9049), .Z(n25105) );
  NAND U14391 ( .A(n9051), .B(n25105), .Z(n9054) );
  NANDN U14392 ( .A(y[2471]), .B(x[2471]), .Z(n9053) );
  NANDN U14393 ( .A(y[2472]), .B(x[2472]), .Z(n9052) );
  AND U14394 ( .A(n9053), .B(n9052), .Z(n25107) );
  NAND U14395 ( .A(n9054), .B(n25107), .Z(n9057) );
  NANDN U14396 ( .A(x[2472]), .B(y[2472]), .Z(n9056) );
  NANDN U14397 ( .A(x[2473]), .B(y[2473]), .Z(n9055) );
  AND U14398 ( .A(n9056), .B(n9055), .Z(n25109) );
  NAND U14399 ( .A(n9057), .B(n25109), .Z(n9058) );
  ANDN U14400 ( .B(x[2474]), .A(y[2474]), .Z(n12005) );
  ANDN U14401 ( .B(n9058), .A(n12005), .Z(n9059) );
  NANDN U14402 ( .A(y[2473]), .B(x[2473]), .Z(n25112) );
  NAND U14403 ( .A(n9059), .B(n25112), .Z(n9060) );
  NANDN U14404 ( .A(x[2475]), .B(y[2475]), .Z(n25117) );
  AND U14405 ( .A(n9060), .B(n25117), .Z(n9061) );
  NANDN U14406 ( .A(x[2474]), .B(y[2474]), .Z(n25113) );
  NAND U14407 ( .A(n9061), .B(n25113), .Z(n9062) );
  NANDN U14408 ( .A(y[2476]), .B(x[2476]), .Z(n25120) );
  NAND U14409 ( .A(n9062), .B(n25120), .Z(n9063) );
  OR U14410 ( .A(n12006), .B(n9063), .Z(n9064) );
  AND U14411 ( .A(n25121), .B(n9064), .Z(n9065) );
  ANDN U14412 ( .B(x[2478]), .A(y[2478]), .Z(n12002) );
  ANDN U14413 ( .B(x[2477]), .A(y[2477]), .Z(n16990) );
  NOR U14414 ( .A(n12002), .B(n16990), .Z(n25123) );
  NANDN U14415 ( .A(n9065), .B(n25123), .Z(n9066) );
  NANDN U14416 ( .A(x[2479]), .B(y[2479]), .Z(n16998) );
  ANDN U14417 ( .B(y[2478]), .A(x[2478]), .Z(n12003) );
  ANDN U14418 ( .B(n16998), .A(n12003), .Z(n25125) );
  NAND U14419 ( .A(n9066), .B(n25125), .Z(n9067) );
  ANDN U14420 ( .B(x[2480]), .A(y[2480]), .Z(n17000) );
  ANDN U14421 ( .B(x[2479]), .A(y[2479]), .Z(n12001) );
  NOR U14422 ( .A(n17000), .B(n12001), .Z(n25128) );
  NAND U14423 ( .A(n9067), .B(n25128), .Z(n9068) );
  NAND U14424 ( .A(n9069), .B(n9068), .Z(n9070) );
  AND U14425 ( .A(n25136), .B(n9070), .Z(n9071) );
  NANDN U14426 ( .A(y[2481]), .B(x[2481]), .Z(n25131) );
  NAND U14427 ( .A(n9071), .B(n25131), .Z(n9072) );
  ANDN U14428 ( .B(y[2482]), .A(x[2482]), .Z(n12000) );
  ANDN U14429 ( .B(n9072), .A(n12000), .Z(n9073) );
  NANDN U14430 ( .A(x[2483]), .B(y[2483]), .Z(n25137) );
  NAND U14431 ( .A(n9073), .B(n25137), .Z(n9075) );
  NANDN U14432 ( .A(y[2483]), .B(x[2483]), .Z(n17005) );
  NANDN U14433 ( .A(y[2484]), .B(x[2484]), .Z(n9074) );
  NAND U14434 ( .A(n17005), .B(n9074), .Z(n25140) );
  ANDN U14435 ( .B(n9075), .A(n25140), .Z(n9077) );
  NANDN U14436 ( .A(x[2484]), .B(y[2484]), .Z(n9076) );
  ANDN U14437 ( .B(y[2485]), .A(x[2485]), .Z(n11996) );
  ANDN U14438 ( .B(n9076), .A(n11996), .Z(n25141) );
  NANDN U14439 ( .A(n9077), .B(n25141), .Z(n9078) );
  AND U14440 ( .A(n25143), .B(n9078), .Z(n9081) );
  NANDN U14441 ( .A(x[2486]), .B(y[2486]), .Z(n9080) );
  NANDN U14442 ( .A(x[2487]), .B(y[2487]), .Z(n9079) );
  AND U14443 ( .A(n9080), .B(n9079), .Z(n25145) );
  NANDN U14444 ( .A(n9081), .B(n25145), .Z(n9082) );
  NAND U14445 ( .A(n9083), .B(n9082), .Z(n9084) );
  NANDN U14446 ( .A(x[2488]), .B(y[2488]), .Z(n25149) );
  NAND U14447 ( .A(n9084), .B(n25149), .Z(n9085) );
  NANDN U14448 ( .A(n11995), .B(n9085), .Z(n9086) );
  AND U14449 ( .A(n25153), .B(n9086), .Z(n9090) );
  NANDN U14450 ( .A(y[2491]), .B(x[2491]), .Z(n9088) );
  NANDN U14451 ( .A(y[2490]), .B(x[2490]), .Z(n9087) );
  AND U14452 ( .A(n9088), .B(n9087), .Z(n9089) );
  XOR U14453 ( .A(x[2492]), .B(y[2492]), .Z(n9091) );
  ANDN U14454 ( .B(n9089), .A(n9091), .Z(n25155) );
  NANDN U14455 ( .A(n9090), .B(n25155), .Z(n9097) );
  NANDN U14456 ( .A(x[2492]), .B(y[2492]), .Z(n9094) );
  NOR U14457 ( .A(n9091), .B(x[2491]), .Z(n9092) );
  NAND U14458 ( .A(n9092), .B(y[2491]), .Z(n9093) );
  AND U14459 ( .A(n9094), .B(n9093), .Z(n9096) );
  NANDN U14460 ( .A(x[2493]), .B(y[2493]), .Z(n9095) );
  AND U14461 ( .A(n9096), .B(n9095), .Z(n25157) );
  NAND U14462 ( .A(n9097), .B(n25157), .Z(n9098) );
  NANDN U14463 ( .A(y[2493]), .B(x[2493]), .Z(n25161) );
  NAND U14464 ( .A(n9098), .B(n25161), .Z(n9099) );
  NANDN U14465 ( .A(n25164), .B(n9099), .Z(n9104) );
  NANDN U14466 ( .A(y[2494]), .B(x[2494]), .Z(n25160) );
  OR U14467 ( .A(n9100), .B(n25160), .Z(n9103) );
  NANDN U14468 ( .A(y[2496]), .B(x[2496]), .Z(n9102) );
  NANDN U14469 ( .A(y[2495]), .B(x[2495]), .Z(n9101) );
  AND U14470 ( .A(n9102), .B(n9101), .Z(n25165) );
  NAND U14471 ( .A(n9103), .B(n25165), .Z(n17023) );
  ANDN U14472 ( .B(n9104), .A(n17023), .Z(n9107) );
  NANDN U14473 ( .A(x[2496]), .B(y[2496]), .Z(n9106) );
  NANDN U14474 ( .A(x[2497]), .B(y[2497]), .Z(n9105) );
  AND U14475 ( .A(n9106), .B(n9105), .Z(n25168) );
  NANDN U14476 ( .A(n9107), .B(n25168), .Z(n9109) );
  XNOR U14477 ( .A(y[2498]), .B(x[2498]), .Z(n9108) );
  ANDN U14478 ( .B(x[2497]), .A(y[2497]), .Z(n17026) );
  ANDN U14479 ( .B(n9108), .A(n17026), .Z(n25169) );
  NAND U14480 ( .A(n9109), .B(n25169), .Z(n9110) );
  NANDN U14481 ( .A(n25172), .B(n9110), .Z(n9111) );
  ANDN U14482 ( .B(x[2500]), .A(y[2500]), .Z(n11993) );
  ANDN U14483 ( .B(x[2499]), .A(y[2499]), .Z(n17030) );
  NOR U14484 ( .A(n11993), .B(n17030), .Z(n25173) );
  NAND U14485 ( .A(n9111), .B(n25173), .Z(n9112) );
  ANDN U14486 ( .B(y[2501]), .A(x[2501]), .Z(n11992) );
  ANDN U14487 ( .B(n9112), .A(n11992), .Z(n9113) );
  NANDN U14488 ( .A(x[2500]), .B(y[2500]), .Z(n25175) );
  NAND U14489 ( .A(n9113), .B(n25175), .Z(n9114) );
  NANDN U14490 ( .A(y[2501]), .B(x[2501]), .Z(n25177) );
  NAND U14491 ( .A(n9114), .B(n25177), .Z(n9116) );
  XNOR U14492 ( .A(y[2502]), .B(n9116), .Z(n9115) );
  NAND U14493 ( .A(n11990), .B(n9115), .Z(n9118) );
  NANDN U14494 ( .A(n9116), .B(y[2502]), .Z(n9117) );
  AND U14495 ( .A(n9118), .B(n9117), .Z(n9119) );
  NAND U14496 ( .A(n9120), .B(n9119), .Z(n9121) );
  NAND U14497 ( .A(n9122), .B(n9121), .Z(n9123) );
  AND U14498 ( .A(n25188), .B(n9123), .Z(n9124) );
  NANDN U14499 ( .A(n11989), .B(n9124), .Z(n9125) );
  ANDN U14500 ( .B(x[2506]), .A(y[2506]), .Z(n11987) );
  ANDN U14501 ( .B(x[2505]), .A(y[2505]), .Z(n17044) );
  NOR U14502 ( .A(n11987), .B(n17044), .Z(n25189) );
  NANDN U14503 ( .A(x[2506]), .B(y[2506]), .Z(n17047) );
  NANDN U14504 ( .A(x[2507]), .B(y[2507]), .Z(n11985) );
  NAND U14505 ( .A(n17047), .B(n11985), .Z(n25192) );
  ANDN U14506 ( .B(x[2508]), .A(y[2508]), .Z(n11982) );
  ANDN U14507 ( .B(x[2507]), .A(y[2507]), .Z(n11986) );
  NOR U14508 ( .A(n11982), .B(n11986), .Z(n25193) );
  ANDN U14509 ( .B(x[2509]), .A(y[2509]), .Z(n11983) );
  NANDN U14510 ( .A(y[2510]), .B(x[2510]), .Z(n9126) );
  NAND U14511 ( .A(n9127), .B(n9126), .Z(n17059) );
  NOR U14512 ( .A(n11983), .B(n17059), .Z(n25197) );
  NANDN U14513 ( .A(y[2512]), .B(x[2512]), .Z(n9129) );
  NANDN U14514 ( .A(y[2513]), .B(x[2513]), .Z(n9128) );
  NAND U14515 ( .A(n9129), .B(n9128), .Z(n25202) );
  NANDN U14516 ( .A(x[2513]), .B(y[2513]), .Z(n25203) );
  NANDN U14517 ( .A(y[2514]), .B(x[2514]), .Z(n25206) );
  NANDN U14518 ( .A(y[2515]), .B(x[2515]), .Z(n20246) );
  NAND U14519 ( .A(n25206), .B(n20246), .Z(n17066) );
  ANDN U14520 ( .B(y[2515]), .A(x[2515]), .Z(n11979) );
  ANDN U14521 ( .B(y[2514]), .A(x[2514]), .Z(n17063) );
  NOR U14522 ( .A(n11979), .B(n17063), .Z(n25207) );
  NANDN U14523 ( .A(x[2516]), .B(y[2516]), .Z(n11978) );
  NAND U14524 ( .A(n11978), .B(n17074), .Z(n25212) );
  NANDN U14525 ( .A(x[2518]), .B(y[2518]), .Z(n17072) );
  ANDN U14526 ( .B(y[2519]), .A(x[2519]), .Z(n11976) );
  ANDN U14527 ( .B(n17072), .A(n11976), .Z(n25218) );
  NANDN U14528 ( .A(y[2519]), .B(x[2519]), .Z(n11977) );
  ANDN U14529 ( .B(x[2520]), .A(y[2520]), .Z(n17080) );
  ANDN U14530 ( .B(n11977), .A(n17080), .Z(n25219) );
  NANDN U14531 ( .A(x[2520]), .B(y[2520]), .Z(n9130) );
  ANDN U14532 ( .B(y[2521]), .A(x[2521]), .Z(n17081) );
  ANDN U14533 ( .B(n9130), .A(n17081), .Z(n25222) );
  NANDN U14534 ( .A(x[2522]), .B(y[2522]), .Z(n25225) );
  NANDN U14535 ( .A(n9131), .B(n25225), .Z(n9132) );
  AND U14536 ( .A(n25227), .B(n9132), .Z(n9133) );
  OR U14537 ( .A(n25230), .B(n9133), .Z(n9134) );
  AND U14538 ( .A(n25231), .B(n9134), .Z(n9135) );
  NANDN U14539 ( .A(x[2525]), .B(y[2525]), .Z(n25234) );
  NANDN U14540 ( .A(n9135), .B(n25234), .Z(n9136) );
  AND U14541 ( .A(n25235), .B(n9136), .Z(n9137) );
  ANDN U14542 ( .B(y[2527]), .A(x[2527]), .Z(n11972) );
  ANDN U14543 ( .B(y[2526]), .A(x[2526]), .Z(n17091) );
  NOR U14544 ( .A(n11972), .B(n17091), .Z(n25237) );
  NANDN U14545 ( .A(n9137), .B(n25237), .Z(n9138) );
  ANDN U14546 ( .B(x[2528]), .A(y[2528]), .Z(n11971) );
  ANDN U14547 ( .B(x[2527]), .A(y[2527]), .Z(n11975) );
  NOR U14548 ( .A(n11971), .B(n11975), .Z(n25239) );
  NAND U14549 ( .A(n9138), .B(n25239), .Z(n9139) );
  NANDN U14550 ( .A(x[2529]), .B(y[2529]), .Z(n17100) );
  ANDN U14551 ( .B(y[2528]), .A(x[2528]), .Z(n11973) );
  ANDN U14552 ( .B(n17100), .A(n11973), .Z(n25241) );
  NAND U14553 ( .A(n9139), .B(n25241), .Z(n9140) );
  AND U14554 ( .A(n25243), .B(n9140), .Z(n9141) );
  NANDN U14555 ( .A(n11969), .B(n9141), .Z(n9142) );
  NANDN U14556 ( .A(x[2530]), .B(y[2530]), .Z(n25246) );
  NAND U14557 ( .A(n9142), .B(n25246), .Z(n9143) );
  NANDN U14558 ( .A(n11970), .B(n9143), .Z(n9144) );
  NANDN U14559 ( .A(n25249), .B(n9144), .Z(n9145) );
  NANDN U14560 ( .A(y[2532]), .B(x[2532]), .Z(n25251) );
  NAND U14561 ( .A(n9145), .B(n25251), .Z(n9146) );
  AND U14562 ( .A(n25254), .B(n9146), .Z(n9147) );
  ANDN U14563 ( .B(x[2534]), .A(y[2534]), .Z(n11968) );
  ANDN U14564 ( .B(x[2533]), .A(y[2533]), .Z(n17105) );
  NOR U14565 ( .A(n11968), .B(n17105), .Z(n25255) );
  NANDN U14566 ( .A(n9147), .B(n25255), .Z(n9148) );
  NANDN U14567 ( .A(n25257), .B(n9148), .Z(n9150) );
  NANDN U14568 ( .A(y[2536]), .B(x[2536]), .Z(n17113) );
  NANDN U14569 ( .A(y[2535]), .B(x[2535]), .Z(n9149) );
  AND U14570 ( .A(n17113), .B(n9149), .Z(n25259) );
  NAND U14571 ( .A(n9150), .B(n25259), .Z(n9153) );
  NANDN U14572 ( .A(x[2537]), .B(y[2537]), .Z(n9152) );
  NANDN U14573 ( .A(x[2536]), .B(y[2536]), .Z(n9151) );
  NAND U14574 ( .A(n9152), .B(n9151), .Z(n25261) );
  ANDN U14575 ( .B(n9153), .A(n25261), .Z(n9156) );
  NANDN U14576 ( .A(y[2537]), .B(x[2537]), .Z(n9155) );
  NANDN U14577 ( .A(y[2538]), .B(x[2538]), .Z(n9154) );
  AND U14578 ( .A(n9155), .B(n9154), .Z(n25263) );
  NANDN U14579 ( .A(y[2539]), .B(x[2539]), .Z(n9158) );
  NANDN U14580 ( .A(y[2540]), .B(x[2540]), .Z(n9157) );
  AND U14581 ( .A(n9158), .B(n9157), .Z(n25267) );
  NANDN U14582 ( .A(x[2541]), .B(y[2541]), .Z(n9160) );
  NANDN U14583 ( .A(x[2540]), .B(y[2540]), .Z(n9159) );
  NAND U14584 ( .A(n9160), .B(n9159), .Z(n25269) );
  NANDN U14585 ( .A(y[2541]), .B(x[2541]), .Z(n9162) );
  NANDN U14586 ( .A(y[2542]), .B(x[2542]), .Z(n9161) );
  AND U14587 ( .A(n9162), .B(n9161), .Z(n25271) );
  NANDN U14588 ( .A(y[2543]), .B(x[2543]), .Z(n25275) );
  NANDN U14589 ( .A(y[2545]), .B(x[2545]), .Z(n17126) );
  NANDN U14590 ( .A(y[2547]), .B(x[2547]), .Z(n9165) );
  NANDN U14591 ( .A(y[2546]), .B(x[2546]), .Z(n9164) );
  NAND U14592 ( .A(n9165), .B(n9164), .Z(n17130) );
  NANDN U14593 ( .A(y[2548]), .B(x[2548]), .Z(n25283) );
  ANDN U14594 ( .B(x[2550]), .A(y[2550]), .Z(n11966) );
  ANDN U14595 ( .B(x[2549]), .A(y[2549]), .Z(n17135) );
  NOR U14596 ( .A(n11966), .B(n17135), .Z(n25287) );
  NANDN U14597 ( .A(y[2551]), .B(x[2551]), .Z(n25291) );
  IV U14598 ( .A(y[2552]), .Z(n11961) );
  NANDN U14599 ( .A(n9166), .B(n11961), .Z(n9169) );
  XOR U14600 ( .A(y[2552]), .B(n9166), .Z(n9167) );
  NAND U14601 ( .A(n9167), .B(x[2552]), .Z(n9168) );
  NAND U14602 ( .A(n9169), .B(n9168), .Z(n9170) );
  AND U14603 ( .A(n25298), .B(n9170), .Z(n9172) );
  NANDN U14604 ( .A(y[2554]), .B(x[2554]), .Z(n25299) );
  ANDN U14605 ( .B(x[2553]), .A(y[2553]), .Z(n11962) );
  ANDN U14606 ( .B(n25299), .A(n11962), .Z(n9171) );
  NANDN U14607 ( .A(n9172), .B(n9171), .Z(n9173) );
  NANDN U14608 ( .A(n25301), .B(n9173), .Z(n9174) );
  AND U14609 ( .A(n25303), .B(n9174), .Z(n9175) );
  OR U14610 ( .A(n25306), .B(n9175), .Z(n9176) );
  AND U14611 ( .A(n25307), .B(n9176), .Z(n9177) );
  NANDN U14612 ( .A(n17158), .B(n9177), .Z(n9178) );
  ANDN U14613 ( .B(y[2559]), .A(x[2559]), .Z(n11956) );
  ANDN U14614 ( .B(n9178), .A(n11956), .Z(n9179) );
  NANDN U14615 ( .A(x[2558]), .B(y[2558]), .Z(n25309) );
  NAND U14616 ( .A(n9179), .B(n25309), .Z(n9180) );
  ANDN U14617 ( .B(x[2559]), .A(y[2559]), .Z(n17159) );
  ANDN U14618 ( .B(n9180), .A(n17159), .Z(n9181) );
  NANDN U14619 ( .A(y[2560]), .B(x[2560]), .Z(n25315) );
  NAND U14620 ( .A(n9181), .B(n25315), .Z(n9182) );
  NANDN U14621 ( .A(x[2561]), .B(y[2561]), .Z(n25317) );
  NAND U14622 ( .A(n9182), .B(n25317), .Z(n9183) );
  OR U14623 ( .A(n11957), .B(n9183), .Z(n9184) );
  AND U14624 ( .A(n25319), .B(n9184), .Z(n9187) );
  NANDN U14625 ( .A(x[2562]), .B(y[2562]), .Z(n9186) );
  NANDN U14626 ( .A(x[2563]), .B(y[2563]), .Z(n9185) );
  AND U14627 ( .A(n9186), .B(n9185), .Z(n25322) );
  NANDN U14628 ( .A(n9187), .B(n25322), .Z(n9188) );
  AND U14629 ( .A(n25323), .B(n9188), .Z(n9191) );
  NANDN U14630 ( .A(x[2564]), .B(y[2564]), .Z(n9190) );
  NANDN U14631 ( .A(x[2565]), .B(y[2565]), .Z(n9189) );
  AND U14632 ( .A(n9190), .B(n9189), .Z(n25325) );
  NANDN U14633 ( .A(n9191), .B(n25325), .Z(n9192) );
  AND U14634 ( .A(n25327), .B(n9192), .Z(n9193) );
  OR U14635 ( .A(n25329), .B(n9193), .Z(n9196) );
  NANDN U14636 ( .A(y[2567]), .B(x[2567]), .Z(n9195) );
  NANDN U14637 ( .A(y[2568]), .B(x[2568]), .Z(n9194) );
  AND U14638 ( .A(n9195), .B(n9194), .Z(n25331) );
  NAND U14639 ( .A(n9196), .B(n25331), .Z(n9199) );
  NANDN U14640 ( .A(x[2569]), .B(y[2569]), .Z(n9198) );
  NANDN U14641 ( .A(x[2568]), .B(y[2568]), .Z(n9197) );
  NAND U14642 ( .A(n9198), .B(n9197), .Z(n25334) );
  ANDN U14643 ( .B(n9199), .A(n25334), .Z(n9202) );
  NANDN U14644 ( .A(y[2569]), .B(x[2569]), .Z(n9201) );
  NANDN U14645 ( .A(y[2570]), .B(x[2570]), .Z(n9200) );
  AND U14646 ( .A(n9201), .B(n9200), .Z(n25335) );
  NANDN U14647 ( .A(n9202), .B(n25335), .Z(n9205) );
  NANDN U14648 ( .A(x[2571]), .B(y[2571]), .Z(n9204) );
  NANDN U14649 ( .A(x[2570]), .B(y[2570]), .Z(n9203) );
  NAND U14650 ( .A(n9204), .B(n9203), .Z(n25338) );
  ANDN U14651 ( .B(n9205), .A(n25338), .Z(n9208) );
  NANDN U14652 ( .A(y[2571]), .B(x[2571]), .Z(n9207) );
  NANDN U14653 ( .A(y[2572]), .B(x[2572]), .Z(n9206) );
  AND U14654 ( .A(n9207), .B(n9206), .Z(n25339) );
  NANDN U14655 ( .A(n9208), .B(n25339), .Z(n9212) );
  XNOR U14656 ( .A(y[2574]), .B(x[2574]), .Z(n9211) );
  NANDN U14657 ( .A(x[2573]), .B(y[2573]), .Z(n9210) );
  NANDN U14658 ( .A(x[2572]), .B(y[2572]), .Z(n9209) );
  AND U14659 ( .A(n9210), .B(n9209), .Z(n25341) );
  NAND U14660 ( .A(n9211), .B(n25341), .Z(n17176) );
  ANDN U14661 ( .B(n9212), .A(n17176), .Z(n9213) );
  OR U14662 ( .A(n17178), .B(n9213), .Z(n9214) );
  NANDN U14663 ( .A(x[2575]), .B(y[2575]), .Z(n25346) );
  NAND U14664 ( .A(n9214), .B(n25346), .Z(n9215) );
  NANDN U14665 ( .A(n25350), .B(n9215), .Z(n9217) );
  IV U14666 ( .A(x[2576]), .Z(n17182) );
  NAND U14667 ( .A(n17182), .B(y[2576]), .Z(n9216) );
  ANDN U14668 ( .B(y[2577]), .A(x[2577]), .Z(n17188) );
  ANDN U14669 ( .B(n9216), .A(n17188), .Z(n25351) );
  NAND U14670 ( .A(n9217), .B(n25351), .Z(n9218) );
  NANDN U14671 ( .A(y[2577]), .B(x[2577]), .Z(n25356) );
  NAND U14672 ( .A(n9218), .B(n25356), .Z(n9219) );
  AND U14673 ( .A(n25357), .B(n9219), .Z(n9220) );
  ANDN U14674 ( .B(x[2578]), .A(y[2578]), .Z(n25353) );
  ANDN U14675 ( .B(x[2579]), .A(y[2579]), .Z(n25360) );
  NOR U14676 ( .A(n25353), .B(n25360), .Z(n17192) );
  NANDN U14677 ( .A(n9220), .B(n17192), .Z(n9221) );
  ANDN U14678 ( .B(y[2579]), .A(x[2579]), .Z(n11954) );
  ANDN U14679 ( .B(n9221), .A(n11954), .Z(n9222) );
  OR U14680 ( .A(n25363), .B(n9222), .Z(n9223) );
  AND U14681 ( .A(n9224), .B(n9223), .Z(n9225) );
  ANDN U14682 ( .B(x[2581]), .A(y[2581]), .Z(n17194) );
  XOR U14683 ( .A(x[2582]), .B(y[2582]), .Z(n17199) );
  NOR U14684 ( .A(n17194), .B(n17199), .Z(n25367) );
  NANDN U14685 ( .A(n9225), .B(n25367), .Z(n9228) );
  NANDN U14686 ( .A(x[2582]), .B(y[2582]), .Z(n9227) );
  NANDN U14687 ( .A(x[2583]), .B(y[2583]), .Z(n9226) );
  AND U14688 ( .A(n9227), .B(n9226), .Z(n25369) );
  NANDN U14689 ( .A(x[2586]), .B(y[2586]), .Z(n9229) );
  ANDN U14690 ( .B(y[2587]), .A(x[2587]), .Z(n11950) );
  ANDN U14691 ( .B(n9229), .A(n11950), .Z(n25377) );
  ANDN U14692 ( .B(x[2587]), .A(y[2587]), .Z(n11952) );
  NANDN U14693 ( .A(y[2588]), .B(x[2588]), .Z(n20244) );
  XNOR U14694 ( .A(x[2590]), .B(y[2590]), .Z(n17216) );
  ANDN U14695 ( .B(x[2589]), .A(y[2589]), .Z(n17213) );
  ANDN U14696 ( .B(n17216), .A(n17213), .Z(n25383) );
  NANDN U14697 ( .A(x[2590]), .B(y[2590]), .Z(n9230) );
  IV U14698 ( .A(x[2591]), .Z(n11948) );
  NAND U14699 ( .A(n11948), .B(y[2591]), .Z(n11946) );
  AND U14700 ( .A(n9230), .B(n11946), .Z(n25385) );
  ANDN U14701 ( .B(x[2592]), .A(y[2592]), .Z(n17227) );
  ANDN U14702 ( .B(x[2596]), .A(y[2596]), .Z(n17245) );
  ANDN U14703 ( .B(x[2595]), .A(y[2595]), .Z(n17241) );
  NOR U14704 ( .A(n17245), .B(n17241), .Z(n25395) );
  NANDN U14705 ( .A(y[2597]), .B(x[2597]), .Z(n25399) );
  IV U14706 ( .A(x[2598]), .Z(n17246) );
  NANDN U14707 ( .A(x[2604]), .B(y[2604]), .Z(n9233) );
  NANDN U14708 ( .A(x[2603]), .B(y[2603]), .Z(n9232) );
  NAND U14709 ( .A(n9233), .B(n9232), .Z(n25414) );
  NANDN U14710 ( .A(y[2604]), .B(x[2604]), .Z(n9235) );
  NANDN U14711 ( .A(y[2605]), .B(x[2605]), .Z(n9234) );
  AND U14712 ( .A(n9235), .B(n9234), .Z(n25415) );
  NANDN U14713 ( .A(x[2606]), .B(y[2606]), .Z(n9237) );
  NANDN U14714 ( .A(x[2605]), .B(y[2605]), .Z(n9236) );
  NAND U14715 ( .A(n9237), .B(n9236), .Z(n25418) );
  NANDN U14716 ( .A(y[2606]), .B(x[2606]), .Z(n9239) );
  NANDN U14717 ( .A(y[2607]), .B(x[2607]), .Z(n9238) );
  AND U14718 ( .A(n9239), .B(n9238), .Z(n25419) );
  NANDN U14719 ( .A(n25421), .B(n9240), .Z(n9243) );
  NANDN U14720 ( .A(y[2608]), .B(x[2608]), .Z(n9242) );
  NANDN U14721 ( .A(y[2609]), .B(x[2609]), .Z(n9241) );
  AND U14722 ( .A(n9242), .B(n9241), .Z(n25423) );
  NAND U14723 ( .A(n9243), .B(n25423), .Z(n9244) );
  NANDN U14724 ( .A(n25425), .B(n9244), .Z(n9245) );
  NANDN U14725 ( .A(y[2610]), .B(x[2610]), .Z(n25427) );
  NAND U14726 ( .A(n9245), .B(n25427), .Z(n9246) );
  ANDN U14727 ( .B(y[2611]), .A(x[2611]), .Z(n25429) );
  ANDN U14728 ( .B(n9246), .A(n25429), .Z(n9248) );
  IV U14729 ( .A(y[2612]), .Z(n17267) );
  NAND U14730 ( .A(n17267), .B(x[2612]), .Z(n9247) );
  ANDN U14731 ( .B(x[2611]), .A(y[2611]), .Z(n11937) );
  ANDN U14732 ( .B(n9247), .A(n11937), .Z(n25431) );
  NANDN U14733 ( .A(n9248), .B(n25431), .Z(n9249) );
  NANDN U14734 ( .A(n25433), .B(n9249), .Z(n9250) );
  NANDN U14735 ( .A(n25435), .B(n9250), .Z(n9251) );
  AND U14736 ( .A(n25438), .B(n9251), .Z(n9252) );
  NANDN U14737 ( .A(y[2615]), .B(x[2615]), .Z(n25439) );
  NANDN U14738 ( .A(n9252), .B(n25439), .Z(n9255) );
  NANDN U14739 ( .A(x[2616]), .B(y[2616]), .Z(n9254) );
  NANDN U14740 ( .A(x[2615]), .B(y[2615]), .Z(n9253) );
  NAND U14741 ( .A(n9254), .B(n9253), .Z(n25441) );
  ANDN U14742 ( .B(n9255), .A(n25441), .Z(n9258) );
  NANDN U14743 ( .A(y[2616]), .B(x[2616]), .Z(n9257) );
  NANDN U14744 ( .A(y[2617]), .B(x[2617]), .Z(n9256) );
  AND U14745 ( .A(n9257), .B(n9256), .Z(n25443) );
  NANDN U14746 ( .A(n9258), .B(n25443), .Z(n9259) );
  AND U14747 ( .A(n25445), .B(n9259), .Z(n9260) );
  OR U14748 ( .A(n25447), .B(n9260), .Z(n9261) );
  ANDN U14749 ( .B(y[2619]), .A(x[2619]), .Z(n11936) );
  ANDN U14750 ( .B(y[2618]), .A(x[2618]), .Z(n17280) );
  NOR U14751 ( .A(n11936), .B(n17280), .Z(n25449) );
  NAND U14752 ( .A(n9261), .B(n25449), .Z(n9262) );
  NANDN U14753 ( .A(y[2619]), .B(x[2619]), .Z(n25454) );
  NAND U14754 ( .A(n9262), .B(n25454), .Z(n9263) );
  ANDN U14755 ( .B(y[2620]), .A(x[2620]), .Z(n25455) );
  ANDN U14756 ( .B(n9263), .A(n25455), .Z(n9265) );
  NANDN U14757 ( .A(y[2621]), .B(x[2621]), .Z(n9264) );
  ANDN U14758 ( .B(x[2620]), .A(y[2620]), .Z(n25451) );
  ANDN U14759 ( .B(n9264), .A(n25451), .Z(n17287) );
  NANDN U14760 ( .A(n9265), .B(n17287), .Z(n9266) );
  ANDN U14761 ( .B(y[2621]), .A(x[2621]), .Z(n11935) );
  ANDN U14762 ( .B(n9266), .A(n11935), .Z(n9267) );
  OR U14763 ( .A(n11933), .B(n9267), .Z(n9268) );
  NAND U14764 ( .A(n9269), .B(n9268), .Z(n9270) );
  AND U14765 ( .A(n25467), .B(n9270), .Z(n9271) );
  NANDN U14766 ( .A(n11934), .B(n9271), .Z(n9272) );
  NANDN U14767 ( .A(n25469), .B(n9272), .Z(n9273) );
  NANDN U14768 ( .A(n25472), .B(n9273), .Z(n9274) );
  NANDN U14769 ( .A(x[2626]), .B(y[2626]), .Z(n11932) );
  NANDN U14770 ( .A(x[2627]), .B(y[2627]), .Z(n17305) );
  NAND U14771 ( .A(n11932), .B(n17305), .Z(n25474) );
  ANDN U14772 ( .B(n9274), .A(n25474), .Z(n9275) );
  NANDN U14773 ( .A(y[2627]), .B(x[2627]), .Z(n17302) );
  ANDN U14774 ( .B(x[2628]), .A(y[2628]), .Z(n11930) );
  ANDN U14775 ( .B(n17302), .A(n11930), .Z(n25475) );
  NANDN U14776 ( .A(n9275), .B(n25475), .Z(n9276) );
  AND U14777 ( .A(n25478), .B(n9276), .Z(n9277) );
  NANDN U14778 ( .A(n11925), .B(n9277), .Z(n9280) );
  NANDN U14779 ( .A(y[2629]), .B(x[2629]), .Z(n9279) );
  ANDN U14780 ( .B(x[2631]), .A(y[2631]), .Z(n9282) );
  NANDN U14781 ( .A(y[2630]), .B(x[2630]), .Z(n9278) );
  NANDN U14782 ( .A(n9282), .B(n9278), .Z(n11927) );
  ANDN U14783 ( .B(n9279), .A(n11927), .Z(n25479) );
  NAND U14784 ( .A(n9280), .B(n25479), .Z(n9281) );
  NANDN U14785 ( .A(n11929), .B(n9281), .Z(n9284) );
  ANDN U14786 ( .B(y[2630]), .A(x[2630]), .Z(n11924) );
  NANDN U14787 ( .A(n9282), .B(n11924), .Z(n9283) );
  NANDN U14788 ( .A(n9284), .B(n9283), .Z(n9285) );
  AND U14789 ( .A(n25483), .B(n9285), .Z(n9286) );
  OR U14790 ( .A(n25486), .B(n9286), .Z(n9287) );
  AND U14791 ( .A(n25487), .B(n9287), .Z(n9290) );
  NANDN U14792 ( .A(x[2634]), .B(y[2634]), .Z(n9289) );
  NANDN U14793 ( .A(x[2635]), .B(y[2635]), .Z(n9288) );
  AND U14794 ( .A(n9289), .B(n9288), .Z(n25490) );
  NANDN U14795 ( .A(n9290), .B(n25490), .Z(n9291) );
  NANDN U14796 ( .A(y[2635]), .B(x[2635]), .Z(n17314) );
  ANDN U14797 ( .B(x[2636]), .A(y[2636]), .Z(n11923) );
  ANDN U14798 ( .B(n17314), .A(n11923), .Z(n25491) );
  NAND U14799 ( .A(n9291), .B(n25491), .Z(n9292) );
  NANDN U14800 ( .A(n9293), .B(n9292), .Z(n9294) );
  AND U14801 ( .A(n25495), .B(n9294), .Z(n9296) );
  NANDN U14802 ( .A(x[2638]), .B(y[2638]), .Z(n17320) );
  NANDN U14803 ( .A(x[2639]), .B(y[2639]), .Z(n25498) );
  AND U14804 ( .A(n17320), .B(n25498), .Z(n9295) );
  NANDN U14805 ( .A(n9296), .B(n9295), .Z(n9297) );
  ANDN U14806 ( .B(x[2640]), .A(y[2640]), .Z(n11920) );
  ANDN U14807 ( .B(x[2639]), .A(y[2639]), .Z(n17322) );
  NOR U14808 ( .A(n11920), .B(n17322), .Z(n25501) );
  NAND U14809 ( .A(n9297), .B(n25501), .Z(n9298) );
  NANDN U14810 ( .A(x[2640]), .B(y[2640]), .Z(n17325) );
  NANDN U14811 ( .A(x[2641]), .B(y[2641]), .Z(n11919) );
  NAND U14812 ( .A(n17325), .B(n11919), .Z(n25503) );
  ANDN U14813 ( .B(n9298), .A(n25503), .Z(n9299) );
  OR U14814 ( .A(n25505), .B(n9299), .Z(n9300) );
  AND U14815 ( .A(n25507), .B(n9300), .Z(n9301) );
  NANDN U14816 ( .A(n11918), .B(n9301), .Z(n9302) );
  ANDN U14817 ( .B(x[2644]), .A(y[2644]), .Z(n11916) );
  ANDN U14818 ( .B(n9302), .A(n11916), .Z(n9303) );
  NANDN U14819 ( .A(y[2643]), .B(x[2643]), .Z(n25510) );
  NAND U14820 ( .A(n9303), .B(n25510), .Z(n9304) );
  ANDN U14821 ( .B(y[2644]), .A(x[2644]), .Z(n11917) );
  ANDN U14822 ( .B(n9304), .A(n11917), .Z(n9305) );
  NAND U14823 ( .A(n9306), .B(n9305), .Z(n9307) );
  NAND U14824 ( .A(n11915), .B(n9307), .Z(n9308) );
  ANDN U14825 ( .B(y[2646]), .A(x[2646]), .Z(n17337) );
  ANDN U14826 ( .B(n9308), .A(n17337), .Z(n9311) );
  NANDN U14827 ( .A(y[2646]), .B(x[2646]), .Z(n9310) );
  NANDN U14828 ( .A(y[2647]), .B(x[2647]), .Z(n9309) );
  AND U14829 ( .A(n9310), .B(n9309), .Z(n25517) );
  NANDN U14830 ( .A(n9311), .B(n25517), .Z(n9314) );
  NANDN U14831 ( .A(x[2648]), .B(y[2648]), .Z(n9313) );
  NANDN U14832 ( .A(x[2647]), .B(y[2647]), .Z(n9312) );
  AND U14833 ( .A(n9313), .B(n9312), .Z(n25519) );
  NAND U14834 ( .A(n9314), .B(n25519), .Z(n9317) );
  NANDN U14835 ( .A(y[2648]), .B(x[2648]), .Z(n9316) );
  NANDN U14836 ( .A(y[2649]), .B(x[2649]), .Z(n9315) );
  AND U14837 ( .A(n9316), .B(n9315), .Z(n25522) );
  NAND U14838 ( .A(n9317), .B(n25522), .Z(n9320) );
  NANDN U14839 ( .A(x[2650]), .B(y[2650]), .Z(n9319) );
  NANDN U14840 ( .A(x[2649]), .B(y[2649]), .Z(n9318) );
  AND U14841 ( .A(n9319), .B(n9318), .Z(n25523) );
  NAND U14842 ( .A(n9320), .B(n25523), .Z(n9323) );
  NANDN U14843 ( .A(y[2650]), .B(x[2650]), .Z(n9322) );
  NANDN U14844 ( .A(y[2651]), .B(x[2651]), .Z(n9321) );
  AND U14845 ( .A(n9322), .B(n9321), .Z(n25526) );
  NAND U14846 ( .A(n9323), .B(n25526), .Z(n9324) );
  ANDN U14847 ( .B(y[2651]), .A(x[2651]), .Z(n11914) );
  ANDN U14848 ( .B(n9324), .A(n11914), .Z(n9325) );
  NANDN U14849 ( .A(y[2653]), .B(x[2653]), .Z(n11912) );
  ANDN U14850 ( .B(x[2654]), .A(y[2654]), .Z(n25534) );
  NANDN U14851 ( .A(x[2656]), .B(y[2656]), .Z(n25540) );
  ANDN U14852 ( .B(y[2657]), .A(x[2657]), .Z(n11909) );
  NANDN U14853 ( .A(y[2657]), .B(x[2657]), .Z(n25541) );
  IV U14854 ( .A(y[2658]), .Z(n11905) );
  NANDN U14855 ( .A(y[2660]), .B(x[2660]), .Z(n25549) );
  ANDN U14856 ( .B(x[2659]), .A(y[2659]), .Z(n11906) );
  ANDN U14857 ( .B(y[2661]), .A(x[2661]), .Z(n11902) );
  ANDN U14858 ( .B(y[2660]), .A(x[2660]), .Z(n11904) );
  NOR U14859 ( .A(n11902), .B(n11904), .Z(n25551) );
  ANDN U14860 ( .B(y[2663]), .A(x[2663]), .Z(n17370) );
  ANDN U14861 ( .B(y[2662]), .A(x[2662]), .Z(n11901) );
  NOR U14862 ( .A(n17370), .B(n11901), .Z(n25556) );
  NANDN U14863 ( .A(n9327), .B(n25556), .Z(n9328) );
  AND U14864 ( .A(n25557), .B(n9328), .Z(n9329) );
  NANDN U14865 ( .A(n11899), .B(n9329), .Z(n9330) );
  ANDN U14866 ( .B(y[2665]), .A(x[2665]), .Z(n11897) );
  ANDN U14867 ( .B(n9330), .A(n11897), .Z(n9331) );
  NANDN U14868 ( .A(x[2664]), .B(y[2664]), .Z(n25559) );
  NAND U14869 ( .A(n9331), .B(n25559), .Z(n9332) );
  AND U14870 ( .A(n25565), .B(n9332), .Z(n9333) );
  NANDN U14871 ( .A(n11900), .B(n9333), .Z(n9334) );
  NANDN U14872 ( .A(x[2667]), .B(y[2667]), .Z(n25567) );
  NAND U14873 ( .A(n9334), .B(n25567), .Z(n9335) );
  OR U14874 ( .A(n11898), .B(n9335), .Z(n9336) );
  AND U14875 ( .A(n25569), .B(n9336), .Z(n9337) );
  NANDN U14876 ( .A(x[2668]), .B(y[2668]), .Z(n17378) );
  ANDN U14877 ( .B(y[2669]), .A(x[2669]), .Z(n11894) );
  ANDN U14878 ( .B(n17378), .A(n11894), .Z(n25572) );
  NANDN U14879 ( .A(n9337), .B(n25572), .Z(n9338) );
  NANDN U14880 ( .A(y[2669]), .B(x[2669]), .Z(n11896) );
  NANDN U14881 ( .A(y[2670]), .B(x[2670]), .Z(n17385) );
  AND U14882 ( .A(n11896), .B(n17385), .Z(n25573) );
  NAND U14883 ( .A(n9338), .B(n25573), .Z(n9339) );
  NANDN U14884 ( .A(n25576), .B(n9339), .Z(n9340) );
  OR U14885 ( .A(n17388), .B(n9340), .Z(n9341) );
  AND U14886 ( .A(n9342), .B(n9341), .Z(n9344) );
  NANDN U14887 ( .A(x[2673]), .B(y[2673]), .Z(n25583) );
  ANDN U14888 ( .B(y[2672]), .A(x[2672]), .Z(n17389) );
  ANDN U14889 ( .B(n25583), .A(n17389), .Z(n9343) );
  NANDN U14890 ( .A(n9344), .B(n9343), .Z(n9345) );
  ANDN U14891 ( .B(x[2673]), .A(y[2673]), .Z(n11892) );
  ANDN U14892 ( .B(n9345), .A(n11892), .Z(n9346) );
  NANDN U14893 ( .A(n25585), .B(n9346), .Z(n9352) );
  NANDN U14894 ( .A(x[2675]), .B(y[2675]), .Z(n11891) );
  NANDN U14895 ( .A(x[2674]), .B(y[2674]), .Z(n17392) );
  NAND U14896 ( .A(n11891), .B(n17392), .Z(n9347) );
  NANDN U14897 ( .A(n9348), .B(n9347), .Z(n9351) );
  NANDN U14898 ( .A(x[2677]), .B(y[2677]), .Z(n9350) );
  NANDN U14899 ( .A(x[2676]), .B(y[2676]), .Z(n9349) );
  NAND U14900 ( .A(n9350), .B(n9349), .Z(n17396) );
  ANDN U14901 ( .B(n9351), .A(n17396), .Z(n25587) );
  NAND U14902 ( .A(n9352), .B(n25587), .Z(n9353) );
  AND U14903 ( .A(n25589), .B(n9353), .Z(n9354) );
  ANDN U14904 ( .B(x[2678]), .A(y[2678]), .Z(n11889) );
  ANDN U14905 ( .B(n9354), .A(n11889), .Z(n9355) );
  ANDN U14906 ( .B(n25591), .A(n9355), .Z(n9356) );
  NAND U14907 ( .A(n9357), .B(n9356), .Z(n9358) );
  NAND U14908 ( .A(n9359), .B(n9358), .Z(n9360) );
  ANDN U14909 ( .B(y[2680]), .A(x[2680]), .Z(n11887) );
  ANDN U14910 ( .B(n9360), .A(n11887), .Z(n9361) );
  NANDN U14911 ( .A(x[2681]), .B(y[2681]), .Z(n25600) );
  NAND U14912 ( .A(n9361), .B(n25600), .Z(n9362) );
  NANDN U14913 ( .A(y[2681]), .B(x[2681]), .Z(n17404) );
  XOR U14914 ( .A(x[2682]), .B(y[2682]), .Z(n17409) );
  ANDN U14915 ( .B(n17404), .A(n17409), .Z(n25601) );
  NAND U14916 ( .A(n9362), .B(n25601), .Z(n9363) );
  NANDN U14917 ( .A(n25603), .B(n9363), .Z(n9366) );
  NANDN U14918 ( .A(y[2684]), .B(x[2684]), .Z(n9365) );
  NANDN U14919 ( .A(y[2683]), .B(x[2683]), .Z(n9364) );
  NAND U14920 ( .A(n9365), .B(n9364), .Z(n25606) );
  ANDN U14921 ( .B(n9366), .A(n25606), .Z(n9369) );
  NANDN U14922 ( .A(x[2684]), .B(y[2684]), .Z(n9368) );
  NANDN U14923 ( .A(x[2685]), .B(y[2685]), .Z(n9367) );
  AND U14924 ( .A(n9368), .B(n9367), .Z(n25607) );
  NANDN U14925 ( .A(n9369), .B(n25607), .Z(n9371) );
  NANDN U14926 ( .A(y[2686]), .B(x[2686]), .Z(n9370) );
  ANDN U14927 ( .B(x[2685]), .A(y[2685]), .Z(n25610) );
  ANDN U14928 ( .B(n9370), .A(n25610), .Z(n17413) );
  NAND U14929 ( .A(n9371), .B(n17413), .Z(n9372) );
  NANDN U14930 ( .A(n17415), .B(n9372), .Z(n9373) );
  AND U14931 ( .A(n17417), .B(n9373), .Z(n9376) );
  NANDN U14932 ( .A(x[2688]), .B(y[2688]), .Z(n9375) );
  NANDN U14933 ( .A(x[2689]), .B(y[2689]), .Z(n9374) );
  AND U14934 ( .A(n9375), .B(n9374), .Z(n25623) );
  NANDN U14935 ( .A(n9376), .B(n25623), .Z(n9379) );
  NANDN U14936 ( .A(y[2690]), .B(x[2690]), .Z(n9378) );
  NANDN U14937 ( .A(y[2689]), .B(x[2689]), .Z(n9377) );
  AND U14938 ( .A(n9378), .B(n9377), .Z(n25624) );
  NAND U14939 ( .A(n9379), .B(n25624), .Z(n9382) );
  NANDN U14940 ( .A(x[2690]), .B(y[2690]), .Z(n9381) );
  NANDN U14941 ( .A(x[2691]), .B(y[2691]), .Z(n9380) );
  AND U14942 ( .A(n9381), .B(n9380), .Z(n25626) );
  NAND U14943 ( .A(n9382), .B(n25626), .Z(n9383) );
  AND U14944 ( .A(n25628), .B(n9383), .Z(n9386) );
  NANDN U14945 ( .A(x[2692]), .B(y[2692]), .Z(n25630) );
  ANDN U14946 ( .B(y[2693]), .A(x[2693]), .Z(n17427) );
  IV U14947 ( .A(n17427), .Z(n9384) );
  AND U14948 ( .A(n25630), .B(n9384), .Z(n9385) );
  NANDN U14949 ( .A(n9386), .B(n9385), .Z(n9387) );
  NANDN U14950 ( .A(y[2694]), .B(x[2694]), .Z(n25634) );
  ANDN U14951 ( .B(x[2693]), .A(y[2693]), .Z(n17424) );
  ANDN U14952 ( .B(n25634), .A(n17424), .Z(n25632) );
  NAND U14953 ( .A(n9387), .B(n25632), .Z(n9388) );
  AND U14954 ( .A(n25637), .B(n9388), .Z(n9389) );
  NANDN U14955 ( .A(n17426), .B(n9389), .Z(n9390) );
  ANDN U14956 ( .B(x[2696]), .A(y[2696]), .Z(n11884) );
  ANDN U14957 ( .B(x[2695]), .A(y[2695]), .Z(n17429) );
  NOR U14958 ( .A(n11884), .B(n17429), .Z(n25640) );
  NAND U14959 ( .A(n9390), .B(n25640), .Z(n9391) );
  NANDN U14960 ( .A(x[2696]), .B(y[2696]), .Z(n17432) );
  NANDN U14961 ( .A(x[2697]), .B(y[2697]), .Z(n11883) );
  NAND U14962 ( .A(n17432), .B(n11883), .Z(n25643) );
  ANDN U14963 ( .B(n9391), .A(n25643), .Z(n9392) );
  OR U14964 ( .A(n25645), .B(n9392), .Z(n9393) );
  AND U14965 ( .A(n25647), .B(n9393), .Z(n9394) );
  NANDN U14966 ( .A(y[2699]), .B(x[2699]), .Z(n25648) );
  NANDN U14967 ( .A(n9394), .B(n25648), .Z(n9397) );
  NANDN U14968 ( .A(x[2700]), .B(y[2700]), .Z(n9396) );
  NANDN U14969 ( .A(x[2699]), .B(y[2699]), .Z(n9395) );
  NAND U14970 ( .A(n9396), .B(n9395), .Z(n25650) );
  ANDN U14971 ( .B(n9397), .A(n25650), .Z(n9400) );
  NANDN U14972 ( .A(y[2700]), .B(x[2700]), .Z(n9399) );
  NANDN U14973 ( .A(y[2701]), .B(x[2701]), .Z(n9398) );
  AND U14974 ( .A(n9399), .B(n9398), .Z(n25652) );
  NANDN U14975 ( .A(n9400), .B(n25652), .Z(n9401) );
  NANDN U14976 ( .A(x[2701]), .B(y[2701]), .Z(n25654) );
  NAND U14977 ( .A(n9401), .B(n25654), .Z(n9402) );
  AND U14978 ( .A(n25656), .B(n9402), .Z(n9403) );
  OR U14979 ( .A(n25658), .B(n9403), .Z(n9404) );
  NANDN U14980 ( .A(y[2703]), .B(x[2703]), .Z(n25661) );
  NAND U14981 ( .A(n9404), .B(n25661), .Z(n9406) );
  NANDN U14982 ( .A(x[2704]), .B(y[2704]), .Z(n9405) );
  NANDN U14983 ( .A(x[2705]), .B(y[2705]), .Z(n9407) );
  AND U14984 ( .A(n9405), .B(n9407), .Z(n25664) );
  NAND U14985 ( .A(n9406), .B(n25664), .Z(n9411) );
  ANDN U14986 ( .B(x[2704]), .A(y[2704]), .Z(n25660) );
  NAND U14987 ( .A(n9407), .B(n25660), .Z(n9409) );
  ANDN U14988 ( .B(x[2707]), .A(y[2707]), .Z(n9412) );
  NANDN U14989 ( .A(y[2706]), .B(x[2706]), .Z(n9408) );
  NANDN U14990 ( .A(n9412), .B(n9408), .Z(n25671) );
  ANDN U14991 ( .B(n9409), .A(n25671), .Z(n9410) );
  ANDN U14992 ( .B(x[2705]), .A(y[2705]), .Z(n25666) );
  ANDN U14993 ( .B(n9410), .A(n25666), .Z(n17449) );
  NAND U14994 ( .A(n9411), .B(n17449), .Z(n9414) );
  NANDN U14995 ( .A(x[2707]), .B(y[2707]), .Z(n25672) );
  NANDN U14996 ( .A(x[2706]), .B(y[2706]), .Z(n25668) );
  OR U14997 ( .A(n9412), .B(n25668), .Z(n9413) );
  NAND U14998 ( .A(n25672), .B(n9413), .Z(n17453) );
  ANDN U14999 ( .B(n9414), .A(n17453), .Z(n9415) );
  OR U15000 ( .A(n11882), .B(n9415), .Z(n9416) );
  NAND U15001 ( .A(n9417), .B(n9416), .Z(n9420) );
  NANDN U15002 ( .A(y[2710]), .B(x[2710]), .Z(n9418) );
  NANDN U15003 ( .A(n9419), .B(n9418), .Z(n25681) );
  ANDN U15004 ( .B(n9420), .A(n25681), .Z(n9421) );
  NANDN U15005 ( .A(n11881), .B(n9421), .Z(n9422) );
  NANDN U15006 ( .A(n25683), .B(n9422), .Z(n9423) );
  NANDN U15007 ( .A(y[2713]), .B(x[2713]), .Z(n25685) );
  NAND U15008 ( .A(n9423), .B(n25685), .Z(n9424) );
  OR U15009 ( .A(n17463), .B(n9424), .Z(n9425) );
  NANDN U15010 ( .A(x[2715]), .B(y[2715]), .Z(n20237) );
  ANDN U15011 ( .B(y[2714]), .A(x[2714]), .Z(n17461) );
  ANDN U15012 ( .B(n20237), .A(n17461), .Z(n25686) );
  NAND U15013 ( .A(n9425), .B(n25686), .Z(n9426) );
  NANDN U15014 ( .A(y[2716]), .B(x[2716]), .Z(n20240) );
  NAND U15015 ( .A(n9426), .B(n20240), .Z(n9427) );
  OR U15016 ( .A(n17464), .B(n9427), .Z(n9428) );
  AND U15017 ( .A(n25690), .B(n9428), .Z(n9429) );
  NANDN U15018 ( .A(y[2717]), .B(x[2717]), .Z(n17470) );
  ANDN U15019 ( .B(x[2718]), .A(y[2718]), .Z(n17476) );
  ANDN U15020 ( .B(n17470), .A(n17476), .Z(n25692) );
  NANDN U15021 ( .A(n9429), .B(n25692), .Z(n9431) );
  NANDN U15022 ( .A(x[2718]), .B(y[2718]), .Z(n11875) );
  NANDN U15023 ( .A(x[2719]), .B(y[2719]), .Z(n9430) );
  AND U15024 ( .A(n11875), .B(n9430), .Z(n25694) );
  NAND U15025 ( .A(n9431), .B(n25694), .Z(n9432) );
  NANDN U15026 ( .A(n25697), .B(n9432), .Z(n9436) );
  NANDN U15027 ( .A(x[2721]), .B(y[2721]), .Z(n9433) );
  NANDN U15028 ( .A(n9434), .B(n9433), .Z(n17489) );
  IV U15029 ( .A(x[2720]), .Z(n17481) );
  NAND U15030 ( .A(n17481), .B(y[2720]), .Z(n9435) );
  NANDN U15031 ( .A(n17489), .B(n9435), .Z(n25698) );
  ANDN U15032 ( .B(n9436), .A(n25698), .Z(n9437) );
  OR U15033 ( .A(n25701), .B(n9437), .Z(n9438) );
  ANDN U15034 ( .B(y[2723]), .A(x[2723]), .Z(n25703) );
  ANDN U15035 ( .B(n9438), .A(n25703), .Z(n9439) );
  OR U15036 ( .A(n25705), .B(n9439), .Z(n9440) );
  AND U15037 ( .A(n25706), .B(n9440), .Z(n9441) );
  NANDN U15038 ( .A(y[2725]), .B(x[2725]), .Z(n17500) );
  ANDN U15039 ( .B(x[2726]), .A(y[2726]), .Z(n11872) );
  ANDN U15040 ( .B(n17500), .A(n11872), .Z(n25709) );
  NANDN U15041 ( .A(n9441), .B(n25709), .Z(n9442) );
  AND U15042 ( .A(n25710), .B(n9442), .Z(n9443) );
  ANDN U15043 ( .B(y[2727]), .A(x[2727]), .Z(n17506) );
  ANDN U15044 ( .B(n9443), .A(n17506), .Z(n9444) );
  ANDN U15045 ( .B(x[2727]), .A(y[2727]), .Z(n25712) );
  NOR U15046 ( .A(n9444), .B(n25712), .Z(n9445) );
  NAND U15047 ( .A(n9446), .B(n9445), .Z(n9447) );
  NAND U15048 ( .A(n9448), .B(n9447), .Z(n9449) );
  AND U15049 ( .A(n25721), .B(n9449), .Z(n9450) );
  NANDN U15050 ( .A(n11871), .B(n9450), .Z(n9451) );
  NANDN U15051 ( .A(x[2731]), .B(y[2731]), .Z(n11867) );
  ANDN U15052 ( .B(y[2730]), .A(x[2730]), .Z(n11869) );
  ANDN U15053 ( .B(n11867), .A(n11869), .Z(n25722) );
  NAND U15054 ( .A(n9451), .B(n25722), .Z(n9453) );
  NANDN U15055 ( .A(y[2731]), .B(x[2731]), .Z(n9452) );
  NANDN U15056 ( .A(y[2732]), .B(x[2732]), .Z(n11866) );
  NAND U15057 ( .A(n9452), .B(n11866), .Z(n25724) );
  ANDN U15058 ( .B(n9453), .A(n25724), .Z(n9454) );
  OR U15059 ( .A(n25726), .B(n9454), .Z(n9455) );
  AND U15060 ( .A(n25729), .B(n9455), .Z(n9456) );
  ANDN U15061 ( .B(x[2734]), .A(y[2734]), .Z(n17523) );
  ANDN U15062 ( .B(n9456), .A(n17523), .Z(n9457) );
  ANDN U15063 ( .B(n25730), .A(n9457), .Z(n9458) );
  IV U15064 ( .A(x[2735]), .Z(n11863) );
  NANDN U15065 ( .A(n9458), .B(n11863), .Z(n9461) );
  XOR U15066 ( .A(x[2735]), .B(n9458), .Z(n9459) );
  NAND U15067 ( .A(n9459), .B(y[2735]), .Z(n9460) );
  NAND U15068 ( .A(n9461), .B(n9460), .Z(n9462) );
  ANDN U15069 ( .B(x[2736]), .A(y[2736]), .Z(n11861) );
  ANDN U15070 ( .B(n9462), .A(n11861), .Z(n9464) );
  NANDN U15071 ( .A(x[2737]), .B(y[2737]), .Z(n25738) );
  ANDN U15072 ( .B(y[2736]), .A(x[2736]), .Z(n11865) );
  ANDN U15073 ( .B(n25738), .A(n11865), .Z(n9463) );
  NANDN U15074 ( .A(n9464), .B(n9463), .Z(n9465) );
  ANDN U15075 ( .B(x[2738]), .A(y[2738]), .Z(n25741) );
  ANDN U15076 ( .B(n9465), .A(n25741), .Z(n9466) );
  ANDN U15077 ( .B(x[2737]), .A(y[2737]), .Z(n11862) );
  ANDN U15078 ( .B(n9466), .A(n11862), .Z(n9467) );
  OR U15079 ( .A(n25743), .B(n9467), .Z(n9468) );
  NANDN U15080 ( .A(n25744), .B(n9468), .Z(n9469) );
  NANDN U15081 ( .A(x[2740]), .B(y[2740]), .Z(n25746) );
  NAND U15082 ( .A(n9469), .B(n25746), .Z(n9470) );
  AND U15083 ( .A(n25748), .B(n9470), .Z(n9473) );
  NANDN U15084 ( .A(x[2741]), .B(y[2741]), .Z(n9472) );
  NANDN U15085 ( .A(x[2742]), .B(y[2742]), .Z(n9471) );
  AND U15086 ( .A(n9472), .B(n9471), .Z(n25750) );
  NANDN U15087 ( .A(n9473), .B(n25750), .Z(n9474) );
  NANDN U15088 ( .A(n25753), .B(n9474), .Z(n9475) );
  NANDN U15089 ( .A(x[2743]), .B(y[2743]), .Z(n25754) );
  NAND U15090 ( .A(n9475), .B(n25754), .Z(n9476) );
  AND U15091 ( .A(n25757), .B(n9476), .Z(n9477) );
  NANDN U15092 ( .A(x[2744]), .B(y[2744]), .Z(n17542) );
  IV U15093 ( .A(x[2745]), .Z(n11859) );
  NAND U15094 ( .A(n11859), .B(y[2745]), .Z(n11857) );
  AND U15095 ( .A(n17542), .B(n11857), .Z(n25758) );
  NANDN U15096 ( .A(n9477), .B(n25758), .Z(n9478) );
  ANDN U15097 ( .B(x[2746]), .A(y[2746]), .Z(n11856) );
  NAND U15098 ( .A(n9478), .B(n25760), .Z(n9479) );
  AND U15099 ( .A(n25762), .B(n9479), .Z(n9481) );
  NANDN U15100 ( .A(y[2747]), .B(x[2747]), .Z(n25765) );
  ANDN U15101 ( .B(x[2748]), .A(y[2748]), .Z(n17555) );
  ANDN U15102 ( .B(n25765), .A(n17555), .Z(n9480) );
  NANDN U15103 ( .A(n9481), .B(n9480), .Z(n9482) );
  AND U15104 ( .A(n25766), .B(n9482), .Z(n9483) );
  NAND U15105 ( .A(n9484), .B(n9483), .Z(n9485) );
  NAND U15106 ( .A(n9486), .B(n9485), .Z(n9487) );
  ANDN U15107 ( .B(y[2750]), .A(x[2750]), .Z(n11855) );
  ANDN U15108 ( .B(n9487), .A(n11855), .Z(n9488) );
  NANDN U15109 ( .A(n11850), .B(n9488), .Z(n9489) );
  NANDN U15110 ( .A(y[2752]), .B(x[2752]), .Z(n25776) );
  NAND U15111 ( .A(n9489), .B(n25776), .Z(n9490) );
  OR U15112 ( .A(n11853), .B(n9490), .Z(n9491) );
  AND U15113 ( .A(n25778), .B(n9491), .Z(n9492) );
  NANDN U15114 ( .A(n11851), .B(n9492), .Z(n9493) );
  AND U15115 ( .A(n25780), .B(n9493), .Z(n9495) );
  NANDN U15116 ( .A(x[2754]), .B(y[2754]), .Z(n25783) );
  ANDN U15117 ( .B(y[2755]), .A(x[2755]), .Z(n11848) );
  ANDN U15118 ( .B(n25783), .A(n11848), .Z(n9494) );
  NANDN U15119 ( .A(n9495), .B(n9494), .Z(n9496) );
  AND U15120 ( .A(n25784), .B(n9496), .Z(n9497) );
  NAND U15121 ( .A(n9498), .B(n9497), .Z(n9499) );
  NAND U15122 ( .A(n9500), .B(n9499), .Z(n9501) );
  AND U15123 ( .A(n25792), .B(n9501), .Z(n9502) );
  NANDN U15124 ( .A(n11846), .B(n9502), .Z(n9503) );
  NANDN U15125 ( .A(n25795), .B(n9503), .Z(n9504) );
  ANDN U15126 ( .B(x[2760]), .A(y[2760]), .Z(n11840) );
  ANDN U15127 ( .B(x[2759]), .A(y[2759]), .Z(n11843) );
  NOR U15128 ( .A(n11840), .B(n11843), .Z(n25796) );
  NAND U15129 ( .A(n9504), .B(n25796), .Z(n9505) );
  NANDN U15130 ( .A(x[2761]), .B(y[2761]), .Z(n17578) );
  NANDN U15131 ( .A(x[2760]), .B(y[2760]), .Z(n11842) );
  NAND U15132 ( .A(n17578), .B(n11842), .Z(n25798) );
  ANDN U15133 ( .B(n9505), .A(n25798), .Z(n9506) );
  ANDN U15134 ( .B(x[2762]), .A(y[2762]), .Z(n17580) );
  ANDN U15135 ( .B(x[2761]), .A(y[2761]), .Z(n11839) );
  NOR U15136 ( .A(n17580), .B(n11839), .Z(n25800) );
  NANDN U15137 ( .A(n9506), .B(n25800), .Z(n9507) );
  AND U15138 ( .A(n25803), .B(n9507), .Z(n9508) );
  NANDN U15139 ( .A(n11837), .B(n9508), .Z(n9510) );
  NANDN U15140 ( .A(y[2764]), .B(x[2764]), .Z(n25809) );
  NANDN U15141 ( .A(y[2763]), .B(x[2763]), .Z(n25804) );
  AND U15142 ( .A(n25809), .B(n25804), .Z(n9509) );
  NAND U15143 ( .A(n9510), .B(n9509), .Z(n9511) );
  NANDN U15144 ( .A(x[2765]), .B(y[2765]), .Z(n25810) );
  NAND U15145 ( .A(n9511), .B(n25810), .Z(n9512) );
  OR U15146 ( .A(n11838), .B(n9512), .Z(n9514) );
  NANDN U15147 ( .A(y[2766]), .B(x[2766]), .Z(n9513) );
  NANDN U15148 ( .A(y[2765]), .B(x[2765]), .Z(n11836) );
  NAND U15149 ( .A(n9513), .B(n11836), .Z(n25812) );
  ANDN U15150 ( .B(n9514), .A(n25812), .Z(n9515) );
  OR U15151 ( .A(n25815), .B(n9515), .Z(n9516) );
  NANDN U15152 ( .A(n25817), .B(n9516), .Z(n9517) );
  NANDN U15153 ( .A(n25819), .B(n9517), .Z(n9518) );
  ANDN U15154 ( .B(x[2770]), .A(y[2770]), .Z(n17600) );
  ANDN U15155 ( .B(n9518), .A(n17600), .Z(n9519) );
  NANDN U15156 ( .A(y[2769]), .B(x[2769]), .Z(n25821) );
  NAND U15157 ( .A(n9519), .B(n25821), .Z(n9521) );
  NANDN U15158 ( .A(x[2770]), .B(y[2770]), .Z(n9520) );
  ANDN U15159 ( .B(y[2771]), .A(x[2771]), .Z(n17601) );
  ANDN U15160 ( .B(n9520), .A(n17601), .Z(n25822) );
  NAND U15161 ( .A(n9521), .B(n25822), .Z(n9524) );
  NANDN U15162 ( .A(y[2772]), .B(x[2772]), .Z(n9523) );
  NANDN U15163 ( .A(y[2771]), .B(x[2771]), .Z(n9522) );
  NAND U15164 ( .A(n9523), .B(n9522), .Z(n17603) );
  ANDN U15165 ( .B(n9524), .A(n17603), .Z(n9527) );
  NANDN U15166 ( .A(x[2772]), .B(y[2772]), .Z(n9526) );
  NANDN U15167 ( .A(x[2773]), .B(y[2773]), .Z(n9525) );
  AND U15168 ( .A(n9526), .B(n9525), .Z(n25827) );
  NANDN U15169 ( .A(n9527), .B(n25827), .Z(n9530) );
  NANDN U15170 ( .A(y[2774]), .B(x[2774]), .Z(n9529) );
  NANDN U15171 ( .A(y[2773]), .B(x[2773]), .Z(n9528) );
  AND U15172 ( .A(n9529), .B(n9528), .Z(n25828) );
  NAND U15173 ( .A(n9530), .B(n25828), .Z(n9533) );
  NANDN U15174 ( .A(x[2775]), .B(y[2775]), .Z(n9532) );
  NANDN U15175 ( .A(x[2774]), .B(y[2774]), .Z(n9531) );
  AND U15176 ( .A(n9532), .B(n9531), .Z(n25831) );
  NAND U15177 ( .A(n9533), .B(n25831), .Z(n9534) );
  ANDN U15178 ( .B(x[2776]), .A(y[2776]), .Z(n20235) );
  NANDN U15179 ( .A(y[2775]), .B(x[2775]), .Z(n25832) );
  NANDN U15180 ( .A(n20235), .B(n25832), .Z(n17608) );
  ANDN U15181 ( .B(n9534), .A(n17608), .Z(n9536) );
  NANDN U15182 ( .A(x[2776]), .B(y[2776]), .Z(n9535) );
  ANDN U15183 ( .B(y[2777]), .A(x[2777]), .Z(n20236) );
  ANDN U15184 ( .B(n9535), .A(n20236), .Z(n25835) );
  NANDN U15185 ( .A(n9536), .B(n25835), .Z(n9539) );
  NANDN U15186 ( .A(y[2778]), .B(x[2778]), .Z(n9538) );
  NANDN U15187 ( .A(y[2777]), .B(x[2777]), .Z(n9537) );
  AND U15188 ( .A(n9538), .B(n9537), .Z(n25838) );
  NAND U15189 ( .A(n9539), .B(n25838), .Z(n9542) );
  NANDN U15190 ( .A(x[2778]), .B(y[2778]), .Z(n9541) );
  NANDN U15191 ( .A(x[2779]), .B(y[2779]), .Z(n9540) );
  AND U15192 ( .A(n9541), .B(n9540), .Z(n25841) );
  NAND U15193 ( .A(n9542), .B(n25841), .Z(n9543) );
  AND U15194 ( .A(n25842), .B(n9543), .Z(n9546) );
  NANDN U15195 ( .A(x[2780]), .B(y[2780]), .Z(n9545) );
  NANDN U15196 ( .A(x[2781]), .B(y[2781]), .Z(n9544) );
  AND U15197 ( .A(n9545), .B(n9544), .Z(n25844) );
  NANDN U15198 ( .A(n9546), .B(n25844), .Z(n9549) );
  XNOR U15199 ( .A(y[2782]), .B(x[2782]), .Z(n9548) );
  NANDN U15200 ( .A(y[2781]), .B(x[2781]), .Z(n9547) );
  AND U15201 ( .A(n9548), .B(n9547), .Z(n25846) );
  NAND U15202 ( .A(n9549), .B(n25846), .Z(n9554) );
  ANDN U15203 ( .B(y[2784]), .A(x[2784]), .Z(n9551) );
  ANDN U15204 ( .B(y[2782]), .A(x[2782]), .Z(n9550) );
  NOR U15205 ( .A(n9551), .B(n9550), .Z(n9553) );
  NANDN U15206 ( .A(x[2783]), .B(y[2783]), .Z(n9552) );
  AND U15207 ( .A(n9553), .B(n9552), .Z(n25849) );
  NAND U15208 ( .A(n9554), .B(n25849), .Z(n9559) );
  NANDN U15209 ( .A(x[2784]), .B(y[2784]), .Z(n9558) );
  XNOR U15210 ( .A(x[2784]), .B(y[2784]), .Z(n9556) );
  NANDN U15211 ( .A(y[2783]), .B(x[2783]), .Z(n9555) );
  NAND U15212 ( .A(n9556), .B(n9555), .Z(n9557) );
  AND U15213 ( .A(n9558), .B(n9557), .Z(n17618) );
  ANDN U15214 ( .B(n9559), .A(n17618), .Z(n9560) );
  IV U15215 ( .A(y[2785]), .Z(n17617) );
  NANDN U15216 ( .A(n9560), .B(n17617), .Z(n9563) );
  XOR U15217 ( .A(y[2785]), .B(n9560), .Z(n9561) );
  NAND U15218 ( .A(n9561), .B(x[2785]), .Z(n9562) );
  NAND U15219 ( .A(n9563), .B(n9562), .Z(n9564) );
  ANDN U15220 ( .B(y[2786]), .A(x[2786]), .Z(n11830) );
  ANDN U15221 ( .B(n9564), .A(n11830), .Z(n9565) );
  NANDN U15222 ( .A(y[2786]), .B(x[2786]), .Z(n25854) );
  ANDN U15223 ( .B(x[2787]), .A(y[2787]), .Z(n25859) );
  ANDN U15224 ( .B(n25854), .A(n25859), .Z(n17622) );
  NANDN U15225 ( .A(n9565), .B(n17622), .Z(n9567) );
  NANDN U15226 ( .A(x[2788]), .B(y[2788]), .Z(n9566) );
  NANDN U15227 ( .A(x[2787]), .B(y[2787]), .Z(n25856) );
  NAND U15228 ( .A(n9566), .B(n25856), .Z(n17624) );
  ANDN U15229 ( .B(n9567), .A(n17624), .Z(n9569) );
  IV U15230 ( .A(y[2788]), .Z(n25860) );
  NAND U15231 ( .A(n25860), .B(x[2788]), .Z(n9568) );
  ANDN U15232 ( .B(x[2789]), .A(y[2789]), .Z(n25866) );
  ANDN U15233 ( .B(n9568), .A(n25866), .Z(n17626) );
  NANDN U15234 ( .A(n9569), .B(n17626), .Z(n9570) );
  NANDN U15235 ( .A(n25868), .B(n9570), .Z(n9573) );
  NANDN U15236 ( .A(y[2790]), .B(x[2790]), .Z(n9572) );
  NANDN U15237 ( .A(y[2791]), .B(x[2791]), .Z(n9571) );
  AND U15238 ( .A(n9572), .B(n9571), .Z(n25869) );
  NAND U15239 ( .A(n9573), .B(n25869), .Z(n9576) );
  NANDN U15240 ( .A(x[2792]), .B(y[2792]), .Z(n9575) );
  NANDN U15241 ( .A(x[2791]), .B(y[2791]), .Z(n9574) );
  NAND U15242 ( .A(n9575), .B(n9574), .Z(n25872) );
  ANDN U15243 ( .B(n9576), .A(n25872), .Z(n9579) );
  NANDN U15244 ( .A(y[2792]), .B(x[2792]), .Z(n9578) );
  NANDN U15245 ( .A(y[2793]), .B(x[2793]), .Z(n9577) );
  AND U15246 ( .A(n9578), .B(n9577), .Z(n25873) );
  NANDN U15247 ( .A(n9579), .B(n25873), .Z(n9580) );
  AND U15248 ( .A(n25876), .B(n9580), .Z(n9581) );
  NANDN U15249 ( .A(y[2794]), .B(x[2794]), .Z(n25877) );
  NANDN U15250 ( .A(n9581), .B(n25877), .Z(n9582) );
  NANDN U15251 ( .A(x[2794]), .B(y[2794]), .Z(n17633) );
  NANDN U15252 ( .A(x[2795]), .B(y[2795]), .Z(n11828) );
  NAND U15253 ( .A(n17633), .B(n11828), .Z(n25879) );
  ANDN U15254 ( .B(n9582), .A(n25879), .Z(n9583) );
  OR U15255 ( .A(n25881), .B(n9583), .Z(n9584) );
  AND U15256 ( .A(n25884), .B(n9584), .Z(n9585) );
  ANDN U15257 ( .B(y[2797]), .A(x[2797]), .Z(n17644) );
  ANDN U15258 ( .B(n9585), .A(n17644), .Z(n9586) );
  ANDN U15259 ( .B(n25885), .A(n9586), .Z(n9587) );
  NAND U15260 ( .A(n9588), .B(n9587), .Z(n9589) );
  NAND U15261 ( .A(n9590), .B(n9589), .Z(n9591) );
  AND U15262 ( .A(n25893), .B(n9591), .Z(n9592) );
  NANDN U15263 ( .A(n11827), .B(n9592), .Z(n9593) );
  NANDN U15264 ( .A(x[2801]), .B(y[2801]), .Z(n17655) );
  ANDN U15265 ( .B(y[2800]), .A(x[2800]), .Z(n17647) );
  ANDN U15266 ( .B(n17655), .A(n17647), .Z(n25896) );
  NAND U15267 ( .A(n9593), .B(n25896), .Z(n9594) );
  AND U15268 ( .A(n25897), .B(n9594), .Z(n9595) );
  OR U15269 ( .A(n25900), .B(n9595), .Z(n9596) );
  AND U15270 ( .A(n25901), .B(n9596), .Z(n9597) );
  ANDN U15271 ( .B(x[2804]), .A(y[2804]), .Z(n11824) );
  ANDN U15272 ( .B(n9597), .A(n11824), .Z(n9598) );
  ANDN U15273 ( .B(n25903), .A(n9598), .Z(n9599) );
  NAND U15274 ( .A(n9600), .B(n9599), .Z(n9601) );
  NAND U15275 ( .A(n9602), .B(n9601), .Z(n9603) );
  AND U15276 ( .A(n25911), .B(n9603), .Z(n9604) );
  NANDN U15277 ( .A(n11822), .B(n9604), .Z(n9606) );
  XNOR U15278 ( .A(x[2808]), .B(y[2808]), .Z(n9605) );
  ANDN U15279 ( .B(x[2807]), .A(y[2807]), .Z(n11820) );
  ANDN U15280 ( .B(n9605), .A(n11820), .Z(n25913) );
  NAND U15281 ( .A(n9606), .B(n25913), .Z(n9608) );
  IV U15282 ( .A(x[2808]), .Z(n11819) );
  NAND U15283 ( .A(n11819), .B(y[2808]), .Z(n9607) );
  ANDN U15284 ( .B(y[2809]), .A(x[2809]), .Z(n11816) );
  ANDN U15285 ( .B(n9607), .A(n11816), .Z(n25916) );
  NAND U15286 ( .A(n9608), .B(n25916), .Z(n9609) );
  AND U15287 ( .A(n25917), .B(n9609), .Z(n9611) );
  NANDN U15288 ( .A(x[2811]), .B(y[2811]), .Z(n11810) );
  ANDN U15289 ( .B(y[2810]), .A(x[2810]), .Z(n25919) );
  ANDN U15290 ( .B(n11810), .A(n25919), .Z(n9610) );
  NANDN U15291 ( .A(n9611), .B(n9610), .Z(n9615) );
  NANDN U15292 ( .A(y[2811]), .B(x[2811]), .Z(n9614) );
  NANDN U15293 ( .A(y[2812]), .B(x[2812]), .Z(n9612) );
  NANDN U15294 ( .A(n9613), .B(n9612), .Z(n11812) );
  ANDN U15295 ( .B(n9614), .A(n11812), .Z(n25921) );
  NAND U15296 ( .A(n9615), .B(n25921), .Z(n9618) );
  NANDN U15297 ( .A(x[2814]), .B(y[2814]), .Z(n9617) );
  NANDN U15298 ( .A(x[2813]), .B(y[2813]), .Z(n9616) );
  NAND U15299 ( .A(n9617), .B(n9616), .Z(n11813) );
  ANDN U15300 ( .B(n9618), .A(n11813), .Z(n9619) );
  NAND U15301 ( .A(n9620), .B(n9619), .Z(n9622) );
  NANDN U15302 ( .A(y[2815]), .B(x[2815]), .Z(n9621) );
  ANDN U15303 ( .B(x[2814]), .A(y[2814]), .Z(n25926) );
  ANDN U15304 ( .B(n9621), .A(n25926), .Z(n17676) );
  NAND U15305 ( .A(n9622), .B(n17676), .Z(n9625) );
  IV U15306 ( .A(x[2815]), .Z(n25929) );
  NAND U15307 ( .A(n25929), .B(y[2815]), .Z(n9624) );
  NANDN U15308 ( .A(x[2816]), .B(y[2816]), .Z(n9623) );
  NAND U15309 ( .A(n9624), .B(n9623), .Z(n17679) );
  ANDN U15310 ( .B(n9625), .A(n17679), .Z(n9626) );
  ANDN U15311 ( .B(x[2817]), .A(y[2817]), .Z(n25939) );
  NANDN U15312 ( .A(n9626), .B(n17680), .Z(n9627) );
  ANDN U15313 ( .B(y[2817]), .A(x[2817]), .Z(n17682) );
  ANDN U15314 ( .B(n9627), .A(n17682), .Z(n9628) );
  OR U15315 ( .A(n17684), .B(n9628), .Z(n9629) );
  NAND U15316 ( .A(n9630), .B(n9629), .Z(n9631) );
  ANDN U15317 ( .B(x[2819]), .A(y[2819]), .Z(n17685) );
  ANDN U15318 ( .B(n9631), .A(n17685), .Z(n9632) );
  NANDN U15319 ( .A(n17688), .B(n9632), .Z(n9633) );
  NANDN U15320 ( .A(x[2821]), .B(y[2821]), .Z(n25948) );
  NAND U15321 ( .A(n9633), .B(n25948), .Z(n9634) );
  OR U15322 ( .A(n11808), .B(n9634), .Z(n9635) );
  AND U15323 ( .A(n25950), .B(n9635), .Z(n9636) );
  ANDN U15324 ( .B(x[2821]), .A(y[2821]), .Z(n17689) );
  ANDN U15325 ( .B(n9636), .A(n17689), .Z(n9637) );
  NANDN U15326 ( .A(x[2822]), .B(y[2822]), .Z(n17691) );
  ANDN U15327 ( .B(y[2823]), .A(x[2823]), .Z(n11805) );
  ANDN U15328 ( .B(n17691), .A(n11805), .Z(n25953) );
  NANDN U15329 ( .A(n9637), .B(n25953), .Z(n9638) );
  NANDN U15330 ( .A(y[2824]), .B(x[2824]), .Z(n17698) );
  ANDN U15331 ( .B(x[2823]), .A(y[2823]), .Z(n11806) );
  ANDN U15332 ( .B(n17698), .A(n11806), .Z(n25954) );
  NAND U15333 ( .A(n9638), .B(n25954), .Z(n9639) );
  NANDN U15334 ( .A(n25956), .B(n9639), .Z(n9640) );
  AND U15335 ( .A(n25958), .B(n9640), .Z(n9643) );
  NANDN U15336 ( .A(x[2825]), .B(y[2825]), .Z(n9642) );
  NANDN U15337 ( .A(x[2826]), .B(y[2826]), .Z(n9641) );
  AND U15338 ( .A(n9642), .B(n9641), .Z(n25960) );
  NANDN U15339 ( .A(n9643), .B(n25960), .Z(n9646) );
  NANDN U15340 ( .A(y[2827]), .B(x[2827]), .Z(n9645) );
  NANDN U15341 ( .A(y[2826]), .B(x[2826]), .Z(n9644) );
  AND U15342 ( .A(n9645), .B(n9644), .Z(n25962) );
  NAND U15343 ( .A(n9646), .B(n25962), .Z(n9647) );
  AND U15344 ( .A(n25964), .B(n9647), .Z(n9648) );
  NAND U15345 ( .A(n9649), .B(n9648), .Z(n9650) );
  NAND U15346 ( .A(n9651), .B(n9650), .Z(n9652) );
  ANDN U15347 ( .B(y[2830]), .A(x[2830]), .Z(n25979) );
  ANDN U15348 ( .B(y[2829]), .A(x[2829]), .Z(n25968) );
  NOR U15349 ( .A(n25979), .B(n25968), .Z(n17707) );
  NAND U15350 ( .A(n9652), .B(n17707), .Z(n9653) );
  AND U15351 ( .A(n17709), .B(n9653), .Z(n9654) );
  OR U15352 ( .A(n17711), .B(n9654), .Z(n9655) );
  ANDN U15353 ( .B(x[2832]), .A(y[2832]), .Z(n11802) );
  NANDN U15354 ( .A(x[2833]), .B(y[2833]), .Z(n25987) );
  NANDN U15355 ( .A(x[2832]), .B(y[2832]), .Z(n25982) );
  NANDN U15356 ( .A(x[2834]), .B(y[2834]), .Z(n17715) );
  NANDN U15357 ( .A(x[2835]), .B(y[2835]), .Z(n11800) );
  NAND U15358 ( .A(n17715), .B(n11800), .Z(n25990) );
  NANDN U15359 ( .A(y[2835]), .B(x[2835]), .Z(n9656) );
  ANDN U15360 ( .B(x[2836]), .A(y[2836]), .Z(n17723) );
  ANDN U15361 ( .B(n9656), .A(n17723), .Z(n25992) );
  IV U15362 ( .A(y[2837]), .Z(n17724) );
  NAND U15363 ( .A(n17724), .B(x[2837]), .Z(n9657) );
  ANDN U15364 ( .B(x[2838]), .A(y[2838]), .Z(n17730) );
  ANDN U15365 ( .B(n9657), .A(n17730), .Z(n25996) );
  NANDN U15366 ( .A(y[2839]), .B(x[2839]), .Z(n26000) );
  XNOR U15367 ( .A(x[2842]), .B(y[2842]), .Z(n26008) );
  ANDN U15368 ( .B(x[2841]), .A(y[2841]), .Z(n17736) );
  NANDN U15369 ( .A(x[2842]), .B(y[2842]), .Z(n9659) );
  NANDN U15370 ( .A(x[2843]), .B(y[2843]), .Z(n9658) );
  NAND U15371 ( .A(n9659), .B(n9658), .Z(n26010) );
  NANDN U15372 ( .A(y[2843]), .B(x[2843]), .Z(n9661) );
  NANDN U15373 ( .A(y[2844]), .B(x[2844]), .Z(n9660) );
  AND U15374 ( .A(n9661), .B(n9660), .Z(n26012) );
  NANDN U15375 ( .A(n9662), .B(n26012), .Z(n9665) );
  NANDN U15376 ( .A(x[2845]), .B(y[2845]), .Z(n9664) );
  NANDN U15377 ( .A(x[2844]), .B(y[2844]), .Z(n9663) );
  NAND U15378 ( .A(n9664), .B(n9663), .Z(n26014) );
  ANDN U15379 ( .B(n9665), .A(n26014), .Z(n9668) );
  NANDN U15380 ( .A(y[2846]), .B(x[2846]), .Z(n9667) );
  NANDN U15381 ( .A(y[2845]), .B(x[2845]), .Z(n9666) );
  AND U15382 ( .A(n9667), .B(n9666), .Z(n26016) );
  NANDN U15383 ( .A(n9668), .B(n26016), .Z(n9669) );
  AND U15384 ( .A(n26019), .B(n9669), .Z(n9670) );
  NANDN U15385 ( .A(n11798), .B(n9670), .Z(n9672) );
  NANDN U15386 ( .A(y[2848]), .B(x[2848]), .Z(n26025) );
  NANDN U15387 ( .A(y[2847]), .B(x[2847]), .Z(n26020) );
  AND U15388 ( .A(n26025), .B(n26020), .Z(n9671) );
  NAND U15389 ( .A(n9672), .B(n9671), .Z(n9673) );
  NANDN U15390 ( .A(x[2849]), .B(y[2849]), .Z(n26026) );
  NAND U15391 ( .A(n9673), .B(n26026), .Z(n9674) );
  OR U15392 ( .A(n11799), .B(n9674), .Z(n9675) );
  NANDN U15393 ( .A(n26028), .B(n9675), .Z(n9676) );
  NANDN U15394 ( .A(n26031), .B(n9676), .Z(n9677) );
  NANDN U15395 ( .A(n26033), .B(n9677), .Z(n9678) );
  ANDN U15396 ( .B(y[2853]), .A(x[2853]), .Z(n11794) );
  ANDN U15397 ( .B(n9678), .A(n11794), .Z(n9679) );
  NANDN U15398 ( .A(x[2852]), .B(y[2852]), .Z(n26034) );
  NAND U15399 ( .A(n9679), .B(n26034), .Z(n9680) );
  NANDN U15400 ( .A(y[2853]), .B(x[2853]), .Z(n26036) );
  NAND U15401 ( .A(n9680), .B(n26036), .Z(n9681) );
  NANDN U15402 ( .A(n9681), .B(y[2854]), .Z(n9684) );
  IV U15403 ( .A(x[2854]), .Z(n11793) );
  XNOR U15404 ( .A(n9681), .B(y[2854]), .Z(n9682) );
  NAND U15405 ( .A(n11793), .B(n9682), .Z(n9683) );
  NAND U15406 ( .A(n9684), .B(n9683), .Z(n9685) );
  NANDN U15407 ( .A(x[2855]), .B(y[2855]), .Z(n26042) );
  NANDN U15408 ( .A(n9685), .B(n26042), .Z(n9686) );
  ANDN U15409 ( .B(x[2855]), .A(y[2855]), .Z(n11792) );
  NANDN U15410 ( .A(y[2856]), .B(x[2856]), .Z(n26044) );
  NANDN U15411 ( .A(x[2857]), .B(y[2857]), .Z(n9688) );
  NANDN U15412 ( .A(x[2856]), .B(y[2856]), .Z(n9687) );
  AND U15413 ( .A(n9688), .B(n9687), .Z(n26046) );
  NANDN U15414 ( .A(y[2857]), .B(x[2857]), .Z(n26050) );
  ANDN U15415 ( .B(x[2858]), .A(y[2858]), .Z(n26048) );
  ANDN U15416 ( .B(x[2859]), .A(y[2859]), .Z(n26054) );
  NOR U15417 ( .A(n26048), .B(n26054), .Z(n17769) );
  NANDN U15418 ( .A(x[2860]), .B(y[2860]), .Z(n9690) );
  NANDN U15419 ( .A(x[2859]), .B(y[2859]), .Z(n9689) );
  AND U15420 ( .A(n9690), .B(n9689), .Z(n26056) );
  NANDN U15421 ( .A(y[2860]), .B(x[2860]), .Z(n9692) );
  NANDN U15422 ( .A(y[2861]), .B(x[2861]), .Z(n9691) );
  AND U15423 ( .A(n9692), .B(n9691), .Z(n26058) );
  ANDN U15424 ( .B(y[2862]), .A(x[2862]), .Z(n17774) );
  NANDN U15425 ( .A(y[2864]), .B(x[2864]), .Z(n26066) );
  ANDN U15426 ( .B(x[2863]), .A(y[2863]), .Z(n17777) );
  ANDN U15427 ( .B(y[2865]), .A(x[2865]), .Z(n11789) );
  ANDN U15428 ( .B(y[2864]), .A(x[2864]), .Z(n11790) );
  NOR U15429 ( .A(n11789), .B(n11790), .Z(n26068) );
  ANDN U15430 ( .B(y[2866]), .A(x[2866]), .Z(n11788) );
  ANDN U15431 ( .B(y[2868]), .A(x[2868]), .Z(n9694) );
  NANDN U15432 ( .A(x[2867]), .B(y[2867]), .Z(n9693) );
  NANDN U15433 ( .A(n9694), .B(n9693), .Z(n17789) );
  NOR U15434 ( .A(n11788), .B(n17789), .Z(n26072) );
  NANDN U15435 ( .A(y[2868]), .B(x[2868]), .Z(n17790) );
  NANDN U15436 ( .A(y[2867]), .B(x[2867]), .Z(n11786) );
  OR U15437 ( .A(n9694), .B(n11786), .Z(n9695) );
  NAND U15438 ( .A(n17790), .B(n9695), .Z(n26074) );
  AND U15439 ( .A(n9697), .B(n9696), .Z(n9698) );
  OR U15440 ( .A(n26082), .B(n9698), .Z(n9700) );
  NANDN U15441 ( .A(y[2871]), .B(x[2871]), .Z(n9699) );
  NANDN U15442 ( .A(y[2872]), .B(x[2872]), .Z(n11783) );
  NAND U15443 ( .A(n9699), .B(n11783), .Z(n26085) );
  ANDN U15444 ( .B(n9700), .A(n26085), .Z(n9702) );
  NANDN U15445 ( .A(x[2872]), .B(y[2872]), .Z(n9701) );
  ANDN U15446 ( .B(y[2873]), .A(x[2873]), .Z(n11782) );
  ANDN U15447 ( .B(n9701), .A(n11782), .Z(n26086) );
  NANDN U15448 ( .A(n9702), .B(n26086), .Z(n9704) );
  NANDN U15449 ( .A(y[2873]), .B(x[2873]), .Z(n26088) );
  ANDN U15450 ( .B(x[2874]), .A(y[2874]), .Z(n11781) );
  ANDN U15451 ( .B(n26088), .A(n11781), .Z(n9703) );
  NAND U15452 ( .A(n9704), .B(n9703), .Z(n9705) );
  ANDN U15453 ( .B(y[2874]), .A(x[2874]), .Z(n26091) );
  ANDN U15454 ( .B(n9705), .A(n26091), .Z(n9706) );
  IV U15455 ( .A(x[2875]), .Z(n17808) );
  NANDN U15456 ( .A(n9706), .B(n17808), .Z(n9709) );
  XOR U15457 ( .A(x[2875]), .B(n9706), .Z(n9707) );
  NAND U15458 ( .A(n9707), .B(y[2875]), .Z(n9708) );
  NAND U15459 ( .A(n9709), .B(n9708), .Z(n9710) );
  AND U15460 ( .A(n26096), .B(n9710), .Z(n9712) );
  NANDN U15461 ( .A(x[2877]), .B(y[2877]), .Z(n26098) );
  ANDN U15462 ( .B(y[2876]), .A(x[2876]), .Z(n17810) );
  ANDN U15463 ( .B(n26098), .A(n17810), .Z(n9711) );
  NANDN U15464 ( .A(n9712), .B(n9711), .Z(n9713) );
  AND U15465 ( .A(n26100), .B(n9713), .Z(n9715) );
  NANDN U15466 ( .A(x[2878]), .B(y[2878]), .Z(n9714) );
  ANDN U15467 ( .B(y[2879]), .A(x[2879]), .Z(n11777) );
  ANDN U15468 ( .B(n9714), .A(n11777), .Z(n26103) );
  NANDN U15469 ( .A(n9715), .B(n26103), .Z(n9716) );
  NANDN U15470 ( .A(y[2879]), .B(x[2879]), .Z(n11779) );
  NANDN U15471 ( .A(y[2880]), .B(x[2880]), .Z(n17823) );
  AND U15472 ( .A(n11779), .B(n17823), .Z(n26104) );
  NAND U15473 ( .A(n9716), .B(n26104), .Z(n9717) );
  NANDN U15474 ( .A(n11776), .B(n9717), .Z(n9718) );
  OR U15475 ( .A(n26107), .B(n9718), .Z(n9719) );
  AND U15476 ( .A(n9720), .B(n9719), .Z(n9722) );
  NANDN U15477 ( .A(x[2883]), .B(y[2883]), .Z(n26114) );
  ANDN U15478 ( .B(y[2882]), .A(x[2882]), .Z(n11775) );
  ANDN U15479 ( .B(n26114), .A(n11775), .Z(n9721) );
  NANDN U15480 ( .A(n9722), .B(n9721), .Z(n9723) );
  ANDN U15481 ( .B(x[2883]), .A(y[2883]), .Z(n11773) );
  ANDN U15482 ( .B(n9723), .A(n11773), .Z(n9724) );
  NANDN U15483 ( .A(n26116), .B(n9724), .Z(n9730) );
  ANDN U15484 ( .B(y[2885]), .A(x[2885]), .Z(n17830) );
  NANDN U15485 ( .A(x[2884]), .B(y[2884]), .Z(n11772) );
  NANDN U15486 ( .A(n17830), .B(n11772), .Z(n9725) );
  NANDN U15487 ( .A(n9726), .B(n9725), .Z(n9729) );
  NANDN U15488 ( .A(x[2887]), .B(y[2887]), .Z(n9728) );
  NANDN U15489 ( .A(x[2886]), .B(y[2886]), .Z(n9727) );
  NAND U15490 ( .A(n9728), .B(n9727), .Z(n17832) );
  ANDN U15491 ( .B(n9729), .A(n17832), .Z(n26118) );
  NAND U15492 ( .A(n9730), .B(n26118), .Z(n9731) );
  AND U15493 ( .A(n26120), .B(n9731), .Z(n9732) );
  ANDN U15494 ( .B(x[2888]), .A(y[2888]), .Z(n17838) );
  ANDN U15495 ( .B(n9732), .A(n17838), .Z(n9733) );
  ANDN U15496 ( .B(n26122), .A(n9733), .Z(n9734) );
  NAND U15497 ( .A(n9735), .B(n9734), .Z(n9736) );
  NAND U15498 ( .A(n9737), .B(n9736), .Z(n9738) );
  AND U15499 ( .A(n26131), .B(n9738), .Z(n9739) );
  NANDN U15500 ( .A(n11771), .B(n9739), .Z(n9740) );
  ANDN U15501 ( .B(x[2892]), .A(y[2892]), .Z(n11766) );
  ANDN U15502 ( .B(x[2891]), .A(y[2891]), .Z(n11769) );
  NOR U15503 ( .A(n11766), .B(n11769), .Z(n26132) );
  NAND U15504 ( .A(n9740), .B(n26132), .Z(n9741) );
  NANDN U15505 ( .A(x[2892]), .B(y[2892]), .Z(n11768) );
  NANDN U15506 ( .A(x[2893]), .B(y[2893]), .Z(n11765) );
  NAND U15507 ( .A(n11768), .B(n11765), .Z(n26134) );
  ANDN U15508 ( .B(n9741), .A(n26134), .Z(n9742) );
  NANDN U15509 ( .A(y[2894]), .B(x[2894]), .Z(n17850) );
  ANDN U15510 ( .B(x[2893]), .A(y[2893]), .Z(n11767) );
  ANDN U15511 ( .B(n17850), .A(n11767), .Z(n26136) );
  NANDN U15512 ( .A(n9742), .B(n26136), .Z(n9743) );
  AND U15513 ( .A(n26139), .B(n9743), .Z(n9744) );
  ANDN U15514 ( .B(y[2895]), .A(x[2895]), .Z(n17854) );
  ANDN U15515 ( .B(n9744), .A(n17854), .Z(n9745) );
  ANDN U15516 ( .B(n26140), .A(n9745), .Z(n9746) );
  NAND U15517 ( .A(n9747), .B(n9746), .Z(n9748) );
  NAND U15518 ( .A(n9749), .B(n9748), .Z(n9750) );
  AND U15519 ( .A(n26148), .B(n9750), .Z(n9751) );
  NANDN U15520 ( .A(n11764), .B(n9751), .Z(n9752) );
  NANDN U15521 ( .A(n26150), .B(n9752), .Z(n9753) );
  AND U15522 ( .A(n26152), .B(n9753), .Z(n9755) );
  NANDN U15523 ( .A(x[2900]), .B(y[2900]), .Z(n9754) );
  ANDN U15524 ( .B(y[2901]), .A(x[2901]), .Z(n11762) );
  ANDN U15525 ( .B(n9754), .A(n11762), .Z(n26154) );
  NANDN U15526 ( .A(n9755), .B(n26154), .Z(n9756) );
  AND U15527 ( .A(n26156), .B(n9756), .Z(n9757) );
  ANDN U15528 ( .B(x[2902]), .A(y[2902]), .Z(n11760) );
  ANDN U15529 ( .B(n9757), .A(n11760), .Z(n9758) );
  ANDN U15530 ( .B(n26158), .A(n9758), .Z(n9759) );
  NAND U15531 ( .A(n9760), .B(n9759), .Z(n9761) );
  NAND U15532 ( .A(n9762), .B(n9761), .Z(n9765) );
  ANDN U15533 ( .B(y[2907]), .A(x[2907]), .Z(n11755) );
  NANDN U15534 ( .A(x[2906]), .B(y[2906]), .Z(n9763) );
  NANDN U15535 ( .A(n11755), .B(n9763), .Z(n9768) );
  NANDN U15536 ( .A(x[2905]), .B(y[2905]), .Z(n9764) );
  NANDN U15537 ( .A(n9768), .B(n9764), .Z(n26167) );
  ANDN U15538 ( .B(n9765), .A(n26167), .Z(n9766) );
  NANDN U15539 ( .A(n11759), .B(n9766), .Z(n9772) );
  ANDN U15540 ( .B(x[2906]), .A(y[2906]), .Z(n11754) );
  NANDN U15541 ( .A(y[2905]), .B(x[2905]), .Z(n17875) );
  NANDN U15542 ( .A(n11754), .B(n17875), .Z(n9767) );
  NANDN U15543 ( .A(n9768), .B(n9767), .Z(n9771) );
  NANDN U15544 ( .A(y[2908]), .B(x[2908]), .Z(n9770) );
  NANDN U15545 ( .A(y[2907]), .B(x[2907]), .Z(n9769) );
  NAND U15546 ( .A(n9770), .B(n9769), .Z(n11756) );
  ANDN U15547 ( .B(n9771), .A(n11756), .Z(n26168) );
  NAND U15548 ( .A(n9772), .B(n26168), .Z(n9773) );
  NANDN U15549 ( .A(x[2908]), .B(y[2908]), .Z(n26170) );
  NAND U15550 ( .A(n9773), .B(n26170), .Z(n9774) );
  NANDN U15551 ( .A(y[2909]), .B(x[2909]), .Z(n26172) );
  NANDN U15552 ( .A(x[2909]), .B(y[2909]), .Z(n9776) );
  NANDN U15553 ( .A(x[2910]), .B(y[2910]), .Z(n9775) );
  AND U15554 ( .A(n9776), .B(n9775), .Z(n26175) );
  ANDN U15555 ( .B(x[2913]), .A(y[2913]), .Z(n26184) );
  NANDN U15556 ( .A(y[2912]), .B(x[2912]), .Z(n26180) );
  NANDN U15557 ( .A(n26184), .B(n26180), .Z(n17888) );
  NANDN U15558 ( .A(x[2913]), .B(y[2913]), .Z(n17889) );
  ANDN U15559 ( .B(y[2912]), .A(x[2912]), .Z(n11753) );
  ANDN U15560 ( .B(n17889), .A(n11753), .Z(n26182) );
  ANDN U15561 ( .B(y[2915]), .A(x[2915]), .Z(n9778) );
  NANDN U15562 ( .A(x[2914]), .B(y[2914]), .Z(n9777) );
  NANDN U15563 ( .A(n9778), .B(n9777), .Z(n26189) );
  NANDN U15564 ( .A(y[2915]), .B(x[2915]), .Z(n26190) );
  NANDN U15565 ( .A(y[2914]), .B(x[2914]), .Z(n26185) );
  OR U15566 ( .A(n9778), .B(n26185), .Z(n9779) );
  NAND U15567 ( .A(n26190), .B(n9779), .Z(n17892) );
  ANDN U15568 ( .B(x[2916]), .A(y[2916]), .Z(n11751) );
  ANDN U15569 ( .B(y[2919]), .A(x[2919]), .Z(n26201) );
  IV U15570 ( .A(x[2920]), .Z(n17901) );
  NANDN U15571 ( .A(y[2921]), .B(x[2921]), .Z(n9780) );
  ANDN U15572 ( .B(x[2922]), .A(y[2922]), .Z(n11748) );
  ANDN U15573 ( .B(n9780), .A(n11748), .Z(n26206) );
  NANDN U15574 ( .A(n9781), .B(n26206), .Z(n9782) );
  AND U15575 ( .A(n26209), .B(n9782), .Z(n9783) );
  ANDN U15576 ( .B(y[2923]), .A(x[2923]), .Z(n17914) );
  ANDN U15577 ( .B(n9783), .A(n17914), .Z(n9784) );
  ANDN U15578 ( .B(n26210), .A(n9784), .Z(n9785) );
  NAND U15579 ( .A(n9786), .B(n9785), .Z(n9787) );
  NAND U15580 ( .A(n9788), .B(n9787), .Z(n9789) );
  AND U15581 ( .A(n26218), .B(n9789), .Z(n9790) );
  NANDN U15582 ( .A(n11747), .B(n9790), .Z(n9791) );
  NANDN U15583 ( .A(n26220), .B(n9791), .Z(n9792) );
  NANDN U15584 ( .A(y[2927]), .B(x[2927]), .Z(n17920) );
  ANDN U15585 ( .B(x[2928]), .A(y[2928]), .Z(n11743) );
  ANDN U15586 ( .B(n17920), .A(n11743), .Z(n26222) );
  NAND U15587 ( .A(n9792), .B(n26222), .Z(n9793) );
  NANDN U15588 ( .A(x[2928]), .B(y[2928]), .Z(n11745) );
  NANDN U15589 ( .A(x[2929]), .B(y[2929]), .Z(n17928) );
  NAND U15590 ( .A(n11745), .B(n17928), .Z(n26225) );
  ANDN U15591 ( .B(n9793), .A(n26225), .Z(n9794) );
  ANDN U15592 ( .B(x[2930]), .A(y[2930]), .Z(n17930) );
  ANDN U15593 ( .B(x[2929]), .A(y[2929]), .Z(n11742) );
  NOR U15594 ( .A(n17930), .B(n11742), .Z(n26226) );
  NANDN U15595 ( .A(n9794), .B(n26226), .Z(n9795) );
  NAND U15596 ( .A(n9796), .B(n9795), .Z(n9797) );
  AND U15597 ( .A(n26234), .B(n9797), .Z(n9798) );
  NANDN U15598 ( .A(y[2931]), .B(x[2931]), .Z(n26230) );
  NAND U15599 ( .A(n9798), .B(n26230), .Z(n9799) );
  NANDN U15600 ( .A(x[2933]), .B(y[2933]), .Z(n26236) );
  NAND U15601 ( .A(n9799), .B(n26236), .Z(n9800) );
  OR U15602 ( .A(n11741), .B(n9800), .Z(n9801) );
  NANDN U15603 ( .A(x[2936]), .B(y[2936]), .Z(n26244) );
  NANDN U15604 ( .A(x[2939]), .B(y[2939]), .Z(n9802) );
  ANDN U15605 ( .B(y[2940]), .A(x[2940]), .Z(n9803) );
  ANDN U15606 ( .B(n9802), .A(n9803), .Z(n26252) );
  ANDN U15607 ( .B(y[2938]), .A(x[2938]), .Z(n17950) );
  NANDN U15608 ( .A(y[2940]), .B(x[2940]), .Z(n26254) );
  NANDN U15609 ( .A(y[2939]), .B(x[2939]), .Z(n17952) );
  NANDN U15610 ( .A(x[2941]), .B(y[2941]), .Z(n26256) );
  NANDN U15611 ( .A(y[2942]), .B(x[2942]), .Z(n11737) );
  NANDN U15612 ( .A(y[2941]), .B(x[2941]), .Z(n17956) );
  NAND U15613 ( .A(n11737), .B(n17956), .Z(n26258) );
  NANDN U15614 ( .A(x[2942]), .B(y[2942]), .Z(n17959) );
  ANDN U15615 ( .B(y[2943]), .A(x[2943]), .Z(n11736) );
  ANDN U15616 ( .B(n17959), .A(n11736), .Z(n26260) );
  ANDN U15617 ( .B(x[2943]), .A(y[2943]), .Z(n26262) );
  ANDN U15618 ( .B(x[2944]), .A(y[2944]), .Z(n11735) );
  NAND U15619 ( .A(n9805), .B(n9804), .Z(n9806) );
  NAND U15620 ( .A(n9807), .B(n9806), .Z(n9810) );
  NANDN U15621 ( .A(x[2948]), .B(y[2948]), .Z(n9808) );
  NANDN U15622 ( .A(x[2949]), .B(y[2949]), .Z(n17974) );
  NAND U15623 ( .A(n9808), .B(n17974), .Z(n9813) );
  NANDN U15624 ( .A(x[2947]), .B(y[2947]), .Z(n9809) );
  NANDN U15625 ( .A(n9813), .B(n9809), .Z(n26273) );
  ANDN U15626 ( .B(n9810), .A(n26273), .Z(n9811) );
  NANDN U15627 ( .A(n11732), .B(n9811), .Z(n9817) );
  ANDN U15628 ( .B(x[2948]), .A(y[2948]), .Z(n17973) );
  NANDN U15629 ( .A(y[2947]), .B(x[2947]), .Z(n11731) );
  NANDN U15630 ( .A(n17973), .B(n11731), .Z(n9812) );
  NANDN U15631 ( .A(n9813), .B(n9812), .Z(n9816) );
  NANDN U15632 ( .A(y[2950]), .B(x[2950]), .Z(n9815) );
  NANDN U15633 ( .A(y[2949]), .B(x[2949]), .Z(n9814) );
  NAND U15634 ( .A(n9815), .B(n9814), .Z(n17972) );
  ANDN U15635 ( .B(n9816), .A(n17972), .Z(n26274) );
  NAND U15636 ( .A(n9817), .B(n26274), .Z(n9818) );
  AND U15637 ( .A(n26277), .B(n9818), .Z(n9819) );
  NANDN U15638 ( .A(n17980), .B(n9819), .Z(n9820) );
  NANDN U15639 ( .A(y[2951]), .B(x[2951]), .Z(n26278) );
  NAND U15640 ( .A(n9820), .B(n26278), .Z(n9821) );
  NAND U15641 ( .A(n9822), .B(n9821), .Z(n9823) );
  NAND U15642 ( .A(n11729), .B(n9823), .Z(n9824) );
  NANDN U15643 ( .A(x[2953]), .B(y[2953]), .Z(n26285) );
  NAND U15644 ( .A(n9824), .B(n26285), .Z(n9825) );
  ANDN U15645 ( .B(x[2953]), .A(y[2953]), .Z(n11730) );
  ANDN U15646 ( .B(n9825), .A(n11730), .Z(n9826) );
  NANDN U15647 ( .A(y[2954]), .B(x[2954]), .Z(n26286) );
  NAND U15648 ( .A(n9826), .B(n26286), .Z(n9827) );
  NANDN U15649 ( .A(x[2955]), .B(y[2955]), .Z(n17991) );
  NANDN U15650 ( .A(x[2954]), .B(y[2954]), .Z(n17984) );
  NAND U15651 ( .A(n17991), .B(n17984), .Z(n26288) );
  ANDN U15652 ( .B(n9827), .A(n26288), .Z(n9828) );
  ANDN U15653 ( .B(x[2956]), .A(y[2956]), .Z(n11728) );
  ANDN U15654 ( .B(x[2955]), .A(y[2955]), .Z(n17986) );
  NOR U15655 ( .A(n11728), .B(n17986), .Z(n26290) );
  NANDN U15656 ( .A(n9828), .B(n26290), .Z(n9829) );
  NANDN U15657 ( .A(n26293), .B(n9829), .Z(n9830) );
  NANDN U15658 ( .A(y[2957]), .B(x[2957]), .Z(n26294) );
  NAND U15659 ( .A(n9830), .B(n26294), .Z(n9831) );
  OR U15660 ( .A(n11727), .B(n9831), .Z(n9832) );
  NANDN U15661 ( .A(y[2960]), .B(x[2960]), .Z(n26303) );
  ANDN U15662 ( .B(x[2959]), .A(y[2959]), .Z(n11726) );
  ANDN U15663 ( .B(x[2962]), .A(y[2962]), .Z(n11721) );
  ANDN U15664 ( .B(x[2961]), .A(y[2961]), .Z(n11723) );
  NOR U15665 ( .A(n11721), .B(n11723), .Z(n26306) );
  NANDN U15666 ( .A(y[2965]), .B(x[2965]), .Z(n26314) );
  ANDN U15667 ( .B(x[2966]), .A(y[2966]), .Z(n18013) );
  ANDN U15668 ( .B(y[2966]), .A(x[2966]), .Z(n11719) );
  NANDN U15669 ( .A(y[2968]), .B(x[2968]), .Z(n26322) );
  ANDN U15670 ( .B(x[2967]), .A(y[2967]), .Z(n18014) );
  NANDN U15671 ( .A(x[2969]), .B(y[2969]), .Z(n18024) );
  ANDN U15672 ( .B(y[2968]), .A(x[2968]), .Z(n18016) );
  ANDN U15673 ( .B(n18024), .A(n18016), .Z(n26324) );
  NANDN U15674 ( .A(y[2969]), .B(x[2969]), .Z(n18020) );
  NANDN U15675 ( .A(y[2970]), .B(x[2970]), .Z(n11717) );
  NAND U15676 ( .A(n18020), .B(n11717), .Z(n26326) );
  NANDN U15677 ( .A(x[2972]), .B(y[2972]), .Z(n26332) );
  ANDN U15678 ( .B(y[2973]), .A(x[2973]), .Z(n18032) );
  ANDN U15679 ( .B(n26332), .A(n18032), .Z(n9836) );
  ANDN U15680 ( .B(x[2973]), .A(y[2973]), .Z(n11716) );
  NANDN U15681 ( .A(x[2975]), .B(y[2975]), .Z(n26341) );
  ANDN U15682 ( .B(y[2974]), .A(x[2974]), .Z(n18033) );
  ANDN U15683 ( .B(x[2976]), .A(y[2976]), .Z(n11712) );
  ANDN U15684 ( .B(x[2975]), .A(y[2975]), .Z(n11714) );
  NOR U15685 ( .A(n11712), .B(n11714), .Z(n26342) );
  NANDN U15686 ( .A(x[2976]), .B(y[2976]), .Z(n18037) );
  NANDN U15687 ( .A(x[2977]), .B(y[2977]), .Z(n11711) );
  NAND U15688 ( .A(n18037), .B(n11711), .Z(n26345) );
  NANDN U15689 ( .A(y[2979]), .B(x[2979]), .Z(n26350) );
  ANDN U15690 ( .B(x[2980]), .A(y[2980]), .Z(n18048) );
  ANDN U15691 ( .B(y[2980]), .A(x[2980]), .Z(n11710) );
  NANDN U15692 ( .A(y[2982]), .B(x[2982]), .Z(n26358) );
  ANDN U15693 ( .B(x[2981]), .A(y[2981]), .Z(n18049) );
  NANDN U15694 ( .A(x[2983]), .B(y[2983]), .Z(n18059) );
  ANDN U15695 ( .B(y[2982]), .A(x[2982]), .Z(n18051) );
  ANDN U15696 ( .B(n18059), .A(n18051), .Z(n26360) );
  NANDN U15697 ( .A(y[2983]), .B(x[2983]), .Z(n18055) );
  NANDN U15698 ( .A(y[2984]), .B(x[2984]), .Z(n11708) );
  NAND U15699 ( .A(n18055), .B(n11708), .Z(n26362) );
  NANDN U15700 ( .A(x[2986]), .B(y[2986]), .Z(n26368) );
  ANDN U15701 ( .B(y[2987]), .A(x[2987]), .Z(n18067) );
  ANDN U15702 ( .B(x[2987]), .A(y[2987]), .Z(n11707) );
  NANDN U15703 ( .A(x[2989]), .B(y[2989]), .Z(n26377) );
  ANDN U15704 ( .B(y[2988]), .A(x[2988]), .Z(n18068) );
  ANDN U15705 ( .B(x[2990]), .A(y[2990]), .Z(n11703) );
  ANDN U15706 ( .B(x[2989]), .A(y[2989]), .Z(n11705) );
  NOR U15707 ( .A(n11703), .B(n11705), .Z(n26378) );
  NANDN U15708 ( .A(x[2990]), .B(y[2990]), .Z(n18072) );
  NANDN U15709 ( .A(x[2991]), .B(y[2991]), .Z(n11702) );
  NAND U15710 ( .A(n18072), .B(n11702), .Z(n26381) );
  NANDN U15711 ( .A(y[2993]), .B(x[2993]), .Z(n26386) );
  ANDN U15712 ( .B(x[2994]), .A(y[2994]), .Z(n18083) );
  ANDN U15713 ( .B(y[2994]), .A(x[2994]), .Z(n11700) );
  NANDN U15714 ( .A(y[2996]), .B(x[2996]), .Z(n26394) );
  ANDN U15715 ( .B(x[2995]), .A(y[2995]), .Z(n18084) );
  NANDN U15716 ( .A(x[2997]), .B(y[2997]), .Z(n18094) );
  ANDN U15717 ( .B(y[2996]), .A(x[2996]), .Z(n18086) );
  ANDN U15718 ( .B(n18094), .A(n18086), .Z(n26396) );
  NANDN U15719 ( .A(y[2997]), .B(x[2997]), .Z(n18090) );
  NANDN U15720 ( .A(y[2998]), .B(x[2998]), .Z(n11699) );
  NAND U15721 ( .A(n18090), .B(n11699), .Z(n26398) );
  NANDN U15722 ( .A(x[3000]), .B(y[3000]), .Z(n26404) );
  ANDN U15723 ( .B(y[3001]), .A(x[3001]), .Z(n18102) );
  ANDN U15724 ( .B(x[3001]), .A(y[3001]), .Z(n11697) );
  NANDN U15725 ( .A(x[3003]), .B(y[3003]), .Z(n26413) );
  ANDN U15726 ( .B(y[3002]), .A(x[3002]), .Z(n18103) );
  ANDN U15727 ( .B(x[3004]), .A(y[3004]), .Z(n11694) );
  ANDN U15728 ( .B(x[3003]), .A(y[3003]), .Z(n11696) );
  NOR U15729 ( .A(n11694), .B(n11696), .Z(n26414) );
  NANDN U15730 ( .A(x[3004]), .B(y[3004]), .Z(n18107) );
  NANDN U15731 ( .A(x[3005]), .B(y[3005]), .Z(n11693) );
  NAND U15732 ( .A(n18107), .B(n11693), .Z(n26417) );
  NANDN U15733 ( .A(y[3007]), .B(x[3007]), .Z(n26422) );
  ANDN U15734 ( .B(x[3008]), .A(y[3008]), .Z(n18118) );
  ANDN U15735 ( .B(y[3008]), .A(x[3008]), .Z(n11692) );
  NANDN U15736 ( .A(y[3010]), .B(x[3010]), .Z(n26430) );
  ANDN U15737 ( .B(x[3009]), .A(y[3009]), .Z(n18119) );
  NANDN U15738 ( .A(x[3011]), .B(y[3011]), .Z(n18129) );
  ANDN U15739 ( .B(y[3010]), .A(x[3010]), .Z(n18121) );
  ANDN U15740 ( .B(n18129), .A(n18121), .Z(n26432) );
  NANDN U15741 ( .A(y[3011]), .B(x[3011]), .Z(n18125) );
  NANDN U15742 ( .A(y[3012]), .B(x[3012]), .Z(n11690) );
  NAND U15743 ( .A(n18125), .B(n11690), .Z(n26434) );
  NANDN U15744 ( .A(x[3014]), .B(y[3014]), .Z(n26440) );
  ANDN U15745 ( .B(y[3015]), .A(x[3015]), .Z(n18137) );
  ANDN U15746 ( .B(x[3015]), .A(y[3015]), .Z(n11689) );
  NANDN U15747 ( .A(x[3017]), .B(y[3017]), .Z(n26449) );
  ANDN U15748 ( .B(y[3016]), .A(x[3016]), .Z(n18138) );
  XNOR U15749 ( .A(x[3018]), .B(y[3018]), .Z(n9841) );
  ANDN U15750 ( .B(x[3017]), .A(y[3017]), .Z(n11687) );
  ANDN U15751 ( .B(n9841), .A(n11687), .Z(n26450) );
  IV U15752 ( .A(x[3018]), .Z(n11686) );
  NAND U15753 ( .A(n11686), .B(y[3018]), .Z(n9842) );
  NANDN U15754 ( .A(x[3019]), .B(y[3019]), .Z(n11685) );
  NAND U15755 ( .A(n9842), .B(n11685), .Z(n26453) );
  NANDN U15756 ( .A(y[3019]), .B(x[3019]), .Z(n18145) );
  ANDN U15757 ( .B(x[3020]), .A(y[3020]), .Z(n11684) );
  ANDN U15758 ( .B(n18145), .A(n11684), .Z(n26454) );
  NANDN U15759 ( .A(y[3021]), .B(x[3021]), .Z(n26458) );
  ANDN U15760 ( .B(x[3022]), .A(y[3022]), .Z(n18155) );
  ANDN U15761 ( .B(y[3022]), .A(x[3022]), .Z(n11683) );
  NANDN U15762 ( .A(y[3023]), .B(x[3023]), .Z(n18154) );
  NANDN U15763 ( .A(y[3024]), .B(x[3024]), .Z(n26466) );
  ANDN U15764 ( .B(y[3025]), .A(x[3025]), .Z(n11679) );
  ANDN U15765 ( .B(y[3024]), .A(x[3024]), .Z(n11681) );
  NOR U15766 ( .A(n11679), .B(n11681), .Z(n26468) );
  NANDN U15767 ( .A(y[3026]), .B(x[3026]), .Z(n18164) );
  NANDN U15768 ( .A(y[3025]), .B(x[3025]), .Z(n11680) );
  NAND U15769 ( .A(n18164), .B(n11680), .Z(n26470) );
  ANDN U15770 ( .B(y[3027]), .A(x[3027]), .Z(n18166) );
  ANDN U15771 ( .B(y[3026]), .A(x[3026]), .Z(n11678) );
  NOR U15772 ( .A(n18166), .B(n11678), .Z(n26472) );
  NANDN U15773 ( .A(x[3028]), .B(y[3028]), .Z(n26476) );
  ANDN U15774 ( .B(y[3029]), .A(x[3029]), .Z(n18172) );
  ANDN U15775 ( .B(x[3029]), .A(y[3029]), .Z(n18170) );
  NANDN U15776 ( .A(x[3031]), .B(y[3031]), .Z(n26485) );
  ANDN U15777 ( .B(y[3030]), .A(x[3030]), .Z(n18173) );
  ANDN U15778 ( .B(x[3031]), .A(y[3031]), .Z(n18175) );
  XOR U15779 ( .A(x[3032]), .B(y[3032]), .Z(n18180) );
  NOR U15780 ( .A(n18175), .B(n18180), .Z(n26486) );
  NANDN U15781 ( .A(x[3032]), .B(y[3032]), .Z(n9845) );
  NANDN U15782 ( .A(x[3033]), .B(y[3033]), .Z(n11675) );
  NAND U15783 ( .A(n9845), .B(n11675), .Z(n26489) );
  NANDN U15784 ( .A(y[3035]), .B(x[3035]), .Z(n26494) );
  ANDN U15785 ( .B(x[3036]), .A(y[3036]), .Z(n18189) );
  ANDN U15786 ( .B(y[3036]), .A(x[3036]), .Z(n11674) );
  ANDN U15787 ( .B(x[3037]), .A(y[3037]), .Z(n18190) );
  ANDN U15788 ( .B(x[3038]), .A(y[3038]), .Z(n26503) );
  IV U15789 ( .A(y[3039]), .Z(n18196) );
  NAND U15790 ( .A(n18196), .B(x[3039]), .Z(n9848) );
  NANDN U15791 ( .A(y[3040]), .B(x[3040]), .Z(n9847) );
  NAND U15792 ( .A(n9848), .B(n9847), .Z(n26506) );
  NANDN U15793 ( .A(x[3042]), .B(y[3042]), .Z(n26512) );
  ANDN U15794 ( .B(y[3043]), .A(x[3043]), .Z(n18212) );
  ANDN U15795 ( .B(x[3043]), .A(y[3043]), .Z(n18210) );
  NANDN U15796 ( .A(x[3045]), .B(y[3045]), .Z(n26521) );
  ANDN U15797 ( .B(y[3044]), .A(x[3044]), .Z(n18213) );
  ANDN U15798 ( .B(x[3045]), .A(y[3045]), .Z(n18215) );
  XOR U15799 ( .A(x[3046]), .B(y[3046]), .Z(n18220) );
  NOR U15800 ( .A(n18215), .B(n18220), .Z(n26522) );
  NANDN U15801 ( .A(x[3046]), .B(y[3046]), .Z(n9851) );
  NANDN U15802 ( .A(x[3047]), .B(y[3047]), .Z(n11669) );
  NAND U15803 ( .A(n9851), .B(n11669), .Z(n26525) );
  NANDN U15804 ( .A(y[3049]), .B(x[3049]), .Z(n26530) );
  ANDN U15805 ( .B(x[3050]), .A(y[3050]), .Z(n18229) );
  ANDN U15806 ( .B(y[3050]), .A(x[3050]), .Z(n11668) );
  NANDN U15807 ( .A(y[3052]), .B(x[3052]), .Z(n26538) );
  ANDN U15808 ( .B(x[3051]), .A(y[3051]), .Z(n18230) );
  ANDN U15809 ( .B(y[3053]), .A(x[3053]), .Z(n11666) );
  ANDN U15810 ( .B(y[3052]), .A(x[3052]), .Z(n18232) );
  NOR U15811 ( .A(n11666), .B(n18232), .Z(n26540) );
  ANDN U15812 ( .B(x[3054]), .A(y[3054]), .Z(n26545) );
  ANDN U15813 ( .B(y[3055]), .A(x[3055]), .Z(n18241) );
  ANDN U15814 ( .B(y[3054]), .A(x[3054]), .Z(n11665) );
  NOR U15815 ( .A(n18241), .B(n11665), .Z(n26546) );
  ANDN U15816 ( .B(x[3056]), .A(y[3056]), .Z(n18245) );
  NAND U15817 ( .A(n9853), .B(n9852), .Z(n9854) );
  NAND U15818 ( .A(n9855), .B(n9854), .Z(n9856) );
  AND U15819 ( .A(n26558), .B(n9856), .Z(n9857) );
  NANDN U15820 ( .A(n11664), .B(n9857), .Z(n9858) );
  ANDN U15821 ( .B(x[3059]), .A(y[3059]), .Z(n18248) );
  XOR U15822 ( .A(x[3060]), .B(y[3060]), .Z(n18251) );
  NOR U15823 ( .A(n18248), .B(n18251), .Z(n26561) );
  NAND U15824 ( .A(n9858), .B(n26561), .Z(n9859) );
  AND U15825 ( .A(n26562), .B(n9859), .Z(n9860) );
  OR U15826 ( .A(n26565), .B(n9860), .Z(n9861) );
  AND U15827 ( .A(n26566), .B(n9861), .Z(n9862) );
  ANDN U15828 ( .B(y[3063]), .A(x[3063]), .Z(n11661) );
  ANDN U15829 ( .B(n9862), .A(n11661), .Z(n9863) );
  ANDN U15830 ( .B(n26568), .A(n9863), .Z(n9864) );
  NAND U15831 ( .A(n9865), .B(n9864), .Z(n9866) );
  NAND U15832 ( .A(n9867), .B(n9866), .Z(n9868) );
  AND U15833 ( .A(n26576), .B(n9868), .Z(n9869) );
  ANDN U15834 ( .B(x[3065]), .A(y[3065]), .Z(n11659) );
  ANDN U15835 ( .B(n9869), .A(n11659), .Z(n9870) );
  ANDN U15836 ( .B(y[3067]), .A(x[3067]), .Z(n11656) );
  ANDN U15837 ( .B(y[3066]), .A(x[3066]), .Z(n11657) );
  NOR U15838 ( .A(n11656), .B(n11657), .Z(n26578) );
  NANDN U15839 ( .A(n9870), .B(n26578), .Z(n9871) );
  AND U15840 ( .A(n26580), .B(n9871), .Z(n9872) );
  NANDN U15841 ( .A(n11654), .B(n9872), .Z(n9873) );
  ANDN U15842 ( .B(y[3069]), .A(x[3069]), .Z(n11652) );
  ANDN U15843 ( .B(y[3074]), .A(x[3074]), .Z(n11648) );
  NANDN U15844 ( .A(x[3076]), .B(y[3076]), .Z(n11643) );
  IV U15845 ( .A(x[3078]), .Z(n18285) );
  ANDN U15846 ( .B(y[3079]), .A(x[3079]), .Z(n18294) );
  IV U15847 ( .A(x[3080]), .Z(n18292) );
  NANDN U15848 ( .A(n9875), .B(y[3082]), .Z(n9878) );
  XNOR U15849 ( .A(n9875), .B(y[3082]), .Z(n9876) );
  NANDN U15850 ( .A(x[3082]), .B(n9876), .Z(n9877) );
  NAND U15851 ( .A(n9878), .B(n9877), .Z(n9879) );
  NAND U15852 ( .A(n9880), .B(n9879), .Z(n9881) );
  NAND U15853 ( .A(n11637), .B(n9881), .Z(n9882) );
  NAND U15854 ( .A(n9883), .B(n9882), .Z(n9884) );
  NAND U15855 ( .A(n9885), .B(n9884), .Z(n9886) );
  NANDN U15856 ( .A(y[3085]), .B(x[3085]), .Z(n18303) );
  NAND U15857 ( .A(n9886), .B(n18303), .Z(n9887) );
  NANDN U15858 ( .A(n9887), .B(y[3086]), .Z(n9890) );
  XNOR U15859 ( .A(n9887), .B(y[3086]), .Z(n9888) );
  NANDN U15860 ( .A(x[3086]), .B(n9888), .Z(n9889) );
  NAND U15861 ( .A(n9890), .B(n9889), .Z(n9891) );
  NAND U15862 ( .A(n9892), .B(n9891), .Z(n9893) );
  AND U15863 ( .A(n11633), .B(n9893), .Z(n9895) );
  XNOR U15864 ( .A(y[3088]), .B(n9895), .Z(n9894) );
  NANDN U15865 ( .A(x[3088]), .B(n9894), .Z(n9897) );
  NANDN U15866 ( .A(n9895), .B(y[3088]), .Z(n9896) );
  AND U15867 ( .A(n9897), .B(n9896), .Z(n9898) );
  NAND U15868 ( .A(n9899), .B(n9898), .Z(n9900) );
  NAND U15869 ( .A(n9901), .B(n9900), .Z(n9902) );
  AND U15870 ( .A(n26634), .B(n9902), .Z(n9903) );
  ANDN U15871 ( .B(y[3090]), .A(x[3090]), .Z(n18312) );
  ANDN U15872 ( .B(n9903), .A(n18312), .Z(n9904) );
  ANDN U15873 ( .B(x[3091]), .A(y[3091]), .Z(n18314) );
  NOR U15874 ( .A(n9904), .B(n18314), .Z(n9906) );
  XNOR U15875 ( .A(x[3092]), .B(y[3092]), .Z(n9905) );
  NAND U15876 ( .A(n9906), .B(n9905), .Z(n9907) );
  IV U15877 ( .A(y[3092]), .Z(n11630) );
  NOR U15878 ( .A(n11630), .B(x[3092]), .Z(n26632) );
  ANDN U15879 ( .B(n9907), .A(n26632), .Z(n9908) );
  NANDN U15880 ( .A(x[3093]), .B(y[3093]), .Z(n26640) );
  NAND U15881 ( .A(n9908), .B(n26640), .Z(n9909) );
  NANDN U15882 ( .A(n9910), .B(n9909), .Z(n9911) );
  OR U15883 ( .A(n11628), .B(n9911), .Z(n9912) );
  NAND U15884 ( .A(n9913), .B(n9912), .Z(n9914) );
  ANDN U15885 ( .B(x[3095]), .A(y[3095]), .Z(n11627) );
  ANDN U15886 ( .B(n9914), .A(n11627), .Z(n9915) );
  NAND U15887 ( .A(n9916), .B(n9915), .Z(n9917) );
  AND U15888 ( .A(n9918), .B(n9917), .Z(n9920) );
  ANDN U15889 ( .B(x[3097]), .A(y[3097]), .Z(n18326) );
  ANDN U15890 ( .B(x[3098]), .A(y[3098]), .Z(n11620) );
  ANDN U15891 ( .B(y[3098]), .A(x[3098]), .Z(n11623) );
  ANDN U15892 ( .B(y[3100]), .A(x[3100]), .Z(n11619) );
  ANDN U15893 ( .B(y[3102]), .A(x[3102]), .Z(n18333) );
  ANDN U15894 ( .B(y[3103]), .A(x[3103]), .Z(n11612) );
  NANDN U15895 ( .A(x[3106]), .B(y[3106]), .Z(n11609) );
  ANDN U15896 ( .B(y[3107]), .A(x[3107]), .Z(n11605) );
  ANDN U15897 ( .B(y[3110]), .A(x[3110]), .Z(n18343) );
  ANDN U15898 ( .B(y[3111]), .A(x[3111]), .Z(n11599) );
  ANDN U15899 ( .B(y[3114]), .A(x[3114]), .Z(n11594) );
  IV U15900 ( .A(n11594), .Z(n9925) );
  ANDN U15901 ( .B(y[3115]), .A(x[3115]), .Z(n11591) );
  ANDN U15902 ( .B(y[3118]), .A(x[3118]), .Z(n18353) );
  ANDN U15903 ( .B(y[3119]), .A(x[3119]), .Z(n11585) );
  AND U15904 ( .A(n9927), .B(n9926), .Z(n9929) );
  ANDN U15905 ( .B(y[3122]), .A(x[3122]), .Z(n18359) );
  ANDN U15906 ( .B(y[3123]), .A(x[3123]), .Z(n11578) );
  NANDN U15907 ( .A(n9929), .B(n9928), .Z(n9930) );
  NANDN U15908 ( .A(n11581), .B(n9930), .Z(n9931) );
  NAND U15909 ( .A(n9932), .B(n9931), .Z(n9933) );
  NAND U15910 ( .A(n11576), .B(n9933), .Z(n9934) );
  NAND U15911 ( .A(n9935), .B(n9934), .Z(n9936) );
  AND U15912 ( .A(n9937), .B(n9936), .Z(n9939) );
  NANDN U15913 ( .A(x[3126]), .B(y[3126]), .Z(n11575) );
  ANDN U15914 ( .B(y[3127]), .A(x[3127]), .Z(n11571) );
  ANDN U15915 ( .B(n11575), .A(n11571), .Z(n9938) );
  NANDN U15916 ( .A(n9939), .B(n9938), .Z(n9940) );
  NANDN U15917 ( .A(n11573), .B(n9940), .Z(n9941) );
  NAND U15918 ( .A(n9942), .B(n9941), .Z(n9943) );
  NAND U15919 ( .A(n11569), .B(n9943), .Z(n9944) );
  OR U15920 ( .A(n11568), .B(n9944), .Z(n9945) );
  NANDN U15921 ( .A(n26713), .B(n9945), .Z(n9948) );
  NANDN U15922 ( .A(y[3130]), .B(x[3130]), .Z(n9947) );
  NANDN U15923 ( .A(y[3131]), .B(x[3131]), .Z(n9946) );
  AND U15924 ( .A(n9947), .B(n9946), .Z(n26714) );
  NAND U15925 ( .A(n9948), .B(n26714), .Z(n9949) );
  NANDN U15926 ( .A(n26716), .B(n9949), .Z(n9952) );
  NANDN U15927 ( .A(y[3132]), .B(x[3132]), .Z(n9951) );
  NANDN U15928 ( .A(y[3133]), .B(x[3133]), .Z(n9950) );
  AND U15929 ( .A(n9951), .B(n9950), .Z(n26718) );
  NANDN U15930 ( .A(x[3134]), .B(y[3134]), .Z(n9954) );
  NANDN U15931 ( .A(x[3133]), .B(y[3133]), .Z(n9953) );
  NAND U15932 ( .A(n9954), .B(n9953), .Z(n26720) );
  NANDN U15933 ( .A(y[3134]), .B(x[3134]), .Z(n9956) );
  NANDN U15934 ( .A(y[3135]), .B(x[3135]), .Z(n9955) );
  AND U15935 ( .A(n9956), .B(n9955), .Z(n26722) );
  NANDN U15936 ( .A(x[3136]), .B(y[3136]), .Z(n9958) );
  NANDN U15937 ( .A(x[3135]), .B(y[3135]), .Z(n9957) );
  NAND U15938 ( .A(n9958), .B(n9957), .Z(n26724) );
  IV U15939 ( .A(y[3141]), .Z(n11561) );
  NAND U15940 ( .A(n9960), .B(n9959), .Z(n9961) );
  AND U15941 ( .A(n11557), .B(n9961), .Z(n9962) );
  NANDN U15942 ( .A(n9962), .B(x[3143]), .Z(n9965) );
  XNOR U15943 ( .A(n9962), .B(x[3143]), .Z(n9963) );
  NANDN U15944 ( .A(y[3143]), .B(n9963), .Z(n9964) );
  NAND U15945 ( .A(n9965), .B(n9964), .Z(n9966) );
  NAND U15946 ( .A(n9967), .B(n9966), .Z(n9968) );
  NAND U15947 ( .A(n11556), .B(n9968), .Z(n9969) );
  NAND U15948 ( .A(n9970), .B(n9969), .Z(n9971) );
  NAND U15949 ( .A(n11555), .B(n9971), .Z(n9972) );
  ANDN U15950 ( .B(y[3146]), .A(x[3146]), .Z(n18391) );
  ANDN U15951 ( .B(n9972), .A(n18391), .Z(n9975) );
  NANDN U15952 ( .A(y[3146]), .B(x[3146]), .Z(n9974) );
  NANDN U15953 ( .A(y[3147]), .B(x[3147]), .Z(n9973) );
  AND U15954 ( .A(n9974), .B(n9973), .Z(n26746) );
  NANDN U15955 ( .A(n9975), .B(n26746), .Z(n9976) );
  NANDN U15956 ( .A(n26749), .B(n9976), .Z(n9979) );
  NANDN U15957 ( .A(y[3148]), .B(x[3148]), .Z(n9978) );
  NANDN U15958 ( .A(y[3149]), .B(x[3149]), .Z(n9977) );
  AND U15959 ( .A(n9978), .B(n9977), .Z(n26750) );
  NAND U15960 ( .A(n9979), .B(n26750), .Z(n9980) );
  NANDN U15961 ( .A(n18398), .B(n9980), .Z(n9981) );
  NANDN U15962 ( .A(n18401), .B(n9981), .Z(n9982) );
  AND U15963 ( .A(n20233), .B(n9982), .Z(n9983) );
  ANDN U15964 ( .B(y[3150]), .A(x[3150]), .Z(n18397) );
  ANDN U15965 ( .B(n9983), .A(n18397), .Z(n9984) );
  XNOR U15966 ( .A(y[3152]), .B(x[3152]), .Z(n18404) );
  ANDN U15967 ( .B(y[3152]), .A(x[3152]), .Z(n20232) );
  ANDN U15968 ( .B(x[3157]), .A(y[3157]), .Z(n11550) );
  ANDN U15969 ( .B(x[3159]), .A(y[3159]), .Z(n18416) );
  IV U15970 ( .A(n18416), .Z(n9987) );
  ANDN U15971 ( .B(x[3160]), .A(y[3160]), .Z(n11546) );
  ANDN U15972 ( .B(x[3163]), .A(y[3163]), .Z(n11541) );
  ANDN U15973 ( .B(x[3164]), .A(y[3164]), .Z(n18426) );
  ANDN U15974 ( .B(x[3167]), .A(y[3167]), .Z(n18430) );
  IV U15975 ( .A(n18430), .Z(n9989) );
  ANDN U15976 ( .B(x[3168]), .A(y[3168]), .Z(n11534) );
  ANDN U15977 ( .B(x[3171]), .A(y[3171]), .Z(n18438) );
  ANDN U15978 ( .B(x[3172]), .A(y[3172]), .Z(n11530) );
  ANDN U15979 ( .B(y[3172]), .A(x[3172]), .Z(n11531) );
  NANDN U15980 ( .A(x[3173]), .B(y[3173]), .Z(n26801) );
  ANDN U15981 ( .B(x[3173]), .A(y[3173]), .Z(n11529) );
  XNOR U15982 ( .A(x[3174]), .B(y[3174]), .Z(n18443) );
  ANDN U15983 ( .B(y[3174]), .A(x[3174]), .Z(n26800) );
  NANDN U15984 ( .A(x[3176]), .B(y[3176]), .Z(n18448) );
  ANDN U15985 ( .B(y[3177]), .A(x[3177]), .Z(n18451) );
  ANDN U15986 ( .B(y[3180]), .A(x[3180]), .Z(n18455) );
  ANDN U15987 ( .B(y[3181]), .A(x[3181]), .Z(n11520) );
  ANDN U15988 ( .B(y[3184]), .A(x[3184]), .Z(n18463) );
  IV U15989 ( .A(n18463), .Z(n9994) );
  ANDN U15990 ( .B(y[3185]), .A(x[3185]), .Z(n11515) );
  ANDN U15991 ( .B(y[3188]), .A(x[3188]), .Z(n18469) );
  ANDN U15992 ( .B(y[3189]), .A(x[3189]), .Z(n11510) );
  ANDN U15993 ( .B(y[3192]), .A(x[3192]), .Z(n18475) );
  IV U15994 ( .A(n18475), .Z(n9997) );
  ANDN U15995 ( .B(y[3193]), .A(x[3193]), .Z(n11506) );
  ANDN U15996 ( .B(y[3196]), .A(x[3196]), .Z(n11501) );
  ANDN U15997 ( .B(y[3197]), .A(x[3197]), .Z(n18485) );
  ANDN U15998 ( .B(y[3200]), .A(x[3200]), .Z(n18489) );
  IV U15999 ( .A(n18489), .Z(n10000) );
  ANDN U16000 ( .B(y[3201]), .A(x[3201]), .Z(n11494) );
  ANDN U16001 ( .B(y[3204]), .A(x[3204]), .Z(n18497) );
  ANDN U16002 ( .B(y[3205]), .A(x[3205]), .Z(n11489) );
  ANDN U16003 ( .B(y[3208]), .A(x[3208]), .Z(n18503) );
  IV U16004 ( .A(n18503), .Z(n10003) );
  ANDN U16005 ( .B(y[3209]), .A(x[3209]), .Z(n11484) );
  ANDN U16006 ( .B(y[3212]), .A(x[3212]), .Z(n18509) );
  ANDN U16007 ( .B(y[3213]), .A(x[3213]), .Z(n11480) );
  ANDN U16008 ( .B(y[3216]), .A(x[3216]), .Z(n11475) );
  IV U16009 ( .A(n11475), .Z(n10006) );
  ANDN U16010 ( .B(y[3217]), .A(x[3217]), .Z(n18519) );
  ANDN U16011 ( .B(y[3220]), .A(x[3220]), .Z(n18523) );
  ANDN U16012 ( .B(y[3221]), .A(x[3221]), .Z(n11468) );
  ANDN U16013 ( .B(y[3224]), .A(x[3224]), .Z(n18531) );
  IV U16014 ( .A(n18531), .Z(n10009) );
  ANDN U16015 ( .B(y[3225]), .A(x[3225]), .Z(n11463) );
  ANDN U16016 ( .B(y[3228]), .A(x[3228]), .Z(n18537) );
  ANDN U16017 ( .B(y[3229]), .A(x[3229]), .Z(n11458) );
  ANDN U16018 ( .B(y[3232]), .A(x[3232]), .Z(n18543) );
  IV U16019 ( .A(n18543), .Z(n10012) );
  ANDN U16020 ( .B(y[3233]), .A(x[3233]), .Z(n11454) );
  ANDN U16021 ( .B(y[3236]), .A(x[3236]), .Z(n11449) );
  ANDN U16022 ( .B(y[3237]), .A(x[3237]), .Z(n18553) );
  ANDN U16023 ( .B(y[3240]), .A(x[3240]), .Z(n18557) );
  ANDN U16024 ( .B(y[3241]), .A(x[3241]), .Z(n11442) );
  ANDN U16025 ( .B(y[3244]), .A(x[3244]), .Z(n18565) );
  ANDN U16026 ( .B(y[3245]), .A(x[3245]), .Z(n11437) );
  ANDN U16027 ( .B(y[3248]), .A(x[3248]), .Z(n18571) );
  ANDN U16028 ( .B(y[3249]), .A(x[3249]), .Z(n11432) );
  ANDN U16029 ( .B(y[3252]), .A(x[3252]), .Z(n18577) );
  ANDN U16030 ( .B(y[3253]), .A(x[3253]), .Z(n11428) );
  ANDN U16031 ( .B(y[3256]), .A(x[3256]), .Z(n11423) );
  ANDN U16032 ( .B(y[3257]), .A(x[3257]), .Z(n18587) );
  IV U16033 ( .A(x[3259]), .Z(n11416) );
  ANDN U16034 ( .B(y[3260]), .A(x[3260]), .Z(n11417) );
  NANDN U16035 ( .A(x[3261]), .B(y[3261]), .Z(n10019) );
  NANDN U16036 ( .A(x[3262]), .B(y[3262]), .Z(n10018) );
  AND U16037 ( .A(n10019), .B(n10018), .Z(n26978) );
  ANDN U16038 ( .B(x[3262]), .A(y[3262]), .Z(n11415) );
  NANDN U16039 ( .A(x[3265]), .B(y[3265]), .Z(n10022) );
  NANDN U16040 ( .A(x[3266]), .B(y[3266]), .Z(n10021) );
  AND U16041 ( .A(n10022), .B(n10021), .Z(n26987) );
  NANDN U16042 ( .A(y[3267]), .B(x[3267]), .Z(n10024) );
  NANDN U16043 ( .A(y[3266]), .B(x[3266]), .Z(n10023) );
  AND U16044 ( .A(n10024), .B(n10023), .Z(n26988) );
  NANDN U16045 ( .A(x[3267]), .B(y[3267]), .Z(n10026) );
  NANDN U16046 ( .A(x[3268]), .B(y[3268]), .Z(n10025) );
  AND U16047 ( .A(n10026), .B(n10025), .Z(n26991) );
  ANDN U16048 ( .B(x[3268]), .A(y[3268]), .Z(n18603) );
  NANDN U16049 ( .A(x[3269]), .B(y[3269]), .Z(n20231) );
  ANDN U16050 ( .B(y[3270]), .A(x[3270]), .Z(n20230) );
  XNOR U16051 ( .A(x[3273]), .B(n10028), .Z(n10027) );
  IV U16052 ( .A(x[3276]), .Z(n11407) );
  IV U16053 ( .A(x[3280]), .Z(n11402) );
  IV U16054 ( .A(x[3286]), .Z(n11393) );
  IV U16055 ( .A(x[3300]), .Z(n11372) );
  IV U16056 ( .A(x[3306]), .Z(n11361) );
  IV U16057 ( .A(x[3310]), .Z(n11356) );
  NAND U16058 ( .A(n10036), .B(n10035), .Z(n10037) );
  NANDN U16059 ( .A(n10037), .B(y[3316]), .Z(n10040) );
  IV U16060 ( .A(x[3316]), .Z(n11347) );
  XNOR U16061 ( .A(n10037), .B(y[3316]), .Z(n10038) );
  NAND U16062 ( .A(n11347), .B(n10038), .Z(n10039) );
  NAND U16063 ( .A(n10040), .B(n10039), .Z(n10041) );
  NAND U16064 ( .A(n10042), .B(n10041), .Z(n10043) );
  AND U16065 ( .A(n18688), .B(n10043), .Z(n10045) );
  XNOR U16066 ( .A(y[3318]), .B(n10045), .Z(n10044) );
  NANDN U16067 ( .A(x[3318]), .B(n10044), .Z(n10047) );
  NANDN U16068 ( .A(n10045), .B(y[3318]), .Z(n10046) );
  AND U16069 ( .A(n10047), .B(n10046), .Z(n10048) );
  NANDN U16070 ( .A(x[3319]), .B(y[3319]), .Z(n20229) );
  NAND U16071 ( .A(n10048), .B(n20229), .Z(n10049) );
  NAND U16072 ( .A(n11342), .B(n10049), .Z(n10050) );
  OR U16073 ( .A(n11344), .B(n10050), .Z(n10051) );
  NAND U16074 ( .A(n10052), .B(n10051), .Z(n10053) );
  ANDN U16075 ( .B(x[3321]), .A(y[3321]), .Z(n11341) );
  ANDN U16076 ( .B(n10053), .A(n11341), .Z(n10054) );
  NAND U16077 ( .A(n10055), .B(n10054), .Z(n10056) );
  ANDN U16078 ( .B(x[3323]), .A(y[3323]), .Z(n18697) );
  IV U16079 ( .A(n18697), .Z(n10057) );
  ANDN U16080 ( .B(x[3324]), .A(y[3324]), .Z(n11339) );
  ANDN U16081 ( .B(y[3324]), .A(x[3324]), .Z(n18700) );
  NANDN U16082 ( .A(x[3325]), .B(y[3325]), .Z(n27107) );
  ANDN U16083 ( .B(x[3325]), .A(y[3325]), .Z(n11338) );
  XNOR U16084 ( .A(x[3326]), .B(y[3326]), .Z(n11337) );
  ANDN U16085 ( .B(y[3326]), .A(x[3326]), .Z(n27106) );
  ANDN U16086 ( .B(y[3328]), .A(x[3328]), .Z(n18707) );
  ANDN U16087 ( .B(y[3329]), .A(x[3329]), .Z(n11334) );
  NANDN U16088 ( .A(x[3334]), .B(y[3334]), .Z(n10061) );
  NANDN U16089 ( .A(x[3333]), .B(y[3333]), .Z(n10060) );
  AND U16090 ( .A(n10061), .B(n10060), .Z(n27124) );
  NANDN U16091 ( .A(x[3332]), .B(y[3332]), .Z(n11329) );
  NANDN U16092 ( .A(n11329), .B(n10062), .Z(n10063) );
  NANDN U16093 ( .A(x[3335]), .B(y[3335]), .Z(n10065) );
  NANDN U16094 ( .A(x[3336]), .B(y[3336]), .Z(n10064) );
  AND U16095 ( .A(n10065), .B(n10064), .Z(n27128) );
  ANDN U16096 ( .B(x[3336]), .A(y[3336]), .Z(n11328) );
  NANDN U16097 ( .A(x[3339]), .B(y[3339]), .Z(n27138) );
  XNOR U16098 ( .A(x[3340]), .B(y[3340]), .Z(n18724) );
  ANDN U16099 ( .B(x[3341]), .A(y[3341]), .Z(n11321) );
  ANDN U16100 ( .B(x[3343]), .A(y[3343]), .Z(n18730) );
  IV U16101 ( .A(n18730), .Z(n10068) );
  ANDN U16102 ( .B(x[3344]), .A(y[3344]), .Z(n11318) );
  ANDN U16103 ( .B(x[3347]), .A(y[3347]), .Z(n18736) );
  ANDN U16104 ( .B(x[3348]), .A(y[3348]), .Z(n11314) );
  ANDN U16105 ( .B(x[3351]), .A(y[3351]), .Z(n11309) );
  ANDN U16106 ( .B(x[3352]), .A(y[3352]), .Z(n18746) );
  ANDN U16107 ( .B(x[3355]), .A(y[3355]), .Z(n18750) );
  XNOR U16108 ( .A(x[3356]), .B(y[3356]), .Z(n18754) );
  ANDN U16109 ( .B(y[3358]), .A(x[3358]), .Z(n27176) );
  IV U16110 ( .A(x[3359]), .Z(n18763) );
  ANDN U16111 ( .B(x[3360]), .A(y[3360]), .Z(n18767) );
  ANDN U16112 ( .B(y[3360]), .A(x[3360]), .Z(n18764) );
  ANDN U16113 ( .B(y[3361]), .A(x[3361]), .Z(n11302) );
  ANDN U16114 ( .B(x[3361]), .A(y[3361]), .Z(n18768) );
  ANDN U16115 ( .B(x[3363]), .A(y[3363]), .Z(n11300) );
  NANDN U16116 ( .A(x[3365]), .B(y[3365]), .Z(n27195) );
  ANDN U16117 ( .B(x[3365]), .A(y[3365]), .Z(n18773) );
  ANDN U16118 ( .B(y[3366]), .A(x[3366]), .Z(n27194) );
  ANDN U16119 ( .B(y[3368]), .A(x[3368]), .Z(n11294) );
  ANDN U16120 ( .B(y[3370]), .A(x[3370]), .Z(n18784) );
  ANDN U16121 ( .B(y[3371]), .A(x[3371]), .Z(n11289) );
  AND U16122 ( .A(n10073), .B(n10072), .Z(n10076) );
  ANDN U16123 ( .B(y[3374]), .A(x[3374]), .Z(n18790) );
  IV U16124 ( .A(n18790), .Z(n10074) );
  ANDN U16125 ( .B(y[3375]), .A(x[3375]), .Z(n11284) );
  ANDN U16126 ( .B(n10074), .A(n11284), .Z(n10075) );
  NANDN U16127 ( .A(n10076), .B(n10075), .Z(n10077) );
  NANDN U16128 ( .A(n11286), .B(n10077), .Z(n10078) );
  NAND U16129 ( .A(n10079), .B(n10078), .Z(n10080) );
  NAND U16130 ( .A(n11281), .B(n10080), .Z(n10082) );
  IV U16131 ( .A(x[3377]), .Z(n11278) );
  NANDN U16132 ( .A(n10082), .B(n11278), .Z(n10081) );
  ANDN U16133 ( .B(y[3378]), .A(x[3378]), .Z(n11280) );
  ANDN U16134 ( .B(n10081), .A(n11280), .Z(n10085) );
  XOR U16135 ( .A(x[3377]), .B(n10082), .Z(n10083) );
  NAND U16136 ( .A(n10083), .B(y[3377]), .Z(n10084) );
  NAND U16137 ( .A(n10085), .B(n10084), .Z(n10088) );
  NANDN U16138 ( .A(y[3379]), .B(x[3379]), .Z(n10087) );
  NANDN U16139 ( .A(y[3378]), .B(x[3378]), .Z(n10086) );
  AND U16140 ( .A(n10087), .B(n10086), .Z(n27222) );
  NAND U16141 ( .A(n10088), .B(n27222), .Z(n10091) );
  NANDN U16142 ( .A(x[3379]), .B(y[3379]), .Z(n10090) );
  NANDN U16143 ( .A(x[3380]), .B(y[3380]), .Z(n10089) );
  AND U16144 ( .A(n10090), .B(n10089), .Z(n27225) );
  NAND U16145 ( .A(n10091), .B(n27225), .Z(n10092) );
  ANDN U16146 ( .B(x[3380]), .A(y[3380]), .Z(n18799) );
  ANDN U16147 ( .B(n10092), .A(n18799), .Z(n10093) );
  NAND U16148 ( .A(n10094), .B(n10093), .Z(n10095) );
  NAND U16149 ( .A(n10096), .B(n10095), .Z(n10097) );
  IV U16150 ( .A(x[3384]), .Z(n11273) );
  ANDN U16151 ( .B(y[3385]), .A(x[3385]), .Z(n11272) );
  ANDN U16152 ( .B(x[3385]), .A(y[3385]), .Z(n18805) );
  ANDN U16153 ( .B(x[3387]), .A(y[3387]), .Z(n18809) );
  ANDN U16154 ( .B(x[3388]), .A(y[3388]), .Z(n18814) );
  ANDN U16155 ( .B(y[3388]), .A(x[3388]), .Z(n11269) );
  NANDN U16156 ( .A(x[3389]), .B(y[3389]), .Z(n27245) );
  ANDN U16157 ( .B(x[3389]), .A(y[3389]), .Z(n18813) );
  ANDN U16158 ( .B(y[3390]), .A(x[3390]), .Z(n27244) );
  ANDN U16159 ( .B(y[3392]), .A(x[3392]), .Z(n18820) );
  ANDN U16160 ( .B(y[3393]), .A(x[3393]), .Z(n11266) );
  ANDN U16161 ( .B(y[3396]), .A(x[3396]), .Z(n11261) );
  ANDN U16162 ( .B(y[3397]), .A(x[3397]), .Z(n18830) );
  ANDN U16163 ( .B(y[3400]), .A(x[3400]), .Z(n18834) );
  ANDN U16164 ( .B(y[3401]), .A(x[3401]), .Z(n11254) );
  ANDN U16165 ( .B(y[3404]), .A(x[3404]), .Z(n18842) );
  ANDN U16166 ( .B(y[3405]), .A(x[3405]), .Z(n11249) );
  NANDN U16167 ( .A(x[3409]), .B(y[3409]), .Z(n27288) );
  ANDN U16168 ( .B(y[3408]), .A(x[3408]), .Z(n18848) );
  XNOR U16169 ( .A(x[3413]), .B(n10103), .Z(n10102) );
  NANDN U16170 ( .A(y[3413]), .B(n10102), .Z(n10105) );
  NANDN U16171 ( .A(n10103), .B(x[3413]), .Z(n10104) );
  IV U16172 ( .A(x[3416]), .Z(n11236) );
  IV U16173 ( .A(x[3420]), .Z(n11231) );
  NANDN U16174 ( .A(n10107), .B(y[3426]), .Z(n10110) );
  IV U16175 ( .A(x[3426]), .Z(n11222) );
  XNOR U16176 ( .A(n10107), .B(y[3426]), .Z(n10108) );
  NAND U16177 ( .A(n11222), .B(n10108), .Z(n10109) );
  NAND U16178 ( .A(n10110), .B(n10109), .Z(n10111) );
  NAND U16179 ( .A(n10112), .B(n10111), .Z(n10113) );
  AND U16180 ( .A(n18885), .B(n10113), .Z(n10115) );
  XNOR U16181 ( .A(y[3428]), .B(n10115), .Z(n10114) );
  NANDN U16182 ( .A(x[3428]), .B(n10114), .Z(n10117) );
  NANDN U16183 ( .A(n10115), .B(y[3428]), .Z(n10116) );
  AND U16184 ( .A(n10117), .B(n10116), .Z(n10118) );
  NAND U16185 ( .A(n10119), .B(n10118), .Z(n10120) );
  NAND U16186 ( .A(n10121), .B(n10120), .Z(n10122) );
  AND U16187 ( .A(n20227), .B(n10122), .Z(n10123) );
  ANDN U16188 ( .B(y[3430]), .A(x[3430]), .Z(n11217) );
  ANDN U16189 ( .B(n10123), .A(n11217), .Z(n10124) );
  ANDN U16190 ( .B(x[3431]), .A(y[3431]), .Z(n18890) );
  NOR U16191 ( .A(n10124), .B(n18890), .Z(n10125) );
  XNOR U16192 ( .A(x[3432]), .B(y[3432]), .Z(n18894) );
  NAND U16193 ( .A(n10125), .B(n18894), .Z(n10126) );
  NANDN U16194 ( .A(x[3432]), .B(y[3432]), .Z(n20226) );
  NAND U16195 ( .A(n10126), .B(n20226), .Z(n10127) );
  ANDN U16196 ( .B(x[3435]), .A(y[3435]), .Z(n11212) );
  ANDN U16197 ( .B(x[3437]), .A(y[3437]), .Z(n18904) );
  ANDN U16198 ( .B(x[3438]), .A(y[3438]), .Z(n18909) );
  ANDN U16199 ( .B(x[3441]), .A(y[3441]), .Z(n18912) );
  IV U16200 ( .A(n18912), .Z(n10130) );
  ANDN U16201 ( .B(x[3442]), .A(y[3442]), .Z(n11204) );
  ANDN U16202 ( .B(x[3445]), .A(y[3445]), .Z(n18920) );
  ANDN U16203 ( .B(x[3446]), .A(y[3446]), .Z(n11202) );
  NANDN U16204 ( .A(y[3449]), .B(x[3449]), .Z(n18929) );
  ANDN U16205 ( .B(x[3450]), .A(y[3450]), .Z(n18932) );
  ANDN U16206 ( .B(x[3453]), .A(y[3453]), .Z(n18936) );
  ANDN U16207 ( .B(x[3454]), .A(y[3454]), .Z(n11194) );
  ANDN U16208 ( .B(x[3457]), .A(y[3457]), .Z(n18946) );
  IV U16209 ( .A(n18946), .Z(n10135) );
  ANDN U16210 ( .B(x[3458]), .A(y[3458]), .Z(n18951) );
  ANDN U16211 ( .B(x[3461]), .A(y[3461]), .Z(n18954) );
  ANDN U16212 ( .B(x[3462]), .A(y[3462]), .Z(n11186) );
  ANDN U16213 ( .B(x[3465]), .A(y[3465]), .Z(n18962) );
  ANDN U16214 ( .B(x[3466]), .A(y[3466]), .Z(n11184) );
  ANDN U16215 ( .B(x[3469]), .A(y[3469]), .Z(n18971) );
  ANDN U16216 ( .B(y[3472]), .A(x[3472]), .Z(n18979) );
  NANDN U16217 ( .A(x[3474]), .B(y[3474]), .Z(n11176) );
  ANDN U16218 ( .B(y[3475]), .A(x[3475]), .Z(n11172) );
  ANDN U16219 ( .B(x[3475]), .A(y[3475]), .Z(n11174) );
  IV U16220 ( .A(y[3476]), .Z(n18985) );
  NANDN U16221 ( .A(x[3477]), .B(y[3477]), .Z(n27427) );
  ANDN U16222 ( .B(y[3479]), .A(x[3479]), .Z(n18997) );
  NANDN U16223 ( .A(y[3485]), .B(x[3485]), .Z(n19008) );
  ANDN U16224 ( .B(y[3487]), .A(x[3487]), .Z(n11160) );
  NANDN U16225 ( .A(y[3488]), .B(x[3488]), .Z(n10143) );
  NANDN U16226 ( .A(y[3489]), .B(x[3489]), .Z(n10142) );
  AND U16227 ( .A(n10143), .B(n10142), .Z(n27450) );
  NANDN U16228 ( .A(y[3490]), .B(x[3490]), .Z(n10145) );
  NANDN U16229 ( .A(y[3491]), .B(x[3491]), .Z(n10144) );
  AND U16230 ( .A(n10145), .B(n10144), .Z(n27455) );
  NANDN U16231 ( .A(x[3492]), .B(y[3492]), .Z(n10147) );
  NANDN U16232 ( .A(x[3491]), .B(y[3491]), .Z(n10146) );
  AND U16233 ( .A(n10147), .B(n10146), .Z(n27456) );
  NANDN U16234 ( .A(y[3492]), .B(x[3492]), .Z(n10149) );
  NANDN U16235 ( .A(y[3493]), .B(x[3493]), .Z(n10148) );
  AND U16236 ( .A(n10149), .B(n10148), .Z(n27459) );
  NANDN U16237 ( .A(x[3498]), .B(y[3498]), .Z(n19027) );
  NANDN U16238 ( .A(x[3501]), .B(y[3501]), .Z(n27478) );
  ANDN U16239 ( .B(y[3500]), .A(x[3500]), .Z(n11152) );
  XNOR U16240 ( .A(x[3502]), .B(y[3502]), .Z(n11148) );
  NANDN U16241 ( .A(x[3502]), .B(y[3502]), .Z(n27476) );
  ANDN U16242 ( .B(y[3503]), .A(x[3503]), .Z(n11144) );
  ANDN U16243 ( .B(y[3504]), .A(x[3504]), .Z(n11145) );
  ANDN U16244 ( .B(y[3506]), .A(x[3506]), .Z(n19037) );
  ANDN U16245 ( .B(y[3507]), .A(x[3507]), .Z(n19041) );
  ANDN U16246 ( .B(y[3508]), .A(x[3508]), .Z(n19042) );
  NANDN U16247 ( .A(y[3513]), .B(x[3513]), .Z(n19053) );
  NANDN U16248 ( .A(y[3515]), .B(x[3515]), .Z(n11132) );
  ANDN U16249 ( .B(y[3521]), .A(x[3521]), .Z(n11124) );
  ANDN U16250 ( .B(x[3521]), .A(y[3521]), .Z(n11126) );
  NANDN U16251 ( .A(y[3522]), .B(x[3522]), .Z(n19071) );
  ANDN U16252 ( .B(y[3522]), .A(x[3522]), .Z(n11123) );
  ANDN U16253 ( .B(x[3523]), .A(y[3523]), .Z(n19072) );
  XNOR U16254 ( .A(x[3524]), .B(y[3524]), .Z(n19075) );
  ANDN U16255 ( .B(y[3524]), .A(x[3524]), .Z(n27522) );
  ANDN U16256 ( .B(y[3529]), .A(x[3529]), .Z(n11118) );
  ANDN U16257 ( .B(x[3529]), .A(y[3529]), .Z(n11120) );
  NANDN U16258 ( .A(y[3530]), .B(x[3530]), .Z(n19090) );
  ANDN U16259 ( .B(y[3532]), .A(x[3532]), .Z(n27540) );
  XNOR U16260 ( .A(y[3538]), .B(n10157), .Z(n10156) );
  ANDN U16261 ( .B(y[3539]), .A(x[3539]), .Z(n11111) );
  ANDN U16262 ( .B(x[3539]), .A(y[3539]), .Z(n19112) );
  NANDN U16263 ( .A(y[3540]), .B(x[3540]), .Z(n11108) );
  ANDN U16264 ( .B(y[3540]), .A(x[3540]), .Z(n11110) );
  ANDN U16265 ( .B(x[3541]), .A(y[3541]), .Z(n11109) );
  NANDN U16266 ( .A(y[3549]), .B(x[3549]), .Z(n11097) );
  ANDN U16267 ( .B(y[3557]), .A(x[3557]), .Z(n11083) );
  ANDN U16268 ( .B(x[3557]), .A(y[3557]), .Z(n11084) );
  NANDN U16269 ( .A(y[3558]), .B(x[3558]), .Z(n11080) );
  NANDN U16270 ( .A(n11084), .B(n11080), .Z(n10161) );
  ANDN U16271 ( .B(y[3558]), .A(x[3558]), .Z(n11082) );
  XNOR U16272 ( .A(x[3560]), .B(y[3560]), .Z(n19147) );
  ANDN U16273 ( .B(x[3559]), .A(y[3559]), .Z(n11081) );
  ANDN U16274 ( .B(y[3563]), .A(x[3563]), .Z(n19156) );
  ANDN U16275 ( .B(x[3563]), .A(y[3563]), .Z(n11078) );
  ANDN U16276 ( .B(x[3564]), .A(y[3564]), .Z(n11076) );
  ANDN U16277 ( .B(y[3564]), .A(x[3564]), .Z(n19157) );
  ANDN U16278 ( .B(y[3565]), .A(x[3565]), .Z(n19160) );
  ANDN U16279 ( .B(x[3565]), .A(y[3565]), .Z(n11077) );
  XNOR U16280 ( .A(x[3567]), .B(n10164), .Z(n10163) );
  NANDN U16281 ( .A(x[3568]), .B(y[3568]), .Z(n19165) );
  NANDN U16282 ( .A(x[3571]), .B(y[3571]), .Z(n27628) );
  ANDN U16283 ( .B(y[3570]), .A(x[3570]), .Z(n11070) );
  XNOR U16284 ( .A(x[3572]), .B(y[3572]), .Z(n11066) );
  NANDN U16285 ( .A(x[3572]), .B(y[3572]), .Z(n27626) );
  ANDN U16286 ( .B(y[3573]), .A(x[3573]), .Z(n19174) );
  ANDN U16287 ( .B(y[3574]), .A(x[3574]), .Z(n19173) );
  ANDN U16288 ( .B(y[3576]), .A(x[3576]), .Z(n19179) );
  IV U16289 ( .A(n19179), .Z(n10167) );
  ANDN U16290 ( .B(y[3577]), .A(x[3577]), .Z(n11060) );
  ANDN U16291 ( .B(y[3578]), .A(x[3578]), .Z(n11061) );
  ANDN U16292 ( .B(y[3581]), .A(x[3581]), .Z(n11055) );
  ANDN U16293 ( .B(x[3581]), .A(y[3581]), .Z(n19186) );
  NANDN U16294 ( .A(y[3582]), .B(x[3582]), .Z(n11052) );
  ANDN U16295 ( .B(y[3583]), .A(x[3583]), .Z(n27653) );
  ANDN U16296 ( .B(y[3582]), .A(x[3582]), .Z(n11054) );
  ANDN U16297 ( .B(x[3583]), .A(y[3583]), .Z(n11053) );
  XOR U16298 ( .A(x[3584]), .B(y[3584]), .Z(n11051) );
  OR U16299 ( .A(n11053), .B(n11051), .Z(n10168) );
  ANDN U16300 ( .B(y[3584]), .A(x[3584]), .Z(n27652) );
  ANDN U16301 ( .B(y[3585]), .A(x[3585]), .Z(n11048) );
  ANDN U16302 ( .B(x[3585]), .A(y[3585]), .Z(n11050) );
  ANDN U16303 ( .B(x[3586]), .A(y[3586]), .Z(n19196) );
  ANDN U16304 ( .B(y[3587]), .A(x[3587]), .Z(n27662) );
  XOR U16305 ( .A(x[3588]), .B(y[3588]), .Z(n11046) );
  ANDN U16306 ( .B(y[3588]), .A(x[3588]), .Z(n27663) );
  NANDN U16307 ( .A(y[3591]), .B(x[3591]), .Z(n11041) );
  XNOR U16308 ( .A(y[3592]), .B(n10171), .Z(n10170) );
  NANDN U16309 ( .A(n10171), .B(y[3592]), .Z(n10172) );
  ANDN U16310 ( .B(y[3595]), .A(x[3595]), .Z(n11035) );
  ANDN U16311 ( .B(x[3595]), .A(y[3595]), .Z(n11037) );
  ANDN U16312 ( .B(x[3596]), .A(y[3596]), .Z(n19214) );
  ANDN U16313 ( .B(y[3597]), .A(x[3597]), .Z(n27687) );
  ANDN U16314 ( .B(y[3596]), .A(x[3596]), .Z(n11034) );
  ANDN U16315 ( .B(x[3597]), .A(y[3597]), .Z(n19213) );
  XOR U16316 ( .A(x[3598]), .B(y[3598]), .Z(n11033) );
  ANDN U16317 ( .B(x[3601]), .A(y[3601]), .Z(n19222) );
  ANDN U16318 ( .B(x[3602]), .A(y[3602]), .Z(n11028) );
  XOR U16319 ( .A(x[3604]), .B(y[3604]), .Z(n11026) );
  ANDN U16320 ( .B(x[3605]), .A(y[3605]), .Z(n19229) );
  NANDN U16321 ( .A(x[3606]), .B(y[3606]), .Z(n27707) );
  ANDN U16322 ( .B(y[3607]), .A(x[3607]), .Z(n19236) );
  ANDN U16323 ( .B(x[3607]), .A(y[3607]), .Z(n11024) );
  XNOR U16324 ( .A(x[3609]), .B(n10175), .Z(n10174) );
  XNOR U16325 ( .A(x[3615]), .B(n10177), .Z(n10176) );
  NANDN U16326 ( .A(n10177), .B(x[3615]), .Z(n10178) );
  IV U16327 ( .A(y[3617]), .Z(n11012) );
  NANDN U16328 ( .A(x[3619]), .B(y[3619]), .Z(n27737) );
  ANDN U16329 ( .B(y[3618]), .A(x[3618]), .Z(n11011) );
  XNOR U16330 ( .A(x[3620]), .B(y[3620]), .Z(n19261) );
  NANDN U16331 ( .A(x[3620]), .B(y[3620]), .Z(n27736) );
  ANDN U16332 ( .B(y[3621]), .A(x[3621]), .Z(n19264) );
  ANDN U16333 ( .B(y[3622]), .A(x[3622]), .Z(n19265) );
  ANDN U16334 ( .B(y[3624]), .A(x[3624]), .Z(n19270) );
  IV U16335 ( .A(n19270), .Z(n10181) );
  ANDN U16336 ( .B(y[3625]), .A(x[3625]), .Z(n11005) );
  ANDN U16337 ( .B(y[3627]), .A(x[3627]), .Z(n27755) );
  XOR U16338 ( .A(x[3628]), .B(y[3628]), .Z(n11001) );
  ANDN U16339 ( .B(x[3629]), .A(y[3629]), .Z(n19278) );
  ANDN U16340 ( .B(x[3630]), .A(y[3630]), .Z(n19285) );
  ANDN U16341 ( .B(y[3633]), .A(x[3633]), .Z(n19291) );
  ANDN U16342 ( .B(x[3633]), .A(y[3633]), .Z(n10999) );
  ANDN U16343 ( .B(x[3634]), .A(y[3634]), .Z(n19294) );
  ANDN U16344 ( .B(y[3634]), .A(x[3634]), .Z(n19292) );
  ANDN U16345 ( .B(y[3635]), .A(x[3635]), .Z(n19297) );
  ANDN U16346 ( .B(x[3635]), .A(y[3635]), .Z(n19295) );
  XNOR U16347 ( .A(x[3639]), .B(n10184), .Z(n10183) );
  NANDN U16348 ( .A(n10184), .B(x[3639]), .Z(n10185) );
  NANDN U16349 ( .A(x[3643]), .B(y[3643]), .Z(n27789) );
  ANDN U16350 ( .B(y[3642]), .A(x[3642]), .Z(n10989) );
  XNOR U16351 ( .A(x[3644]), .B(y[3644]), .Z(n19309) );
  NANDN U16352 ( .A(x[3644]), .B(y[3644]), .Z(n27788) );
  ANDN U16353 ( .B(y[3645]), .A(x[3645]), .Z(n19313) );
  ANDN U16354 ( .B(y[3646]), .A(x[3646]), .Z(n19314) );
  ANDN U16355 ( .B(y[3648]), .A(x[3648]), .Z(n19319) );
  ANDN U16356 ( .B(y[3649]), .A(x[3649]), .Z(n10981) );
  ANDN U16357 ( .B(y[3650]), .A(x[3650]), .Z(n10980) );
  ANDN U16358 ( .B(x[3651]), .A(y[3651]), .Z(n10978) );
  XNOR U16359 ( .A(x[3652]), .B(y[3652]), .Z(n19326) );
  ANDN U16360 ( .B(x[3655]), .A(y[3655]), .Z(n19332) );
  ANDN U16361 ( .B(x[3656]), .A(y[3656]), .Z(n10975) );
  NAND U16362 ( .A(n10188), .B(n10187), .Z(n10189) );
  NANDN U16363 ( .A(n10190), .B(n10189), .Z(n10191) );
  AND U16364 ( .A(n19341), .B(n10191), .Z(n10192) );
  NANDN U16365 ( .A(n10974), .B(n10192), .Z(n10193) );
  ANDN U16366 ( .B(y[3659]), .A(x[3659]), .Z(n10970) );
  ANDN U16367 ( .B(n10193), .A(n10970), .Z(n10194) );
  NANDN U16368 ( .A(n27822), .B(n10194), .Z(n10195) );
  ANDN U16369 ( .B(x[3659]), .A(y[3659]), .Z(n10973) );
  ANDN U16370 ( .B(n10195), .A(n10973), .Z(n10196) );
  OR U16371 ( .A(n10971), .B(n10196), .Z(n10197) );
  NANDN U16372 ( .A(n27830), .B(n10197), .Z(n10198) );
  NANDN U16373 ( .A(n10969), .B(n10198), .Z(n10199) );
  NANDN U16374 ( .A(n10967), .B(n10199), .Z(n10200) );
  AND U16375 ( .A(n27838), .B(n10200), .Z(n10201) );
  ANDN U16376 ( .B(y[3662]), .A(x[3662]), .Z(n10968) );
  ANDN U16377 ( .B(n10201), .A(n10968), .Z(n10202) );
  ANDN U16378 ( .B(x[3663]), .A(y[3663]), .Z(n10966) );
  NOR U16379 ( .A(n10202), .B(n10966), .Z(n10204) );
  XNOR U16380 ( .A(x[3664]), .B(y[3664]), .Z(n10203) );
  NAND U16381 ( .A(n10204), .B(n10203), .Z(n10205) );
  AND U16382 ( .A(n27836), .B(n10205), .Z(n10206) );
  NAND U16383 ( .A(n10207), .B(n10206), .Z(n10208) );
  NANDN U16384 ( .A(x[3666]), .B(y[3666]), .Z(n19353) );
  ANDN U16385 ( .B(y[3667]), .A(x[3667]), .Z(n10960) );
  ANDN U16386 ( .B(y[3668]), .A(x[3668]), .Z(n10961) );
  NANDN U16387 ( .A(y[3671]), .B(x[3671]), .Z(n19362) );
  NANDN U16388 ( .A(y[3673]), .B(x[3673]), .Z(n10954) );
  NANDN U16389 ( .A(y[3681]), .B(x[3681]), .Z(n19383) );
  NANDN U16390 ( .A(y[3683]), .B(x[3683]), .Z(n10943) );
  NANDN U16391 ( .A(y[3691]), .B(x[3691]), .Z(n19404) );
  NANDN U16392 ( .A(y[3693]), .B(x[3693]), .Z(n10932) );
  ANDN U16393 ( .B(y[3697]), .A(x[3697]), .Z(n10926) );
  ANDN U16394 ( .B(x[3697]), .A(y[3697]), .Z(n19413) );
  ANDN U16395 ( .B(x[3698]), .A(y[3698]), .Z(n10924) );
  ANDN U16396 ( .B(y[3699]), .A(x[3699]), .Z(n27913) );
  XOR U16397 ( .A(x[3700]), .B(y[3700]), .Z(n19418) );
  ANDN U16398 ( .B(y[3709]), .A(x[3709]), .Z(n19450) );
  ANDN U16399 ( .B(x[3709]), .A(y[3709]), .Z(n10922) );
  ANDN U16400 ( .B(x[3710]), .A(y[3710]), .Z(n19453) );
  ANDN U16401 ( .B(y[3711]), .A(x[3711]), .Z(n27937) );
  ANDN U16402 ( .B(y[3710]), .A(x[3710]), .Z(n19449) );
  ANDN U16403 ( .B(x[3711]), .A(y[3711]), .Z(n19452) );
  XOR U16404 ( .A(x[3712]), .B(y[3712]), .Z(n10920) );
  OR U16405 ( .A(n19452), .B(n10920), .Z(n10216) );
  ANDN U16406 ( .B(y[3712]), .A(x[3712]), .Z(n27936) );
  ANDN U16407 ( .B(y[3717]), .A(x[3717]), .Z(n10915) );
  ANDN U16408 ( .B(x[3717]), .A(y[3717]), .Z(n10917) );
  ANDN U16409 ( .B(x[3718]), .A(y[3718]), .Z(n19471) );
  ANDN U16410 ( .B(y[3719]), .A(x[3719]), .Z(n27954) );
  XOR U16411 ( .A(x[3720]), .B(y[3720]), .Z(n10913) );
  ANDN U16412 ( .B(y[3720]), .A(x[3720]), .Z(n27955) );
  ANDN U16413 ( .B(y[3723]), .A(x[3723]), .Z(n19481) );
  ANDN U16414 ( .B(x[3723]), .A(y[3723]), .Z(n10910) );
  ANDN U16415 ( .B(x[3724]), .A(y[3724]), .Z(n19484) );
  ANDN U16416 ( .B(y[3725]), .A(x[3725]), .Z(n27971) );
  ANDN U16417 ( .B(y[3724]), .A(x[3724]), .Z(n19480) );
  ANDN U16418 ( .B(x[3725]), .A(y[3725]), .Z(n19483) );
  XOR U16419 ( .A(x[3726]), .B(y[3726]), .Z(n10908) );
  ANDN U16420 ( .B(y[3727]), .A(x[3727]), .Z(n27977) );
  XOR U16421 ( .A(x[3728]), .B(y[3728]), .Z(n10907) );
  NANDN U16422 ( .A(y[3735]), .B(x[3735]), .Z(n19502) );
  ANDN U16423 ( .B(y[3737]), .A(x[3737]), .Z(n10890) );
  ANDN U16424 ( .B(x[3737]), .A(y[3737]), .Z(n10892) );
  NANDN U16425 ( .A(y[3738]), .B(x[3738]), .Z(n19507) );
  ANDN U16426 ( .B(y[3739]), .A(x[3739]), .Z(n20220) );
  ANDN U16427 ( .B(y[3738]), .A(x[3738]), .Z(n10889) );
  ANDN U16428 ( .B(x[3739]), .A(y[3739]), .Z(n19508) );
  XOR U16429 ( .A(x[3740]), .B(y[3740]), .Z(n19510) );
  ANDN U16430 ( .B(y[3740]), .A(x[3740]), .Z(n20221) );
  ANDN U16431 ( .B(y[3743]), .A(x[3743]), .Z(n10884) );
  ANDN U16432 ( .B(x[3743]), .A(y[3743]), .Z(n19515) );
  NANDN U16433 ( .A(y[3744]), .B(x[3744]), .Z(n19519) );
  ANDN U16434 ( .B(y[3745]), .A(x[3745]), .Z(n20219) );
  ANDN U16435 ( .B(y[3744]), .A(x[3744]), .Z(n10883) );
  XOR U16436 ( .A(x[3746]), .B(y[3746]), .Z(n19522) );
  ANDN U16437 ( .B(x[3745]), .A(y[3745]), .Z(n19520) );
  XOR U16438 ( .A(x[3748]), .B(y[3748]), .Z(n10880) );
  ANDN U16439 ( .B(y[3749]), .A(x[3749]), .Z(n19531) );
  ANDN U16440 ( .B(x[3749]), .A(y[3749]), .Z(n19528) );
  ANDN U16441 ( .B(x[3750]), .A(y[3750]), .Z(n19535) );
  ANDN U16442 ( .B(y[3750]), .A(x[3750]), .Z(n19532) );
  IV U16443 ( .A(n19532), .Z(n10223) );
  ANDN U16444 ( .B(y[3751]), .A(x[3751]), .Z(n19537) );
  ANDN U16445 ( .B(x[3751]), .A(y[3751]), .Z(n19534) );
  NANDN U16446 ( .A(x[3763]), .B(y[3763]), .Z(n20217) );
  ANDN U16447 ( .B(y[3762]), .A(x[3762]), .Z(n19557) );
  ANDN U16448 ( .B(n20217), .A(n19557), .Z(n10226) );
  XNOR U16449 ( .A(x[3764]), .B(y[3764]), .Z(n10864) );
  NANDN U16450 ( .A(x[3764]), .B(y[3764]), .Z(n20216) );
  ANDN U16451 ( .B(y[3765]), .A(x[3765]), .Z(n19564) );
  ANDN U16452 ( .B(y[3766]), .A(x[3766]), .Z(n19565) );
  ANDN U16453 ( .B(y[3768]), .A(x[3768]), .Z(n19570) );
  ANDN U16454 ( .B(y[3769]), .A(x[3769]), .Z(n10859) );
  ANDN U16455 ( .B(y[3770]), .A(x[3770]), .Z(n10858) );
  ANDN U16456 ( .B(x[3771]), .A(y[3771]), .Z(n19575) );
  XOR U16457 ( .A(x[3772]), .B(y[3772]), .Z(n10857) );
  OR U16458 ( .A(n19575), .B(n10857), .Z(n10229) );
  ANDN U16459 ( .B(y[3775]), .A(x[3775]), .Z(n19586) );
  ANDN U16460 ( .B(x[3775]), .A(y[3775]), .Z(n10854) );
  ANDN U16461 ( .B(x[3776]), .A(y[3776]), .Z(n19589) );
  ANDN U16462 ( .B(y[3777]), .A(x[3777]), .Z(n28083) );
  XOR U16463 ( .A(x[3778]), .B(y[3778]), .Z(n10852) );
  NANDN U16464 ( .A(y[3789]), .B(x[3789]), .Z(n19617) );
  ANDN U16465 ( .B(y[3791]), .A(x[3791]), .Z(n10839) );
  ANDN U16466 ( .B(x[3791]), .A(y[3791]), .Z(n19621) );
  NANDN U16467 ( .A(y[3792]), .B(x[3792]), .Z(n10836) );
  NANDN U16468 ( .A(n19621), .B(n10836), .Z(n10233) );
  ANDN U16469 ( .B(y[3793]), .A(x[3793]), .Z(n20214) );
  ANDN U16470 ( .B(y[3792]), .A(x[3792]), .Z(n10838) );
  ANDN U16471 ( .B(x[3793]), .A(y[3793]), .Z(n10837) );
  XOR U16472 ( .A(x[3794]), .B(y[3794]), .Z(n10835) );
  ANDN U16473 ( .B(y[3796]), .A(x[3796]), .Z(n28118) );
  XNOR U16474 ( .A(y[3800]), .B(n10236), .Z(n10235) );
  IV U16475 ( .A(x[3806]), .Z(n10818) );
  XNOR U16476 ( .A(n10237), .B(y[3806]), .Z(n10238) );
  NAND U16477 ( .A(n10818), .B(n10238), .Z(n10239) );
  IV U16478 ( .A(x[3807]), .Z(n10815) );
  ANDN U16479 ( .B(y[3808]), .A(x[3808]), .Z(n10817) );
  NANDN U16480 ( .A(y[3808]), .B(x[3808]), .Z(n10241) );
  NANDN U16481 ( .A(y[3809]), .B(x[3809]), .Z(n10240) );
  AND U16482 ( .A(n10241), .B(n10240), .Z(n28147) );
  NANDN U16483 ( .A(x[3810]), .B(y[3810]), .Z(n10243) );
  NANDN U16484 ( .A(x[3809]), .B(y[3809]), .Z(n10242) );
  AND U16485 ( .A(n10243), .B(n10242), .Z(n28148) );
  NANDN U16486 ( .A(y[3811]), .B(x[3811]), .Z(n10245) );
  NANDN U16487 ( .A(y[3810]), .B(x[3810]), .Z(n10244) );
  NAND U16488 ( .A(n10245), .B(n10244), .Z(n28150) );
  XOR U16489 ( .A(x[3814]), .B(y[3814]), .Z(n10812) );
  XNOR U16490 ( .A(y[3816]), .B(n10247), .Z(n10246) );
  NAND U16491 ( .A(n10809), .B(n10246), .Z(n10249) );
  NANDN U16492 ( .A(n10247), .B(y[3816]), .Z(n10248) );
  AND U16493 ( .A(n10249), .B(n10248), .Z(n10250) );
  ANDN U16494 ( .B(y[3817]), .A(x[3817]), .Z(n19668) );
  ANDN U16495 ( .B(n10250), .A(n19668), .Z(n10253) );
  ANDN U16496 ( .B(x[3817]), .A(y[3817]), .Z(n10807) );
  ANDN U16497 ( .B(x[3818]), .A(y[3818]), .Z(n19671) );
  IV U16498 ( .A(n19671), .Z(n10251) );
  NANDN U16499 ( .A(n10807), .B(n10251), .Z(n10252) );
  OR U16500 ( .A(n10253), .B(n10252), .Z(n10254) );
  AND U16501 ( .A(n28172), .B(n10254), .Z(n10255) );
  ANDN U16502 ( .B(y[3818]), .A(x[3818]), .Z(n19667) );
  ANDN U16503 ( .B(n10255), .A(n19667), .Z(n10257) );
  ANDN U16504 ( .B(x[3819]), .A(y[3819]), .Z(n19670) );
  XOR U16505 ( .A(x[3820]), .B(y[3820]), .Z(n19675) );
  OR U16506 ( .A(n19670), .B(n19675), .Z(n10256) );
  OR U16507 ( .A(n10257), .B(n10256), .Z(n10258) );
  ANDN U16508 ( .B(y[3821]), .A(x[3821]), .Z(n28178) );
  ANDN U16509 ( .B(n10258), .A(n28178), .Z(n10259) );
  ANDN U16510 ( .B(y[3820]), .A(x[3820]), .Z(n28170) );
  ANDN U16511 ( .B(n10259), .A(n28170), .Z(n10261) );
  XOR U16512 ( .A(x[3822]), .B(y[3822]), .Z(n10804) );
  ANDN U16513 ( .B(x[3821]), .A(y[3821]), .Z(n10806) );
  NOR U16514 ( .A(n10804), .B(n10806), .Z(n10260) );
  NANDN U16515 ( .A(n10261), .B(n10260), .Z(n10262) );
  NAND U16516 ( .A(n10263), .B(n10262), .Z(n10264) );
  XOR U16517 ( .A(x[3824]), .B(y[3824]), .Z(n19680) );
  ANDN U16518 ( .B(n10264), .A(n19680), .Z(n10265) );
  NANDN U16519 ( .A(n10803), .B(n10265), .Z(n10266) );
  ANDN U16520 ( .B(y[3825]), .A(x[3825]), .Z(n10799) );
  ANDN U16521 ( .B(n10266), .A(n10799), .Z(n10267) );
  NANDN U16522 ( .A(n28182), .B(n10267), .Z(n10268) );
  ANDN U16523 ( .B(x[3825]), .A(y[3825]), .Z(n10801) );
  ANDN U16524 ( .B(n10268), .A(n10801), .Z(n10269) );
  NANDN U16525 ( .A(n10797), .B(n10269), .Z(n10270) );
  XOR U16526 ( .A(x[3828]), .B(y[3828]), .Z(n10795) );
  NANDN U16527 ( .A(x[3828]), .B(y[3828]), .Z(n20213) );
  NANDN U16528 ( .A(x[3831]), .B(y[3831]), .Z(n28202) );
  ANDN U16529 ( .B(y[3830]), .A(x[3830]), .Z(n10792) );
  XNOR U16530 ( .A(x[3832]), .B(y[3832]), .Z(n10788) );
  NANDN U16531 ( .A(x[3832]), .B(y[3832]), .Z(n28200) );
  ANDN U16532 ( .B(y[3833]), .A(x[3833]), .Z(n19694) );
  ANDN U16533 ( .B(y[3834]), .A(x[3834]), .Z(n19695) );
  ANDN U16534 ( .B(y[3836]), .A(x[3836]), .Z(n19700) );
  ANDN U16535 ( .B(y[3837]), .A(x[3837]), .Z(n19704) );
  ANDN U16536 ( .B(y[3838]), .A(x[3838]), .Z(n19705) );
  NANDN U16537 ( .A(n10272), .B(y[3842]), .Z(n10275) );
  XNOR U16538 ( .A(n10272), .B(y[3842]), .Z(n10273) );
  NANDN U16539 ( .A(x[3842]), .B(n10273), .Z(n10274) );
  NAND U16540 ( .A(n10275), .B(n10274), .Z(n10276) );
  ANDN U16541 ( .B(x[3843]), .A(y[3843]), .Z(n10781) );
  ANDN U16542 ( .B(n10276), .A(n10781), .Z(n10279) );
  NANDN U16543 ( .A(x[3843]), .B(y[3843]), .Z(n10278) );
  NANDN U16544 ( .A(x[3844]), .B(y[3844]), .Z(n10277) );
  AND U16545 ( .A(n10278), .B(n10277), .Z(n28226) );
  NANDN U16546 ( .A(n10279), .B(n28226), .Z(n10280) );
  NANDN U16547 ( .A(n28228), .B(n10280), .Z(n10281) );
  NANDN U16548 ( .A(n10778), .B(n10281), .Z(n10282) );
  NANDN U16549 ( .A(n19723), .B(n10282), .Z(n10283) );
  ANDN U16550 ( .B(y[3846]), .A(x[3846]), .Z(n10779) );
  ANDN U16551 ( .B(n10283), .A(n10779), .Z(n10284) );
  NAND U16552 ( .A(n10285), .B(n10284), .Z(n10286) );
  NAND U16553 ( .A(n10287), .B(n10286), .Z(n10288) );
  ANDN U16554 ( .B(y[3848]), .A(x[3848]), .Z(n10777) );
  ANDN U16555 ( .B(n10288), .A(n10777), .Z(n10289) );
  NAND U16556 ( .A(n10290), .B(n10289), .Z(n10291) );
  AND U16557 ( .A(n10292), .B(n10291), .Z(n10294) );
  NANDN U16558 ( .A(x[3851]), .B(y[3851]), .Z(n28244) );
  ANDN U16559 ( .B(y[3850]), .A(x[3850]), .Z(n10773) );
  ANDN U16560 ( .B(n28244), .A(n10773), .Z(n10293) );
  NANDN U16561 ( .A(n10294), .B(n10293), .Z(n10295) );
  ANDN U16562 ( .B(y[3852]), .A(x[3852]), .Z(n28242) );
  XNOR U16563 ( .A(y[3858]), .B(n10297), .Z(n10296) );
  ANDN U16564 ( .B(y[3859]), .A(x[3859]), .Z(n10755) );
  ANDN U16565 ( .B(x[3859]), .A(y[3859]), .Z(n10756) );
  ANDN U16566 ( .B(x[3860]), .A(y[3860]), .Z(n19743) );
  ANDN U16567 ( .B(y[3861]), .A(x[3861]), .Z(n28267) );
  ANDN U16568 ( .B(y[3860]), .A(x[3860]), .Z(n10754) );
  ANDN U16569 ( .B(x[3861]), .A(y[3861]), .Z(n19742) );
  XOR U16570 ( .A(x[3862]), .B(y[3862]), .Z(n10753) );
  ANDN U16571 ( .B(y[3862]), .A(x[3862]), .Z(n28264) );
  NANDN U16572 ( .A(n10728), .B(n10303), .Z(n10304) );
  NANDN U16573 ( .A(y[3883]), .B(x[3883]), .Z(n19789) );
  NAND U16574 ( .A(n10304), .B(n19789), .Z(n10306) );
  XNOR U16575 ( .A(y[3884]), .B(n10306), .Z(n10305) );
  NAND U16576 ( .A(n10726), .B(n10305), .Z(n10308) );
  NANDN U16577 ( .A(n10306), .B(y[3884]), .Z(n10307) );
  AND U16578 ( .A(n10308), .B(n10307), .Z(n10309) );
  NANDN U16579 ( .A(n10725), .B(n10309), .Z(n10310) );
  NANDN U16580 ( .A(y[3885]), .B(x[3885]), .Z(n19793) );
  NAND U16581 ( .A(n10310), .B(n19793), .Z(n10312) );
  XNOR U16582 ( .A(y[3886]), .B(n10312), .Z(n10311) );
  NANDN U16583 ( .A(x[3886]), .B(n10311), .Z(n10314) );
  NANDN U16584 ( .A(n10312), .B(y[3886]), .Z(n10313) );
  AND U16585 ( .A(n10314), .B(n10313), .Z(n10315) );
  NANDN U16586 ( .A(n10721), .B(n10315), .Z(n10316) );
  NANDN U16587 ( .A(y[3887]), .B(x[3887]), .Z(n10723) );
  NAND U16588 ( .A(n10316), .B(n10723), .Z(n10318) );
  XNOR U16589 ( .A(y[3888]), .B(n10318), .Z(n10317) );
  NAND U16590 ( .A(n10719), .B(n10317), .Z(n10320) );
  NANDN U16591 ( .A(n10318), .B(y[3888]), .Z(n10319) );
  AND U16592 ( .A(n10320), .B(n10319), .Z(n10321) );
  NANDN U16593 ( .A(n10716), .B(n10321), .Z(n10322) );
  ANDN U16594 ( .B(x[3889]), .A(y[3889]), .Z(n10717) );
  ANDN U16595 ( .B(n10322), .A(n10717), .Z(n10323) );
  XOR U16596 ( .A(x[3892]), .B(y[3892]), .Z(n10712) );
  ANDN U16597 ( .B(x[3891]), .A(y[3891]), .Z(n10713) );
  ANDN U16598 ( .B(x[3893]), .A(y[3893]), .Z(n19803) );
  IV U16599 ( .A(y[3894]), .Z(n10707) );
  XOR U16600 ( .A(x[3896]), .B(y[3896]), .Z(n19808) );
  ANDN U16601 ( .B(y[3897]), .A(x[3897]), .Z(n28341) );
  XOR U16602 ( .A(x[3898]), .B(y[3898]), .Z(n10704) );
  XOR U16603 ( .A(x[3900]), .B(y[3900]), .Z(n10701) );
  NANDN U16604 ( .A(x[3900]), .B(y[3900]), .Z(n28347) );
  NANDN U16605 ( .A(x[3903]), .B(y[3903]), .Z(n28357) );
  ANDN U16606 ( .B(y[3902]), .A(x[3902]), .Z(n10700) );
  XNOR U16607 ( .A(x[3904]), .B(y[3904]), .Z(n10698) );
  NANDN U16608 ( .A(x[3904]), .B(y[3904]), .Z(n28356) );
  ANDN U16609 ( .B(y[3905]), .A(x[3905]), .Z(n10695) );
  ANDN U16610 ( .B(y[3906]), .A(x[3906]), .Z(n10694) );
  ANDN U16611 ( .B(x[3907]), .A(y[3907]), .Z(n19828) );
  XNOR U16612 ( .A(x[3908]), .B(y[3908]), .Z(n10327) );
  IV U16613 ( .A(y[3908]), .Z(n10692) );
  NOR U16614 ( .A(n10692), .B(x[3908]), .Z(n20208) );
  ANDN U16615 ( .B(x[3909]), .A(y[3909]), .Z(n10690) );
  ANDN U16616 ( .B(y[3910]), .A(x[3910]), .Z(n28370) );
  ANDN U16617 ( .B(y[3911]), .A(x[3911]), .Z(n10687) );
  ANDN U16618 ( .B(x[3911]), .A(y[3911]), .Z(n10689) );
  ANDN U16619 ( .B(x[3912]), .A(y[3912]), .Z(n19840) );
  ANDN U16620 ( .B(y[3913]), .A(x[3913]), .Z(n20206) );
  XOR U16621 ( .A(x[3914]), .B(y[3914]), .Z(n10685) );
  ANDN U16622 ( .B(y[3914]), .A(x[3914]), .Z(n20207) );
  XNOR U16623 ( .A(y[3916]), .B(n10329), .Z(n10328) );
  NAND U16624 ( .A(n19847), .B(n10328), .Z(n10331) );
  NANDN U16625 ( .A(n10329), .B(y[3916]), .Z(n10330) );
  ANDN U16626 ( .B(y[3917]), .A(x[3917]), .Z(n10682) );
  ANDN U16627 ( .B(x[3917]), .A(y[3917]), .Z(n10684) );
  ANDN U16628 ( .B(x[3918]), .A(y[3918]), .Z(n19854) );
  ANDN U16629 ( .B(y[3919]), .A(x[3919]), .Z(n20205) );
  ANDN U16630 ( .B(y[3918]), .A(x[3918]), .Z(n10681) );
  ANDN U16631 ( .B(x[3919]), .A(y[3919]), .Z(n19853) );
  XOR U16632 ( .A(x[3920]), .B(y[3920]), .Z(n10680) );
  ANDN U16633 ( .B(y[3920]), .A(x[3920]), .Z(n20204) );
  XNOR U16634 ( .A(y[3924]), .B(n10333), .Z(n10332) );
  NANDN U16635 ( .A(n10333), .B(y[3924]), .Z(n10334) );
  ANDN U16636 ( .B(y[3925]), .A(x[3925]), .Z(n19871) );
  ANDN U16637 ( .B(x[3925]), .A(y[3925]), .Z(n10677) );
  ANDN U16638 ( .B(x[3926]), .A(y[3926]), .Z(n19874) );
  ANDN U16639 ( .B(y[3927]), .A(x[3927]), .Z(n28409) );
  XOR U16640 ( .A(x[3928]), .B(y[3928]), .Z(n10675) );
  ANDN U16641 ( .B(x[3929]), .A(y[3929]), .Z(n19878) );
  ANDN U16642 ( .B(x[3930]), .A(y[3930]), .Z(n10672) );
  XOR U16643 ( .A(x[3932]), .B(y[3932]), .Z(n10670) );
  ANDN U16644 ( .B(y[3933]), .A(x[3933]), .Z(n19887) );
  NANDN U16645 ( .A(n20202), .B(n10335), .Z(n10336) );
  ANDN U16646 ( .B(x[3933]), .A(y[3933]), .Z(n10669) );
  ANDN U16647 ( .B(n10336), .A(n10669), .Z(n10337) );
  ANDN U16648 ( .B(x[3934]), .A(y[3934]), .Z(n10666) );
  ANDN U16649 ( .B(n10337), .A(n10666), .Z(n10339) );
  NANDN U16650 ( .A(x[3934]), .B(y[3934]), .Z(n19886) );
  ANDN U16651 ( .B(y[3935]), .A(x[3935]), .Z(n10665) );
  ANDN U16652 ( .B(n19886), .A(n10665), .Z(n10338) );
  NANDN U16653 ( .A(n10339), .B(n10338), .Z(n10340) );
  ANDN U16654 ( .B(x[3935]), .A(y[3935]), .Z(n10667) );
  ANDN U16655 ( .B(n10340), .A(n10667), .Z(n10341) );
  NANDN U16656 ( .A(n10663), .B(n10341), .Z(n10342) );
  NANDN U16657 ( .A(x[3936]), .B(y[3936]), .Z(n10664) );
  NAND U16658 ( .A(n10342), .B(n10664), .Z(n10344) );
  XNOR U16659 ( .A(x[3937]), .B(n10344), .Z(n10343) );
  NAND U16660 ( .A(n10661), .B(n10343), .Z(n10346) );
  NANDN U16661 ( .A(n10344), .B(x[3937]), .Z(n10345) );
  AND U16662 ( .A(n10346), .B(n10345), .Z(n10347) );
  NANDN U16663 ( .A(n10660), .B(n10347), .Z(n10348) );
  NANDN U16664 ( .A(x[3938]), .B(y[3938]), .Z(n19893) );
  NAND U16665 ( .A(n10348), .B(n19893), .Z(n10350) );
  XNOR U16666 ( .A(x[3939]), .B(n10350), .Z(n10349) );
  NAND U16667 ( .A(n10658), .B(n10349), .Z(n10352) );
  NANDN U16668 ( .A(n10350), .B(x[3939]), .Z(n10351) );
  AND U16669 ( .A(n10352), .B(n10351), .Z(n10353) );
  NANDN U16670 ( .A(n10657), .B(n10353), .Z(n10354) );
  NANDN U16671 ( .A(x[3940]), .B(y[3940]), .Z(n19897) );
  NAND U16672 ( .A(n10354), .B(n19897), .Z(n10356) );
  XNOR U16673 ( .A(x[3941]), .B(n10356), .Z(n10355) );
  NANDN U16674 ( .A(n10356), .B(x[3941]), .Z(n10357) );
  NANDN U16675 ( .A(x[3942]), .B(y[3942]), .Z(n10655) );
  IV U16676 ( .A(y[3943]), .Z(n10651) );
  NANDN U16677 ( .A(x[3945]), .B(y[3945]), .Z(n28448) );
  ANDN U16678 ( .B(y[3944]), .A(x[3944]), .Z(n19903) );
  XNOR U16679 ( .A(x[3946]), .B(y[3946]), .Z(n10648) );
  NANDN U16680 ( .A(x[3946]), .B(y[3946]), .Z(n28447) );
  ANDN U16681 ( .B(y[3947]), .A(x[3947]), .Z(n10645) );
  ANDN U16682 ( .B(y[3948]), .A(x[3948]), .Z(n10644) );
  ANDN U16683 ( .B(x[3949]), .A(y[3949]), .Z(n19910) );
  IV U16684 ( .A(y[3950]), .Z(n19915) );
  NOR U16685 ( .A(n19915), .B(x[3950]), .Z(n28456) );
  ANDN U16686 ( .B(x[3951]), .A(y[3951]), .Z(n19916) );
  XOR U16687 ( .A(x[3952]), .B(y[3952]), .Z(n10642) );
  ANDN U16688 ( .B(y[3953]), .A(x[3953]), .Z(n28470) );
  ANDN U16689 ( .B(y[3952]), .A(x[3952]), .Z(n28462) );
  ANDN U16690 ( .B(x[3953]), .A(y[3953]), .Z(n10641) );
  XOR U16691 ( .A(x[3954]), .B(y[3954]), .Z(n19922) );
  ANDN U16692 ( .B(y[3954]), .A(x[3954]), .Z(n28468) );
  ANDN U16693 ( .B(x[3955]), .A(y[3955]), .Z(n10639) );
  NANDN U16694 ( .A(x[3957]), .B(y[3957]), .Z(n28479) );
  XOR U16695 ( .A(x[3958]), .B(y[3958]), .Z(n19930) );
  ANDN U16696 ( .B(x[3957]), .A(y[3957]), .Z(n10636) );
  XOR U16697 ( .A(x[3960]), .B(y[3960]), .Z(n10633) );
  ANDN U16698 ( .B(y[3961]), .A(x[3961]), .Z(n10630) );
  ANDN U16699 ( .B(x[3961]), .A(y[3961]), .Z(n10632) );
  ANDN U16700 ( .B(x[3962]), .A(y[3962]), .Z(n10627) );
  NANDN U16701 ( .A(x[3962]), .B(y[3962]), .Z(n10629) );
  ANDN U16702 ( .B(y[3963]), .A(x[3963]), .Z(n19940) );
  ANDN U16703 ( .B(x[3963]), .A(y[3963]), .Z(n10628) );
  NANDN U16704 ( .A(x[3964]), .B(y[3964]), .Z(n19939) );
  XNOR U16705 ( .A(x[3967]), .B(n10361), .Z(n10360) );
  NANDN U16706 ( .A(n10361), .B(x[3967]), .Z(n10362) );
  ANDN U16707 ( .B(x[3968]), .A(y[3968]), .Z(n19953) );
  ANDN U16708 ( .B(y[3969]), .A(x[3969]), .Z(n28507) );
  ANDN U16709 ( .B(y[3968]), .A(x[3968]), .Z(n19949) );
  XOR U16710 ( .A(x[3970]), .B(y[3970]), .Z(n10623) );
  ANDN U16711 ( .B(y[3971]), .A(x[3971]), .Z(n28514) );
  XOR U16712 ( .A(x[3972]), .B(y[3972]), .Z(n10622) );
  NANDN U16713 ( .A(x[3972]), .B(y[3972]), .Z(n28513) );
  XNOR U16714 ( .A(x[3975]), .B(n10364), .Z(n10363) );
  NANDN U16715 ( .A(x[3981]), .B(y[3981]), .Z(n28535) );
  ANDN U16716 ( .B(y[3980]), .A(x[3980]), .Z(n19978) );
  XNOR U16717 ( .A(x[3982]), .B(y[3982]), .Z(n10611) );
  NANDN U16718 ( .A(x[3982]), .B(y[3982]), .Z(n28534) );
  ANDN U16719 ( .B(y[3983]), .A(x[3983]), .Z(n10607) );
  ANDN U16720 ( .B(y[3984]), .A(x[3984]), .Z(n10608) );
  NANDN U16721 ( .A(x[3986]), .B(y[3986]), .Z(n19989) );
  ANDN U16722 ( .B(y[3987]), .A(x[3987]), .Z(n19992) );
  ANDN U16723 ( .B(y[3988]), .A(x[3988]), .Z(n19993) );
  XNOR U16724 ( .A(y[3990]), .B(n10367), .Z(n10366) );
  NANDN U16725 ( .A(x[3990]), .B(n10366), .Z(n10369) );
  NANDN U16726 ( .A(n10367), .B(y[3990]), .Z(n10368) );
  NANDN U16727 ( .A(y[3993]), .B(x[3993]), .Z(n20004) );
  NANDN U16728 ( .A(y[3995]), .B(x[3995]), .Z(n20008) );
  NANDN U16729 ( .A(n10593), .B(n10370), .Z(n10371) );
  NANDN U16730 ( .A(y[3997]), .B(x[3997]), .Z(n10595) );
  NAND U16731 ( .A(n10371), .B(n10595), .Z(n10373) );
  XNOR U16732 ( .A(y[3998]), .B(n10373), .Z(n10372) );
  NAND U16733 ( .A(n10591), .B(n10372), .Z(n10375) );
  NANDN U16734 ( .A(n10373), .B(y[3998]), .Z(n10374) );
  AND U16735 ( .A(n10375), .B(n10374), .Z(n10376) );
  NANDN U16736 ( .A(n10590), .B(n10376), .Z(n10377) );
  NANDN U16737 ( .A(y[3999]), .B(x[3999]), .Z(n20014) );
  NAND U16738 ( .A(n10377), .B(n20014), .Z(n10379) );
  XNOR U16739 ( .A(y[4000]), .B(n10379), .Z(n10378) );
  NAND U16740 ( .A(n10588), .B(n10378), .Z(n10381) );
  NANDN U16741 ( .A(n10379), .B(y[4000]), .Z(n10380) );
  AND U16742 ( .A(n10381), .B(n10380), .Z(n10382) );
  NANDN U16743 ( .A(n10587), .B(n10382), .Z(n10383) );
  NANDN U16744 ( .A(y[4001]), .B(x[4001]), .Z(n20018) );
  NAND U16745 ( .A(n10383), .B(n20018), .Z(n10385) );
  XNOR U16746 ( .A(y[4002]), .B(n10385), .Z(n10384) );
  NANDN U16747 ( .A(x[4002]), .B(n10384), .Z(n10387) );
  NANDN U16748 ( .A(n10385), .B(y[4002]), .Z(n10386) );
  AND U16749 ( .A(n10387), .B(n10386), .Z(n10388) );
  ANDN U16750 ( .B(y[4003]), .A(x[4003]), .Z(n10582) );
  ANDN U16751 ( .B(n10388), .A(n10582), .Z(n10389) );
  OR U16752 ( .A(n10585), .B(n10389), .Z(n10390) );
  NANDN U16753 ( .A(n10583), .B(n10390), .Z(n10393) );
  NANDN U16754 ( .A(y[4004]), .B(x[4004]), .Z(n10392) );
  NANDN U16755 ( .A(y[4005]), .B(x[4005]), .Z(n10391) );
  AND U16756 ( .A(n10392), .B(n10391), .Z(n28582) );
  NAND U16757 ( .A(n10393), .B(n28582), .Z(n10394) );
  AND U16758 ( .A(n28584), .B(n10394), .Z(n10397) );
  NANDN U16759 ( .A(y[4006]), .B(x[4006]), .Z(n10396) );
  NANDN U16760 ( .A(y[4007]), .B(x[4007]), .Z(n10395) );
  AND U16761 ( .A(n10396), .B(n10395), .Z(n28587) );
  NANDN U16762 ( .A(n10397), .B(n28587), .Z(n10400) );
  NANDN U16763 ( .A(x[4008]), .B(y[4008]), .Z(n10399) );
  NANDN U16764 ( .A(x[4007]), .B(y[4007]), .Z(n10398) );
  AND U16765 ( .A(n10399), .B(n10398), .Z(n28588) );
  NAND U16766 ( .A(n10400), .B(n28588), .Z(n10403) );
  NANDN U16767 ( .A(y[4008]), .B(x[4008]), .Z(n10402) );
  NANDN U16768 ( .A(y[4009]), .B(x[4009]), .Z(n10401) );
  AND U16769 ( .A(n10402), .B(n10401), .Z(n28590) );
  NAND U16770 ( .A(n10403), .B(n28590), .Z(n10404) );
  ANDN U16771 ( .B(y[4009]), .A(x[4009]), .Z(n10580) );
  ANDN U16772 ( .B(n10404), .A(n10580), .Z(n10405) );
  NAND U16773 ( .A(n10406), .B(n10405), .Z(n10407) );
  NAND U16774 ( .A(n10578), .B(n10407), .Z(n10408) );
  NANDN U16775 ( .A(n20031), .B(n10408), .Z(n10409) );
  ANDN U16776 ( .B(x[4011]), .A(y[4011]), .Z(n10579) );
  ANDN U16777 ( .B(n10409), .A(n10579), .Z(n10410) );
  NANDN U16778 ( .A(n10577), .B(n10410), .Z(n10411) );
  NANDN U16779 ( .A(x[4012]), .B(y[4012]), .Z(n20030) );
  NAND U16780 ( .A(n10411), .B(n20030), .Z(n10413) );
  XNOR U16781 ( .A(x[4013]), .B(n10413), .Z(n10412) );
  NANDN U16782 ( .A(y[4013]), .B(n10412), .Z(n10415) );
  NANDN U16783 ( .A(n10413), .B(x[4013]), .Z(n10414) );
  AND U16784 ( .A(n10415), .B(n10414), .Z(n10416) );
  NANDN U16785 ( .A(n10573), .B(n10416), .Z(n10417) );
  NANDN U16786 ( .A(x[4014]), .B(y[4014]), .Z(n10575) );
  NAND U16787 ( .A(n10417), .B(n10575), .Z(n10418) );
  NANDN U16788 ( .A(x[4016]), .B(y[4016]), .Z(n20037) );
  NANDN U16789 ( .A(n10419), .B(x[4021]), .Z(n10422) );
  XNOR U16790 ( .A(n10419), .B(x[4021]), .Z(n10420) );
  NANDN U16791 ( .A(y[4021]), .B(n10420), .Z(n10421) );
  NAND U16792 ( .A(n10422), .B(n10421), .Z(n10423) );
  OR U16793 ( .A(n20054), .B(n10423), .Z(n10425) );
  NANDN U16794 ( .A(x[4023]), .B(y[4023]), .Z(n28623) );
  ANDN U16795 ( .B(y[4022]), .A(x[4022]), .Z(n10567) );
  ANDN U16796 ( .B(n28623), .A(n10567), .Z(n10424) );
  NAND U16797 ( .A(n10425), .B(n10424), .Z(n10426) );
  NANDN U16798 ( .A(n20053), .B(n10426), .Z(n10427) );
  XNOR U16799 ( .A(x[4024]), .B(y[4024]), .Z(n10565) );
  NANDN U16800 ( .A(n10427), .B(n10565), .Z(n10428) );
  ANDN U16801 ( .B(y[4024]), .A(x[4024]), .Z(n28620) );
  ANDN U16802 ( .B(n10428), .A(n28620), .Z(n10429) );
  NAND U16803 ( .A(n10430), .B(n10429), .Z(n10431) );
  AND U16804 ( .A(n10432), .B(n10431), .Z(n10434) );
  NANDN U16805 ( .A(x[4027]), .B(y[4027]), .Z(n28632) );
  ANDN U16806 ( .B(y[4026]), .A(x[4026]), .Z(n10562) );
  ANDN U16807 ( .B(n28632), .A(n10562), .Z(n10433) );
  NANDN U16808 ( .A(n10434), .B(n10433), .Z(n10435) );
  NANDN U16809 ( .A(n10436), .B(n10435), .Z(n10437) );
  ANDN U16810 ( .B(y[4028]), .A(x[4028]), .Z(n28630) );
  ANDN U16811 ( .B(n10437), .A(n28630), .Z(n10438) );
  NANDN U16812 ( .A(n10555), .B(n10438), .Z(n10439) );
  ANDN U16813 ( .B(x[4029]), .A(y[4029]), .Z(n10556) );
  ANDN U16814 ( .B(y[4030]), .A(x[4030]), .Z(n10554) );
  NAND U16815 ( .A(n10440), .B(n10554), .Z(n10443) );
  NANDN U16816 ( .A(x[4032]), .B(y[4032]), .Z(n10442) );
  NANDN U16817 ( .A(x[4031]), .B(y[4031]), .Z(n10441) );
  NAND U16818 ( .A(n10442), .B(n10441), .Z(n28640) );
  NANDN U16819 ( .A(y[4033]), .B(x[4033]), .Z(n10445) );
  NANDN U16820 ( .A(y[4032]), .B(x[4032]), .Z(n10444) );
  AND U16821 ( .A(n10445), .B(n10444), .Z(n28642) );
  ANDN U16822 ( .B(x[4034]), .A(y[4034]), .Z(n10553) );
  NANDN U16823 ( .A(x[4035]), .B(y[4035]), .Z(n28651) );
  ANDN U16824 ( .B(y[4034]), .A(x[4034]), .Z(n20068) );
  IV U16825 ( .A(y[4036]), .Z(n20075) );
  NOR U16826 ( .A(n20075), .B(x[4036]), .Z(n28648) );
  XNOR U16827 ( .A(x[4038]), .B(y[4038]), .Z(n10551) );
  ANDN U16828 ( .B(x[4037]), .A(y[4037]), .Z(n20076) );
  ANDN U16829 ( .B(y[4038]), .A(x[4038]), .Z(n28654) );
  XNOR U16830 ( .A(y[4040]), .B(n10447), .Z(n10446) );
  XNOR U16831 ( .A(y[4046]), .B(n10449), .Z(n10448) );
  ANDN U16832 ( .B(y[4049]), .A(x[4049]), .Z(n10543) );
  ANDN U16833 ( .B(x[4049]), .A(y[4049]), .Z(n10545) );
  ANDN U16834 ( .B(x[4050]), .A(y[4050]), .Z(n20112) );
  ANDN U16835 ( .B(y[4051]), .A(x[4051]), .Z(n20200) );
  ANDN U16836 ( .B(y[4050]), .A(x[4050]), .Z(n10542) );
  ANDN U16837 ( .B(x[4051]), .A(y[4051]), .Z(n20111) );
  XOR U16838 ( .A(x[4052]), .B(y[4052]), .Z(n10541) );
  ANDN U16839 ( .B(y[4053]), .A(x[4053]), .Z(n28690) );
  XOR U16840 ( .A(x[4054]), .B(y[4054]), .Z(n20117) );
  XNOR U16841 ( .A(y[4060]), .B(n10452), .Z(n10451) );
  NANDN U16842 ( .A(x[4060]), .B(n10451), .Z(n10454) );
  NANDN U16843 ( .A(n10452), .B(y[4060]), .Z(n10453) );
  ANDN U16844 ( .B(y[4063]), .A(x[4063]), .Z(n20140) );
  ANDN U16845 ( .B(x[4063]), .A(y[4063]), .Z(n10529) );
  ANDN U16846 ( .B(x[4064]), .A(y[4064]), .Z(n20143) );
  ANDN U16847 ( .B(y[4064]), .A(x[4064]), .Z(n20139) );
  ANDN U16848 ( .B(x[4065]), .A(y[4065]), .Z(n20142) );
  XOR U16849 ( .A(x[4066]), .B(y[4066]), .Z(n10527) );
  ANDN U16850 ( .B(y[4066]), .A(x[4066]), .Z(n28714) );
  XNOR U16851 ( .A(y[4068]), .B(n10456), .Z(n10455) );
  NAND U16852 ( .A(n10524), .B(n10455), .Z(n10458) );
  NANDN U16853 ( .A(n10456), .B(y[4068]), .Z(n10457) );
  AND U16854 ( .A(n10458), .B(n10457), .Z(n10459) );
  ANDN U16855 ( .B(y[4069]), .A(x[4069]), .Z(n20152) );
  ANDN U16856 ( .B(n10459), .A(n20152), .Z(n10460) );
  NAND U16857 ( .A(n10461), .B(n10460), .Z(n10462) );
  NAND U16858 ( .A(n10520), .B(n10462), .Z(n10463) );
  NANDN U16859 ( .A(n10519), .B(n10463), .Z(n10464) );
  ANDN U16860 ( .B(x[4071]), .A(y[4071]), .Z(n10521) );
  ANDN U16861 ( .B(n10464), .A(n10521), .Z(n10465) );
  NANDN U16862 ( .A(n10517), .B(n10465), .Z(n10466) );
  NANDN U16863 ( .A(n10467), .B(n10466), .Z(n10468) );
  XOR U16864 ( .A(x[4074]), .B(y[4074]), .Z(n10515) );
  ANDN U16865 ( .B(n10468), .A(n10515), .Z(n10469) );
  NANDN U16866 ( .A(n10516), .B(n10469), .Z(n10470) );
  NANDN U16867 ( .A(x[4074]), .B(y[4074]), .Z(n28733) );
  NAND U16868 ( .A(n10470), .B(n28733), .Z(n10472) );
  XNOR U16869 ( .A(x[4075]), .B(n10472), .Z(n10471) );
  NANDN U16870 ( .A(y[4075]), .B(n10471), .Z(n10474) );
  NANDN U16871 ( .A(n10472), .B(x[4075]), .Z(n10473) );
  AND U16872 ( .A(n10474), .B(n10473), .Z(n10475) );
  NANDN U16873 ( .A(n10510), .B(n10475), .Z(n10476) );
  NANDN U16874 ( .A(x[4076]), .B(y[4076]), .Z(n10512) );
  NAND U16875 ( .A(n10476), .B(n10512), .Z(n10478) );
  XNOR U16876 ( .A(x[4077]), .B(n10478), .Z(n10477) );
  NAND U16877 ( .A(n10508), .B(n10477), .Z(n10480) );
  NANDN U16878 ( .A(n10478), .B(x[4077]), .Z(n10479) );
  AND U16879 ( .A(n10480), .B(n10479), .Z(n10481) );
  NANDN U16880 ( .A(n10507), .B(n10481), .Z(n10482) );
  NANDN U16881 ( .A(x[4078]), .B(y[4078]), .Z(n20163) );
  NAND U16882 ( .A(n10482), .B(n20163), .Z(n10484) );
  XNOR U16883 ( .A(x[4079]), .B(n10484), .Z(n10483) );
  NAND U16884 ( .A(n10505), .B(n10483), .Z(n10486) );
  NANDN U16885 ( .A(n10484), .B(x[4079]), .Z(n10485) );
  AND U16886 ( .A(n10486), .B(n10485), .Z(n10487) );
  ANDN U16887 ( .B(x[4080]), .A(y[4080]), .Z(n10504) );
  ANDN U16888 ( .B(n10487), .A(n10504), .Z(n10489) );
  NANDN U16889 ( .A(x[4081]), .B(y[4081]), .Z(n20199) );
  ANDN U16890 ( .B(y[4080]), .A(x[4080]), .Z(n20168) );
  ANDN U16891 ( .B(n20199), .A(n20168), .Z(n10488) );
  NANDN U16892 ( .A(n10489), .B(n10488), .Z(n10490) );
  NANDN U16893 ( .A(n20171), .B(n10490), .Z(n10491) );
  ANDN U16894 ( .B(y[4083]), .A(x[4083]), .Z(n20197) );
  ANDN U16895 ( .B(n10491), .A(n20197), .Z(n10492) );
  ANDN U16896 ( .B(y[4082]), .A(x[4082]), .Z(n20198) );
  ANDN U16897 ( .B(n10492), .A(n20198), .Z(n10494) );
  ANDN U16898 ( .B(x[4083]), .A(y[4083]), .Z(n10502) );
  XOR U16899 ( .A(x[4084]), .B(y[4084]), .Z(n10500) );
  OR U16900 ( .A(n10502), .B(n10500), .Z(n10493) );
  OR U16901 ( .A(n10494), .B(n10493), .Z(n10495) );
  ANDN U16902 ( .B(y[4085]), .A(x[4085]), .Z(n20195) );
  ANDN U16903 ( .B(n10495), .A(n20195), .Z(n10496) );
  NANDN U16904 ( .A(n20196), .B(n10496), .Z(n10497) );
  NAND U16905 ( .A(n10497), .B(n28761), .Z(n10498) );
  AND U16906 ( .A(n10499), .B(n10498), .Z(n20178) );
  NOR U16907 ( .A(n20197), .B(n10500), .Z(n20176) );
  NANDN U16908 ( .A(y[4082]), .B(x[4082]), .Z(n10501) );
  NANDN U16909 ( .A(n10502), .B(n10501), .Z(n28753) );
  NANDN U16910 ( .A(y[4081]), .B(x[4081]), .Z(n10503) );
  NANDN U16911 ( .A(n10504), .B(n10503), .Z(n28749) );
  NAND U16912 ( .A(n10505), .B(x[4079]), .Z(n10506) );
  NANDN U16913 ( .A(n10507), .B(n10506), .Z(n28745) );
  NAND U16914 ( .A(n10508), .B(x[4077]), .Z(n10509) );
  NANDN U16915 ( .A(n10510), .B(n10509), .Z(n28741) );
  NANDN U16916 ( .A(x[4075]), .B(y[4075]), .Z(n10511) );
  NAND U16917 ( .A(n10512), .B(n10511), .Z(n28738) );
  NANDN U16918 ( .A(y[4075]), .B(x[4075]), .Z(n10514) );
  NANDN U16919 ( .A(y[4074]), .B(x[4074]), .Z(n10513) );
  NAND U16920 ( .A(n10514), .B(n10513), .Z(n28736) );
  NOR U16921 ( .A(n28734), .B(n10515), .Z(n20159) );
  OR U16922 ( .A(n10517), .B(n10516), .Z(n28731) );
  NANDN U16923 ( .A(n10519), .B(n10518), .Z(n28729) );
  NANDN U16924 ( .A(n10521), .B(n10520), .Z(n28726) );
  NANDN U16925 ( .A(y[4068]), .B(x[4068]), .Z(n10523) );
  NANDN U16926 ( .A(y[4069]), .B(x[4069]), .Z(n10522) );
  NAND U16927 ( .A(n10523), .B(n10522), .Z(n28723) );
  NAND U16928 ( .A(n10524), .B(y[4068]), .Z(n10526) );
  ANDN U16929 ( .B(n10526), .A(n10525), .Z(n28720) );
  ANDN U16930 ( .B(n28716), .A(n10527), .Z(n20146) );
  NANDN U16931 ( .A(y[4062]), .B(x[4062]), .Z(n10528) );
  NANDN U16932 ( .A(n10529), .B(n10528), .Z(n28709) );
  NAND U16933 ( .A(n10530), .B(y[4062]), .Z(n10532) );
  ANDN U16934 ( .B(n10532), .A(n10531), .Z(n28706) );
  NAND U16935 ( .A(n10533), .B(y[4058]), .Z(n10535) );
  ANDN U16936 ( .B(n10535), .A(n10534), .Z(n28698) );
  NAND U16937 ( .A(n10536), .B(y[4056]), .Z(n10538) );
  ANDN U16938 ( .B(n10538), .A(n10537), .Z(n28694) );
  NANDN U16939 ( .A(y[4052]), .B(x[4052]), .Z(n10539) );
  NANDN U16940 ( .A(n10540), .B(n10539), .Z(n28687) );
  NOR U16941 ( .A(n20200), .B(n10541), .Z(n20115) );
  NOR U16942 ( .A(n10543), .B(n10542), .Z(n28680) );
  NANDN U16943 ( .A(y[4048]), .B(x[4048]), .Z(n10544) );
  NANDN U16944 ( .A(n10545), .B(n10544), .Z(n28679) );
  NAND U16945 ( .A(n10546), .B(y[4046]), .Z(n10548) );
  ANDN U16946 ( .B(n10548), .A(n10547), .Z(n28672) );
  NANDN U16947 ( .A(x[4042]), .B(y[4042]), .Z(n10549) );
  NANDN U16948 ( .A(n10550), .B(n10549), .Z(n28665) );
  AND U16949 ( .A(n10551), .B(n28657), .Z(n20080) );
  NANDN U16950 ( .A(y[4035]), .B(x[4035]), .Z(n10552) );
  NANDN U16951 ( .A(n10553), .B(n10552), .Z(n28647) );
  OR U16952 ( .A(n10555), .B(n10554), .Z(n28637) );
  NANDN U16953 ( .A(y[4028]), .B(x[4028]), .Z(n10557) );
  ANDN U16954 ( .B(n10557), .A(n10556), .Z(n28634) );
  NANDN U16955 ( .A(n10558), .B(n28632), .Z(n20062) );
  OR U16956 ( .A(n10560), .B(n10559), .Z(n28629) );
  NANDN U16957 ( .A(x[4025]), .B(y[4025]), .Z(n10561) );
  NANDN U16958 ( .A(n10562), .B(n10561), .Z(n28627) );
  NANDN U16959 ( .A(y[4024]), .B(x[4024]), .Z(n10563) );
  AND U16960 ( .A(n10564), .B(n10563), .Z(n28624) );
  NAND U16961 ( .A(n10565), .B(n28623), .Z(n20057) );
  NANDN U16962 ( .A(x[4021]), .B(y[4021]), .Z(n10566) );
  NANDN U16963 ( .A(n10567), .B(n10566), .Z(n28617) );
  NAND U16964 ( .A(n10568), .B(x[4019]), .Z(n10570) );
  ANDN U16965 ( .B(n10570), .A(n10569), .Z(n28610) );
  NAND U16966 ( .A(n10571), .B(x[4015]), .Z(n10572) );
  NANDN U16967 ( .A(n10573), .B(n10572), .Z(n28603) );
  NANDN U16968 ( .A(x[4013]), .B(y[4013]), .Z(n10574) );
  NAND U16969 ( .A(n10575), .B(n10574), .Z(n28600) );
  NANDN U16970 ( .A(y[4013]), .B(x[4013]), .Z(n10576) );
  NANDN U16971 ( .A(n10577), .B(n10576), .Z(n28599) );
  NANDN U16972 ( .A(n10579), .B(n10578), .Z(n28594) );
  NANDN U16973 ( .A(x[4010]), .B(y[4010]), .Z(n10581) );
  ANDN U16974 ( .B(n10581), .A(n10580), .Z(n28592) );
  OR U16975 ( .A(n10583), .B(n10582), .Z(n28581) );
  NANDN U16976 ( .A(y[4002]), .B(x[4002]), .Z(n10584) );
  NANDN U16977 ( .A(n10585), .B(n10584), .Z(n28578) );
  NANDN U16978 ( .A(x[4002]), .B(y[4002]), .Z(n10586) );
  NANDN U16979 ( .A(n10587), .B(n10586), .Z(n28577) );
  NAND U16980 ( .A(n10588), .B(y[4000]), .Z(n10589) );
  NANDN U16981 ( .A(n10590), .B(n10589), .Z(n28573) );
  NAND U16982 ( .A(n10591), .B(y[3998]), .Z(n10592) );
  NANDN U16983 ( .A(n10593), .B(n10592), .Z(n28568) );
  NANDN U16984 ( .A(y[3996]), .B(x[3996]), .Z(n10594) );
  NAND U16985 ( .A(n10595), .B(n10594), .Z(n28566) );
  NANDN U16986 ( .A(x[3996]), .B(y[3996]), .Z(n10596) );
  NANDN U16987 ( .A(n10597), .B(n10596), .Z(n28565) );
  NAND U16988 ( .A(n10598), .B(y[3994]), .Z(n10599) );
  NANDN U16989 ( .A(n10600), .B(n10599), .Z(n28561) );
  NANDN U16990 ( .A(x[3992]), .B(y[3992]), .Z(n10602) );
  ANDN U16991 ( .B(n10602), .A(n10601), .Z(n28556) );
  NANDN U16992 ( .A(x[3990]), .B(y[3990]), .Z(n10603) );
  NANDN U16993 ( .A(n10604), .B(n10603), .Z(n28552) );
  OR U16994 ( .A(n10606), .B(n10605), .Z(n28547) );
  OR U16995 ( .A(n10608), .B(n10607), .Z(n28540) );
  NANDN U16996 ( .A(y[3982]), .B(x[3982]), .Z(n10609) );
  NANDN U16997 ( .A(n10610), .B(n10609), .Z(n28539) );
  AND U16998 ( .A(n10611), .B(n28535), .Z(n19982) );
  OR U16999 ( .A(n10613), .B(n10612), .Z(n28533) );
  NANDN U17000 ( .A(y[3979]), .B(x[3979]), .Z(n10615) );
  ANDN U17001 ( .B(n10615), .A(n10614), .Z(n28528) );
  NAND U17002 ( .A(n10616), .B(x[3977]), .Z(n10618) );
  ANDN U17003 ( .B(n10618), .A(n10617), .Z(n28524) );
  NAND U17004 ( .A(n10619), .B(x[3973]), .Z(n10621) );
  NANDN U17005 ( .A(y[3972]), .B(x[3972]), .Z(n10620) );
  AND U17006 ( .A(n10621), .B(n10620), .Z(n28516) );
  OR U17007 ( .A(n10622), .B(n28514), .Z(n19961) );
  OR U17008 ( .A(n10623), .B(n28507), .Z(n19956) );
  NAND U17009 ( .A(n10624), .B(x[3967]), .Z(n10626) );
  ANDN U17010 ( .B(n10626), .A(n10625), .Z(n28500) );
  OR U17011 ( .A(n10628), .B(n10627), .Z(n28493) );
  NANDN U17012 ( .A(n10630), .B(n10629), .Z(n28490) );
  NANDN U17013 ( .A(y[3960]), .B(x[3960]), .Z(n10631) );
  NANDN U17014 ( .A(n10632), .B(n10631), .Z(n28488) );
  NOR U17015 ( .A(n28486), .B(n10633), .Z(n19935) );
  NANDN U17016 ( .A(y[3958]), .B(x[3958]), .Z(n10634) );
  NANDN U17017 ( .A(n10635), .B(n10634), .Z(n28483) );
  OR U17018 ( .A(n10637), .B(n10636), .Z(n28477) );
  NANDN U17019 ( .A(y[3954]), .B(x[3954]), .Z(n10638) );
  NANDN U17020 ( .A(n10639), .B(n10638), .Z(n28472) );
  NANDN U17021 ( .A(y[3952]), .B(x[3952]), .Z(n10640) );
  NANDN U17022 ( .A(n10641), .B(n10640), .Z(n28466) );
  ANDN U17023 ( .B(n28465), .A(n10642), .Z(n19920) );
  XOR U17024 ( .A(x[3950]), .B(n19915), .Z(n10643) );
  AND U17025 ( .A(n28457), .B(n10643), .Z(n19914) );
  OR U17026 ( .A(n10645), .B(n10644), .Z(n28452) );
  NANDN U17027 ( .A(y[3946]), .B(x[3946]), .Z(n10646) );
  NANDN U17028 ( .A(n10647), .B(n10646), .Z(n28451) );
  AND U17029 ( .A(n10648), .B(n28448), .Z(n19907) );
  OR U17030 ( .A(n10650), .B(n10649), .Z(n28445) );
  NAND U17031 ( .A(n10651), .B(x[3943]), .Z(n10652) );
  NANDN U17032 ( .A(n10653), .B(n10652), .Z(n28441) );
  NANDN U17033 ( .A(x[3941]), .B(y[3941]), .Z(n10654) );
  NAND U17034 ( .A(n10655), .B(n10654), .Z(n28438) );
  NANDN U17035 ( .A(y[3941]), .B(x[3941]), .Z(n10656) );
  NANDN U17036 ( .A(n10657), .B(n10656), .Z(n28437) );
  NAND U17037 ( .A(n10658), .B(x[3939]), .Z(n10659) );
  NANDN U17038 ( .A(n10660), .B(n10659), .Z(n28433) );
  NAND U17039 ( .A(n10661), .B(x[3937]), .Z(n10662) );
  NANDN U17040 ( .A(n10663), .B(n10662), .Z(n28428) );
  NANDN U17041 ( .A(n10665), .B(n10664), .Z(n28426) );
  OR U17042 ( .A(n10667), .B(n10666), .Z(n28425) );
  NANDN U17043 ( .A(y[3932]), .B(x[3932]), .Z(n10668) );
  NANDN U17044 ( .A(n10669), .B(n10668), .Z(n28421) );
  NOR U17045 ( .A(n20203), .B(n10670), .Z(n19884) );
  OR U17046 ( .A(n10672), .B(n10671), .Z(n28416) );
  NANDN U17047 ( .A(n10674), .B(n10673), .Z(n28414) );
  NOR U17048 ( .A(n28409), .B(n10675), .Z(n19877) );
  NANDN U17049 ( .A(y[3924]), .B(x[3924]), .Z(n10676) );
  NANDN U17050 ( .A(n10677), .B(n10676), .Z(n28402) );
  NANDN U17051 ( .A(x[3924]), .B(y[3924]), .Z(n10678) );
  NANDN U17052 ( .A(n10679), .B(n10678), .Z(n28400) );
  NOR U17053 ( .A(n20205), .B(n10680), .Z(n19857) );
  OR U17054 ( .A(n10682), .B(n10681), .Z(n28388) );
  NANDN U17055 ( .A(y[3916]), .B(x[3916]), .Z(n10683) );
  NANDN U17056 ( .A(n10684), .B(n10683), .Z(n28387) );
  NOR U17057 ( .A(n20206), .B(n10685), .Z(n19843) );
  OR U17058 ( .A(n10687), .B(n10686), .Z(n28376) );
  NANDN U17059 ( .A(y[3910]), .B(x[3910]), .Z(n10688) );
  NANDN U17060 ( .A(n10689), .B(n10688), .Z(n28375) );
  NAND U17061 ( .A(n10692), .B(x[3908]), .Z(n10691) );
  ANDN U17062 ( .B(n10691), .A(n10690), .Z(n28368) );
  XOR U17063 ( .A(x[3908]), .B(n10692), .Z(n10693) );
  NAND U17064 ( .A(n10693), .B(n20209), .Z(n19832) );
  OR U17065 ( .A(n10695), .B(n10694), .Z(n28362) );
  NANDN U17066 ( .A(y[3904]), .B(x[3904]), .Z(n10697) );
  ANDN U17067 ( .B(n10697), .A(n10696), .Z(n28360) );
  NAND U17068 ( .A(n28357), .B(n10698), .Z(n19825) );
  NANDN U17069 ( .A(x[3901]), .B(y[3901]), .Z(n10699) );
  NANDN U17070 ( .A(n10700), .B(n10699), .Z(n28352) );
  NANDN U17071 ( .A(n10701), .B(n28348), .Z(n19816) );
  NANDN U17072 ( .A(y[3898]), .B(x[3898]), .Z(n10703) );
  ANDN U17073 ( .B(n10703), .A(n10702), .Z(n28344) );
  NOR U17074 ( .A(n28341), .B(n10704), .Z(n19813) );
  NANDN U17075 ( .A(y[3896]), .B(x[3896]), .Z(n10705) );
  NANDN U17076 ( .A(n10706), .B(n10705), .Z(n28339) );
  NAND U17077 ( .A(n10707), .B(x[3894]), .Z(n10708) );
  NANDN U17078 ( .A(n10709), .B(n10708), .Z(n28335) );
  NANDN U17079 ( .A(x[3894]), .B(y[3894]), .Z(n10711) );
  ANDN U17080 ( .B(n10711), .A(n10710), .Z(n28333) );
  OR U17081 ( .A(n10712), .B(n28327), .Z(n19802) );
  NOR U17082 ( .A(n10714), .B(n10713), .Z(n28324) );
  OR U17083 ( .A(n10716), .B(n10715), .Z(n28322) );
  NANDN U17084 ( .A(y[3888]), .B(x[3888]), .Z(n10718) );
  ANDN U17085 ( .B(n10718), .A(n10717), .Z(n28320) );
  NAND U17086 ( .A(n10719), .B(y[3888]), .Z(n10720) );
  NANDN U17087 ( .A(n10721), .B(n10720), .Z(n28318) );
  NANDN U17088 ( .A(y[3886]), .B(x[3886]), .Z(n10722) );
  NAND U17089 ( .A(n10723), .B(n10722), .Z(n28316) );
  NANDN U17090 ( .A(x[3886]), .B(y[3886]), .Z(n10724) );
  NANDN U17091 ( .A(n10725), .B(n10724), .Z(n28315) );
  NAND U17092 ( .A(n10726), .B(y[3884]), .Z(n10727) );
  NANDN U17093 ( .A(n10728), .B(n10727), .Z(n28311) );
  NANDN U17094 ( .A(x[3882]), .B(y[3882]), .Z(n10730) );
  ANDN U17095 ( .B(n10730), .A(n10729), .Z(n28306) );
  NAND U17096 ( .A(n10731), .B(y[3878]), .Z(n10733) );
  ANDN U17097 ( .B(n10733), .A(n10732), .Z(n28298) );
  NAND U17098 ( .A(n10734), .B(y[3876]), .Z(n10736) );
  ANDN U17099 ( .B(n10736), .A(n10735), .Z(n28294) );
  NANDN U17100 ( .A(x[3874]), .B(y[3874]), .Z(n10737) );
  NANDN U17101 ( .A(n10738), .B(n10737), .Z(n28290) );
  NANDN U17102 ( .A(y[3868]), .B(x[3868]), .Z(n10740) );
  ANDN U17103 ( .B(n10740), .A(n10739), .Z(n28280) );
  NAND U17104 ( .A(n10741), .B(y[3868]), .Z(n10742) );
  NANDN U17105 ( .A(n10743), .B(n10742), .Z(n28278) );
  NANDN U17106 ( .A(x[3866]), .B(y[3866]), .Z(n10744) );
  NANDN U17107 ( .A(n10745), .B(n10744), .Z(n28275) );
  NANDN U17108 ( .A(y[3864]), .B(x[3864]), .Z(n10747) );
  ANDN U17109 ( .B(n10747), .A(n10746), .Z(n28272) );
  NAND U17110 ( .A(n10748), .B(y[3864]), .Z(n10749) );
  NANDN U17111 ( .A(n10750), .B(n10749), .Z(n28270) );
  NANDN U17112 ( .A(y[3862]), .B(x[3862]), .Z(n10752) );
  ANDN U17113 ( .B(n10752), .A(n10751), .Z(n28268) );
  OR U17114 ( .A(n10753), .B(n28267), .Z(n19746) );
  OR U17115 ( .A(n10755), .B(n10754), .Z(n28261) );
  NANDN U17116 ( .A(y[3858]), .B(x[3858]), .Z(n10757) );
  ANDN U17117 ( .B(n10757), .A(n10756), .Z(n28258) );
  NAND U17118 ( .A(n10758), .B(y[3858]), .Z(n10759) );
  NANDN U17119 ( .A(n10760), .B(n10759), .Z(n28256) );
  NANDN U17120 ( .A(y[3856]), .B(x[3856]), .Z(n10762) );
  ANDN U17121 ( .B(n10762), .A(n10761), .Z(n28254) );
  NAND U17122 ( .A(n10763), .B(y[3856]), .Z(n10764) );
  NANDN U17123 ( .A(n10765), .B(n10764), .Z(n28253) );
  NANDN U17124 ( .A(x[3854]), .B(y[3854]), .Z(n10766) );
  NANDN U17125 ( .A(n10767), .B(n10766), .Z(n28248) );
  NANDN U17126 ( .A(y[3852]), .B(x[3852]), .Z(n10769) );
  ANDN U17127 ( .B(n10769), .A(n10768), .Z(n28246) );
  NOR U17128 ( .A(n10771), .B(n10770), .Z(n28240) );
  NANDN U17129 ( .A(x[3849]), .B(y[3849]), .Z(n10772) );
  NANDN U17130 ( .A(n10773), .B(n10772), .Z(n28238) );
  NANDN U17131 ( .A(n10775), .B(n10774), .Z(n28236) );
  NANDN U17132 ( .A(x[3847]), .B(y[3847]), .Z(n10776) );
  NANDN U17133 ( .A(n10777), .B(n10776), .Z(n28235) );
  OR U17134 ( .A(n10779), .B(n10778), .Z(n28231) );
  NANDN U17135 ( .A(y[3842]), .B(x[3842]), .Z(n10780) );
  NANDN U17136 ( .A(n10781), .B(n10780), .Z(n28224) );
  NANDN U17137 ( .A(x[3842]), .B(y[3842]), .Z(n10782) );
  NANDN U17138 ( .A(n10783), .B(n10782), .Z(n28222) );
  OR U17139 ( .A(n10785), .B(n10784), .Z(n28213) );
  NANDN U17140 ( .A(y[3832]), .B(x[3832]), .Z(n10786) );
  NANDN U17141 ( .A(n10787), .B(n10786), .Z(n28205) );
  AND U17142 ( .A(n10788), .B(n28202), .Z(n19692) );
  OR U17143 ( .A(n10790), .B(n10789), .Z(n28199) );
  NANDN U17144 ( .A(x[3829]), .B(y[3829]), .Z(n10791) );
  NANDN U17145 ( .A(n10792), .B(n10791), .Z(n28197) );
  NANDN U17146 ( .A(y[3828]), .B(x[3828]), .Z(n10794) );
  NANDN U17147 ( .A(y[3829]), .B(x[3829]), .Z(n10793) );
  NAND U17148 ( .A(n10794), .B(n10793), .Z(n28195) );
  NOR U17149 ( .A(n20212), .B(n10795), .Z(n19687) );
  OR U17150 ( .A(n10797), .B(n10796), .Z(n28191) );
  NANDN U17151 ( .A(n10799), .B(n10798), .Z(n28188) );
  NANDN U17152 ( .A(y[3824]), .B(x[3824]), .Z(n10800) );
  NANDN U17153 ( .A(n10801), .B(n10800), .Z(n28187) );
  NANDN U17154 ( .A(y[3822]), .B(x[3822]), .Z(n10802) );
  NANDN U17155 ( .A(n10803), .B(n10802), .Z(n28181) );
  NOR U17156 ( .A(n28178), .B(n10804), .Z(n19678) );
  NANDN U17157 ( .A(y[3820]), .B(x[3820]), .Z(n10805) );
  NANDN U17158 ( .A(n10806), .B(n10805), .Z(n28175) );
  NANDN U17159 ( .A(y[3816]), .B(x[3816]), .Z(n10808) );
  ANDN U17160 ( .B(n10808), .A(n10807), .Z(n28164) );
  NAND U17161 ( .A(n10809), .B(y[3816]), .Z(n10810) );
  NANDN U17162 ( .A(n10811), .B(n10810), .Z(n28162) );
  NANDN U17163 ( .A(n10812), .B(n28158), .Z(n19661) );
  OR U17164 ( .A(n10814), .B(n10813), .Z(n28153) );
  NAND U17165 ( .A(n10815), .B(y[3807]), .Z(n10816) );
  NANDN U17166 ( .A(n10817), .B(n10816), .Z(n28144) );
  NAND U17167 ( .A(n10818), .B(y[3806]), .Z(n10819) );
  NANDN U17168 ( .A(n10820), .B(n10819), .Z(n28141) );
  NANDN U17169 ( .A(x[3804]), .B(y[3804]), .Z(n10821) );
  NANDN U17170 ( .A(n10822), .B(n10821), .Z(n28137) );
  NANDN U17171 ( .A(y[3802]), .B(x[3802]), .Z(n10824) );
  ANDN U17172 ( .B(n10824), .A(n10823), .Z(n28134) );
  NAND U17173 ( .A(n10825), .B(y[3802]), .Z(n10826) );
  NANDN U17174 ( .A(n10827), .B(n10826), .Z(n28132) );
  NAND U17175 ( .A(n10828), .B(y[3800]), .Z(n10830) );
  ANDN U17176 ( .B(n10830), .A(n10829), .Z(n28128) );
  NANDN U17177 ( .A(x[3798]), .B(y[3798]), .Z(n10831) );
  NANDN U17178 ( .A(n10832), .B(n10831), .Z(n28125) );
  NANDN U17179 ( .A(y[3794]), .B(x[3794]), .Z(n10834) );
  ANDN U17180 ( .B(n10834), .A(n10833), .Z(n28116) );
  OR U17181 ( .A(n10835), .B(n20214), .Z(n19626) );
  NANDN U17182 ( .A(n10837), .B(n10836), .Z(n28113) );
  OR U17183 ( .A(n10839), .B(n10838), .Z(n28111) );
  NAND U17184 ( .A(n10840), .B(y[3790]), .Z(n10841) );
  NANDN U17185 ( .A(n10842), .B(n10841), .Z(n28107) );
  NANDN U17186 ( .A(x[3788]), .B(y[3788]), .Z(n10844) );
  ANDN U17187 ( .B(n10844), .A(n10843), .Z(n28102) );
  NANDN U17188 ( .A(x[3786]), .B(y[3786]), .Z(n10845) );
  NANDN U17189 ( .A(n10846), .B(n10845), .Z(n28099) );
  NAND U17190 ( .A(n10847), .B(y[3782]), .Z(n10849) );
  ANDN U17191 ( .B(n10849), .A(n10848), .Z(n28090) );
  NANDN U17192 ( .A(x[3780]), .B(y[3780]), .Z(n10850) );
  NANDN U17193 ( .A(n10851), .B(n10850), .Z(n28087) );
  NOR U17194 ( .A(n28083), .B(n10852), .Z(n19592) );
  NANDN U17195 ( .A(y[3774]), .B(x[3774]), .Z(n10853) );
  NANDN U17196 ( .A(n10854), .B(n10853), .Z(n28075) );
  NANDN U17197 ( .A(x[3774]), .B(y[3774]), .Z(n10855) );
  NANDN U17198 ( .A(n10856), .B(n10855), .Z(n28072) );
  ANDN U17199 ( .B(n28068), .A(n10857), .Z(n19579) );
  NOR U17200 ( .A(n10859), .B(n10858), .Z(n28062) );
  OR U17201 ( .A(n10861), .B(n10860), .Z(n28060) );
  NANDN U17202 ( .A(y[3764]), .B(x[3764]), .Z(n10862) );
  NANDN U17203 ( .A(n10863), .B(n10862), .Z(n28053) );
  AND U17204 ( .A(n10864), .B(n20217), .Z(n19562) );
  OR U17205 ( .A(n10866), .B(n10865), .Z(n28049) );
  NANDN U17206 ( .A(y[3761]), .B(x[3761]), .Z(n10867) );
  NANDN U17207 ( .A(n10868), .B(n10867), .Z(n28045) );
  NANDN U17208 ( .A(x[3759]), .B(y[3759]), .Z(n10870) );
  ANDN U17209 ( .B(n10870), .A(n10869), .Z(n28042) );
  NAND U17210 ( .A(n10871), .B(x[3759]), .Z(n10872) );
  NANDN U17211 ( .A(n10873), .B(n10872), .Z(n28040) );
  NAND U17212 ( .A(n10874), .B(x[3757]), .Z(n10876) );
  ANDN U17213 ( .B(n10876), .A(n10875), .Z(n28036) );
  NAND U17214 ( .A(n10877), .B(x[3753]), .Z(n10879) );
  ANDN U17215 ( .B(n10879), .A(n10878), .Z(n28028) );
  NANDN U17216 ( .A(n10880), .B(n28017), .Z(n19527) );
  NANDN U17217 ( .A(y[3746]), .B(x[3746]), .Z(n10882) );
  ANDN U17218 ( .B(n10882), .A(n10881), .Z(n28014) );
  OR U17219 ( .A(n10884), .B(n10883), .Z(n28009) );
  NANDN U17220 ( .A(x[3742]), .B(y[3742]), .Z(n10885) );
  NANDN U17221 ( .A(n10886), .B(n10885), .Z(n28005) );
  NANDN U17222 ( .A(y[3740]), .B(x[3740]), .Z(n10888) );
  ANDN U17223 ( .B(n10888), .A(n10887), .Z(n28002) );
  OR U17224 ( .A(n10890), .B(n10889), .Z(n27997) );
  NANDN U17225 ( .A(y[3736]), .B(x[3736]), .Z(n10891) );
  NANDN U17226 ( .A(n10892), .B(n10891), .Z(n27995) );
  NANDN U17227 ( .A(x[3736]), .B(y[3736]), .Z(n10893) );
  NANDN U17228 ( .A(n10894), .B(n10893), .Z(n27993) );
  NAND U17229 ( .A(n10895), .B(y[3734]), .Z(n10896) );
  NANDN U17230 ( .A(n10897), .B(n10896), .Z(n27989) );
  NANDN U17231 ( .A(y[3732]), .B(x[3732]), .Z(n10899) );
  ANDN U17232 ( .B(n10899), .A(n10898), .Z(n27986) );
  NAND U17233 ( .A(n10900), .B(y[3732]), .Z(n10901) );
  NANDN U17234 ( .A(n10902), .B(n10901), .Z(n27985) );
  NANDN U17235 ( .A(x[3730]), .B(y[3730]), .Z(n10903) );
  NANDN U17236 ( .A(n10904), .B(n10903), .Z(n27980) );
  NANDN U17237 ( .A(y[3728]), .B(x[3728]), .Z(n10906) );
  ANDN U17238 ( .B(n10906), .A(n10905), .Z(n27978) );
  OR U17239 ( .A(n10907), .B(n27977), .Z(n19492) );
  NOR U17240 ( .A(n27971), .B(n10908), .Z(n19487) );
  NANDN U17241 ( .A(y[3722]), .B(x[3722]), .Z(n10909) );
  NANDN U17242 ( .A(n10910), .B(n10909), .Z(n27963) );
  NANDN U17243 ( .A(x[3722]), .B(y[3722]), .Z(n10911) );
  NANDN U17244 ( .A(n10912), .B(n10911), .Z(n27960) );
  NOR U17245 ( .A(n27954), .B(n10913), .Z(n19474) );
  NOR U17246 ( .A(n10915), .B(n10914), .Z(n27950) );
  NANDN U17247 ( .A(y[3716]), .B(x[3716]), .Z(n10916) );
  NANDN U17248 ( .A(n10917), .B(n10916), .Z(n27949) );
  NANDN U17249 ( .A(x[3716]), .B(y[3716]), .Z(n10918) );
  NANDN U17250 ( .A(n10919), .B(n10918), .Z(n27947) );
  NOR U17251 ( .A(n27937), .B(n10920), .Z(n19456) );
  NANDN U17252 ( .A(y[3708]), .B(x[3708]), .Z(n10921) );
  NANDN U17253 ( .A(n10922), .B(n10921), .Z(n27931) );
  NOR U17254 ( .A(n10924), .B(n10923), .Z(n27908) );
  OR U17255 ( .A(n10926), .B(n10925), .Z(n27907) );
  NANDN U17256 ( .A(x[3696]), .B(y[3696]), .Z(n10927) );
  NANDN U17257 ( .A(n10928), .B(n10927), .Z(n27902) );
  NANDN U17258 ( .A(x[3694]), .B(y[3694]), .Z(n10929) );
  NANDN U17259 ( .A(n10930), .B(n10929), .Z(n27899) );
  NANDN U17260 ( .A(y[3692]), .B(x[3692]), .Z(n10931) );
  NAND U17261 ( .A(n10932), .B(n10931), .Z(n27897) );
  NANDN U17262 ( .A(x[3692]), .B(y[3692]), .Z(n10933) );
  NANDN U17263 ( .A(n10934), .B(n10933), .Z(n27895) );
  NAND U17264 ( .A(n10935), .B(y[3690]), .Z(n10936) );
  NANDN U17265 ( .A(n10937), .B(n10936), .Z(n27891) );
  NANDN U17266 ( .A(x[3688]), .B(y[3688]), .Z(n10938) );
  NANDN U17267 ( .A(n10939), .B(n10938), .Z(n27887) );
  NANDN U17268 ( .A(x[3684]), .B(y[3684]), .Z(n10940) );
  NANDN U17269 ( .A(n10941), .B(n10940), .Z(n27879) );
  NANDN U17270 ( .A(y[3682]), .B(x[3682]), .Z(n10942) );
  NAND U17271 ( .A(n10943), .B(n10942), .Z(n27877) );
  NANDN U17272 ( .A(x[3682]), .B(y[3682]), .Z(n10944) );
  NANDN U17273 ( .A(n10945), .B(n10944), .Z(n27875) );
  NAND U17274 ( .A(n10946), .B(y[3680]), .Z(n10947) );
  NANDN U17275 ( .A(n10948), .B(n10947), .Z(n27871) );
  NANDN U17276 ( .A(x[3678]), .B(y[3678]), .Z(n10949) );
  NANDN U17277 ( .A(n10950), .B(n10949), .Z(n27867) );
  NANDN U17278 ( .A(x[3674]), .B(y[3674]), .Z(n10951) );
  NANDN U17279 ( .A(n10952), .B(n10951), .Z(n27859) );
  NANDN U17280 ( .A(y[3672]), .B(x[3672]), .Z(n10953) );
  NAND U17281 ( .A(n10954), .B(n10953), .Z(n27857) );
  NANDN U17282 ( .A(x[3672]), .B(y[3672]), .Z(n10955) );
  NANDN U17283 ( .A(n10956), .B(n10955), .Z(n27855) );
  NAND U17284 ( .A(n10957), .B(y[3670]), .Z(n10958) );
  NANDN U17285 ( .A(n10959), .B(n10958), .Z(n27851) );
  OR U17286 ( .A(n10961), .B(n10960), .Z(n27847) );
  OR U17287 ( .A(n10963), .B(n10962), .Z(n27845) );
  NANDN U17288 ( .A(y[3664]), .B(x[3664]), .Z(n10964) );
  NAND U17289 ( .A(n10965), .B(n10964), .Z(n27841) );
  OR U17290 ( .A(n10967), .B(n10966), .Z(n27835) );
  OR U17291 ( .A(n10969), .B(n10968), .Z(n27833) );
  OR U17292 ( .A(n10971), .B(n10970), .Z(n27829) );
  NANDN U17293 ( .A(y[3658]), .B(x[3658]), .Z(n10972) );
  NANDN U17294 ( .A(n10973), .B(n10972), .Z(n27827) );
  OR U17295 ( .A(n10975), .B(n10974), .Z(n27821) );
  NANDN U17296 ( .A(y[3652]), .B(x[3652]), .Z(n10977) );
  ANDN U17297 ( .B(n10977), .A(n10976), .Z(n27810) );
  NOR U17298 ( .A(n10979), .B(n10978), .Z(n27804) );
  OR U17299 ( .A(n10981), .B(n10980), .Z(n27802) );
  OR U17300 ( .A(n10983), .B(n10982), .Z(n27801) );
  NANDN U17301 ( .A(y[3644]), .B(x[3644]), .Z(n10984) );
  NANDN U17302 ( .A(n10985), .B(n10984), .Z(n27793) );
  NOR U17303 ( .A(n10987), .B(n10986), .Z(n27786) );
  NANDN U17304 ( .A(x[3641]), .B(y[3641]), .Z(n10988) );
  NANDN U17305 ( .A(n10989), .B(n10988), .Z(n27784) );
  NANDN U17306 ( .A(y[3641]), .B(x[3641]), .Z(n10990) );
  NANDN U17307 ( .A(n10991), .B(n10990), .Z(n27783) );
  NANDN U17308 ( .A(y[3639]), .B(x[3639]), .Z(n10992) );
  NANDN U17309 ( .A(n10993), .B(n10992), .Z(n27779) );
  NANDN U17310 ( .A(x[3637]), .B(y[3637]), .Z(n10995) );
  ANDN U17311 ( .B(n10995), .A(n10994), .Z(n27776) );
  NAND U17312 ( .A(n10996), .B(x[3637]), .Z(n10997) );
  NANDN U17313 ( .A(n10998), .B(n10997), .Z(n27774) );
  NANDN U17314 ( .A(y[3632]), .B(x[3632]), .Z(n11000) );
  ANDN U17315 ( .B(n11000), .A(n10999), .Z(n27766) );
  OR U17316 ( .A(n11001), .B(n27755), .Z(n19277) );
  NOR U17317 ( .A(n11003), .B(n11002), .Z(n27752) );
  OR U17318 ( .A(n11005), .B(n11004), .Z(n27750) );
  OR U17319 ( .A(n11007), .B(n11006), .Z(n27749) );
  NANDN U17320 ( .A(y[3620]), .B(x[3620]), .Z(n11008) );
  NANDN U17321 ( .A(n11009), .B(n11008), .Z(n27741) );
  NANDN U17322 ( .A(x[3617]), .B(y[3617]), .Z(n11010) );
  NANDN U17323 ( .A(n11011), .B(n11010), .Z(n27732) );
  NAND U17324 ( .A(n11012), .B(x[3617]), .Z(n11014) );
  ANDN U17325 ( .B(n11014), .A(n11013), .Z(n27730) );
  NANDN U17326 ( .A(y[3615]), .B(x[3615]), .Z(n11015) );
  NANDN U17327 ( .A(n11016), .B(n11015), .Z(n27727) );
  NANDN U17328 ( .A(y[3613]), .B(x[3613]), .Z(n11017) );
  NANDN U17329 ( .A(n11018), .B(n11017), .Z(n27722) );
  NANDN U17330 ( .A(x[3611]), .B(y[3611]), .Z(n11020) );
  ANDN U17331 ( .B(n11020), .A(n11019), .Z(n27720) );
  NAND U17332 ( .A(n11021), .B(x[3611]), .Z(n11022) );
  NANDN U17333 ( .A(n11023), .B(n11022), .Z(n27719) );
  NANDN U17334 ( .A(y[3606]), .B(x[3606]), .Z(n11025) );
  ANDN U17335 ( .B(n11025), .A(n11024), .Z(n27710) );
  NOR U17336 ( .A(n27701), .B(n11026), .Z(n19228) );
  OR U17337 ( .A(n11028), .B(n11027), .Z(n27699) );
  NANDN U17338 ( .A(n11030), .B(n11029), .Z(n27696) );
  NANDN U17339 ( .A(y[3598]), .B(x[3598]), .Z(n11032) );
  ANDN U17340 ( .B(n11032), .A(n11031), .Z(n27688) );
  NOR U17341 ( .A(n27687), .B(n11033), .Z(n19217) );
  OR U17342 ( .A(n11035), .B(n11034), .Z(n27681) );
  NANDN U17343 ( .A(y[3594]), .B(x[3594]), .Z(n11036) );
  NANDN U17344 ( .A(n11037), .B(n11036), .Z(n27679) );
  NANDN U17345 ( .A(x[3592]), .B(y[3592]), .Z(n11038) );
  NANDN U17346 ( .A(n11039), .B(n11038), .Z(n27673) );
  NANDN U17347 ( .A(y[3590]), .B(x[3590]), .Z(n11040) );
  NAND U17348 ( .A(n11041), .B(n11040), .Z(n27671) );
  NANDN U17349 ( .A(x[3590]), .B(y[3590]), .Z(n11042) );
  NANDN U17350 ( .A(n11043), .B(n11042), .Z(n27669) );
  NANDN U17351 ( .A(y[3588]), .B(x[3588]), .Z(n11045) );
  ANDN U17352 ( .B(n11045), .A(n11044), .Z(n27666) );
  NOR U17353 ( .A(n27662), .B(n11046), .Z(n19199) );
  OR U17354 ( .A(n11048), .B(n11047), .Z(n27658) );
  NANDN U17355 ( .A(y[3584]), .B(x[3584]), .Z(n11049) );
  NANDN U17356 ( .A(n11050), .B(n11049), .Z(n27657) );
  NOR U17357 ( .A(n27653), .B(n11051), .Z(n19192) );
  NANDN U17358 ( .A(n11053), .B(n11052), .Z(n27650) );
  OR U17359 ( .A(n11055), .B(n11054), .Z(n27649) );
  NANDN U17360 ( .A(x[3580]), .B(y[3580]), .Z(n11056) );
  NANDN U17361 ( .A(n11057), .B(n11056), .Z(n27645) );
  ANDN U17362 ( .B(n11059), .A(n11058), .Z(n27642) );
  OR U17363 ( .A(n11061), .B(n11060), .Z(n27640) );
  OR U17364 ( .A(n11063), .B(n11062), .Z(n27639) );
  NANDN U17365 ( .A(y[3572]), .B(x[3572]), .Z(n11064) );
  NANDN U17366 ( .A(n11065), .B(n11064), .Z(n27631) );
  AND U17367 ( .A(n11066), .B(n27628), .Z(n19171) );
  OR U17368 ( .A(n11068), .B(n11067), .Z(n27625) );
  NANDN U17369 ( .A(x[3569]), .B(y[3569]), .Z(n11069) );
  NANDN U17370 ( .A(n11070), .B(n11069), .Z(n27623) );
  NANDN U17371 ( .A(y[3569]), .B(x[3569]), .Z(n11071) );
  NANDN U17372 ( .A(n11072), .B(n11071), .Z(n27621) );
  NAND U17373 ( .A(n11073), .B(x[3567]), .Z(n11074) );
  NANDN U17374 ( .A(n11075), .B(n11074), .Z(n27617) );
  OR U17375 ( .A(n11077), .B(n11076), .Z(n27613) );
  NANDN U17376 ( .A(y[3562]), .B(x[3562]), .Z(n11079) );
  ANDN U17377 ( .B(n11079), .A(n11078), .Z(n27608) );
  NANDN U17378 ( .A(n11081), .B(n11080), .Z(n27598) );
  OR U17379 ( .A(n11083), .B(n11082), .Z(n27597) );
  NANDN U17380 ( .A(y[3556]), .B(x[3556]), .Z(n11085) );
  ANDN U17381 ( .B(n11085), .A(n11084), .Z(n27594) );
  NAND U17382 ( .A(n11086), .B(y[3556]), .Z(n11087) );
  NANDN U17383 ( .A(n11088), .B(n11087), .Z(n27593) );
  NANDN U17384 ( .A(x[3554]), .B(y[3554]), .Z(n11089) );
  NANDN U17385 ( .A(n11090), .B(n11089), .Z(n27588) );
  NAND U17386 ( .A(n11091), .B(y[3552]), .Z(n11093) );
  ANDN U17387 ( .B(n11093), .A(n11092), .Z(n27584) );
  NANDN U17388 ( .A(x[3550]), .B(y[3550]), .Z(n11094) );
  NANDN U17389 ( .A(n11095), .B(n11094), .Z(n27581) );
  NANDN U17390 ( .A(y[3548]), .B(x[3548]), .Z(n11096) );
  NAND U17391 ( .A(n11097), .B(n11096), .Z(n27578) );
  NANDN U17392 ( .A(x[3548]), .B(y[3548]), .Z(n11098) );
  NANDN U17393 ( .A(n11099), .B(n11098), .Z(n27577) );
  NANDN U17394 ( .A(y[3546]), .B(x[3546]), .Z(n11101) );
  ANDN U17395 ( .B(n11101), .A(n11100), .Z(n27574) );
  NAND U17396 ( .A(n11102), .B(y[3546]), .Z(n11103) );
  NANDN U17397 ( .A(n11104), .B(n11103), .Z(n27573) );
  NANDN U17398 ( .A(x[3544]), .B(y[3544]), .Z(n11105) );
  NANDN U17399 ( .A(n11106), .B(n11105), .Z(n27568) );
  XOR U17400 ( .A(n11107), .B(y[3542]), .Z(n19118) );
  NANDN U17401 ( .A(n11109), .B(n11108), .Z(n27561) );
  OR U17402 ( .A(n11111), .B(n11110), .Z(n27559) );
  NAND U17403 ( .A(n11112), .B(y[3538]), .Z(n11113) );
  NANDN U17404 ( .A(n11114), .B(n11113), .Z(n27555) );
  NANDN U17405 ( .A(x[3536]), .B(y[3536]), .Z(n11115) );
  NANDN U17406 ( .A(n11116), .B(n11115), .Z(n27551) );
  OR U17407 ( .A(n11118), .B(n11117), .Z(n27537) );
  NANDN U17408 ( .A(y[3528]), .B(x[3528]), .Z(n11119) );
  NANDN U17409 ( .A(n11120), .B(n11119), .Z(n27535) );
  NANDN U17410 ( .A(x[3528]), .B(y[3528]), .Z(n11121) );
  NANDN U17411 ( .A(n11122), .B(n11121), .Z(n27533) );
  OR U17412 ( .A(n11124), .B(n11123), .Z(n27519) );
  NANDN U17413 ( .A(y[3520]), .B(x[3520]), .Z(n11125) );
  NANDN U17414 ( .A(n11126), .B(n11125), .Z(n27517) );
  NANDN U17415 ( .A(x[3520]), .B(y[3520]), .Z(n11127) );
  NANDN U17416 ( .A(n11128), .B(n11127), .Z(n27515) );
  NANDN U17417 ( .A(x[3516]), .B(y[3516]), .Z(n11129) );
  NANDN U17418 ( .A(n11130), .B(n11129), .Z(n27507) );
  NANDN U17419 ( .A(y[3514]), .B(x[3514]), .Z(n11131) );
  NAND U17420 ( .A(n11132), .B(n11131), .Z(n27505) );
  NANDN U17421 ( .A(x[3514]), .B(y[3514]), .Z(n11133) );
  NANDN U17422 ( .A(n11134), .B(n11133), .Z(n27503) );
  NAND U17423 ( .A(n11135), .B(y[3512]), .Z(n11136) );
  NANDN U17424 ( .A(n11137), .B(n11136), .Z(n27499) );
  NANDN U17425 ( .A(x[3510]), .B(y[3510]), .Z(n11138) );
  NANDN U17426 ( .A(n11139), .B(n11138), .Z(n27495) );
  OR U17427 ( .A(n11141), .B(n11140), .Z(n27489) );
  NAND U17428 ( .A(n11143), .B(n11142), .Z(n27485) );
  OR U17429 ( .A(n11145), .B(n11144), .Z(n27483) );
  NANDN U17430 ( .A(y[3502]), .B(x[3502]), .Z(n11147) );
  ANDN U17431 ( .B(n11147), .A(n11146), .Z(n27480) );
  AND U17432 ( .A(n11148), .B(n27478), .Z(n19033) );
  OR U17433 ( .A(n11150), .B(n11149), .Z(n27475) );
  NANDN U17434 ( .A(x[3499]), .B(y[3499]), .Z(n11151) );
  NANDN U17435 ( .A(n11152), .B(n11151), .Z(n27473) );
  NANDN U17436 ( .A(y[3499]), .B(x[3499]), .Z(n11153) );
  NANDN U17437 ( .A(n11154), .B(n11153), .Z(n27471) );
  NAND U17438 ( .A(n11155), .B(x[3497]), .Z(n11156) );
  NANDN U17439 ( .A(n11157), .B(n11156), .Z(n27467) );
  NANDN U17440 ( .A(y[3495]), .B(x[3495]), .Z(n11158) );
  NANDN U17441 ( .A(n11159), .B(n11158), .Z(n27463) );
  OR U17442 ( .A(n11161), .B(n11160), .Z(n27449) );
  NANDN U17443 ( .A(y[3486]), .B(x[3486]), .Z(n11162) );
  NANDN U17444 ( .A(n11163), .B(n11162), .Z(n27447) );
  NANDN U17445 ( .A(x[3486]), .B(y[3486]), .Z(n11164) );
  NANDN U17446 ( .A(n11165), .B(n11164), .Z(n27445) );
  NAND U17447 ( .A(n11166), .B(y[3484]), .Z(n11167) );
  NANDN U17448 ( .A(n11168), .B(n11167), .Z(n27441) );
  NANDN U17449 ( .A(x[3482]), .B(y[3482]), .Z(n11169) );
  NANDN U17450 ( .A(n11170), .B(n11169), .Z(n27437) );
  NANDN U17451 ( .A(x[3476]), .B(y[3476]), .Z(n11171) );
  NANDN U17452 ( .A(n11172), .B(n11171), .Z(n27423) );
  OR U17453 ( .A(n11174), .B(n11173), .Z(n27421) );
  NANDN U17454 ( .A(x[3473]), .B(y[3473]), .Z(n11175) );
  NAND U17455 ( .A(n11176), .B(n11175), .Z(n27419) );
  NANDN U17456 ( .A(n11178), .B(n11177), .Z(n27417) );
  NANDN U17457 ( .A(y[3470]), .B(x[3470]), .Z(n11180) );
  NAND U17458 ( .A(n11180), .B(n11179), .Z(n27413) );
  NAND U17459 ( .A(n11182), .B(n11181), .Z(n27405) );
  NANDN U17460 ( .A(y[3467]), .B(x[3467]), .Z(n11183) );
  NANDN U17461 ( .A(n11184), .B(n11183), .Z(n27402) );
  NANDN U17462 ( .A(y[3463]), .B(x[3463]), .Z(n11185) );
  NANDN U17463 ( .A(n11186), .B(n11185), .Z(n27395) );
  OR U17464 ( .A(n11188), .B(n11187), .Z(n27392) );
  NAND U17465 ( .A(n11190), .B(n11189), .Z(n27389) );
  OR U17466 ( .A(n11192), .B(n11191), .Z(n27385) );
  NANDN U17467 ( .A(y[3455]), .B(x[3455]), .Z(n11193) );
  NANDN U17468 ( .A(n11194), .B(n11193), .Z(n27379) );
  NAND U17469 ( .A(n11196), .B(n11195), .Z(n27372) );
  OR U17470 ( .A(n11198), .B(n11197), .Z(n27369) );
  NAND U17471 ( .A(n11200), .B(n11199), .Z(n27365) );
  NANDN U17472 ( .A(y[3447]), .B(x[3447]), .Z(n11201) );
  NANDN U17473 ( .A(n11202), .B(n11201), .Z(n27362) );
  NANDN U17474 ( .A(y[3443]), .B(x[3443]), .Z(n11203) );
  NANDN U17475 ( .A(n11204), .B(n11203), .Z(n27355) );
  OR U17476 ( .A(n11206), .B(n11205), .Z(n27352) );
  NAND U17477 ( .A(n11208), .B(n11207), .Z(n27349) );
  OR U17478 ( .A(n11210), .B(n11209), .Z(n27345) );
  NANDN U17479 ( .A(y[3434]), .B(x[3434]), .Z(n11211) );
  NANDN U17480 ( .A(n11212), .B(n11211), .Z(n27339) );
  NAND U17481 ( .A(n11213), .B(x[3433]), .Z(n11215) );
  NANDN U17482 ( .A(y[3432]), .B(x[3432]), .Z(n11214) );
  NAND U17483 ( .A(n11215), .B(n11214), .Z(n27335) );
  NANDN U17484 ( .A(x[3429]), .B(y[3429]), .Z(n11216) );
  NANDN U17485 ( .A(n11217), .B(n11216), .Z(n27329) );
  NANDN U17486 ( .A(y[3428]), .B(x[3428]), .Z(n11218) );
  NAND U17487 ( .A(n11219), .B(n11218), .Z(n27327) );
  NANDN U17488 ( .A(y[3427]), .B(x[3427]), .Z(n11221) );
  NANDN U17489 ( .A(y[3426]), .B(x[3426]), .Z(n11220) );
  NAND U17490 ( .A(n11221), .B(n11220), .Z(n27322) );
  NAND U17491 ( .A(n11222), .B(y[3426]), .Z(n11224) );
  ANDN U17492 ( .B(n11224), .A(n11223), .Z(n27320) );
  NAND U17493 ( .A(n11226), .B(n11225), .Z(n27317) );
  NANDN U17494 ( .A(x[3422]), .B(y[3422]), .Z(n11228) );
  NAND U17495 ( .A(n11228), .B(n11227), .Z(n27312) );
  NANDN U17496 ( .A(y[3421]), .B(x[3421]), .Z(n11230) );
  NANDN U17497 ( .A(y[3420]), .B(x[3420]), .Z(n11229) );
  AND U17498 ( .A(n11230), .B(n11229), .Z(n27310) );
  NAND U17499 ( .A(n11231), .B(y[3420]), .Z(n11232) );
  NANDN U17500 ( .A(n11233), .B(n11232), .Z(n27309) );
  NANDN U17501 ( .A(y[3417]), .B(x[3417]), .Z(n11235) );
  NANDN U17502 ( .A(y[3416]), .B(x[3416]), .Z(n11234) );
  NAND U17503 ( .A(n11235), .B(n11234), .Z(n27302) );
  NAND U17504 ( .A(n11236), .B(y[3416]), .Z(n11238) );
  ANDN U17505 ( .B(n11238), .A(n11237), .Z(n27300) );
  NANDN U17506 ( .A(x[3413]), .B(y[3413]), .Z(n11239) );
  NAND U17507 ( .A(n11240), .B(n11239), .Z(n27297) );
  NANDN U17508 ( .A(y[3410]), .B(x[3410]), .Z(n11241) );
  AND U17509 ( .A(n11242), .B(n11241), .Z(n27290) );
  XOR U17510 ( .A(n11243), .B(y[3410]), .Z(n11244) );
  AND U17511 ( .A(n27288), .B(n11244), .Z(n18853) );
  OR U17512 ( .A(n11246), .B(n11245), .Z(n27285) );
  NAND U17513 ( .A(n11248), .B(n11247), .Z(n27280) );
  NANDN U17514 ( .A(x[3406]), .B(y[3406]), .Z(n11250) );
  ANDN U17515 ( .B(n11250), .A(n11249), .Z(n27278) );
  OR U17516 ( .A(n11252), .B(n11251), .Z(n27277) );
  NANDN U17517 ( .A(x[3402]), .B(y[3402]), .Z(n11253) );
  NANDN U17518 ( .A(n11254), .B(n11253), .Z(n27270) );
  NOR U17519 ( .A(n11256), .B(n11255), .Z(n27268) );
  NAND U17520 ( .A(n11258), .B(n11257), .Z(n27265) );
  OR U17521 ( .A(n11260), .B(n11259), .Z(n27260) );
  NANDN U17522 ( .A(x[3395]), .B(y[3395]), .Z(n11262) );
  ANDN U17523 ( .B(n11262), .A(n11261), .Z(n27258) );
  NAND U17524 ( .A(n11264), .B(n11263), .Z(n27257) );
  NANDN U17525 ( .A(x[3394]), .B(y[3394]), .Z(n11265) );
  NANDN U17526 ( .A(n11266), .B(n11265), .Z(n27255) );
  NANDN U17527 ( .A(y[3390]), .B(x[3390]), .Z(n11267) );
  AND U17528 ( .A(n11268), .B(n11267), .Z(n27248) );
  XNOR U17529 ( .A(y[3390]), .B(x[3390]), .Z(n18817) );
  NOR U17530 ( .A(n11270), .B(n11269), .Z(n27240) );
  NANDN U17531 ( .A(n11272), .B(n11271), .Z(n27237) );
  NAND U17532 ( .A(n11273), .B(y[3384]), .Z(n11274) );
  NANDN U17533 ( .A(n11275), .B(n11274), .Z(n27232) );
  NANDN U17534 ( .A(n11277), .B(n11276), .Z(n27228) );
  NAND U17535 ( .A(n11278), .B(y[3377]), .Z(n11279) );
  NANDN U17536 ( .A(n11280), .B(n11279), .Z(n27220) );
  NANDN U17537 ( .A(y[3377]), .B(x[3377]), .Z(n11282) );
  AND U17538 ( .A(n11282), .B(n11281), .Z(n27218) );
  NANDN U17539 ( .A(x[3376]), .B(y[3376]), .Z(n11283) );
  NANDN U17540 ( .A(n11284), .B(n11283), .Z(n27217) );
  OR U17541 ( .A(n11286), .B(n11285), .Z(n27215) );
  NAND U17542 ( .A(n11288), .B(n11287), .Z(n27210) );
  NANDN U17543 ( .A(x[3372]), .B(y[3372]), .Z(n11290) );
  ANDN U17544 ( .B(n11290), .A(n11289), .Z(n27208) );
  OR U17545 ( .A(n11292), .B(n11291), .Z(n27207) );
  NANDN U17546 ( .A(x[3367]), .B(y[3367]), .Z(n11293) );
  NANDN U17547 ( .A(n11294), .B(n11293), .Z(n27200) );
  NANDN U17548 ( .A(y[3366]), .B(x[3366]), .Z(n11295) );
  AND U17549 ( .A(n11296), .B(n11295), .Z(n27198) );
  NOR U17550 ( .A(n11298), .B(n11297), .Z(n27190) );
  NANDN U17551 ( .A(y[3362]), .B(x[3362]), .Z(n11299) );
  NANDN U17552 ( .A(n11300), .B(n11299), .Z(n27189) );
  NANDN U17553 ( .A(n11302), .B(n11301), .Z(n27187) );
  NANDN U17554 ( .A(y[3359]), .B(x[3359]), .Z(n11304) );
  NANDN U17555 ( .A(y[3358]), .B(x[3358]), .Z(n11303) );
  AND U17556 ( .A(n11304), .B(n11303), .Z(n27180) );
  NAND U17557 ( .A(n11306), .B(n11305), .Z(n27167) );
  OR U17558 ( .A(n11308), .B(n11307), .Z(n27162) );
  NANDN U17559 ( .A(y[3350]), .B(x[3350]), .Z(n11310) );
  ANDN U17560 ( .B(n11310), .A(n11309), .Z(n27160) );
  NAND U17561 ( .A(n11312), .B(n11311), .Z(n27159) );
  NANDN U17562 ( .A(y[3349]), .B(x[3349]), .Z(n11313) );
  NANDN U17563 ( .A(n11314), .B(n11313), .Z(n27157) );
  AND U17564 ( .A(n11316), .B(n11315), .Z(n27150) );
  NANDN U17565 ( .A(y[3345]), .B(x[3345]), .Z(n11317) );
  NANDN U17566 ( .A(n11318), .B(n11317), .Z(n27149) );
  OR U17567 ( .A(n11320), .B(n11319), .Z(n27147) );
  NANDN U17568 ( .A(y[3340]), .B(x[3340]), .Z(n11322) );
  ANDN U17569 ( .B(n11322), .A(n11321), .Z(n27140) );
  OR U17570 ( .A(n11324), .B(n11323), .Z(n27135) );
  NANDN U17571 ( .A(n11326), .B(n11325), .Z(n27133) );
  NANDN U17572 ( .A(y[3337]), .B(x[3337]), .Z(n11327) );
  NANDN U17573 ( .A(n11328), .B(n11327), .Z(n27130) );
  NANDN U17574 ( .A(x[3331]), .B(y[3331]), .Z(n11330) );
  NAND U17575 ( .A(n11330), .B(n11329), .Z(n27121) );
  AND U17576 ( .A(n11332), .B(n11331), .Z(n27118) );
  NANDN U17577 ( .A(x[3330]), .B(y[3330]), .Z(n11333) );
  NANDN U17578 ( .A(n11334), .B(n11333), .Z(n27117) );
  NANDN U17579 ( .A(y[3326]), .B(x[3326]), .Z(n11335) );
  AND U17580 ( .A(n11336), .B(n11335), .Z(n27110) );
  AND U17581 ( .A(n11337), .B(n27107), .Z(n18705) );
  OR U17582 ( .A(n11339), .B(n11338), .Z(n27104) );
  NANDN U17583 ( .A(y[3320]), .B(x[3320]), .Z(n11340) );
  NANDN U17584 ( .A(n11341), .B(n11340), .Z(n27097) );
  AND U17585 ( .A(n20229), .B(n11342), .Z(n18692) );
  NANDN U17586 ( .A(y[3318]), .B(x[3318]), .Z(n11343) );
  NANDN U17587 ( .A(n11344), .B(n11343), .Z(n27093) );
  NANDN U17588 ( .A(y[3317]), .B(x[3317]), .Z(n11346) );
  NANDN U17589 ( .A(y[3316]), .B(x[3316]), .Z(n11345) );
  NAND U17590 ( .A(n11346), .B(n11345), .Z(n27089) );
  NAND U17591 ( .A(n11347), .B(y[3316]), .Z(n11349) );
  ANDN U17592 ( .B(n11349), .A(n11348), .Z(n27086) );
  NAND U17593 ( .A(n11351), .B(n11350), .Z(n27083) );
  NANDN U17594 ( .A(x[3312]), .B(y[3312]), .Z(n11353) );
  NAND U17595 ( .A(n11353), .B(n11352), .Z(n27079) );
  NANDN U17596 ( .A(y[3311]), .B(x[3311]), .Z(n11355) );
  NANDN U17597 ( .A(y[3310]), .B(x[3310]), .Z(n11354) );
  AND U17598 ( .A(n11355), .B(n11354), .Z(n27076) );
  NAND U17599 ( .A(n11356), .B(y[3310]), .Z(n11357) );
  NANDN U17600 ( .A(n11358), .B(n11357), .Z(n27074) );
  NANDN U17601 ( .A(y[3307]), .B(x[3307]), .Z(n11360) );
  NANDN U17602 ( .A(y[3306]), .B(x[3306]), .Z(n11359) );
  NAND U17603 ( .A(n11360), .B(n11359), .Z(n27069) );
  NAND U17604 ( .A(n11361), .B(y[3306]), .Z(n11363) );
  AND U17605 ( .A(n11363), .B(n11362), .Z(n27066) );
  NANDN U17606 ( .A(y[3305]), .B(x[3305]), .Z(n11365) );
  NANDN U17607 ( .A(y[3304]), .B(x[3304]), .Z(n11364) );
  NAND U17608 ( .A(n11365), .B(n11364), .Z(n27064) );
  NANDN U17609 ( .A(x[3304]), .B(y[3304]), .Z(n11366) );
  NANDN U17610 ( .A(n11367), .B(n11366), .Z(n27063) );
  NAND U17611 ( .A(n11369), .B(n11368), .Z(n27059) );
  NANDN U17612 ( .A(y[3300]), .B(x[3300]), .Z(n11371) );
  NANDN U17613 ( .A(y[3301]), .B(x[3301]), .Z(n11370) );
  AND U17614 ( .A(n11371), .B(n11370), .Z(n27056) );
  NAND U17615 ( .A(n11372), .B(y[3300]), .Z(n11374) );
  NAND U17616 ( .A(n11374), .B(n11373), .Z(n27054) );
  NANDN U17617 ( .A(y[3299]), .B(x[3299]), .Z(n11376) );
  NANDN U17618 ( .A(y[3298]), .B(x[3298]), .Z(n11375) );
  NAND U17619 ( .A(n11376), .B(n11375), .Z(n27053) );
  AND U17620 ( .A(n11378), .B(n11377), .Z(n27046) );
  NANDN U17621 ( .A(y[3295]), .B(x[3295]), .Z(n11380) );
  NANDN U17622 ( .A(y[3294]), .B(x[3294]), .Z(n11379) );
  NAND U17623 ( .A(n11380), .B(n11379), .Z(n27044) );
  NANDN U17624 ( .A(x[3294]), .B(y[3294]), .Z(n11382) );
  NAND U17625 ( .A(n11382), .B(n11381), .Z(n27043) );
  NANDN U17626 ( .A(x[3292]), .B(y[3292]), .Z(n11383) );
  NANDN U17627 ( .A(n11384), .B(n11383), .Z(n27039) );
  NANDN U17628 ( .A(y[3290]), .B(x[3290]), .Z(n11386) );
  ANDN U17629 ( .B(n11386), .A(n11385), .Z(n27036) );
  NAND U17630 ( .A(n11388), .B(n11387), .Z(n27034) );
  NANDN U17631 ( .A(y[3289]), .B(x[3289]), .Z(n11390) );
  NANDN U17632 ( .A(y[3288]), .B(x[3288]), .Z(n11389) );
  NAND U17633 ( .A(n11390), .B(n11389), .Z(n27033) );
  NANDN U17634 ( .A(y[3287]), .B(x[3287]), .Z(n11392) );
  NANDN U17635 ( .A(y[3286]), .B(x[3286]), .Z(n11391) );
  NAND U17636 ( .A(n11392), .B(n11391), .Z(n27029) );
  NAND U17637 ( .A(n11393), .B(y[3286]), .Z(n11395) );
  ANDN U17638 ( .B(n11395), .A(n11394), .Z(n27026) );
  NAND U17639 ( .A(n11397), .B(n11396), .Z(n27023) );
  NANDN U17640 ( .A(x[3282]), .B(y[3282]), .Z(n11399) );
  NAND U17641 ( .A(n11399), .B(n11398), .Z(n27019) );
  NANDN U17642 ( .A(y[3281]), .B(x[3281]), .Z(n11401) );
  NANDN U17643 ( .A(y[3280]), .B(x[3280]), .Z(n11400) );
  AND U17644 ( .A(n11401), .B(n11400), .Z(n27016) );
  NAND U17645 ( .A(n11402), .B(y[3280]), .Z(n11403) );
  NANDN U17646 ( .A(n11404), .B(n11403), .Z(n27014) );
  NANDN U17647 ( .A(y[3277]), .B(x[3277]), .Z(n11406) );
  NANDN U17648 ( .A(y[3276]), .B(x[3276]), .Z(n11405) );
  NAND U17649 ( .A(n11406), .B(n11405), .Z(n27009) );
  NAND U17650 ( .A(n11407), .B(y[3276]), .Z(n11409) );
  ANDN U17651 ( .B(n11409), .A(n11408), .Z(n27006) );
  NANDN U17652 ( .A(x[3273]), .B(y[3273]), .Z(n11410) );
  NAND U17653 ( .A(n11411), .B(n11410), .Z(n27003) );
  NANDN U17654 ( .A(y[3270]), .B(x[3270]), .Z(n11412) );
  AND U17655 ( .A(n11413), .B(n11412), .Z(n26996) );
  NANDN U17656 ( .A(y[3263]), .B(x[3263]), .Z(n11414) );
  NANDN U17657 ( .A(n11415), .B(n11414), .Z(n26981) );
  NAND U17658 ( .A(n11416), .B(y[3259]), .Z(n11418) );
  ANDN U17659 ( .B(n11418), .A(n11417), .Z(n26974) );
  NANDN U17660 ( .A(y[3259]), .B(x[3259]), .Z(n11419) );
  NAND U17661 ( .A(n11420), .B(n11419), .Z(n26972) );
  OR U17662 ( .A(n11422), .B(n11421), .Z(n26969) );
  NANDN U17663 ( .A(x[3255]), .B(y[3255]), .Z(n11424) );
  ANDN U17664 ( .B(n11424), .A(n11423), .Z(n26966) );
  NAND U17665 ( .A(n11426), .B(n11425), .Z(n26964) );
  NANDN U17666 ( .A(x[3254]), .B(y[3254]), .Z(n11427) );
  NANDN U17667 ( .A(n11428), .B(n11427), .Z(n26963) );
  AND U17668 ( .A(n11430), .B(n11429), .Z(n26956) );
  NANDN U17669 ( .A(x[3250]), .B(y[3250]), .Z(n11431) );
  NANDN U17670 ( .A(n11432), .B(n11431), .Z(n26954) );
  OR U17671 ( .A(n11434), .B(n11433), .Z(n26953) );
  NAND U17672 ( .A(n11436), .B(n11435), .Z(n26949) );
  NANDN U17673 ( .A(x[3246]), .B(y[3246]), .Z(n11438) );
  ANDN U17674 ( .B(n11438), .A(n11437), .Z(n26946) );
  OR U17675 ( .A(n11440), .B(n11439), .Z(n26944) );
  NANDN U17676 ( .A(x[3242]), .B(y[3242]), .Z(n11441) );
  NANDN U17677 ( .A(n11442), .B(n11441), .Z(n26939) );
  NOR U17678 ( .A(n11444), .B(n11443), .Z(n26936) );
  NAND U17679 ( .A(n11446), .B(n11445), .Z(n26933) );
  OR U17680 ( .A(n11448), .B(n11447), .Z(n26929) );
  NANDN U17681 ( .A(x[3235]), .B(y[3235]), .Z(n11450) );
  ANDN U17682 ( .B(n11450), .A(n11449), .Z(n26926) );
  NAND U17683 ( .A(n11452), .B(n11451), .Z(n26924) );
  NANDN U17684 ( .A(x[3234]), .B(y[3234]), .Z(n11453) );
  NANDN U17685 ( .A(n11454), .B(n11453), .Z(n26923) );
  AND U17686 ( .A(n11456), .B(n11455), .Z(n26916) );
  NANDN U17687 ( .A(x[3230]), .B(y[3230]), .Z(n11457) );
  NANDN U17688 ( .A(n11458), .B(n11457), .Z(n26914) );
  OR U17689 ( .A(n11460), .B(n11459), .Z(n26913) );
  NAND U17690 ( .A(n11462), .B(n11461), .Z(n26909) );
  NANDN U17691 ( .A(x[3226]), .B(y[3226]), .Z(n11464) );
  ANDN U17692 ( .B(n11464), .A(n11463), .Z(n26906) );
  OR U17693 ( .A(n11466), .B(n11465), .Z(n26904) );
  NANDN U17694 ( .A(x[3222]), .B(y[3222]), .Z(n11467) );
  NANDN U17695 ( .A(n11468), .B(n11467), .Z(n26899) );
  NOR U17696 ( .A(n11470), .B(n11469), .Z(n26896) );
  NAND U17697 ( .A(n11472), .B(n11471), .Z(n26893) );
  OR U17698 ( .A(n11474), .B(n11473), .Z(n26889) );
  NANDN U17699 ( .A(x[3215]), .B(y[3215]), .Z(n11476) );
  ANDN U17700 ( .B(n11476), .A(n11475), .Z(n26886) );
  NAND U17701 ( .A(n11478), .B(n11477), .Z(n26884) );
  NANDN U17702 ( .A(x[3214]), .B(y[3214]), .Z(n11479) );
  NANDN U17703 ( .A(n11480), .B(n11479), .Z(n26883) );
  AND U17704 ( .A(n11482), .B(n11481), .Z(n26876) );
  NANDN U17705 ( .A(x[3210]), .B(y[3210]), .Z(n11483) );
  NANDN U17706 ( .A(n11484), .B(n11483), .Z(n26874) );
  OR U17707 ( .A(n11486), .B(n11485), .Z(n26873) );
  NAND U17708 ( .A(n11488), .B(n11487), .Z(n26869) );
  NANDN U17709 ( .A(x[3206]), .B(y[3206]), .Z(n11490) );
  ANDN U17710 ( .B(n11490), .A(n11489), .Z(n26866) );
  OR U17711 ( .A(n11492), .B(n11491), .Z(n26864) );
  NANDN U17712 ( .A(x[3202]), .B(y[3202]), .Z(n11493) );
  NANDN U17713 ( .A(n11494), .B(n11493), .Z(n26859) );
  NOR U17714 ( .A(n11496), .B(n11495), .Z(n26856) );
  NAND U17715 ( .A(n11498), .B(n11497), .Z(n26853) );
  OR U17716 ( .A(n11500), .B(n11499), .Z(n26849) );
  NANDN U17717 ( .A(x[3195]), .B(y[3195]), .Z(n11502) );
  ANDN U17718 ( .B(n11502), .A(n11501), .Z(n26846) );
  NAND U17719 ( .A(n11504), .B(n11503), .Z(n26844) );
  NANDN U17720 ( .A(x[3194]), .B(y[3194]), .Z(n11505) );
  NANDN U17721 ( .A(n11506), .B(n11505), .Z(n26843) );
  AND U17722 ( .A(n11508), .B(n11507), .Z(n26836) );
  NANDN U17723 ( .A(x[3190]), .B(y[3190]), .Z(n11509) );
  NANDN U17724 ( .A(n11510), .B(n11509), .Z(n26834) );
  OR U17725 ( .A(n11512), .B(n11511), .Z(n26833) );
  NAND U17726 ( .A(n11514), .B(n11513), .Z(n26829) );
  NANDN U17727 ( .A(x[3186]), .B(y[3186]), .Z(n11516) );
  ANDN U17728 ( .B(n11516), .A(n11515), .Z(n26826) );
  OR U17729 ( .A(n11518), .B(n11517), .Z(n26824) );
  NANDN U17730 ( .A(x[3182]), .B(y[3182]), .Z(n11519) );
  NANDN U17731 ( .A(n11520), .B(n11519), .Z(n26819) );
  NOR U17732 ( .A(n11522), .B(n11521), .Z(n26816) );
  NAND U17733 ( .A(n11524), .B(n11523), .Z(n26813) );
  OR U17734 ( .A(n11526), .B(n11525), .Z(n26809) );
  NANDN U17735 ( .A(y[3174]), .B(x[3174]), .Z(n11528) );
  NAND U17736 ( .A(n11528), .B(n11527), .Z(n26805) );
  NOR U17737 ( .A(n11530), .B(n11529), .Z(n26798) );
  OR U17738 ( .A(n11532), .B(n11531), .Z(n26796) );
  NANDN U17739 ( .A(y[3169]), .B(x[3169]), .Z(n11533) );
  NANDN U17740 ( .A(n11534), .B(n11533), .Z(n26791) );
  NOR U17741 ( .A(n11536), .B(n11535), .Z(n26788) );
  NAND U17742 ( .A(n11538), .B(n11537), .Z(n26785) );
  OR U17743 ( .A(n11540), .B(n11539), .Z(n26781) );
  NANDN U17744 ( .A(y[3162]), .B(x[3162]), .Z(n11542) );
  ANDN U17745 ( .B(n11542), .A(n11541), .Z(n26778) );
  NAND U17746 ( .A(n11544), .B(n11543), .Z(n26776) );
  NANDN U17747 ( .A(y[3161]), .B(x[3161]), .Z(n11545) );
  NANDN U17748 ( .A(n11546), .B(n11545), .Z(n26775) );
  ANDN U17749 ( .B(n11548), .A(n11547), .Z(n26768) );
  NANDN U17750 ( .A(y[3156]), .B(x[3156]), .Z(n11549) );
  NANDN U17751 ( .A(n11550), .B(n11549), .Z(n26766) );
  NANDN U17752 ( .A(x[3155]), .B(y[3155]), .Z(n11551) );
  NAND U17753 ( .A(n11552), .B(n11551), .Z(n26765) );
  NANDN U17754 ( .A(y[3152]), .B(x[3152]), .Z(n11553) );
  AND U17755 ( .A(n11554), .B(n11553), .Z(n26758) );
  NAND U17756 ( .A(n11556), .B(n11555), .Z(n26743) );
  NANDN U17757 ( .A(y[3143]), .B(x[3143]), .Z(n11558) );
  NAND U17758 ( .A(n11558), .B(n11557), .Z(n26738) );
  NANDN U17759 ( .A(x[3142]), .B(y[3142]), .Z(n11560) );
  NANDN U17760 ( .A(x[3141]), .B(y[3141]), .Z(n11559) );
  AND U17761 ( .A(n11560), .B(n11559), .Z(n26736) );
  NAND U17762 ( .A(n11561), .B(x[3141]), .Z(n11562) );
  NANDN U17763 ( .A(n11563), .B(n11562), .Z(n26735) );
  NANDN U17764 ( .A(x[3138]), .B(y[3138]), .Z(n11564) );
  NANDN U17765 ( .A(n11565), .B(n11564), .Z(n26728) );
  NOR U17766 ( .A(n11567), .B(n11566), .Z(n26726) );
  ANDN U17767 ( .B(n11569), .A(n11568), .Z(n26710) );
  NANDN U17768 ( .A(x[3128]), .B(y[3128]), .Z(n11570) );
  NANDN U17769 ( .A(n11571), .B(n11570), .Z(n26709) );
  OR U17770 ( .A(n11573), .B(n11572), .Z(n26707) );
  NANDN U17771 ( .A(x[3125]), .B(y[3125]), .Z(n11574) );
  NAND U17772 ( .A(n11575), .B(n11574), .Z(n26704) );
  NAND U17773 ( .A(n11577), .B(n11576), .Z(n26703) );
  NANDN U17774 ( .A(x[3124]), .B(y[3124]), .Z(n11579) );
  ANDN U17775 ( .B(n11579), .A(n11578), .Z(n26700) );
  OR U17776 ( .A(n11581), .B(n11580), .Z(n26699) );
  NAND U17777 ( .A(n11583), .B(n11582), .Z(n26694) );
  NANDN U17778 ( .A(x[3120]), .B(y[3120]), .Z(n11584) );
  NANDN U17779 ( .A(n11585), .B(n11584), .Z(n26693) );
  NOR U17780 ( .A(n11587), .B(n11586), .Z(n26690) );
  NAND U17781 ( .A(n11589), .B(n11588), .Z(n26687) );
  NANDN U17782 ( .A(x[3116]), .B(y[3116]), .Z(n11590) );
  NANDN U17783 ( .A(n11591), .B(n11590), .Z(n26684) );
  OR U17784 ( .A(n11593), .B(n11592), .Z(n26683) );
  NANDN U17785 ( .A(x[3113]), .B(y[3113]), .Z(n11595) );
  ANDN U17786 ( .B(n11595), .A(n11594), .Z(n26680) );
  NAND U17787 ( .A(n11597), .B(n11596), .Z(n26679) );
  NANDN U17788 ( .A(x[3112]), .B(y[3112]), .Z(n11598) );
  NANDN U17789 ( .A(n11599), .B(n11598), .Z(n26677) );
  OR U17790 ( .A(n11601), .B(n11600), .Z(n26674) );
  AND U17791 ( .A(n11603), .B(n11602), .Z(n26670) );
  NANDN U17792 ( .A(x[3108]), .B(y[3108]), .Z(n11604) );
  NANDN U17793 ( .A(n11605), .B(n11604), .Z(n26669) );
  OR U17794 ( .A(n11607), .B(n11606), .Z(n26667) );
  NANDN U17795 ( .A(x[3105]), .B(y[3105]), .Z(n11608) );
  NAND U17796 ( .A(n11609), .B(n11608), .Z(n26664) );
  NAND U17797 ( .A(n11611), .B(n11610), .Z(n26663) );
  NANDN U17798 ( .A(x[3104]), .B(y[3104]), .Z(n11613) );
  ANDN U17799 ( .B(n11613), .A(n11612), .Z(n26660) );
  OR U17800 ( .A(n11615), .B(n11614), .Z(n26659) );
  NANDN U17801 ( .A(n11617), .B(n11616), .Z(n26654) );
  NANDN U17802 ( .A(x[3099]), .B(y[3099]), .Z(n11618) );
  NANDN U17803 ( .A(n11619), .B(n11618), .Z(n26653) );
  ANDN U17804 ( .B(n11621), .A(n11620), .Z(n26650) );
  OR U17805 ( .A(n11623), .B(n11622), .Z(n26649) );
  NANDN U17806 ( .A(n11625), .B(n11624), .Z(n26644) );
  NANDN U17807 ( .A(y[3094]), .B(x[3094]), .Z(n11626) );
  NANDN U17808 ( .A(n11627), .B(n11626), .Z(n26643) );
  NAND U17809 ( .A(n11630), .B(x[3092]), .Z(n11629) );
  ANDN U17810 ( .B(n11629), .A(n11628), .Z(n26636) );
  XOR U17811 ( .A(n11630), .B(x[3092]), .Z(n18318) );
  NANDN U17812 ( .A(y[3088]), .B(x[3088]), .Z(n11632) );
  NAND U17813 ( .A(n11632), .B(n11631), .Z(n26627) );
  NANDN U17814 ( .A(x[3088]), .B(y[3088]), .Z(n11634) );
  NAND U17815 ( .A(n11634), .B(n11633), .Z(n26624) );
  NANDN U17816 ( .A(x[3086]), .B(y[3086]), .Z(n11635) );
  NANDN U17817 ( .A(n11636), .B(n11635), .Z(n26621) );
  NAND U17818 ( .A(n11638), .B(n11637), .Z(n26617) );
  NANDN U17819 ( .A(y[3083]), .B(x[3083]), .Z(n11640) );
  NANDN U17820 ( .A(y[3082]), .B(x[3082]), .Z(n11639) );
  NAND U17821 ( .A(n11640), .B(n11639), .Z(n26614) );
  NANDN U17822 ( .A(y[3081]), .B(x[3081]), .Z(n11642) );
  NANDN U17823 ( .A(y[3080]), .B(x[3080]), .Z(n11641) );
  NAND U17824 ( .A(n11642), .B(n11641), .Z(n26611) );
  NANDN U17825 ( .A(x[3075]), .B(y[3075]), .Z(n11644) );
  NAND U17826 ( .A(n11644), .B(n11643), .Z(n26601) );
  NANDN U17827 ( .A(n11646), .B(n11645), .Z(n26599) );
  NANDN U17828 ( .A(x[3073]), .B(y[3073]), .Z(n11647) );
  NANDN U17829 ( .A(n11648), .B(n11647), .Z(n26597) );
  NAND U17830 ( .A(n11649), .B(y[3072]), .Z(n11650) );
  NANDN U17831 ( .A(n11651), .B(n11650), .Z(n26593) );
  OR U17832 ( .A(n11653), .B(n11652), .Z(n26588) );
  NANDN U17833 ( .A(n11654), .B(n26583), .Z(n18272) );
  NOR U17834 ( .A(n11656), .B(n11655), .Z(n18270) );
  ANDN U17835 ( .B(n26575), .A(n11657), .Z(n18266) );
  NANDN U17836 ( .A(y[3064]), .B(x[3064]), .Z(n11658) );
  NANDN U17837 ( .A(n11659), .B(n11658), .Z(n26573) );
  NANDN U17838 ( .A(n11661), .B(n11660), .Z(n26571) );
  ANDN U17839 ( .B(n26566), .A(n11662), .Z(n18259) );
  NANDN U17840 ( .A(x[3057]), .B(y[3057]), .Z(n11663) );
  NANDN U17841 ( .A(n11664), .B(n11663), .Z(n26554) );
  NOR U17842 ( .A(n11666), .B(n11665), .Z(n18238) );
  NOR U17843 ( .A(n11668), .B(n11667), .Z(n26532) );
  AND U17844 ( .A(n11669), .B(n26528), .Z(n18224) );
  ANDN U17845 ( .B(x[3046]), .A(y[3046]), .Z(n11670) );
  ANDN U17846 ( .B(n11671), .A(n11670), .Z(n18222) );
  AND U17847 ( .A(n11672), .B(n26512), .Z(n18208) );
  NOR U17848 ( .A(n11674), .B(n11673), .Z(n26496) );
  AND U17849 ( .A(n11675), .B(n26492), .Z(n18184) );
  ANDN U17850 ( .B(x[3032]), .A(y[3032]), .Z(n11676) );
  ANDN U17851 ( .B(n11677), .A(n11676), .Z(n18182) );
  NOR U17852 ( .A(n11679), .B(n11678), .Z(n18162) );
  AND U17853 ( .A(n26466), .B(n11680), .Z(n18160) );
  NANDN U17854 ( .A(n11681), .B(n26464), .Z(n18158) );
  OR U17855 ( .A(n11683), .B(n11682), .Z(n26461) );
  ANDN U17856 ( .B(n26458), .A(n11684), .Z(n18152) );
  AND U17857 ( .A(n26456), .B(n11685), .Z(n18150) );
  XOR U17858 ( .A(n11686), .B(y[3018]), .Z(n18144) );
  ANDN U17859 ( .B(n26446), .A(n11687), .Z(n18141) );
  OR U17860 ( .A(n11689), .B(n11688), .Z(n26442) );
  AND U17861 ( .A(n26438), .B(n11690), .Z(n18132) );
  NOR U17862 ( .A(n11692), .B(n11691), .Z(n26424) );
  AND U17863 ( .A(n11693), .B(n26420), .Z(n18113) );
  ANDN U17864 ( .B(n11695), .A(n11694), .Z(n18111) );
  ANDN U17865 ( .B(n26410), .A(n11696), .Z(n18106) );
  OR U17866 ( .A(n11698), .B(n11697), .Z(n26406) );
  AND U17867 ( .A(n26402), .B(n11699), .Z(n18097) );
  NOR U17868 ( .A(n11701), .B(n11700), .Z(n26388) );
  AND U17869 ( .A(n11702), .B(n26384), .Z(n18078) );
  ANDN U17870 ( .B(n11704), .A(n11703), .Z(n18076) );
  ANDN U17871 ( .B(n26374), .A(n11705), .Z(n18071) );
  OR U17872 ( .A(n11707), .B(n11706), .Z(n26370) );
  AND U17873 ( .A(n26366), .B(n11708), .Z(n18062) );
  NOR U17874 ( .A(n11710), .B(n11709), .Z(n26352) );
  AND U17875 ( .A(n11711), .B(n26348), .Z(n18043) );
  ANDN U17876 ( .B(n11713), .A(n11712), .Z(n18041) );
  ANDN U17877 ( .B(n26338), .A(n11714), .Z(n18036) );
  OR U17878 ( .A(n11716), .B(n11715), .Z(n26334) );
  AND U17879 ( .A(n26330), .B(n11717), .Z(n18027) );
  NOR U17880 ( .A(n11719), .B(n11718), .Z(n26316) );
  ANDN U17881 ( .B(n26312), .A(n11720), .Z(n18008) );
  ANDN U17882 ( .B(n11722), .A(n11721), .Z(n18006) );
  ANDN U17883 ( .B(n26303), .A(n11723), .Z(n18001) );
  OR U17884 ( .A(n11725), .B(n11724), .Z(n26301) );
  OR U17885 ( .A(n11727), .B(n11726), .Z(n26299) );
  ANDN U17886 ( .B(n26294), .A(n11728), .Z(n17994) );
  NANDN U17887 ( .A(n11730), .B(n11729), .Z(n26282) );
  NAND U17888 ( .A(n11731), .B(n26270), .Z(n17969) );
  NANDN U17889 ( .A(x[2945]), .B(y[2945]), .Z(n11733) );
  ANDN U17890 ( .B(n11733), .A(n11732), .Z(n26268) );
  NANDN U17891 ( .A(n11735), .B(n11734), .Z(n26266) );
  ANDN U17892 ( .B(n26264), .A(n11736), .Z(n17965) );
  ANDN U17893 ( .B(n11737), .A(n26262), .Z(n17963) );
  AND U17894 ( .A(n26247), .B(n11738), .Z(n17948) );
  NANDN U17895 ( .A(y[2934]), .B(x[2934]), .Z(n17940) );
  ANDN U17896 ( .B(n26234), .A(n11739), .Z(n17935) );
  OR U17897 ( .A(n11741), .B(n11740), .Z(n26232) );
  NOR U17898 ( .A(n11743), .B(n11742), .Z(n17926) );
  ANDN U17899 ( .B(n11745), .A(n11744), .Z(n17924) );
  NANDN U17900 ( .A(y[2924]), .B(x[2924]), .Z(n11746) );
  NANDN U17901 ( .A(n11747), .B(n11746), .Z(n26214) );
  ANDN U17902 ( .B(n26210), .A(n11748), .Z(n17912) );
  NANDN U17903 ( .A(x[2917]), .B(y[2917]), .Z(n11749) );
  NANDN U17904 ( .A(n11750), .B(n11749), .Z(n26197) );
  ANDN U17905 ( .B(n11752), .A(n11751), .Z(n26194) );
  OR U17906 ( .A(n11753), .B(n26178), .Z(n17886) );
  NANDN U17907 ( .A(n11755), .B(n11754), .Z(n11757) );
  ANDN U17908 ( .B(n11757), .A(n11756), .Z(n17880) );
  NANDN U17909 ( .A(x[2903]), .B(y[2903]), .Z(n11758) );
  NANDN U17910 ( .A(n11759), .B(n11758), .Z(n26162) );
  ANDN U17911 ( .B(n11761), .A(n11760), .Z(n26160) );
  ANDN U17912 ( .B(n26158), .A(n11762), .Z(n17872) );
  NANDN U17913 ( .A(y[2896]), .B(x[2896]), .Z(n11763) );
  NANDN U17914 ( .A(n11764), .B(n11763), .Z(n26144) );
  AND U17915 ( .A(n26139), .B(n11765), .Z(n17849) );
  NOR U17916 ( .A(n11767), .B(n11766), .Z(n17847) );
  NAND U17917 ( .A(n11768), .B(n26131), .Z(n17845) );
  ANDN U17918 ( .B(n26128), .A(n11769), .Z(n17843) );
  NANDN U17919 ( .A(x[2889]), .B(y[2889]), .Z(n11770) );
  NANDN U17920 ( .A(n11771), .B(n11770), .Z(n26126) );
  AND U17921 ( .A(n11772), .B(n26114), .Z(n17828) );
  OR U17922 ( .A(n11774), .B(n11773), .Z(n26112) );
  OR U17923 ( .A(n11776), .B(n11775), .Z(n26110) );
  NOR U17924 ( .A(n26107), .B(n11777), .Z(n17821) );
  AND U17925 ( .A(n11779), .B(n11778), .Z(n17819) );
  XNOR U17926 ( .A(x[2878]), .B(y[2878]), .Z(n17817) );
  NANDN U17927 ( .A(y[2875]), .B(x[2875]), .Z(n11780) );
  NANDN U17928 ( .A(n11781), .B(n11780), .Z(n26093) );
  NOR U17929 ( .A(n26091), .B(n11782), .Z(n17806) );
  AND U17930 ( .A(n26088), .B(n11783), .Z(n17804) );
  XNOR U17931 ( .A(x[2872]), .B(y[2872]), .Z(n17802) );
  ANDN U17932 ( .B(n11785), .A(n11784), .Z(n17795) );
  NAND U17933 ( .A(n11787), .B(n11786), .Z(n17787) );
  NOR U17934 ( .A(n11789), .B(n11788), .Z(n17785) );
  ANDN U17935 ( .B(n26064), .A(n11790), .Z(n17780) );
  NANDN U17936 ( .A(y[2854]), .B(x[2854]), .Z(n11791) );
  NANDN U17937 ( .A(n11792), .B(n11791), .Z(n26040) );
  NAND U17938 ( .A(n11793), .B(y[2854]), .Z(n11795) );
  ANDN U17939 ( .B(n11795), .A(n11794), .Z(n26038) );
  AND U17940 ( .A(n11797), .B(n11796), .Z(n17755) );
  OR U17941 ( .A(n11799), .B(n11798), .Z(n26023) );
  AND U17942 ( .A(n11801), .B(n11800), .Z(n17721) );
  XNOR U17943 ( .A(y[2835]), .B(x[2835]), .Z(n17719) );
  NOR U17944 ( .A(n11803), .B(n11802), .Z(n25980) );
  NAND U17945 ( .A(n25966), .B(n25974), .Z(n17706) );
  OR U17946 ( .A(x[2828]), .B(n11804), .Z(n25970) );
  AND U17947 ( .A(n25970), .B(n25964), .Z(n17704) );
  NOR U17948 ( .A(n25956), .B(n11805), .Z(n17697) );
  ANDN U17949 ( .B(n25950), .A(n11806), .Z(n17695) );
  OR U17950 ( .A(n11808), .B(n11807), .Z(n25944) );
  NAND U17951 ( .A(n11810), .B(n11809), .Z(n11811) );
  NANDN U17952 ( .A(n11812), .B(n11811), .Z(n11814) );
  ANDN U17953 ( .B(n11814), .A(n11813), .Z(n25923) );
  NANDN U17954 ( .A(n11815), .B(n25921), .Z(n17674) );
  NOR U17955 ( .A(n25919), .B(n11816), .Z(n17672) );
  ANDN U17956 ( .B(x[2808]), .A(y[2808]), .Z(n11817) );
  ANDN U17957 ( .B(n11818), .A(n11817), .Z(n17670) );
  XOR U17958 ( .A(n11819), .B(y[2808]), .Z(n17667) );
  NOR U17959 ( .A(n25909), .B(n11820), .Z(n17665) );
  NANDN U17960 ( .A(x[2805]), .B(y[2805]), .Z(n11821) );
  NANDN U17961 ( .A(n11822), .B(n11821), .Z(n25908) );
  NANDN U17962 ( .A(n11824), .B(n11823), .Z(n25906) );
  ANDN U17963 ( .B(n25901), .A(n11825), .Z(n17658) );
  NANDN U17964 ( .A(y[2798]), .B(x[2798]), .Z(n11826) );
  NANDN U17965 ( .A(n11827), .B(n11826), .Z(n25889) );
  AND U17966 ( .A(n25884), .B(n11828), .Z(n17639) );
  NANDN U17967 ( .A(x[2785]), .B(y[2785]), .Z(n11829) );
  NANDN U17968 ( .A(n11830), .B(n11829), .Z(n25852) );
  AND U17969 ( .A(n25821), .B(n11831), .Z(n17596) );
  AND U17970 ( .A(n11833), .B(n11832), .Z(n17594) );
  XOR U17971 ( .A(y[2767]), .B(n11834), .Z(n17592) );
  XOR U17972 ( .A(n11835), .B(y[2766]), .Z(n17588) );
  AND U17973 ( .A(n25809), .B(n11836), .Z(n17585) );
  OR U17974 ( .A(n11838), .B(n11837), .Z(n25807) );
  NOR U17975 ( .A(n11840), .B(n11839), .Z(n17576) );
  AND U17976 ( .A(n11842), .B(n11841), .Z(n17574) );
  NANDN U17977 ( .A(n11843), .B(n25792), .Z(n17572) );
  AND U17978 ( .A(n25791), .B(n11844), .Z(n17570) );
  NANDN U17979 ( .A(y[2756]), .B(x[2756]), .Z(n11845) );
  NANDN U17980 ( .A(n11846), .B(n11845), .Z(n25789) );
  NANDN U17981 ( .A(n11848), .B(n11847), .Z(n25787) );
  ANDN U17982 ( .B(n25776), .A(n11849), .Z(n17561) );
  OR U17983 ( .A(n11851), .B(n11850), .Z(n25775) );
  OR U17984 ( .A(n11853), .B(n11852), .Z(n25773) );
  NANDN U17985 ( .A(x[2749]), .B(y[2749]), .Z(n11854) );
  NANDN U17986 ( .A(n11855), .B(n11854), .Z(n25771) );
  ANDN U17987 ( .B(n25765), .A(n11856), .Z(n17550) );
  AND U17988 ( .A(n11858), .B(n11857), .Z(n17548) );
  XOR U17989 ( .A(y[2745]), .B(n11859), .Z(n17546) );
  NANDN U17990 ( .A(y[2740]), .B(x[2740]), .Z(n11860) );
  AND U17991 ( .A(n25748), .B(n11860), .Z(n17538) );
  OR U17992 ( .A(n11862), .B(n11861), .Z(n25737) );
  NAND U17993 ( .A(n11863), .B(y[2735]), .Z(n11864) );
  NANDN U17994 ( .A(n11865), .B(n11864), .Z(n25735) );
  AND U17995 ( .A(n25729), .B(n11866), .Z(n17518) );
  AND U17996 ( .A(n11868), .B(n11867), .Z(n17516) );
  XNOR U17997 ( .A(y[2731]), .B(x[2731]), .Z(n17514) );
  ANDN U17998 ( .B(n25718), .A(n11869), .Z(n17511) );
  NANDN U17999 ( .A(y[2728]), .B(x[2728]), .Z(n11870) );
  NANDN U18000 ( .A(n11871), .B(n11870), .Z(n25716) );
  OR U18001 ( .A(n11872), .B(n25712), .Z(n17505) );
  ANDN U18002 ( .B(n25710), .A(n11873), .Z(n17503) );
  ANDN U18003 ( .B(n11875), .A(n11874), .Z(n17474) );
  NANDN U18004 ( .A(n11877), .B(n11876), .Z(n11879) );
  ANDN U18005 ( .B(n11879), .A(n11878), .Z(n17459) );
  AND U18006 ( .A(n25678), .B(n11880), .Z(n17456) );
  OR U18007 ( .A(n11882), .B(n11881), .Z(n25677) );
  AND U18008 ( .A(n25647), .B(n11883), .Z(n17438) );
  ANDN U18009 ( .B(n11885), .A(n11884), .Z(n17436) );
  NANDN U18010 ( .A(x[2679]), .B(y[2679]), .Z(n11886) );
  NANDN U18011 ( .A(n11887), .B(n11886), .Z(n25595) );
  NANDN U18012 ( .A(n11889), .B(n11888), .Z(n25594) );
  NANDN U18013 ( .A(n11891), .B(n11890), .Z(n17399) );
  OR U18014 ( .A(n11893), .B(n11892), .Z(n25581) );
  NOR U18015 ( .A(n25576), .B(n11894), .Z(n17384) );
  ANDN U18016 ( .B(n11896), .A(n11895), .Z(n17382) );
  OR U18017 ( .A(n11898), .B(n11897), .Z(n25563) );
  NOR U18018 ( .A(n11900), .B(n11899), .Z(n25561) );
  NOR U18019 ( .A(n11902), .B(n11901), .Z(n17366) );
  ANDN U18020 ( .B(n25549), .A(n11903), .Z(n17364) );
  NANDN U18021 ( .A(n11904), .B(n25548), .Z(n17362) );
  NAND U18022 ( .A(n11905), .B(x[2658]), .Z(n11907) );
  ANDN U18023 ( .B(n11907), .A(n11906), .Z(n25545) );
  NANDN U18024 ( .A(x[2658]), .B(y[2658]), .Z(n11908) );
  NANDN U18025 ( .A(n11909), .B(n11908), .Z(n25544) );
  ANDN U18026 ( .B(n25541), .A(n11910), .Z(n17358) );
  NAND U18027 ( .A(n11912), .B(n11911), .Z(n25530) );
  NANDN U18028 ( .A(x[2652]), .B(y[2652]), .Z(n11913) );
  NANDN U18029 ( .A(n11914), .B(n11913), .Z(n25528) );
  NANDN U18030 ( .A(n11916), .B(n11915), .Z(n25514) );
  NOR U18031 ( .A(n11918), .B(n11917), .Z(n25511) );
  AND U18032 ( .A(n25507), .B(n11919), .Z(n17331) );
  ANDN U18033 ( .B(n11921), .A(n11920), .Z(n17329) );
  NOR U18034 ( .A(n11923), .B(n11922), .Z(n17318) );
  OR U18035 ( .A(n11925), .B(n11924), .Z(n11926) );
  NANDN U18036 ( .A(n11927), .B(n11926), .Z(n11928) );
  NANDN U18037 ( .A(n11929), .B(n11928), .Z(n25481) );
  NANDN U18038 ( .A(n11930), .B(n25479), .Z(n17308) );
  AND U18039 ( .A(n11932), .B(n11931), .Z(n17299) );
  OR U18040 ( .A(n11934), .B(n11933), .Z(n25464) );
  ANDN U18041 ( .B(n25462), .A(n11935), .Z(n17290) );
  NOR U18042 ( .A(n25455), .B(n11936), .Z(n17286) );
  NANDN U18043 ( .A(n25447), .B(n25454), .Z(n17284) );
  ANDN U18044 ( .B(n25427), .A(n11937), .Z(n17263) );
  OR U18045 ( .A(n11939), .B(n11938), .Z(n25409) );
  NANDN U18046 ( .A(y[2600]), .B(x[2600]), .Z(n11941) );
  ANDN U18047 ( .B(n11941), .A(n11940), .Z(n25407) );
  NAND U18048 ( .A(n11943), .B(n11942), .Z(n25406) );
  NANDN U18049 ( .A(y[2599]), .B(x[2599]), .Z(n11945) );
  NANDN U18050 ( .A(y[2598]), .B(x[2598]), .Z(n11944) );
  AND U18051 ( .A(n11945), .B(n11944), .Z(n25403) );
  AND U18052 ( .A(n11947), .B(n11946), .Z(n17225) );
  XOR U18053 ( .A(y[2591]), .B(n11948), .Z(n17223) );
  NANDN U18054 ( .A(y[2590]), .B(x[2590]), .Z(n17221) );
  NANDN U18055 ( .A(n11950), .B(n11949), .Z(n11951) );
  NANDN U18056 ( .A(n11952), .B(n11951), .Z(n20243) );
  AND U18057 ( .A(n25377), .B(n11953), .Z(n17209) );
  OR U18058 ( .A(n11955), .B(n11954), .Z(n25362) );
  OR U18059 ( .A(n11957), .B(n11956), .Z(n25313) );
  ANDN U18060 ( .B(n25307), .A(n11958), .Z(n17154) );
  AND U18061 ( .A(n11960), .B(n11959), .Z(n17152) );
  XNOR U18062 ( .A(y[2555]), .B(x[2555]), .Z(n17150) );
  NAND U18063 ( .A(n11961), .B(x[2552]), .Z(n11963) );
  ANDN U18064 ( .B(n11963), .A(n11962), .Z(n25295) );
  NANDN U18065 ( .A(x[2552]), .B(y[2552]), .Z(n11964) );
  NANDN U18066 ( .A(n11965), .B(n11964), .Z(n25293) );
  ANDN U18067 ( .B(n25291), .A(n11966), .Z(n17142) );
  ANDN U18068 ( .B(n25282), .A(n11967), .Z(n17134) );
  ANDN U18069 ( .B(n25259), .A(n11968), .Z(n17112) );
  NOR U18070 ( .A(n11970), .B(n11969), .Z(n25247) );
  ANDN U18071 ( .B(n25243), .A(n11971), .Z(n17099) );
  NOR U18072 ( .A(n11973), .B(n11972), .Z(n17097) );
  OR U18073 ( .A(n11975), .B(n11974), .Z(n17095) );
  ANDN U18074 ( .B(n25222), .A(n11976), .Z(n17079) );
  AND U18075 ( .A(n25215), .B(n11977), .Z(n17077) );
  NANDN U18076 ( .A(n11979), .B(n11978), .Z(n17069) );
  AND U18077 ( .A(n11981), .B(n11980), .Z(n17057) );
  NOR U18078 ( .A(n11983), .B(n11982), .Z(n17055) );
  NAND U18079 ( .A(n11985), .B(n11984), .Z(n17053) );
  NOR U18080 ( .A(n11987), .B(n11986), .Z(n17051) );
  NANDN U18081 ( .A(x[2503]), .B(y[2503]), .Z(n11988) );
  NANDN U18082 ( .A(n11989), .B(n11988), .Z(n25183) );
  NAND U18083 ( .A(n11990), .B(y[2502]), .Z(n11991) );
  NANDN U18084 ( .A(n11992), .B(n11991), .Z(n25180) );
  ANDN U18085 ( .B(n25177), .A(n11993), .Z(n17038) );
  OR U18086 ( .A(n11995), .B(n11994), .Z(n25151) );
  NANDN U18087 ( .A(n11997), .B(n11996), .Z(n11998) );
  AND U18088 ( .A(n25145), .B(n11998), .Z(n17014) );
  NOR U18089 ( .A(n12000), .B(n11999), .Z(n25133) );
  NOR U18090 ( .A(n12002), .B(n12001), .Z(n16996) );
  OR U18091 ( .A(n12004), .B(n12003), .Z(n16994) );
  OR U18092 ( .A(n12006), .B(n12005), .Z(n25116) );
  ANDN U18093 ( .B(n25096), .A(n12007), .Z(n16972) );
  NANDN U18094 ( .A(x[2460]), .B(y[2460]), .Z(n12008) );
  NANDN U18095 ( .A(n12009), .B(n12008), .Z(n25082) );
  NOR U18096 ( .A(n25080), .B(n12010), .Z(n16958) );
  AND U18097 ( .A(n25077), .B(n12011), .Z(n16956) );
  XOR U18098 ( .A(y[2457]), .B(n12012), .Z(n16954) );
  OR U18099 ( .A(n12013), .B(n25067), .Z(n16947) );
  AND U18100 ( .A(n12015), .B(n12014), .Z(n16936) );
  XOR U18101 ( .A(x[2450]), .B(n12016), .Z(n16934) );
  NANDN U18102 ( .A(n12018), .B(n12017), .Z(n12019) );
  NANDN U18103 ( .A(n12020), .B(n12019), .Z(n25049) );
  ANDN U18104 ( .B(n25047), .A(n12021), .Z(n16924) );
  ANDN U18105 ( .B(n25033), .A(n12022), .Z(n16911) );
  OR U18106 ( .A(n12024), .B(n12023), .Z(n25032) );
  NANDN U18107 ( .A(n12026), .B(n12025), .Z(n12027) );
  NANDN U18108 ( .A(n12028), .B(n12027), .Z(n24984) );
  NANDN U18109 ( .A(x[2419]), .B(y[2419]), .Z(n12029) );
  NANDN U18110 ( .A(n12030), .B(n12029), .Z(n24982) );
  ANDN U18111 ( .B(n24971), .A(n12031), .Z(n16860) );
  ANDN U18112 ( .B(n24966), .A(n12032), .Z(n16858) );
  NANDN U18113 ( .A(n12033), .B(n24963), .Z(n16856) );
  NOR U18114 ( .A(n24937), .B(n12034), .Z(n16836) );
  AND U18115 ( .A(n12036), .B(n12035), .Z(n16834) );
  XOR U18116 ( .A(y[2401]), .B(n12037), .Z(n16832) );
  NANDN U18117 ( .A(y[2400]), .B(x[2400]), .Z(n16830) );
  OR U18118 ( .A(n12038), .B(n24925), .Z(n16825) );
  NAND U18119 ( .A(n12040), .B(n12039), .Z(n24907) );
  NANDN U18120 ( .A(y[2391]), .B(x[2391]), .Z(n12041) );
  NANDN U18121 ( .A(n12042), .B(n12041), .Z(n24905) );
  NAND U18122 ( .A(n12043), .B(n24903), .Z(n16810) );
  NANDN U18123 ( .A(n12045), .B(n12044), .Z(n12046) );
  NANDN U18124 ( .A(n12047), .B(n12046), .Z(n24878) );
  NANDN U18125 ( .A(n12048), .B(n24873), .Z(n16759) );
  ANDN U18126 ( .B(n24872), .A(n12049), .Z(n16757) );
  OR U18127 ( .A(n12051), .B(n12050), .Z(n24857) );
  NOR U18128 ( .A(n24852), .B(n12052), .Z(n16738) );
  AND U18129 ( .A(n12054), .B(n12053), .Z(n16736) );
  XOR U18130 ( .A(y[2365]), .B(n12055), .Z(n16734) );
  NAND U18131 ( .A(n12057), .B(n12056), .Z(n16732) );
  XOR U18132 ( .A(y[2360]), .B(n12058), .Z(n16719) );
  NAND U18133 ( .A(n12060), .B(n12059), .Z(n12062) );
  ANDN U18134 ( .B(n12062), .A(n12061), .Z(n16711) );
  NOR U18135 ( .A(n12064), .B(n12063), .Z(n16692) );
  ANDN U18136 ( .B(n24803), .A(n12065), .Z(n16687) );
  NANDN U18137 ( .A(y[2342]), .B(x[2342]), .Z(n12066) );
  NANDN U18138 ( .A(n12067), .B(n12066), .Z(n24802) );
  ANDN U18139 ( .B(n24795), .A(n12068), .Z(n16678) );
  NANDN U18140 ( .A(n12070), .B(n12069), .Z(n12071) );
  NANDN U18141 ( .A(n12072), .B(n12071), .Z(n12073) );
  NANDN U18142 ( .A(n12074), .B(n12073), .Z(n24786) );
  NANDN U18143 ( .A(n12076), .B(n12075), .Z(n12078) );
  ANDN U18144 ( .B(n12078), .A(n12077), .Z(n16658) );
  NOR U18145 ( .A(n24749), .B(n12079), .Z(n16645) );
  AND U18146 ( .A(n12081), .B(n12080), .Z(n16643) );
  XNOR U18147 ( .A(y[2317]), .B(x[2317]), .Z(n16641) );
  NANDN U18148 ( .A(n12082), .B(n24736), .Z(n16634) );
  OR U18149 ( .A(n12084), .B(n12083), .Z(n24735) );
  NANDN U18150 ( .A(n12086), .B(n12085), .Z(n12087) );
  AND U18151 ( .A(n24730), .B(n12087), .Z(n16630) );
  XOR U18152 ( .A(n12088), .B(x[2309]), .Z(n16621) );
  NOR U18153 ( .A(n12090), .B(n12089), .Z(n16618) );
  NOR U18154 ( .A(n12092), .B(n12091), .Z(n16607) );
  OR U18155 ( .A(n12094), .B(n12093), .Z(n16605) );
  NAND U18156 ( .A(n12095), .B(n24697), .Z(n16594) );
  ANDN U18157 ( .B(n24694), .A(n12096), .Z(n16592) );
  ANDN U18158 ( .B(n24684), .A(n12097), .Z(n16583) );
  OR U18159 ( .A(n12099), .B(n12098), .Z(n24682) );
  NANDN U18160 ( .A(n12101), .B(n12100), .Z(n24679) );
  NANDN U18161 ( .A(n12103), .B(n12102), .Z(n12104) );
  AND U18162 ( .A(n24626), .B(n12104), .Z(n16537) );
  AND U18163 ( .A(n12106), .B(n12105), .Z(n16525) );
  XNOR U18164 ( .A(y[2260]), .B(x[2260]), .Z(n16523) );
  XNOR U18165 ( .A(x[2254]), .B(y[2254]), .Z(n16511) );
  ANDN U18166 ( .B(n24592), .A(n12107), .Z(n16499) );
  AND U18167 ( .A(n24580), .B(n12108), .Z(n16485) );
  NANDN U18168 ( .A(n12109), .B(n24574), .Z(n16477) );
  AND U18169 ( .A(n24573), .B(n12110), .Z(n16475) );
  XNOR U18170 ( .A(n12112), .B(n12111), .Z(n16473) );
  NANDN U18171 ( .A(y[2240]), .B(x[2240]), .Z(n16471) );
  ANDN U18172 ( .B(n24562), .A(n12113), .Z(n12118) );
  OR U18173 ( .A(n12115), .B(n12114), .Z(n24558) );
  NANDN U18174 ( .A(n12116), .B(n24558), .Z(n12117) );
  NAND U18175 ( .A(n12118), .B(n12117), .Z(n16466) );
  ANDN U18176 ( .B(n12120), .A(n12119), .Z(n16464) );
  XNOR U18177 ( .A(y[2234]), .B(x[2234]), .Z(n16459) );
  XOR U18178 ( .A(x[2212]), .B(n12121), .Z(n12123) );
  AND U18179 ( .A(n12123), .B(n12122), .Z(n12127) );
  NANDN U18180 ( .A(n12125), .B(n12124), .Z(n12126) );
  NAND U18181 ( .A(n12127), .B(n12126), .Z(n24495) );
  NAND U18182 ( .A(n12128), .B(y[2209]), .Z(n12129) );
  NANDN U18183 ( .A(n12130), .B(n12129), .Z(n24493) );
  NANDN U18184 ( .A(y[2209]), .B(x[2209]), .Z(n12131) );
  NANDN U18185 ( .A(n12132), .B(n12131), .Z(n24490) );
  NAND U18186 ( .A(n12133), .B(n24478), .Z(n16406) );
  OR U18187 ( .A(n12135), .B(n12134), .Z(n24457) );
  ANDN U18188 ( .B(n24442), .A(n12136), .Z(n16379) );
  NAND U18189 ( .A(n12137), .B(y[2181]), .Z(n12138) );
  NANDN U18190 ( .A(n12139), .B(n12138), .Z(n24425) );
  NANDN U18191 ( .A(y[2181]), .B(x[2181]), .Z(n12140) );
  NANDN U18192 ( .A(n12141), .B(n12140), .Z(n24422) );
  AND U18193 ( .A(n12143), .B(n12142), .Z(n16328) );
  XNOR U18194 ( .A(x[2170]), .B(y[2170]), .Z(n16326) );
  NANDN U18195 ( .A(y[2167]), .B(x[2167]), .Z(n12144) );
  NANDN U18196 ( .A(n12145), .B(n12144), .Z(n24390) );
  XNOR U18197 ( .A(y[2164]), .B(x[2164]), .Z(n16309) );
  AND U18198 ( .A(n24366), .B(n12146), .Z(n16292) );
  AND U18199 ( .A(n12148), .B(n12147), .Z(n16290) );
  XOR U18200 ( .A(y[2155]), .B(n12149), .Z(n16288) );
  NANDN U18201 ( .A(n12151), .B(n12150), .Z(n12152) );
  NANDN U18202 ( .A(n12153), .B(n12152), .Z(n12154) );
  NANDN U18203 ( .A(n12155), .B(n12154), .Z(n24329) );
  ANDN U18204 ( .B(n24314), .A(n12156), .Z(n16248) );
  OR U18205 ( .A(n12158), .B(n12157), .Z(n24312) );
  NAND U18206 ( .A(n12159), .B(n24308), .Z(n16242) );
  OR U18207 ( .A(n12161), .B(n12160), .Z(n24260) );
  ANDN U18208 ( .B(n12162), .A(n24240), .Z(n16171) );
  AND U18209 ( .A(n12164), .B(n12163), .Z(n16169) );
  XOR U18210 ( .A(y[2099]), .B(n12165), .Z(n16167) );
  XNOR U18211 ( .A(n12167), .B(n12166), .Z(n16163) );
  NANDN U18212 ( .A(y[2096]), .B(x[2096]), .Z(n20262) );
  ANDN U18213 ( .B(n20262), .A(n12168), .Z(n16160) );
  ANDN U18214 ( .B(y[2096]), .A(x[2096]), .Z(n20260) );
  OR U18215 ( .A(n20261), .B(n12169), .Z(n12171) );
  ANDN U18216 ( .B(n12171), .A(n12170), .Z(n16157) );
  OR U18217 ( .A(n12172), .B(x[2093]), .Z(n12175) );
  XOR U18218 ( .A(n12172), .B(x[2093]), .Z(n12173) );
  NAND U18219 ( .A(n12173), .B(y[2093]), .Z(n12174) );
  NAND U18220 ( .A(n12175), .B(n12174), .Z(n16154) );
  AND U18221 ( .A(n24214), .B(n12176), .Z(n16141) );
  XNOR U18222 ( .A(x[2087]), .B(y[2087]), .Z(n16139) );
  NANDN U18223 ( .A(y[2086]), .B(x[2086]), .Z(n16137) );
  NANDN U18224 ( .A(x[2083]), .B(y[2083]), .Z(n12177) );
  NANDN U18225 ( .A(n12178), .B(n12177), .Z(n24202) );
  NANDN U18226 ( .A(n12180), .B(n12179), .Z(n24200) );
  XOR U18227 ( .A(x[2079]), .B(n12181), .Z(n16118) );
  OR U18228 ( .A(n12183), .B(n12182), .Z(n24166) );
  XOR U18229 ( .A(y[2064]), .B(n12184), .Z(n16085) );
  ANDN U18230 ( .B(n24149), .A(n12185), .Z(n16082) );
  OR U18231 ( .A(n12187), .B(n12186), .Z(n24148) );
  AND U18232 ( .A(n24145), .B(n12188), .Z(n16079) );
  AND U18233 ( .A(n24143), .B(n12189), .Z(n16077) );
  XOR U18234 ( .A(y[2059]), .B(n12190), .Z(n16075) );
  ANDN U18235 ( .B(n24105), .A(n12191), .Z(n16032) );
  AND U18236 ( .A(n24103), .B(n12192), .Z(n16030) );
  XOR U18237 ( .A(x[2038]), .B(n12193), .Z(n16028) );
  XOR U18238 ( .A(n12194), .B(x[2037]), .Z(n16024) );
  ANDN U18239 ( .B(n24093), .A(n12195), .Z(n16021) );
  OR U18240 ( .A(n12197), .B(n12196), .Z(n24092) );
  OR U18241 ( .A(n12198), .B(n24087), .Z(n16015) );
  OR U18242 ( .A(n12200), .B(n12199), .Z(n24071) );
  NOR U18243 ( .A(n24055), .B(n12201), .Z(n15985) );
  OR U18244 ( .A(n12203), .B(n12202), .Z(n24054) );
  NANDN U18245 ( .A(x[1999]), .B(y[1999]), .Z(n12204) );
  NANDN U18246 ( .A(n12205), .B(n12204), .Z(n24010) );
  ANDN U18247 ( .B(n24004), .A(n12206), .Z(n15941) );
  AND U18248 ( .A(n12208), .B(n12207), .Z(n15939) );
  XOR U18249 ( .A(y[1995]), .B(n12209), .Z(n15937) );
  XNOR U18250 ( .A(x[1994]), .B(y[1994]), .Z(n15933) );
  AND U18251 ( .A(n23992), .B(n12210), .Z(n15930) );
  OR U18252 ( .A(n12212), .B(n12211), .Z(n23990) );
  OR U18253 ( .A(n12214), .B(n12213), .Z(n23969) );
  AND U18254 ( .A(n23966), .B(n12215), .Z(n15914) );
  AND U18255 ( .A(n12217), .B(n12216), .Z(n15912) );
  XNOR U18256 ( .A(y[1981]), .B(x[1981]), .Z(n15910) );
  NANDN U18257 ( .A(n12219), .B(n12218), .Z(n23931) );
  XNOR U18258 ( .A(x[1960]), .B(n12220), .Z(n23908) );
  NANDN U18259 ( .A(n12222), .B(n12221), .Z(n12223) );
  NANDN U18260 ( .A(n12224), .B(n12223), .Z(n23904) );
  NANDN U18261 ( .A(n12226), .B(n12225), .Z(n15859) );
  NANDN U18262 ( .A(n23886), .B(n23890), .Z(n15856) );
  NANDN U18263 ( .A(n12228), .B(n12227), .Z(n23841) );
  OR U18264 ( .A(n12230), .B(n12229), .Z(n23820) );
  NANDN U18265 ( .A(n12232), .B(n12231), .Z(n12233) );
  NANDN U18266 ( .A(n12234), .B(n12233), .Z(n23804) );
  NANDN U18267 ( .A(y[1902]), .B(x[1902]), .Z(n12235) );
  NANDN U18268 ( .A(n12236), .B(n12235), .Z(n23771) );
  NANDN U18269 ( .A(y[1901]), .B(x[1901]), .Z(n12237) );
  NANDN U18270 ( .A(n12238), .B(n12237), .Z(n23768) );
  NOR U18271 ( .A(n23766), .B(n12239), .Z(n15768) );
  AND U18272 ( .A(n23763), .B(n12240), .Z(n15766) );
  XOR U18273 ( .A(x[1898]), .B(n12241), .Z(n15764) );
  AND U18274 ( .A(n12243), .B(n12242), .Z(n15760) );
  XOR U18275 ( .A(x[1896]), .B(n12244), .Z(n15758) );
  NANDN U18276 ( .A(n12246), .B(n12245), .Z(n12247) );
  NANDN U18277 ( .A(n12248), .B(n12247), .Z(n15727) );
  NANDN U18278 ( .A(n12250), .B(n12249), .Z(n23722) );
  AND U18279 ( .A(n23719), .B(n12251), .Z(n15717) );
  AND U18280 ( .A(n23717), .B(n12252), .Z(n15715) );
  XOR U18281 ( .A(y[1877]), .B(n12253), .Z(n15713) );
  NANDN U18282 ( .A(n12255), .B(n12254), .Z(n15680) );
  NAND U18283 ( .A(n12257), .B(n12256), .Z(n23676) );
  NANDN U18284 ( .A(y[1859]), .B(x[1859]), .Z(n12258) );
  NANDN U18285 ( .A(n12259), .B(n12258), .Z(n23674) );
  ANDN U18286 ( .B(n23671), .A(n12260), .Z(n15667) );
  NANDN U18287 ( .A(n12262), .B(n12261), .Z(n12263) );
  NANDN U18288 ( .A(n12264), .B(n12263), .Z(n23660) );
  AND U18289 ( .A(n23658), .B(n12265), .Z(n15655) );
  ANDN U18290 ( .B(n23647), .A(n12266), .Z(n15646) );
  NOR U18291 ( .A(n23644), .B(n12267), .Z(n15637) );
  NANDN U18292 ( .A(x[1837]), .B(y[1837]), .Z(n12269) );
  ANDN U18293 ( .B(n12269), .A(n12268), .Z(n23623) );
  NANDN U18294 ( .A(n12271), .B(n12270), .Z(n23622) );
  OR U18295 ( .A(n12273), .B(n12272), .Z(n23603) );
  AND U18296 ( .A(n23589), .B(n12274), .Z(n15606) );
  NANDN U18297 ( .A(x[1824]), .B(y[1824]), .Z(n12275) );
  NANDN U18298 ( .A(n12276), .B(n12275), .Z(n23579) );
  NANDN U18299 ( .A(n12278), .B(n12277), .Z(n12279) );
  AND U18300 ( .A(n23573), .B(n12279), .Z(n15595) );
  ANDN U18301 ( .B(x[1816]), .A(y[1816]), .Z(n23559) );
  OR U18302 ( .A(x[1816]), .B(n12280), .Z(n23561) );
  ANDN U18303 ( .B(n23561), .A(n12281), .Z(n15580) );
  ANDN U18304 ( .B(n12282), .A(n23556), .Z(n15578) );
  XOR U18305 ( .A(x[1814]), .B(n12283), .Z(n15576) );
  XNOR U18306 ( .A(y[1813]), .B(x[1813]), .Z(n15572) );
  ANDN U18307 ( .B(n23544), .A(n12284), .Z(n15564) );
  OR U18308 ( .A(n12286), .B(n12285), .Z(n23542) );
  ANDN U18309 ( .B(n23540), .A(n12287), .Z(n15561) );
  ANDN U18310 ( .B(n23528), .A(n12288), .Z(n15549) );
  OR U18311 ( .A(n12290), .B(n12289), .Z(n23527) );
  XOR U18312 ( .A(x[1792]), .B(y[1792]), .Z(n23499) );
  NANDN U18313 ( .A(y[1790]), .B(x[1790]), .Z(n12291) );
  NANDN U18314 ( .A(n12292), .B(n12291), .Z(n23495) );
  NAND U18315 ( .A(n12294), .B(n12293), .Z(n23493) );
  NANDN U18316 ( .A(y[1789]), .B(x[1789]), .Z(n12295) );
  NANDN U18317 ( .A(n12296), .B(n12295), .Z(n23491) );
  OR U18318 ( .A(n12298), .B(n12297), .Z(n23472) );
  NANDN U18319 ( .A(n12300), .B(n12299), .Z(n12301) );
  NANDN U18320 ( .A(n12302), .B(n12301), .Z(n23459) );
  NANDN U18321 ( .A(n12304), .B(n12303), .Z(n15504) );
  NANDN U18322 ( .A(n12306), .B(n12305), .Z(n12307) );
  NANDN U18323 ( .A(n12308), .B(n12307), .Z(n23415) );
  AND U18324 ( .A(n12310), .B(n12309), .Z(n15476) );
  XNOR U18325 ( .A(y[1751]), .B(x[1751]), .Z(n15474) );
  XNOR U18326 ( .A(x[1730]), .B(y[1730]), .Z(n15435) );
  OR U18327 ( .A(n12312), .B(n12311), .Z(n23338) );
  NANDN U18328 ( .A(x[1713]), .B(y[1713]), .Z(n12313) );
  NANDN U18329 ( .A(n12314), .B(n12313), .Z(n23329) );
  NAND U18330 ( .A(n12316), .B(n12315), .Z(n23327) );
  NANDN U18331 ( .A(x[1711]), .B(y[1711]), .Z(n12318) );
  NANDN U18332 ( .A(x[1712]), .B(y[1712]), .Z(n12317) );
  NAND U18333 ( .A(n12318), .B(n12317), .Z(n23324) );
  NANDN U18334 ( .A(n12320), .B(n12319), .Z(n23323) );
  NANDN U18335 ( .A(n12322), .B(n12321), .Z(n12323) );
  NANDN U18336 ( .A(n12324), .B(n12323), .Z(n23309) );
  AND U18337 ( .A(n23306), .B(n12325), .Z(n15401) );
  XOR U18338 ( .A(x[1700]), .B(n12326), .Z(n15391) );
  AND U18339 ( .A(n12328), .B(n12327), .Z(n15387) );
  XNOR U18340 ( .A(x[1698]), .B(y[1698]), .Z(n15385) );
  XNOR U18341 ( .A(y[1697]), .B(x[1697]), .Z(n15381) );
  ANDN U18342 ( .B(n23280), .A(n12329), .Z(n15366) );
  NANDN U18343 ( .A(x[1691]), .B(y[1691]), .Z(n12330) );
  NANDN U18344 ( .A(n12331), .B(n12330), .Z(n23278) );
  NAND U18345 ( .A(n12332), .B(n23274), .Z(n15360) );
  AND U18346 ( .A(n12334), .B(n12333), .Z(n15351) );
  XOR U18347 ( .A(x[1686]), .B(n12335), .Z(n15349) );
  NOR U18348 ( .A(n12337), .B(n12336), .Z(n23258) );
  AND U18349 ( .A(n12339), .B(n12338), .Z(n15332) );
  XNOR U18350 ( .A(y[1679]), .B(x[1679]), .Z(n15330) );
  NOR U18351 ( .A(n12341), .B(n12340), .Z(n15319) );
  AND U18352 ( .A(n23240), .B(n12342), .Z(n15317) );
  XNOR U18353 ( .A(x[1674]), .B(y[1674]), .Z(n15315) );
  NOR U18354 ( .A(n12344), .B(n12343), .Z(n23230) );
  NANDN U18355 ( .A(y[1670]), .B(x[1670]), .Z(n12345) );
  NANDN U18356 ( .A(n12346), .B(n12345), .Z(n23228) );
  NANDN U18357 ( .A(n12348), .B(n12347), .Z(n23227) );
  AND U18358 ( .A(n23224), .B(n12349), .Z(n15306) );
  AND U18359 ( .A(n23222), .B(n12350), .Z(n15304) );
  XOR U18360 ( .A(y[1667]), .B(n12351), .Z(n15302) );
  NANDN U18361 ( .A(x[1651]), .B(y[1651]), .Z(n12352) );
  NANDN U18362 ( .A(n12353), .B(n12352), .Z(n23190) );
  NANDN U18363 ( .A(x[1649]), .B(y[1649]), .Z(n12354) );
  NANDN U18364 ( .A(n12355), .B(n12354), .Z(n23187) );
  NANDN U18365 ( .A(n12357), .B(n12356), .Z(n12358) );
  NANDN U18366 ( .A(n12359), .B(n12358), .Z(n23171) );
  ANDN U18367 ( .B(n20276), .A(n12360), .Z(n15235) );
  ANDN U18368 ( .B(n23146), .A(n12361), .Z(n15226) );
  OR U18369 ( .A(n12363), .B(n12362), .Z(n23141) );
  NANDN U18370 ( .A(x[1622]), .B(y[1622]), .Z(n12365) );
  NANDN U18371 ( .A(x[1621]), .B(y[1621]), .Z(n12364) );
  NAND U18372 ( .A(n12365), .B(n12364), .Z(n23118) );
  ANDN U18373 ( .B(n12367), .A(n12366), .Z(n23115) );
  NOR U18374 ( .A(n12369), .B(n12368), .Z(n23103) );
  ANDN U18375 ( .B(n23089), .A(n12370), .Z(n15185) );
  NANDN U18376 ( .A(y[1608]), .B(x[1608]), .Z(n12371) );
  NANDN U18377 ( .A(n12372), .B(n12371), .Z(n23087) );
  NANDN U18378 ( .A(y[1607]), .B(x[1607]), .Z(n12373) );
  NANDN U18379 ( .A(n12374), .B(n12373), .Z(n23084) );
  NANDN U18380 ( .A(x[1596]), .B(y[1596]), .Z(n12375) );
  NAND U18381 ( .A(n12376), .B(n12375), .Z(n23061) );
  NANDN U18382 ( .A(y[1595]), .B(x[1595]), .Z(n12377) );
  NANDN U18383 ( .A(n12378), .B(n12377), .Z(n23059) );
  ANDN U18384 ( .B(n23057), .A(n12379), .Z(n15163) );
  NANDN U18385 ( .A(n23055), .B(n23051), .Z(n15161) );
  NANDN U18386 ( .A(n12381), .B(n12380), .Z(n23032) );
  NANDN U18387 ( .A(n12383), .B(n12382), .Z(n12385) );
  ANDN U18388 ( .B(n12385), .A(n12384), .Z(n23028) );
  OR U18389 ( .A(n12387), .B(n12386), .Z(n12388) );
  NANDN U18390 ( .A(n12389), .B(n12388), .Z(n12391) );
  ANDN U18391 ( .B(n12391), .A(n12390), .Z(n23011) );
  AND U18392 ( .A(n23001), .B(n12392), .Z(n15126) );
  NANDN U18393 ( .A(n12394), .B(n12393), .Z(n22997) );
  NANDN U18394 ( .A(y[1560]), .B(x[1560]), .Z(n12395) );
  NANDN U18395 ( .A(n12396), .B(n12395), .Z(n22988) );
  NANDN U18396 ( .A(y[1558]), .B(x[1558]), .Z(n12398) );
  NANDN U18397 ( .A(y[1559]), .B(x[1559]), .Z(n12397) );
  NAND U18398 ( .A(n12398), .B(n12397), .Z(n22984) );
  NAND U18399 ( .A(n12399), .B(y[1558]), .Z(n12401) );
  ANDN U18400 ( .B(n12401), .A(n12400), .Z(n22981) );
  NANDN U18401 ( .A(n22976), .B(n22980), .Z(n15112) );
  ANDN U18402 ( .B(n22977), .A(n22974), .Z(n15110) );
  NANDN U18403 ( .A(y[1554]), .B(x[1554]), .Z(n12402) );
  NANDN U18404 ( .A(n12403), .B(n12402), .Z(n22971) );
  NANDN U18405 ( .A(x[1547]), .B(y[1547]), .Z(n12404) );
  NANDN U18406 ( .A(n12405), .B(n12404), .Z(n22957) );
  NANDN U18407 ( .A(x[1546]), .B(y[1546]), .Z(n12406) );
  NANDN U18408 ( .A(n12407), .B(n12406), .Z(n22954) );
  OR U18409 ( .A(n12408), .B(n22947), .Z(n15090) );
  OR U18410 ( .A(n12410), .B(n12409), .Z(n22944) );
  OR U18411 ( .A(n12412), .B(n12411), .Z(n12413) );
  NANDN U18412 ( .A(n12414), .B(n12413), .Z(n12416) );
  ANDN U18413 ( .B(n12416), .A(n12415), .Z(n22933) );
  ANDN U18414 ( .B(n22930), .A(n22926), .Z(n15076) );
  ANDN U18415 ( .B(n22923), .A(n12417), .Z(n15074) );
  NANDN U18416 ( .A(n12419), .B(n12418), .Z(n22922) );
  NANDN U18417 ( .A(n12421), .B(n12420), .Z(n22896) );
  NANDN U18418 ( .A(x[1511]), .B(y[1511]), .Z(n12422) );
  NANDN U18419 ( .A(n12423), .B(n12422), .Z(n22884) );
  OR U18420 ( .A(n12425), .B(n12424), .Z(n20282) );
  IV U18421 ( .A(n20282), .Z(n15035) );
  NAND U18422 ( .A(n12426), .B(x[1500]), .Z(n12427) );
  NANDN U18423 ( .A(n12428), .B(n12427), .Z(n22866) );
  NANDN U18424 ( .A(x[1500]), .B(y[1500]), .Z(n12429) );
  NAND U18425 ( .A(n12430), .B(n12429), .Z(n22863) );
  NANDN U18426 ( .A(y[1499]), .B(x[1499]), .Z(n12432) );
  ANDN U18427 ( .B(n12432), .A(n12431), .Z(n22861) );
  AND U18428 ( .A(n22857), .B(n22853), .Z(n15021) );
  NAND U18429 ( .A(n12434), .B(n12433), .Z(n22840) );
  NANDN U18430 ( .A(y[1488]), .B(x[1488]), .Z(n12436) );
  NANDN U18431 ( .A(y[1489]), .B(x[1489]), .Z(n12435) );
  NAND U18432 ( .A(n12436), .B(n12435), .Z(n22838) );
  NANDN U18433 ( .A(x[1488]), .B(y[1488]), .Z(n12437) );
  NAND U18434 ( .A(n12438), .B(n12437), .Z(n22836) );
  NANDN U18435 ( .A(y[1487]), .B(x[1487]), .Z(n12439) );
  NANDN U18436 ( .A(n12440), .B(n12439), .Z(n22833) );
  ANDN U18437 ( .B(n22823), .A(n12441), .Z(n15000) );
  NANDN U18438 ( .A(y[1482]), .B(x[1482]), .Z(n12442) );
  NANDN U18439 ( .A(n12443), .B(n12442), .Z(n22821) );
  NANDN U18440 ( .A(x[1477]), .B(y[1477]), .Z(n12444) );
  NANDN U18441 ( .A(n12445), .B(n12444), .Z(n22812) );
  NANDN U18442 ( .A(n12447), .B(n12446), .Z(n22810) );
  NANDN U18443 ( .A(y[1474]), .B(x[1474]), .Z(n12448) );
  NAND U18444 ( .A(n12449), .B(n12448), .Z(n22806) );
  NAND U18445 ( .A(n12450), .B(y[1474]), .Z(n12452) );
  ANDN U18446 ( .B(n12452), .A(n12451), .Z(n22803) );
  NANDN U18447 ( .A(n12453), .B(n22802), .Z(n14983) );
  NANDN U18448 ( .A(y[1470]), .B(x[1470]), .Z(n12454) );
  NANDN U18449 ( .A(n12455), .B(n12454), .Z(n22793) );
  ANDN U18450 ( .B(n22771), .A(n12456), .Z(n22768) );
  NANDN U18451 ( .A(x[1453]), .B(y[1453]), .Z(n12457) );
  NANDN U18452 ( .A(n12458), .B(n12457), .Z(n22755) );
  ANDN U18453 ( .B(n12460), .A(n12459), .Z(n22752) );
  NANDN U18454 ( .A(x[1451]), .B(y[1451]), .Z(n12461) );
  NANDN U18455 ( .A(n12462), .B(n12461), .Z(n22750) );
  ANDN U18456 ( .B(n12464), .A(n12463), .Z(n22748) );
  ANDN U18457 ( .B(n22741), .A(n22744), .Z(n14943) );
  NANDN U18458 ( .A(y[1442]), .B(x[1442]), .Z(n12465) );
  NANDN U18459 ( .A(n12466), .B(n12465), .Z(n22729) );
  NANDN U18460 ( .A(n12468), .B(n12467), .Z(n22727) );
  NANDN U18461 ( .A(y[1440]), .B(x[1440]), .Z(n12469) );
  NANDN U18462 ( .A(n12470), .B(n12469), .Z(n22725) );
  NANDN U18463 ( .A(y[1439]), .B(x[1439]), .Z(n12471) );
  NANDN U18464 ( .A(n12472), .B(n12471), .Z(n22721) );
  NANDN U18465 ( .A(x[1429]), .B(y[1429]), .Z(n12473) );
  NANDN U18466 ( .A(n12474), .B(n12473), .Z(n22702) );
  NAND U18467 ( .A(n12476), .B(n12475), .Z(n22700) );
  NANDN U18468 ( .A(x[1427]), .B(y[1427]), .Z(n12478) );
  NANDN U18469 ( .A(x[1428]), .B(y[1428]), .Z(n12477) );
  NAND U18470 ( .A(n12478), .B(n12477), .Z(n22698) );
  AND U18471 ( .A(n12479), .B(n22694), .Z(n14909) );
  NAND U18472 ( .A(n22688), .B(n22693), .Z(n14907) );
  NOR U18473 ( .A(n22687), .B(n12480), .Z(n14905) );
  NANDN U18474 ( .A(x[1417]), .B(y[1417]), .Z(n12481) );
  NANDN U18475 ( .A(n12482), .B(n12481), .Z(n22675) );
  NANDN U18476 ( .A(x[1415]), .B(y[1415]), .Z(n12483) );
  NANDN U18477 ( .A(n12484), .B(n12483), .Z(n22671) );
  NANDN U18478 ( .A(n12486), .B(n12485), .Z(n22669) );
  NANDN U18479 ( .A(y[1404]), .B(x[1404]), .Z(n12487) );
  NANDN U18480 ( .A(n12488), .B(n12487), .Z(n22652) );
  ANDN U18481 ( .B(n12490), .A(n12489), .Z(n22650) );
  OR U18482 ( .A(n12492), .B(n12491), .Z(n22649) );
  NANDN U18483 ( .A(y[1394]), .B(x[1394]), .Z(n12493) );
  NANDN U18484 ( .A(n12494), .B(n12493), .Z(n22633) );
  NANDN U18485 ( .A(n12496), .B(n12495), .Z(n22631) );
  NANDN U18486 ( .A(y[1392]), .B(x[1392]), .Z(n12497) );
  NANDN U18487 ( .A(n12498), .B(n12497), .Z(n22629) );
  NANDN U18488 ( .A(n12500), .B(n12499), .Z(n22627) );
  NANDN U18489 ( .A(n12502), .B(n12501), .Z(n22623) );
  NANDN U18490 ( .A(n12504), .B(n12503), .Z(n22607) );
  NANDN U18491 ( .A(y[1378]), .B(x[1378]), .Z(n12505) );
  NANDN U18492 ( .A(n12506), .B(n12505), .Z(n22605) );
  OR U18493 ( .A(n12507), .B(n12510), .Z(n12508) );
  NAND U18494 ( .A(n12509), .B(n12508), .Z(n22603) );
  OR U18495 ( .A(n12511), .B(n12510), .Z(n22600) );
  ANDN U18496 ( .B(n22578), .A(n12512), .Z(n14821) );
  AND U18497 ( .A(n12514), .B(n12513), .Z(n22560) );
  NANDN U18498 ( .A(x[1354]), .B(y[1354]), .Z(n12517) );
  NANDN U18499 ( .A(n12519), .B(n12515), .Z(n12516) );
  NAND U18500 ( .A(n12517), .B(n12516), .Z(n22559) );
  OR U18501 ( .A(n12519), .B(n12518), .Z(n22557) );
  NANDN U18502 ( .A(n12521), .B(n12520), .Z(n12522) );
  NANDN U18503 ( .A(n12523), .B(n12522), .Z(n22554) );
  NANDN U18504 ( .A(x[1345]), .B(y[1345]), .Z(n12524) );
  NANDN U18505 ( .A(n12525), .B(n12524), .Z(n22547) );
  NANDN U18506 ( .A(x[1343]), .B(y[1343]), .Z(n12526) );
  NANDN U18507 ( .A(n12527), .B(n12526), .Z(n22543) );
  NANDN U18508 ( .A(n12529), .B(n12528), .Z(n22541) );
  AND U18509 ( .A(n22530), .B(n12530), .Z(n14791) );
  AND U18510 ( .A(n12532), .B(n12531), .Z(n22512) );
  NANDN U18511 ( .A(x[1330]), .B(y[1330]), .Z(n12533) );
  NANDN U18512 ( .A(n12534), .B(n12533), .Z(n22511) );
  OR U18513 ( .A(n12535), .B(n22504), .Z(n14772) );
  NANDN U18514 ( .A(x[1321]), .B(y[1321]), .Z(n12536) );
  NANDN U18515 ( .A(n12537), .B(n12536), .Z(n22492) );
  NANDN U18516 ( .A(y[1321]), .B(x[1321]), .Z(n12538) );
  AND U18517 ( .A(n12539), .B(n12538), .Z(n22490) );
  NANDN U18518 ( .A(x[1319]), .B(y[1319]), .Z(n12541) );
  NANDN U18519 ( .A(x[1320]), .B(y[1320]), .Z(n12540) );
  NAND U18520 ( .A(n12541), .B(n12540), .Z(n22489) );
  NAND U18521 ( .A(n12542), .B(x[1319]), .Z(n12544) );
  ANDN U18522 ( .B(n12544), .A(n12543), .Z(n22486) );
  ANDN U18523 ( .B(n22482), .A(n22479), .Z(n14756) );
  ANDN U18524 ( .B(n22476), .A(n12545), .Z(n14754) );
  NOR U18525 ( .A(n12547), .B(n12546), .Z(n22472) );
  NANDN U18526 ( .A(y[1308]), .B(x[1308]), .Z(n12549) );
  ANDN U18527 ( .B(n12549), .A(n12548), .Z(n22462) );
  NANDN U18528 ( .A(y[1307]), .B(x[1307]), .Z(n12550) );
  NANDN U18529 ( .A(n12551), .B(n12550), .Z(n22459) );
  NANDN U18530 ( .A(n12553), .B(n12552), .Z(n12555) );
  ANDN U18531 ( .B(n12555), .A(n12554), .Z(n22455) );
  NANDN U18532 ( .A(n12557), .B(n12556), .Z(n22452) );
  OR U18533 ( .A(n12559), .B(n12558), .Z(n22434) );
  ANDN U18534 ( .B(n22432), .A(n12560), .Z(n14727) );
  NANDN U18535 ( .A(y[1290]), .B(x[1290]), .Z(n12561) );
  NANDN U18536 ( .A(n12562), .B(n12561), .Z(n22422) );
  NAND U18537 ( .A(n12563), .B(y[1290]), .Z(n12564) );
  NANDN U18538 ( .A(n12565), .B(n12564), .Z(n22421) );
  ANDN U18539 ( .B(n12567), .A(n12566), .Z(n22410) );
  NANDN U18540 ( .A(x[1283]), .B(y[1283]), .Z(n12568) );
  NANDN U18541 ( .A(n12569), .B(n12568), .Z(n22408) );
  NANDN U18542 ( .A(n12571), .B(n12570), .Z(n22407) );
  NANDN U18543 ( .A(n12573), .B(n12572), .Z(n12575) );
  ANDN U18544 ( .B(n12575), .A(n12574), .Z(n22403) );
  NANDN U18545 ( .A(x[1273]), .B(y[1273]), .Z(n12576) );
  NANDN U18546 ( .A(n12577), .B(n12576), .Z(n22388) );
  NAND U18547 ( .A(n12578), .B(x[1273]), .Z(n12579) );
  NANDN U18548 ( .A(n12580), .B(n12579), .Z(n22387) );
  NANDN U18549 ( .A(y[1271]), .B(x[1271]), .Z(n12581) );
  NANDN U18550 ( .A(n12582), .B(n12581), .Z(n22382) );
  ANDN U18551 ( .B(n22380), .A(n12583), .Z(n14690) );
  NANDN U18552 ( .A(n22378), .B(n22374), .Z(n14688) );
  OR U18553 ( .A(n12585), .B(n12584), .Z(n22371) );
  NANDN U18554 ( .A(x[1261]), .B(y[1261]), .Z(n12586) );
  NANDN U18555 ( .A(n12587), .B(n12586), .Z(n22361) );
  NANDN U18556 ( .A(n12589), .B(n12588), .Z(n22359) );
  NANDN U18557 ( .A(n12591), .B(n12590), .Z(n22355) );
  AND U18558 ( .A(n22346), .B(n22350), .Z(n14667) );
  NANDN U18559 ( .A(n12593), .B(n12592), .Z(n22341) );
  NANDN U18560 ( .A(x[1247]), .B(y[1247]), .Z(n12594) );
  NANDN U18561 ( .A(n12595), .B(n12594), .Z(n22329) );
  NAND U18562 ( .A(n12597), .B(n12596), .Z(n22327) );
  NANDN U18563 ( .A(x[1246]), .B(y[1246]), .Z(n12600) );
  OR U18564 ( .A(n12598), .B(n12601), .Z(n12599) );
  NAND U18565 ( .A(n12600), .B(n12599), .Z(n22325) );
  OR U18566 ( .A(n12602), .B(n12601), .Z(n22323) );
  NANDN U18567 ( .A(x[1237]), .B(y[1237]), .Z(n12603) );
  NANDN U18568 ( .A(n12604), .B(n12603), .Z(n22313) );
  NANDN U18569 ( .A(n12606), .B(n12605), .Z(n22311) );
  NANDN U18570 ( .A(n12608), .B(n12607), .Z(n22307) );
  AND U18571 ( .A(n22296), .B(n12609), .Z(n14635) );
  NOR U18572 ( .A(n12611), .B(n12610), .Z(n22292) );
  NANDN U18573 ( .A(n12613), .B(n12612), .Z(n12614) );
  NANDN U18574 ( .A(n12615), .B(n12614), .Z(n22279) );
  OR U18575 ( .A(n12617), .B(n12616), .Z(n22259) );
  ANDN U18576 ( .B(n22256), .A(n12618), .Z(n14606) );
  NOR U18577 ( .A(n12620), .B(n12619), .Z(n22244) );
  NAND U18578 ( .A(n22230), .B(n22226), .Z(n14583) );
  NANDN U18579 ( .A(x[1194]), .B(y[1194]), .Z(n12622) );
  NAND U18580 ( .A(n12622), .B(n12621), .Z(n22220) );
  NAND U18581 ( .A(n12624), .B(n12623), .Z(n22211) );
  OR U18582 ( .A(n12626), .B(n12625), .Z(n22207) );
  ANDN U18583 ( .B(n22204), .A(n12627), .Z(n14562) );
  NANDN U18584 ( .A(y[1176]), .B(x[1176]), .Z(n12628) );
  NANDN U18585 ( .A(n12629), .B(n12628), .Z(n22183) );
  NANDN U18586 ( .A(y[1175]), .B(x[1175]), .Z(n12630) );
  NANDN U18587 ( .A(n12631), .B(n12630), .Z(n22178) );
  ANDN U18588 ( .B(n22175), .A(n12632), .Z(n14544) );
  AND U18589 ( .A(n12634), .B(n12633), .Z(n14540) );
  NOR U18590 ( .A(n12636), .B(n12635), .Z(n14521) );
  NANDN U18591 ( .A(n12638), .B(n12637), .Z(n22139) );
  OR U18592 ( .A(n14501), .B(n12639), .Z(n22133) );
  OR U18593 ( .A(n12641), .B(n12640), .Z(n22117) );
  ANDN U18594 ( .B(n22114), .A(n12642), .Z(n14490) );
  NAND U18595 ( .A(n22108), .B(n22113), .Z(n14488) );
  ANDN U18596 ( .B(n22106), .A(n12643), .Z(n14486) );
  NANDN U18597 ( .A(y[1128]), .B(x[1128]), .Z(n12644) );
  NANDN U18598 ( .A(n12645), .B(n12644), .Z(n22093) );
  NANDN U18599 ( .A(y[1127]), .B(x[1127]), .Z(n12646) );
  NANDN U18600 ( .A(n12647), .B(n12646), .Z(n22089) );
  ANDN U18601 ( .B(n22086), .A(n12648), .Z(n14469) );
  NANDN U18602 ( .A(n22084), .B(n22080), .Z(n14467) );
  ANDN U18603 ( .B(n22078), .A(n12649), .Z(n14465) );
  NANDN U18604 ( .A(y[1122]), .B(x[1122]), .Z(n12650) );
  NANDN U18605 ( .A(n12651), .B(n12650), .Z(n22077) );
  NAND U18606 ( .A(n12652), .B(y[1122]), .Z(n12654) );
  ANDN U18607 ( .B(n12654), .A(n12653), .Z(n22074) );
  ANDN U18608 ( .B(n22054), .A(n12655), .Z(n14451) );
  OR U18609 ( .A(n12657), .B(n12656), .Z(n22053) );
  AND U18610 ( .A(n22049), .B(n22050), .Z(n14448) );
  NANDN U18611 ( .A(n12659), .B(n12658), .Z(n12660) );
  NANDN U18612 ( .A(n12661), .B(n12660), .Z(n12663) );
  NAND U18613 ( .A(n12663), .B(n12662), .Z(n22039) );
  ANDN U18614 ( .B(n22028), .A(n12664), .Z(n14436) );
  NANDN U18615 ( .A(y[1098]), .B(x[1098]), .Z(n12665) );
  NANDN U18616 ( .A(n12666), .B(n12665), .Z(n22027) );
  NANDN U18617 ( .A(n12668), .B(n12667), .Z(n22009) );
  OR U18618 ( .A(n12670), .B(n12669), .Z(n22005) );
  NANDN U18619 ( .A(x[1081]), .B(y[1081]), .Z(n12671) );
  NANDN U18620 ( .A(n12672), .B(n12671), .Z(n21997) );
  ANDN U18621 ( .B(n12674), .A(n12673), .Z(n21994) );
  NANDN U18622 ( .A(x[1079]), .B(y[1079]), .Z(n12675) );
  NANDN U18623 ( .A(n12676), .B(n12675), .Z(n21993) );
  ANDN U18624 ( .B(n21989), .A(n12677), .Z(n14400) );
  OR U18625 ( .A(n12679), .B(n12678), .Z(n21977) );
  NANDN U18626 ( .A(y[1062]), .B(x[1062]), .Z(n12680) );
  NANDN U18627 ( .A(n12681), .B(n12680), .Z(n21954) );
  NANDN U18628 ( .A(n12683), .B(n12682), .Z(n21953) );
  NANDN U18629 ( .A(n12685), .B(n12684), .Z(n12686) );
  NANDN U18630 ( .A(n12687), .B(n12686), .Z(n12689) );
  NAND U18631 ( .A(n12689), .B(n12688), .Z(n21943) );
  NOR U18632 ( .A(n21941), .B(n12690), .Z(n14371) );
  ANDN U18633 ( .B(n21932), .A(n12691), .Z(n14367) );
  NANDN U18634 ( .A(y[1050]), .B(x[1050]), .Z(n12692) );
  NANDN U18635 ( .A(n12693), .B(n12692), .Z(n21931) );
  NAND U18636 ( .A(n12694), .B(y[1050]), .Z(n12695) );
  NANDN U18637 ( .A(n12696), .B(n12695), .Z(n21929) );
  ANDN U18638 ( .B(n21916), .A(n12697), .Z(n14352) );
  ANDN U18639 ( .B(n21914), .A(n21911), .Z(n14350) );
  NANDN U18640 ( .A(y[1038]), .B(x[1038]), .Z(n12698) );
  NANDN U18641 ( .A(n12699), .B(n12698), .Z(n21906) );
  NAND U18642 ( .A(n12701), .B(n12700), .Z(n21894) );
  NANDN U18643 ( .A(y[1031]), .B(x[1031]), .Z(n12702) );
  NANDN U18644 ( .A(n12703), .B(n12702), .Z(n21891) );
  ANDN U18645 ( .B(n21888), .A(n12704), .Z(n14329) );
  AND U18646 ( .A(n21883), .B(n21886), .Z(n14327) );
  NANDN U18647 ( .A(n12706), .B(n12705), .Z(n21879) );
  ANDN U18648 ( .B(n21872), .A(n12707), .Z(n14317) );
  AND U18649 ( .A(n21871), .B(n12708), .Z(n14315) );
  XOR U18650 ( .A(x[1022]), .B(n12709), .Z(n14313) );
  NANDN U18651 ( .A(n12711), .B(n12710), .Z(n12712) );
  NANDN U18652 ( .A(n12713), .B(n12712), .Z(n21803) );
  OR U18653 ( .A(n12715), .B(n12714), .Z(n21718) );
  ANDN U18654 ( .B(n21696), .A(n12716), .Z(n14214) );
  ANDN U18655 ( .B(n21633), .A(n12717), .Z(n14173) );
  ANDN U18656 ( .B(n21539), .A(n12718), .Z(n14117) );
  NOR U18657 ( .A(n12720), .B(n12719), .Z(n21473) );
  NANDN U18658 ( .A(n12722), .B(n12721), .Z(n12723) );
  NANDN U18659 ( .A(n12724), .B(n12723), .Z(n21400) );
  NANDN U18660 ( .A(n12726), .B(n12725), .Z(n12727) );
  NANDN U18661 ( .A(n12728), .B(n12727), .Z(n21364) );
  OR U18662 ( .A(n12730), .B(n12729), .Z(n21362) );
  AND U18663 ( .A(n12732), .B(n12731), .Z(n13968) );
  XNOR U18664 ( .A(x[766]), .B(y[766]), .Z(n13966) );
  OR U18665 ( .A(n12734), .B(n12733), .Z(n12736) );
  NAND U18666 ( .A(n12736), .B(n12735), .Z(n12737) );
  NANDN U18667 ( .A(n12738), .B(n12737), .Z(n21226) );
  NANDN U18668 ( .A(n12740), .B(n12739), .Z(n12741) );
  NANDN U18669 ( .A(n12742), .B(n12741), .Z(n21154) );
  NANDN U18670 ( .A(n12744), .B(n12743), .Z(n12745) );
  NANDN U18671 ( .A(n12746), .B(n12745), .Z(n21047) );
  XOR U18672 ( .A(n12747), .B(x[603]), .Z(n13764) );
  NAND U18673 ( .A(n12749), .B(n12748), .Z(n12750) );
  NANDN U18674 ( .A(n12751), .B(n12750), .Z(n20889) );
  NANDN U18675 ( .A(n12753), .B(n12752), .Z(n12754) );
  NANDN U18676 ( .A(n12755), .B(n12754), .Z(n20809) );
  ANDN U18677 ( .B(n12757), .A(n12756), .Z(n12758) );
  NANDN U18678 ( .A(n12759), .B(n12758), .Z(n12760) );
  NAND U18679 ( .A(n12760), .B(n20792), .Z(n13669) );
  NANDN U18680 ( .A(n12762), .B(n12761), .Z(n12763) );
  NANDN U18681 ( .A(n12764), .B(n12763), .Z(n20781) );
  NAND U18682 ( .A(n12765), .B(y[376]), .Z(n12767) );
  ANDN U18683 ( .B(n12767), .A(n12766), .Z(n12769) );
  NANDN U18684 ( .A(n12769), .B(n12768), .Z(n12770) );
  NANDN U18685 ( .A(n12771), .B(n12770), .Z(n20500) );
  OR U18686 ( .A(n12773), .B(n12772), .Z(n20400) );
  NANDN U18687 ( .A(n12775), .B(n12774), .Z(n12777) );
  ANDN U18688 ( .B(n12777), .A(n12776), .Z(n13250) );
  NAND U18689 ( .A(n12779), .B(n12778), .Z(n13035) );
  NAND U18690 ( .A(n12780), .B(y[98]), .Z(n12782) );
  ANDN U18691 ( .B(n12782), .A(n12781), .Z(n13033) );
  NANDN U18692 ( .A(y[97]), .B(x[97]), .Z(n12783) );
  AND U18693 ( .A(n12784), .B(n12783), .Z(n13031) );
  XNOR U18694 ( .A(x[97]), .B(y[97]), .Z(n13029) );
  ANDN U18695 ( .B(n12786), .A(n12785), .Z(n12854) );
  OR U18696 ( .A(n12788), .B(n12787), .Z(n12844) );
  NOR U18697 ( .A(n12790), .B(n12789), .Z(n12828) );
  NOR U18698 ( .A(n12792), .B(n12791), .Z(n12814) );
  ANDN U18699 ( .B(n12793), .A(y[0]), .Z(n12794) );
  NAND U18700 ( .A(n12794), .B(x[0]), .Z(n12795) );
  NANDN U18701 ( .A(n12796), .B(n12795), .Z(n12797) );
  NANDN U18702 ( .A(n12798), .B(n12797), .Z(n12801) );
  OR U18703 ( .A(n12801), .B(y[3]), .Z(n12799) );
  AND U18704 ( .A(n12800), .B(n12799), .Z(n12804) );
  XOR U18705 ( .A(n12801), .B(y[3]), .Z(n12802) );
  NAND U18706 ( .A(n12802), .B(x[3]), .Z(n12803) );
  NAND U18707 ( .A(n12804), .B(n12803), .Z(n12805) );
  NANDN U18708 ( .A(n12806), .B(n12805), .Z(n12807) );
  NANDN U18709 ( .A(n12808), .B(n12807), .Z(n12810) );
  ANDN U18710 ( .B(n12810), .A(n12809), .Z(n12811) );
  OR U18711 ( .A(n12812), .B(n12811), .Z(n12813) );
  AND U18712 ( .A(n12814), .B(n12813), .Z(n12816) );
  NOR U18713 ( .A(n12816), .B(n12815), .Z(n12817) );
  NANDN U18714 ( .A(n12818), .B(n12817), .Z(n12820) );
  ANDN U18715 ( .B(n12820), .A(n12819), .Z(n12822) );
  NAND U18716 ( .A(n12822), .B(n12821), .Z(n12824) );
  ANDN U18717 ( .B(n12824), .A(n12823), .Z(n12825) );
  NANDN U18718 ( .A(n12826), .B(n12825), .Z(n12827) );
  NAND U18719 ( .A(n12828), .B(n12827), .Z(n12830) );
  NAND U18720 ( .A(n12830), .B(n12829), .Z(n12831) );
  OR U18721 ( .A(n12832), .B(n12831), .Z(n12834) );
  ANDN U18722 ( .B(n12834), .A(n12833), .Z(n12835) );
  OR U18723 ( .A(n12836), .B(n12835), .Z(n12837) );
  NANDN U18724 ( .A(n12838), .B(n12837), .Z(n12839) );
  NANDN U18725 ( .A(n12840), .B(n12839), .Z(n12841) );
  NAND U18726 ( .A(n12842), .B(n12841), .Z(n12843) );
  NANDN U18727 ( .A(n12844), .B(n12843), .Z(n12846) );
  ANDN U18728 ( .B(n12846), .A(n12845), .Z(n12848) );
  OR U18729 ( .A(n12848), .B(n12847), .Z(n12849) );
  NANDN U18730 ( .A(n12850), .B(n12849), .Z(n12851) );
  NANDN U18731 ( .A(n12852), .B(n12851), .Z(n12853) );
  NAND U18732 ( .A(n12854), .B(n12853), .Z(n12856) );
  NAND U18733 ( .A(n12856), .B(n12855), .Z(n12859) );
  AND U18734 ( .A(x[22]), .B(n12857), .Z(n12858) );
  OR U18735 ( .A(n12859), .B(n12858), .Z(n12863) );
  ANDN U18736 ( .B(n12861), .A(n12860), .Z(n12862) );
  NAND U18737 ( .A(n12863), .B(n12862), .Z(n12865) );
  NAND U18738 ( .A(n12865), .B(n12864), .Z(n12866) );
  NANDN U18739 ( .A(n12867), .B(n12866), .Z(n12868) );
  NANDN U18740 ( .A(n12869), .B(n12868), .Z(n12871) );
  ANDN U18741 ( .B(n12871), .A(n12870), .Z(n12872) );
  OR U18742 ( .A(n12873), .B(n12872), .Z(n12874) );
  NANDN U18743 ( .A(n12875), .B(n12874), .Z(n12876) );
  NANDN U18744 ( .A(n12877), .B(n12876), .Z(n12878) );
  NANDN U18745 ( .A(n12879), .B(n12878), .Z(n12880) );
  NANDN U18746 ( .A(n12881), .B(n12880), .Z(n12883) );
  ANDN U18747 ( .B(n12883), .A(n12882), .Z(n12884) );
  OR U18748 ( .A(n12885), .B(n12884), .Z(n12886) );
  NANDN U18749 ( .A(n12887), .B(n12886), .Z(n12888) );
  NANDN U18750 ( .A(n12889), .B(n12888), .Z(n12890) );
  NANDN U18751 ( .A(n12891), .B(n12890), .Z(n12892) );
  NANDN U18752 ( .A(n12893), .B(n12892), .Z(n12895) );
  ANDN U18753 ( .B(n12895), .A(n12894), .Z(n12896) );
  OR U18754 ( .A(n12897), .B(n12896), .Z(n12898) );
  NANDN U18755 ( .A(n12899), .B(n12898), .Z(n12900) );
  NANDN U18756 ( .A(n12901), .B(n12900), .Z(n12902) );
  NANDN U18757 ( .A(n12903), .B(n12902), .Z(n12904) );
  NANDN U18758 ( .A(n12905), .B(n12904), .Z(n12907) );
  ANDN U18759 ( .B(n12907), .A(n12906), .Z(n12908) );
  OR U18760 ( .A(n12909), .B(n12908), .Z(n12910) );
  NANDN U18761 ( .A(n12911), .B(n12910), .Z(n12912) );
  NANDN U18762 ( .A(n12913), .B(n12912), .Z(n12914) );
  NANDN U18763 ( .A(n12915), .B(n12914), .Z(n12916) );
  NANDN U18764 ( .A(n12917), .B(n12916), .Z(n12919) );
  ANDN U18765 ( .B(n12919), .A(n12918), .Z(n12920) );
  OR U18766 ( .A(n12921), .B(n12920), .Z(n12922) );
  NANDN U18767 ( .A(n12923), .B(n12922), .Z(n12924) );
  NANDN U18768 ( .A(n12925), .B(n12924), .Z(n12926) );
  NANDN U18769 ( .A(n12927), .B(n12926), .Z(n12928) );
  NANDN U18770 ( .A(n12929), .B(n12928), .Z(n12931) );
  ANDN U18771 ( .B(n12931), .A(n12930), .Z(n12934) );
  AND U18772 ( .A(x[56]), .B(n12932), .Z(n12933) );
  OR U18773 ( .A(n12934), .B(n12933), .Z(n12938) );
  ANDN U18774 ( .B(n12936), .A(n12935), .Z(n12937) );
  NAND U18775 ( .A(n12938), .B(n12937), .Z(n12940) );
  NAND U18776 ( .A(n12940), .B(n12939), .Z(n12941) );
  NANDN U18777 ( .A(n12942), .B(n12941), .Z(n12943) );
  NANDN U18778 ( .A(n12944), .B(n12943), .Z(n12946) );
  ANDN U18779 ( .B(n12946), .A(n12945), .Z(n12947) );
  OR U18780 ( .A(n12948), .B(n12947), .Z(n12949) );
  NANDN U18781 ( .A(n12950), .B(n12949), .Z(n12951) );
  NANDN U18782 ( .A(n12952), .B(n12951), .Z(n12953) );
  NANDN U18783 ( .A(n12954), .B(n12953), .Z(n12955) );
  NANDN U18784 ( .A(n12956), .B(n12955), .Z(n12958) );
  ANDN U18785 ( .B(n12958), .A(n12957), .Z(n12960) );
  OR U18786 ( .A(n12960), .B(n12959), .Z(n12961) );
  NANDN U18787 ( .A(n12962), .B(n12961), .Z(n12965) );
  OR U18788 ( .A(n12965), .B(y[68]), .Z(n12963) );
  AND U18789 ( .A(n12964), .B(n12963), .Z(n12968) );
  XOR U18790 ( .A(n12965), .B(y[68]), .Z(n12966) );
  NAND U18791 ( .A(x[68]), .B(n12966), .Z(n12967) );
  NAND U18792 ( .A(n12968), .B(n12967), .Z(n12969) );
  NANDN U18793 ( .A(n12970), .B(n12969), .Z(n12971) );
  NANDN U18794 ( .A(n12972), .B(n12971), .Z(n12974) );
  ANDN U18795 ( .B(n12974), .A(n12973), .Z(n12975) );
  OR U18796 ( .A(n12976), .B(n12975), .Z(n12977) );
  NANDN U18797 ( .A(n12978), .B(n12977), .Z(n12979) );
  NANDN U18798 ( .A(n12980), .B(n12979), .Z(n12981) );
  NANDN U18799 ( .A(n12982), .B(n12981), .Z(n12983) );
  NANDN U18800 ( .A(n12984), .B(n12983), .Z(n12986) );
  ANDN U18801 ( .B(n12986), .A(n12985), .Z(n12987) );
  OR U18802 ( .A(n12988), .B(n12987), .Z(n12989) );
  NANDN U18803 ( .A(n12990), .B(n12989), .Z(n12991) );
  NANDN U18804 ( .A(n12992), .B(n12991), .Z(n12993) );
  NANDN U18805 ( .A(n12994), .B(n12993), .Z(n12995) );
  NANDN U18806 ( .A(n12996), .B(n12995), .Z(n12998) );
  ANDN U18807 ( .B(n12998), .A(n12997), .Z(n12999) );
  OR U18808 ( .A(n13000), .B(n12999), .Z(n13001) );
  NANDN U18809 ( .A(n13002), .B(n13001), .Z(n13003) );
  NANDN U18810 ( .A(n13004), .B(n13003), .Z(n13005) );
  NANDN U18811 ( .A(n13006), .B(n13005), .Z(n13007) );
  NANDN U18812 ( .A(n13008), .B(n13007), .Z(n13010) );
  ANDN U18813 ( .B(n13010), .A(n13009), .Z(n13011) );
  OR U18814 ( .A(n13012), .B(n13011), .Z(n13013) );
  NANDN U18815 ( .A(n13014), .B(n13013), .Z(n13015) );
  NANDN U18816 ( .A(n13016), .B(n13015), .Z(n13017) );
  NANDN U18817 ( .A(n13018), .B(n13017), .Z(n13019) );
  NANDN U18818 ( .A(n13020), .B(n13019), .Z(n13021) );
  NANDN U18819 ( .A(n13022), .B(n13021), .Z(n13024) );
  NANDN U18820 ( .A(n13024), .B(x[96]), .Z(n13027) );
  XOR U18821 ( .A(n13024), .B(n13023), .Z(n13025) );
  NANDN U18822 ( .A(y[96]), .B(n13025), .Z(n13026) );
  NAND U18823 ( .A(n13027), .B(n13026), .Z(n13028) );
  NAND U18824 ( .A(n13029), .B(n13028), .Z(n13030) );
  NAND U18825 ( .A(n13031), .B(n13030), .Z(n13032) );
  NAND U18826 ( .A(n13033), .B(n13032), .Z(n13034) );
  NAND U18827 ( .A(n13035), .B(n13034), .Z(n13037) );
  NANDN U18828 ( .A(n13037), .B(n13036), .Z(n13038) );
  NANDN U18829 ( .A(n13039), .B(n13038), .Z(n13041) );
  NAND U18830 ( .A(n13041), .B(n13040), .Z(n13042) );
  NANDN U18831 ( .A(n13043), .B(n13042), .Z(n13045) );
  NAND U18832 ( .A(n13045), .B(n13044), .Z(n13047) );
  ANDN U18833 ( .B(n13047), .A(n13046), .Z(n13049) );
  NANDN U18834 ( .A(n13049), .B(n13048), .Z(n13050) );
  NANDN U18835 ( .A(n13051), .B(n13050), .Z(n13053) );
  NAND U18836 ( .A(n13053), .B(n13052), .Z(n13054) );
  NANDN U18837 ( .A(n13055), .B(n13054), .Z(n13057) );
  NAND U18838 ( .A(n13057), .B(n13056), .Z(n13059) );
  ANDN U18839 ( .B(n13059), .A(n13058), .Z(n13061) );
  NANDN U18840 ( .A(n13061), .B(n13060), .Z(n13062) );
  NANDN U18841 ( .A(n13063), .B(n13062), .Z(n13065) );
  NAND U18842 ( .A(n13065), .B(n13064), .Z(n13066) );
  NANDN U18843 ( .A(n13067), .B(n13066), .Z(n13069) );
  NAND U18844 ( .A(n13069), .B(n13068), .Z(n13071) );
  ANDN U18845 ( .B(n13071), .A(n13070), .Z(n13073) );
  NANDN U18846 ( .A(n13073), .B(n13072), .Z(n13074) );
  NANDN U18847 ( .A(n13075), .B(n13074), .Z(n13077) );
  NAND U18848 ( .A(n13077), .B(n13076), .Z(n13078) );
  NANDN U18849 ( .A(n13079), .B(n13078), .Z(n13081) );
  NAND U18850 ( .A(n13081), .B(n13080), .Z(n13083) );
  ANDN U18851 ( .B(n13083), .A(n13082), .Z(n13085) );
  NANDN U18852 ( .A(n13085), .B(n13084), .Z(n13086) );
  NANDN U18853 ( .A(n13087), .B(n13086), .Z(n13089) );
  NAND U18854 ( .A(n13089), .B(n13088), .Z(n13090) );
  NANDN U18855 ( .A(n13091), .B(n13090), .Z(n13093) );
  NAND U18856 ( .A(n13093), .B(n13092), .Z(n13095) );
  ANDN U18857 ( .B(n13095), .A(n13094), .Z(n13097) );
  NANDN U18858 ( .A(n13097), .B(n13096), .Z(n13098) );
  NANDN U18859 ( .A(n13099), .B(n13098), .Z(n13101) );
  NAND U18860 ( .A(n13101), .B(n13100), .Z(n13102) );
  NANDN U18861 ( .A(n13103), .B(n13102), .Z(n13105) );
  NAND U18862 ( .A(n13105), .B(n13104), .Z(n13107) );
  ANDN U18863 ( .B(n13107), .A(n13106), .Z(n13109) );
  NANDN U18864 ( .A(n13109), .B(n13108), .Z(n13110) );
  NANDN U18865 ( .A(n13111), .B(n13110), .Z(n13113) );
  NAND U18866 ( .A(n13113), .B(n13112), .Z(n13114) );
  NANDN U18867 ( .A(n13115), .B(n13114), .Z(n13117) );
  NAND U18868 ( .A(n13117), .B(n13116), .Z(n13119) );
  ANDN U18869 ( .B(n13119), .A(n13118), .Z(n13121) );
  NANDN U18870 ( .A(n13121), .B(n13120), .Z(n13122) );
  NANDN U18871 ( .A(n13123), .B(n13122), .Z(n13125) );
  NAND U18872 ( .A(n13125), .B(n13124), .Z(n13126) );
  NANDN U18873 ( .A(n13127), .B(n13126), .Z(n13129) );
  NAND U18874 ( .A(n13129), .B(n13128), .Z(n13131) );
  ANDN U18875 ( .B(n13131), .A(n13130), .Z(n13133) );
  NANDN U18876 ( .A(n13133), .B(n13132), .Z(n13134) );
  NANDN U18877 ( .A(n13135), .B(n13134), .Z(n13137) );
  NAND U18878 ( .A(n13137), .B(n13136), .Z(n13138) );
  NANDN U18879 ( .A(n13139), .B(n13138), .Z(n13141) );
  NAND U18880 ( .A(n13141), .B(n13140), .Z(n13143) );
  ANDN U18881 ( .B(n13143), .A(n13142), .Z(n13145) );
  NANDN U18882 ( .A(n13145), .B(n13144), .Z(n13146) );
  NANDN U18883 ( .A(n13147), .B(n13146), .Z(n13149) );
  NAND U18884 ( .A(n13149), .B(n13148), .Z(n13150) );
  NANDN U18885 ( .A(n13151), .B(n13150), .Z(n13153) );
  NAND U18886 ( .A(n13153), .B(n13152), .Z(n13154) );
  NANDN U18887 ( .A(n13155), .B(n13154), .Z(n13158) );
  OR U18888 ( .A(n13158), .B(y[160]), .Z(n13156) );
  AND U18889 ( .A(n13157), .B(n13156), .Z(n13161) );
  XOR U18890 ( .A(n13158), .B(y[160]), .Z(n13159) );
  NAND U18891 ( .A(n13159), .B(x[160]), .Z(n13160) );
  NAND U18892 ( .A(n13161), .B(n13160), .Z(n13162) );
  NANDN U18893 ( .A(n13163), .B(n13162), .Z(n13165) );
  NAND U18894 ( .A(n13165), .B(n13164), .Z(n13167) );
  ANDN U18895 ( .B(n13167), .A(n13166), .Z(n13169) );
  NANDN U18896 ( .A(n13169), .B(n13168), .Z(n13170) );
  NANDN U18897 ( .A(n13171), .B(n13170), .Z(n13173) );
  NAND U18898 ( .A(n13173), .B(n13172), .Z(n13174) );
  NANDN U18899 ( .A(n13175), .B(n13174), .Z(n13177) );
  NAND U18900 ( .A(n13177), .B(n13176), .Z(n13179) );
  ANDN U18901 ( .B(n13179), .A(n13178), .Z(n13181) );
  NANDN U18902 ( .A(n13181), .B(n13180), .Z(n13182) );
  NANDN U18903 ( .A(n13183), .B(n13182), .Z(n13185) );
  NAND U18904 ( .A(n13185), .B(n13184), .Z(n13186) );
  NANDN U18905 ( .A(n13187), .B(n13186), .Z(n13189) );
  NAND U18906 ( .A(n13189), .B(n13188), .Z(n13191) );
  ANDN U18907 ( .B(n13191), .A(n13190), .Z(n13193) );
  NANDN U18908 ( .A(n13193), .B(n13192), .Z(n13194) );
  NANDN U18909 ( .A(n13195), .B(n13194), .Z(n13197) );
  NAND U18910 ( .A(n13197), .B(n13196), .Z(n13198) );
  NANDN U18911 ( .A(n13199), .B(n13198), .Z(n13201) );
  NAND U18912 ( .A(n13201), .B(n13200), .Z(n13203) );
  ANDN U18913 ( .B(n13203), .A(n13202), .Z(n13205) );
  NANDN U18914 ( .A(n13205), .B(n13204), .Z(n13206) );
  NANDN U18915 ( .A(n13207), .B(n13206), .Z(n13209) );
  NAND U18916 ( .A(n13209), .B(n13208), .Z(n13210) );
  NANDN U18917 ( .A(n13211), .B(n13210), .Z(n13213) );
  NAND U18918 ( .A(n13212), .B(n13213), .Z(n13216) );
  XOR U18919 ( .A(n13213), .B(n13212), .Z(n13214) );
  NAND U18920 ( .A(n13214), .B(y[186]), .Z(n13215) );
  NAND U18921 ( .A(n13216), .B(n13215), .Z(n13218) );
  ANDN U18922 ( .B(n13218), .A(n13217), .Z(n13219) );
  OR U18923 ( .A(n13220), .B(n13219), .Z(n13221) );
  NANDN U18924 ( .A(n13222), .B(n13221), .Z(n13223) );
  NANDN U18925 ( .A(n13224), .B(n13223), .Z(n13225) );
  NANDN U18926 ( .A(n13226), .B(n13225), .Z(n13227) );
  NANDN U18927 ( .A(n13228), .B(n13227), .Z(n13230) );
  ANDN U18928 ( .B(n13230), .A(n13229), .Z(n13231) );
  OR U18929 ( .A(n13232), .B(n13231), .Z(n13233) );
  NANDN U18930 ( .A(n13234), .B(n13233), .Z(n13235) );
  NANDN U18931 ( .A(n13236), .B(n13235), .Z(n13237) );
  NANDN U18932 ( .A(n13238), .B(n13237), .Z(n13239) );
  NANDN U18933 ( .A(n13240), .B(n13239), .Z(n13242) );
  ANDN U18934 ( .B(n13242), .A(n13241), .Z(n13243) );
  OR U18935 ( .A(n13244), .B(n13243), .Z(n13245) );
  NANDN U18936 ( .A(n13246), .B(n13245), .Z(n13247) );
  NANDN U18937 ( .A(n13248), .B(n13247), .Z(n13249) );
  NAND U18938 ( .A(n13250), .B(n13249), .Z(n13251) );
  NANDN U18939 ( .A(n13252), .B(n13251), .Z(n13253) );
  NANDN U18940 ( .A(n13254), .B(n13253), .Z(n13255) );
  NANDN U18941 ( .A(n13256), .B(n13255), .Z(n13258) );
  ANDN U18942 ( .B(n13258), .A(n13257), .Z(n13259) );
  OR U18943 ( .A(n13260), .B(n13259), .Z(n13261) );
  NANDN U18944 ( .A(n13262), .B(n13261), .Z(n13264) );
  ANDN U18945 ( .B(n13264), .A(n13263), .Z(n13265) );
  OR U18946 ( .A(n13265), .B(x[216]), .Z(n13268) );
  XOR U18947 ( .A(n13265), .B(x[216]), .Z(n13266) );
  NAND U18948 ( .A(n13266), .B(y[216]), .Z(n13267) );
  NAND U18949 ( .A(n13268), .B(n13267), .Z(n13270) );
  ANDN U18950 ( .B(n13270), .A(n13269), .Z(n13271) );
  OR U18951 ( .A(n13272), .B(n13271), .Z(n13273) );
  NANDN U18952 ( .A(n13274), .B(n13273), .Z(n13275) );
  NANDN U18953 ( .A(n13276), .B(n13275), .Z(n13277) );
  NANDN U18954 ( .A(n13278), .B(n13277), .Z(n13279) );
  NANDN U18955 ( .A(n13280), .B(n13279), .Z(n13282) );
  ANDN U18956 ( .B(n13282), .A(n13281), .Z(n13284) );
  NAND U18957 ( .A(n13284), .B(n13283), .Z(n13288) );
  ANDN U18958 ( .B(n13286), .A(n13285), .Z(n13287) );
  NAND U18959 ( .A(n13288), .B(n13287), .Z(n13289) );
  NANDN U18960 ( .A(n13290), .B(n13289), .Z(n13292) );
  NANDN U18961 ( .A(n13292), .B(n13291), .Z(n13295) );
  XNOR U18962 ( .A(n13292), .B(n13291), .Z(n13293) );
  NAND U18963 ( .A(n13293), .B(y[226]), .Z(n13294) );
  NAND U18964 ( .A(n13295), .B(n13294), .Z(n13297) );
  ANDN U18965 ( .B(n13297), .A(n13296), .Z(n13299) );
  NANDN U18966 ( .A(n13299), .B(n13298), .Z(n13300) );
  NANDN U18967 ( .A(n13301), .B(n13300), .Z(n13303) );
  NAND U18968 ( .A(n13303), .B(n13302), .Z(n13304) );
  NANDN U18969 ( .A(n13305), .B(n13304), .Z(n13307) );
  NAND U18970 ( .A(n13307), .B(n13306), .Z(n13309) );
  ANDN U18971 ( .B(n13309), .A(n13308), .Z(n13311) );
  NANDN U18972 ( .A(n13311), .B(n13310), .Z(n13312) );
  NANDN U18973 ( .A(n13313), .B(n13312), .Z(n13315) );
  NAND U18974 ( .A(n13315), .B(n13314), .Z(n13316) );
  NANDN U18975 ( .A(n13317), .B(n13316), .Z(n13319) );
  NAND U18976 ( .A(n13319), .B(n13318), .Z(n13321) );
  ANDN U18977 ( .B(n13321), .A(n13320), .Z(n13323) );
  NANDN U18978 ( .A(n13323), .B(n13322), .Z(n13324) );
  NANDN U18979 ( .A(n13325), .B(n13324), .Z(n13327) );
  NAND U18980 ( .A(n13327), .B(n13326), .Z(n13328) );
  NANDN U18981 ( .A(n13329), .B(n13328), .Z(n13331) );
  NAND U18982 ( .A(n13331), .B(n13330), .Z(n13333) );
  ANDN U18983 ( .B(n13333), .A(n13332), .Z(n13335) );
  NANDN U18984 ( .A(n13335), .B(n13334), .Z(n13336) );
  NANDN U18985 ( .A(n13337), .B(n13336), .Z(n13339) );
  NAND U18986 ( .A(n13339), .B(n13338), .Z(n13340) );
  NANDN U18987 ( .A(n13341), .B(n13340), .Z(n13343) );
  NAND U18988 ( .A(n13343), .B(n13342), .Z(n13345) );
  ANDN U18989 ( .B(n13345), .A(n13344), .Z(n13347) );
  NANDN U18990 ( .A(n13347), .B(n13346), .Z(n13348) );
  NANDN U18991 ( .A(n13349), .B(n13348), .Z(n13351) );
  NAND U18992 ( .A(n13351), .B(n13350), .Z(n13352) );
  NANDN U18993 ( .A(n13353), .B(n13352), .Z(n13355) );
  NAND U18994 ( .A(n13355), .B(n13354), .Z(n13357) );
  ANDN U18995 ( .B(n13357), .A(n13356), .Z(n13359) );
  NANDN U18996 ( .A(n13359), .B(n13358), .Z(n13360) );
  NANDN U18997 ( .A(n13361), .B(n13360), .Z(n13363) );
  NAND U18998 ( .A(n13363), .B(n13362), .Z(n13364) );
  NANDN U18999 ( .A(n13365), .B(n13364), .Z(n13367) );
  NAND U19000 ( .A(n13367), .B(n13366), .Z(n13369) );
  ANDN U19001 ( .B(n13369), .A(n13368), .Z(n13371) );
  NANDN U19002 ( .A(n13371), .B(n13370), .Z(n13372) );
  NANDN U19003 ( .A(n13373), .B(n13372), .Z(n13375) );
  NAND U19004 ( .A(n13375), .B(n13374), .Z(n13376) );
  NANDN U19005 ( .A(x[270]), .B(n13376), .Z(n13379) );
  XNOR U19006 ( .A(n13376), .B(x[270]), .Z(n13377) );
  NAND U19007 ( .A(n13377), .B(y[270]), .Z(n13378) );
  NAND U19008 ( .A(n13379), .B(n13378), .Z(n13381) );
  ANDN U19009 ( .B(n13381), .A(n13380), .Z(n13383) );
  NANDN U19010 ( .A(n13383), .B(n13382), .Z(n13384) );
  NANDN U19011 ( .A(n13385), .B(n13384), .Z(n13387) );
  NAND U19012 ( .A(n13387), .B(n13386), .Z(n13388) );
  NANDN U19013 ( .A(n13389), .B(n13388), .Z(n13391) );
  NAND U19014 ( .A(n13391), .B(n13390), .Z(n13393) );
  ANDN U19015 ( .B(n13393), .A(n13392), .Z(n13395) );
  NANDN U19016 ( .A(n13395), .B(n13394), .Z(n13396) );
  NANDN U19017 ( .A(n13397), .B(n13396), .Z(n13399) );
  NAND U19018 ( .A(n13399), .B(n13398), .Z(n13400) );
  NANDN U19019 ( .A(n13401), .B(n13400), .Z(n13403) );
  NAND U19020 ( .A(n13403), .B(n13402), .Z(n13405) );
  ANDN U19021 ( .B(n13405), .A(n13404), .Z(n13407) );
  NANDN U19022 ( .A(n13407), .B(n13406), .Z(n13409) );
  ANDN U19023 ( .B(n13409), .A(n13408), .Z(n20308) );
  NAND U19024 ( .A(n13410), .B(n20308), .Z(n13411) );
  NAND U19025 ( .A(n13411), .B(n20307), .Z(n13413) );
  ANDN U19026 ( .B(n13413), .A(n13412), .Z(n13414) );
  NANDN U19027 ( .A(n13414), .B(n20313), .Z(n13415) );
  NANDN U19028 ( .A(n13416), .B(n13415), .Z(n13417) );
  NANDN U19029 ( .A(n20317), .B(n13417), .Z(n13418) );
  NAND U19030 ( .A(n13418), .B(n20319), .Z(n13419) );
  NANDN U19031 ( .A(n20322), .B(n13419), .Z(n13420) );
  AND U19032 ( .A(n20323), .B(n13420), .Z(n13421) );
  OR U19033 ( .A(n20326), .B(n13421), .Z(n13422) );
  NAND U19034 ( .A(n13422), .B(n20327), .Z(n13423) );
  NANDN U19035 ( .A(n20329), .B(n13423), .Z(n13424) );
  NAND U19036 ( .A(n13424), .B(n20331), .Z(n13425) );
  NANDN U19037 ( .A(n20334), .B(n13425), .Z(n13426) );
  AND U19038 ( .A(n20335), .B(n13426), .Z(n13427) );
  OR U19039 ( .A(n20338), .B(n13427), .Z(n13428) );
  NAND U19040 ( .A(n13428), .B(n20339), .Z(n13429) );
  NANDN U19041 ( .A(n20341), .B(n13429), .Z(n13430) );
  NAND U19042 ( .A(n13430), .B(n20343), .Z(n13431) );
  NANDN U19043 ( .A(n20346), .B(n13431), .Z(n13432) );
  AND U19044 ( .A(n20347), .B(n13432), .Z(n13433) );
  OR U19045 ( .A(n20350), .B(n13433), .Z(n13434) );
  NAND U19046 ( .A(n13434), .B(n20351), .Z(n13435) );
  NANDN U19047 ( .A(n20353), .B(n13435), .Z(n13436) );
  NAND U19048 ( .A(n13436), .B(n20355), .Z(n13438) );
  NAND U19049 ( .A(n13438), .B(n13437), .Z(n13440) );
  ANDN U19050 ( .B(n13440), .A(n13439), .Z(n13441) );
  NANDN U19051 ( .A(n13441), .B(n20365), .Z(n13442) );
  NAND U19052 ( .A(n13442), .B(n20367), .Z(n13443) );
  NAND U19053 ( .A(n13443), .B(n20370), .Z(n13444) );
  NAND U19054 ( .A(n13444), .B(n20371), .Z(n13445) );
  NAND U19055 ( .A(n13445), .B(n20373), .Z(n13446) );
  AND U19056 ( .A(n20375), .B(n13446), .Z(n13447) );
  NANDN U19057 ( .A(n13447), .B(n20377), .Z(n13448) );
  NAND U19058 ( .A(n13448), .B(n20379), .Z(n13449) );
  NAND U19059 ( .A(n13449), .B(n20383), .Z(n13450) );
  NANDN U19060 ( .A(n20386), .B(n13450), .Z(n13451) );
  NANDN U19061 ( .A(n13452), .B(n13451), .Z(n13453) );
  ANDN U19062 ( .B(n13453), .A(n20390), .Z(n13454) );
  NANDN U19063 ( .A(n13454), .B(n20391), .Z(n13455) );
  NANDN U19064 ( .A(n13456), .B(n13455), .Z(n13457) );
  NAND U19065 ( .A(n13457), .B(n20395), .Z(n13458) );
  NAND U19066 ( .A(n13458), .B(n20306), .Z(n13459) );
  NANDN U19067 ( .A(n20400), .B(n13459), .Z(n13460) );
  AND U19068 ( .A(n20304), .B(n13460), .Z(n13461) );
  OR U19069 ( .A(n13461), .B(n20404), .Z(n13462) );
  NANDN U19070 ( .A(n13463), .B(n13462), .Z(n13464) );
  NAND U19071 ( .A(n13464), .B(n20407), .Z(n13465) );
  NAND U19072 ( .A(n13465), .B(n20409), .Z(n13466) );
  NAND U19073 ( .A(n13466), .B(n20411), .Z(n13467) );
  AND U19074 ( .A(n20414), .B(n13467), .Z(n13468) );
  NANDN U19075 ( .A(n13468), .B(n20415), .Z(n13469) );
  NAND U19076 ( .A(n13469), .B(n20417), .Z(n13470) );
  NAND U19077 ( .A(n13470), .B(n20419), .Z(n13471) );
  NAND U19078 ( .A(n13471), .B(n20421), .Z(n13472) );
  NAND U19079 ( .A(n13472), .B(n20423), .Z(n13473) );
  AND U19080 ( .A(n20426), .B(n13473), .Z(n13474) );
  NANDN U19081 ( .A(n13474), .B(n20427), .Z(n13475) );
  NAND U19082 ( .A(n13475), .B(n20429), .Z(n13476) );
  NAND U19083 ( .A(n13476), .B(n20431), .Z(n13477) );
  NAND U19084 ( .A(n13477), .B(n20433), .Z(n13478) );
  NAND U19085 ( .A(n13478), .B(n20435), .Z(n13479) );
  AND U19086 ( .A(n20438), .B(n13479), .Z(n13480) );
  NANDN U19087 ( .A(n13480), .B(n20439), .Z(n13481) );
  NAND U19088 ( .A(n13481), .B(n20441), .Z(n13482) );
  NAND U19089 ( .A(n13482), .B(n20443), .Z(n13483) );
  NAND U19090 ( .A(n13483), .B(n20445), .Z(n13484) );
  NAND U19091 ( .A(n13484), .B(n20447), .Z(n13485) );
  AND U19092 ( .A(n20450), .B(n13485), .Z(n13490) );
  NANDN U19093 ( .A(n13487), .B(n13486), .Z(n13488) );
  NANDN U19094 ( .A(n13489), .B(n13488), .Z(n20452) );
  OR U19095 ( .A(n13490), .B(n20452), .Z(n13491) );
  NAND U19096 ( .A(n13491), .B(n20453), .Z(n13492) );
  NAND U19097 ( .A(n13492), .B(n20455), .Z(n13493) );
  NAND U19098 ( .A(n13493), .B(n20457), .Z(n13494) );
  NAND U19099 ( .A(n13494), .B(n20459), .Z(n13495) );
  AND U19100 ( .A(n20462), .B(n13495), .Z(n13496) );
  NANDN U19101 ( .A(n13496), .B(n20463), .Z(n13497) );
  NAND U19102 ( .A(n13497), .B(n20466), .Z(n13498) );
  NAND U19103 ( .A(n13498), .B(n20467), .Z(n13499) );
  NAND U19104 ( .A(n13499), .B(n20469), .Z(n13500) );
  NANDN U19105 ( .A(n13501), .B(n13500), .Z(n13503) );
  ANDN U19106 ( .B(n13503), .A(n13502), .Z(n13504) );
  NANDN U19107 ( .A(n13504), .B(n20479), .Z(n13505) );
  NAND U19108 ( .A(n13505), .B(n20481), .Z(n13506) );
  NAND U19109 ( .A(n13506), .B(n20483), .Z(n13507) );
  NANDN U19110 ( .A(n20486), .B(n13507), .Z(n13508) );
  NAND U19111 ( .A(n13508), .B(n20487), .Z(n13509) );
  AND U19112 ( .A(n20490), .B(n13509), .Z(n13510) );
  NANDN U19113 ( .A(n13510), .B(n20491), .Z(n13511) );
  NAND U19114 ( .A(n13511), .B(n20493), .Z(n13512) );
  NAND U19115 ( .A(n13512), .B(n20495), .Z(n13513) );
  NANDN U19116 ( .A(n20498), .B(n13513), .Z(n13514) );
  NANDN U19117 ( .A(n20500), .B(n13514), .Z(n13515) );
  AND U19118 ( .A(n20502), .B(n13515), .Z(n13516) );
  NANDN U19119 ( .A(n13516), .B(n20503), .Z(n13517) );
  NAND U19120 ( .A(n13517), .B(n20505), .Z(n13518) );
  NAND U19121 ( .A(n13518), .B(n20507), .Z(n13519) );
  NAND U19122 ( .A(n13519), .B(n20509), .Z(n13520) );
  NAND U19123 ( .A(n13520), .B(n20511), .Z(n13521) );
  AND U19124 ( .A(n20514), .B(n13521), .Z(n13522) );
  NANDN U19125 ( .A(n13522), .B(n20515), .Z(n13523) );
  NAND U19126 ( .A(n13523), .B(n20517), .Z(n13524) );
  NAND U19127 ( .A(n13524), .B(n20519), .Z(n13525) );
  NAND U19128 ( .A(n13525), .B(n20521), .Z(n13526) );
  NAND U19129 ( .A(n13526), .B(n20523), .Z(n13527) );
  AND U19130 ( .A(n20526), .B(n13527), .Z(n13528) );
  NANDN U19131 ( .A(n13528), .B(n20527), .Z(n13529) );
  NAND U19132 ( .A(n13529), .B(n20529), .Z(n13530) );
  NAND U19133 ( .A(n13530), .B(n20531), .Z(n13531) );
  NAND U19134 ( .A(n13531), .B(n20533), .Z(n13532) );
  NAND U19135 ( .A(n13532), .B(n20535), .Z(n13533) );
  AND U19136 ( .A(n20538), .B(n13533), .Z(n13534) );
  NANDN U19137 ( .A(n13534), .B(n20539), .Z(n13535) );
  NAND U19138 ( .A(n13535), .B(n20541), .Z(n13536) );
  NAND U19139 ( .A(n13536), .B(n20543), .Z(n13537) );
  NAND U19140 ( .A(n13537), .B(n20545), .Z(n13538) );
  NAND U19141 ( .A(n13538), .B(n20547), .Z(n13539) );
  AND U19142 ( .A(n20550), .B(n13539), .Z(n13540) );
  NANDN U19143 ( .A(n13540), .B(n20551), .Z(n13541) );
  NAND U19144 ( .A(n13541), .B(n20553), .Z(n13542) );
  NAND U19145 ( .A(n13542), .B(n20555), .Z(n13543) );
  NAND U19146 ( .A(n13543), .B(n20557), .Z(n13544) );
  NAND U19147 ( .A(n13544), .B(n20559), .Z(n13545) );
  AND U19148 ( .A(n20562), .B(n13545), .Z(n13546) );
  NANDN U19149 ( .A(n13546), .B(n20563), .Z(n13547) );
  NAND U19150 ( .A(n13547), .B(n20565), .Z(n13548) );
  NAND U19151 ( .A(n13548), .B(n20567), .Z(n13549) );
  NAND U19152 ( .A(n13549), .B(n20569), .Z(n13550) );
  NAND U19153 ( .A(n13550), .B(n20571), .Z(n13551) );
  AND U19154 ( .A(n20574), .B(n13551), .Z(n13552) );
  NANDN U19155 ( .A(n13552), .B(n20575), .Z(n13553) );
  NAND U19156 ( .A(n13553), .B(n20577), .Z(n13554) );
  NAND U19157 ( .A(n13554), .B(n20579), .Z(n13555) );
  NAND U19158 ( .A(n13555), .B(n20581), .Z(n13556) );
  NAND U19159 ( .A(n13556), .B(n20583), .Z(n13557) );
  AND U19160 ( .A(n20586), .B(n13557), .Z(n13558) );
  NANDN U19161 ( .A(n13558), .B(n20587), .Z(n13559) );
  NAND U19162 ( .A(n13559), .B(n20590), .Z(n13560) );
  NAND U19163 ( .A(n13560), .B(n20591), .Z(n13561) );
  NAND U19164 ( .A(n13561), .B(n20593), .Z(n13562) );
  NANDN U19165 ( .A(n13563), .B(n13562), .Z(n13565) );
  ANDN U19166 ( .B(n13565), .A(n13564), .Z(n13566) );
  NANDN U19167 ( .A(n13566), .B(n20603), .Z(n13567) );
  NAND U19168 ( .A(n13567), .B(n20605), .Z(n13568) );
  NAND U19169 ( .A(n13568), .B(n20607), .Z(n13569) );
  NAND U19170 ( .A(n13569), .B(n20609), .Z(n13570) );
  NAND U19171 ( .A(n13570), .B(n20611), .Z(n13571) );
  AND U19172 ( .A(n20614), .B(n13571), .Z(n13572) );
  NANDN U19173 ( .A(n13572), .B(n20615), .Z(n13573) );
  NAND U19174 ( .A(n13573), .B(n20617), .Z(n13575) );
  NAND U19175 ( .A(n13575), .B(n13574), .Z(n13576) );
  NANDN U19176 ( .A(n13577), .B(n13576), .Z(n13578) );
  NAND U19177 ( .A(n13578), .B(n20628), .Z(n13579) );
  AND U19178 ( .A(n20630), .B(n13579), .Z(n13580) );
  NANDN U19179 ( .A(n13580), .B(n20632), .Z(n13581) );
  NAND U19180 ( .A(n13581), .B(n20634), .Z(n13582) );
  NAND U19181 ( .A(n13582), .B(n20636), .Z(n13583) );
  NAND U19182 ( .A(n13583), .B(n20639), .Z(n13584) );
  NAND U19183 ( .A(n13584), .B(n20640), .Z(n13585) );
  AND U19184 ( .A(n20642), .B(n13585), .Z(n13586) );
  NANDN U19185 ( .A(n13586), .B(n20644), .Z(n13587) );
  NAND U19186 ( .A(n13587), .B(n20646), .Z(n13588) );
  NAND U19187 ( .A(n13588), .B(n20648), .Z(n13589) );
  NAND U19188 ( .A(n13589), .B(n20651), .Z(n13590) );
  NAND U19189 ( .A(n13590), .B(n20652), .Z(n13591) );
  AND U19190 ( .A(n20654), .B(n13591), .Z(n13592) );
  NANDN U19191 ( .A(n13592), .B(n20656), .Z(n13593) );
  NANDN U19192 ( .A(n20659), .B(n13593), .Z(n13594) );
  NAND U19193 ( .A(n13594), .B(n20660), .Z(n13595) );
  NAND U19194 ( .A(n13595), .B(n20663), .Z(n13596) );
  NAND U19195 ( .A(n13596), .B(n20664), .Z(n13597) );
  AND U19196 ( .A(n20666), .B(n13597), .Z(n13598) );
  NANDN U19197 ( .A(n13598), .B(n20668), .Z(n13599) );
  NAND U19198 ( .A(n13599), .B(n20670), .Z(n13600) );
  NAND U19199 ( .A(n13600), .B(n20672), .Z(n13601) );
  NAND U19200 ( .A(n13601), .B(n20675), .Z(n13602) );
  NAND U19201 ( .A(n13602), .B(n20676), .Z(n13603) );
  AND U19202 ( .A(n20678), .B(n13603), .Z(n13604) );
  NANDN U19203 ( .A(n13604), .B(n20680), .Z(n13605) );
  NAND U19204 ( .A(n13605), .B(n20682), .Z(n13606) );
  NAND U19205 ( .A(n13606), .B(n20684), .Z(n13607) );
  NAND U19206 ( .A(n13607), .B(n20687), .Z(n13608) );
  NAND U19207 ( .A(n13608), .B(n20688), .Z(n13609) );
  AND U19208 ( .A(n20690), .B(n13609), .Z(n13610) );
  NANDN U19209 ( .A(n13610), .B(n20692), .Z(n13611) );
  NAND U19210 ( .A(n13611), .B(n20694), .Z(n13612) );
  NAND U19211 ( .A(n13612), .B(n20696), .Z(n13613) );
  NAND U19212 ( .A(n13613), .B(n20699), .Z(n13614) );
  NAND U19213 ( .A(n13614), .B(n20700), .Z(n13615) );
  AND U19214 ( .A(n20702), .B(n13615), .Z(n13616) );
  NANDN U19215 ( .A(n13616), .B(n20704), .Z(n13617) );
  NAND U19216 ( .A(n13617), .B(n20706), .Z(n13618) );
  NAND U19217 ( .A(n13618), .B(n20708), .Z(n13619) );
  NAND U19218 ( .A(n13619), .B(n20711), .Z(n13620) );
  NAND U19219 ( .A(n13620), .B(n20712), .Z(n13621) );
  ANDN U19220 ( .B(n13621), .A(n20715), .Z(n13629) );
  NAND U19221 ( .A(n13622), .B(y[482]), .Z(n13624) );
  ANDN U19222 ( .B(n13624), .A(n13623), .Z(n13626) );
  NANDN U19223 ( .A(n13626), .B(n13625), .Z(n13627) );
  NANDN U19224 ( .A(n13628), .B(n13627), .Z(n20717) );
  OR U19225 ( .A(n13629), .B(n20717), .Z(n13630) );
  NANDN U19226 ( .A(n20719), .B(n13630), .Z(n13631) );
  NAND U19227 ( .A(n13631), .B(n20720), .Z(n13632) );
  NANDN U19228 ( .A(n20722), .B(n13632), .Z(n13633) );
  NAND U19229 ( .A(n13633), .B(n20724), .Z(n13634) );
  ANDN U19230 ( .B(n13634), .A(n20727), .Z(n13635) );
  NANDN U19231 ( .A(n13635), .B(n20728), .Z(n13636) );
  NANDN U19232 ( .A(n20731), .B(n13636), .Z(n13637) );
  NAND U19233 ( .A(n13637), .B(n20732), .Z(n13638) );
  NANDN U19234 ( .A(n20734), .B(n13638), .Z(n13639) );
  NAND U19235 ( .A(n13639), .B(n20736), .Z(n13640) );
  ANDN U19236 ( .B(n13640), .A(n20739), .Z(n13641) );
  NANDN U19237 ( .A(n13641), .B(n20740), .Z(n13642) );
  NANDN U19238 ( .A(n20743), .B(n13642), .Z(n13643) );
  NAND U19239 ( .A(n13643), .B(n20744), .Z(n13644) );
  NANDN U19240 ( .A(n20746), .B(n13644), .Z(n13645) );
  NAND U19241 ( .A(n13645), .B(n20748), .Z(n13646) );
  ANDN U19242 ( .B(n13646), .A(n20751), .Z(n13647) );
  NANDN U19243 ( .A(n13647), .B(n20752), .Z(n13648) );
  NANDN U19244 ( .A(n20755), .B(n13648), .Z(n13649) );
  NAND U19245 ( .A(n13649), .B(n20756), .Z(n13650) );
  NANDN U19246 ( .A(n20758), .B(n13650), .Z(n13651) );
  NAND U19247 ( .A(n13651), .B(n20760), .Z(n13652) );
  ANDN U19248 ( .B(n13652), .A(n20763), .Z(n13653) );
  NANDN U19249 ( .A(n13653), .B(n20764), .Z(n13654) );
  NANDN U19250 ( .A(n20767), .B(n13654), .Z(n13655) );
  NAND U19251 ( .A(n13655), .B(n20768), .Z(n13656) );
  NANDN U19252 ( .A(n20770), .B(n13656), .Z(n13657) );
  NAND U19253 ( .A(n13657), .B(n20772), .Z(n13658) );
  ANDN U19254 ( .B(n13658), .A(n20775), .Z(n13659) );
  NANDN U19255 ( .A(n13659), .B(n20776), .Z(n13660) );
  NAND U19256 ( .A(n13660), .B(n20778), .Z(n13661) );
  NANDN U19257 ( .A(n20781), .B(n13661), .Z(n13662) );
  NANDN U19258 ( .A(n20782), .B(n13662), .Z(n13663) );
  NAND U19259 ( .A(n13663), .B(n20784), .Z(n13664) );
  ANDN U19260 ( .B(n13664), .A(n20787), .Z(n13665) );
  OR U19261 ( .A(n13666), .B(n13665), .Z(n13667) );
  NANDN U19262 ( .A(n20791), .B(n13667), .Z(n13668) );
  NANDN U19263 ( .A(n13669), .B(n13668), .Z(n13670) );
  NANDN U19264 ( .A(n20794), .B(n13670), .Z(n13671) );
  NAND U19265 ( .A(n13671), .B(n20796), .Z(n13672) );
  ANDN U19266 ( .B(n13672), .A(n20799), .Z(n13673) );
  NANDN U19267 ( .A(n13673), .B(n20800), .Z(n13674) );
  NANDN U19268 ( .A(n20803), .B(n13674), .Z(n13675) );
  NAND U19269 ( .A(n13675), .B(n20804), .Z(n13676) );
  NAND U19270 ( .A(n13676), .B(n20807), .Z(n13677) );
  NANDN U19271 ( .A(n20809), .B(n13677), .Z(n13678) );
  ANDN U19272 ( .B(n13678), .A(n20811), .Z(n13679) );
  NANDN U19273 ( .A(n13679), .B(n20812), .Z(n13680) );
  NANDN U19274 ( .A(n20815), .B(n13680), .Z(n13681) );
  NAND U19275 ( .A(n13681), .B(n20816), .Z(n13682) );
  NANDN U19276 ( .A(n20818), .B(n13682), .Z(n13683) );
  NAND U19277 ( .A(n13683), .B(n20820), .Z(n13684) );
  ANDN U19278 ( .B(n13684), .A(n20823), .Z(n13685) );
  NANDN U19279 ( .A(n13685), .B(n20824), .Z(n13686) );
  NANDN U19280 ( .A(n20827), .B(n13686), .Z(n13687) );
  NAND U19281 ( .A(n13687), .B(n20828), .Z(n13688) );
  NANDN U19282 ( .A(n20830), .B(n13688), .Z(n13689) );
  NAND U19283 ( .A(n13689), .B(n20832), .Z(n13690) );
  ANDN U19284 ( .B(n13690), .A(n20835), .Z(n13691) );
  NANDN U19285 ( .A(n13691), .B(n20836), .Z(n13692) );
  NANDN U19286 ( .A(n20839), .B(n13692), .Z(n13693) );
  NAND U19287 ( .A(n13693), .B(n20840), .Z(n13694) );
  NANDN U19288 ( .A(n20842), .B(n13694), .Z(n13695) );
  NAND U19289 ( .A(n13695), .B(n20844), .Z(n13696) );
  ANDN U19290 ( .B(n13696), .A(n20847), .Z(n13697) );
  NANDN U19291 ( .A(n13697), .B(n20848), .Z(n13698) );
  NANDN U19292 ( .A(n20851), .B(n13698), .Z(n13699) );
  NAND U19293 ( .A(n13699), .B(n20852), .Z(n13700) );
  NANDN U19294 ( .A(n20854), .B(n13700), .Z(n13701) );
  NAND U19295 ( .A(n13701), .B(n20856), .Z(n13702) );
  ANDN U19296 ( .B(n13702), .A(n20859), .Z(n13704) );
  NANDN U19297 ( .A(n13704), .B(n13703), .Z(n13706) );
  NAND U19298 ( .A(n13706), .B(n13705), .Z(n13707) );
  NAND U19299 ( .A(n13707), .B(n20864), .Z(n13711) );
  NANDN U19300 ( .A(n13709), .B(n13708), .Z(n13710) );
  NANDN U19301 ( .A(n13711), .B(n13710), .Z(n13712) );
  ANDN U19302 ( .B(n13712), .A(n20866), .Z(n13713) );
  NANDN U19303 ( .A(n13713), .B(n20868), .Z(n13714) );
  NANDN U19304 ( .A(n20871), .B(n13714), .Z(n13715) );
  NAND U19305 ( .A(n13715), .B(n20872), .Z(n13716) );
  NANDN U19306 ( .A(n20875), .B(n13716), .Z(n13717) );
  NANDN U19307 ( .A(n13718), .B(n13717), .Z(n13719) );
  AND U19308 ( .A(n20879), .B(n13719), .Z(n13720) );
  NANDN U19309 ( .A(n13720), .B(n20880), .Z(n13721) );
  NANDN U19310 ( .A(n20887), .B(n13721), .Z(n13722) );
  NANDN U19311 ( .A(n20889), .B(n13722), .Z(n13723) );
  NAND U19312 ( .A(n13723), .B(n20891), .Z(n13724) );
  NAND U19313 ( .A(n13724), .B(n20892), .Z(n13725) );
  AND U19314 ( .A(n20894), .B(n13725), .Z(n13726) );
  NANDN U19315 ( .A(n13726), .B(n20896), .Z(n13727) );
  NAND U19316 ( .A(n13727), .B(n20898), .Z(n13728) );
  NAND U19317 ( .A(n13728), .B(n20900), .Z(n13729) );
  NAND U19318 ( .A(n13729), .B(n20903), .Z(n13730) );
  NANDN U19319 ( .A(n20905), .B(n13730), .Z(n13731) );
  AND U19320 ( .A(n20906), .B(n13731), .Z(n13732) );
  OR U19321 ( .A(n20908), .B(n13732), .Z(n13733) );
  NAND U19322 ( .A(n13733), .B(n20910), .Z(n13734) );
  NAND U19323 ( .A(n13734), .B(n20912), .Z(n13735) );
  NAND U19324 ( .A(n13735), .B(n20914), .Z(n13736) );
  NANDN U19325 ( .A(n20917), .B(n13736), .Z(n13737) );
  AND U19326 ( .A(n20918), .B(n13737), .Z(n13738) );
  OR U19327 ( .A(n13738), .B(n20920), .Z(n13739) );
  AND U19328 ( .A(n20922), .B(n13739), .Z(n13740) );
  OR U19329 ( .A(n20925), .B(n13740), .Z(n13741) );
  NAND U19330 ( .A(n13741), .B(n20926), .Z(n13743) );
  NAND U19331 ( .A(n13743), .B(n13742), .Z(n13744) );
  NAND U19332 ( .A(n13745), .B(n13744), .Z(n13746) );
  NANDN U19333 ( .A(n13747), .B(n13746), .Z(n13749) );
  ANDN U19334 ( .B(n13749), .A(n13748), .Z(n13750) );
  NANDN U19335 ( .A(n13750), .B(n20933), .Z(n13751) );
  NAND U19336 ( .A(n13751), .B(n20934), .Z(n13752) );
  ANDN U19337 ( .B(n13752), .A(n20937), .Z(n13753) );
  NANDN U19338 ( .A(n13753), .B(n20938), .Z(n13754) );
  NANDN U19339 ( .A(n20941), .B(n13754), .Z(n13755) );
  NAND U19340 ( .A(n13755), .B(n20942), .Z(n13756) );
  NANDN U19341 ( .A(n20944), .B(n13756), .Z(n13757) );
  NAND U19342 ( .A(n13757), .B(n20946), .Z(n13758) );
  ANDN U19343 ( .B(n13758), .A(n20949), .Z(n13759) );
  NANDN U19344 ( .A(n13759), .B(n20950), .Z(n13760) );
  NANDN U19345 ( .A(n20953), .B(n13760), .Z(n13762) );
  NAND U19346 ( .A(n13762), .B(n13761), .Z(n13763) );
  NAND U19347 ( .A(n13764), .B(n13763), .Z(n13765) );
  AND U19348 ( .A(n13766), .B(n13765), .Z(n13769) );
  OR U19349 ( .A(n13769), .B(y[604]), .Z(n13767) );
  AND U19350 ( .A(n13768), .B(n13767), .Z(n13772) );
  XOR U19351 ( .A(y[604]), .B(n13769), .Z(n13770) );
  NAND U19352 ( .A(n13770), .B(x[604]), .Z(n13771) );
  NAND U19353 ( .A(n13772), .B(n13771), .Z(n13773) );
  NANDN U19354 ( .A(n20961), .B(n13773), .Z(n13774) );
  NAND U19355 ( .A(n13774), .B(n20962), .Z(n13775) );
  ANDN U19356 ( .B(n13775), .A(n20965), .Z(n13776) );
  NANDN U19357 ( .A(n13776), .B(n20966), .Z(n13777) );
  NANDN U19358 ( .A(n20968), .B(n13777), .Z(n13778) );
  NAND U19359 ( .A(n13778), .B(n20970), .Z(n13779) );
  NANDN U19360 ( .A(n20973), .B(n13779), .Z(n13780) );
  NAND U19361 ( .A(n13780), .B(n20974), .Z(n13781) );
  ANDN U19362 ( .B(n13781), .A(n20977), .Z(n13782) );
  NANDN U19363 ( .A(n13782), .B(n20978), .Z(n13783) );
  NANDN U19364 ( .A(n20980), .B(n13783), .Z(n13784) );
  NAND U19365 ( .A(n13784), .B(n20982), .Z(n13785) );
  NANDN U19366 ( .A(n20985), .B(n13785), .Z(n13786) );
  NAND U19367 ( .A(n13786), .B(n20986), .Z(n13787) );
  ANDN U19368 ( .B(n13787), .A(n20989), .Z(n13788) );
  NANDN U19369 ( .A(n13788), .B(n20990), .Z(n13789) );
  NANDN U19370 ( .A(n20992), .B(n13789), .Z(n13790) );
  NAND U19371 ( .A(n13790), .B(n20994), .Z(n13791) );
  NANDN U19372 ( .A(n20997), .B(n13791), .Z(n13792) );
  NAND U19373 ( .A(n13792), .B(n20998), .Z(n13793) );
  AND U19374 ( .A(n21000), .B(n13793), .Z(n13794) );
  NANDN U19375 ( .A(n13794), .B(n21002), .Z(n13795) );
  NANDN U19376 ( .A(n21004), .B(n13795), .Z(n13796) );
  NAND U19377 ( .A(n13796), .B(n21006), .Z(n13797) );
  NANDN U19378 ( .A(n21009), .B(n13797), .Z(n13798) );
  NAND U19379 ( .A(n13798), .B(n21010), .Z(n13799) );
  AND U19380 ( .A(n13800), .B(n13799), .Z(n13803) );
  AND U19381 ( .A(x[632]), .B(n13801), .Z(n13802) );
  OR U19382 ( .A(n13803), .B(n13802), .Z(n13804) );
  NANDN U19383 ( .A(n13805), .B(n13804), .Z(n13807) );
  NAND U19384 ( .A(n13807), .B(n13806), .Z(n13808) );
  NANDN U19385 ( .A(n21019), .B(n13808), .Z(n13809) );
  NANDN U19386 ( .A(n13810), .B(n13809), .Z(n13811) );
  NAND U19387 ( .A(n13811), .B(n21023), .Z(n13812) );
  NAND U19388 ( .A(n13812), .B(n21024), .Z(n13813) );
  NANDN U19389 ( .A(n21027), .B(n13813), .Z(n13814) );
  AND U19390 ( .A(n21028), .B(n13814), .Z(n13815) );
  OR U19391 ( .A(n21031), .B(n13815), .Z(n13816) );
  NAND U19392 ( .A(n13816), .B(n21032), .Z(n13817) );
  NANDN U19393 ( .A(n21034), .B(n13817), .Z(n13818) );
  NAND U19394 ( .A(n13818), .B(n21036), .Z(n13819) );
  NAND U19395 ( .A(n13819), .B(n21039), .Z(n13820) );
  AND U19396 ( .A(n21040), .B(n13820), .Z(n13825) );
  NANDN U19397 ( .A(n13822), .B(n13821), .Z(n13823) );
  NANDN U19398 ( .A(n13824), .B(n13823), .Z(n21043) );
  OR U19399 ( .A(n13825), .B(n21043), .Z(n13826) );
  NAND U19400 ( .A(n13826), .B(n21044), .Z(n13827) );
  NANDN U19401 ( .A(n21047), .B(n13827), .Z(n13828) );
  NANDN U19402 ( .A(n21049), .B(n13828), .Z(n13829) );
  NAND U19403 ( .A(n13829), .B(n21050), .Z(n13830) );
  ANDN U19404 ( .B(n13830), .A(n21053), .Z(n13831) );
  NANDN U19405 ( .A(n13831), .B(n21054), .Z(n13832) );
  NANDN U19406 ( .A(n21056), .B(n13832), .Z(n13833) );
  NAND U19407 ( .A(n13833), .B(n21058), .Z(n13834) );
  NANDN U19408 ( .A(n21061), .B(n13834), .Z(n13835) );
  NAND U19409 ( .A(n13835), .B(n21062), .Z(n13836) );
  ANDN U19410 ( .B(n13836), .A(n21065), .Z(n13837) );
  NANDN U19411 ( .A(n13837), .B(n21066), .Z(n13838) );
  NANDN U19412 ( .A(n21068), .B(n13838), .Z(n13839) );
  NAND U19413 ( .A(n13839), .B(n21070), .Z(n13840) );
  NANDN U19414 ( .A(n21073), .B(n13840), .Z(n13841) );
  NAND U19415 ( .A(n13841), .B(n21074), .Z(n13842) );
  AND U19416 ( .A(n21076), .B(n13842), .Z(n13847) );
  NANDN U19417 ( .A(n13844), .B(n13843), .Z(n13845) );
  NANDN U19418 ( .A(n13846), .B(n13845), .Z(n21079) );
  OR U19419 ( .A(n13847), .B(n21079), .Z(n13848) );
  NANDN U19420 ( .A(n21080), .B(n13848), .Z(n13849) );
  NAND U19421 ( .A(n13849), .B(n21082), .Z(n13850) );
  NANDN U19422 ( .A(n21085), .B(n13850), .Z(n13851) );
  NAND U19423 ( .A(n13851), .B(n21086), .Z(n13852) );
  ANDN U19424 ( .B(n13852), .A(n21089), .Z(n13853) );
  NANDN U19425 ( .A(n13853), .B(n21090), .Z(n13854) );
  NANDN U19426 ( .A(n21092), .B(n13854), .Z(n13856) );
  NAND U19427 ( .A(n13856), .B(n13855), .Z(n13857) );
  NANDN U19428 ( .A(n13857), .B(n21094), .Z(n13859) );
  AND U19429 ( .A(n21096), .B(n21101), .Z(n13858) );
  NAND U19430 ( .A(n13859), .B(n13858), .Z(n13860) );
  NAND U19431 ( .A(n13860), .B(n21104), .Z(n13862) );
  NANDN U19432 ( .A(n13862), .B(n13861), .Z(n13863) );
  NANDN U19433 ( .A(n13864), .B(n13863), .Z(n13865) );
  NANDN U19434 ( .A(n13866), .B(n13865), .Z(n13867) );
  NANDN U19435 ( .A(n13868), .B(n13867), .Z(n13869) );
  NAND U19436 ( .A(n13869), .B(n21117), .Z(n13870) );
  AND U19437 ( .A(n21119), .B(n13870), .Z(n13871) );
  NANDN U19438 ( .A(n13871), .B(n21122), .Z(n13872) );
  NAND U19439 ( .A(n13872), .B(n21123), .Z(n13873) );
  NAND U19440 ( .A(n13873), .B(n21125), .Z(n13874) );
  NAND U19441 ( .A(n13874), .B(n21127), .Z(n13875) );
  NAND U19442 ( .A(n13875), .B(n21129), .Z(n13876) );
  AND U19443 ( .A(n21131), .B(n13876), .Z(n13877) );
  NANDN U19444 ( .A(n13877), .B(n21134), .Z(n13878) );
  NAND U19445 ( .A(n13878), .B(n21135), .Z(n13879) );
  NAND U19446 ( .A(n13879), .B(n21137), .Z(n13880) );
  NAND U19447 ( .A(n13880), .B(n21139), .Z(n13881) );
  NAND U19448 ( .A(n13881), .B(n21141), .Z(n13882) );
  AND U19449 ( .A(n21143), .B(n13882), .Z(n13884) );
  NANDN U19450 ( .A(n13884), .B(n13883), .Z(n13885) );
  NAND U19451 ( .A(n13885), .B(n21147), .Z(n13886) );
  NAND U19452 ( .A(n13886), .B(n20299), .Z(n13887) );
  NAND U19453 ( .A(n13887), .B(n21151), .Z(n13888) );
  NANDN U19454 ( .A(n21154), .B(n13888), .Z(n13889) );
  ANDN U19455 ( .B(n13889), .A(n21156), .Z(n13890) );
  NANDN U19456 ( .A(n13890), .B(n21157), .Z(n13891) );
  NANDN U19457 ( .A(n21160), .B(n13891), .Z(n13892) );
  NAND U19458 ( .A(n13892), .B(n21161), .Z(n13893) );
  NANDN U19459 ( .A(n21163), .B(n13893), .Z(n13894) );
  NAND U19460 ( .A(n13894), .B(n21165), .Z(n13895) );
  NANDN U19461 ( .A(n21168), .B(n13895), .Z(n13896) );
  NAND U19462 ( .A(n13896), .B(n21169), .Z(n13897) );
  NANDN U19463 ( .A(n21172), .B(n13897), .Z(n13898) );
  AND U19464 ( .A(n21173), .B(n13898), .Z(n13899) );
  OR U19465 ( .A(n21175), .B(n13899), .Z(n13900) );
  NAND U19466 ( .A(n13900), .B(n21177), .Z(n13901) );
  NANDN U19467 ( .A(n21180), .B(n13901), .Z(n13902) );
  NAND U19468 ( .A(n13902), .B(n21181), .Z(n13903) );
  NAND U19469 ( .A(n13903), .B(n21183), .Z(n13908) );
  NANDN U19470 ( .A(n13905), .B(n13904), .Z(n13906) );
  NANDN U19471 ( .A(n13907), .B(n13906), .Z(n21186) );
  ANDN U19472 ( .B(n13908), .A(n21186), .Z(n13909) );
  OR U19473 ( .A(n13909), .B(n21187), .Z(n13910) );
  NAND U19474 ( .A(n13910), .B(n21189), .Z(n13911) );
  ANDN U19475 ( .B(n13911), .A(n21192), .Z(n13912) );
  NANDN U19476 ( .A(n13912), .B(n21193), .Z(n13913) );
  NANDN U19477 ( .A(n21196), .B(n13913), .Z(n13914) );
  NAND U19478 ( .A(n13914), .B(n21197), .Z(n13915) );
  NANDN U19479 ( .A(n21199), .B(n13915), .Z(n13916) );
  NAND U19480 ( .A(n13916), .B(n21201), .Z(n13917) );
  ANDN U19481 ( .B(n13917), .A(n21204), .Z(n13918) );
  NANDN U19482 ( .A(n13918), .B(n21205), .Z(n13919) );
  NANDN U19483 ( .A(n21208), .B(n13919), .Z(n13920) );
  NAND U19484 ( .A(n13920), .B(n21209), .Z(n13921) );
  NANDN U19485 ( .A(n21211), .B(n13921), .Z(n13922) );
  NAND U19486 ( .A(n13922), .B(n21213), .Z(n13923) );
  ANDN U19487 ( .B(n13923), .A(n21216), .Z(n13924) );
  NANDN U19488 ( .A(n13924), .B(n21217), .Z(n13925) );
  NANDN U19489 ( .A(n21220), .B(n13925), .Z(n13926) );
  NAND U19490 ( .A(n13926), .B(n21221), .Z(n13927) );
  NAND U19491 ( .A(n13927), .B(n21224), .Z(n13928) );
  NANDN U19492 ( .A(n21226), .B(n13928), .Z(n13929) );
  ANDN U19493 ( .B(n13929), .A(n21228), .Z(n13930) );
  NANDN U19494 ( .A(n13930), .B(n21229), .Z(n13931) );
  NANDN U19495 ( .A(n21232), .B(n13931), .Z(n13932) );
  AND U19496 ( .A(n21233), .B(n13932), .Z(n13933) );
  NANDN U19497 ( .A(n13933), .B(n21236), .Z(n13934) );
  NAND U19498 ( .A(n13934), .B(n21237), .Z(n13935) );
  NAND U19499 ( .A(n13935), .B(n21239), .Z(n13936) );
  NAND U19500 ( .A(n13936), .B(n21241), .Z(n13937) );
  NAND U19501 ( .A(n13937), .B(n21243), .Z(n13938) );
  AND U19502 ( .A(n21245), .B(n13938), .Z(n13939) );
  NANDN U19503 ( .A(n13939), .B(n21248), .Z(n13940) );
  NAND U19504 ( .A(n13940), .B(n21249), .Z(n13941) );
  NAND U19505 ( .A(n13941), .B(n21251), .Z(n13942) );
  NANDN U19506 ( .A(n13943), .B(n13942), .Z(n13944) );
  NAND U19507 ( .A(n13945), .B(n13944), .Z(n13947) );
  NAND U19508 ( .A(n13947), .B(n13946), .Z(n13949) );
  ANDN U19509 ( .B(n13949), .A(n13948), .Z(n13950) );
  OR U19510 ( .A(n13950), .B(n21260), .Z(n13952) );
  NAND U19511 ( .A(n13952), .B(n13951), .Z(n13953) );
  AND U19512 ( .A(n21267), .B(n13953), .Z(n13954) );
  NANDN U19513 ( .A(n13954), .B(n21269), .Z(n13955) );
  NAND U19514 ( .A(n13955), .B(n21271), .Z(n13956) );
  NAND U19515 ( .A(n13956), .B(n21273), .Z(n13957) );
  NAND U19516 ( .A(n13957), .B(n21275), .Z(n13958) );
  NAND U19517 ( .A(n13958), .B(n21278), .Z(n13959) );
  AND U19518 ( .A(n21279), .B(n13959), .Z(n13960) );
  NANDN U19519 ( .A(n13960), .B(n21281), .Z(n13961) );
  NAND U19520 ( .A(n13961), .B(n21283), .Z(n13962) );
  NAND U19521 ( .A(n13962), .B(n21285), .Z(n13964) );
  ANDN U19522 ( .B(n13964), .A(n13963), .Z(n13965) );
  NAND U19523 ( .A(n13966), .B(n13965), .Z(n13967) );
  NAND U19524 ( .A(n13968), .B(n13967), .Z(n13969) );
  NAND U19525 ( .A(n13969), .B(n21291), .Z(n13970) );
  NAND U19526 ( .A(n13970), .B(n21293), .Z(n13971) );
  AND U19527 ( .A(n21295), .B(n13971), .Z(n13972) );
  NANDN U19528 ( .A(n13972), .B(n21297), .Z(n13973) );
  NAND U19529 ( .A(n13973), .B(n21299), .Z(n13974) );
  NAND U19530 ( .A(n13974), .B(n21302), .Z(n13975) );
  NAND U19531 ( .A(n13975), .B(n21303), .Z(n13976) );
  NANDN U19532 ( .A(n21305), .B(n13976), .Z(n13984) );
  NAND U19533 ( .A(n13977), .B(y[774]), .Z(n13979) );
  ANDN U19534 ( .B(n13979), .A(n13978), .Z(n13981) );
  NANDN U19535 ( .A(n13981), .B(n13980), .Z(n13982) );
  NANDN U19536 ( .A(n13983), .B(n13982), .Z(n21308) );
  ANDN U19537 ( .B(n13984), .A(n21308), .Z(n13985) );
  NANDN U19538 ( .A(n13985), .B(n21309), .Z(n13986) );
  NAND U19539 ( .A(n13986), .B(n21312), .Z(n13987) );
  NAND U19540 ( .A(n13987), .B(n21313), .Z(n13988) );
  NAND U19541 ( .A(n13988), .B(n21315), .Z(n13989) );
  NAND U19542 ( .A(n13989), .B(n21317), .Z(n13990) );
  AND U19543 ( .A(n21319), .B(n13990), .Z(n13991) );
  NANDN U19544 ( .A(n13991), .B(n21321), .Z(n13992) );
  NAND U19545 ( .A(n13992), .B(n21324), .Z(n13993) );
  NAND U19546 ( .A(n13993), .B(n21325), .Z(n13994) );
  NAND U19547 ( .A(n13994), .B(n21327), .Z(n13995) );
  NAND U19548 ( .A(n13995), .B(n21329), .Z(n13996) );
  AND U19549 ( .A(n21331), .B(n13996), .Z(n13997) );
  NANDN U19550 ( .A(n13997), .B(n21333), .Z(n13998) );
  NAND U19551 ( .A(n13998), .B(n21336), .Z(n13999) );
  NAND U19552 ( .A(n13999), .B(n21337), .Z(n14000) );
  NAND U19553 ( .A(n14000), .B(n21339), .Z(n14001) );
  NAND U19554 ( .A(n14001), .B(n21341), .Z(n14002) );
  AND U19555 ( .A(n21343), .B(n14002), .Z(n14003) );
  NANDN U19556 ( .A(n14003), .B(n21345), .Z(n14004) );
  NAND U19557 ( .A(n14004), .B(n21348), .Z(n14005) );
  NAND U19558 ( .A(n14005), .B(n21349), .Z(n14006) );
  NAND U19559 ( .A(n14006), .B(n21351), .Z(n14007) );
  NAND U19560 ( .A(n14007), .B(n21353), .Z(n14008) );
  AND U19561 ( .A(n21355), .B(n14008), .Z(n14009) );
  NANDN U19562 ( .A(n14009), .B(n21357), .Z(n14010) );
  NAND U19563 ( .A(n14010), .B(n21360), .Z(n14011) );
  NANDN U19564 ( .A(n21362), .B(n14011), .Z(n14012) );
  NANDN U19565 ( .A(n21364), .B(n14012), .Z(n14013) );
  NAND U19566 ( .A(n14013), .B(n21365), .Z(n14014) );
  AND U19567 ( .A(n21367), .B(n14014), .Z(n14015) );
  OR U19568 ( .A(n21370), .B(n14015), .Z(n14016) );
  NAND U19569 ( .A(n14016), .B(n21371), .Z(n14017) );
  NANDN U19570 ( .A(n21374), .B(n14017), .Z(n14018) );
  NAND U19571 ( .A(n14018), .B(n21375), .Z(n14019) );
  NANDN U19572 ( .A(n21377), .B(n14019), .Z(n14020) );
  AND U19573 ( .A(n21379), .B(n14020), .Z(n14021) );
  OR U19574 ( .A(n21382), .B(n14021), .Z(n14022) );
  NAND U19575 ( .A(n14022), .B(n21383), .Z(n14023) );
  NANDN U19576 ( .A(n21386), .B(n14023), .Z(n14024) );
  NAND U19577 ( .A(n14024), .B(n21387), .Z(n14025) );
  NANDN U19578 ( .A(n21389), .B(n14025), .Z(n14026) );
  AND U19579 ( .A(n21391), .B(n14026), .Z(n14027) );
  OR U19580 ( .A(n21394), .B(n14027), .Z(n14028) );
  NAND U19581 ( .A(n14028), .B(n21395), .Z(n14029) );
  NAND U19582 ( .A(n14029), .B(n21397), .Z(n14030) );
  NANDN U19583 ( .A(n21400), .B(n14030), .Z(n14031) );
  NANDN U19584 ( .A(n21401), .B(n14031), .Z(n14032) );
  AND U19585 ( .A(n21403), .B(n14032), .Z(n14033) );
  OR U19586 ( .A(n21406), .B(n14033), .Z(n14034) );
  NAND U19587 ( .A(n14034), .B(n21407), .Z(n14035) );
  NANDN U19588 ( .A(n21410), .B(n14035), .Z(n14036) );
  NAND U19589 ( .A(n14036), .B(n21411), .Z(n14037) );
  NANDN U19590 ( .A(n21413), .B(n14037), .Z(n14038) );
  AND U19591 ( .A(n21415), .B(n14038), .Z(n14039) );
  OR U19592 ( .A(n21418), .B(n14039), .Z(n14040) );
  NAND U19593 ( .A(n14040), .B(n21419), .Z(n14041) );
  NANDN U19594 ( .A(n21422), .B(n14041), .Z(n14042) );
  NAND U19595 ( .A(n14042), .B(n21423), .Z(n14043) );
  NANDN U19596 ( .A(n21425), .B(n14043), .Z(n14045) );
  NAND U19597 ( .A(n14045), .B(n14044), .Z(n14046) );
  NANDN U19598 ( .A(n14046), .B(n21427), .Z(n14047) );
  NANDN U19599 ( .A(n21430), .B(n14047), .Z(n14049) );
  NAND U19600 ( .A(n14049), .B(n14048), .Z(n14050) );
  NANDN U19601 ( .A(n21434), .B(n14050), .Z(n14051) );
  NAND U19602 ( .A(n14051), .B(n21435), .Z(n14052) );
  ANDN U19603 ( .B(n14052), .A(n21437), .Z(n14053) );
  NANDN U19604 ( .A(n14053), .B(n21439), .Z(n14054) );
  ANDN U19605 ( .B(n14054), .A(n21442), .Z(n14055) );
  OR U19606 ( .A(n14056), .B(n14055), .Z(n14057) );
  NANDN U19607 ( .A(n14058), .B(n14057), .Z(n14060) );
  ANDN U19608 ( .B(n14060), .A(n14059), .Z(n14061) );
  OR U19609 ( .A(n14061), .B(x[850]), .Z(n14064) );
  XOR U19610 ( .A(x[850]), .B(n14061), .Z(n14062) );
  NAND U19611 ( .A(n14062), .B(y[850]), .Z(n14063) );
  NAND U19612 ( .A(n14064), .B(n14063), .Z(n14065) );
  AND U19613 ( .A(n21450), .B(n14065), .Z(n14066) );
  ANDN U19614 ( .B(n21451), .A(n14066), .Z(n14068) );
  NAND U19615 ( .A(n14068), .B(n14067), .Z(n14069) );
  AND U19616 ( .A(n21453), .B(n14069), .Z(n14070) );
  NANDN U19617 ( .A(n14070), .B(n21455), .Z(n14071) );
  NAND U19618 ( .A(n14071), .B(n21457), .Z(n14072) );
  NAND U19619 ( .A(n14072), .B(n21459), .Z(n14073) );
  NAND U19620 ( .A(n14073), .B(n21462), .Z(n14074) );
  NAND U19621 ( .A(n14074), .B(n21464), .Z(n14075) );
  ANDN U19622 ( .B(n14075), .A(n21467), .Z(n14076) );
  ANDN U19623 ( .B(n21471), .A(n14076), .Z(n14077) );
  NANDN U19624 ( .A(n14078), .B(n14077), .Z(n14079) );
  AND U19625 ( .A(n21473), .B(n14079), .Z(n14080) );
  ANDN U19626 ( .B(n21476), .A(n14080), .Z(n14082) );
  NAND U19627 ( .A(n14082), .B(n14081), .Z(n14083) );
  ANDN U19628 ( .B(n14083), .A(n21478), .Z(n14085) );
  NANDN U19629 ( .A(n14085), .B(n14084), .Z(n14086) );
  NANDN U19630 ( .A(n21482), .B(n14086), .Z(n14087) );
  NANDN U19631 ( .A(n21484), .B(n14087), .Z(n14088) );
  NANDN U19632 ( .A(n21486), .B(n14088), .Z(n14089) );
  NAND U19633 ( .A(n14089), .B(n21487), .Z(n14090) );
  ANDN U19634 ( .B(n14090), .A(n21490), .Z(n14091) );
  NANDN U19635 ( .A(n14091), .B(n21491), .Z(n14092) );
  NAND U19636 ( .A(n14092), .B(n21494), .Z(n14093) );
  NAND U19637 ( .A(n14093), .B(n21495), .Z(n14094) );
  NANDN U19638 ( .A(n21498), .B(n14094), .Z(n14095) );
  NAND U19639 ( .A(n14095), .B(n21499), .Z(n14096) );
  ANDN U19640 ( .B(n14096), .A(n21502), .Z(n14097) );
  NANDN U19641 ( .A(n14097), .B(n21503), .Z(n14098) );
  NAND U19642 ( .A(n14098), .B(n21506), .Z(n14099) );
  AND U19643 ( .A(n21507), .B(n14099), .Z(n14100) );
  OR U19644 ( .A(n21510), .B(n14100), .Z(n14101) );
  NAND U19645 ( .A(n14101), .B(n21511), .Z(n14102) );
  NANDN U19646 ( .A(n21514), .B(n14102), .Z(n14103) );
  NAND U19647 ( .A(n14103), .B(n21515), .Z(n14104) );
  NANDN U19648 ( .A(n21517), .B(n14104), .Z(n14105) );
  AND U19649 ( .A(n21520), .B(n14105), .Z(n14106) );
  NANDN U19650 ( .A(n14106), .B(n21523), .Z(n14108) );
  NAND U19651 ( .A(n14108), .B(n14107), .Z(n14109) );
  NANDN U19652 ( .A(n14110), .B(n14109), .Z(n14111) );
  NAND U19653 ( .A(n14111), .B(n21531), .Z(n14112) );
  NANDN U19654 ( .A(n21534), .B(n14112), .Z(n14114) );
  ANDN U19655 ( .B(n14114), .A(n14113), .Z(n14115) );
  NANDN U19656 ( .A(n14115), .B(n21537), .Z(n14116) );
  AND U19657 ( .A(n14117), .B(n14116), .Z(n14118) );
  OR U19658 ( .A(n21541), .B(n14118), .Z(n14119) );
  NAND U19659 ( .A(n14119), .B(n21543), .Z(n14120) );
  NANDN U19660 ( .A(n21546), .B(n14120), .Z(n14121) );
  NAND U19661 ( .A(n14121), .B(n21547), .Z(n14122) );
  NANDN U19662 ( .A(n21550), .B(n14122), .Z(n14123) );
  AND U19663 ( .A(n21552), .B(n14123), .Z(n14124) );
  NANDN U19664 ( .A(n14124), .B(n21555), .Z(n14125) );
  NANDN U19665 ( .A(n14126), .B(n14125), .Z(n14127) );
  NANDN U19666 ( .A(n21559), .B(n14127), .Z(n14128) );
  NAND U19667 ( .A(n14128), .B(n21561), .Z(n14129) );
  NANDN U19668 ( .A(n21564), .B(n14129), .Z(n14130) );
  AND U19669 ( .A(n21565), .B(n14130), .Z(n14131) );
  NANDN U19670 ( .A(n14131), .B(n21567), .Z(n14132) );
  NAND U19671 ( .A(n14132), .B(n21569), .Z(n14133) );
  NAND U19672 ( .A(n14133), .B(n21572), .Z(n14134) );
  NAND U19673 ( .A(n14134), .B(n21573), .Z(n14135) );
  NAND U19674 ( .A(n14135), .B(n21575), .Z(n14136) );
  AND U19675 ( .A(n21577), .B(n14136), .Z(n14137) );
  NANDN U19676 ( .A(n14137), .B(n21579), .Z(n14138) );
  NAND U19677 ( .A(n14138), .B(n21582), .Z(n14139) );
  NAND U19678 ( .A(n14139), .B(n21585), .Z(n14140) );
  NANDN U19679 ( .A(n14141), .B(n14140), .Z(n14142) );
  NANDN U19680 ( .A(n14143), .B(n14142), .Z(n14145) );
  ANDN U19681 ( .B(n14145), .A(n14144), .Z(n14146) );
  NANDN U19682 ( .A(n14146), .B(n21599), .Z(n14147) );
  NAND U19683 ( .A(n14147), .B(n21601), .Z(n14148) );
  NAND U19684 ( .A(n14148), .B(n21604), .Z(n14149) );
  NAND U19685 ( .A(n14149), .B(n21605), .Z(n14150) );
  NAND U19686 ( .A(n14150), .B(n21607), .Z(n14151) );
  AND U19687 ( .A(n21609), .B(n14151), .Z(n14152) );
  NANDN U19688 ( .A(n14152), .B(n21611), .Z(n14153) );
  NAND U19689 ( .A(n14153), .B(n21613), .Z(n14154) );
  NAND U19690 ( .A(n14154), .B(n21616), .Z(n14155) );
  NAND U19691 ( .A(n14155), .B(n21617), .Z(n14156) );
  NAND U19692 ( .A(n14156), .B(n21619), .Z(n14157) );
  AND U19693 ( .A(n21621), .B(n14157), .Z(n14159) );
  NANDN U19694 ( .A(n14159), .B(n14158), .Z(n14160) );
  ANDN U19695 ( .B(n14160), .A(n21626), .Z(n14161) );
  ANDN U19696 ( .B(n14162), .A(n14161), .Z(n14166) );
  XNOR U19697 ( .A(x[921]), .B(y[921]), .Z(n14163) );
  NAND U19698 ( .A(n14164), .B(n14163), .Z(n14165) );
  AND U19699 ( .A(n14166), .B(n14165), .Z(n14168) );
  OR U19700 ( .A(n14168), .B(y[922]), .Z(n14167) );
  AND U19701 ( .A(n21631), .B(n14167), .Z(n14171) );
  XOR U19702 ( .A(y[922]), .B(n14168), .Z(n14169) );
  NAND U19703 ( .A(x[922]), .B(n14169), .Z(n14170) );
  NAND U19704 ( .A(n14171), .B(n14170), .Z(n14172) );
  NAND U19705 ( .A(n14173), .B(n14172), .Z(n14174) );
  NAND U19706 ( .A(n14174), .B(n21635), .Z(n14175) );
  NAND U19707 ( .A(n14175), .B(n21637), .Z(n14176) );
  NAND U19708 ( .A(n14176), .B(n21640), .Z(n14177) );
  AND U19709 ( .A(n21641), .B(n14177), .Z(n14178) );
  NANDN U19710 ( .A(n14178), .B(n21643), .Z(n14179) );
  NAND U19711 ( .A(n14179), .B(n21647), .Z(n14180) );
  NAND U19712 ( .A(n14180), .B(n21649), .Z(n14181) );
  NANDN U19713 ( .A(n14182), .B(n14181), .Z(n14183) );
  NANDN U19714 ( .A(n14184), .B(n14183), .Z(n14186) );
  ANDN U19715 ( .B(n14186), .A(n14185), .Z(n14187) );
  NANDN U19716 ( .A(n14187), .B(n21662), .Z(n14188) );
  NAND U19717 ( .A(n14188), .B(n21664), .Z(n14189) );
  NAND U19718 ( .A(n14189), .B(n21667), .Z(n14190) );
  NAND U19719 ( .A(n14190), .B(n21668), .Z(n14191) );
  NAND U19720 ( .A(n14191), .B(n21670), .Z(n14192) );
  AND U19721 ( .A(n21672), .B(n14192), .Z(n14193) );
  NANDN U19722 ( .A(n14193), .B(n21674), .Z(n14194) );
  NAND U19723 ( .A(n14194), .B(n21676), .Z(n14195) );
  NAND U19724 ( .A(n14195), .B(n21679), .Z(n14196) );
  NAND U19725 ( .A(n14196), .B(n21681), .Z(n14197) );
  NAND U19726 ( .A(n14197), .B(n20297), .Z(n14199) );
  ANDN U19727 ( .B(n14199), .A(n14198), .Z(n14201) );
  NANDN U19728 ( .A(n14201), .B(n14200), .Z(n14202) );
  AND U19729 ( .A(n21688), .B(n14202), .Z(n14203) );
  ANDN U19730 ( .B(n14204), .A(n14203), .Z(n14207) );
  XNOR U19731 ( .A(x[945]), .B(y[945]), .Z(n14205) );
  NAND U19732 ( .A(n14205), .B(n20296), .Z(n14206) );
  AND U19733 ( .A(n14207), .B(n14206), .Z(n14209) );
  OR U19734 ( .A(n14209), .B(y[946]), .Z(n14208) );
  AND U19735 ( .A(n21695), .B(n14208), .Z(n14212) );
  XOR U19736 ( .A(y[946]), .B(n14209), .Z(n14210) );
  NAND U19737 ( .A(n14210), .B(x[946]), .Z(n14211) );
  NAND U19738 ( .A(n14212), .B(n14211), .Z(n14213) );
  NAND U19739 ( .A(n14214), .B(n14213), .Z(n14215) );
  NAND U19740 ( .A(n14215), .B(n21698), .Z(n14216) );
  NAND U19741 ( .A(n14216), .B(n21700), .Z(n14217) );
  NAND U19742 ( .A(n14217), .B(n21702), .Z(n14218) );
  AND U19743 ( .A(n21704), .B(n14218), .Z(n14219) );
  NANDN U19744 ( .A(n14219), .B(n21707), .Z(n14220) );
  ANDN U19745 ( .B(n14220), .A(n21708), .Z(n14221) );
  NANDN U19746 ( .A(n14221), .B(n20293), .Z(n14222) );
  NANDN U19747 ( .A(n14223), .B(n14222), .Z(n14224) );
  NAND U19748 ( .A(n14224), .B(n20294), .Z(n14225) );
  NANDN U19749 ( .A(n21714), .B(n14225), .Z(n14226) );
  NANDN U19750 ( .A(n21718), .B(n14226), .Z(n14227) );
  AND U19751 ( .A(n14228), .B(n14227), .Z(n14229) );
  NAND U19752 ( .A(n14229), .B(n21720), .Z(n14230) );
  NANDN U19753 ( .A(n21722), .B(n14230), .Z(n14232) );
  ANDN U19754 ( .B(n14232), .A(n14231), .Z(n14233) );
  OR U19755 ( .A(n21727), .B(n14233), .Z(n14234) );
  NAND U19756 ( .A(n14234), .B(n21728), .Z(n14235) );
  NANDN U19757 ( .A(n21731), .B(n14235), .Z(n14236) );
  NAND U19758 ( .A(n14236), .B(n21732), .Z(n14237) );
  NANDN U19759 ( .A(n21734), .B(n14237), .Z(n14238) );
  NAND U19760 ( .A(n14238), .B(n21736), .Z(n14239) );
  NAND U19761 ( .A(n14239), .B(n21738), .Z(n14240) );
  NAND U19762 ( .A(n14240), .B(n21740), .Z(n14241) );
  ANDN U19763 ( .B(n14241), .A(n21743), .Z(n14242) );
  NANDN U19764 ( .A(n14242), .B(n21744), .Z(n14243) );
  NANDN U19765 ( .A(n21746), .B(n14243), .Z(n14244) );
  NAND U19766 ( .A(n14244), .B(n21748), .Z(n14245) );
  NAND U19767 ( .A(n14245), .B(n21750), .Z(n14246) );
  NAND U19768 ( .A(n14246), .B(n21752), .Z(n14247) );
  ANDN U19769 ( .B(n14247), .A(n21755), .Z(n14248) );
  NANDN U19770 ( .A(n14248), .B(n21756), .Z(n14249) );
  NANDN U19771 ( .A(n21758), .B(n14249), .Z(n14250) );
  NAND U19772 ( .A(n14250), .B(n21760), .Z(n14251) );
  NANDN U19773 ( .A(n21763), .B(n14251), .Z(n14252) );
  NAND U19774 ( .A(n14252), .B(n21764), .Z(n14253) );
  AND U19775 ( .A(n21766), .B(n14253), .Z(n14254) );
  NANDN U19776 ( .A(n14254), .B(n21768), .Z(n14255) );
  NANDN U19777 ( .A(n21770), .B(n14255), .Z(n14256) );
  NAND U19778 ( .A(n14256), .B(n21772), .Z(n14257) );
  NANDN U19779 ( .A(n21775), .B(n14257), .Z(n14258) );
  NAND U19780 ( .A(n14258), .B(n21776), .Z(n14259) );
  AND U19781 ( .A(n21778), .B(n14259), .Z(n14260) );
  NANDN U19782 ( .A(n14260), .B(n21780), .Z(n14261) );
  NANDN U19783 ( .A(n21782), .B(n14261), .Z(n14262) );
  NAND U19784 ( .A(n14262), .B(n21784), .Z(n14263) );
  NANDN U19785 ( .A(n21787), .B(n14263), .Z(n14264) );
  NAND U19786 ( .A(n14264), .B(n21788), .Z(n14265) );
  ANDN U19787 ( .B(n14265), .A(n21791), .Z(n14266) );
  NANDN U19788 ( .A(n14266), .B(n21793), .Z(n14267) );
  NAND U19789 ( .A(n14267), .B(n21796), .Z(n14268) );
  NAND U19790 ( .A(n14268), .B(n21799), .Z(n14270) );
  OR U19791 ( .A(n14270), .B(n14269), .Z(n14271) );
  NANDN U19792 ( .A(n21803), .B(n14271), .Z(n14272) );
  NAND U19793 ( .A(n14272), .B(n21804), .Z(n14273) );
  NAND U19794 ( .A(n14273), .B(n21807), .Z(n14274) );
  NAND U19795 ( .A(n14274), .B(n21808), .Z(n14275) );
  AND U19796 ( .A(n21810), .B(n14275), .Z(n14276) );
  NANDN U19797 ( .A(n14276), .B(n21812), .Z(n14277) );
  NAND U19798 ( .A(n14277), .B(n21814), .Z(n14278) );
  NAND U19799 ( .A(n14278), .B(n21816), .Z(n14279) );
  NAND U19800 ( .A(n14279), .B(n21819), .Z(n14280) );
  NAND U19801 ( .A(n14280), .B(n21821), .Z(n14281) );
  ANDN U19802 ( .B(n14281), .A(n21824), .Z(n14283) );
  NANDN U19803 ( .A(n14283), .B(n14282), .Z(n14284) );
  NAND U19804 ( .A(n14284), .B(n21830), .Z(n14285) );
  NAND U19805 ( .A(n14285), .B(n21832), .Z(n14286) );
  NAND U19806 ( .A(n14286), .B(n21835), .Z(n14287) );
  NAND U19807 ( .A(n14287), .B(n21836), .Z(n14288) );
  AND U19808 ( .A(n21838), .B(n14288), .Z(n14289) );
  NANDN U19809 ( .A(n14289), .B(n21840), .Z(n14290) );
  AND U19810 ( .A(n21842), .B(n14290), .Z(n14291) );
  NANDN U19811 ( .A(n14291), .B(n21844), .Z(n14292) );
  NAND U19812 ( .A(n14292), .B(n21847), .Z(n14293) );
  NAND U19813 ( .A(n14293), .B(n21849), .Z(n14294) );
  NAND U19814 ( .A(n14294), .B(n20289), .Z(n14296) );
  NAND U19815 ( .A(n14296), .B(n14295), .Z(n14297) );
  AND U19816 ( .A(n20290), .B(n14297), .Z(n14298) );
  NANDN U19817 ( .A(n14298), .B(n21856), .Z(n14303) );
  NANDN U19818 ( .A(n14300), .B(n14299), .Z(n14301) );
  NANDN U19819 ( .A(n14302), .B(n14301), .Z(n21858) );
  ANDN U19820 ( .B(n14303), .A(n21858), .Z(n14304) );
  NANDN U19821 ( .A(n14304), .B(n21860), .Z(n14305) );
  NAND U19822 ( .A(n14305), .B(n21862), .Z(n14306) );
  NANDN U19823 ( .A(n14307), .B(n14306), .Z(n14308) );
  NANDN U19824 ( .A(n14308), .B(x[1021]), .Z(n14311) );
  XNOR U19825 ( .A(n14308), .B(x[1021]), .Z(n14309) );
  NANDN U19826 ( .A(y[1021]), .B(n14309), .Z(n14310) );
  NAND U19827 ( .A(n14311), .B(n14310), .Z(n14312) );
  NAND U19828 ( .A(n14313), .B(n14312), .Z(n14314) );
  NAND U19829 ( .A(n14315), .B(n14314), .Z(n14316) );
  NAND U19830 ( .A(n14317), .B(n14316), .Z(n14318) );
  NAND U19831 ( .A(n14318), .B(n21874), .Z(n14321) );
  NANDN U19832 ( .A(x[1026]), .B(y[1026]), .Z(n14320) );
  ANDN U19833 ( .B(n14320), .A(n14319), .Z(n21876) );
  NAND U19834 ( .A(n14321), .B(n21876), .Z(n14322) );
  NANDN U19835 ( .A(n21879), .B(n14322), .Z(n14324) );
  ANDN U19836 ( .B(n14324), .A(n14323), .Z(n14325) );
  NAND U19837 ( .A(n14325), .B(n21880), .Z(n14326) );
  NAND U19838 ( .A(n14327), .B(n14326), .Z(n14328) );
  NAND U19839 ( .A(n14329), .B(n14328), .Z(n14330) );
  NANDN U19840 ( .A(n21891), .B(n14330), .Z(n14333) );
  NANDN U19841 ( .A(x[1031]), .B(y[1031]), .Z(n14332) );
  NANDN U19842 ( .A(x[1032]), .B(y[1032]), .Z(n14331) );
  AND U19843 ( .A(n14332), .B(n14331), .Z(n21892) );
  NAND U19844 ( .A(n14333), .B(n21892), .Z(n14334) );
  NANDN U19845 ( .A(n21894), .B(n14334), .Z(n14337) );
  NANDN U19846 ( .A(x[1033]), .B(y[1033]), .Z(n14335) );
  NANDN U19847 ( .A(n14336), .B(n14335), .Z(n21897) );
  ANDN U19848 ( .B(n14337), .A(n21897), .Z(n14338) );
  NANDN U19849 ( .A(n14338), .B(n21898), .Z(n14339) );
  NAND U19850 ( .A(n14339), .B(n21900), .Z(n14340) );
  NAND U19851 ( .A(n14340), .B(n21902), .Z(n14344) );
  NAND U19852 ( .A(n14341), .B(y[1038]), .Z(n14343) );
  ANDN U19853 ( .B(n14343), .A(n14342), .Z(n21904) );
  NAND U19854 ( .A(n14344), .B(n21904), .Z(n14345) );
  NANDN U19855 ( .A(n21906), .B(n14345), .Z(n14347) );
  ANDN U19856 ( .B(n14347), .A(n14346), .Z(n14348) );
  NAND U19857 ( .A(n14348), .B(n21908), .Z(n14349) );
  NAND U19858 ( .A(n14350), .B(n14349), .Z(n14351) );
  NAND U19859 ( .A(n14352), .B(n14351), .Z(n14359) );
  NANDN U19860 ( .A(n14354), .B(n14353), .Z(n14355) );
  NANDN U19861 ( .A(n14356), .B(n14355), .Z(n14358) );
  ANDN U19862 ( .B(n14358), .A(n14357), .Z(n21919) );
  NAND U19863 ( .A(n14359), .B(n21919), .Z(n14360) );
  NAND U19864 ( .A(n14360), .B(n21920), .Z(n14361) );
  NANDN U19865 ( .A(n21923), .B(n14361), .Z(n14362) );
  AND U19866 ( .A(n21924), .B(n14362), .Z(n14363) );
  OR U19867 ( .A(n21927), .B(n14363), .Z(n14364) );
  NANDN U19868 ( .A(n21929), .B(n14364), .Z(n14365) );
  NANDN U19869 ( .A(n21931), .B(n14365), .Z(n14366) );
  NAND U19870 ( .A(n14367), .B(n14366), .Z(n14368) );
  NAND U19871 ( .A(n14368), .B(n21934), .Z(n14369) );
  NANDN U19872 ( .A(n14369), .B(n21938), .Z(n14370) );
  AND U19873 ( .A(n14371), .B(n14370), .Z(n14372) );
  OR U19874 ( .A(n21943), .B(n14372), .Z(n14373) );
  NAND U19875 ( .A(n14373), .B(n21944), .Z(n14374) );
  NAND U19876 ( .A(n14374), .B(n21946), .Z(n14375) );
  NAND U19877 ( .A(n14375), .B(n21949), .Z(n14376) );
  NANDN U19878 ( .A(n21951), .B(n14376), .Z(n14377) );
  NANDN U19879 ( .A(n21953), .B(n14377), .Z(n14378) );
  NANDN U19880 ( .A(n21954), .B(n14378), .Z(n14379) );
  AND U19881 ( .A(n21956), .B(n14379), .Z(n14381) );
  NAND U19882 ( .A(n14381), .B(n14380), .Z(n14382) );
  NAND U19883 ( .A(n14382), .B(n21959), .Z(n14384) );
  NAND U19884 ( .A(n14384), .B(n14383), .Z(n14385) );
  AND U19885 ( .A(n21962), .B(n14385), .Z(n14386) );
  NANDN U19886 ( .A(n14386), .B(n21964), .Z(n14387) );
  NAND U19887 ( .A(n14387), .B(n21966), .Z(n14388) );
  NAND U19888 ( .A(n14388), .B(n21968), .Z(n14389) );
  NAND U19889 ( .A(n14389), .B(n21971), .Z(n14390) );
  NAND U19890 ( .A(n14390), .B(n21972), .Z(n14391) );
  AND U19891 ( .A(n21974), .B(n14391), .Z(n14392) );
  OR U19892 ( .A(n21977), .B(n14392), .Z(n14393) );
  NANDN U19893 ( .A(n21979), .B(n14393), .Z(n14395) );
  NAND U19894 ( .A(n14395), .B(n14394), .Z(n14396) );
  NANDN U19895 ( .A(n14396), .B(n21980), .Z(n14397) );
  AND U19896 ( .A(n21982), .B(n14397), .Z(n14398) );
  NAND U19897 ( .A(n14398), .B(n21986), .Z(n14399) );
  NAND U19898 ( .A(n14400), .B(n14399), .Z(n14403) );
  ANDN U19899 ( .B(n14402), .A(n14401), .Z(n21990) );
  NAND U19900 ( .A(n14403), .B(n21990), .Z(n14404) );
  NANDN U19901 ( .A(n21993), .B(n14404), .Z(n14405) );
  AND U19902 ( .A(n21994), .B(n14405), .Z(n14406) );
  OR U19903 ( .A(n21997), .B(n14406), .Z(n14407) );
  NAND U19904 ( .A(n14407), .B(n21998), .Z(n14408) );
  NANDN U19905 ( .A(n22000), .B(n14408), .Z(n14409) );
  NAND U19906 ( .A(n14409), .B(n22002), .Z(n14410) );
  NANDN U19907 ( .A(n22005), .B(n14410), .Z(n14411) );
  ANDN U19908 ( .B(n14411), .A(n22007), .Z(n14412) );
  OR U19909 ( .A(n22009), .B(n14412), .Z(n14417) );
  NANDN U19910 ( .A(n14414), .B(n14413), .Z(n14416) );
  ANDN U19911 ( .B(n14416), .A(n14415), .Z(n22010) );
  NAND U19912 ( .A(n14417), .B(n22010), .Z(n14418) );
  NAND U19913 ( .A(n14418), .B(n22013), .Z(n14425) );
  OR U19914 ( .A(n14420), .B(n14419), .Z(n14421) );
  NANDN U19915 ( .A(n14422), .B(n14421), .Z(n14424) );
  ANDN U19916 ( .B(n14424), .A(n14423), .Z(n22014) );
  NAND U19917 ( .A(n14425), .B(n22014), .Z(n14426) );
  NAND U19918 ( .A(n14426), .B(n22016), .Z(n14427) );
  NAND U19919 ( .A(n14427), .B(n22018), .Z(n14428) );
  NAND U19920 ( .A(n14428), .B(n22020), .Z(n14429) );
  NAND U19921 ( .A(n14429), .B(n22022), .Z(n14433) );
  NAND U19922 ( .A(n14430), .B(y[1098]), .Z(n14431) );
  NANDN U19923 ( .A(n14432), .B(n14431), .Z(n22024) );
  ANDN U19924 ( .B(n14433), .A(n22024), .Z(n14434) );
  OR U19925 ( .A(n22027), .B(n14434), .Z(n14435) );
  AND U19926 ( .A(n14436), .B(n14435), .Z(n14437) );
  ANDN U19927 ( .B(n22034), .A(n14437), .Z(n14438) );
  NAND U19928 ( .A(n14438), .B(n22030), .Z(n14439) );
  ANDN U19929 ( .B(n14439), .A(n22036), .Z(n14440) );
  NANDN U19930 ( .A(n14441), .B(n14440), .Z(n14442) );
  NANDN U19931 ( .A(n22039), .B(n14442), .Z(n14443) );
  AND U19932 ( .A(n22040), .B(n14443), .Z(n14444) );
  NANDN U19933 ( .A(n14444), .B(n22042), .Z(n14445) );
  NAND U19934 ( .A(n14445), .B(n22044), .Z(n14446) );
  NAND U19935 ( .A(n14446), .B(n22046), .Z(n14447) );
  NAND U19936 ( .A(n14448), .B(n14447), .Z(n14449) );
  NANDN U19937 ( .A(n22053), .B(n14449), .Z(n14450) );
  NAND U19938 ( .A(n14451), .B(n14450), .Z(n14452) );
  NANDN U19939 ( .A(n22057), .B(n14452), .Z(n14453) );
  NANDN U19940 ( .A(n14454), .B(n14453), .Z(n14455) );
  NANDN U19941 ( .A(n22060), .B(n14455), .Z(n14456) );
  AND U19942 ( .A(n22062), .B(n14456), .Z(n14457) );
  OR U19943 ( .A(n22065), .B(n14457), .Z(n14458) );
  NAND U19944 ( .A(n14458), .B(n22066), .Z(n14459) );
  NANDN U19945 ( .A(n22069), .B(n14459), .Z(n14460) );
  NAND U19946 ( .A(n14460), .B(n22070), .Z(n14461) );
  NANDN U19947 ( .A(n22072), .B(n14461), .Z(n14462) );
  AND U19948 ( .A(n22074), .B(n14462), .Z(n14463) );
  OR U19949 ( .A(n22077), .B(n14463), .Z(n14464) );
  AND U19950 ( .A(n14465), .B(n14464), .Z(n14466) );
  OR U19951 ( .A(n14467), .B(n14466), .Z(n14468) );
  AND U19952 ( .A(n14469), .B(n14468), .Z(n14470) );
  OR U19953 ( .A(n22089), .B(n14470), .Z(n14473) );
  AND U19954 ( .A(n14472), .B(n14471), .Z(n22090) );
  NAND U19955 ( .A(n14473), .B(n22090), .Z(n14474) );
  NANDN U19956 ( .A(n22093), .B(n14474), .Z(n14475) );
  NAND U19957 ( .A(n14475), .B(n22094), .Z(n14476) );
  NANDN U19958 ( .A(n22096), .B(n14476), .Z(n14477) );
  AND U19959 ( .A(n22098), .B(n14477), .Z(n14478) );
  OR U19960 ( .A(n22100), .B(n14478), .Z(n14481) );
  NANDN U19961 ( .A(x[1134]), .B(y[1134]), .Z(n14480) );
  ANDN U19962 ( .B(n14480), .A(n14479), .Z(n22102) );
  NAND U19963 ( .A(n14481), .B(n22102), .Z(n14484) );
  NANDN U19964 ( .A(y[1134]), .B(x[1134]), .Z(n14483) );
  ANDN U19965 ( .B(n14483), .A(n14482), .Z(n22104) );
  NAND U19966 ( .A(n14484), .B(n22104), .Z(n14485) );
  NAND U19967 ( .A(n14486), .B(n14485), .Z(n14487) );
  NANDN U19968 ( .A(n14488), .B(n14487), .Z(n14489) );
  NAND U19969 ( .A(n14490), .B(n14489), .Z(n14491) );
  NANDN U19970 ( .A(n22117), .B(n14491), .Z(n14492) );
  NAND U19971 ( .A(n14492), .B(n22118), .Z(n14493) );
  NAND U19972 ( .A(n14493), .B(n22120), .Z(n14494) );
  AND U19973 ( .A(n22122), .B(n14494), .Z(n14495) );
  NANDN U19974 ( .A(n14495), .B(n22125), .Z(n14496) );
  NAND U19975 ( .A(n14496), .B(n22126), .Z(n14497) );
  NAND U19976 ( .A(n14497), .B(n22128), .Z(n14498) );
  NAND U19977 ( .A(n14498), .B(n22130), .Z(n14499) );
  NANDN U19978 ( .A(n22133), .B(n14499), .Z(n14504) );
  NANDN U19979 ( .A(n14501), .B(n14500), .Z(n14502) );
  NAND U19980 ( .A(n14503), .B(n14502), .Z(n22135) );
  ANDN U19981 ( .B(n14504), .A(n22135), .Z(n14507) );
  NANDN U19982 ( .A(y[1150]), .B(x[1150]), .Z(n14505) );
  NANDN U19983 ( .A(n14506), .B(n14505), .Z(n22136) );
  OR U19984 ( .A(n14507), .B(n22136), .Z(n14508) );
  NANDN U19985 ( .A(n22139), .B(n14508), .Z(n14511) );
  NANDN U19986 ( .A(y[1152]), .B(x[1152]), .Z(n14509) );
  NANDN U19987 ( .A(n14510), .B(n14509), .Z(n22141) );
  ANDN U19988 ( .B(n14511), .A(n22141), .Z(n14512) );
  NANDN U19989 ( .A(n14512), .B(n22142), .Z(n14513) );
  NANDN U19990 ( .A(n22145), .B(n14513), .Z(n14514) );
  NAND U19991 ( .A(n14514), .B(n22146), .Z(n14515) );
  NANDN U19992 ( .A(n22148), .B(n14515), .Z(n14517) );
  ANDN U19993 ( .B(n14517), .A(n14516), .Z(n14518) );
  OR U19994 ( .A(n14519), .B(n14518), .Z(n14520) );
  AND U19995 ( .A(n14521), .B(n14520), .Z(n14525) );
  NAND U19996 ( .A(n14523), .B(n14522), .Z(n14524) );
  NANDN U19997 ( .A(n14525), .B(n14524), .Z(n14526) );
  AND U19998 ( .A(n14527), .B(n14526), .Z(n14528) );
  OR U19999 ( .A(n22157), .B(n14528), .Z(n14529) );
  NAND U20000 ( .A(n14529), .B(n22158), .Z(n14530) );
  NANDN U20001 ( .A(n22160), .B(n14530), .Z(n14531) );
  NAND U20002 ( .A(n14531), .B(n22162), .Z(n14532) );
  NANDN U20003 ( .A(n22165), .B(n14532), .Z(n14533) );
  AND U20004 ( .A(n22166), .B(n14533), .Z(n14534) );
  OR U20005 ( .A(n22169), .B(n14534), .Z(n14535) );
  NANDN U20006 ( .A(n14536), .B(n14535), .Z(n14537) );
  NANDN U20007 ( .A(n14538), .B(n14537), .Z(n14539) );
  NAND U20008 ( .A(n14540), .B(n14539), .Z(n14541) );
  NANDN U20009 ( .A(n14542), .B(n14541), .Z(n14543) );
  NAND U20010 ( .A(n14544), .B(n14543), .Z(n14545) );
  NANDN U20011 ( .A(n22178), .B(n14545), .Z(n14548) );
  AND U20012 ( .A(n14547), .B(n14546), .Z(n22180) );
  NAND U20013 ( .A(n14548), .B(n22180), .Z(n14549) );
  NANDN U20014 ( .A(n22183), .B(n14549), .Z(n14550) );
  AND U20015 ( .A(n22184), .B(n14550), .Z(n14551) );
  OR U20016 ( .A(n22187), .B(n14551), .Z(n14552) );
  NAND U20017 ( .A(n14552), .B(n22188), .Z(n14553) );
  NANDN U20018 ( .A(n22190), .B(n14553), .Z(n14554) );
  NAND U20019 ( .A(n14554), .B(n22192), .Z(n14555) );
  NANDN U20020 ( .A(n22195), .B(n14555), .Z(n14557) );
  ANDN U20021 ( .B(n14557), .A(n14556), .Z(n14558) );
  NAND U20022 ( .A(n14558), .B(n22196), .Z(n14559) );
  AND U20023 ( .A(n22198), .B(n14559), .Z(n14560) );
  NAND U20024 ( .A(n14560), .B(n22203), .Z(n14561) );
  NAND U20025 ( .A(n14562), .B(n14561), .Z(n14563) );
  NANDN U20026 ( .A(n22207), .B(n14563), .Z(n14566) );
  NANDN U20027 ( .A(x[1188]), .B(y[1188]), .Z(n14565) );
  ANDN U20028 ( .B(n14565), .A(n14564), .Z(n22208) );
  NAND U20029 ( .A(n14566), .B(n22208), .Z(n14567) );
  NANDN U20030 ( .A(n22211), .B(n14567), .Z(n14570) );
  NANDN U20031 ( .A(x[1189]), .B(y[1189]), .Z(n14568) );
  NANDN U20032 ( .A(n14569), .B(n14568), .Z(n22213) );
  ANDN U20033 ( .B(n14570), .A(n22213), .Z(n14571) );
  NANDN U20034 ( .A(n14571), .B(n22214), .Z(n14572) );
  NANDN U20035 ( .A(n22217), .B(n14572), .Z(n14573) );
  NAND U20036 ( .A(n14573), .B(n22218), .Z(n14574) );
  NANDN U20037 ( .A(n22220), .B(n14574), .Z(n14578) );
  NAND U20038 ( .A(n14575), .B(x[1194]), .Z(n14577) );
  ANDN U20039 ( .B(n14577), .A(n14576), .Z(n22222) );
  NAND U20040 ( .A(n14578), .B(n22222), .Z(n14579) );
  AND U20041 ( .A(n14580), .B(n14579), .Z(n14581) );
  NAND U20042 ( .A(n14581), .B(n22225), .Z(n14582) );
  NANDN U20043 ( .A(n14583), .B(n14582), .Z(n14584) );
  ANDN U20044 ( .B(n14584), .A(n22232), .Z(n14586) );
  AND U20045 ( .A(n14586), .B(n14585), .Z(n14593) );
  NANDN U20046 ( .A(n14588), .B(n14587), .Z(n14589) );
  NANDN U20047 ( .A(n14590), .B(n14589), .Z(n14592) );
  ANDN U20048 ( .B(n14592), .A(n14591), .Z(n22234) );
  NANDN U20049 ( .A(n14593), .B(n22234), .Z(n14594) );
  NAND U20050 ( .A(n14594), .B(n22236), .Z(n14595) );
  NAND U20051 ( .A(n14595), .B(n22239), .Z(n14596) );
  AND U20052 ( .A(n22240), .B(n14596), .Z(n14597) );
  OR U20053 ( .A(n14597), .B(n22243), .Z(n14598) );
  AND U20054 ( .A(n22244), .B(n14598), .Z(n14599) );
  NANDN U20055 ( .A(n14599), .B(n22246), .Z(n14601) );
  ANDN U20056 ( .B(n14601), .A(n14600), .Z(n14602) );
  NAND U20057 ( .A(n14602), .B(n22248), .Z(n14603) );
  AND U20058 ( .A(n22251), .B(n14603), .Z(n14604) );
  NAND U20059 ( .A(n14604), .B(n22255), .Z(n14605) );
  NAND U20060 ( .A(n14606), .B(n14605), .Z(n14607) );
  NANDN U20061 ( .A(n22259), .B(n14607), .Z(n14608) );
  NANDN U20062 ( .A(n22260), .B(n14608), .Z(n14609) );
  NAND U20063 ( .A(n14609), .B(n22262), .Z(n14610) );
  ANDN U20064 ( .B(n14610), .A(n22265), .Z(n14611) );
  NANDN U20065 ( .A(n14611), .B(n22266), .Z(n14612) );
  AND U20066 ( .A(n22268), .B(n14612), .Z(n14613) );
  NANDN U20067 ( .A(n14613), .B(n22271), .Z(n14614) );
  NAND U20068 ( .A(n14614), .B(n22272), .Z(n14615) );
  NANDN U20069 ( .A(n22275), .B(n14615), .Z(n14618) );
  NOR U20070 ( .A(n14617), .B(n14616), .Z(n22276) );
  NAND U20071 ( .A(n14618), .B(n22276), .Z(n14619) );
  NANDN U20072 ( .A(n22279), .B(n14619), .Z(n14620) );
  AND U20073 ( .A(n22280), .B(n14620), .Z(n14627) );
  NANDN U20074 ( .A(n14622), .B(n14621), .Z(n14623) );
  NANDN U20075 ( .A(n14624), .B(n14623), .Z(n14626) );
  ANDN U20076 ( .B(n14626), .A(n14625), .Z(n22283) );
  NANDN U20077 ( .A(n14627), .B(n22283), .Z(n14628) );
  NAND U20078 ( .A(n14628), .B(n22284), .Z(n14629) );
  NANDN U20079 ( .A(n22286), .B(n14629), .Z(n14630) );
  NAND U20080 ( .A(n14630), .B(n22288), .Z(n14631) );
  NANDN U20081 ( .A(n22291), .B(n14631), .Z(n14632) );
  AND U20082 ( .A(n22292), .B(n14632), .Z(n14633) );
  NANDN U20083 ( .A(n14633), .B(n22294), .Z(n14634) );
  AND U20084 ( .A(n14635), .B(n14634), .Z(n14638) );
  NOR U20085 ( .A(n14637), .B(n14636), .Z(n22298) );
  NANDN U20086 ( .A(n14638), .B(n22298), .Z(n14639) );
  AND U20087 ( .A(n14640), .B(n14639), .Z(n14641) );
  NAND U20088 ( .A(n14641), .B(n22304), .Z(n14642) );
  NANDN U20089 ( .A(n22307), .B(n14642), .Z(n14645) );
  NANDN U20090 ( .A(x[1235]), .B(y[1235]), .Z(n14643) );
  NANDN U20091 ( .A(n14644), .B(n14643), .Z(n22308) );
  ANDN U20092 ( .B(n14645), .A(n22308), .Z(n14646) );
  OR U20093 ( .A(n22311), .B(n14646), .Z(n14647) );
  NANDN U20094 ( .A(n22313), .B(n14647), .Z(n14648) );
  NAND U20095 ( .A(n14648), .B(n22314), .Z(n14649) );
  NANDN U20096 ( .A(n22317), .B(n14649), .Z(n14650) );
  NAND U20097 ( .A(n14650), .B(n22318), .Z(n14651) );
  AND U20098 ( .A(n22321), .B(n14651), .Z(n14652) );
  OR U20099 ( .A(n22323), .B(n14652), .Z(n14653) );
  NANDN U20100 ( .A(n22325), .B(n14653), .Z(n14654) );
  NANDN U20101 ( .A(n22327), .B(n14654), .Z(n14655) );
  NANDN U20102 ( .A(n22329), .B(n14655), .Z(n14656) );
  NAND U20103 ( .A(n14656), .B(n22330), .Z(n14657) );
  ANDN U20104 ( .B(n14657), .A(n22332), .Z(n14658) );
  NANDN U20105 ( .A(n14658), .B(n22334), .Z(n14659) );
  NANDN U20106 ( .A(n22337), .B(n14659), .Z(n14660) );
  NAND U20107 ( .A(n14660), .B(n22338), .Z(n14661) );
  NANDN U20108 ( .A(n22341), .B(n14661), .Z(n14662) );
  NAND U20109 ( .A(n14662), .B(n22342), .Z(n14664) );
  NAND U20110 ( .A(n14664), .B(n14663), .Z(n14665) );
  NANDN U20111 ( .A(n14665), .B(n22345), .Z(n14666) );
  AND U20112 ( .A(n14667), .B(n14666), .Z(n14670) );
  NOR U20113 ( .A(n22352), .B(n14668), .Z(n14669) );
  NANDN U20114 ( .A(n14670), .B(n14669), .Z(n14671) );
  NANDN U20115 ( .A(n22355), .B(n14671), .Z(n14674) );
  NANDN U20116 ( .A(x[1259]), .B(y[1259]), .Z(n14672) );
  NANDN U20117 ( .A(n14673), .B(n14672), .Z(n22357) );
  ANDN U20118 ( .B(n14674), .A(n22357), .Z(n14675) );
  OR U20119 ( .A(n22359), .B(n14675), .Z(n14676) );
  NANDN U20120 ( .A(n22361), .B(n14676), .Z(n14677) );
  NAND U20121 ( .A(n14677), .B(n22362), .Z(n14678) );
  NANDN U20122 ( .A(n22364), .B(n14678), .Z(n14679) );
  NAND U20123 ( .A(n14679), .B(n22366), .Z(n14682) );
  OR U20124 ( .A(n14681), .B(n14680), .Z(n22369) );
  ANDN U20125 ( .B(n14682), .A(n22369), .Z(n14683) );
  OR U20126 ( .A(n22371), .B(n14683), .Z(n14686) );
  ANDN U20127 ( .B(n22372), .A(n14684), .Z(n14685) );
  NAND U20128 ( .A(n14686), .B(n14685), .Z(n14687) );
  NANDN U20129 ( .A(n14688), .B(n14687), .Z(n14689) );
  NAND U20130 ( .A(n14690), .B(n14689), .Z(n14691) );
  NANDN U20131 ( .A(n22382), .B(n14691), .Z(n14695) );
  NAND U20132 ( .A(n14692), .B(y[1271]), .Z(n14693) );
  NANDN U20133 ( .A(n14694), .B(n14693), .Z(n22385) );
  ANDN U20134 ( .B(n14695), .A(n22385), .Z(n14696) );
  OR U20135 ( .A(n22387), .B(n14696), .Z(n14697) );
  NANDN U20136 ( .A(n22388), .B(n14697), .Z(n14698) );
  NAND U20137 ( .A(n14698), .B(n22390), .Z(n14699) );
  NANDN U20138 ( .A(n22392), .B(n14699), .Z(n14700) );
  NAND U20139 ( .A(n14700), .B(n22394), .Z(n14703) );
  NANDN U20140 ( .A(n14702), .B(n14701), .Z(n22396) );
  ANDN U20141 ( .B(n14703), .A(n22396), .Z(n14704) );
  OR U20142 ( .A(n14704), .B(n22399), .Z(n14707) );
  NANDN U20143 ( .A(x[1279]), .B(y[1279]), .Z(n14705) );
  NANDN U20144 ( .A(n14706), .B(n14705), .Z(n22400) );
  ANDN U20145 ( .B(n14707), .A(n22400), .Z(n14708) );
  OR U20146 ( .A(n22403), .B(n14708), .Z(n14709) );
  NAND U20147 ( .A(n14709), .B(n22404), .Z(n14710) );
  NANDN U20148 ( .A(n22407), .B(n14710), .Z(n14711) );
  NANDN U20149 ( .A(n22408), .B(n14711), .Z(n14712) );
  AND U20150 ( .A(n22410), .B(n14712), .Z(n14715) );
  NANDN U20151 ( .A(x[1285]), .B(y[1285]), .Z(n14713) );
  NANDN U20152 ( .A(n14714), .B(n14713), .Z(n22413) );
  OR U20153 ( .A(n14715), .B(n22413), .Z(n14716) );
  AND U20154 ( .A(n22414), .B(n14716), .Z(n14717) );
  OR U20155 ( .A(n22417), .B(n14717), .Z(n14718) );
  NANDN U20156 ( .A(n22419), .B(n14718), .Z(n14719) );
  NANDN U20157 ( .A(n22421), .B(n14719), .Z(n14720) );
  NANDN U20158 ( .A(n22422), .B(n14720), .Z(n14722) );
  ANDN U20159 ( .B(n14722), .A(n14721), .Z(n14723) );
  NAND U20160 ( .A(n14723), .B(n22424), .Z(n14724) );
  AND U20161 ( .A(n22426), .B(n14724), .Z(n14725) );
  NAND U20162 ( .A(n14725), .B(n22430), .Z(n14726) );
  NAND U20163 ( .A(n14727), .B(n14726), .Z(n14728) );
  NANDN U20164 ( .A(n22434), .B(n14728), .Z(n14729) );
  NAND U20165 ( .A(n14729), .B(n22436), .Z(n14730) );
  NAND U20166 ( .A(n14730), .B(n22439), .Z(n14731) );
  AND U20167 ( .A(n22440), .B(n14731), .Z(n14732) );
  NANDN U20168 ( .A(n14732), .B(n22443), .Z(n14733) );
  AND U20169 ( .A(n22444), .B(n14733), .Z(n14734) );
  NANDN U20170 ( .A(n14734), .B(n22446), .Z(n14737) );
  OR U20171 ( .A(n14736), .B(n14735), .Z(n22449) );
  ANDN U20172 ( .B(n14737), .A(n22449), .Z(n14738) );
  NANDN U20173 ( .A(n14738), .B(n22450), .Z(n14739) );
  NANDN U20174 ( .A(n22452), .B(n14739), .Z(n14740) );
  NANDN U20175 ( .A(n22455), .B(n14740), .Z(n14741) );
  NAND U20176 ( .A(n14741), .B(n22456), .Z(n14742) );
  NANDN U20177 ( .A(n22459), .B(n14742), .Z(n14745) );
  NAND U20178 ( .A(n14744), .B(n14743), .Z(n22460) );
  ANDN U20179 ( .B(n14745), .A(n22460), .Z(n14746) );
  ANDN U20180 ( .B(n22462), .A(n14746), .Z(n14747) );
  NANDN U20181 ( .A(n14747), .B(n22465), .Z(n14748) );
  NAND U20182 ( .A(n14748), .B(n22466), .Z(n14749) );
  NAND U20183 ( .A(n14749), .B(n22468), .Z(n14750) );
  NAND U20184 ( .A(n14750), .B(n22470), .Z(n14751) );
  AND U20185 ( .A(n22472), .B(n14751), .Z(n14752) );
  NANDN U20186 ( .A(n14752), .B(n22475), .Z(n14753) );
  NAND U20187 ( .A(n14754), .B(n14753), .Z(n14755) );
  NAND U20188 ( .A(n14756), .B(n14755), .Z(n14757) );
  NAND U20189 ( .A(n14757), .B(n22484), .Z(n14759) );
  NANDN U20190 ( .A(n14759), .B(n14758), .Z(n14760) );
  AND U20191 ( .A(n22486), .B(n14760), .Z(n14761) );
  OR U20192 ( .A(n22489), .B(n14761), .Z(n14762) );
  AND U20193 ( .A(n22490), .B(n14762), .Z(n14763) );
  OR U20194 ( .A(n22492), .B(n14763), .Z(n14764) );
  NANDN U20195 ( .A(n22494), .B(n14764), .Z(n14765) );
  NAND U20196 ( .A(n14765), .B(n22496), .Z(n14766) );
  ANDN U20197 ( .B(n14766), .A(n22499), .Z(n14769) );
  NOR U20198 ( .A(n14768), .B(n14767), .Z(n22500) );
  NANDN U20199 ( .A(n14769), .B(n22500), .Z(n14770) );
  AND U20200 ( .A(n22502), .B(n14770), .Z(n14771) );
  OR U20201 ( .A(n14772), .B(n14771), .Z(n14775) );
  ANDN U20202 ( .B(n20287), .A(n14773), .Z(n14774) );
  NAND U20203 ( .A(n14775), .B(n14774), .Z(n14776) );
  NANDN U20204 ( .A(n22511), .B(n14776), .Z(n14777) );
  AND U20205 ( .A(n22512), .B(n14777), .Z(n14780) );
  NANDN U20206 ( .A(x[1331]), .B(y[1331]), .Z(n14778) );
  NANDN U20207 ( .A(n14779), .B(n14778), .Z(n22514) );
  OR U20208 ( .A(n14780), .B(n22514), .Z(n14781) );
  AND U20209 ( .A(n22516), .B(n14781), .Z(n14782) );
  OR U20210 ( .A(n22518), .B(n14782), .Z(n14783) );
  NAND U20211 ( .A(n14783), .B(n22520), .Z(n14784) );
  NANDN U20212 ( .A(n22522), .B(n14784), .Z(n14785) );
  NAND U20213 ( .A(n14785), .B(n22524), .Z(n14788) );
  OR U20214 ( .A(n14787), .B(n14786), .Z(n22526) );
  ANDN U20215 ( .B(n14788), .A(n22526), .Z(n14789) );
  NANDN U20216 ( .A(n14789), .B(n22528), .Z(n14790) );
  NAND U20217 ( .A(n14791), .B(n14790), .Z(n14795) );
  OR U20218 ( .A(n14792), .B(n22535), .Z(n22533) );
  NAND U20219 ( .A(n14793), .B(n22533), .Z(n14794) );
  AND U20220 ( .A(n14795), .B(n14794), .Z(n14796) );
  NANDN U20221 ( .A(n14796), .B(n22538), .Z(n14797) );
  NANDN U20222 ( .A(n22541), .B(n14797), .Z(n14798) );
  NANDN U20223 ( .A(n22543), .B(n14798), .Z(n14801) );
  ANDN U20224 ( .B(n14800), .A(n14799), .Z(n22544) );
  NAND U20225 ( .A(n14801), .B(n22544), .Z(n14802) );
  NANDN U20226 ( .A(n22547), .B(n14802), .Z(n14803) );
  AND U20227 ( .A(n22548), .B(n14803), .Z(n14804) );
  NANDN U20228 ( .A(n14804), .B(n22551), .Z(n14805) );
  NAND U20229 ( .A(n14805), .B(n22552), .Z(n14806) );
  NANDN U20230 ( .A(n22554), .B(n14806), .Z(n14807) );
  NANDN U20231 ( .A(n22557), .B(n14807), .Z(n14808) );
  NANDN U20232 ( .A(n22559), .B(n14808), .Z(n14809) );
  AND U20233 ( .A(n22560), .B(n14809), .Z(n14812) );
  NANDN U20234 ( .A(x[1355]), .B(y[1355]), .Z(n14810) );
  NANDN U20235 ( .A(n14811), .B(n14810), .Z(n22563) );
  OR U20236 ( .A(n14812), .B(n22563), .Z(n14813) );
  AND U20237 ( .A(n22564), .B(n14813), .Z(n14814) );
  OR U20238 ( .A(n14814), .B(n22566), .Z(n14815) );
  AND U20239 ( .A(n22568), .B(n14815), .Z(n14816) );
  OR U20240 ( .A(n22570), .B(n14816), .Z(n14817) );
  NAND U20241 ( .A(n14817), .B(n22572), .Z(n14818) );
  NANDN U20242 ( .A(n22575), .B(n14818), .Z(n14819) );
  NAND U20243 ( .A(n14819), .B(n22576), .Z(n14820) );
  AND U20244 ( .A(n14821), .B(n14820), .Z(n14822) );
  ANDN U20245 ( .B(n22584), .A(n14822), .Z(n14823) );
  NAND U20246 ( .A(n14823), .B(n22580), .Z(n14824) );
  AND U20247 ( .A(n22586), .B(n14824), .Z(n14825) );
  NANDN U20248 ( .A(n14826), .B(n14825), .Z(n14833) );
  NANDN U20249 ( .A(n14828), .B(n14827), .Z(n14829) );
  NANDN U20250 ( .A(n14830), .B(n14829), .Z(n14832) );
  ANDN U20251 ( .B(n14832), .A(n14831), .Z(n22588) );
  NAND U20252 ( .A(n14833), .B(n22588), .Z(n14834) );
  AND U20253 ( .A(n22590), .B(n14834), .Z(n14835) );
  OR U20254 ( .A(n22593), .B(n14835), .Z(n14836) );
  NAND U20255 ( .A(n14836), .B(n22594), .Z(n14837) );
  NANDN U20256 ( .A(n22597), .B(n14837), .Z(n14838) );
  NAND U20257 ( .A(n14838), .B(n22598), .Z(n14839) );
  NANDN U20258 ( .A(n22600), .B(n14839), .Z(n14840) );
  NANDN U20259 ( .A(n22603), .B(n14840), .Z(n14841) );
  NANDN U20260 ( .A(n22605), .B(n14841), .Z(n14842) );
  NANDN U20261 ( .A(n22607), .B(n14842), .Z(n14845) );
  NANDN U20262 ( .A(y[1380]), .B(x[1380]), .Z(n14843) );
  NANDN U20263 ( .A(n14844), .B(n14843), .Z(n22608) );
  ANDN U20264 ( .B(n14845), .A(n22608), .Z(n14846) );
  NANDN U20265 ( .A(n14846), .B(n22610), .Z(n14847) );
  NANDN U20266 ( .A(n22613), .B(n14847), .Z(n14848) );
  NAND U20267 ( .A(n14848), .B(n22614), .Z(n14849) );
  NAND U20268 ( .A(n14849), .B(n22616), .Z(n14850) );
  AND U20269 ( .A(n22619), .B(n14850), .Z(n14851) );
  OR U20270 ( .A(n14851), .B(n22621), .Z(n14852) );
  NANDN U20271 ( .A(n22623), .B(n14852), .Z(n14855) );
  NANDN U20272 ( .A(y[1390]), .B(x[1390]), .Z(n14853) );
  NANDN U20273 ( .A(n14854), .B(n14853), .Z(n22624) );
  ANDN U20274 ( .B(n14855), .A(n22624), .Z(n14856) );
  OR U20275 ( .A(n22627), .B(n14856), .Z(n14857) );
  NANDN U20276 ( .A(n22629), .B(n14857), .Z(n14858) );
  NANDN U20277 ( .A(n22631), .B(n14858), .Z(n14859) );
  NANDN U20278 ( .A(n22633), .B(n14859), .Z(n14860) );
  NAND U20279 ( .A(n14860), .B(n22634), .Z(n14861) );
  NAND U20280 ( .A(n14861), .B(n22636), .Z(n14862) );
  NANDN U20281 ( .A(n14863), .B(n14862), .Z(n14864) );
  NANDN U20282 ( .A(n14865), .B(n14864), .Z(n14866) );
  NANDN U20283 ( .A(n14867), .B(n14866), .Z(n14868) );
  NANDN U20284 ( .A(n14868), .B(x[1400]), .Z(n14872) );
  XNOR U20285 ( .A(n14868), .B(x[1400]), .Z(n14869) );
  NAND U20286 ( .A(n14870), .B(n14869), .Z(n14871) );
  NAND U20287 ( .A(n14872), .B(n14871), .Z(n14873) );
  NANDN U20288 ( .A(n14873), .B(n22644), .Z(n14874) );
  AND U20289 ( .A(n14875), .B(n14874), .Z(n14876) );
  NAND U20290 ( .A(n14876), .B(n22646), .Z(n14877) );
  NANDN U20291 ( .A(n22649), .B(n14877), .Z(n14878) );
  AND U20292 ( .A(n22650), .B(n14878), .Z(n14879) );
  OR U20293 ( .A(n22652), .B(n14879), .Z(n14880) );
  NAND U20294 ( .A(n14880), .B(n22654), .Z(n14881) );
  NANDN U20295 ( .A(n22657), .B(n14881), .Z(n14882) );
  AND U20296 ( .A(n22658), .B(n14882), .Z(n14883) );
  OR U20297 ( .A(n14883), .B(n22661), .Z(n14884) );
  AND U20298 ( .A(n22662), .B(n14884), .Z(n14887) );
  NOR U20299 ( .A(n14886), .B(n14885), .Z(n22665) );
  NANDN U20300 ( .A(n14887), .B(n22665), .Z(n14892) );
  NANDN U20301 ( .A(n14889), .B(n14888), .Z(n14891) );
  ANDN U20302 ( .B(n14891), .A(n14890), .Z(n22666) );
  NAND U20303 ( .A(n14892), .B(n22666), .Z(n14893) );
  NANDN U20304 ( .A(n22669), .B(n14893), .Z(n14894) );
  NANDN U20305 ( .A(n22671), .B(n14894), .Z(n14897) );
  NANDN U20306 ( .A(n14896), .B(n14895), .Z(n22673) );
  ANDN U20307 ( .B(n14897), .A(n22673), .Z(n14898) );
  OR U20308 ( .A(n22675), .B(n14898), .Z(n14899) );
  NAND U20309 ( .A(n14899), .B(n22677), .Z(n14900) );
  NAND U20310 ( .A(n14900), .B(n22678), .Z(n14901) );
  NAND U20311 ( .A(n14901), .B(n22680), .Z(n14902) );
  NAND U20312 ( .A(n14902), .B(n22682), .Z(n14903) );
  NANDN U20313 ( .A(n22685), .B(n14903), .Z(n14904) );
  NAND U20314 ( .A(n14905), .B(n14904), .Z(n14906) );
  NANDN U20315 ( .A(n14907), .B(n14906), .Z(n14908) );
  NAND U20316 ( .A(n14909), .B(n14908), .Z(n14913) );
  NAND U20317 ( .A(n14910), .B(x[1427]), .Z(n14911) );
  NANDN U20318 ( .A(n14912), .B(n14911), .Z(n22696) );
  ANDN U20319 ( .B(n14913), .A(n22696), .Z(n14914) );
  OR U20320 ( .A(n22698), .B(n14914), .Z(n14915) );
  NANDN U20321 ( .A(n22700), .B(n14915), .Z(n14916) );
  NANDN U20322 ( .A(n22702), .B(n14916), .Z(n14917) );
  NAND U20323 ( .A(n14917), .B(n22705), .Z(n14918) );
  NAND U20324 ( .A(n14918), .B(n22706), .Z(n14919) );
  AND U20325 ( .A(n22708), .B(n14919), .Z(n14920) );
  NANDN U20326 ( .A(n14920), .B(n22710), .Z(n14921) );
  AND U20327 ( .A(n22712), .B(n14921), .Z(n14923) );
  NANDN U20328 ( .A(n14923), .B(n14922), .Z(n14924) );
  NAND U20329 ( .A(n14924), .B(n22716), .Z(n14925) );
  AND U20330 ( .A(n14926), .B(n14925), .Z(n14927) );
  NAND U20331 ( .A(n14927), .B(n22718), .Z(n14928) );
  NANDN U20332 ( .A(n22721), .B(n14928), .Z(n14931) );
  NAND U20333 ( .A(n14930), .B(n14929), .Z(n22722) );
  ANDN U20334 ( .B(n14931), .A(n22722), .Z(n14932) );
  OR U20335 ( .A(n22725), .B(n14932), .Z(n14933) );
  NANDN U20336 ( .A(n22727), .B(n14933), .Z(n14934) );
  NANDN U20337 ( .A(n22729), .B(n14934), .Z(n14935) );
  NAND U20338 ( .A(n14935), .B(n22730), .Z(n14936) );
  NANDN U20339 ( .A(n22733), .B(n14936), .Z(n14937) );
  NAND U20340 ( .A(n14937), .B(n22734), .Z(n14938) );
  NANDN U20341 ( .A(n22737), .B(n14938), .Z(n14939) );
  AND U20342 ( .A(n22738), .B(n14939), .Z(n14941) );
  NAND U20343 ( .A(n14941), .B(n14940), .Z(n14942) );
  NAND U20344 ( .A(n14943), .B(n14942), .Z(n14945) );
  NAND U20345 ( .A(n14945), .B(n14944), .Z(n14946) );
  NANDN U20346 ( .A(n14946), .B(n22746), .Z(n14947) );
  AND U20347 ( .A(n22748), .B(n14947), .Z(n14948) );
  OR U20348 ( .A(n22750), .B(n14948), .Z(n14949) );
  AND U20349 ( .A(n22752), .B(n14949), .Z(n14950) );
  OR U20350 ( .A(n22755), .B(n14950), .Z(n14951) );
  NAND U20351 ( .A(n14951), .B(n22756), .Z(n14952) );
  NANDN U20352 ( .A(n22759), .B(n14952), .Z(n14953) );
  AND U20353 ( .A(n22760), .B(n14953), .Z(n14956) );
  NOR U20354 ( .A(n14955), .B(n14954), .Z(n22763) );
  NANDN U20355 ( .A(n14956), .B(n22763), .Z(n14957) );
  AND U20356 ( .A(n22764), .B(n14957), .Z(n14960) );
  NAND U20357 ( .A(n14958), .B(n22766), .Z(n14959) );
  OR U20358 ( .A(n14960), .B(n14959), .Z(n14961) );
  AND U20359 ( .A(n22768), .B(n14961), .Z(n14964) );
  OR U20360 ( .A(n14962), .B(n22775), .Z(n14963) );
  OR U20361 ( .A(n14964), .B(n14963), .Z(n14967) );
  OR U20362 ( .A(n14966), .B(n14965), .Z(n22777) );
  ANDN U20363 ( .B(n14967), .A(n22777), .Z(n14968) );
  NANDN U20364 ( .A(n14968), .B(n22778), .Z(n14969) );
  NAND U20365 ( .A(n14969), .B(n22781), .Z(n14970) );
  NAND U20366 ( .A(n14970), .B(n22782), .Z(n14971) );
  NANDN U20367 ( .A(n22784), .B(n14971), .Z(n14972) );
  NAND U20368 ( .A(n14972), .B(n22786), .Z(n14973) );
  NANDN U20369 ( .A(n22789), .B(n14973), .Z(n14977) );
  NAND U20370 ( .A(n14974), .B(y[1470]), .Z(n14976) );
  ANDN U20371 ( .B(n14976), .A(n14975), .Z(n22790) );
  NAND U20372 ( .A(n14977), .B(n22790), .Z(n14978) );
  NANDN U20373 ( .A(n22793), .B(n14978), .Z(n14980) );
  ANDN U20374 ( .B(n14980), .A(n14979), .Z(n14981) );
  NAND U20375 ( .A(n14981), .B(n22794), .Z(n14982) );
  NANDN U20376 ( .A(n14983), .B(n14982), .Z(n14984) );
  AND U20377 ( .A(n22803), .B(n14984), .Z(n14985) );
  OR U20378 ( .A(n22806), .B(n14985), .Z(n14988) );
  NANDN U20379 ( .A(x[1475]), .B(y[1475]), .Z(n14987) );
  ANDN U20380 ( .B(n14987), .A(n14986), .Z(n22808) );
  NAND U20381 ( .A(n14988), .B(n22808), .Z(n14989) );
  NANDN U20382 ( .A(n22810), .B(n14989), .Z(n14990) );
  NANDN U20383 ( .A(n22812), .B(n14990), .Z(n14991) );
  NAND U20384 ( .A(n14991), .B(n22813), .Z(n14992) );
  ANDN U20385 ( .B(n14992), .A(n22816), .Z(n14993) );
  OR U20386 ( .A(n22818), .B(n14993), .Z(n14997) );
  NAND U20387 ( .A(n14994), .B(y[1482]), .Z(n14996) );
  ANDN U20388 ( .B(n14996), .A(n14995), .Z(n22819) );
  NAND U20389 ( .A(n14997), .B(n22819), .Z(n14998) );
  NANDN U20390 ( .A(n22821), .B(n14998), .Z(n14999) );
  NAND U20391 ( .A(n15000), .B(n14999), .Z(n15001) );
  NAND U20392 ( .A(n15001), .B(n22825), .Z(n15002) );
  NANDN U20393 ( .A(n15002), .B(n22829), .Z(n15004) );
  ANDN U20394 ( .B(n15004), .A(n15003), .Z(n15005) );
  NAND U20395 ( .A(n15005), .B(n22831), .Z(n15006) );
  NANDN U20396 ( .A(n22833), .B(n15006), .Z(n15007) );
  NANDN U20397 ( .A(n22836), .B(n15007), .Z(n15008) );
  NANDN U20398 ( .A(n22838), .B(n15008), .Z(n15009) );
  NANDN U20399 ( .A(n22840), .B(n15009), .Z(n15012) );
  NANDN U20400 ( .A(y[1490]), .B(x[1490]), .Z(n15010) );
  NANDN U20401 ( .A(n15011), .B(n15010), .Z(n22842) );
  ANDN U20402 ( .B(n15012), .A(n22842), .Z(n15013) );
  NANDN U20403 ( .A(n15013), .B(n22843), .Z(n15014) );
  ANDN U20404 ( .B(n15014), .A(n22845), .Z(n15015) );
  NANDN U20405 ( .A(n15015), .B(n22847), .Z(n15016) );
  ANDN U20406 ( .B(n15016), .A(n22849), .Z(n15019) );
  NANDN U20407 ( .A(n15017), .B(n22852), .Z(n15018) );
  OR U20408 ( .A(n15019), .B(n15018), .Z(n15020) );
  AND U20409 ( .A(n15021), .B(n15020), .Z(n15024) );
  OR U20410 ( .A(n15022), .B(n22860), .Z(n15023) );
  OR U20411 ( .A(n15024), .B(n15023), .Z(n15025) );
  AND U20412 ( .A(n22861), .B(n15025), .Z(n15026) );
  OR U20413 ( .A(n22863), .B(n15026), .Z(n15027) );
  NANDN U20414 ( .A(n22866), .B(n15027), .Z(n15028) );
  NAND U20415 ( .A(n15028), .B(n22867), .Z(n15029) );
  NAND U20416 ( .A(n15029), .B(n22870), .Z(n15030) );
  NAND U20417 ( .A(n15030), .B(n22871), .Z(n15031) );
  NAND U20418 ( .A(n15031), .B(n22873), .Z(n15032) );
  NANDN U20419 ( .A(n15033), .B(n15032), .Z(n15034) );
  NAND U20420 ( .A(n15035), .B(n15034), .Z(n15036) );
  AND U20421 ( .A(n15037), .B(n15036), .Z(n15038) );
  NANDN U20422 ( .A(n20283), .B(n15038), .Z(n15039) );
  NANDN U20423 ( .A(n20284), .B(n15039), .Z(n15041) );
  NAND U20424 ( .A(n15041), .B(n15040), .Z(n15045) );
  NAND U20425 ( .A(n15042), .B(x[1511]), .Z(n15043) );
  NANDN U20426 ( .A(n15044), .B(n15043), .Z(n22882) );
  ANDN U20427 ( .B(n15045), .A(n22882), .Z(n15046) );
  NOR U20428 ( .A(n22884), .B(n15046), .Z(n15047) );
  NANDN U20429 ( .A(n15047), .B(n22886), .Z(n15048) );
  NAND U20430 ( .A(n15048), .B(n22887), .Z(n15049) );
  NAND U20431 ( .A(n15049), .B(n22890), .Z(n15050) );
  NAND U20432 ( .A(n15050), .B(n22891), .Z(n15051) );
  NAND U20433 ( .A(n15051), .B(n22894), .Z(n15052) );
  NANDN U20434 ( .A(n22896), .B(n15052), .Z(n15055) );
  NANDN U20435 ( .A(y[1518]), .B(x[1518]), .Z(n15053) );
  NANDN U20436 ( .A(n15054), .B(n15053), .Z(n22898) );
  ANDN U20437 ( .B(n15055), .A(n22898), .Z(n15058) );
  NANDN U20438 ( .A(n15056), .B(n22899), .Z(n15057) );
  OR U20439 ( .A(n15058), .B(n15057), .Z(n15059) );
  ANDN U20440 ( .B(n15059), .A(n22902), .Z(n15061) );
  NANDN U20441 ( .A(n15061), .B(n15060), .Z(n15062) );
  AND U20442 ( .A(n22906), .B(n15062), .Z(n15063) );
  NANDN U20443 ( .A(n15063), .B(n22907), .Z(n15064) );
  AND U20444 ( .A(n22910), .B(n15064), .Z(n15065) );
  NANDN U20445 ( .A(n15065), .B(n22911), .Z(n15066) );
  NAND U20446 ( .A(n15066), .B(n22914), .Z(n15067) );
  AND U20447 ( .A(n22915), .B(n15067), .Z(n15068) );
  NANDN U20448 ( .A(n15068), .B(n22917), .Z(n15071) );
  NANDN U20449 ( .A(x[1530]), .B(y[1530]), .Z(n15070) );
  ANDN U20450 ( .B(n15070), .A(n15069), .Z(n22919) );
  NAND U20451 ( .A(n15071), .B(n22919), .Z(n15072) );
  NANDN U20452 ( .A(n22922), .B(n15072), .Z(n15073) );
  NAND U20453 ( .A(n15074), .B(n15073), .Z(n15075) );
  AND U20454 ( .A(n15076), .B(n15075), .Z(n15077) );
  ANDN U20455 ( .B(n22932), .A(n15077), .Z(n15079) );
  NAND U20456 ( .A(n15079), .B(n15078), .Z(n15080) );
  AND U20457 ( .A(n22933), .B(n15080), .Z(n15081) );
  NANDN U20458 ( .A(n15081), .B(n22936), .Z(n15082) );
  NAND U20459 ( .A(n15082), .B(n22937), .Z(n15083) );
  NAND U20460 ( .A(n15083), .B(n22939), .Z(n15084) );
  AND U20461 ( .A(n22941), .B(n15084), .Z(n15085) );
  OR U20462 ( .A(n22944), .B(n15085), .Z(n15088) );
  OR U20463 ( .A(n15087), .B(n15086), .Z(n22945) );
  ANDN U20464 ( .B(n15088), .A(n22945), .Z(n15089) );
  OR U20465 ( .A(n15090), .B(n15089), .Z(n15093) );
  ANDN U20466 ( .B(n20281), .A(n15091), .Z(n15092) );
  NAND U20467 ( .A(n15093), .B(n15092), .Z(n15094) );
  NANDN U20468 ( .A(n22954), .B(n15094), .Z(n15097) );
  AND U20469 ( .A(n15096), .B(n15095), .Z(n22955) );
  NAND U20470 ( .A(n15097), .B(n22955), .Z(n15098) );
  NANDN U20471 ( .A(n22957), .B(n15098), .Z(n15099) );
  AND U20472 ( .A(n22959), .B(n15099), .Z(n15100) );
  OR U20473 ( .A(n22961), .B(n15100), .Z(n15101) );
  NAND U20474 ( .A(n15101), .B(n22963), .Z(n15102) );
  AND U20475 ( .A(n22965), .B(n15102), .Z(n15103) );
  NANDN U20476 ( .A(n15103), .B(n22967), .Z(n15107) );
  NAND U20477 ( .A(n15104), .B(y[1554]), .Z(n15106) );
  ANDN U20478 ( .B(n15106), .A(n15105), .Z(n22969) );
  NAND U20479 ( .A(n15107), .B(n22969), .Z(n15108) );
  NANDN U20480 ( .A(n22971), .B(n15108), .Z(n15109) );
  NAND U20481 ( .A(n15110), .B(n15109), .Z(n15111) );
  NANDN U20482 ( .A(n15112), .B(n15111), .Z(n15113) );
  AND U20483 ( .A(n22981), .B(n15113), .Z(n15114) );
  OR U20484 ( .A(n22984), .B(n15114), .Z(n15117) );
  AND U20485 ( .A(n15116), .B(n15115), .Z(n22985) );
  NAND U20486 ( .A(n15117), .B(n22985), .Z(n15118) );
  NANDN U20487 ( .A(n22988), .B(n15118), .Z(n15119) );
  NAND U20488 ( .A(n15119), .B(n22989), .Z(n15120) );
  NAND U20489 ( .A(n15120), .B(n22991), .Z(n15121) );
  AND U20490 ( .A(n22993), .B(n15121), .Z(n15122) );
  NANDN U20491 ( .A(n15122), .B(n22995), .Z(n15123) );
  NANDN U20492 ( .A(n22997), .B(n15123), .Z(n15124) );
  NAND U20493 ( .A(n15124), .B(n22999), .Z(n15125) );
  NAND U20494 ( .A(n15126), .B(n15125), .Z(n15127) );
  NAND U20495 ( .A(n15127), .B(n23003), .Z(n15128) );
  NANDN U20496 ( .A(n15128), .B(n23007), .Z(n15129) );
  AND U20497 ( .A(n23010), .B(n15129), .Z(n15131) );
  NAND U20498 ( .A(n15131), .B(n15130), .Z(n15132) );
  AND U20499 ( .A(n23011), .B(n15132), .Z(n15133) );
  NANDN U20500 ( .A(n15133), .B(n23014), .Z(n15134) );
  AND U20501 ( .A(n23015), .B(n15134), .Z(n15135) );
  NANDN U20502 ( .A(n15135), .B(n23018), .Z(n15136) );
  NAND U20503 ( .A(n15136), .B(n23019), .Z(n15137) );
  NAND U20504 ( .A(n15137), .B(n23022), .Z(n15140) );
  NOR U20505 ( .A(n15139), .B(n15138), .Z(n23023) );
  NAND U20506 ( .A(n15140), .B(n23023), .Z(n15141) );
  NANDN U20507 ( .A(n23025), .B(n15141), .Z(n15142) );
  NANDN U20508 ( .A(n23028), .B(n15142), .Z(n15143) );
  AND U20509 ( .A(n23029), .B(n15143), .Z(n15144) );
  OR U20510 ( .A(n23032), .B(n15144), .Z(n15147) );
  NANDN U20511 ( .A(x[1583]), .B(y[1583]), .Z(n15145) );
  NANDN U20512 ( .A(n15146), .B(n15145), .Z(n23034) );
  ANDN U20513 ( .B(n15147), .A(n23034), .Z(n15148) );
  NANDN U20514 ( .A(n15148), .B(n23035), .Z(n15149) );
  ANDN U20515 ( .B(n15149), .A(n23037), .Z(n15150) );
  NANDN U20516 ( .A(n15150), .B(n23039), .Z(n15151) );
  NANDN U20517 ( .A(n23042), .B(n15151), .Z(n15152) );
  NAND U20518 ( .A(n15152), .B(n23043), .Z(n15155) );
  NANDN U20519 ( .A(n15154), .B(n15153), .Z(n23046) );
  ANDN U20520 ( .B(n15155), .A(n23046), .Z(n15156) );
  NANDN U20521 ( .A(n15156), .B(n23047), .Z(n15159) );
  ANDN U20522 ( .B(n23049), .A(n15157), .Z(n15158) );
  NAND U20523 ( .A(n15159), .B(n15158), .Z(n15160) );
  NANDN U20524 ( .A(n15161), .B(n15160), .Z(n15162) );
  NAND U20525 ( .A(n15163), .B(n15162), .Z(n15164) );
  NANDN U20526 ( .A(n23059), .B(n15164), .Z(n15165) );
  NANDN U20527 ( .A(n23061), .B(n15165), .Z(n15169) );
  NAND U20528 ( .A(n15166), .B(x[1596]), .Z(n15167) );
  NANDN U20529 ( .A(n15168), .B(n15167), .Z(n23063) );
  ANDN U20530 ( .B(n15169), .A(n23063), .Z(n15170) );
  NANDN U20531 ( .A(n15170), .B(n23065), .Z(n15171) );
  NAND U20532 ( .A(n15171), .B(n23067), .Z(n15172) );
  NAND U20533 ( .A(n15172), .B(n23069), .Z(n15173) );
  NAND U20534 ( .A(n15173), .B(n23071), .Z(n15174) );
  NAND U20535 ( .A(n15174), .B(n23073), .Z(n15175) );
  NAND U20536 ( .A(n15175), .B(n23076), .Z(n15176) );
  NAND U20537 ( .A(n15176), .B(n23077), .Z(n15177) );
  NAND U20538 ( .A(n15177), .B(n23079), .Z(n15178) );
  AND U20539 ( .A(n23081), .B(n15178), .Z(n15179) );
  OR U20540 ( .A(n23084), .B(n15179), .Z(n15182) );
  AND U20541 ( .A(n15181), .B(n15180), .Z(n23085) );
  NAND U20542 ( .A(n15182), .B(n23085), .Z(n15183) );
  NANDN U20543 ( .A(n23087), .B(n15183), .Z(n15184) );
  NAND U20544 ( .A(n15185), .B(n15184), .Z(n15186) );
  NAND U20545 ( .A(n15186), .B(n23091), .Z(n15188) );
  NANDN U20546 ( .A(n15188), .B(y[1611]), .Z(n15191) );
  XOR U20547 ( .A(n15188), .B(n15187), .Z(n15189) );
  NANDN U20548 ( .A(x[1611]), .B(n15189), .Z(n15190) );
  AND U20549 ( .A(n15191), .B(n15190), .Z(n15192) );
  NANDN U20550 ( .A(n15192), .B(n15193), .Z(n15196) );
  XNOR U20551 ( .A(n15193), .B(n15192), .Z(n15194) );
  NAND U20552 ( .A(n15194), .B(y[1612]), .Z(n15195) );
  NAND U20553 ( .A(n15196), .B(n15195), .Z(n15197) );
  AND U20554 ( .A(n23099), .B(n15197), .Z(n15200) );
  NAND U20555 ( .A(n15198), .B(n23101), .Z(n15199) );
  OR U20556 ( .A(n15200), .B(n15199), .Z(n15201) );
  AND U20557 ( .A(n23103), .B(n15201), .Z(n15202) );
  OR U20558 ( .A(n23106), .B(n15202), .Z(n15203) );
  NAND U20559 ( .A(n15203), .B(n23107), .Z(n15204) );
  NANDN U20560 ( .A(n23109), .B(n15204), .Z(n15205) );
  NAND U20561 ( .A(n15205), .B(n23111), .Z(n15206) );
  NANDN U20562 ( .A(n23114), .B(n15206), .Z(n15207) );
  AND U20563 ( .A(n23115), .B(n15207), .Z(n15208) );
  OR U20564 ( .A(n23118), .B(n15208), .Z(n15211) );
  ANDN U20565 ( .B(n15210), .A(n15209), .Z(n23119) );
  NAND U20566 ( .A(n15211), .B(n23119), .Z(n15213) );
  NAND U20567 ( .A(n15213), .B(n15212), .Z(n15215) );
  NAND U20568 ( .A(n15215), .B(n15214), .Z(n15216) );
  AND U20569 ( .A(n15217), .B(n15216), .Z(n15218) );
  NANDN U20570 ( .A(n15218), .B(n20279), .Z(n15219) );
  NAND U20571 ( .A(n15219), .B(n23133), .Z(n15220) );
  NAND U20572 ( .A(n15220), .B(n23136), .Z(n15221) );
  NAND U20573 ( .A(n15221), .B(n23138), .Z(n15222) );
  NANDN U20574 ( .A(n23141), .B(n15222), .Z(n15223) );
  AND U20575 ( .A(n23143), .B(n15223), .Z(n15224) );
  NANDN U20576 ( .A(n15224), .B(n23144), .Z(n15225) );
  AND U20577 ( .A(n15226), .B(n15225), .Z(n15227) );
  NANDN U20578 ( .A(n15227), .B(n23148), .Z(n15229) );
  ANDN U20579 ( .B(n15229), .A(n15228), .Z(n15230) );
  NANDN U20580 ( .A(n15230), .B(n23154), .Z(n15231) );
  NAND U20581 ( .A(n15231), .B(n20277), .Z(n15233) );
  NAND U20582 ( .A(n15233), .B(n15232), .Z(n15234) );
  NAND U20583 ( .A(n15235), .B(n15234), .Z(n15236) );
  NANDN U20584 ( .A(n23158), .B(n15236), .Z(n15238) );
  NANDN U20585 ( .A(n15238), .B(y[1639]), .Z(n15241) );
  XOR U20586 ( .A(n15238), .B(n15237), .Z(n15239) );
  NANDN U20587 ( .A(x[1639]), .B(n15239), .Z(n15240) );
  NAND U20588 ( .A(n15241), .B(n15240), .Z(n15242) );
  NANDN U20589 ( .A(n15242), .B(n23166), .Z(n15243) );
  AND U20590 ( .A(n23169), .B(n15243), .Z(n15245) );
  NAND U20591 ( .A(n15245), .B(n15244), .Z(n15246) );
  NANDN U20592 ( .A(n23171), .B(n15246), .Z(n15247) );
  ANDN U20593 ( .B(n15247), .A(n23173), .Z(n15248) );
  NANDN U20594 ( .A(n15248), .B(n23174), .Z(n15249) );
  NANDN U20595 ( .A(n15250), .B(n15249), .Z(n15252) );
  XNOR U20596 ( .A(y[1646]), .B(n15252), .Z(n15251) );
  NANDN U20597 ( .A(x[1646]), .B(n15251), .Z(n15254) );
  NANDN U20598 ( .A(n15252), .B(y[1646]), .Z(n15253) );
  AND U20599 ( .A(n15254), .B(n15253), .Z(n15255) );
  NANDN U20600 ( .A(n15255), .B(n23180), .Z(n15257) );
  ANDN U20601 ( .B(n15257), .A(n15256), .Z(n15258) );
  NAND U20602 ( .A(n15258), .B(n23182), .Z(n15261) );
  ANDN U20603 ( .B(n15260), .A(n15259), .Z(n23184) );
  NAND U20604 ( .A(n15261), .B(n23184), .Z(n15262) );
  NANDN U20605 ( .A(n23187), .B(n15262), .Z(n15265) );
  ANDN U20606 ( .B(n15264), .A(n15263), .Z(n23188) );
  NAND U20607 ( .A(n15265), .B(n23188), .Z(n15266) );
  NANDN U20608 ( .A(n23190), .B(n15266), .Z(n15268) );
  ANDN U20609 ( .B(n15268), .A(n15267), .Z(n15269) );
  NAND U20610 ( .A(n15269), .B(n23192), .Z(n15270) );
  NAND U20611 ( .A(n15270), .B(n23194), .Z(n15272) );
  ANDN U20612 ( .B(n15272), .A(n15271), .Z(n15273) );
  OR U20613 ( .A(n23199), .B(n15273), .Z(n15274) );
  NANDN U20614 ( .A(n23201), .B(n15274), .Z(n15276) );
  NAND U20615 ( .A(n15276), .B(n15275), .Z(n15277) );
  NANDN U20616 ( .A(n15278), .B(n15277), .Z(n15279) );
  AND U20617 ( .A(n15280), .B(n15279), .Z(n15281) );
  NAND U20618 ( .A(n15281), .B(n23208), .Z(n15282) );
  NANDN U20619 ( .A(n23213), .B(n15282), .Z(n15286) );
  NAND U20620 ( .A(n15284), .B(n15283), .Z(n15285) );
  NAND U20621 ( .A(n15286), .B(n15285), .Z(n15288) );
  NANDN U20622 ( .A(n15288), .B(n15287), .Z(n15290) );
  ANDN U20623 ( .B(n15290), .A(n15289), .Z(n15291) );
  OR U20624 ( .A(n15292), .B(n15291), .Z(n15295) );
  NANDN U20625 ( .A(x[1665]), .B(n15295), .Z(n15293) );
  AND U20626 ( .A(n15294), .B(n15293), .Z(n15298) );
  XNOR U20627 ( .A(x[1665]), .B(n15295), .Z(n15296) );
  NAND U20628 ( .A(n15296), .B(y[1665]), .Z(n15297) );
  NAND U20629 ( .A(n15298), .B(n15297), .Z(n15300) );
  ANDN U20630 ( .B(n15300), .A(n15299), .Z(n15301) );
  NAND U20631 ( .A(n15302), .B(n15301), .Z(n15303) );
  NAND U20632 ( .A(n15304), .B(n15303), .Z(n15305) );
  NAND U20633 ( .A(n15306), .B(n15305), .Z(n15307) );
  NANDN U20634 ( .A(n23227), .B(n15307), .Z(n15308) );
  NANDN U20635 ( .A(n23228), .B(n15308), .Z(n15309) );
  AND U20636 ( .A(n23230), .B(n15309), .Z(n15310) );
  ANDN U20637 ( .B(n23233), .A(n15310), .Z(n15312) );
  NAND U20638 ( .A(n15312), .B(n15311), .Z(n15313) );
  AND U20639 ( .A(n23234), .B(n15313), .Z(n15314) );
  NAND U20640 ( .A(n15315), .B(n15314), .Z(n15316) );
  NAND U20641 ( .A(n15317), .B(n15316), .Z(n15318) );
  NAND U20642 ( .A(n15319), .B(n15318), .Z(n15320) );
  NAND U20643 ( .A(n15321), .B(n15320), .Z(n15323) );
  NANDN U20644 ( .A(n15323), .B(n15322), .Z(n15324) );
  NANDN U20645 ( .A(n20271), .B(n15324), .Z(n15326) );
  XNOR U20646 ( .A(x[1678]), .B(n15326), .Z(n15325) );
  NANDN U20647 ( .A(y[1678]), .B(n15325), .Z(n15328) );
  NANDN U20648 ( .A(n15326), .B(x[1678]), .Z(n15327) );
  AND U20649 ( .A(n15328), .B(n15327), .Z(n15329) );
  NAND U20650 ( .A(n15330), .B(n15329), .Z(n15331) );
  NAND U20651 ( .A(n15332), .B(n15331), .Z(n15333) );
  NANDN U20652 ( .A(n15334), .B(n15333), .Z(n15335) );
  NANDN U20653 ( .A(y[1681]), .B(n15335), .Z(n15338) );
  XNOR U20654 ( .A(y[1681]), .B(n15335), .Z(n15336) );
  NAND U20655 ( .A(n15336), .B(x[1681]), .Z(n15337) );
  NAND U20656 ( .A(n15338), .B(n15337), .Z(n15339) );
  AND U20657 ( .A(n23254), .B(n15339), .Z(n15342) );
  OR U20658 ( .A(n15340), .B(n23256), .Z(n15341) );
  OR U20659 ( .A(n15342), .B(n15341), .Z(n15343) );
  AND U20660 ( .A(n23258), .B(n15343), .Z(n15344) );
  ANDN U20661 ( .B(n23261), .A(n15344), .Z(n15346) );
  NAND U20662 ( .A(n15346), .B(n15345), .Z(n15347) );
  AND U20663 ( .A(n23262), .B(n15347), .Z(n15348) );
  NAND U20664 ( .A(n15349), .B(n15348), .Z(n15350) );
  NAND U20665 ( .A(n15351), .B(n15350), .Z(n15353) );
  AND U20666 ( .A(n15353), .B(n15352), .Z(n15354) );
  OR U20667 ( .A(n15354), .B(x[1688]), .Z(n15357) );
  XOR U20668 ( .A(x[1688]), .B(n15354), .Z(n15355) );
  NAND U20669 ( .A(n15355), .B(y[1688]), .Z(n15356) );
  NAND U20670 ( .A(n15357), .B(n15356), .Z(n15358) );
  AND U20671 ( .A(n23272), .B(n15358), .Z(n15359) );
  OR U20672 ( .A(n15360), .B(n15359), .Z(n15363) );
  ANDN U20673 ( .B(n15362), .A(n15361), .Z(n23276) );
  NAND U20674 ( .A(n15363), .B(n23276), .Z(n15364) );
  NANDN U20675 ( .A(n23278), .B(n15364), .Z(n15365) );
  NAND U20676 ( .A(n15366), .B(n15365), .Z(n15368) );
  ANDN U20677 ( .B(n15368), .A(n15367), .Z(n15369) );
  OR U20678 ( .A(n15369), .B(x[1694]), .Z(n15372) );
  XOR U20679 ( .A(x[1694]), .B(n15369), .Z(n15370) );
  NAND U20680 ( .A(n15370), .B(y[1694]), .Z(n15371) );
  NAND U20681 ( .A(n15372), .B(n15371), .Z(n15373) );
  AND U20682 ( .A(n23288), .B(n15373), .Z(n15374) );
  ANDN U20683 ( .B(n15375), .A(n15374), .Z(n15379) );
  XNOR U20684 ( .A(y[1696]), .B(x[1696]), .Z(n15376) );
  NAND U20685 ( .A(n15377), .B(n15376), .Z(n15378) );
  NAND U20686 ( .A(n15379), .B(n15378), .Z(n15380) );
  NAND U20687 ( .A(n15381), .B(n15380), .Z(n15383) );
  AND U20688 ( .A(n15383), .B(n15382), .Z(n15384) );
  NAND U20689 ( .A(n15385), .B(n15384), .Z(n15386) );
  NAND U20690 ( .A(n15387), .B(n15386), .Z(n15389) );
  ANDN U20691 ( .B(n15389), .A(n15388), .Z(n15390) );
  NAND U20692 ( .A(n15391), .B(n15390), .Z(n15392) );
  NAND U20693 ( .A(n15393), .B(n15392), .Z(n15395) );
  ANDN U20694 ( .B(n15395), .A(n15394), .Z(n15396) );
  NANDN U20695 ( .A(n15396), .B(n23300), .Z(n15397) );
  AND U20696 ( .A(n15398), .B(n15397), .Z(n15399) );
  NANDN U20697 ( .A(n15399), .B(n23304), .Z(n15400) );
  AND U20698 ( .A(n15401), .B(n15400), .Z(n15402) );
  OR U20699 ( .A(n23309), .B(n15402), .Z(n15403) );
  NAND U20700 ( .A(n15403), .B(n23310), .Z(n15404) );
  NAND U20701 ( .A(n15404), .B(n23313), .Z(n15405) );
  NAND U20702 ( .A(n15405), .B(n23315), .Z(n15406) );
  NAND U20703 ( .A(n15406), .B(n23318), .Z(n15408) );
  ANDN U20704 ( .B(n15408), .A(n15407), .Z(n15409) );
  OR U20705 ( .A(n23323), .B(n15409), .Z(n15410) );
  NANDN U20706 ( .A(n23324), .B(n15410), .Z(n15411) );
  NANDN U20707 ( .A(n23327), .B(n15411), .Z(n15412) );
  NANDN U20708 ( .A(n23329), .B(n15412), .Z(n15413) );
  NAND U20709 ( .A(n15413), .B(n23330), .Z(n15414) );
  ANDN U20710 ( .B(n15414), .A(n23333), .Z(n15415) );
  NANDN U20711 ( .A(n15415), .B(n23334), .Z(n15416) );
  NAND U20712 ( .A(n15416), .B(n23337), .Z(n15417) );
  NANDN U20713 ( .A(n23338), .B(n15417), .Z(n15418) );
  NANDN U20714 ( .A(n23340), .B(n15418), .Z(n15420) );
  ANDN U20715 ( .B(n15420), .A(n15419), .Z(n15421) );
  NAND U20716 ( .A(n15421), .B(n23342), .Z(n15422) );
  AND U20717 ( .A(n23344), .B(n15422), .Z(n15423) );
  OR U20718 ( .A(n15424), .B(n15423), .Z(n15425) );
  ANDN U20719 ( .B(n15425), .A(n23349), .Z(n15426) );
  NANDN U20720 ( .A(n15426), .B(n23350), .Z(n15427) );
  ANDN U20721 ( .B(n15427), .A(n23352), .Z(n15428) );
  NANDN U20722 ( .A(n15428), .B(n23354), .Z(n15429) );
  NANDN U20723 ( .A(n23356), .B(n15429), .Z(n15430) );
  NAND U20724 ( .A(n15430), .B(n23358), .Z(n15431) );
  NAND U20725 ( .A(n15431), .B(n23360), .Z(n15433) );
  ANDN U20726 ( .B(n15433), .A(n15432), .Z(n15434) );
  NAND U20727 ( .A(n15435), .B(n15434), .Z(n15436) );
  AND U20728 ( .A(n23364), .B(n15436), .Z(n15437) );
  NANDN U20729 ( .A(n15437), .B(n23366), .Z(n15438) );
  AND U20730 ( .A(n23368), .B(n15438), .Z(n15439) );
  NANDN U20731 ( .A(n15439), .B(n23370), .Z(n15440) );
  NAND U20732 ( .A(n15440), .B(n23372), .Z(n15441) );
  NAND U20733 ( .A(n15441), .B(n23375), .Z(n15442) );
  NAND U20734 ( .A(n15442), .B(n23376), .Z(n15443) );
  AND U20735 ( .A(n23379), .B(n15443), .Z(n15444) );
  NANDN U20736 ( .A(n15444), .B(n23380), .Z(n15445) );
  AND U20737 ( .A(n23382), .B(n15445), .Z(n15450) );
  NANDN U20738 ( .A(n15447), .B(n15446), .Z(n15448) );
  NANDN U20739 ( .A(n15449), .B(n15448), .Z(n23384) );
  OR U20740 ( .A(n15450), .B(n23384), .Z(n15451) );
  NAND U20741 ( .A(n15451), .B(n23386), .Z(n15452) );
  ANDN U20742 ( .B(n15452), .A(n23388), .Z(n15453) );
  NANDN U20743 ( .A(n15453), .B(n23390), .Z(n15454) );
  AND U20744 ( .A(n23392), .B(n15454), .Z(n15455) );
  OR U20745 ( .A(n15456), .B(n15455), .Z(n15457) );
  NAND U20746 ( .A(n15458), .B(n15457), .Z(n15461) );
  XOR U20747 ( .A(n15458), .B(n15457), .Z(n15459) );
  NAND U20748 ( .A(n15459), .B(x[1746]), .Z(n15460) );
  NAND U20749 ( .A(n15461), .B(n15460), .Z(n15463) );
  ANDN U20750 ( .B(n15463), .A(n15462), .Z(n15464) );
  NANDN U20751 ( .A(n15464), .B(n23398), .Z(n15465) );
  AND U20752 ( .A(n23400), .B(n15465), .Z(n15467) );
  OR U20753 ( .A(n15467), .B(n15466), .Z(n15468) );
  NANDN U20754 ( .A(n15468), .B(y[1750]), .Z(n15472) );
  XNOR U20755 ( .A(n15468), .B(y[1750]), .Z(n15469) );
  NAND U20756 ( .A(n15470), .B(n15469), .Z(n15471) );
  NAND U20757 ( .A(n15472), .B(n15471), .Z(n15473) );
  NAND U20758 ( .A(n15474), .B(n15473), .Z(n15475) );
  NAND U20759 ( .A(n15476), .B(n15475), .Z(n15478) );
  ANDN U20760 ( .B(n15478), .A(n15477), .Z(n15479) );
  NAND U20761 ( .A(n15479), .B(n23410), .Z(n15480) );
  NAND U20762 ( .A(n15480), .B(n23413), .Z(n15482) );
  NANDN U20763 ( .A(n15482), .B(n15481), .Z(n15483) );
  NANDN U20764 ( .A(n23415), .B(n15483), .Z(n15484) );
  NANDN U20765 ( .A(n23417), .B(n15484), .Z(n15485) );
  NAND U20766 ( .A(n15485), .B(n23418), .Z(n15486) );
  NANDN U20767 ( .A(n23421), .B(n15486), .Z(n15487) );
  AND U20768 ( .A(n23422), .B(n15487), .Z(n15488) );
  NANDN U20769 ( .A(n15488), .B(n23425), .Z(n15491) );
  NOR U20770 ( .A(n15490), .B(n15489), .Z(n23426) );
  NAND U20771 ( .A(n15491), .B(n23426), .Z(n15492) );
  NANDN U20772 ( .A(n23429), .B(n15492), .Z(n15494) );
  ANDN U20773 ( .B(n15494), .A(n15493), .Z(n15495) );
  NAND U20774 ( .A(n15495), .B(n23430), .Z(n15497) );
  NAND U20775 ( .A(n15497), .B(n15496), .Z(n15498) );
  NANDN U20776 ( .A(n15498), .B(n23432), .Z(n15499) );
  AND U20777 ( .A(n23438), .B(n15499), .Z(n15502) );
  NAND U20778 ( .A(n15500), .B(x[1764]), .Z(n15501) );
  NAND U20779 ( .A(n15502), .B(n15501), .Z(n15503) );
  NAND U20780 ( .A(n15504), .B(n15503), .Z(n15505) );
  OR U20781 ( .A(n23440), .B(n15505), .Z(n15506) );
  AND U20782 ( .A(n23442), .B(n15506), .Z(n15507) );
  OR U20783 ( .A(n15507), .B(n23445), .Z(n15508) );
  AND U20784 ( .A(n23446), .B(n15508), .Z(n15509) );
  OR U20785 ( .A(n23449), .B(n15509), .Z(n15510) );
  NAND U20786 ( .A(n15510), .B(n23450), .Z(n15511) );
  NAND U20787 ( .A(n15511), .B(n23453), .Z(n15512) );
  NAND U20788 ( .A(n15512), .B(n23454), .Z(n15513) );
  AND U20789 ( .A(n23456), .B(n15513), .Z(n15514) );
  OR U20790 ( .A(n23459), .B(n15514), .Z(n15515) );
  NANDN U20791 ( .A(n23461), .B(n15515), .Z(n15517) );
  NAND U20792 ( .A(n15517), .B(n15516), .Z(n15518) );
  NAND U20793 ( .A(n15519), .B(n15518), .Z(n15522) );
  XOR U20794 ( .A(n15519), .B(n15518), .Z(n15520) );
  NAND U20795 ( .A(n15520), .B(x[1778]), .Z(n15521) );
  NAND U20796 ( .A(n15522), .B(n15521), .Z(n15523) );
  NANDN U20797 ( .A(n23500), .B(n15528), .Z(n15529) );
  NAND U20798 ( .A(n15529), .B(n23502), .Z(n15530) );
  NAND U20799 ( .A(n15530), .B(n23504), .Z(n15531) );
  NAND U20800 ( .A(n15531), .B(n23506), .Z(n15536) );
  NANDN U20801 ( .A(n15533), .B(n15532), .Z(n15534) );
  NANDN U20802 ( .A(n15535), .B(n15534), .Z(n23509) );
  ANDN U20803 ( .B(n15536), .A(n23509), .Z(n15537) );
  NANDN U20804 ( .A(n15537), .B(n23511), .Z(n15538) );
  ANDN U20805 ( .B(n15538), .A(n23515), .Z(n15539) );
  OR U20806 ( .A(n15540), .B(n15539), .Z(n15541) );
  NAND U20807 ( .A(n15541), .B(n23519), .Z(n15542) );
  AND U20808 ( .A(n23520), .B(n15542), .Z(n15543) );
  NANDN U20809 ( .A(n15543), .B(n23522), .Z(n15546) );
  NOR U20810 ( .A(n15545), .B(n15544), .Z(n23524) );
  NAND U20811 ( .A(n15546), .B(n23524), .Z(n15547) );
  NANDN U20812 ( .A(n23527), .B(n15547), .Z(n15548) );
  NAND U20813 ( .A(n15549), .B(n15548), .Z(n15550) );
  NANDN U20814 ( .A(n23530), .B(n15550), .Z(n15551) );
  NANDN U20815 ( .A(n15551), .B(x[1806]), .Z(n15554) );
  XNOR U20816 ( .A(n15551), .B(x[1806]), .Z(n15552) );
  NANDN U20817 ( .A(y[1806]), .B(n15552), .Z(n15553) );
  AND U20818 ( .A(n15554), .B(n15553), .Z(n15556) );
  NANDN U20819 ( .A(x[1807]), .B(n15556), .Z(n15555) );
  AND U20820 ( .A(n23538), .B(n15555), .Z(n15559) );
  XNOR U20821 ( .A(n15556), .B(x[1807]), .Z(n15557) );
  NAND U20822 ( .A(n15557), .B(y[1807]), .Z(n15558) );
  NAND U20823 ( .A(n15559), .B(n15558), .Z(n15560) );
  NAND U20824 ( .A(n15561), .B(n15560), .Z(n15562) );
  NANDN U20825 ( .A(n23542), .B(n15562), .Z(n15563) );
  NAND U20826 ( .A(n15564), .B(n15563), .Z(n15565) );
  NAND U20827 ( .A(n15565), .B(n23546), .Z(n15566) );
  NANDN U20828 ( .A(n15566), .B(x[1812]), .Z(n15570) );
  XNOR U20829 ( .A(n15566), .B(x[1812]), .Z(n15567) );
  NAND U20830 ( .A(n15568), .B(n15567), .Z(n15569) );
  NAND U20831 ( .A(n15570), .B(n15569), .Z(n15571) );
  NAND U20832 ( .A(n15572), .B(n15571), .Z(n15573) );
  NAND U20833 ( .A(n15574), .B(n15573), .Z(n15575) );
  NAND U20834 ( .A(n15576), .B(n15575), .Z(n15577) );
  NAND U20835 ( .A(n15578), .B(n15577), .Z(n15579) );
  NAND U20836 ( .A(n15580), .B(n15579), .Z(n15582) );
  NAND U20837 ( .A(n15582), .B(n15581), .Z(n15583) );
  OR U20838 ( .A(n23559), .B(n15583), .Z(n15584) );
  NANDN U20839 ( .A(n23560), .B(n15584), .Z(n15586) );
  XNOR U20840 ( .A(x[1818]), .B(n15586), .Z(n15585) );
  NANDN U20841 ( .A(y[1818]), .B(n15585), .Z(n15588) );
  NANDN U20842 ( .A(n15586), .B(x[1818]), .Z(n15587) );
  NAND U20843 ( .A(n15588), .B(n15587), .Z(n15590) );
  OR U20844 ( .A(n15590), .B(x[1819]), .Z(n15589) );
  AND U20845 ( .A(n23570), .B(n15589), .Z(n15593) );
  XOR U20846 ( .A(n15590), .B(x[1819]), .Z(n15591) );
  NAND U20847 ( .A(n15591), .B(y[1819]), .Z(n15592) );
  NAND U20848 ( .A(n15593), .B(n15592), .Z(n15594) );
  NAND U20849 ( .A(n15595), .B(n15594), .Z(n15596) );
  NAND U20850 ( .A(n15596), .B(n23574), .Z(n15597) );
  ANDN U20851 ( .B(n15597), .A(n23577), .Z(n15598) );
  OR U20852 ( .A(n23579), .B(n15598), .Z(n15600) );
  ANDN U20853 ( .B(x[1824]), .A(y[1824]), .Z(n23581) );
  NOR U20854 ( .A(n23587), .B(n23581), .Z(n15599) );
  NAND U20855 ( .A(n15600), .B(n15599), .Z(n15602) );
  NAND U20856 ( .A(n15602), .B(n15601), .Z(n15604) );
  NAND U20857 ( .A(n15604), .B(n15603), .Z(n15605) );
  AND U20858 ( .A(n15606), .B(n15605), .Z(n15608) );
  NANDN U20859 ( .A(n23598), .B(n23594), .Z(n15607) );
  OR U20860 ( .A(n15608), .B(n15607), .Z(n15609) );
  AND U20861 ( .A(n15610), .B(n15609), .Z(n15611) );
  NAND U20862 ( .A(n15611), .B(n23600), .Z(n15612) );
  NANDN U20863 ( .A(n23603), .B(n15612), .Z(n15613) );
  AND U20864 ( .A(n23604), .B(n15613), .Z(n15615) );
  NANDN U20865 ( .A(n15615), .B(n15614), .Z(n15616) );
  NANDN U20866 ( .A(n15617), .B(n15616), .Z(n15619) );
  NAND U20867 ( .A(n15619), .B(n15618), .Z(n15620) );
  AND U20868 ( .A(n23619), .B(n15620), .Z(n15621) );
  OR U20869 ( .A(n23622), .B(n15621), .Z(n15622) );
  AND U20870 ( .A(n23623), .B(n15622), .Z(n15623) );
  ANDN U20871 ( .B(n23625), .A(n15623), .Z(n15624) );
  NAND U20872 ( .A(n15624), .B(n23630), .Z(n15626) );
  ANDN U20873 ( .B(n15626), .A(n15625), .Z(n15627) );
  NAND U20874 ( .A(n15627), .B(n23627), .Z(n15628) );
  NAND U20875 ( .A(n15629), .B(n15628), .Z(n15631) );
  ANDN U20876 ( .B(n15631), .A(n15630), .Z(n15632) );
  NANDN U20877 ( .A(n15633), .B(n15632), .Z(n15634) );
  AND U20878 ( .A(n23637), .B(n15634), .Z(n15635) );
  NAND U20879 ( .A(n15635), .B(n23641), .Z(n15636) );
  NAND U20880 ( .A(n15637), .B(n15636), .Z(n15644) );
  NANDN U20881 ( .A(n15639), .B(n15638), .Z(n15640) );
  NANDN U20882 ( .A(n15641), .B(n15640), .Z(n15643) );
  ANDN U20883 ( .B(n15643), .A(n15642), .Z(n23645) );
  NAND U20884 ( .A(n15644), .B(n23645), .Z(n15645) );
  NAND U20885 ( .A(n15646), .B(n15645), .Z(n15647) );
  NANDN U20886 ( .A(n23650), .B(n15647), .Z(n15648) );
  NANDN U20887 ( .A(n15648), .B(y[1849]), .Z(n15652) );
  XNOR U20888 ( .A(n15648), .B(y[1849]), .Z(n15649) );
  NAND U20889 ( .A(n15650), .B(n15649), .Z(n15651) );
  NAND U20890 ( .A(n15652), .B(n15651), .Z(n15653) );
  NANDN U20891 ( .A(n15653), .B(n23655), .Z(n15654) );
  NAND U20892 ( .A(n15655), .B(n15654), .Z(n15656) );
  NANDN U20893 ( .A(n23660), .B(n15656), .Z(n15657) );
  NANDN U20894 ( .A(n23662), .B(n15657), .Z(n15658) );
  NAND U20895 ( .A(n15658), .B(n23663), .Z(n15659) );
  AND U20896 ( .A(n15660), .B(n15659), .Z(n15662) );
  OR U20897 ( .A(n15662), .B(y[1856]), .Z(n15661) );
  AND U20898 ( .A(n23670), .B(n15661), .Z(n15665) );
  XOR U20899 ( .A(y[1856]), .B(n15662), .Z(n15663) );
  NAND U20900 ( .A(x[1856]), .B(n15663), .Z(n15664) );
  NAND U20901 ( .A(n15665), .B(n15664), .Z(n15666) );
  NAND U20902 ( .A(n15667), .B(n15666), .Z(n15668) );
  NANDN U20903 ( .A(n23674), .B(n15668), .Z(n15669) );
  NANDN U20904 ( .A(n23676), .B(n15669), .Z(n15672) );
  NANDN U20905 ( .A(y[1860]), .B(x[1860]), .Z(n15670) );
  NANDN U20906 ( .A(n15671), .B(n15670), .Z(n23678) );
  ANDN U20907 ( .B(n15672), .A(n23678), .Z(n15675) );
  AND U20908 ( .A(n23679), .B(n15673), .Z(n15674) );
  NANDN U20909 ( .A(n15675), .B(n15674), .Z(n15676) );
  NANDN U20910 ( .A(n23681), .B(n15676), .Z(n15678) );
  ANDN U20911 ( .B(n15678), .A(n15677), .Z(n15679) );
  NAND U20912 ( .A(n15680), .B(n15679), .Z(n15681) );
  NANDN U20913 ( .A(n23685), .B(n15681), .Z(n15682) );
  NANDN U20914 ( .A(n23688), .B(n15682), .Z(n15683) );
  NAND U20915 ( .A(n15683), .B(n23690), .Z(n15684) );
  AND U20916 ( .A(n20269), .B(n15684), .Z(n15686) );
  NANDN U20917 ( .A(n15686), .B(n15685), .Z(n15689) );
  AND U20918 ( .A(n20268), .B(n15687), .Z(n15688) );
  NAND U20919 ( .A(n15689), .B(n15688), .Z(n15691) );
  NAND U20920 ( .A(n15691), .B(n15690), .Z(n15692) );
  NANDN U20921 ( .A(n15692), .B(n23697), .Z(n15695) );
  NANDN U20922 ( .A(n15693), .B(n20267), .Z(n15694) );
  AND U20923 ( .A(n15695), .B(n15694), .Z(n15696) );
  NANDN U20924 ( .A(n15697), .B(n15696), .Z(n15698) );
  NANDN U20925 ( .A(x[1873]), .B(n15698), .Z(n15701) );
  XNOR U20926 ( .A(x[1873]), .B(n15698), .Z(n15699) );
  NAND U20927 ( .A(n15699), .B(y[1873]), .Z(n15700) );
  NAND U20928 ( .A(n15701), .B(n15700), .Z(n15702) );
  AND U20929 ( .A(n15703), .B(n15702), .Z(n15704) );
  NANDN U20930 ( .A(n15704), .B(n23709), .Z(n15705) );
  NAND U20931 ( .A(n15706), .B(n15705), .Z(n15707) );
  NANDN U20932 ( .A(n15707), .B(y[1876]), .Z(n15711) );
  XNOR U20933 ( .A(n15707), .B(y[1876]), .Z(n15708) );
  NAND U20934 ( .A(n15709), .B(n15708), .Z(n15710) );
  NAND U20935 ( .A(n15711), .B(n15710), .Z(n15712) );
  NAND U20936 ( .A(n15713), .B(n15712), .Z(n15714) );
  NAND U20937 ( .A(n15715), .B(n15714), .Z(n15716) );
  NAND U20938 ( .A(n15717), .B(n15716), .Z(n15718) );
  NANDN U20939 ( .A(n23722), .B(n15718), .Z(n15721) );
  NANDN U20940 ( .A(y[1880]), .B(x[1880]), .Z(n15719) );
  NANDN U20941 ( .A(n15720), .B(n15719), .Z(n23724) );
  ANDN U20942 ( .B(n15721), .A(n23724), .Z(n15724) );
  NAND U20943 ( .A(n15722), .B(n23725), .Z(n15723) );
  OR U20944 ( .A(n15724), .B(n15723), .Z(n15725) );
  ANDN U20945 ( .B(n15725), .A(n23728), .Z(n15726) );
  OR U20946 ( .A(n15727), .B(n15726), .Z(n15728) );
  NAND U20947 ( .A(n15728), .B(n23731), .Z(n15729) );
  NAND U20948 ( .A(n15729), .B(n23734), .Z(n15730) );
  NAND U20949 ( .A(n15730), .B(n23735), .Z(n15731) );
  NANDN U20950 ( .A(n15732), .B(n15731), .Z(n15735) );
  NAND U20951 ( .A(n15736), .B(n15735), .Z(n15733) );
  AND U20952 ( .A(n15734), .B(n15733), .Z(n15739) );
  XOR U20953 ( .A(n15736), .B(n15735), .Z(n15737) );
  NAND U20954 ( .A(n15737), .B(y[1889]), .Z(n15738) );
  NAND U20955 ( .A(n15739), .B(n15738), .Z(n15740) );
  NANDN U20956 ( .A(n15741), .B(n15740), .Z(n15742) );
  NANDN U20957 ( .A(y[1891]), .B(n15742), .Z(n15745) );
  XNOR U20958 ( .A(y[1891]), .B(n15742), .Z(n15743) );
  NAND U20959 ( .A(n15743), .B(x[1891]), .Z(n15744) );
  NAND U20960 ( .A(n15745), .B(n15744), .Z(n15746) );
  AND U20961 ( .A(n23746), .B(n15746), .Z(n15749) );
  NANDN U20962 ( .A(n15747), .B(n23747), .Z(n15748) );
  OR U20963 ( .A(n15749), .B(n15748), .Z(n15752) );
  OR U20964 ( .A(n15751), .B(n15750), .Z(n23750) );
  ANDN U20965 ( .B(n15752), .A(n23750), .Z(n15753) );
  ANDN U20966 ( .B(n23751), .A(n15753), .Z(n15755) );
  NAND U20967 ( .A(n15755), .B(n15754), .Z(n15756) );
  AND U20968 ( .A(n23754), .B(n15756), .Z(n15757) );
  NAND U20969 ( .A(n15758), .B(n15757), .Z(n15759) );
  NAND U20970 ( .A(n15760), .B(n15759), .Z(n15762) );
  AND U20971 ( .A(n15762), .B(n15761), .Z(n15763) );
  NAND U20972 ( .A(n15764), .B(n15763), .Z(n15765) );
  NAND U20973 ( .A(n15766), .B(n15765), .Z(n15767) );
  NAND U20974 ( .A(n15768), .B(n15767), .Z(n15769) );
  NANDN U20975 ( .A(n23768), .B(n15769), .Z(n15772) );
  NAND U20976 ( .A(n15771), .B(n15770), .Z(n23769) );
  ANDN U20977 ( .B(n15772), .A(n23769), .Z(n15773) );
  OR U20978 ( .A(n23771), .B(n15773), .Z(n15775) );
  ANDN U20979 ( .B(n15775), .A(n15774), .Z(n15776) );
  AND U20980 ( .A(n23774), .B(n15776), .Z(n15777) );
  NANDN U20981 ( .A(n15777), .B(n23775), .Z(n15779) );
  ANDN U20982 ( .B(n15779), .A(n15778), .Z(n15780) );
  NANDN U20983 ( .A(n15780), .B(n23779), .Z(n15782) );
  ANDN U20984 ( .B(n15782), .A(n15781), .Z(n15784) );
  NANDN U20985 ( .A(n15784), .B(n15783), .Z(n15785) );
  AND U20986 ( .A(n23789), .B(n15785), .Z(n15786) );
  OR U20987 ( .A(n23792), .B(n15786), .Z(n15787) );
  NAND U20988 ( .A(n15787), .B(n23793), .Z(n15788) );
  NANDN U20989 ( .A(n23796), .B(n15788), .Z(n15789) );
  NANDN U20990 ( .A(n15790), .B(n15789), .Z(n15791) );
  NAND U20991 ( .A(n15791), .B(n23800), .Z(n15792) );
  AND U20992 ( .A(n23801), .B(n15792), .Z(n15793) );
  NANDN U20993 ( .A(n15794), .B(n15793), .Z(n15795) );
  NANDN U20994 ( .A(n23804), .B(n15795), .Z(n15796) );
  AND U20995 ( .A(n23805), .B(n15796), .Z(n15797) );
  OR U20996 ( .A(n15797), .B(n23808), .Z(n15798) );
  AND U20997 ( .A(n23811), .B(n15798), .Z(n15799) );
  OR U20998 ( .A(n15799), .B(n23814), .Z(n15800) );
  NANDN U20999 ( .A(n15801), .B(n15800), .Z(n15802) );
  AND U21000 ( .A(n23818), .B(n15802), .Z(n15803) );
  OR U21001 ( .A(n23820), .B(n15803), .Z(n15804) );
  ANDN U21002 ( .B(n15804), .A(n23822), .Z(n15805) );
  OR U21003 ( .A(n15806), .B(n15805), .Z(n15807) );
  NANDN U21004 ( .A(n15808), .B(n15807), .Z(n15809) );
  NAND U21005 ( .A(n15809), .B(n23829), .Z(n15810) );
  NAND U21006 ( .A(n15810), .B(n23833), .Z(n15811) );
  NAND U21007 ( .A(n15811), .B(n23835), .Z(n15812) );
  AND U21008 ( .A(n23838), .B(n15812), .Z(n15813) );
  NANDN U21009 ( .A(n15813), .B(n23839), .Z(n15814) );
  NANDN U21010 ( .A(n23841), .B(n15814), .Z(n15816) );
  NAND U21011 ( .A(n15816), .B(n15815), .Z(n15817) );
  ANDN U21012 ( .B(n15817), .A(n23846), .Z(n15822) );
  XOR U21013 ( .A(n15818), .B(y[1932]), .Z(n15820) );
  NAND U21014 ( .A(n15820), .B(n15819), .Z(n15821) );
  NANDN U21015 ( .A(n15822), .B(n15821), .Z(n15824) );
  NANDN U21016 ( .A(n15824), .B(n15823), .Z(n15826) );
  ANDN U21017 ( .B(n15826), .A(n15825), .Z(n15827) );
  ANDN U21018 ( .B(n15828), .A(n15827), .Z(n15832) );
  NANDN U21019 ( .A(n15832), .B(n15831), .Z(n15829) );
  AND U21020 ( .A(n15830), .B(n15829), .Z(n15835) );
  XNOR U21021 ( .A(n15832), .B(n15831), .Z(n15833) );
  NAND U21022 ( .A(n15833), .B(y[1934]), .Z(n15834) );
  NAND U21023 ( .A(n15835), .B(n15834), .Z(n15836) );
  NAND U21024 ( .A(n15836), .B(n23854), .Z(n15837) );
  NAND U21025 ( .A(n15837), .B(n23855), .Z(n15838) );
  AND U21026 ( .A(n23857), .B(n15838), .Z(n15839) );
  NANDN U21027 ( .A(n15839), .B(n23859), .Z(n15840) );
  AND U21028 ( .A(n23861), .B(n15840), .Z(n15841) );
  NANDN U21029 ( .A(n15841), .B(n23863), .Z(n15842) );
  AND U21030 ( .A(n23866), .B(n15842), .Z(n15843) );
  NANDN U21031 ( .A(n15843), .B(n23867), .Z(n15844) );
  NAND U21032 ( .A(n15844), .B(n23870), .Z(n15845) );
  NAND U21033 ( .A(n15845), .B(n23871), .Z(n15846) );
  NAND U21034 ( .A(n15846), .B(n23874), .Z(n15847) );
  AND U21035 ( .A(n23875), .B(n15847), .Z(n15848) );
  OR U21036 ( .A(n23878), .B(n15848), .Z(n15850) );
  NAND U21037 ( .A(n15850), .B(n15849), .Z(n15852) );
  NAND U21038 ( .A(n15852), .B(n15851), .Z(n15854) );
  NAND U21039 ( .A(n15854), .B(n15853), .Z(n15855) );
  NANDN U21040 ( .A(n15856), .B(n15855), .Z(n15857) );
  AND U21041 ( .A(n23891), .B(n15857), .Z(n15858) );
  NAND U21042 ( .A(n15859), .B(n15858), .Z(n15860) );
  NANDN U21043 ( .A(n23894), .B(n15860), .Z(n15861) );
  NAND U21044 ( .A(n15861), .B(n23895), .Z(n15862) );
  AND U21045 ( .A(n23897), .B(n15862), .Z(n15863) );
  NANDN U21046 ( .A(n15863), .B(n23899), .Z(n15864) );
  NANDN U21047 ( .A(n23904), .B(n15864), .Z(n15865) );
  AND U21048 ( .A(n15866), .B(n15865), .Z(n15868) );
  NANDN U21049 ( .A(n15868), .B(n15867), .Z(n15870) );
  ANDN U21050 ( .B(n15870), .A(n15869), .Z(n15871) );
  NANDN U21051 ( .A(n23908), .B(n15871), .Z(n15873) );
  NAND U21052 ( .A(n15873), .B(n15872), .Z(n15875) );
  ANDN U21053 ( .B(n15875), .A(n15874), .Z(n15879) );
  NANDN U21054 ( .A(n15877), .B(n15876), .Z(n15878) );
  AND U21055 ( .A(n15879), .B(n15878), .Z(n15880) );
  NANDN U21056 ( .A(n15880), .B(n23915), .Z(n15881) );
  ANDN U21057 ( .B(n15881), .A(n23918), .Z(n15882) );
  NANDN U21058 ( .A(n15882), .B(n23919), .Z(n15883) );
  NANDN U21059 ( .A(n23922), .B(n15883), .Z(n15884) );
  NAND U21060 ( .A(n15884), .B(n23923), .Z(n15885) );
  NANDN U21061 ( .A(n23925), .B(n15885), .Z(n15886) );
  AND U21062 ( .A(n23927), .B(n15886), .Z(n15887) );
  NANDN U21063 ( .A(n15887), .B(n23929), .Z(n15888) );
  NANDN U21064 ( .A(n23931), .B(n15888), .Z(n15891) );
  NANDN U21065 ( .A(x[1971]), .B(y[1971]), .Z(n15890) );
  NAND U21066 ( .A(n15890), .B(n15889), .Z(n23934) );
  ANDN U21067 ( .B(n15891), .A(n23934), .Z(n15893) );
  NANDN U21068 ( .A(n15893), .B(n15892), .Z(n15894) );
  NANDN U21069 ( .A(n15895), .B(n15894), .Z(n15897) );
  NAND U21070 ( .A(n15897), .B(n15896), .Z(n15898) );
  NAND U21071 ( .A(n15898), .B(n23948), .Z(n15899) );
  NANDN U21072 ( .A(n23950), .B(n15899), .Z(n15900) );
  AND U21073 ( .A(n23951), .B(n15900), .Z(n15901) );
  ANDN U21074 ( .B(n23954), .A(n15901), .Z(n15903) );
  NAND U21075 ( .A(n15903), .B(n15902), .Z(n15905) );
  ANDN U21076 ( .B(n15905), .A(n15904), .Z(n15906) );
  NAND U21077 ( .A(n15906), .B(n23955), .Z(n15908) );
  NANDN U21078 ( .A(y[1980]), .B(x[1980]), .Z(n15907) );
  AND U21079 ( .A(n15908), .B(n15907), .Z(n15909) );
  NAND U21080 ( .A(n15910), .B(n15909), .Z(n15911) );
  NAND U21081 ( .A(n15912), .B(n15911), .Z(n15913) );
  NAND U21082 ( .A(n15914), .B(n15913), .Z(n15916) );
  NAND U21083 ( .A(n15916), .B(n15915), .Z(n15917) );
  NANDN U21084 ( .A(n15917), .B(n23967), .Z(n15918) );
  NANDN U21085 ( .A(n23969), .B(n15918), .Z(n15919) );
  NAND U21086 ( .A(n15919), .B(n23971), .Z(n15920) );
  NAND U21087 ( .A(n15920), .B(n23973), .Z(n15921) );
  NAND U21088 ( .A(n15921), .B(n23976), .Z(n15922) );
  ANDN U21089 ( .B(n15922), .A(n23978), .Z(n15923) );
  NANDN U21090 ( .A(n15923), .B(n23980), .Z(n15924) );
  AND U21091 ( .A(n23982), .B(n15924), .Z(n15925) );
  NANDN U21092 ( .A(n15925), .B(n23985), .Z(n15926) );
  NANDN U21093 ( .A(n15927), .B(n15926), .Z(n15928) );
  NANDN U21094 ( .A(n23990), .B(n15928), .Z(n15929) );
  NAND U21095 ( .A(n15930), .B(n15929), .Z(n15931) );
  NAND U21096 ( .A(n15931), .B(n23993), .Z(n15932) );
  NAND U21097 ( .A(n15933), .B(n15932), .Z(n15934) );
  NAND U21098 ( .A(n15935), .B(n15934), .Z(n15936) );
  NAND U21099 ( .A(n15937), .B(n15936), .Z(n15938) );
  NAND U21100 ( .A(n15939), .B(n15938), .Z(n15940) );
  NAND U21101 ( .A(n15941), .B(n15940), .Z(n15943) );
  NAND U21102 ( .A(n15943), .B(n15942), .Z(n15944) );
  NANDN U21103 ( .A(n15944), .B(n24005), .Z(n15947) );
  NANDN U21104 ( .A(n15946), .B(n15945), .Z(n24008) );
  ANDN U21105 ( .B(n15947), .A(n24008), .Z(n15948) );
  OR U21106 ( .A(n24010), .B(n15948), .Z(n15951) );
  OR U21107 ( .A(n15950), .B(n15949), .Z(n24012) );
  ANDN U21108 ( .B(n15951), .A(n24012), .Z(n15956) );
  NANDN U21109 ( .A(n15953), .B(n15952), .Z(n15955) );
  ANDN U21110 ( .B(n15955), .A(n15954), .Z(n24013) );
  NANDN U21111 ( .A(n15956), .B(n24013), .Z(n15957) );
  AND U21112 ( .A(n15958), .B(n15957), .Z(n15959) );
  NANDN U21113 ( .A(n15959), .B(n15960), .Z(n15963) );
  XNOR U21114 ( .A(n15960), .B(n15959), .Z(n15961) );
  NAND U21115 ( .A(n15961), .B(x[2004]), .Z(n15962) );
  NAND U21116 ( .A(n15963), .B(n15962), .Z(n15964) );
  AND U21117 ( .A(n15965), .B(n15964), .Z(n15966) );
  NANDN U21118 ( .A(n15966), .B(n24020), .Z(n15967) );
  AND U21119 ( .A(n24021), .B(n15967), .Z(n15968) );
  NANDN U21120 ( .A(n15968), .B(n24023), .Z(n15969) );
  NAND U21121 ( .A(n15969), .B(n24025), .Z(n15970) );
  AND U21122 ( .A(n24027), .B(n15970), .Z(n15971) );
  NANDN U21123 ( .A(n15971), .B(n24029), .Z(n15973) );
  NAND U21124 ( .A(n15973), .B(n15972), .Z(n15975) );
  NAND U21125 ( .A(n15975), .B(n15974), .Z(n15976) );
  AND U21126 ( .A(n15977), .B(n15976), .Z(n15978) );
  NANDN U21127 ( .A(n15978), .B(n24043), .Z(n15979) );
  AND U21128 ( .A(n24046), .B(n15979), .Z(n15980) );
  NANDN U21129 ( .A(n15980), .B(n24050), .Z(n15982) );
  NAND U21130 ( .A(n15982), .B(n15981), .Z(n15983) );
  NANDN U21131 ( .A(n24054), .B(n15983), .Z(n15984) );
  NAND U21132 ( .A(n15985), .B(n15984), .Z(n15986) );
  NAND U21133 ( .A(n15986), .B(n24058), .Z(n15987) );
  NAND U21134 ( .A(n15988), .B(n15987), .Z(n15989) );
  NANDN U21135 ( .A(n24062), .B(n15989), .Z(n15990) );
  NAND U21136 ( .A(n15990), .B(n24063), .Z(n15991) );
  NANDN U21137 ( .A(n24066), .B(n15991), .Z(n15992) );
  NAND U21138 ( .A(n15992), .B(n24067), .Z(n15993) );
  NAND U21139 ( .A(n15993), .B(n24070), .Z(n15994) );
  NANDN U21140 ( .A(n24071), .B(n15994), .Z(n15996) );
  ANDN U21141 ( .B(n15996), .A(n15995), .Z(n15997) );
  NAND U21142 ( .A(n15997), .B(n24074), .Z(n15998) );
  AND U21143 ( .A(n15999), .B(n15998), .Z(n16000) );
  NAND U21144 ( .A(n16000), .B(n24075), .Z(n16001) );
  NANDN U21145 ( .A(n16002), .B(n16001), .Z(n16004) );
  NANDN U21146 ( .A(n16004), .B(x[2030]), .Z(n16007) );
  XOR U21147 ( .A(n16004), .B(n16003), .Z(n16005) );
  NANDN U21148 ( .A(y[2030]), .B(n16005), .Z(n16006) );
  AND U21149 ( .A(n16007), .B(n16006), .Z(n16008) );
  OR U21150 ( .A(n16008), .B(y[2031]), .Z(n16011) );
  XOR U21151 ( .A(y[2031]), .B(n16008), .Z(n16009) );
  NAND U21152 ( .A(n16009), .B(x[2031]), .Z(n16010) );
  NAND U21153 ( .A(n16011), .B(n16010), .Z(n16013) );
  ANDN U21154 ( .B(n16013), .A(n16012), .Z(n16014) );
  OR U21155 ( .A(n16015), .B(n16014), .Z(n16018) );
  ANDN U21156 ( .B(n24089), .A(n16016), .Z(n16017) );
  NAND U21157 ( .A(n16018), .B(n16017), .Z(n16019) );
  NANDN U21158 ( .A(n24092), .B(n16019), .Z(n16020) );
  NAND U21159 ( .A(n16021), .B(n16020), .Z(n16022) );
  NAND U21160 ( .A(n16022), .B(n24095), .Z(n16023) );
  NAND U21161 ( .A(n16024), .B(n16023), .Z(n16025) );
  NAND U21162 ( .A(n16026), .B(n16025), .Z(n16027) );
  NAND U21163 ( .A(n16028), .B(n16027), .Z(n16029) );
  NAND U21164 ( .A(n16030), .B(n16029), .Z(n16031) );
  NAND U21165 ( .A(n16032), .B(n16031), .Z(n16034) );
  NAND U21166 ( .A(n16034), .B(n16033), .Z(n16041) );
  OR U21167 ( .A(n16036), .B(n16035), .Z(n16037) );
  NANDN U21168 ( .A(n16038), .B(n16037), .Z(n16040) );
  ANDN U21169 ( .B(n16040), .A(n16039), .Z(n24107) );
  NANDN U21170 ( .A(n16041), .B(n24107), .Z(n16042) );
  NAND U21171 ( .A(n16042), .B(n24109), .Z(n16043) );
  NANDN U21172 ( .A(n16044), .B(n16043), .Z(n16048) );
  NANDN U21173 ( .A(n16046), .B(n16045), .Z(n16047) );
  NANDN U21174 ( .A(n16048), .B(n16047), .Z(n16049) );
  NAND U21175 ( .A(n16049), .B(n24113), .Z(n16050) );
  AND U21176 ( .A(n24115), .B(n16050), .Z(n16051) );
  NANDN U21177 ( .A(n16051), .B(n24117), .Z(n16052) );
  NANDN U21178 ( .A(n24120), .B(n16052), .Z(n16053) );
  NAND U21179 ( .A(n16053), .B(n24121), .Z(n16054) );
  NANDN U21180 ( .A(n24123), .B(n16054), .Z(n16055) );
  NAND U21181 ( .A(n16055), .B(n24125), .Z(n16056) );
  AND U21182 ( .A(n24128), .B(n16056), .Z(n16057) );
  NANDN U21183 ( .A(n16057), .B(n24129), .Z(n16060) );
  NANDN U21184 ( .A(y[2055]), .B(x[2055]), .Z(n16058) );
  NANDN U21185 ( .A(n16059), .B(n16058), .Z(n24132) );
  ANDN U21186 ( .B(n16060), .A(n24132), .Z(n16064) );
  NAND U21187 ( .A(n16061), .B(y[2055]), .Z(n16063) );
  AND U21188 ( .A(n16063), .B(n16062), .Z(n24133) );
  NANDN U21189 ( .A(n16064), .B(n24133), .Z(n16067) );
  ANDN U21190 ( .B(n16066), .A(n16065), .Z(n24138) );
  ANDN U21191 ( .B(n16067), .A(n24138), .Z(n16069) );
  NAND U21192 ( .A(n16069), .B(n16068), .Z(n16070) );
  NANDN U21193 ( .A(n16070), .B(y[2058]), .Z(n16073) );
  XNOR U21194 ( .A(n16070), .B(y[2058]), .Z(n16071) );
  NANDN U21195 ( .A(x[2058]), .B(n16071), .Z(n16072) );
  NAND U21196 ( .A(n16073), .B(n16072), .Z(n16074) );
  NAND U21197 ( .A(n16075), .B(n16074), .Z(n16076) );
  NAND U21198 ( .A(n16077), .B(n16076), .Z(n16078) );
  NAND U21199 ( .A(n16079), .B(n16078), .Z(n16080) );
  NANDN U21200 ( .A(n24148), .B(n16080), .Z(n16081) );
  NAND U21201 ( .A(n16082), .B(n16081), .Z(n16083) );
  NAND U21202 ( .A(n16083), .B(n24151), .Z(n16084) );
  NAND U21203 ( .A(n16085), .B(n16084), .Z(n16087) );
  NAND U21204 ( .A(n16087), .B(n16086), .Z(n16088) );
  NANDN U21205 ( .A(n16088), .B(n16089), .Z(n16092) );
  XNOR U21206 ( .A(n16089), .B(n16088), .Z(n16090) );
  NAND U21207 ( .A(n16090), .B(x[2065]), .Z(n16091) );
  NAND U21208 ( .A(n16092), .B(n16091), .Z(n16093) );
  AND U21209 ( .A(n24159), .B(n16093), .Z(n16098) );
  NANDN U21210 ( .A(n24162), .B(n16094), .Z(n16095) );
  NANDN U21211 ( .A(n16096), .B(n16095), .Z(n16097) );
  NANDN U21212 ( .A(n16098), .B(n16097), .Z(n16099) );
  NAND U21213 ( .A(n16099), .B(n24163), .Z(n16100) );
  NANDN U21214 ( .A(n24166), .B(n16100), .Z(n16101) );
  ANDN U21215 ( .B(n16101), .A(n24168), .Z(n16102) );
  ANDN U21216 ( .B(n24169), .A(n16102), .Z(n16104) );
  NAND U21217 ( .A(n16104), .B(n16103), .Z(n16105) );
  AND U21218 ( .A(n24172), .B(n16105), .Z(n16107) );
  OR U21219 ( .A(n16107), .B(n16106), .Z(n16108) );
  ANDN U21220 ( .B(n16108), .A(n24176), .Z(n16109) );
  NANDN U21221 ( .A(n16109), .B(n24179), .Z(n16110) );
  ANDN U21222 ( .B(n16110), .A(n24181), .Z(n16112) );
  NANDN U21223 ( .A(n16112), .B(n16111), .Z(n16113) );
  NAND U21224 ( .A(n16113), .B(n24185), .Z(n16114) );
  NAND U21225 ( .A(n16114), .B(n24187), .Z(n16116) );
  ANDN U21226 ( .B(n16116), .A(n16115), .Z(n16117) );
  NAND U21227 ( .A(n16118), .B(n16117), .Z(n16119) );
  NAND U21228 ( .A(n16120), .B(n16119), .Z(n16121) );
  AND U21229 ( .A(n24193), .B(n16121), .Z(n16126) );
  NAND U21230 ( .A(n16122), .B(n24195), .Z(n16123) );
  AND U21231 ( .A(n16124), .B(n16123), .Z(n16125) );
  OR U21232 ( .A(n16126), .B(n16125), .Z(n16127) );
  NAND U21233 ( .A(n16127), .B(n24198), .Z(n16128) );
  NANDN U21234 ( .A(n24200), .B(n16128), .Z(n16129) );
  NANDN U21235 ( .A(n24202), .B(n16129), .Z(n16130) );
  AND U21236 ( .A(n24203), .B(n16130), .Z(n16131) );
  NANDN U21237 ( .A(n16132), .B(n16131), .Z(n16133) );
  AND U21238 ( .A(n24205), .B(n16133), .Z(n16135) );
  NAND U21239 ( .A(n16135), .B(n16134), .Z(n16136) );
  AND U21240 ( .A(n16137), .B(n16136), .Z(n16138) );
  NAND U21241 ( .A(n16139), .B(n16138), .Z(n16140) );
  AND U21242 ( .A(n16141), .B(n16140), .Z(n16142) );
  ANDN U21243 ( .B(n16143), .A(n16142), .Z(n16144) );
  NAND U21244 ( .A(n16144), .B(n24215), .Z(n16149) );
  NANDN U21245 ( .A(n16146), .B(n16145), .Z(n16147) );
  NANDN U21246 ( .A(n16148), .B(n16147), .Z(n24218) );
  ANDN U21247 ( .B(n16149), .A(n24218), .Z(n16151) );
  NANDN U21248 ( .A(n16151), .B(n16150), .Z(n16152) );
  ANDN U21249 ( .B(n16152), .A(n24222), .Z(n16153) );
  ANDN U21250 ( .B(n16154), .A(n16153), .Z(n16155) );
  NANDN U21251 ( .A(n16155), .B(n24225), .Z(n16156) );
  NANDN U21252 ( .A(n16157), .B(n16156), .Z(n16158) );
  NANDN U21253 ( .A(n20260), .B(n16158), .Z(n16159) );
  NAND U21254 ( .A(n16160), .B(n16159), .Z(n16161) );
  NAND U21255 ( .A(n16161), .B(n20259), .Z(n16162) );
  NAND U21256 ( .A(n16163), .B(n16162), .Z(n16164) );
  NAND U21257 ( .A(n16165), .B(n16164), .Z(n16166) );
  NAND U21258 ( .A(n16167), .B(n16166), .Z(n16168) );
  NAND U21259 ( .A(n16169), .B(n16168), .Z(n16170) );
  NAND U21260 ( .A(n16171), .B(n16170), .Z(n16172) );
  AND U21261 ( .A(n24241), .B(n16172), .Z(n16176) );
  NANDN U21262 ( .A(n16174), .B(n16173), .Z(n16175) );
  NAND U21263 ( .A(n16176), .B(n16175), .Z(n16177) );
  ANDN U21264 ( .B(n16177), .A(n24243), .Z(n16178) );
  NANDN U21265 ( .A(n16178), .B(n24245), .Z(n16179) );
  NANDN U21266 ( .A(n24248), .B(n16179), .Z(n16180) );
  NAND U21267 ( .A(n16180), .B(n24249), .Z(n16181) );
  NANDN U21268 ( .A(n16182), .B(n16181), .Z(n16184) );
  XNOR U21269 ( .A(y[2108]), .B(n16184), .Z(n16183) );
  NANDN U21270 ( .A(x[2108]), .B(n16183), .Z(n16186) );
  NANDN U21271 ( .A(n16184), .B(y[2108]), .Z(n16185) );
  AND U21272 ( .A(n16186), .B(n16185), .Z(n16187) );
  NANDN U21273 ( .A(n16187), .B(n24255), .Z(n16190) );
  AND U21274 ( .A(n24257), .B(n16188), .Z(n16189) );
  NAND U21275 ( .A(n16190), .B(n16189), .Z(n16191) );
  NANDN U21276 ( .A(n24260), .B(n16191), .Z(n16192) );
  NAND U21277 ( .A(n16192), .B(n24261), .Z(n16193) );
  AND U21278 ( .A(n24264), .B(n16193), .Z(n16195) );
  NAND U21279 ( .A(n16195), .B(n16194), .Z(n16197) );
  ANDN U21280 ( .B(n16197), .A(n16196), .Z(n16198) );
  NAND U21281 ( .A(n16198), .B(n24265), .Z(n16201) );
  NAND U21282 ( .A(n16199), .B(n24271), .Z(n16200) );
  ANDN U21283 ( .B(n16201), .A(n16200), .Z(n16207) );
  NANDN U21284 ( .A(n16203), .B(n16202), .Z(n16205) );
  ANDN U21285 ( .B(n16205), .A(n16204), .Z(n16206) );
  NANDN U21286 ( .A(n16207), .B(n16206), .Z(n16209) );
  ANDN U21287 ( .B(n16209), .A(n16208), .Z(n16210) );
  NANDN U21288 ( .A(n16210), .B(n24282), .Z(n16211) );
  AND U21289 ( .A(n24285), .B(n16211), .Z(n16212) );
  OR U21290 ( .A(n16212), .B(n24287), .Z(n16213) );
  NANDN U21291 ( .A(n16214), .B(n16213), .Z(n16215) );
  NANDN U21292 ( .A(n16215), .B(y[2122]), .Z(n16219) );
  XNOR U21293 ( .A(n16215), .B(y[2122]), .Z(n16216) );
  NAND U21294 ( .A(n16217), .B(n16216), .Z(n16218) );
  NAND U21295 ( .A(n16219), .B(n16218), .Z(n16220) );
  NAND U21296 ( .A(n16220), .B(n24292), .Z(n16221) );
  AND U21297 ( .A(n16222), .B(n16221), .Z(n16223) );
  NAND U21298 ( .A(n16223), .B(n24294), .Z(n16230) );
  NAND U21299 ( .A(n16225), .B(n16224), .Z(n16226) );
  NANDN U21300 ( .A(n16227), .B(n16226), .Z(n16229) );
  ANDN U21301 ( .B(n16229), .A(n16228), .Z(n24296) );
  NAND U21302 ( .A(n16230), .B(n24296), .Z(n16233) );
  ANDN U21303 ( .B(n24298), .A(n16231), .Z(n16232) );
  NAND U21304 ( .A(n16233), .B(n16232), .Z(n16235) );
  ANDN U21305 ( .B(n16235), .A(n16234), .Z(n16236) );
  OR U21306 ( .A(n16236), .B(y[2129]), .Z(n16239) );
  XOR U21307 ( .A(y[2129]), .B(n16236), .Z(n16237) );
  NAND U21308 ( .A(n16237), .B(x[2129]), .Z(n16238) );
  NAND U21309 ( .A(n16239), .B(n16238), .Z(n16240) );
  AND U21310 ( .A(n24306), .B(n16240), .Z(n16241) );
  OR U21311 ( .A(n16242), .B(n16241), .Z(n16245) );
  NOR U21312 ( .A(n16244), .B(n16243), .Z(n24310) );
  NAND U21313 ( .A(n16245), .B(n24310), .Z(n16246) );
  NANDN U21314 ( .A(n24312), .B(n16246), .Z(n16247) );
  NAND U21315 ( .A(n16248), .B(n16247), .Z(n16250) );
  ANDN U21316 ( .B(n16250), .A(n16249), .Z(n16251) );
  NANDN U21317 ( .A(n16251), .B(n16252), .Z(n16255) );
  XNOR U21318 ( .A(n16252), .B(n16251), .Z(n16253) );
  NAND U21319 ( .A(n16253), .B(x[2135]), .Z(n16254) );
  NAND U21320 ( .A(n16255), .B(n16254), .Z(n16256) );
  AND U21321 ( .A(n16257), .B(n16256), .Z(n16258) );
  ANDN U21322 ( .B(n24325), .A(n16258), .Z(n16260) );
  NAND U21323 ( .A(n16260), .B(n16259), .Z(n16261) );
  AND U21324 ( .A(n16262), .B(n16261), .Z(n16263) );
  NAND U21325 ( .A(n16263), .B(n24326), .Z(n16264) );
  NANDN U21326 ( .A(n24329), .B(n16264), .Z(n16265) );
  AND U21327 ( .A(n24330), .B(n16265), .Z(n16267) );
  NOR U21328 ( .A(n16267), .B(n16266), .Z(n16268) );
  NAND U21329 ( .A(n16268), .B(n24333), .Z(n16269) );
  NAND U21330 ( .A(n16269), .B(n24334), .Z(n16271) );
  ANDN U21331 ( .B(n16271), .A(n16270), .Z(n16272) );
  NANDN U21332 ( .A(n16272), .B(n24338), .Z(n16273) );
  NAND U21333 ( .A(n16273), .B(n24341), .Z(n16274) );
  NAND U21334 ( .A(n16274), .B(n24342), .Z(n16275) );
  AND U21335 ( .A(n24344), .B(n16275), .Z(n16276) );
  NANDN U21336 ( .A(n16276), .B(n24346), .Z(n16277) );
  NAND U21337 ( .A(n16277), .B(n24348), .Z(n16278) );
  NANDN U21338 ( .A(n24351), .B(n16278), .Z(n16279) );
  NAND U21339 ( .A(n16279), .B(n24352), .Z(n16281) );
  AND U21340 ( .A(n16281), .B(n16280), .Z(n16282) );
  NAND U21341 ( .A(n16282), .B(n24355), .Z(n16286) );
  NANDN U21342 ( .A(n16284), .B(n16283), .Z(n16285) );
  AND U21343 ( .A(n16286), .B(n16285), .Z(n16287) );
  NAND U21344 ( .A(n16288), .B(n16287), .Z(n16289) );
  NAND U21345 ( .A(n16290), .B(n16289), .Z(n16291) );
  NAND U21346 ( .A(n16292), .B(n16291), .Z(n16294) );
  NAND U21347 ( .A(n16294), .B(n16293), .Z(n16295) );
  NANDN U21348 ( .A(n16295), .B(n24368), .Z(n16297) );
  ANDN U21349 ( .B(n16297), .A(n16296), .Z(n16298) );
  NANDN U21350 ( .A(n16298), .B(n24372), .Z(n16300) );
  ANDN U21351 ( .B(n16300), .A(n16299), .Z(n16301) );
  NAND U21352 ( .A(n16301), .B(n24374), .Z(n16302) );
  NAND U21353 ( .A(n16302), .B(n24377), .Z(n16304) );
  ANDN U21354 ( .B(n16304), .A(n16303), .Z(n16305) );
  OR U21355 ( .A(n16305), .B(n24381), .Z(n16307) );
  ANDN U21356 ( .B(n16307), .A(n16306), .Z(n16308) );
  NAND U21357 ( .A(n16309), .B(n16308), .Z(n16310) );
  NAND U21358 ( .A(n16311), .B(n16310), .Z(n16312) );
  AND U21359 ( .A(n24386), .B(n16312), .Z(n16315) );
  ANDN U21360 ( .B(n24388), .A(n16313), .Z(n16314) );
  NANDN U21361 ( .A(n16315), .B(n16314), .Z(n16316) );
  NANDN U21362 ( .A(n24390), .B(n16316), .Z(n16320) );
  NAND U21363 ( .A(n16317), .B(y[2167]), .Z(n16318) );
  NANDN U21364 ( .A(n16319), .B(n16318), .Z(n24393) );
  ANDN U21365 ( .B(n16320), .A(n24393), .Z(n16321) );
  ANDN U21366 ( .B(n24394), .A(n16321), .Z(n16323) );
  NAND U21367 ( .A(n16323), .B(n16322), .Z(n16324) );
  AND U21368 ( .A(n24397), .B(n16324), .Z(n16325) );
  NAND U21369 ( .A(n16326), .B(n16325), .Z(n16327) );
  NAND U21370 ( .A(n16328), .B(n16327), .Z(n16330) );
  NAND U21371 ( .A(n16330), .B(n16329), .Z(n16332) );
  XNOR U21372 ( .A(x[2172]), .B(n16332), .Z(n16331) );
  NANDN U21373 ( .A(y[2172]), .B(n16331), .Z(n16334) );
  NANDN U21374 ( .A(n16332), .B(x[2172]), .Z(n16333) );
  NAND U21375 ( .A(n16334), .B(n16333), .Z(n16336) );
  NANDN U21376 ( .A(n16336), .B(y[2173]), .Z(n16339) );
  XOR U21377 ( .A(n16336), .B(n16335), .Z(n16337) );
  NANDN U21378 ( .A(x[2173]), .B(n16337), .Z(n16338) );
  AND U21379 ( .A(n16339), .B(n16338), .Z(n16340) );
  OR U21380 ( .A(n16340), .B(x[2174]), .Z(n16343) );
  XOR U21381 ( .A(x[2174]), .B(n16340), .Z(n16341) );
  NAND U21382 ( .A(n16341), .B(y[2174]), .Z(n16342) );
  NAND U21383 ( .A(n16343), .B(n16342), .Z(n16344) );
  NAND U21384 ( .A(n16345), .B(n16344), .Z(n16346) );
  NANDN U21385 ( .A(n16347), .B(n16346), .Z(n16349) );
  NANDN U21386 ( .A(n16349), .B(x[2176]), .Z(n16352) );
  XOR U21387 ( .A(n16349), .B(n16348), .Z(n16350) );
  NANDN U21388 ( .A(y[2176]), .B(n16350), .Z(n16351) );
  AND U21389 ( .A(n16352), .B(n16351), .Z(n16353) );
  OR U21390 ( .A(n16353), .B(y[2177]), .Z(n16356) );
  XOR U21391 ( .A(y[2177]), .B(n16353), .Z(n16354) );
  NAND U21392 ( .A(n16354), .B(x[2177]), .Z(n16355) );
  NAND U21393 ( .A(n16356), .B(n16355), .Z(n16358) );
  ANDN U21394 ( .B(n16358), .A(n16357), .Z(n16359) );
  ANDN U21395 ( .B(n24418), .A(n16359), .Z(n16361) );
  NAND U21396 ( .A(n16361), .B(n16360), .Z(n16362) );
  ANDN U21397 ( .B(n16362), .A(n24420), .Z(n16364) );
  ANDN U21398 ( .B(n16364), .A(n16363), .Z(n16365) );
  OR U21399 ( .A(n24422), .B(n16365), .Z(n16366) );
  NANDN U21400 ( .A(n24425), .B(n16366), .Z(n16367) );
  NANDN U21401 ( .A(n24426), .B(n16367), .Z(n16368) );
  AND U21402 ( .A(n24428), .B(n16368), .Z(n16369) );
  OR U21403 ( .A(n16370), .B(n16369), .Z(n16371) );
  NANDN U21404 ( .A(n16372), .B(n16371), .Z(n16373) );
  ANDN U21405 ( .B(n16373), .A(n24437), .Z(n16374) );
  NANDN U21406 ( .A(n16374), .B(n24438), .Z(n16375) );
  AND U21407 ( .A(n16376), .B(n16375), .Z(n16377) );
  NAND U21408 ( .A(n16377), .B(n24441), .Z(n16378) );
  NAND U21409 ( .A(n16379), .B(n16378), .Z(n16380) );
  AND U21410 ( .A(n16381), .B(n16380), .Z(n16383) );
  NANDN U21411 ( .A(y[2190]), .B(x[2190]), .Z(n16382) );
  NAND U21412 ( .A(n16383), .B(n16382), .Z(n16387) );
  OR U21413 ( .A(n16385), .B(n16384), .Z(n16386) );
  ANDN U21414 ( .B(n16387), .A(n16386), .Z(n16388) );
  ANDN U21415 ( .B(n24452), .A(n16388), .Z(n16390) );
  NAND U21416 ( .A(n16390), .B(n16389), .Z(n16391) );
  AND U21417 ( .A(n24454), .B(n16391), .Z(n16393) );
  ANDN U21418 ( .B(n16393), .A(n16392), .Z(n16394) );
  OR U21419 ( .A(n24457), .B(n16394), .Z(n16395) );
  NANDN U21420 ( .A(n24459), .B(n16395), .Z(n16396) );
  NAND U21421 ( .A(n16396), .B(n24460), .Z(n16397) );
  ANDN U21422 ( .B(n16397), .A(n24462), .Z(n16398) );
  OR U21423 ( .A(n24465), .B(n16398), .Z(n16399) );
  NANDN U21424 ( .A(n24466), .B(n16399), .Z(n16400) );
  NAND U21425 ( .A(n16400), .B(n24469), .Z(n16401) );
  NAND U21426 ( .A(n16401), .B(n24473), .Z(n16402) );
  NANDN U21427 ( .A(n16403), .B(n16402), .Z(n16404) );
  ANDN U21428 ( .B(n16404), .A(n24476), .Z(n16405) );
  OR U21429 ( .A(n16406), .B(n16405), .Z(n16407) );
  NANDN U21430 ( .A(n24480), .B(n16407), .Z(n16408) );
  NANDN U21431 ( .A(n16409), .B(n16408), .Z(n16413) );
  NAND U21432 ( .A(n16411), .B(n16410), .Z(n16412) );
  NANDN U21433 ( .A(n16413), .B(n16412), .Z(n16414) );
  ANDN U21434 ( .B(n16414), .A(n24485), .Z(n16415) );
  NANDN U21435 ( .A(n16415), .B(n24486), .Z(n16416) );
  NANDN U21436 ( .A(n24488), .B(n16416), .Z(n16417) );
  NANDN U21437 ( .A(n24490), .B(n16417), .Z(n16418) );
  NANDN U21438 ( .A(n24493), .B(n16418), .Z(n16419) );
  NANDN U21439 ( .A(n24495), .B(n16419), .Z(n16420) );
  ANDN U21440 ( .B(n16420), .A(n24496), .Z(n16421) );
  NANDN U21441 ( .A(n16421), .B(n24498), .Z(n16422) );
  ANDN U21442 ( .B(n16422), .A(n24500), .Z(n16423) );
  NANDN U21443 ( .A(n16423), .B(n24502), .Z(n16425) );
  ANDN U21444 ( .B(n16425), .A(n16424), .Z(n16426) );
  OR U21445 ( .A(n16427), .B(n16426), .Z(n16428) );
  ANDN U21446 ( .B(n16428), .A(n24510), .Z(n16430) );
  NANDN U21447 ( .A(n16430), .B(n16429), .Z(n16431) );
  AND U21448 ( .A(n24514), .B(n16431), .Z(n16436) );
  NANDN U21449 ( .A(n16433), .B(n16432), .Z(n16434) );
  AND U21450 ( .A(n24516), .B(n16434), .Z(n16435) );
  NANDN U21451 ( .A(n16436), .B(n16435), .Z(n16437) );
  NAND U21452 ( .A(n16437), .B(n24518), .Z(n16438) );
  ANDN U21453 ( .B(n16438), .A(n24521), .Z(n16439) );
  NANDN U21454 ( .A(n16439), .B(n24522), .Z(n16440) );
  AND U21455 ( .A(n24526), .B(n16440), .Z(n16441) );
  NANDN U21456 ( .A(n16441), .B(n24528), .Z(n16443) );
  ANDN U21457 ( .B(n16443), .A(n16442), .Z(n16445) );
  OR U21458 ( .A(n16445), .B(n16444), .Z(n16447) );
  ANDN U21459 ( .B(n16447), .A(n16446), .Z(n16448) );
  NANDN U21460 ( .A(n16448), .B(n24540), .Z(n16450) );
  ANDN U21461 ( .B(n16450), .A(n16449), .Z(n16451) );
  NAND U21462 ( .A(n16451), .B(n24542), .Z(n16452) );
  NAND U21463 ( .A(n16452), .B(n24544), .Z(n16454) );
  ANDN U21464 ( .B(n16454), .A(n16453), .Z(n16455) );
  OR U21465 ( .A(n16455), .B(n24549), .Z(n16457) );
  ANDN U21466 ( .B(n16457), .A(n16456), .Z(n16458) );
  NAND U21467 ( .A(n16459), .B(n16458), .Z(n16460) );
  NAND U21468 ( .A(n16461), .B(n16460), .Z(n16462) );
  NAND U21469 ( .A(n16462), .B(n24554), .Z(n16463) );
  NAND U21470 ( .A(n16464), .B(n16463), .Z(n16465) );
  NANDN U21471 ( .A(n16466), .B(n16465), .Z(n16467) );
  AND U21472 ( .A(n20251), .B(n16467), .Z(n16469) );
  NAND U21473 ( .A(n16469), .B(n16468), .Z(n16470) );
  AND U21474 ( .A(n16471), .B(n16470), .Z(n16472) );
  NAND U21475 ( .A(n16473), .B(n16472), .Z(n16474) );
  AND U21476 ( .A(n16475), .B(n16474), .Z(n16476) );
  OR U21477 ( .A(n16477), .B(n16476), .Z(n16480) );
  NOR U21478 ( .A(n16479), .B(n16478), .Z(n24576) );
  NAND U21479 ( .A(n16480), .B(n24576), .Z(n16482) );
  NAND U21480 ( .A(n16482), .B(n16481), .Z(n16483) );
  NANDN U21481 ( .A(n16483), .B(n24579), .Z(n16484) );
  NAND U21482 ( .A(n16485), .B(n16484), .Z(n16486) );
  NANDN U21483 ( .A(n16487), .B(n16486), .Z(n16489) );
  XNOR U21484 ( .A(y[2247]), .B(n16489), .Z(n16488) );
  NANDN U21485 ( .A(x[2247]), .B(n16488), .Z(n16491) );
  NANDN U21486 ( .A(n16489), .B(y[2247]), .Z(n16490) );
  NAND U21487 ( .A(n16491), .B(n16490), .Z(n16493) );
  NANDN U21488 ( .A(n16493), .B(x[2248]), .Z(n16496) );
  XOR U21489 ( .A(n16493), .B(n16492), .Z(n16494) );
  NANDN U21490 ( .A(y[2248]), .B(n16494), .Z(n16495) );
  NAND U21491 ( .A(n16496), .B(n16495), .Z(n16497) );
  NANDN U21492 ( .A(n16497), .B(n24591), .Z(n16498) );
  AND U21493 ( .A(n16499), .B(n16498), .Z(n16508) );
  NANDN U21494 ( .A(y[2252]), .B(x[2252]), .Z(n16505) );
  NANDN U21495 ( .A(n16501), .B(n16500), .Z(n16502) );
  NANDN U21496 ( .A(n16503), .B(n16502), .Z(n16504) );
  NAND U21497 ( .A(n16505), .B(n16504), .Z(n24595) );
  NANDN U21498 ( .A(n24595), .B(n16506), .Z(n16507) );
  OR U21499 ( .A(n16508), .B(n16507), .Z(n16509) );
  AND U21500 ( .A(n24596), .B(n16509), .Z(n16510) );
  NAND U21501 ( .A(n16511), .B(n16510), .Z(n16512) );
  NAND U21502 ( .A(n16513), .B(n16512), .Z(n16515) );
  ANDN U21503 ( .B(n16515), .A(n16514), .Z(n16516) );
  OR U21504 ( .A(n16516), .B(n24603), .Z(n16517) );
  NAND U21505 ( .A(n16517), .B(n24604), .Z(n16518) );
  ANDN U21506 ( .B(n16518), .A(n24606), .Z(n16519) );
  NANDN U21507 ( .A(n16519), .B(n24608), .Z(n16521) );
  ANDN U21508 ( .B(n16521), .A(n16520), .Z(n16522) );
  NAND U21509 ( .A(n16523), .B(n16522), .Z(n16524) );
  NAND U21510 ( .A(n16525), .B(n16524), .Z(n16526) );
  NAND U21511 ( .A(n16526), .B(n24614), .Z(n16527) );
  NAND U21512 ( .A(n16527), .B(n24616), .Z(n16528) );
  AND U21513 ( .A(n24618), .B(n16528), .Z(n16529) );
  NANDN U21514 ( .A(n16529), .B(n24621), .Z(n16534) );
  AND U21515 ( .A(n16531), .B(n16530), .Z(n20250) );
  NOR U21516 ( .A(n20250), .B(n16532), .Z(n16533) );
  NAND U21517 ( .A(n16534), .B(n16533), .Z(n16535) );
  NAND U21518 ( .A(n16535), .B(n24624), .Z(n16536) );
  AND U21519 ( .A(n16537), .B(n16536), .Z(n16538) );
  OR U21520 ( .A(n24628), .B(n16538), .Z(n16542) );
  NANDN U21521 ( .A(y[2270]), .B(x[2270]), .Z(n16539) );
  AND U21522 ( .A(n16540), .B(n16539), .Z(n16541) );
  NAND U21523 ( .A(n16542), .B(n16541), .Z(n16544) );
  NAND U21524 ( .A(n16544), .B(n16543), .Z(n16545) );
  NANDN U21525 ( .A(x[2271]), .B(n16545), .Z(n16548) );
  XNOR U21526 ( .A(x[2271]), .B(n16545), .Z(n16546) );
  NAND U21527 ( .A(n16546), .B(y[2271]), .Z(n16547) );
  NAND U21528 ( .A(n16548), .B(n16547), .Z(n16550) );
  ANDN U21529 ( .B(n16550), .A(n16549), .Z(n16551) );
  OR U21530 ( .A(n24636), .B(n16551), .Z(n16552) );
  AND U21531 ( .A(n24638), .B(n16552), .Z(n16553) );
  OR U21532 ( .A(n24641), .B(n16553), .Z(n16554) );
  NAND U21533 ( .A(n16554), .B(n24642), .Z(n16555) );
  NANDN U21534 ( .A(n24645), .B(n16555), .Z(n16556) );
  AND U21535 ( .A(n24646), .B(n16556), .Z(n16557) );
  NANDN U21536 ( .A(n16557), .B(n24649), .Z(n16560) );
  NOR U21537 ( .A(n16559), .B(n16558), .Z(n24650) );
  NAND U21538 ( .A(n16560), .B(n24650), .Z(n16561) );
  NANDN U21539 ( .A(n24652), .B(n16561), .Z(n16562) );
  NAND U21540 ( .A(n16562), .B(n24654), .Z(n16564) );
  ANDN U21541 ( .B(n16564), .A(n16563), .Z(n16565) );
  NANDN U21542 ( .A(n16565), .B(n24660), .Z(n16566) );
  ANDN U21543 ( .B(n16566), .A(n24663), .Z(n16568) );
  NAND U21544 ( .A(n16568), .B(n16567), .Z(n16570) );
  ANDN U21545 ( .B(n16570), .A(n16569), .Z(n16571) );
  NANDN U21546 ( .A(n16571), .B(n24667), .Z(n16572) );
  NAND U21547 ( .A(n16572), .B(n24668), .Z(n16573) );
  NAND U21548 ( .A(n16573), .B(n24670), .Z(n16574) );
  NAND U21549 ( .A(n16574), .B(n24672), .Z(n16575) );
  NAND U21550 ( .A(n16575), .B(n24675), .Z(n16576) );
  AND U21551 ( .A(n24676), .B(n16576), .Z(n16577) );
  OR U21552 ( .A(n24679), .B(n16577), .Z(n16580) );
  NANDN U21553 ( .A(y[2292]), .B(x[2292]), .Z(n16579) );
  ANDN U21554 ( .B(n16579), .A(n16578), .Z(n24680) );
  NAND U21555 ( .A(n16580), .B(n24680), .Z(n16581) );
  NANDN U21556 ( .A(n24682), .B(n16581), .Z(n16582) );
  NAND U21557 ( .A(n16583), .B(n16582), .Z(n16585) );
  NAND U21558 ( .A(n16585), .B(n16584), .Z(n16586) );
  NANDN U21559 ( .A(n16586), .B(n24686), .Z(n16587) );
  AND U21560 ( .A(n16588), .B(n16587), .Z(n16590) );
  NAND U21561 ( .A(n16590), .B(n16589), .Z(n16591) );
  AND U21562 ( .A(n16592), .B(n16591), .Z(n16593) );
  OR U21563 ( .A(n16594), .B(n16593), .Z(n16597) );
  NOR U21564 ( .A(n16596), .B(n16595), .Z(n24698) );
  NAND U21565 ( .A(n16597), .B(n24698), .Z(n16599) );
  NAND U21566 ( .A(n16599), .B(n16598), .Z(n16600) );
  NANDN U21567 ( .A(n16600), .B(n24701), .Z(n16603) );
  ANDN U21568 ( .B(n24702), .A(n16601), .Z(n16602) );
  NAND U21569 ( .A(n16603), .B(n16602), .Z(n16604) );
  NANDN U21570 ( .A(n16605), .B(n16604), .Z(n16606) );
  NAND U21571 ( .A(n16607), .B(n16606), .Z(n16608) );
  NAND U21572 ( .A(n16608), .B(n24713), .Z(n16610) );
  NANDN U21573 ( .A(n16610), .B(n16609), .Z(n16614) );
  NOR U21574 ( .A(n16612), .B(n16611), .Z(n16613) );
  NAND U21575 ( .A(n16614), .B(n16613), .Z(n16615) );
  NAND U21576 ( .A(n16616), .B(n16615), .Z(n16617) );
  NAND U21577 ( .A(n16618), .B(n16617), .Z(n16619) );
  NAND U21578 ( .A(n16619), .B(n24719), .Z(n16620) );
  NAND U21579 ( .A(n16621), .B(n16620), .Z(n16622) );
  AND U21580 ( .A(n16623), .B(n16622), .Z(n16625) );
  OR U21581 ( .A(n16625), .B(y[2310]), .Z(n16624) );
  AND U21582 ( .A(n24729), .B(n16624), .Z(n16628) );
  XOR U21583 ( .A(n16625), .B(y[2310]), .Z(n16626) );
  NAND U21584 ( .A(n16626), .B(x[2310]), .Z(n16627) );
  NAND U21585 ( .A(n16628), .B(n16627), .Z(n16629) );
  AND U21586 ( .A(n16630), .B(n16629), .Z(n16631) );
  NANDN U21587 ( .A(n16631), .B(n24733), .Z(n16632) );
  NANDN U21588 ( .A(n24735), .B(n16632), .Z(n16633) );
  NANDN U21589 ( .A(n16634), .B(n16633), .Z(n16635) );
  NANDN U21590 ( .A(n24738), .B(n16635), .Z(n16637) );
  XNOR U21591 ( .A(x[2316]), .B(n16637), .Z(n16636) );
  NANDN U21592 ( .A(y[2316]), .B(n16636), .Z(n16639) );
  NANDN U21593 ( .A(n16637), .B(x[2316]), .Z(n16638) );
  AND U21594 ( .A(n16639), .B(n16638), .Z(n16640) );
  NAND U21595 ( .A(n16641), .B(n16640), .Z(n16642) );
  NAND U21596 ( .A(n16643), .B(n16642), .Z(n16644) );
  NAND U21597 ( .A(n16645), .B(n16644), .Z(n16647) );
  NAND U21598 ( .A(n16647), .B(n16646), .Z(n16648) );
  NANDN U21599 ( .A(n16648), .B(n24750), .Z(n16651) );
  OR U21600 ( .A(n16650), .B(n16649), .Z(n24752) );
  ANDN U21601 ( .B(n16651), .A(n24752), .Z(n16652) );
  OR U21602 ( .A(n24755), .B(n16652), .Z(n16655) );
  AND U21603 ( .A(n24756), .B(n16653), .Z(n16654) );
  NAND U21604 ( .A(n16655), .B(n16654), .Z(n16656) );
  NANDN U21605 ( .A(n24758), .B(n16656), .Z(n16657) );
  AND U21606 ( .A(n16658), .B(n16657), .Z(n16659) );
  OR U21607 ( .A(n16659), .B(n24763), .Z(n16660) );
  NANDN U21608 ( .A(n16661), .B(n16660), .Z(n16663) );
  ANDN U21609 ( .B(n16663), .A(n16662), .Z(n16664) );
  NANDN U21610 ( .A(n16664), .B(n24773), .Z(n16665) );
  AND U21611 ( .A(n24775), .B(n16665), .Z(n16666) );
  OR U21612 ( .A(n24777), .B(n16666), .Z(n16667) );
  NAND U21613 ( .A(n16667), .B(n24779), .Z(n16668) );
  NAND U21614 ( .A(n16668), .B(n24782), .Z(n16669) );
  NAND U21615 ( .A(n16669), .B(n24783), .Z(n16670) );
  NANDN U21616 ( .A(n24786), .B(n16670), .Z(n16672) );
  ANDN U21617 ( .B(n16672), .A(n16671), .Z(n16673) );
  NAND U21618 ( .A(n16673), .B(n24787), .Z(n16674) );
  AND U21619 ( .A(n16675), .B(n16674), .Z(n16676) );
  NAND U21620 ( .A(n16676), .B(n24790), .Z(n16677) );
  NAND U21621 ( .A(n16678), .B(n16677), .Z(n16679) );
  NAND U21622 ( .A(n16679), .B(n24798), .Z(n16681) );
  NANDN U21623 ( .A(n16681), .B(n16680), .Z(n16684) );
  ANDN U21624 ( .B(n16683), .A(n16682), .Z(n24799) );
  NAND U21625 ( .A(n16684), .B(n24799), .Z(n16685) );
  NANDN U21626 ( .A(n24802), .B(n16685), .Z(n16686) );
  NAND U21627 ( .A(n16687), .B(n16686), .Z(n16689) );
  NAND U21628 ( .A(n16689), .B(n16688), .Z(n16690) );
  NANDN U21629 ( .A(n16690), .B(n24806), .Z(n16691) );
  AND U21630 ( .A(n16692), .B(n16691), .Z(n16693) );
  ANDN U21631 ( .B(n24813), .A(n16693), .Z(n16695) );
  NAND U21632 ( .A(n16695), .B(n16694), .Z(n16697) );
  ANDN U21633 ( .B(n16697), .A(n16696), .Z(n16698) );
  AND U21634 ( .A(n24815), .B(n16698), .Z(n16705) );
  NANDN U21635 ( .A(n16700), .B(n16699), .Z(n16701) );
  NANDN U21636 ( .A(n16702), .B(n16701), .Z(n16704) );
  ANDN U21637 ( .B(n16704), .A(n16703), .Z(n24818) );
  NANDN U21638 ( .A(n16705), .B(n24818), .Z(n16708) );
  ANDN U21639 ( .B(n24819), .A(n16706), .Z(n16707) );
  NAND U21640 ( .A(n16708), .B(n16707), .Z(n16709) );
  NANDN U21641 ( .A(n24822), .B(n16709), .Z(n16710) );
  AND U21642 ( .A(n16711), .B(n16710), .Z(n16712) );
  NANDN U21643 ( .A(n16712), .B(n24826), .Z(n16713) );
  NAND U21644 ( .A(n16713), .B(n24827), .Z(n16714) );
  NAND U21645 ( .A(n16714), .B(n24829), .Z(n16715) );
  AND U21646 ( .A(n24831), .B(n16715), .Z(n16717) );
  NOR U21647 ( .A(n16717), .B(n16716), .Z(n16718) );
  NAND U21648 ( .A(n16719), .B(n16718), .Z(n16720) );
  NAND U21649 ( .A(n16721), .B(n16720), .Z(n16723) );
  ANDN U21650 ( .B(n16723), .A(n16722), .Z(n16725) );
  NANDN U21651 ( .A(n16725), .B(n16724), .Z(n16727) );
  ANDN U21652 ( .B(n16727), .A(n16726), .Z(n16730) );
  NAND U21653 ( .A(n16728), .B(n24840), .Z(n16729) );
  OR U21654 ( .A(n16730), .B(n16729), .Z(n16731) );
  AND U21655 ( .A(n16732), .B(n16731), .Z(n16733) );
  NAND U21656 ( .A(n16734), .B(n16733), .Z(n16735) );
  NAND U21657 ( .A(n16736), .B(n16735), .Z(n16737) );
  NAND U21658 ( .A(n16738), .B(n16737), .Z(n16740) );
  NAND U21659 ( .A(n16740), .B(n16739), .Z(n16741) );
  NANDN U21660 ( .A(n16741), .B(n24853), .Z(n16742) );
  AND U21661 ( .A(n16743), .B(n16742), .Z(n16744) );
  OR U21662 ( .A(n24857), .B(n16744), .Z(n16747) );
  NOR U21663 ( .A(n24859), .B(n16745), .Z(n16746) );
  NAND U21664 ( .A(n16747), .B(n16746), .Z(n16748) );
  NAND U21665 ( .A(n16748), .B(n24861), .Z(n16750) );
  ANDN U21666 ( .B(n16750), .A(n16749), .Z(n16751) );
  NANDN U21667 ( .A(n16751), .B(n24865), .Z(n16752) );
  NANDN U21668 ( .A(n16753), .B(n16752), .Z(n16755) );
  NAND U21669 ( .A(n16755), .B(n16754), .Z(n16756) );
  AND U21670 ( .A(n16757), .B(n16756), .Z(n16758) );
  OR U21671 ( .A(n16759), .B(n16758), .Z(n16760) );
  NANDN U21672 ( .A(n24878), .B(n16760), .Z(n16762) );
  NAND U21673 ( .A(n16762), .B(n16761), .Z(n16763) );
  NANDN U21674 ( .A(n24875), .B(n16763), .Z(n16765) );
  XNOR U21675 ( .A(y[2379]), .B(n16765), .Z(n16764) );
  NANDN U21676 ( .A(x[2379]), .B(n16764), .Z(n16767) );
  NANDN U21677 ( .A(n16765), .B(y[2379]), .Z(n16766) );
  NAND U21678 ( .A(n16767), .B(n16766), .Z(n16768) );
  NANDN U21679 ( .A(n16768), .B(x[2380]), .Z(n16772) );
  XNOR U21680 ( .A(n16768), .B(x[2380]), .Z(n16769) );
  NAND U21681 ( .A(n16770), .B(n16769), .Z(n16771) );
  AND U21682 ( .A(n16772), .B(n16771), .Z(n16773) );
  OR U21683 ( .A(n16773), .B(y[2381]), .Z(n16776) );
  XOR U21684 ( .A(y[2381]), .B(n16773), .Z(n16774) );
  NAND U21685 ( .A(n16774), .B(x[2381]), .Z(n16775) );
  NAND U21686 ( .A(n16776), .B(n16775), .Z(n16778) );
  ANDN U21687 ( .B(n16778), .A(n16777), .Z(n16782) );
  OR U21688 ( .A(n16780), .B(n16779), .Z(n16781) );
  OR U21689 ( .A(n16782), .B(n16781), .Z(n16783) );
  NANDN U21690 ( .A(n16784), .B(n16783), .Z(n16786) );
  NANDN U21691 ( .A(n16786), .B(x[2384]), .Z(n16789) );
  XOR U21692 ( .A(n16786), .B(n16785), .Z(n16787) );
  NANDN U21693 ( .A(y[2384]), .B(n16787), .Z(n16788) );
  AND U21694 ( .A(n16789), .B(n16788), .Z(n16790) );
  OR U21695 ( .A(n16790), .B(y[2385]), .Z(n16793) );
  XOR U21696 ( .A(y[2385]), .B(n16790), .Z(n16791) );
  NAND U21697 ( .A(n16791), .B(x[2385]), .Z(n16792) );
  NAND U21698 ( .A(n16793), .B(n16792), .Z(n16794) );
  NANDN U21699 ( .A(n16795), .B(n16794), .Z(n16796) );
  NANDN U21700 ( .A(n16797), .B(n16796), .Z(n16799) );
  NANDN U21701 ( .A(n16799), .B(y[2387]), .Z(n16802) );
  XOR U21702 ( .A(n16799), .B(n16798), .Z(n16800) );
  NANDN U21703 ( .A(x[2387]), .B(n16800), .Z(n16801) );
  AND U21704 ( .A(n16802), .B(n16801), .Z(n16803) );
  NANDN U21705 ( .A(n16803), .B(n16804), .Z(n16807) );
  XNOR U21706 ( .A(n16804), .B(n16803), .Z(n16805) );
  NAND U21707 ( .A(n16805), .B(y[2388]), .Z(n16806) );
  NAND U21708 ( .A(n16807), .B(n16806), .Z(n16808) );
  AND U21709 ( .A(n24901), .B(n16808), .Z(n16809) );
  OR U21710 ( .A(n16810), .B(n16809), .Z(n16811) );
  NANDN U21711 ( .A(n24905), .B(n16811), .Z(n16812) );
  NANDN U21712 ( .A(n24907), .B(n16812), .Z(n16815) );
  NANDN U21713 ( .A(y[2392]), .B(x[2392]), .Z(n16813) );
  NANDN U21714 ( .A(n16814), .B(n16813), .Z(n24909) );
  ANDN U21715 ( .B(n16815), .A(n24909), .Z(n16817) );
  NANDN U21716 ( .A(n16817), .B(n16816), .Z(n16818) );
  NAND U21717 ( .A(n16818), .B(n24914), .Z(n16819) );
  ANDN U21718 ( .B(n16819), .A(n24917), .Z(n16820) );
  NANDN U21719 ( .A(n16820), .B(n24921), .Z(n16823) );
  NOR U21720 ( .A(n16822), .B(n16821), .Z(n24923) );
  NAND U21721 ( .A(n16823), .B(n24923), .Z(n16824) );
  NANDN U21722 ( .A(n16825), .B(n16824), .Z(n16826) );
  AND U21723 ( .A(n16826), .B(n24927), .Z(n16827) );
  NANDN U21724 ( .A(n16828), .B(n16827), .Z(n16829) );
  AND U21725 ( .A(n16830), .B(n16829), .Z(n16831) );
  NAND U21726 ( .A(n16832), .B(n16831), .Z(n16833) );
  NAND U21727 ( .A(n16834), .B(n16833), .Z(n16835) );
  NAND U21728 ( .A(n16836), .B(n16835), .Z(n16838) );
  NAND U21729 ( .A(n16838), .B(n16837), .Z(n16839) );
  NANDN U21730 ( .A(n16839), .B(n24939), .Z(n16842) );
  OR U21731 ( .A(n16841), .B(n16840), .Z(n24942) );
  ANDN U21732 ( .B(n16842), .A(n24942), .Z(n16843) );
  NANDN U21733 ( .A(n16843), .B(n24943), .Z(n16844) );
  AND U21734 ( .A(n24946), .B(n16844), .Z(n16845) );
  NANDN U21735 ( .A(n16845), .B(n24947), .Z(n16846) );
  NANDN U21736 ( .A(n24950), .B(n16846), .Z(n16847) );
  NAND U21737 ( .A(n16847), .B(n24951), .Z(n16848) );
  AND U21738 ( .A(n24955), .B(n16848), .Z(n16849) );
  NANDN U21739 ( .A(n16849), .B(n24957), .Z(n16851) );
  NAND U21740 ( .A(n16851), .B(n16850), .Z(n16854) );
  OR U21741 ( .A(n16853), .B(n16852), .Z(n24961) );
  ANDN U21742 ( .B(n16854), .A(n24961), .Z(n16855) );
  OR U21743 ( .A(n16856), .B(n16855), .Z(n16857) );
  NAND U21744 ( .A(n16858), .B(n16857), .Z(n16859) );
  NAND U21745 ( .A(n16860), .B(n16859), .Z(n16865) );
  NANDN U21746 ( .A(n16862), .B(n16861), .Z(n16863) );
  AND U21747 ( .A(n24973), .B(n16863), .Z(n16864) );
  NAND U21748 ( .A(n16865), .B(n16864), .Z(n16866) );
  AND U21749 ( .A(n24976), .B(n16866), .Z(n16867) );
  NANDN U21750 ( .A(n16867), .B(n24977), .Z(n16871) );
  NAND U21751 ( .A(n16868), .B(x[2419]), .Z(n16869) );
  NANDN U21752 ( .A(n16870), .B(n16869), .Z(n24979) );
  ANDN U21753 ( .B(n16871), .A(n24979), .Z(n16872) );
  OR U21754 ( .A(n24982), .B(n16872), .Z(n16873) );
  NANDN U21755 ( .A(n24984), .B(n16873), .Z(n16874) );
  NAND U21756 ( .A(n16874), .B(n24985), .Z(n16875) );
  ANDN U21757 ( .B(n16875), .A(n24987), .Z(n16876) );
  NANDN U21758 ( .A(n16876), .B(n24989), .Z(n16878) );
  NAND U21759 ( .A(n16878), .B(n16877), .Z(n16880) );
  ANDN U21760 ( .B(n16880), .A(n16879), .Z(n16881) );
  NANDN U21761 ( .A(n16881), .B(n24997), .Z(n16882) );
  NANDN U21762 ( .A(n16883), .B(n16882), .Z(n16885) );
  ANDN U21763 ( .B(n16885), .A(n16884), .Z(n16886) );
  OR U21764 ( .A(n16886), .B(y[2429]), .Z(n16889) );
  XOR U21765 ( .A(y[2429]), .B(n16886), .Z(n16887) );
  NAND U21766 ( .A(n16887), .B(x[2429]), .Z(n16888) );
  NAND U21767 ( .A(n16889), .B(n16888), .Z(n16890) );
  AND U21768 ( .A(n25008), .B(n16890), .Z(n16896) );
  NANDN U21769 ( .A(n16892), .B(n16891), .Z(n16894) );
  ANDN U21770 ( .B(n16894), .A(n16893), .Z(n16895) );
  NANDN U21771 ( .A(n16896), .B(n16895), .Z(n16897) );
  NAND U21772 ( .A(n16897), .B(n25011), .Z(n16898) );
  NAND U21773 ( .A(n16898), .B(n25015), .Z(n16901) );
  OR U21774 ( .A(n16900), .B(n16899), .Z(n25017) );
  ANDN U21775 ( .B(n16901), .A(n25017), .Z(n16902) );
  NANDN U21776 ( .A(n16902), .B(n25019), .Z(n16903) );
  NANDN U21777 ( .A(n25021), .B(n16903), .Z(n16904) );
  AND U21778 ( .A(n25023), .B(n16904), .Z(n16906) );
  NANDN U21779 ( .A(n16906), .B(n16905), .Z(n16907) );
  NANDN U21780 ( .A(n16908), .B(n16907), .Z(n16909) );
  NANDN U21781 ( .A(n25032), .B(n16909), .Z(n16910) );
  NAND U21782 ( .A(n16911), .B(n16910), .Z(n16912) );
  NAND U21783 ( .A(n16912), .B(n25036), .Z(n16913) );
  NANDN U21784 ( .A(n16914), .B(n16913), .Z(n16915) );
  NANDN U21785 ( .A(n25040), .B(n16915), .Z(n16917) );
  NAND U21786 ( .A(n16917), .B(n16916), .Z(n16919) );
  NANDN U21787 ( .A(y[2444]), .B(n16919), .Z(n16918) );
  AND U21788 ( .A(n25045), .B(n16918), .Z(n16922) );
  XNOR U21789 ( .A(y[2444]), .B(n16919), .Z(n16920) );
  NAND U21790 ( .A(n16920), .B(x[2444]), .Z(n16921) );
  NAND U21791 ( .A(n16922), .B(n16921), .Z(n16923) );
  NAND U21792 ( .A(n16924), .B(n16923), .Z(n16925) );
  NANDN U21793 ( .A(n25049), .B(n16925), .Z(n16927) );
  NAND U21794 ( .A(n16927), .B(n16926), .Z(n16928) );
  NANDN U21795 ( .A(n25052), .B(n16928), .Z(n16930) );
  XNOR U21796 ( .A(y[2449]), .B(n16930), .Z(n16929) );
  NANDN U21797 ( .A(x[2449]), .B(n16929), .Z(n16932) );
  NANDN U21798 ( .A(n16930), .B(y[2449]), .Z(n16931) );
  AND U21799 ( .A(n16932), .B(n16931), .Z(n16933) );
  NAND U21800 ( .A(n16934), .B(n16933), .Z(n16935) );
  NAND U21801 ( .A(n16936), .B(n16935), .Z(n16938) );
  ANDN U21802 ( .B(n16938), .A(n16937), .Z(n16939) );
  NAND U21803 ( .A(n16939), .B(n25061), .Z(n16940) );
  NAND U21804 ( .A(n16940), .B(n25064), .Z(n16942) );
  NANDN U21805 ( .A(n16942), .B(n16941), .Z(n16945) );
  NOR U21806 ( .A(n16944), .B(n16943), .Z(n25065) );
  NAND U21807 ( .A(n16945), .B(n25065), .Z(n16946) );
  NANDN U21808 ( .A(n16947), .B(n16946), .Z(n16948) );
  NAND U21809 ( .A(n16948), .B(n25069), .Z(n16950) );
  XNOR U21810 ( .A(x[2456]), .B(n16950), .Z(n16949) );
  NANDN U21811 ( .A(y[2456]), .B(n16949), .Z(n16952) );
  NANDN U21812 ( .A(n16950), .B(x[2456]), .Z(n16951) );
  AND U21813 ( .A(n16952), .B(n16951), .Z(n16953) );
  NAND U21814 ( .A(n16954), .B(n16953), .Z(n16955) );
  NAND U21815 ( .A(n16956), .B(n16955), .Z(n16957) );
  NAND U21816 ( .A(n16958), .B(n16957), .Z(n16959) );
  NANDN U21817 ( .A(n25082), .B(n16959), .Z(n16963) );
  NAND U21818 ( .A(n16960), .B(x[2460]), .Z(n16962) );
  NAND U21819 ( .A(n16962), .B(n16961), .Z(n25083) );
  ANDN U21820 ( .B(n16963), .A(n25083), .Z(n16964) );
  NANDN U21821 ( .A(n16964), .B(n25085), .Z(n16967) );
  ANDN U21822 ( .B(n25087), .A(n16965), .Z(n16966) );
  NAND U21823 ( .A(n16967), .B(n16966), .Z(n16969) );
  NAND U21824 ( .A(n16969), .B(n16968), .Z(n16970) );
  NANDN U21825 ( .A(n16970), .B(n25089), .Z(n16971) );
  AND U21826 ( .A(n16972), .B(n16971), .Z(n16977) );
  NANDN U21827 ( .A(n16974), .B(n16973), .Z(n16975) );
  AND U21828 ( .A(n25097), .B(n16975), .Z(n16976) );
  NANDN U21829 ( .A(n16977), .B(n16976), .Z(n16978) );
  NAND U21830 ( .A(n16978), .B(n25099), .Z(n16979) );
  NAND U21831 ( .A(n16979), .B(n25101), .Z(n16980) );
  AND U21832 ( .A(n25104), .B(n16980), .Z(n16981) );
  NANDN U21833 ( .A(n16981), .B(n25105), .Z(n16982) );
  NAND U21834 ( .A(n16982), .B(n25107), .Z(n16983) );
  NAND U21835 ( .A(n16983), .B(n25109), .Z(n16984) );
  AND U21836 ( .A(n25112), .B(n16984), .Z(n16985) );
  NANDN U21837 ( .A(n16985), .B(n25113), .Z(n16986) );
  NANDN U21838 ( .A(n25116), .B(n16986), .Z(n16988) );
  NAND U21839 ( .A(n16988), .B(n16987), .Z(n16989) );
  NANDN U21840 ( .A(n16989), .B(n25117), .Z(n16992) );
  ANDN U21841 ( .B(n25120), .A(n16990), .Z(n16991) );
  NAND U21842 ( .A(n16992), .B(n16991), .Z(n16993) );
  NANDN U21843 ( .A(n16994), .B(n16993), .Z(n16995) );
  NAND U21844 ( .A(n16996), .B(n16995), .Z(n16997) );
  NAND U21845 ( .A(n16997), .B(n25129), .Z(n16999) );
  NANDN U21846 ( .A(n16999), .B(n16998), .Z(n17001) );
  ANDN U21847 ( .B(n17001), .A(n17000), .Z(n17002) );
  NAND U21848 ( .A(n17002), .B(n25131), .Z(n17003) );
  AND U21849 ( .A(n25133), .B(n17003), .Z(n17004) );
  ANDN U21850 ( .B(n25136), .A(n17004), .Z(n17006) );
  NAND U21851 ( .A(n17006), .B(n17005), .Z(n17007) );
  NAND U21852 ( .A(n17007), .B(n25137), .Z(n17009) );
  OR U21853 ( .A(n17009), .B(y[2484]), .Z(n17008) );
  AND U21854 ( .A(n25143), .B(n17008), .Z(n17012) );
  XOR U21855 ( .A(n17009), .B(y[2484]), .Z(n17010) );
  NAND U21856 ( .A(n17010), .B(x[2484]), .Z(n17011) );
  NAND U21857 ( .A(n17012), .B(n17011), .Z(n17013) );
  NAND U21858 ( .A(n17014), .B(n17013), .Z(n17015) );
  NAND U21859 ( .A(n17015), .B(n25148), .Z(n17016) );
  AND U21860 ( .A(n25149), .B(n17016), .Z(n17017) );
  OR U21861 ( .A(n25151), .B(n17017), .Z(n17018) );
  AND U21862 ( .A(n25153), .B(n17018), .Z(n17019) );
  NANDN U21863 ( .A(n17019), .B(n25155), .Z(n17020) );
  NAND U21864 ( .A(n17020), .B(n25157), .Z(n17021) );
  NAND U21865 ( .A(n17021), .B(n25161), .Z(n17022) );
  NANDN U21866 ( .A(n25164), .B(n17022), .Z(n17024) );
  ANDN U21867 ( .B(n17024), .A(n17023), .Z(n17025) );
  NANDN U21868 ( .A(n17025), .B(n25168), .Z(n17027) );
  ANDN U21869 ( .B(n17027), .A(n17026), .Z(n17029) );
  NANDN U21870 ( .A(n17029), .B(n17028), .Z(n17031) );
  ANDN U21871 ( .B(n17031), .A(n17030), .Z(n17033) );
  NANDN U21872 ( .A(y[2498]), .B(x[2498]), .Z(n17032) );
  NAND U21873 ( .A(n17033), .B(n17032), .Z(n17034) );
  AND U21874 ( .A(n17035), .B(n17034), .Z(n17036) );
  NAND U21875 ( .A(n17036), .B(n25175), .Z(n17037) );
  NAND U21876 ( .A(n17038), .B(n17037), .Z(n17039) );
  NANDN U21877 ( .A(n25180), .B(n17039), .Z(n17042) );
  NANDN U21878 ( .A(y[2502]), .B(x[2502]), .Z(n17041) );
  NAND U21879 ( .A(n17041), .B(n17040), .Z(n25181) );
  ANDN U21880 ( .B(n17042), .A(n25181), .Z(n17043) );
  OR U21881 ( .A(n25183), .B(n17043), .Z(n17046) );
  ANDN U21882 ( .B(n25185), .A(n17044), .Z(n17045) );
  NAND U21883 ( .A(n17046), .B(n17045), .Z(n17048) );
  NAND U21884 ( .A(n17048), .B(n17047), .Z(n17049) );
  NANDN U21885 ( .A(n17049), .B(n25188), .Z(n17050) );
  AND U21886 ( .A(n17051), .B(n17050), .Z(n17052) );
  OR U21887 ( .A(n17053), .B(n17052), .Z(n17054) );
  NAND U21888 ( .A(n17055), .B(n17054), .Z(n17056) );
  NAND U21889 ( .A(n17057), .B(n17056), .Z(n17058) );
  NANDN U21890 ( .A(n17059), .B(n17058), .Z(n17061) );
  ANDN U21891 ( .B(n17061), .A(n17060), .Z(n17062) );
  OR U21892 ( .A(n17062), .B(n25202), .Z(n17064) );
  ANDN U21893 ( .B(n17064), .A(n17063), .Z(n17065) );
  NAND U21894 ( .A(n17065), .B(n25203), .Z(n17067) );
  ANDN U21895 ( .B(n17067), .A(n17066), .Z(n17068) );
  OR U21896 ( .A(n17069), .B(n17068), .Z(n17070) );
  NAND U21897 ( .A(n17071), .B(n17070), .Z(n17073) );
  NAND U21898 ( .A(n17073), .B(n17072), .Z(n17075) );
  NANDN U21899 ( .A(n17075), .B(n17074), .Z(n17076) );
  NAND U21900 ( .A(n17077), .B(n17076), .Z(n17078) );
  NAND U21901 ( .A(n17079), .B(n17078), .Z(n17084) );
  NANDN U21902 ( .A(n17081), .B(n17080), .Z(n17082) );
  AND U21903 ( .A(n25223), .B(n17082), .Z(n17083) );
  NAND U21904 ( .A(n17084), .B(n17083), .Z(n17085) );
  NAND U21905 ( .A(n17085), .B(n25225), .Z(n17086) );
  NAND U21906 ( .A(n17086), .B(n25227), .Z(n17087) );
  NANDN U21907 ( .A(n25230), .B(n17087), .Z(n17089) );
  ANDN U21908 ( .B(n17089), .A(n17088), .Z(n17090) );
  NAND U21909 ( .A(n17090), .B(n25231), .Z(n17093) );
  NANDN U21910 ( .A(n17091), .B(n25234), .Z(n17092) );
  ANDN U21911 ( .B(n17093), .A(n17092), .Z(n17094) );
  OR U21912 ( .A(n17095), .B(n17094), .Z(n17096) );
  NAND U21913 ( .A(n17097), .B(n17096), .Z(n17098) );
  NAND U21914 ( .A(n17099), .B(n17098), .Z(n17101) );
  NAND U21915 ( .A(n17101), .B(n17100), .Z(n17102) );
  NANDN U21916 ( .A(n17102), .B(n25246), .Z(n17103) );
  AND U21917 ( .A(n25247), .B(n17103), .Z(n17104) );
  OR U21918 ( .A(n25249), .B(n17104), .Z(n17107) );
  ANDN U21919 ( .B(n25251), .A(n17105), .Z(n17106) );
  NAND U21920 ( .A(n17107), .B(n17106), .Z(n17109) );
  NAND U21921 ( .A(n17109), .B(n17108), .Z(n17110) );
  NANDN U21922 ( .A(n17110), .B(n25254), .Z(n17111) );
  AND U21923 ( .A(n17112), .B(n17111), .Z(n17117) );
  NAND U21924 ( .A(n17114), .B(n17113), .Z(n17115) );
  ANDN U21925 ( .B(n17115), .A(n25261), .Z(n17116) );
  NANDN U21926 ( .A(n17117), .B(n17116), .Z(n17118) );
  NAND U21927 ( .A(n17118), .B(n25263), .Z(n17119) );
  ANDN U21928 ( .B(n17119), .A(n25265), .Z(n17120) );
  NANDN U21929 ( .A(n17120), .B(n25267), .Z(n17121) );
  ANDN U21930 ( .B(n17121), .A(n25269), .Z(n17122) );
  NANDN U21931 ( .A(n17122), .B(n25271), .Z(n17123) );
  ANDN U21932 ( .B(n17123), .A(n25274), .Z(n17124) );
  NANDN U21933 ( .A(n17124), .B(n25275), .Z(n17125) );
  NANDN U21934 ( .A(n25278), .B(n17125), .Z(n17132) );
  NANDN U21935 ( .A(n17127), .B(n17126), .Z(n17128) );
  NANDN U21936 ( .A(n17129), .B(n17128), .Z(n17131) );
  ANDN U21937 ( .B(n17131), .A(n17130), .Z(n25279) );
  NAND U21938 ( .A(n17132), .B(n25279), .Z(n17133) );
  NAND U21939 ( .A(n17134), .B(n17133), .Z(n17136) );
  ANDN U21940 ( .B(n17136), .A(n17135), .Z(n17137) );
  NAND U21941 ( .A(n17137), .B(n25283), .Z(n17138) );
  AND U21942 ( .A(n17139), .B(n17138), .Z(n17140) );
  NAND U21943 ( .A(n17140), .B(n25290), .Z(n17141) );
  NAND U21944 ( .A(n17142), .B(n17141), .Z(n17143) );
  NANDN U21945 ( .A(n25293), .B(n17143), .Z(n17144) );
  AND U21946 ( .A(n25295), .B(n17144), .Z(n17145) );
  ANDN U21947 ( .B(n25298), .A(n17145), .Z(n17147) );
  NAND U21948 ( .A(n17147), .B(n17146), .Z(n17148) );
  AND U21949 ( .A(n25299), .B(n17148), .Z(n17149) );
  NAND U21950 ( .A(n17150), .B(n17149), .Z(n17151) );
  NAND U21951 ( .A(n17152), .B(n17151), .Z(n17153) );
  NAND U21952 ( .A(n17154), .B(n17153), .Z(n17155) );
  NAND U21953 ( .A(n17155), .B(n25309), .Z(n17157) );
  NANDN U21954 ( .A(n17157), .B(n17156), .Z(n17160) );
  NOR U21955 ( .A(n17159), .B(n17158), .Z(n25311) );
  NAND U21956 ( .A(n17160), .B(n25311), .Z(n17161) );
  NANDN U21957 ( .A(n25313), .B(n17161), .Z(n17162) );
  AND U21958 ( .A(n25315), .B(n17162), .Z(n17163) );
  NANDN U21959 ( .A(n17163), .B(n25317), .Z(n17164) );
  AND U21960 ( .A(n25319), .B(n17164), .Z(n17165) );
  NANDN U21961 ( .A(n17165), .B(n25322), .Z(n17166) );
  AND U21962 ( .A(n25323), .B(n17166), .Z(n17167) );
  NANDN U21963 ( .A(n17167), .B(n25325), .Z(n17168) );
  AND U21964 ( .A(n25327), .B(n17168), .Z(n17169) );
  OR U21965 ( .A(n17169), .B(n25329), .Z(n17170) );
  NAND U21966 ( .A(n17170), .B(n25331), .Z(n17171) );
  ANDN U21967 ( .B(n17171), .A(n25334), .Z(n17172) );
  NANDN U21968 ( .A(n17172), .B(n25335), .Z(n17173) );
  ANDN U21969 ( .B(n17173), .A(n25338), .Z(n17174) );
  NANDN U21970 ( .A(n17174), .B(n25339), .Z(n17175) );
  NANDN U21971 ( .A(n17176), .B(n17175), .Z(n17177) );
  NANDN U21972 ( .A(n17178), .B(n17177), .Z(n17180) );
  NANDN U21973 ( .A(n17180), .B(n17179), .Z(n17181) );
  NAND U21974 ( .A(n17181), .B(n25346), .Z(n17183) );
  NANDN U21975 ( .A(n17183), .B(x[2576]), .Z(n17186) );
  XOR U21976 ( .A(n17183), .B(n17182), .Z(n17184) );
  NANDN U21977 ( .A(y[2576]), .B(n17184), .Z(n17185) );
  NAND U21978 ( .A(n17186), .B(n17185), .Z(n17187) );
  NANDN U21979 ( .A(n17187), .B(n25356), .Z(n17189) );
  ANDN U21980 ( .B(n17189), .A(n17188), .Z(n17190) );
  NAND U21981 ( .A(n17190), .B(n25357), .Z(n17191) );
  AND U21982 ( .A(n17192), .B(n17191), .Z(n17193) );
  OR U21983 ( .A(n25362), .B(n17193), .Z(n17196) );
  NOR U21984 ( .A(n25363), .B(n17194), .Z(n17195) );
  NAND U21985 ( .A(n17196), .B(n17195), .Z(n17197) );
  NAND U21986 ( .A(n17197), .B(n25365), .Z(n17198) );
  NANDN U21987 ( .A(n17199), .B(n17198), .Z(n17200) );
  NAND U21988 ( .A(n17200), .B(n25369), .Z(n17202) );
  NAND U21989 ( .A(n17202), .B(n17201), .Z(n17204) );
  NANDN U21990 ( .A(y[2584]), .B(n17204), .Z(n17203) );
  AND U21991 ( .A(n25375), .B(n17203), .Z(n17207) );
  XNOR U21992 ( .A(y[2584]), .B(n17204), .Z(n17205) );
  NAND U21993 ( .A(x[2584]), .B(n17205), .Z(n17206) );
  NAND U21994 ( .A(n17207), .B(n17206), .Z(n17208) );
  NAND U21995 ( .A(n17209), .B(n17208), .Z(n17210) );
  NANDN U21996 ( .A(n20243), .B(n17210), .Z(n17212) );
  NAND U21997 ( .A(n17212), .B(n17211), .Z(n17214) );
  ANDN U21998 ( .B(n17214), .A(n17213), .Z(n17215) );
  NAND U21999 ( .A(n17215), .B(n20244), .Z(n17217) );
  NAND U22000 ( .A(n17217), .B(n17216), .Z(n17219) );
  NANDN U22001 ( .A(n17219), .B(n17218), .Z(n17220) );
  AND U22002 ( .A(n17221), .B(n17220), .Z(n17222) );
  NAND U22003 ( .A(n17223), .B(n17222), .Z(n17224) );
  NAND U22004 ( .A(n17225), .B(n17224), .Z(n17226) );
  NANDN U22005 ( .A(n17227), .B(n17226), .Z(n17229) );
  NANDN U22006 ( .A(n17229), .B(y[2593]), .Z(n17232) );
  XOR U22007 ( .A(n17229), .B(n17228), .Z(n17230) );
  NANDN U22008 ( .A(x[2593]), .B(n17230), .Z(n17231) );
  AND U22009 ( .A(n17232), .B(n17231), .Z(n17236) );
  NANDN U22010 ( .A(n17236), .B(n17235), .Z(n17233) );
  AND U22011 ( .A(n17234), .B(n17233), .Z(n17239) );
  XNOR U22012 ( .A(n17236), .B(n17235), .Z(n17237) );
  NAND U22013 ( .A(n17237), .B(y[2594]), .Z(n17238) );
  NAND U22014 ( .A(n17239), .B(n17238), .Z(n17240) );
  NANDN U22015 ( .A(n17241), .B(n17240), .Z(n17242) );
  NAND U22016 ( .A(n17242), .B(n25397), .Z(n17243) );
  AND U22017 ( .A(n25399), .B(n17243), .Z(n17244) );
  NANDN U22018 ( .A(n17245), .B(n17244), .Z(n17249) );
  NAND U22019 ( .A(n17246), .B(y[2598]), .Z(n17248) );
  ANDN U22020 ( .B(n17248), .A(n17247), .Z(n25402) );
  NAND U22021 ( .A(n17249), .B(n25402), .Z(n17250) );
  AND U22022 ( .A(n25403), .B(n17250), .Z(n17251) );
  OR U22023 ( .A(n25406), .B(n17251), .Z(n17252) );
  AND U22024 ( .A(n25407), .B(n17252), .Z(n17253) );
  OR U22025 ( .A(n25409), .B(n17253), .Z(n17254) );
  AND U22026 ( .A(n25411), .B(n17254), .Z(n17255) );
  OR U22027 ( .A(n17255), .B(n25414), .Z(n17256) );
  AND U22028 ( .A(n25415), .B(n17256), .Z(n17257) );
  OR U22029 ( .A(n17257), .B(n25418), .Z(n17258) );
  AND U22030 ( .A(n25419), .B(n17258), .Z(n17259) );
  OR U22031 ( .A(n17259), .B(n25421), .Z(n17260) );
  AND U22032 ( .A(n25423), .B(n17260), .Z(n17261) );
  OR U22033 ( .A(n17261), .B(n25425), .Z(n17262) );
  NAND U22034 ( .A(n17263), .B(n17262), .Z(n17264) );
  NANDN U22035 ( .A(n25429), .B(n17264), .Z(n17265) );
  NANDN U22036 ( .A(n17265), .B(x[2612]), .Z(n17269) );
  XNOR U22037 ( .A(n17265), .B(x[2612]), .Z(n17266) );
  NAND U22038 ( .A(n17267), .B(n17266), .Z(n17268) );
  AND U22039 ( .A(n17269), .B(n17268), .Z(n17270) );
  OR U22040 ( .A(n17270), .B(y[2613]), .Z(n17273) );
  XOR U22041 ( .A(y[2613]), .B(n17270), .Z(n17271) );
  NAND U22042 ( .A(n17271), .B(x[2613]), .Z(n17272) );
  NAND U22043 ( .A(n17273), .B(n17272), .Z(n17274) );
  AND U22044 ( .A(n25438), .B(n17274), .Z(n17275) );
  ANDN U22045 ( .B(n25439), .A(n17275), .Z(n17277) );
  NAND U22046 ( .A(n17277), .B(n17276), .Z(n17278) );
  ANDN U22047 ( .B(n17278), .A(n25441), .Z(n17279) );
  NANDN U22048 ( .A(n17279), .B(n25443), .Z(n17282) );
  ANDN U22049 ( .B(n25445), .A(n17280), .Z(n17281) );
  NAND U22050 ( .A(n17282), .B(n17281), .Z(n17283) );
  NANDN U22051 ( .A(n17284), .B(n17283), .Z(n17285) );
  NAND U22052 ( .A(n17286), .B(n17285), .Z(n17288) );
  NAND U22053 ( .A(n17288), .B(n17287), .Z(n17289) );
  AND U22054 ( .A(n17290), .B(n17289), .Z(n17291) );
  OR U22055 ( .A(n25464), .B(n17291), .Z(n17294) );
  AND U22056 ( .A(n25466), .B(n17292), .Z(n17293) );
  NAND U22057 ( .A(n17294), .B(n17293), .Z(n17296) );
  NAND U22058 ( .A(n17296), .B(n17295), .Z(n17297) );
  NANDN U22059 ( .A(n17297), .B(n25467), .Z(n17298) );
  AND U22060 ( .A(n17299), .B(n17298), .Z(n17300) );
  ANDN U22061 ( .B(n17301), .A(n17300), .Z(n17303) );
  NAND U22062 ( .A(n17303), .B(n17302), .Z(n17304) );
  AND U22063 ( .A(n25478), .B(n17304), .Z(n17306) );
  AND U22064 ( .A(n17306), .B(n17305), .Z(n17307) );
  OR U22065 ( .A(n17308), .B(n17307), .Z(n17309) );
  NANDN U22066 ( .A(n25481), .B(n17309), .Z(n17310) );
  NAND U22067 ( .A(n17310), .B(n25483), .Z(n17311) );
  ANDN U22068 ( .B(n17311), .A(n25486), .Z(n17312) );
  NANDN U22069 ( .A(n17312), .B(n25487), .Z(n17313) );
  NAND U22070 ( .A(n17313), .B(n25490), .Z(n17315) );
  NAND U22071 ( .A(n17315), .B(n17314), .Z(n17316) );
  NAND U22072 ( .A(n17316), .B(n25493), .Z(n17317) );
  AND U22073 ( .A(n17318), .B(n17317), .Z(n17321) );
  AND U22074 ( .A(n17320), .B(n17319), .Z(n20242) );
  NANDN U22075 ( .A(n17321), .B(n20242), .Z(n17324) );
  ANDN U22076 ( .B(n20241), .A(n17322), .Z(n17323) );
  NAND U22077 ( .A(n17324), .B(n17323), .Z(n17326) );
  NAND U22078 ( .A(n17326), .B(n17325), .Z(n17327) );
  NANDN U22079 ( .A(n17327), .B(n25498), .Z(n17328) );
  NAND U22080 ( .A(n17329), .B(n17328), .Z(n17330) );
  NAND U22081 ( .A(n17331), .B(n17330), .Z(n17333) );
  NAND U22082 ( .A(n17333), .B(n17332), .Z(n17334) );
  NANDN U22083 ( .A(n17334), .B(n25510), .Z(n17335) );
  AND U22084 ( .A(n25511), .B(n17335), .Z(n17336) );
  OR U22085 ( .A(n25514), .B(n17336), .Z(n17339) );
  NANDN U22086 ( .A(x[2645]), .B(y[2645]), .Z(n17338) );
  ANDN U22087 ( .B(n17338), .A(n17337), .Z(n25515) );
  NAND U22088 ( .A(n17339), .B(n25515), .Z(n17340) );
  AND U22089 ( .A(n25517), .B(n17340), .Z(n17341) );
  NANDN U22090 ( .A(n17341), .B(n25519), .Z(n17342) );
  NAND U22091 ( .A(n17342), .B(n25522), .Z(n17343) );
  NAND U22092 ( .A(n17343), .B(n25523), .Z(n17344) );
  AND U22093 ( .A(n25526), .B(n17344), .Z(n17345) );
  OR U22094 ( .A(n25528), .B(n17345), .Z(n17346) );
  NANDN U22095 ( .A(n25530), .B(n17346), .Z(n17347) );
  NAND U22096 ( .A(n17347), .B(n25531), .Z(n17349) );
  NANDN U22097 ( .A(n17349), .B(n17348), .Z(n17350) );
  NANDN U22098 ( .A(n25534), .B(n17350), .Z(n17352) );
  NANDN U22099 ( .A(n17352), .B(y[2655]), .Z(n17355) );
  XOR U22100 ( .A(n17352), .B(n17351), .Z(n17353) );
  NANDN U22101 ( .A(x[2655]), .B(n17353), .Z(n17354) );
  NAND U22102 ( .A(n17355), .B(n17354), .Z(n17356) );
  NANDN U22103 ( .A(n17356), .B(n25540), .Z(n17357) );
  NAND U22104 ( .A(n17358), .B(n17357), .Z(n17359) );
  NANDN U22105 ( .A(n25544), .B(n17359), .Z(n17360) );
  AND U22106 ( .A(n25545), .B(n17360), .Z(n17361) );
  OR U22107 ( .A(n17362), .B(n17361), .Z(n17363) );
  NAND U22108 ( .A(n17364), .B(n17363), .Z(n17365) );
  NAND U22109 ( .A(n17366), .B(n17365), .Z(n17367) );
  NAND U22110 ( .A(n17367), .B(n25557), .Z(n17369) );
  NANDN U22111 ( .A(n17369), .B(n17368), .Z(n17371) );
  ANDN U22112 ( .B(n17371), .A(n17370), .Z(n17372) );
  NAND U22113 ( .A(n17372), .B(n25559), .Z(n17373) );
  AND U22114 ( .A(n25561), .B(n17373), .Z(n17374) );
  OR U22115 ( .A(n25563), .B(n17374), .Z(n17377) );
  ANDN U22116 ( .B(n25565), .A(n17375), .Z(n17376) );
  NAND U22117 ( .A(n17377), .B(n17376), .Z(n17379) );
  NAND U22118 ( .A(n17379), .B(n17378), .Z(n17380) );
  NANDN U22119 ( .A(n17380), .B(n25567), .Z(n17381) );
  NAND U22120 ( .A(n17382), .B(n17381), .Z(n17383) );
  NAND U22121 ( .A(n17384), .B(n17383), .Z(n17386) );
  NAND U22122 ( .A(n17386), .B(n17385), .Z(n17387) );
  NANDN U22123 ( .A(n17387), .B(n25577), .Z(n17390) );
  OR U22124 ( .A(n17389), .B(n17388), .Z(n25579) );
  ANDN U22125 ( .B(n17390), .A(n25579), .Z(n17391) );
  OR U22126 ( .A(n25581), .B(n17391), .Z(n17394) );
  AND U22127 ( .A(n25583), .B(n17392), .Z(n17393) );
  NAND U22128 ( .A(n17394), .B(n17393), .Z(n17395) );
  NANDN U22129 ( .A(n25585), .B(n17395), .Z(n17397) );
  ANDN U22130 ( .B(n17397), .A(n17396), .Z(n17398) );
  NAND U22131 ( .A(n17399), .B(n17398), .Z(n17400) );
  NAND U22132 ( .A(n17400), .B(n25589), .Z(n17401) );
  AND U22133 ( .A(n25591), .B(n17401), .Z(n17402) );
  OR U22134 ( .A(n25594), .B(n17402), .Z(n17403) );
  NANDN U22135 ( .A(n25595), .B(n17403), .Z(n17405) );
  NAND U22136 ( .A(n17405), .B(n17404), .Z(n17406) );
  NANDN U22137 ( .A(n17406), .B(n25597), .Z(n17407) );
  NAND U22138 ( .A(n17407), .B(n25600), .Z(n17408) );
  NANDN U22139 ( .A(n17409), .B(n17408), .Z(n17410) );
  ANDN U22140 ( .B(n17410), .A(n25603), .Z(n17411) );
  OR U22141 ( .A(n25606), .B(n17411), .Z(n17412) );
  NAND U22142 ( .A(n17412), .B(n25607), .Z(n17414) );
  NAND U22143 ( .A(n17414), .B(n17413), .Z(n17416) );
  ANDN U22144 ( .B(n17416), .A(n17415), .Z(n17418) );
  NANDN U22145 ( .A(n17418), .B(n17417), .Z(n17419) );
  AND U22146 ( .A(n25623), .B(n17419), .Z(n17420) );
  NANDN U22147 ( .A(n17420), .B(n25624), .Z(n17421) );
  NAND U22148 ( .A(n17421), .B(n25626), .Z(n17422) );
  AND U22149 ( .A(n25628), .B(n17422), .Z(n17423) );
  NANDN U22150 ( .A(n17423), .B(n25630), .Z(n17425) );
  ANDN U22151 ( .B(n17425), .A(n17424), .Z(n17428) );
  NOR U22152 ( .A(n17427), .B(n17426), .Z(n25635) );
  NANDN U22153 ( .A(n17428), .B(n25635), .Z(n17431) );
  ANDN U22154 ( .B(n25634), .A(n17429), .Z(n17430) );
  NAND U22155 ( .A(n17431), .B(n17430), .Z(n17433) );
  NAND U22156 ( .A(n17433), .B(n17432), .Z(n17434) );
  NANDN U22157 ( .A(n17434), .B(n25637), .Z(n17435) );
  NAND U22158 ( .A(n17436), .B(n17435), .Z(n17437) );
  NAND U22159 ( .A(n17438), .B(n17437), .Z(n17440) );
  NAND U22160 ( .A(n17440), .B(n17439), .Z(n17441) );
  NANDN U22161 ( .A(n17441), .B(n25648), .Z(n17442) );
  ANDN U22162 ( .B(n17442), .A(n25650), .Z(n17443) );
  NANDN U22163 ( .A(n17443), .B(n25652), .Z(n17444) );
  NAND U22164 ( .A(n17444), .B(n25654), .Z(n17445) );
  NAND U22165 ( .A(n17445), .B(n25656), .Z(n17446) );
  ANDN U22166 ( .B(n17446), .A(n25658), .Z(n17447) );
  ANDN U22167 ( .B(n25661), .A(n17447), .Z(n17448) );
  NANDN U22168 ( .A(n17448), .B(n25664), .Z(n17450) );
  NAND U22169 ( .A(n17450), .B(n17449), .Z(n17451) );
  NAND U22170 ( .A(n17451), .B(n25674), .Z(n17452) );
  OR U22171 ( .A(n17453), .B(n17452), .Z(n17454) );
  NANDN U22172 ( .A(n25677), .B(n17454), .Z(n17455) );
  AND U22173 ( .A(n17456), .B(n17455), .Z(n17457) );
  OR U22174 ( .A(n17457), .B(n25681), .Z(n17458) );
  AND U22175 ( .A(n17459), .B(n17458), .Z(n17460) );
  NANDN U22176 ( .A(n17460), .B(n25685), .Z(n17462) );
  ANDN U22177 ( .B(n17462), .A(n17461), .Z(n17466) );
  OR U22178 ( .A(n17464), .B(n17463), .Z(n20238) );
  IV U22179 ( .A(n20238), .Z(n17465) );
  NANDN U22180 ( .A(n17466), .B(n17465), .Z(n17469) );
  ANDN U22181 ( .B(n20237), .A(n17467), .Z(n17468) );
  NAND U22182 ( .A(n17469), .B(n17468), .Z(n17471) );
  NAND U22183 ( .A(n17471), .B(n17470), .Z(n17472) );
  NANDN U22184 ( .A(n17472), .B(n20240), .Z(n17473) );
  NAND U22185 ( .A(n17474), .B(n17473), .Z(n17475) );
  NANDN U22186 ( .A(n17476), .B(n17475), .Z(n17478) );
  XNOR U22187 ( .A(y[2719]), .B(n17478), .Z(n17477) );
  NANDN U22188 ( .A(x[2719]), .B(n17477), .Z(n17480) );
  NANDN U22189 ( .A(n17478), .B(y[2719]), .Z(n17479) );
  NAND U22190 ( .A(n17480), .B(n17479), .Z(n17482) );
  NANDN U22191 ( .A(n17482), .B(x[2720]), .Z(n17485) );
  XOR U22192 ( .A(n17482), .B(n17481), .Z(n17483) );
  NANDN U22193 ( .A(y[2720]), .B(n17483), .Z(n17484) );
  NAND U22194 ( .A(n17485), .B(n17484), .Z(n17487) );
  NANDN U22195 ( .A(n17487), .B(n17486), .Z(n17488) );
  NANDN U22196 ( .A(n17489), .B(n17488), .Z(n17491) );
  NAND U22197 ( .A(n17491), .B(n17490), .Z(n17492) );
  OR U22198 ( .A(n17493), .B(n17492), .Z(n17494) );
  NANDN U22199 ( .A(n25703), .B(n17494), .Z(n17496) );
  NANDN U22200 ( .A(n17496), .B(x[2724]), .Z(n17499) );
  XOR U22201 ( .A(n17496), .B(n17495), .Z(n17497) );
  NANDN U22202 ( .A(y[2724]), .B(n17497), .Z(n17498) );
  NAND U22203 ( .A(n17499), .B(n17498), .Z(n17501) );
  NANDN U22204 ( .A(n17501), .B(n17500), .Z(n17502) );
  AND U22205 ( .A(n17503), .B(n17502), .Z(n17504) );
  OR U22206 ( .A(n17505), .B(n17504), .Z(n17508) );
  ANDN U22207 ( .B(n17507), .A(n17506), .Z(n25714) );
  NAND U22208 ( .A(n17508), .B(n25714), .Z(n17509) );
  NANDN U22209 ( .A(n25716), .B(n17509), .Z(n17510) );
  NAND U22210 ( .A(n17511), .B(n17510), .Z(n17512) );
  AND U22211 ( .A(n25721), .B(n17512), .Z(n17513) );
  NAND U22212 ( .A(n17514), .B(n17513), .Z(n17515) );
  NAND U22213 ( .A(n17516), .B(n17515), .Z(n17517) );
  NAND U22214 ( .A(n17518), .B(n17517), .Z(n17520) );
  NAND U22215 ( .A(n17520), .B(n17519), .Z(n17521) );
  NANDN U22216 ( .A(n17521), .B(n25730), .Z(n17524) );
  NANDN U22217 ( .A(y[2735]), .B(x[2735]), .Z(n17522) );
  NANDN U22218 ( .A(n17523), .B(n17522), .Z(n25732) );
  ANDN U22219 ( .B(n17524), .A(n25732), .Z(n17525) );
  OR U22220 ( .A(n25735), .B(n17525), .Z(n17526) );
  NANDN U22221 ( .A(n25737), .B(n17526), .Z(n17528) );
  NAND U22222 ( .A(n17528), .B(n17527), .Z(n17529) );
  NANDN U22223 ( .A(n17529), .B(n25738), .Z(n17530) );
  NANDN U22224 ( .A(n25741), .B(n17530), .Z(n17531) );
  NANDN U22225 ( .A(n17531), .B(y[2739]), .Z(n17535) );
  XNOR U22226 ( .A(n17531), .B(y[2739]), .Z(n17532) );
  NAND U22227 ( .A(n17533), .B(n17532), .Z(n17534) );
  NAND U22228 ( .A(n17535), .B(n17534), .Z(n17536) );
  NANDN U22229 ( .A(n17536), .B(n25746), .Z(n17537) );
  AND U22230 ( .A(n17538), .B(n17537), .Z(n17539) );
  NANDN U22231 ( .A(n17539), .B(n25750), .Z(n17540) );
  ANDN U22232 ( .B(n17540), .A(n25753), .Z(n17541) );
  ANDN U22233 ( .B(n25754), .A(n17541), .Z(n17543) );
  NAND U22234 ( .A(n17543), .B(n17542), .Z(n17544) );
  AND U22235 ( .A(n25757), .B(n17544), .Z(n17545) );
  NAND U22236 ( .A(n17546), .B(n17545), .Z(n17547) );
  NAND U22237 ( .A(n17548), .B(n17547), .Z(n17549) );
  NAND U22238 ( .A(n17550), .B(n17549), .Z(n17552) );
  NAND U22239 ( .A(n17552), .B(n17551), .Z(n17553) );
  NANDN U22240 ( .A(n17553), .B(n25766), .Z(n17556) );
  NANDN U22241 ( .A(n17555), .B(n17554), .Z(n25768) );
  ANDN U22242 ( .B(n17556), .A(n25768), .Z(n17557) );
  OR U22243 ( .A(n25771), .B(n17557), .Z(n17558) );
  NANDN U22244 ( .A(n25773), .B(n17558), .Z(n17559) );
  NANDN U22245 ( .A(n25775), .B(n17559), .Z(n17560) );
  NAND U22246 ( .A(n17561), .B(n17560), .Z(n17562) );
  AND U22247 ( .A(n25778), .B(n17562), .Z(n17563) );
  NAND U22248 ( .A(n17563), .B(n25783), .Z(n17564) );
  AND U22249 ( .A(n17565), .B(n17564), .Z(n17566) );
  NAND U22250 ( .A(n17566), .B(n25784), .Z(n17567) );
  NANDN U22251 ( .A(n25787), .B(n17567), .Z(n17568) );
  NANDN U22252 ( .A(n25789), .B(n17568), .Z(n17569) );
  AND U22253 ( .A(n17570), .B(n17569), .Z(n17571) );
  OR U22254 ( .A(n17572), .B(n17571), .Z(n17573) );
  NAND U22255 ( .A(n17574), .B(n17573), .Z(n17575) );
  NAND U22256 ( .A(n17576), .B(n17575), .Z(n17577) );
  NAND U22257 ( .A(n17577), .B(n25803), .Z(n17579) );
  NANDN U22258 ( .A(n17579), .B(n17578), .Z(n17582) );
  ANDN U22259 ( .B(n25804), .A(n17580), .Z(n17581) );
  NAND U22260 ( .A(n17582), .B(n17581), .Z(n17583) );
  NANDN U22261 ( .A(n25807), .B(n17583), .Z(n17584) );
  NAND U22262 ( .A(n17585), .B(n17584), .Z(n17586) );
  NAND U22263 ( .A(n17586), .B(n25810), .Z(n17587) );
  NAND U22264 ( .A(n17588), .B(n17587), .Z(n17589) );
  NAND U22265 ( .A(n17590), .B(n17589), .Z(n17591) );
  NAND U22266 ( .A(n17592), .B(n17591), .Z(n17593) );
  NAND U22267 ( .A(n17594), .B(n17593), .Z(n17595) );
  NAND U22268 ( .A(n17596), .B(n17595), .Z(n17598) );
  NAND U22269 ( .A(n17598), .B(n17597), .Z(n17599) );
  NANDN U22270 ( .A(n17599), .B(n25822), .Z(n17604) );
  NANDN U22271 ( .A(n17601), .B(n17600), .Z(n17602) );
  NANDN U22272 ( .A(n17603), .B(n17602), .Z(n25825) );
  ANDN U22273 ( .B(n17604), .A(n25825), .Z(n17605) );
  NANDN U22274 ( .A(n17605), .B(n25827), .Z(n17606) );
  AND U22275 ( .A(n25828), .B(n17606), .Z(n17607) );
  NANDN U22276 ( .A(n17607), .B(n25831), .Z(n17609) );
  ANDN U22277 ( .B(n17609), .A(n17608), .Z(n17610) );
  NANDN U22278 ( .A(n17610), .B(n25835), .Z(n17611) );
  AND U22279 ( .A(n25838), .B(n17611), .Z(n17612) );
  NANDN U22280 ( .A(n17612), .B(n25841), .Z(n17613) );
  AND U22281 ( .A(n25842), .B(n17613), .Z(n17614) );
  NANDN U22282 ( .A(n17614), .B(n25844), .Z(n17615) );
  AND U22283 ( .A(n25846), .B(n17615), .Z(n17616) );
  NANDN U22284 ( .A(n17616), .B(n25849), .Z(n17620) );
  NAND U22285 ( .A(n17617), .B(x[2785]), .Z(n17619) );
  ANDN U22286 ( .B(n17619), .A(n17618), .Z(n25850) );
  NAND U22287 ( .A(n17620), .B(n25850), .Z(n17621) );
  NANDN U22288 ( .A(n25852), .B(n17621), .Z(n17623) );
  NAND U22289 ( .A(n17623), .B(n17622), .Z(n17625) );
  ANDN U22290 ( .B(n17625), .A(n17624), .Z(n17627) );
  NANDN U22291 ( .A(n17627), .B(n17626), .Z(n17628) );
  ANDN U22292 ( .B(n17628), .A(n25868), .Z(n17629) );
  NANDN U22293 ( .A(n17629), .B(n25869), .Z(n17630) );
  ANDN U22294 ( .B(n17630), .A(n25872), .Z(n17631) );
  NANDN U22295 ( .A(n17631), .B(n25873), .Z(n17632) );
  AND U22296 ( .A(n17633), .B(n17632), .Z(n17634) );
  NAND U22297 ( .A(n17634), .B(n25876), .Z(n17635) );
  AND U22298 ( .A(n17636), .B(n17635), .Z(n17637) );
  NAND U22299 ( .A(n17637), .B(n25877), .Z(n17638) );
  NAND U22300 ( .A(n17639), .B(n17638), .Z(n17641) );
  NAND U22301 ( .A(n17641), .B(n17640), .Z(n17642) );
  NANDN U22302 ( .A(n17642), .B(n25885), .Z(n17645) );
  NANDN U22303 ( .A(n17644), .B(n17643), .Z(n25887) );
  ANDN U22304 ( .B(n17645), .A(n25887), .Z(n17646) );
  OR U22305 ( .A(n25889), .B(n17646), .Z(n17648) );
  ANDN U22306 ( .B(n17648), .A(n17647), .Z(n17649) );
  NAND U22307 ( .A(n17649), .B(n25892), .Z(n17651) );
  ANDN U22308 ( .B(n17651), .A(n17650), .Z(n17652) );
  NAND U22309 ( .A(n17652), .B(n25893), .Z(n17653) );
  AND U22310 ( .A(n17654), .B(n17653), .Z(n17656) );
  NAND U22311 ( .A(n17656), .B(n17655), .Z(n17657) );
  NAND U22312 ( .A(n17658), .B(n17657), .Z(n17659) );
  NAND U22313 ( .A(n17659), .B(n25903), .Z(n17661) );
  NANDN U22314 ( .A(n17661), .B(n17660), .Z(n17662) );
  NANDN U22315 ( .A(n25906), .B(n17662), .Z(n17663) );
  NANDN U22316 ( .A(n25908), .B(n17663), .Z(n17664) );
  NAND U22317 ( .A(n17665), .B(n17664), .Z(n17666) );
  NAND U22318 ( .A(n17667), .B(n17666), .Z(n17668) );
  NANDN U22319 ( .A(n17668), .B(n25911), .Z(n17669) );
  NAND U22320 ( .A(n17670), .B(n17669), .Z(n17671) );
  NAND U22321 ( .A(n17672), .B(n17671), .Z(n17673) );
  NANDN U22322 ( .A(n17674), .B(n17673), .Z(n17675) );
  AND U22323 ( .A(n25923), .B(n17675), .Z(n17677) );
  NANDN U22324 ( .A(n17677), .B(n17676), .Z(n17678) );
  NANDN U22325 ( .A(n17679), .B(n17678), .Z(n17681) );
  NAND U22326 ( .A(n17681), .B(n17680), .Z(n17683) );
  ANDN U22327 ( .B(n25938), .A(n17682), .Z(n25933) );
  NAND U22328 ( .A(n17683), .B(n25933), .Z(n17686) );
  OR U22329 ( .A(n17685), .B(n17684), .Z(n25943) );
  ANDN U22330 ( .B(n17686), .A(n25943), .Z(n17687) );
  OR U22331 ( .A(n25944), .B(n17687), .Z(n17690) );
  NOR U22332 ( .A(n17689), .B(n17688), .Z(n25946) );
  NAND U22333 ( .A(n17690), .B(n25946), .Z(n17692) );
  NAND U22334 ( .A(n17692), .B(n17691), .Z(n17693) );
  NANDN U22335 ( .A(n17693), .B(n25948), .Z(n17694) );
  NAND U22336 ( .A(n17695), .B(n17694), .Z(n17696) );
  NAND U22337 ( .A(n17697), .B(n17696), .Z(n17699) );
  NAND U22338 ( .A(n17699), .B(n17698), .Z(n17700) );
  NANDN U22339 ( .A(n17700), .B(n25958), .Z(n17701) );
  AND U22340 ( .A(n25960), .B(n17701), .Z(n17702) );
  NANDN U22341 ( .A(n17702), .B(n25962), .Z(n17703) );
  AND U22342 ( .A(n17704), .B(n17703), .Z(n17705) );
  OR U22343 ( .A(n17706), .B(n17705), .Z(n17708) );
  NAND U22344 ( .A(n17708), .B(n17707), .Z(n17710) );
  NAND U22345 ( .A(n17710), .B(n17709), .Z(n17712) );
  ANDN U22346 ( .B(n25982), .A(n17711), .Z(n25977) );
  NAND U22347 ( .A(n17712), .B(n25977), .Z(n17713) );
  AND U22348 ( .A(n25980), .B(n17713), .Z(n17714) );
  ANDN U22349 ( .B(n25987), .A(n17714), .Z(n17716) );
  NAND U22350 ( .A(n17716), .B(n17715), .Z(n17717) );
  AND U22351 ( .A(n25988), .B(n17717), .Z(n17718) );
  NAND U22352 ( .A(n17719), .B(n17718), .Z(n17720) );
  NAND U22353 ( .A(n17721), .B(n17720), .Z(n17722) );
  NANDN U22354 ( .A(n17723), .B(n17722), .Z(n17725) );
  NANDN U22355 ( .A(n17725), .B(y[2837]), .Z(n17728) );
  XOR U22356 ( .A(n17725), .B(n17724), .Z(n17726) );
  NANDN U22357 ( .A(x[2837]), .B(n17726), .Z(n17727) );
  NAND U22358 ( .A(n17728), .B(n17727), .Z(n17729) );
  NANDN U22359 ( .A(n17729), .B(n25999), .Z(n17731) );
  ANDN U22360 ( .B(n17731), .A(n17730), .Z(n17732) );
  NAND U22361 ( .A(n17732), .B(n26000), .Z(n17735) );
  NANDN U22362 ( .A(x[2840]), .B(y[2840]), .Z(n17733) );
  NANDN U22363 ( .A(n17734), .B(n17733), .Z(n26002) );
  ANDN U22364 ( .B(n17735), .A(n26002), .Z(n17738) );
  ANDN U22365 ( .B(n17737), .A(n17736), .Z(n26004) );
  NANDN U22366 ( .A(n17738), .B(n26004), .Z(n17739) );
  AND U22367 ( .A(n26007), .B(n17739), .Z(n17740) );
  NANDN U22368 ( .A(n17740), .B(n26008), .Z(n17741) );
  ANDN U22369 ( .B(n17741), .A(n26010), .Z(n17742) );
  NANDN U22370 ( .A(n17742), .B(n26012), .Z(n17743) );
  NANDN U22371 ( .A(n26014), .B(n17743), .Z(n17744) );
  NAND U22372 ( .A(n17744), .B(n26016), .Z(n17745) );
  AND U22373 ( .A(n26019), .B(n17745), .Z(n17746) );
  NANDN U22374 ( .A(n17746), .B(n26020), .Z(n17747) );
  NANDN U22375 ( .A(n26023), .B(n17747), .Z(n17748) );
  AND U22376 ( .A(n17749), .B(n17748), .Z(n17750) );
  NAND U22377 ( .A(n17750), .B(n26025), .Z(n17751) );
  AND U22378 ( .A(n17752), .B(n17751), .Z(n17753) );
  NAND U22379 ( .A(n17753), .B(n26026), .Z(n17754) );
  NAND U22380 ( .A(n17755), .B(n17754), .Z(n17756) );
  NAND U22381 ( .A(n17756), .B(n26034), .Z(n17758) );
  NANDN U22382 ( .A(n17758), .B(n17757), .Z(n17759) );
  AND U22383 ( .A(n17760), .B(n17759), .Z(n17761) );
  NAND U22384 ( .A(n17761), .B(n26036), .Z(n17762) );
  AND U22385 ( .A(n26038), .B(n17762), .Z(n17763) );
  OR U22386 ( .A(n26040), .B(n17763), .Z(n17764) );
  AND U22387 ( .A(n26042), .B(n17764), .Z(n17765) );
  NANDN U22388 ( .A(n17765), .B(n26044), .Z(n17766) );
  NAND U22389 ( .A(n17766), .B(n26046), .Z(n17767) );
  NAND U22390 ( .A(n17767), .B(n26050), .Z(n17768) );
  AND U22391 ( .A(n26052), .B(n17768), .Z(n17770) );
  NANDN U22392 ( .A(n17770), .B(n17769), .Z(n17771) );
  NAND U22393 ( .A(n17771), .B(n26056), .Z(n17772) );
  NAND U22394 ( .A(n17772), .B(n26058), .Z(n17775) );
  NOR U22395 ( .A(n17774), .B(n17773), .Z(n26060) );
  NAND U22396 ( .A(n17775), .B(n26060), .Z(n17778) );
  NOR U22397 ( .A(n17777), .B(n17776), .Z(n26063) );
  NAND U22398 ( .A(n17778), .B(n26063), .Z(n17779) );
  AND U22399 ( .A(n17780), .B(n17779), .Z(n17783) );
  NAND U22400 ( .A(n17781), .B(n26066), .Z(n17782) );
  OR U22401 ( .A(n17783), .B(n17782), .Z(n17784) );
  AND U22402 ( .A(n17785), .B(n17784), .Z(n17786) );
  OR U22403 ( .A(n17787), .B(n17786), .Z(n17788) );
  NANDN U22404 ( .A(n17789), .B(n17788), .Z(n17791) );
  NAND U22405 ( .A(n17791), .B(n17790), .Z(n17793) );
  NANDN U22406 ( .A(n17793), .B(n17792), .Z(n17794) );
  NAND U22407 ( .A(n17795), .B(n17794), .Z(n17796) );
  NANDN U22408 ( .A(n26080), .B(n17796), .Z(n17798) );
  XNOR U22409 ( .A(y[2871]), .B(n17798), .Z(n17797) );
  NANDN U22410 ( .A(x[2871]), .B(n17797), .Z(n17800) );
  NANDN U22411 ( .A(n17798), .B(y[2871]), .Z(n17799) );
  AND U22412 ( .A(n17800), .B(n17799), .Z(n17801) );
  NAND U22413 ( .A(n17802), .B(n17801), .Z(n17803) );
  NAND U22414 ( .A(n17804), .B(n17803), .Z(n17805) );
  NAND U22415 ( .A(n17806), .B(n17805), .Z(n17807) );
  NANDN U22416 ( .A(n26093), .B(n17807), .Z(n17811) );
  NAND U22417 ( .A(n17808), .B(y[2875]), .Z(n17809) );
  NANDN U22418 ( .A(n17810), .B(n17809), .Z(n26094) );
  ANDN U22419 ( .B(n17811), .A(n26094), .Z(n17812) );
  ANDN U22420 ( .B(n26096), .A(n17812), .Z(n17814) );
  NAND U22421 ( .A(n17814), .B(n17813), .Z(n17815) );
  AND U22422 ( .A(n26098), .B(n17815), .Z(n17816) );
  NAND U22423 ( .A(n17817), .B(n17816), .Z(n17818) );
  NAND U22424 ( .A(n17819), .B(n17818), .Z(n17820) );
  NAND U22425 ( .A(n17821), .B(n17820), .Z(n17822) );
  NAND U22426 ( .A(n17822), .B(n26108), .Z(n17824) );
  NANDN U22427 ( .A(n17824), .B(n17823), .Z(n17825) );
  NANDN U22428 ( .A(n26110), .B(n17825), .Z(n17826) );
  NANDN U22429 ( .A(n26112), .B(n17826), .Z(n17827) );
  NAND U22430 ( .A(n17828), .B(n17827), .Z(n17829) );
  ANDN U22431 ( .B(n17829), .A(n26116), .Z(n17835) );
  NANDN U22432 ( .A(n17831), .B(n17830), .Z(n17833) );
  ANDN U22433 ( .B(n17833), .A(n17832), .Z(n17834) );
  NANDN U22434 ( .A(n17835), .B(n17834), .Z(n17836) );
  NAND U22435 ( .A(n17836), .B(n26120), .Z(n17837) );
  NAND U22436 ( .A(n17837), .B(n26122), .Z(n17840) );
  ANDN U22437 ( .B(n17839), .A(n17838), .Z(n26124) );
  NAND U22438 ( .A(n17840), .B(n26124), .Z(n17841) );
  NANDN U22439 ( .A(n26126), .B(n17841), .Z(n17842) );
  AND U22440 ( .A(n17843), .B(n17842), .Z(n17844) );
  OR U22441 ( .A(n17845), .B(n17844), .Z(n17846) );
  NAND U22442 ( .A(n17847), .B(n17846), .Z(n17848) );
  NAND U22443 ( .A(n17849), .B(n17848), .Z(n17851) );
  NAND U22444 ( .A(n17851), .B(n17850), .Z(n17852) );
  NANDN U22445 ( .A(n17852), .B(n26140), .Z(n17855) );
  NANDN U22446 ( .A(n17854), .B(n17853), .Z(n26142) );
  ANDN U22447 ( .B(n17855), .A(n26142), .Z(n17856) );
  OR U22448 ( .A(n26144), .B(n17856), .Z(n17857) );
  AND U22449 ( .A(n26147), .B(n17857), .Z(n17859) );
  NAND U22450 ( .A(n17859), .B(n17858), .Z(n17860) );
  NAND U22451 ( .A(n17860), .B(n26148), .Z(n17862) );
  NANDN U22452 ( .A(n17862), .B(y[2899]), .Z(n17865) );
  XOR U22453 ( .A(n17862), .B(n17861), .Z(n17863) );
  NANDN U22454 ( .A(x[2899]), .B(n17863), .Z(n17864) );
  AND U22455 ( .A(n17865), .B(n17864), .Z(n17866) );
  OR U22456 ( .A(n17866), .B(x[2900]), .Z(n17869) );
  XOR U22457 ( .A(x[2900]), .B(n17866), .Z(n17867) );
  NAND U22458 ( .A(y[2900]), .B(n17867), .Z(n17868) );
  NAND U22459 ( .A(n17869), .B(n17868), .Z(n17870) );
  NAND U22460 ( .A(n17870), .B(n26156), .Z(n17871) );
  NAND U22461 ( .A(n17872), .B(n17871), .Z(n17873) );
  AND U22462 ( .A(n26160), .B(n17873), .Z(n17874) );
  OR U22463 ( .A(n26162), .B(n17874), .Z(n17877) );
  AND U22464 ( .A(n26164), .B(n17875), .Z(n17876) );
  NAND U22465 ( .A(n17877), .B(n17876), .Z(n17878) );
  NANDN U22466 ( .A(n26167), .B(n17878), .Z(n17879) );
  NAND U22467 ( .A(n17880), .B(n17879), .Z(n17881) );
  NAND U22468 ( .A(n17881), .B(n26170), .Z(n17882) );
  AND U22469 ( .A(n26172), .B(n17882), .Z(n17883) );
  NANDN U22470 ( .A(n17883), .B(n26175), .Z(n17884) );
  AND U22471 ( .A(n26176), .B(n17884), .Z(n17885) );
  OR U22472 ( .A(n17886), .B(n17885), .Z(n17887) );
  NANDN U22473 ( .A(n17888), .B(n17887), .Z(n17890) );
  NAND U22474 ( .A(n17890), .B(n17889), .Z(n17891) );
  OR U22475 ( .A(n17891), .B(n26189), .Z(n17893) );
  ANDN U22476 ( .B(n17893), .A(n17892), .Z(n17894) );
  NANDN U22477 ( .A(n17894), .B(n26193), .Z(n17895) );
  AND U22478 ( .A(n26194), .B(n17895), .Z(n17896) );
  OR U22479 ( .A(n26197), .B(n17896), .Z(n17897) );
  AND U22480 ( .A(n26198), .B(n17897), .Z(n17899) );
  NAND U22481 ( .A(n17899), .B(n17898), .Z(n17900) );
  NANDN U22482 ( .A(n26201), .B(n17900), .Z(n17902) );
  NANDN U22483 ( .A(n17902), .B(x[2920]), .Z(n17905) );
  XOR U22484 ( .A(n17902), .B(n17901), .Z(n17903) );
  NANDN U22485 ( .A(y[2920]), .B(n17903), .Z(n17904) );
  AND U22486 ( .A(n17905), .B(n17904), .Z(n17906) );
  OR U22487 ( .A(n17906), .B(y[2921]), .Z(n17909) );
  XOR U22488 ( .A(y[2921]), .B(n17906), .Z(n17907) );
  NAND U22489 ( .A(x[2921]), .B(n17907), .Z(n17908) );
  NAND U22490 ( .A(n17909), .B(n17908), .Z(n17910) );
  NAND U22491 ( .A(n17910), .B(n26209), .Z(n17911) );
  NAND U22492 ( .A(n17912), .B(n17911), .Z(n17915) );
  NANDN U22493 ( .A(n17914), .B(n17913), .Z(n26212) );
  ANDN U22494 ( .B(n17915), .A(n26212), .Z(n17916) );
  OR U22495 ( .A(n26214), .B(n17916), .Z(n17919) );
  AND U22496 ( .A(n26217), .B(n17917), .Z(n17918) );
  NAND U22497 ( .A(n17919), .B(n17918), .Z(n17921) );
  NAND U22498 ( .A(n17921), .B(n17920), .Z(n17922) );
  NANDN U22499 ( .A(n17922), .B(n26218), .Z(n17923) );
  NAND U22500 ( .A(n17924), .B(n17923), .Z(n17925) );
  NAND U22501 ( .A(n17926), .B(n17925), .Z(n17927) );
  NAND U22502 ( .A(n17927), .B(n26228), .Z(n17929) );
  NANDN U22503 ( .A(n17929), .B(n17928), .Z(n17932) );
  ANDN U22504 ( .B(n26230), .A(n17930), .Z(n17931) );
  NAND U22505 ( .A(n17932), .B(n17931), .Z(n17933) );
  NANDN U22506 ( .A(n26232), .B(n17933), .Z(n17934) );
  NAND U22507 ( .A(n17935), .B(n17934), .Z(n17937) );
  NAND U22508 ( .A(n17937), .B(n17936), .Z(n17938) );
  NANDN U22509 ( .A(n17938), .B(n26236), .Z(n17939) );
  NAND U22510 ( .A(n17940), .B(n17939), .Z(n17941) );
  NANDN U22511 ( .A(n17941), .B(y[2935]), .Z(n17945) );
  XNOR U22512 ( .A(n17941), .B(y[2935]), .Z(n17942) );
  NAND U22513 ( .A(n17943), .B(n17942), .Z(n17944) );
  NAND U22514 ( .A(n17945), .B(n17944), .Z(n17946) );
  NANDN U22515 ( .A(n17946), .B(n26244), .Z(n17947) );
  NAND U22516 ( .A(n17948), .B(n17947), .Z(n17951) );
  NOR U22517 ( .A(n17950), .B(n17949), .Z(n26248) );
  NAND U22518 ( .A(n17951), .B(n26248), .Z(n17954) );
  NANDN U22519 ( .A(n17953), .B(n17952), .Z(n26251) );
  ANDN U22520 ( .B(n17954), .A(n26251), .Z(n17955) );
  NANDN U22521 ( .A(n17955), .B(n26252), .Z(n17958) );
  AND U22522 ( .A(n26254), .B(n17956), .Z(n17957) );
  NAND U22523 ( .A(n17958), .B(n17957), .Z(n17960) );
  NAND U22524 ( .A(n17960), .B(n17959), .Z(n17961) );
  NANDN U22525 ( .A(n17961), .B(n26256), .Z(n17962) );
  NAND U22526 ( .A(n17963), .B(n17962), .Z(n17964) );
  NAND U22527 ( .A(n17965), .B(n17964), .Z(n17966) );
  NANDN U22528 ( .A(n26266), .B(n17966), .Z(n17967) );
  AND U22529 ( .A(n26268), .B(n17967), .Z(n17968) );
  OR U22530 ( .A(n17969), .B(n17968), .Z(n17970) );
  NANDN U22531 ( .A(n26273), .B(n17970), .Z(n17971) );
  NANDN U22532 ( .A(n17972), .B(n17971), .Z(n17976) );
  NAND U22533 ( .A(n17974), .B(n17973), .Z(n17975) );
  NANDN U22534 ( .A(n17976), .B(n17975), .Z(n17977) );
  AND U22535 ( .A(n26277), .B(n17977), .Z(n17978) );
  NANDN U22536 ( .A(n17978), .B(n26278), .Z(n17981) );
  NANDN U22537 ( .A(x[2952]), .B(y[2952]), .Z(n17979) );
  NANDN U22538 ( .A(n17980), .B(n17979), .Z(n26280) );
  ANDN U22539 ( .B(n17981), .A(n26280), .Z(n17982) );
  OR U22540 ( .A(n26282), .B(n17982), .Z(n17983) );
  AND U22541 ( .A(n17984), .B(n17983), .Z(n17985) );
  NAND U22542 ( .A(n17985), .B(n26285), .Z(n17987) );
  ANDN U22543 ( .B(n17987), .A(n17986), .Z(n17988) );
  NAND U22544 ( .A(n17988), .B(n26286), .Z(n17989) );
  AND U22545 ( .A(n17990), .B(n17989), .Z(n17992) );
  NAND U22546 ( .A(n17992), .B(n17991), .Z(n17993) );
  NAND U22547 ( .A(n17994), .B(n17993), .Z(n17995) );
  NAND U22548 ( .A(n17995), .B(n26296), .Z(n17997) );
  NANDN U22549 ( .A(n17997), .B(n17996), .Z(n17998) );
  NANDN U22550 ( .A(n26299), .B(n17998), .Z(n17999) );
  NANDN U22551 ( .A(n26301), .B(n17999), .Z(n18000) );
  NAND U22552 ( .A(n18001), .B(n18000), .Z(n18003) );
  NAND U22553 ( .A(n18003), .B(n18002), .Z(n18004) );
  NANDN U22554 ( .A(n18004), .B(n26304), .Z(n18005) );
  NAND U22555 ( .A(n18006), .B(n18005), .Z(n18007) );
  NAND U22556 ( .A(n18008), .B(n18007), .Z(n18010) );
  NAND U22557 ( .A(n18010), .B(n18009), .Z(n18011) );
  NANDN U22558 ( .A(n18011), .B(n26314), .Z(n18012) );
  AND U22559 ( .A(n26316), .B(n18012), .Z(n18015) );
  NOR U22560 ( .A(n18014), .B(n18013), .Z(n26319) );
  NANDN U22561 ( .A(n18015), .B(n26319), .Z(n18017) );
  ANDN U22562 ( .B(n18017), .A(n18016), .Z(n18018) );
  NAND U22563 ( .A(n18018), .B(n26320), .Z(n18019) );
  AND U22564 ( .A(n18020), .B(n18019), .Z(n18021) );
  NAND U22565 ( .A(n18021), .B(n26322), .Z(n18022) );
  AND U22566 ( .A(n18023), .B(n18022), .Z(n18025) );
  NAND U22567 ( .A(n18025), .B(n18024), .Z(n18026) );
  NAND U22568 ( .A(n18027), .B(n18026), .Z(n18028) );
  NAND U22569 ( .A(n18028), .B(n26332), .Z(n18030) );
  NANDN U22570 ( .A(n18030), .B(n18029), .Z(n18031) );
  NANDN U22571 ( .A(n26334), .B(n18031), .Z(n18034) );
  NOR U22572 ( .A(n18033), .B(n18032), .Z(n26336) );
  NAND U22573 ( .A(n18034), .B(n26336), .Z(n18035) );
  NAND U22574 ( .A(n18036), .B(n18035), .Z(n18038) );
  NAND U22575 ( .A(n18038), .B(n18037), .Z(n18039) );
  NANDN U22576 ( .A(n18039), .B(n26341), .Z(n18040) );
  NAND U22577 ( .A(n18041), .B(n18040), .Z(n18042) );
  NAND U22578 ( .A(n18043), .B(n18042), .Z(n18045) );
  NAND U22579 ( .A(n18045), .B(n18044), .Z(n18046) );
  NANDN U22580 ( .A(n18046), .B(n26350), .Z(n18047) );
  AND U22581 ( .A(n26352), .B(n18047), .Z(n18050) );
  NOR U22582 ( .A(n18049), .B(n18048), .Z(n26355) );
  NANDN U22583 ( .A(n18050), .B(n26355), .Z(n18052) );
  ANDN U22584 ( .B(n18052), .A(n18051), .Z(n18053) );
  NAND U22585 ( .A(n18053), .B(n26356), .Z(n18054) );
  AND U22586 ( .A(n18055), .B(n18054), .Z(n18056) );
  NAND U22587 ( .A(n18056), .B(n26358), .Z(n18057) );
  AND U22588 ( .A(n18058), .B(n18057), .Z(n18060) );
  NAND U22589 ( .A(n18060), .B(n18059), .Z(n18061) );
  NAND U22590 ( .A(n18062), .B(n18061), .Z(n18063) );
  NAND U22591 ( .A(n18063), .B(n26368), .Z(n18065) );
  NANDN U22592 ( .A(n18065), .B(n18064), .Z(n18066) );
  NANDN U22593 ( .A(n26370), .B(n18066), .Z(n18069) );
  NOR U22594 ( .A(n18068), .B(n18067), .Z(n26372) );
  NAND U22595 ( .A(n18069), .B(n26372), .Z(n18070) );
  NAND U22596 ( .A(n18071), .B(n18070), .Z(n18073) );
  NAND U22597 ( .A(n18073), .B(n18072), .Z(n18074) );
  NANDN U22598 ( .A(n18074), .B(n26377), .Z(n18075) );
  NAND U22599 ( .A(n18076), .B(n18075), .Z(n18077) );
  NAND U22600 ( .A(n18078), .B(n18077), .Z(n18080) );
  NAND U22601 ( .A(n18080), .B(n18079), .Z(n18081) );
  NANDN U22602 ( .A(n18081), .B(n26386), .Z(n18082) );
  AND U22603 ( .A(n26388), .B(n18082), .Z(n18085) );
  NOR U22604 ( .A(n18084), .B(n18083), .Z(n26391) );
  NANDN U22605 ( .A(n18085), .B(n26391), .Z(n18087) );
  ANDN U22606 ( .B(n18087), .A(n18086), .Z(n18088) );
  NAND U22607 ( .A(n18088), .B(n26392), .Z(n18089) );
  AND U22608 ( .A(n18090), .B(n18089), .Z(n18091) );
  NAND U22609 ( .A(n18091), .B(n26394), .Z(n18092) );
  AND U22610 ( .A(n18093), .B(n18092), .Z(n18095) );
  NAND U22611 ( .A(n18095), .B(n18094), .Z(n18096) );
  NAND U22612 ( .A(n18097), .B(n18096), .Z(n18098) );
  NAND U22613 ( .A(n18098), .B(n26404), .Z(n18100) );
  NANDN U22614 ( .A(n18100), .B(n18099), .Z(n18101) );
  NANDN U22615 ( .A(n26406), .B(n18101), .Z(n18104) );
  NOR U22616 ( .A(n18103), .B(n18102), .Z(n26408) );
  NAND U22617 ( .A(n18104), .B(n26408), .Z(n18105) );
  NAND U22618 ( .A(n18106), .B(n18105), .Z(n18108) );
  NAND U22619 ( .A(n18108), .B(n18107), .Z(n18109) );
  NANDN U22620 ( .A(n18109), .B(n26413), .Z(n18110) );
  NAND U22621 ( .A(n18111), .B(n18110), .Z(n18112) );
  NAND U22622 ( .A(n18113), .B(n18112), .Z(n18115) );
  NAND U22623 ( .A(n18115), .B(n18114), .Z(n18116) );
  NANDN U22624 ( .A(n18116), .B(n26422), .Z(n18117) );
  AND U22625 ( .A(n26424), .B(n18117), .Z(n18120) );
  NOR U22626 ( .A(n18119), .B(n18118), .Z(n26427) );
  NANDN U22627 ( .A(n18120), .B(n26427), .Z(n18122) );
  ANDN U22628 ( .B(n18122), .A(n18121), .Z(n18123) );
  NAND U22629 ( .A(n18123), .B(n26428), .Z(n18124) );
  AND U22630 ( .A(n18125), .B(n18124), .Z(n18126) );
  NAND U22631 ( .A(n18126), .B(n26430), .Z(n18127) );
  AND U22632 ( .A(n18128), .B(n18127), .Z(n18130) );
  NAND U22633 ( .A(n18130), .B(n18129), .Z(n18131) );
  NAND U22634 ( .A(n18132), .B(n18131), .Z(n18133) );
  NAND U22635 ( .A(n18133), .B(n26440), .Z(n18135) );
  NANDN U22636 ( .A(n18135), .B(n18134), .Z(n18136) );
  NANDN U22637 ( .A(n26442), .B(n18136), .Z(n18139) );
  NOR U22638 ( .A(n18138), .B(n18137), .Z(n26444) );
  NAND U22639 ( .A(n18139), .B(n26444), .Z(n18140) );
  NAND U22640 ( .A(n18141), .B(n18140), .Z(n18142) );
  AND U22641 ( .A(n26449), .B(n18142), .Z(n18143) );
  NAND U22642 ( .A(n18144), .B(n18143), .Z(n18146) );
  NAND U22643 ( .A(n18146), .B(n18145), .Z(n18148) );
  ANDN U22644 ( .B(x[3018]), .A(y[3018]), .Z(n18147) );
  OR U22645 ( .A(n18148), .B(n18147), .Z(n18149) );
  NAND U22646 ( .A(n18150), .B(n18149), .Z(n18151) );
  NAND U22647 ( .A(n18152), .B(n18151), .Z(n18153) );
  NANDN U22648 ( .A(n26461), .B(n18153), .Z(n18156) );
  NANDN U22649 ( .A(n18155), .B(n18154), .Z(n26462) );
  ANDN U22650 ( .B(n18156), .A(n26462), .Z(n18157) );
  OR U22651 ( .A(n18158), .B(n18157), .Z(n18159) );
  NAND U22652 ( .A(n18160), .B(n18159), .Z(n18161) );
  NAND U22653 ( .A(n18162), .B(n18161), .Z(n18163) );
  NAND U22654 ( .A(n18163), .B(n26474), .Z(n18165) );
  NANDN U22655 ( .A(n18165), .B(n18164), .Z(n18167) );
  ANDN U22656 ( .B(n18167), .A(n18166), .Z(n18168) );
  NAND U22657 ( .A(n18168), .B(n26476), .Z(n18171) );
  OR U22658 ( .A(n18170), .B(n18169), .Z(n26478) );
  ANDN U22659 ( .B(n18171), .A(n26478), .Z(n18174) );
  NOR U22660 ( .A(n18173), .B(n18172), .Z(n26480) );
  NANDN U22661 ( .A(n18174), .B(n26480), .Z(n18177) );
  ANDN U22662 ( .B(n26482), .A(n18175), .Z(n18176) );
  NAND U22663 ( .A(n18177), .B(n18176), .Z(n18178) );
  NAND U22664 ( .A(n18178), .B(n26485), .Z(n18179) );
  OR U22665 ( .A(n18180), .B(n18179), .Z(n18181) );
  NAND U22666 ( .A(n18182), .B(n18181), .Z(n18183) );
  NAND U22667 ( .A(n18184), .B(n18183), .Z(n18186) );
  NAND U22668 ( .A(n18186), .B(n18185), .Z(n18187) );
  NANDN U22669 ( .A(n18187), .B(n26494), .Z(n18188) );
  AND U22670 ( .A(n26496), .B(n18188), .Z(n18191) );
  NOR U22671 ( .A(n18190), .B(n18189), .Z(n26499) );
  NANDN U22672 ( .A(n18191), .B(n26499), .Z(n18192) );
  AND U22673 ( .A(n26500), .B(n18192), .Z(n18194) );
  NAND U22674 ( .A(n18194), .B(n18193), .Z(n18195) );
  NANDN U22675 ( .A(n26503), .B(n18195), .Z(n18197) );
  NANDN U22676 ( .A(n18197), .B(y[3039]), .Z(n18200) );
  XOR U22677 ( .A(n18197), .B(n18196), .Z(n18198) );
  NANDN U22678 ( .A(x[3039]), .B(n18198), .Z(n18199) );
  AND U22679 ( .A(n18200), .B(n18199), .Z(n18201) );
  NANDN U22680 ( .A(n18201), .B(n18202), .Z(n18205) );
  XNOR U22681 ( .A(n18202), .B(n18201), .Z(n18203) );
  NAND U22682 ( .A(n18203), .B(y[3040]), .Z(n18204) );
  NAND U22683 ( .A(n18205), .B(n18204), .Z(n18206) );
  NAND U22684 ( .A(n18206), .B(n26510), .Z(n18207) );
  NAND U22685 ( .A(n18208), .B(n18207), .Z(n18211) );
  OR U22686 ( .A(n18210), .B(n18209), .Z(n26514) );
  ANDN U22687 ( .B(n18211), .A(n26514), .Z(n18214) );
  NOR U22688 ( .A(n18213), .B(n18212), .Z(n26516) );
  NANDN U22689 ( .A(n18214), .B(n26516), .Z(n18217) );
  ANDN U22690 ( .B(n26518), .A(n18215), .Z(n18216) );
  NAND U22691 ( .A(n18217), .B(n18216), .Z(n18218) );
  NAND U22692 ( .A(n18218), .B(n26521), .Z(n18219) );
  OR U22693 ( .A(n18220), .B(n18219), .Z(n18221) );
  NAND U22694 ( .A(n18222), .B(n18221), .Z(n18223) );
  NAND U22695 ( .A(n18224), .B(n18223), .Z(n18226) );
  NAND U22696 ( .A(n18226), .B(n18225), .Z(n18227) );
  NANDN U22697 ( .A(n18227), .B(n26530), .Z(n18228) );
  AND U22698 ( .A(n26532), .B(n18228), .Z(n18231) );
  NOR U22699 ( .A(n18230), .B(n18229), .Z(n26535) );
  NANDN U22700 ( .A(n18231), .B(n26535), .Z(n18234) );
  ANDN U22701 ( .B(n26536), .A(n18232), .Z(n18233) );
  NAND U22702 ( .A(n18234), .B(n18233), .Z(n18235) );
  NAND U22703 ( .A(n18235), .B(n26543), .Z(n18236) );
  NANDN U22704 ( .A(n18236), .B(n26538), .Z(n18237) );
  AND U22705 ( .A(n18238), .B(n18237), .Z(n18240) );
  NANDN U22706 ( .A(n26545), .B(n26549), .Z(n18239) );
  OR U22707 ( .A(n18240), .B(n18239), .Z(n18242) );
  ANDN U22708 ( .B(n18242), .A(n18241), .Z(n18243) );
  NAND U22709 ( .A(n18243), .B(n26550), .Z(n18246) );
  NANDN U22710 ( .A(n18245), .B(n18244), .Z(n26552) );
  ANDN U22711 ( .B(n18246), .A(n26552), .Z(n18247) );
  OR U22712 ( .A(n26554), .B(n18247), .Z(n18249) );
  ANDN U22713 ( .B(n18249), .A(n18248), .Z(n18250) );
  NAND U22714 ( .A(n18250), .B(n26557), .Z(n18252) );
  ANDN U22715 ( .B(n18252), .A(n18251), .Z(n18253) );
  NAND U22716 ( .A(n18253), .B(n26558), .Z(n18255) );
  ANDN U22717 ( .B(x[3060]), .A(y[3060]), .Z(n18254) );
  ANDN U22718 ( .B(n18255), .A(n18254), .Z(n18257) );
  NAND U22719 ( .A(n18257), .B(n18256), .Z(n18258) );
  NAND U22720 ( .A(n18259), .B(n18258), .Z(n18260) );
  NAND U22721 ( .A(n18260), .B(n26568), .Z(n18262) );
  NANDN U22722 ( .A(n18262), .B(n18261), .Z(n18263) );
  NANDN U22723 ( .A(n26571), .B(n18263), .Z(n18264) );
  NANDN U22724 ( .A(n26573), .B(n18264), .Z(n18265) );
  NAND U22725 ( .A(n18266), .B(n18265), .Z(n18267) );
  NAND U22726 ( .A(n18267), .B(n26580), .Z(n18268) );
  NANDN U22727 ( .A(n18268), .B(n26576), .Z(n18269) );
  AND U22728 ( .A(n18270), .B(n18269), .Z(n18271) );
  OR U22729 ( .A(n18272), .B(n18271), .Z(n18273) );
  NANDN U22730 ( .A(n26588), .B(n18273), .Z(n18276) );
  NANDN U22731 ( .A(y[3070]), .B(x[3070]), .Z(n18275) );
  ANDN U22732 ( .B(n18275), .A(n18274), .Z(n26590) );
  NAND U22733 ( .A(n18276), .B(n26590), .Z(n18277) );
  NANDN U22734 ( .A(n26593), .B(n18277), .Z(n18280) );
  NANDN U22735 ( .A(y[3072]), .B(x[3072]), .Z(n18278) );
  NAND U22736 ( .A(n18279), .B(n18278), .Z(n26594) );
  ANDN U22737 ( .B(n18280), .A(n26594), .Z(n18281) );
  OR U22738 ( .A(n26597), .B(n18281), .Z(n18282) );
  NANDN U22739 ( .A(n26599), .B(n18282), .Z(n18283) );
  NANDN U22740 ( .A(n26601), .B(n18283), .Z(n18284) );
  AND U22741 ( .A(n26602), .B(n18284), .Z(n18288) );
  NAND U22742 ( .A(n18285), .B(y[3078]), .Z(n18287) );
  NAND U22743 ( .A(n18287), .B(n18286), .Z(n26604) );
  OR U22744 ( .A(n18288), .B(n26604), .Z(n18291) );
  NANDN U22745 ( .A(y[3078]), .B(x[3078]), .Z(n18290) );
  ANDN U22746 ( .B(n18290), .A(n18289), .Z(n26606) );
  NAND U22747 ( .A(n18291), .B(n26606), .Z(n18295) );
  NAND U22748 ( .A(n18292), .B(y[3080]), .Z(n18293) );
  NANDN U22749 ( .A(n18294), .B(n18293), .Z(n26609) );
  ANDN U22750 ( .B(n18295), .A(n26609), .Z(n18296) );
  OR U22751 ( .A(n26611), .B(n18296), .Z(n18299) );
  NANDN U22752 ( .A(x[3082]), .B(y[3082]), .Z(n18298) );
  AND U22753 ( .A(n18298), .B(n18297), .Z(n26612) );
  NAND U22754 ( .A(n18299), .B(n26612), .Z(n18300) );
  NANDN U22755 ( .A(n26614), .B(n18300), .Z(n18301) );
  NANDN U22756 ( .A(n26617), .B(n18301), .Z(n18304) );
  NANDN U22757 ( .A(y[3084]), .B(x[3084]), .Z(n18302) );
  NAND U22758 ( .A(n18303), .B(n18302), .Z(n26619) );
  ANDN U22759 ( .B(n18304), .A(n26619), .Z(n18305) );
  OR U22760 ( .A(n26621), .B(n18305), .Z(n18308) );
  NANDN U22761 ( .A(y[3087]), .B(x[3087]), .Z(n18307) );
  NANDN U22762 ( .A(y[3086]), .B(x[3086]), .Z(n18306) );
  AND U22763 ( .A(n18307), .B(n18306), .Z(n26622) );
  NAND U22764 ( .A(n18308), .B(n26622), .Z(n18309) );
  NANDN U22765 ( .A(n26624), .B(n18309), .Z(n18310) );
  NANDN U22766 ( .A(n26627), .B(n18310), .Z(n18313) );
  NANDN U22767 ( .A(x[3089]), .B(y[3089]), .Z(n18311) );
  NANDN U22768 ( .A(n18312), .B(n18311), .Z(n26629) );
  ANDN U22769 ( .B(n18313), .A(n26629), .Z(n18316) );
  NOR U22770 ( .A(n18315), .B(n18314), .Z(n26630) );
  NANDN U22771 ( .A(n18316), .B(n26630), .Z(n18317) );
  NAND U22772 ( .A(n18318), .B(n18317), .Z(n18319) );
  NANDN U22773 ( .A(n18319), .B(n26634), .Z(n18320) );
  AND U22774 ( .A(n26636), .B(n18320), .Z(n18321) );
  ANDN U22775 ( .B(n26640), .A(n18321), .Z(n18323) );
  XNOR U22776 ( .A(x[3094]), .B(y[3094]), .Z(n18322) );
  AND U22777 ( .A(n18323), .B(n18322), .Z(n18324) );
  OR U22778 ( .A(n26643), .B(n18324), .Z(n18325) );
  NANDN U22779 ( .A(n26644), .B(n18325), .Z(n18328) );
  NANDN U22780 ( .A(y[3096]), .B(x[3096]), .Z(n18327) );
  ANDN U22781 ( .B(n18327), .A(n18326), .Z(n26646) );
  NAND U22782 ( .A(n18328), .B(n26646), .Z(n18329) );
  NANDN U22783 ( .A(n26649), .B(n18329), .Z(n18330) );
  AND U22784 ( .A(n26650), .B(n18330), .Z(n18331) );
  OR U22785 ( .A(n26653), .B(n18331), .Z(n18332) );
  NANDN U22786 ( .A(n26654), .B(n18332), .Z(n18335) );
  NANDN U22787 ( .A(x[3101]), .B(y[3101]), .Z(n18334) );
  ANDN U22788 ( .B(n18334), .A(n18333), .Z(n26656) );
  NAND U22789 ( .A(n18335), .B(n26656), .Z(n18336) );
  NANDN U22790 ( .A(n26659), .B(n18336), .Z(n18337) );
  AND U22791 ( .A(n26660), .B(n18337), .Z(n18338) );
  OR U22792 ( .A(n26663), .B(n18338), .Z(n18339) );
  NANDN U22793 ( .A(n26664), .B(n18339), .Z(n18340) );
  NANDN U22794 ( .A(n26667), .B(n18340), .Z(n18341) );
  NANDN U22795 ( .A(n26669), .B(n18341), .Z(n18342) );
  AND U22796 ( .A(n26670), .B(n18342), .Z(n18345) );
  NANDN U22797 ( .A(x[3109]), .B(y[3109]), .Z(n18344) );
  ANDN U22798 ( .B(n18344), .A(n18343), .Z(n26672) );
  NANDN U22799 ( .A(n18345), .B(n26672), .Z(n18346) );
  NANDN U22800 ( .A(n26674), .B(n18346), .Z(n18347) );
  NANDN U22801 ( .A(n26677), .B(n18347), .Z(n18348) );
  NANDN U22802 ( .A(n26679), .B(n18348), .Z(n18349) );
  AND U22803 ( .A(n26680), .B(n18349), .Z(n18350) );
  OR U22804 ( .A(n26683), .B(n18350), .Z(n18351) );
  NANDN U22805 ( .A(n26684), .B(n18351), .Z(n18352) );
  NANDN U22806 ( .A(n26687), .B(n18352), .Z(n18355) );
  NANDN U22807 ( .A(x[3117]), .B(y[3117]), .Z(n18354) );
  ANDN U22808 ( .B(n18354), .A(n18353), .Z(n26688) );
  NAND U22809 ( .A(n18355), .B(n26688), .Z(n18356) );
  AND U22810 ( .A(n26690), .B(n18356), .Z(n18357) );
  OR U22811 ( .A(n26693), .B(n18357), .Z(n18358) );
  NANDN U22812 ( .A(n26694), .B(n18358), .Z(n18361) );
  NANDN U22813 ( .A(x[3121]), .B(y[3121]), .Z(n18360) );
  ANDN U22814 ( .B(n18360), .A(n18359), .Z(n26696) );
  NAND U22815 ( .A(n18361), .B(n26696), .Z(n18362) );
  NANDN U22816 ( .A(n26699), .B(n18362), .Z(n18363) );
  AND U22817 ( .A(n26700), .B(n18363), .Z(n18364) );
  OR U22818 ( .A(n26703), .B(n18364), .Z(n18365) );
  NANDN U22819 ( .A(n26704), .B(n18365), .Z(n18366) );
  NANDN U22820 ( .A(n26707), .B(n18366), .Z(n18367) );
  NANDN U22821 ( .A(n26709), .B(n18367), .Z(n18368) );
  AND U22822 ( .A(n26710), .B(n18368), .Z(n18369) );
  OR U22823 ( .A(n18369), .B(n26713), .Z(n18370) );
  AND U22824 ( .A(n26714), .B(n18370), .Z(n18371) );
  OR U22825 ( .A(n18371), .B(n26716), .Z(n18372) );
  AND U22826 ( .A(n26718), .B(n18372), .Z(n18373) );
  OR U22827 ( .A(n18373), .B(n26720), .Z(n18374) );
  AND U22828 ( .A(n26722), .B(n18374), .Z(n18375) );
  OR U22829 ( .A(n18375), .B(n26724), .Z(n18376) );
  AND U22830 ( .A(n26726), .B(n18376), .Z(n18377) );
  OR U22831 ( .A(n26728), .B(n18377), .Z(n18380) );
  AND U22832 ( .A(n18379), .B(n18378), .Z(n26730) );
  NAND U22833 ( .A(n18380), .B(n26730), .Z(n18383) );
  NANDN U22834 ( .A(x[3139]), .B(y[3139]), .Z(n18382) );
  ANDN U22835 ( .B(n18382), .A(n18381), .Z(n26732) );
  NAND U22836 ( .A(n18383), .B(n26732), .Z(n18384) );
  NANDN U22837 ( .A(n26735), .B(n18384), .Z(n18385) );
  AND U22838 ( .A(n26736), .B(n18385), .Z(n18386) );
  OR U22839 ( .A(n26738), .B(n18386), .Z(n18389) );
  NANDN U22840 ( .A(x[3143]), .B(y[3143]), .Z(n18388) );
  NANDN U22841 ( .A(x[3144]), .B(y[3144]), .Z(n18387) );
  AND U22842 ( .A(n18388), .B(n18387), .Z(n26740) );
  NAND U22843 ( .A(n18389), .B(n26740), .Z(n18390) );
  NANDN U22844 ( .A(n26743), .B(n18390), .Z(n18393) );
  NANDN U22845 ( .A(x[3145]), .B(y[3145]), .Z(n18392) );
  ANDN U22846 ( .B(n18392), .A(n18391), .Z(n26744) );
  NAND U22847 ( .A(n18393), .B(n26744), .Z(n18394) );
  NAND U22848 ( .A(n18394), .B(n26746), .Z(n18395) );
  ANDN U22849 ( .B(n18395), .A(n26749), .Z(n18396) );
  NANDN U22850 ( .A(n18396), .B(n26750), .Z(n18399) );
  OR U22851 ( .A(n18398), .B(n18397), .Z(n26752) );
  ANDN U22852 ( .B(n18399), .A(n26752), .Z(n18402) );
  NOR U22853 ( .A(n18401), .B(n18400), .Z(n26754) );
  NANDN U22854 ( .A(n18402), .B(n26754), .Z(n18403) );
  NAND U22855 ( .A(n18404), .B(n18403), .Z(n18405) );
  NANDN U22856 ( .A(n18405), .B(n20233), .Z(n18406) );
  AND U22857 ( .A(n26758), .B(n18406), .Z(n18409) );
  NANDN U22858 ( .A(x[3153]), .B(y[3153]), .Z(n18408) );
  ANDN U22859 ( .B(n18408), .A(n18407), .Z(n26760) );
  NANDN U22860 ( .A(n18409), .B(n26760), .Z(n18412) );
  NANDN U22861 ( .A(y[3155]), .B(x[3155]), .Z(n18411) );
  ANDN U22862 ( .B(n18411), .A(n18410), .Z(n26762) );
  NAND U22863 ( .A(n18412), .B(n26762), .Z(n18413) );
  NANDN U22864 ( .A(n26765), .B(n18413), .Z(n18414) );
  NANDN U22865 ( .A(n26766), .B(n18414), .Z(n18415) );
  AND U22866 ( .A(n26768), .B(n18415), .Z(n18418) );
  NANDN U22867 ( .A(y[3158]), .B(x[3158]), .Z(n18417) );
  ANDN U22868 ( .B(n18417), .A(n18416), .Z(n26770) );
  NANDN U22869 ( .A(n18418), .B(n26770), .Z(n18421) );
  NOR U22870 ( .A(n18420), .B(n18419), .Z(n26772) );
  NAND U22871 ( .A(n18421), .B(n26772), .Z(n18422) );
  NANDN U22872 ( .A(n26775), .B(n18422), .Z(n18423) );
  NANDN U22873 ( .A(n26776), .B(n18423), .Z(n18424) );
  AND U22874 ( .A(n26778), .B(n18424), .Z(n18425) );
  OR U22875 ( .A(n26781), .B(n18425), .Z(n18428) );
  NANDN U22876 ( .A(y[3165]), .B(x[3165]), .Z(n18427) );
  ANDN U22877 ( .B(n18427), .A(n18426), .Z(n26782) );
  NAND U22878 ( .A(n18428), .B(n26782), .Z(n18429) );
  NANDN U22879 ( .A(n26785), .B(n18429), .Z(n18432) );
  NANDN U22880 ( .A(y[3166]), .B(x[3166]), .Z(n18431) );
  ANDN U22881 ( .B(n18431), .A(n18430), .Z(n26787) );
  NAND U22882 ( .A(n18432), .B(n26787), .Z(n18433) );
  AND U22883 ( .A(n26788), .B(n18433), .Z(n18434) );
  OR U22884 ( .A(n26791), .B(n18434), .Z(n18437) );
  AND U22885 ( .A(n18436), .B(n18435), .Z(n26792) );
  NAND U22886 ( .A(n18437), .B(n26792), .Z(n18440) );
  NANDN U22887 ( .A(y[3170]), .B(x[3170]), .Z(n18439) );
  ANDN U22888 ( .B(n18439), .A(n18438), .Z(n26794) );
  NAND U22889 ( .A(n18440), .B(n26794), .Z(n18441) );
  NANDN U22890 ( .A(n26796), .B(n18441), .Z(n18442) );
  AND U22891 ( .A(n26798), .B(n18442), .Z(n18445) );
  AND U22892 ( .A(n18443), .B(n26801), .Z(n18444) );
  NANDN U22893 ( .A(n18445), .B(n18444), .Z(n18446) );
  NANDN U22894 ( .A(n26805), .B(n18446), .Z(n18449) );
  NANDN U22895 ( .A(x[3175]), .B(y[3175]), .Z(n18447) );
  NAND U22896 ( .A(n18448), .B(n18447), .Z(n26807) );
  ANDN U22897 ( .B(n18449), .A(n26807), .Z(n18450) );
  OR U22898 ( .A(n26809), .B(n18450), .Z(n18453) );
  NANDN U22899 ( .A(x[3178]), .B(y[3178]), .Z(n18452) );
  ANDN U22900 ( .B(n18452), .A(n18451), .Z(n26810) );
  NAND U22901 ( .A(n18453), .B(n26810), .Z(n18454) );
  NANDN U22902 ( .A(n26813), .B(n18454), .Z(n18457) );
  NANDN U22903 ( .A(x[3179]), .B(y[3179]), .Z(n18456) );
  ANDN U22904 ( .B(n18456), .A(n18455), .Z(n26815) );
  NAND U22905 ( .A(n18457), .B(n26815), .Z(n18458) );
  AND U22906 ( .A(n26816), .B(n18458), .Z(n18459) );
  OR U22907 ( .A(n26819), .B(n18459), .Z(n18462) );
  AND U22908 ( .A(n18461), .B(n18460), .Z(n26820) );
  NAND U22909 ( .A(n18462), .B(n26820), .Z(n18465) );
  NANDN U22910 ( .A(x[3183]), .B(y[3183]), .Z(n18464) );
  ANDN U22911 ( .B(n18464), .A(n18463), .Z(n26822) );
  NAND U22912 ( .A(n18465), .B(n26822), .Z(n18466) );
  NANDN U22913 ( .A(n26824), .B(n18466), .Z(n18467) );
  AND U22914 ( .A(n26826), .B(n18467), .Z(n18468) );
  OR U22915 ( .A(n26829), .B(n18468), .Z(n18471) );
  NANDN U22916 ( .A(x[3187]), .B(y[3187]), .Z(n18470) );
  ANDN U22917 ( .B(n18470), .A(n18469), .Z(n26830) );
  NAND U22918 ( .A(n18471), .B(n26830), .Z(n18472) );
  NANDN U22919 ( .A(n26833), .B(n18472), .Z(n18473) );
  NANDN U22920 ( .A(n26834), .B(n18473), .Z(n18474) );
  AND U22921 ( .A(n26836), .B(n18474), .Z(n18477) );
  NANDN U22922 ( .A(x[3191]), .B(y[3191]), .Z(n18476) );
  ANDN U22923 ( .B(n18476), .A(n18475), .Z(n26838) );
  NANDN U22924 ( .A(n18477), .B(n26838), .Z(n18480) );
  NOR U22925 ( .A(n18479), .B(n18478), .Z(n26840) );
  NAND U22926 ( .A(n18480), .B(n26840), .Z(n18481) );
  NANDN U22927 ( .A(n26843), .B(n18481), .Z(n18482) );
  NANDN U22928 ( .A(n26844), .B(n18482), .Z(n18483) );
  AND U22929 ( .A(n26846), .B(n18483), .Z(n18484) );
  OR U22930 ( .A(n26849), .B(n18484), .Z(n18487) );
  NANDN U22931 ( .A(x[3198]), .B(y[3198]), .Z(n18486) );
  ANDN U22932 ( .B(n18486), .A(n18485), .Z(n26850) );
  NAND U22933 ( .A(n18487), .B(n26850), .Z(n18488) );
  NANDN U22934 ( .A(n26853), .B(n18488), .Z(n18491) );
  NANDN U22935 ( .A(x[3199]), .B(y[3199]), .Z(n18490) );
  ANDN U22936 ( .B(n18490), .A(n18489), .Z(n26855) );
  NAND U22937 ( .A(n18491), .B(n26855), .Z(n18492) );
  AND U22938 ( .A(n26856), .B(n18492), .Z(n18493) );
  OR U22939 ( .A(n26859), .B(n18493), .Z(n18496) );
  AND U22940 ( .A(n18495), .B(n18494), .Z(n26860) );
  NAND U22941 ( .A(n18496), .B(n26860), .Z(n18499) );
  NANDN U22942 ( .A(x[3203]), .B(y[3203]), .Z(n18498) );
  ANDN U22943 ( .B(n18498), .A(n18497), .Z(n26862) );
  NAND U22944 ( .A(n18499), .B(n26862), .Z(n18500) );
  NANDN U22945 ( .A(n26864), .B(n18500), .Z(n18501) );
  AND U22946 ( .A(n26866), .B(n18501), .Z(n18502) );
  OR U22947 ( .A(n26869), .B(n18502), .Z(n18505) );
  NANDN U22948 ( .A(x[3207]), .B(y[3207]), .Z(n18504) );
  ANDN U22949 ( .B(n18504), .A(n18503), .Z(n26870) );
  NAND U22950 ( .A(n18505), .B(n26870), .Z(n18506) );
  NANDN U22951 ( .A(n26873), .B(n18506), .Z(n18507) );
  NANDN U22952 ( .A(n26874), .B(n18507), .Z(n18508) );
  AND U22953 ( .A(n26876), .B(n18508), .Z(n18511) );
  NANDN U22954 ( .A(x[3211]), .B(y[3211]), .Z(n18510) );
  ANDN U22955 ( .B(n18510), .A(n18509), .Z(n26878) );
  NANDN U22956 ( .A(n18511), .B(n26878), .Z(n18514) );
  NOR U22957 ( .A(n18513), .B(n18512), .Z(n26880) );
  NAND U22958 ( .A(n18514), .B(n26880), .Z(n18515) );
  NANDN U22959 ( .A(n26883), .B(n18515), .Z(n18516) );
  NANDN U22960 ( .A(n26884), .B(n18516), .Z(n18517) );
  AND U22961 ( .A(n26886), .B(n18517), .Z(n18518) );
  OR U22962 ( .A(n26889), .B(n18518), .Z(n18521) );
  NANDN U22963 ( .A(x[3218]), .B(y[3218]), .Z(n18520) );
  ANDN U22964 ( .B(n18520), .A(n18519), .Z(n26890) );
  NAND U22965 ( .A(n18521), .B(n26890), .Z(n18522) );
  NANDN U22966 ( .A(n26893), .B(n18522), .Z(n18525) );
  NANDN U22967 ( .A(x[3219]), .B(y[3219]), .Z(n18524) );
  ANDN U22968 ( .B(n18524), .A(n18523), .Z(n26895) );
  NAND U22969 ( .A(n18525), .B(n26895), .Z(n18526) );
  AND U22970 ( .A(n26896), .B(n18526), .Z(n18527) );
  OR U22971 ( .A(n26899), .B(n18527), .Z(n18530) );
  AND U22972 ( .A(n18529), .B(n18528), .Z(n26900) );
  NAND U22973 ( .A(n18530), .B(n26900), .Z(n18533) );
  NANDN U22974 ( .A(x[3223]), .B(y[3223]), .Z(n18532) );
  ANDN U22975 ( .B(n18532), .A(n18531), .Z(n26902) );
  NAND U22976 ( .A(n18533), .B(n26902), .Z(n18534) );
  NANDN U22977 ( .A(n26904), .B(n18534), .Z(n18535) );
  AND U22978 ( .A(n26906), .B(n18535), .Z(n18536) );
  OR U22979 ( .A(n26909), .B(n18536), .Z(n18539) );
  NANDN U22980 ( .A(x[3227]), .B(y[3227]), .Z(n18538) );
  ANDN U22981 ( .B(n18538), .A(n18537), .Z(n26910) );
  NAND U22982 ( .A(n18539), .B(n26910), .Z(n18540) );
  NANDN U22983 ( .A(n26913), .B(n18540), .Z(n18541) );
  NANDN U22984 ( .A(n26914), .B(n18541), .Z(n18542) );
  AND U22985 ( .A(n26916), .B(n18542), .Z(n18545) );
  NANDN U22986 ( .A(x[3231]), .B(y[3231]), .Z(n18544) );
  ANDN U22987 ( .B(n18544), .A(n18543), .Z(n26918) );
  NANDN U22988 ( .A(n18545), .B(n26918), .Z(n18548) );
  NOR U22989 ( .A(n18547), .B(n18546), .Z(n26920) );
  NAND U22990 ( .A(n18548), .B(n26920), .Z(n18549) );
  NANDN U22991 ( .A(n26923), .B(n18549), .Z(n18550) );
  NANDN U22992 ( .A(n26924), .B(n18550), .Z(n18551) );
  AND U22993 ( .A(n26926), .B(n18551), .Z(n18552) );
  OR U22994 ( .A(n26929), .B(n18552), .Z(n18555) );
  NANDN U22995 ( .A(x[3238]), .B(y[3238]), .Z(n18554) );
  ANDN U22996 ( .B(n18554), .A(n18553), .Z(n26930) );
  NAND U22997 ( .A(n18555), .B(n26930), .Z(n18556) );
  NANDN U22998 ( .A(n26933), .B(n18556), .Z(n18559) );
  NANDN U22999 ( .A(x[3239]), .B(y[3239]), .Z(n18558) );
  ANDN U23000 ( .B(n18558), .A(n18557), .Z(n26935) );
  NAND U23001 ( .A(n18559), .B(n26935), .Z(n18560) );
  AND U23002 ( .A(n26936), .B(n18560), .Z(n18561) );
  OR U23003 ( .A(n26939), .B(n18561), .Z(n18564) );
  AND U23004 ( .A(n18563), .B(n18562), .Z(n26940) );
  NAND U23005 ( .A(n18564), .B(n26940), .Z(n18567) );
  NANDN U23006 ( .A(x[3243]), .B(y[3243]), .Z(n18566) );
  ANDN U23007 ( .B(n18566), .A(n18565), .Z(n26942) );
  NAND U23008 ( .A(n18567), .B(n26942), .Z(n18568) );
  NANDN U23009 ( .A(n26944), .B(n18568), .Z(n18569) );
  AND U23010 ( .A(n26946), .B(n18569), .Z(n18570) );
  OR U23011 ( .A(n26949), .B(n18570), .Z(n18573) );
  NANDN U23012 ( .A(x[3247]), .B(y[3247]), .Z(n18572) );
  ANDN U23013 ( .B(n18572), .A(n18571), .Z(n26950) );
  NAND U23014 ( .A(n18573), .B(n26950), .Z(n18574) );
  NANDN U23015 ( .A(n26953), .B(n18574), .Z(n18575) );
  NANDN U23016 ( .A(n26954), .B(n18575), .Z(n18576) );
  AND U23017 ( .A(n26956), .B(n18576), .Z(n18579) );
  NANDN U23018 ( .A(x[3251]), .B(y[3251]), .Z(n18578) );
  ANDN U23019 ( .B(n18578), .A(n18577), .Z(n26958) );
  NANDN U23020 ( .A(n18579), .B(n26958), .Z(n18582) );
  NOR U23021 ( .A(n18581), .B(n18580), .Z(n26960) );
  NAND U23022 ( .A(n18582), .B(n26960), .Z(n18583) );
  NANDN U23023 ( .A(n26963), .B(n18583), .Z(n18584) );
  NANDN U23024 ( .A(n26964), .B(n18584), .Z(n18585) );
  AND U23025 ( .A(n26966), .B(n18585), .Z(n18586) );
  OR U23026 ( .A(n26969), .B(n18586), .Z(n18589) );
  NANDN U23027 ( .A(x[3258]), .B(y[3258]), .Z(n18588) );
  ANDN U23028 ( .B(n18588), .A(n18587), .Z(n26970) );
  NAND U23029 ( .A(n18589), .B(n26970), .Z(n18590) );
  NANDN U23030 ( .A(n26972), .B(n18590), .Z(n18591) );
  AND U23031 ( .A(n26974), .B(n18591), .Z(n18592) );
  OR U23032 ( .A(n26977), .B(n18592), .Z(n18593) );
  NAND U23033 ( .A(n18593), .B(n26978), .Z(n18594) );
  NANDN U23034 ( .A(n26981), .B(n18594), .Z(n18597) );
  NANDN U23035 ( .A(n18596), .B(n18595), .Z(n26982) );
  ANDN U23036 ( .B(n18597), .A(n26982), .Z(n18598) );
  NANDN U23037 ( .A(n18598), .B(n26984), .Z(n18599) );
  NAND U23038 ( .A(n18599), .B(n26987), .Z(n18600) );
  NAND U23039 ( .A(n18600), .B(n26988), .Z(n18601) );
  NAND U23040 ( .A(n18601), .B(n26991), .Z(n18604) );
  NOR U23041 ( .A(n18603), .B(n18602), .Z(n26992) );
  NAND U23042 ( .A(n18604), .B(n26992), .Z(n18605) );
  NAND U23043 ( .A(n18605), .B(n20231), .Z(n18607) );
  NANDN U23044 ( .A(n18607), .B(n18606), .Z(n18608) );
  AND U23045 ( .A(n26996), .B(n18608), .Z(n18611) );
  NANDN U23046 ( .A(x[3271]), .B(y[3271]), .Z(n18610) );
  ANDN U23047 ( .B(n18610), .A(n18609), .Z(n26998) );
  NANDN U23048 ( .A(n18611), .B(n26998), .Z(n18614) );
  NANDN U23049 ( .A(y[3273]), .B(x[3273]), .Z(n18613) );
  ANDN U23050 ( .B(n18613), .A(n18612), .Z(n27000) );
  NAND U23051 ( .A(n18614), .B(n27000), .Z(n18615) );
  NANDN U23052 ( .A(n27003), .B(n18615), .Z(n18618) );
  NANDN U23053 ( .A(y[3274]), .B(x[3274]), .Z(n18617) );
  ANDN U23054 ( .B(n18617), .A(n18616), .Z(n27005) );
  NAND U23055 ( .A(n18618), .B(n27005), .Z(n18619) );
  AND U23056 ( .A(n27006), .B(n18619), .Z(n18620) );
  OR U23057 ( .A(n27009), .B(n18620), .Z(n18623) );
  AND U23058 ( .A(n18622), .B(n18621), .Z(n27010) );
  NAND U23059 ( .A(n18623), .B(n27010), .Z(n18626) );
  NANDN U23060 ( .A(y[3278]), .B(x[3278]), .Z(n18625) );
  ANDN U23061 ( .B(n18625), .A(n18624), .Z(n27012) );
  NAND U23062 ( .A(n18626), .B(n27012), .Z(n18627) );
  NANDN U23063 ( .A(n27014), .B(n18627), .Z(n18628) );
  AND U23064 ( .A(n27016), .B(n18628), .Z(n18629) );
  OR U23065 ( .A(n27019), .B(n18629), .Z(n18632) );
  NANDN U23066 ( .A(y[3283]), .B(x[3283]), .Z(n18631) );
  NANDN U23067 ( .A(y[3282]), .B(x[3282]), .Z(n18630) );
  AND U23068 ( .A(n18631), .B(n18630), .Z(n27020) );
  NAND U23069 ( .A(n18632), .B(n27020), .Z(n18633) );
  NANDN U23070 ( .A(n27023), .B(n18633), .Z(n18636) );
  NANDN U23071 ( .A(y[3284]), .B(x[3284]), .Z(n18635) );
  ANDN U23072 ( .B(n18635), .A(n18634), .Z(n27025) );
  NAND U23073 ( .A(n18636), .B(n27025), .Z(n18637) );
  AND U23074 ( .A(n27026), .B(n18637), .Z(n18638) );
  OR U23075 ( .A(n27029), .B(n18638), .Z(n18641) );
  NANDN U23076 ( .A(x[3288]), .B(y[3288]), .Z(n18640) );
  AND U23077 ( .A(n18640), .B(n18639), .Z(n27030) );
  NAND U23078 ( .A(n18641), .B(n27030), .Z(n18642) );
  NANDN U23079 ( .A(n27033), .B(n18642), .Z(n18643) );
  NANDN U23080 ( .A(n27034), .B(n18643), .Z(n18644) );
  AND U23081 ( .A(n27036), .B(n18644), .Z(n18645) );
  OR U23082 ( .A(n27039), .B(n18645), .Z(n18648) );
  NANDN U23083 ( .A(y[3293]), .B(x[3293]), .Z(n18647) );
  NANDN U23084 ( .A(y[3292]), .B(x[3292]), .Z(n18646) );
  AND U23085 ( .A(n18647), .B(n18646), .Z(n27040) );
  NAND U23086 ( .A(n18648), .B(n27040), .Z(n18649) );
  NANDN U23087 ( .A(n27043), .B(n18649), .Z(n18650) );
  NANDN U23088 ( .A(n27044), .B(n18650), .Z(n18651) );
  AND U23089 ( .A(n27046), .B(n18651), .Z(n18654) );
  NANDN U23090 ( .A(y[3296]), .B(x[3296]), .Z(n18653) );
  ANDN U23091 ( .B(n18653), .A(n18652), .Z(n27048) );
  NANDN U23092 ( .A(n18654), .B(n27048), .Z(n18657) );
  NANDN U23093 ( .A(x[3298]), .B(y[3298]), .Z(n18656) );
  ANDN U23094 ( .B(n18656), .A(n18655), .Z(n27050) );
  NAND U23095 ( .A(n18657), .B(n27050), .Z(n18658) );
  NANDN U23096 ( .A(n27053), .B(n18658), .Z(n18659) );
  NANDN U23097 ( .A(n27054), .B(n18659), .Z(n18660) );
  AND U23098 ( .A(n27056), .B(n18660), .Z(n18661) );
  OR U23099 ( .A(n27059), .B(n18661), .Z(n18664) );
  NANDN U23100 ( .A(y[3302]), .B(x[3302]), .Z(n18663) );
  ANDN U23101 ( .B(n18663), .A(n18662), .Z(n27060) );
  NAND U23102 ( .A(n18664), .B(n27060), .Z(n18665) );
  NANDN U23103 ( .A(n27063), .B(n18665), .Z(n18666) );
  NANDN U23104 ( .A(n27064), .B(n18666), .Z(n18667) );
  AND U23105 ( .A(n27066), .B(n18667), .Z(n18668) );
  OR U23106 ( .A(n27069), .B(n18668), .Z(n18671) );
  AND U23107 ( .A(n18670), .B(n18669), .Z(n27070) );
  NAND U23108 ( .A(n18671), .B(n27070), .Z(n18674) );
  NANDN U23109 ( .A(y[3308]), .B(x[3308]), .Z(n18673) );
  ANDN U23110 ( .B(n18673), .A(n18672), .Z(n27072) );
  NAND U23111 ( .A(n18674), .B(n27072), .Z(n18675) );
  NANDN U23112 ( .A(n27074), .B(n18675), .Z(n18676) );
  AND U23113 ( .A(n27076), .B(n18676), .Z(n18677) );
  OR U23114 ( .A(n27079), .B(n18677), .Z(n18680) );
  NANDN U23115 ( .A(y[3313]), .B(x[3313]), .Z(n18679) );
  NANDN U23116 ( .A(y[3312]), .B(x[3312]), .Z(n18678) );
  AND U23117 ( .A(n18679), .B(n18678), .Z(n27080) );
  NAND U23118 ( .A(n18680), .B(n27080), .Z(n18681) );
  NANDN U23119 ( .A(n27083), .B(n18681), .Z(n18684) );
  NANDN U23120 ( .A(y[3314]), .B(x[3314]), .Z(n18683) );
  ANDN U23121 ( .B(n18683), .A(n18682), .Z(n27085) );
  NAND U23122 ( .A(n18684), .B(n27085), .Z(n18685) );
  AND U23123 ( .A(n27086), .B(n18685), .Z(n18686) );
  OR U23124 ( .A(n27089), .B(n18686), .Z(n18689) );
  NANDN U23125 ( .A(x[3318]), .B(y[3318]), .Z(n18687) );
  AND U23126 ( .A(n18688), .B(n18687), .Z(n27090) );
  NAND U23127 ( .A(n18689), .B(n27090), .Z(n18690) );
  NANDN U23128 ( .A(n27093), .B(n18690), .Z(n18691) );
  NAND U23129 ( .A(n18692), .B(n18691), .Z(n18693) );
  NANDN U23130 ( .A(n27097), .B(n18693), .Z(n18696) );
  NANDN U23131 ( .A(n18695), .B(n18694), .Z(n27099) );
  ANDN U23132 ( .B(n18696), .A(n27099), .Z(n18699) );
  NANDN U23133 ( .A(y[3322]), .B(x[3322]), .Z(n18698) );
  ANDN U23134 ( .B(n18698), .A(n18697), .Z(n27100) );
  NANDN U23135 ( .A(n18699), .B(n27100), .Z(n18702) );
  NOR U23136 ( .A(n18701), .B(n18700), .Z(n27102) );
  NAND U23137 ( .A(n18702), .B(n27102), .Z(n18703) );
  NANDN U23138 ( .A(n27104), .B(n18703), .Z(n18704) );
  NAND U23139 ( .A(n18705), .B(n18704), .Z(n18706) );
  AND U23140 ( .A(n27110), .B(n18706), .Z(n18709) );
  NANDN U23141 ( .A(x[3327]), .B(y[3327]), .Z(n18708) );
  ANDN U23142 ( .B(n18708), .A(n18707), .Z(n27113) );
  NANDN U23143 ( .A(n18709), .B(n27113), .Z(n18712) );
  NOR U23144 ( .A(n18711), .B(n18710), .Z(n27114) );
  NAND U23145 ( .A(n18712), .B(n27114), .Z(n18713) );
  NANDN U23146 ( .A(n27117), .B(n18713), .Z(n18714) );
  AND U23147 ( .A(n27118), .B(n18714), .Z(n18715) );
  OR U23148 ( .A(n27121), .B(n18715), .Z(n18716) );
  NANDN U23149 ( .A(n27122), .B(n18716), .Z(n18717) );
  NAND U23150 ( .A(n18717), .B(n27124), .Z(n18718) );
  ANDN U23151 ( .B(n18718), .A(n27126), .Z(n18719) );
  NANDN U23152 ( .A(n18719), .B(n27128), .Z(n18720) );
  NANDN U23153 ( .A(n27130), .B(n18720), .Z(n18721) );
  NANDN U23154 ( .A(n27133), .B(n18721), .Z(n18722) );
  NANDN U23155 ( .A(n27135), .B(n18722), .Z(n18723) );
  NAND U23156 ( .A(n18724), .B(n18723), .Z(n18725) );
  NANDN U23157 ( .A(n18725), .B(n27138), .Z(n18726) );
  AND U23158 ( .A(n27140), .B(n18726), .Z(n18729) );
  ANDN U23159 ( .B(n18728), .A(n18727), .Z(n27143) );
  NANDN U23160 ( .A(n18729), .B(n27143), .Z(n18732) );
  NANDN U23161 ( .A(y[3342]), .B(x[3342]), .Z(n18731) );
  ANDN U23162 ( .B(n18731), .A(n18730), .Z(n27144) );
  NAND U23163 ( .A(n18732), .B(n27144), .Z(n18733) );
  NANDN U23164 ( .A(n27147), .B(n18733), .Z(n18734) );
  NANDN U23165 ( .A(n27149), .B(n18734), .Z(n18735) );
  AND U23166 ( .A(n27150), .B(n18735), .Z(n18738) );
  NANDN U23167 ( .A(y[3346]), .B(x[3346]), .Z(n18737) );
  ANDN U23168 ( .B(n18737), .A(n18736), .Z(n27153) );
  NANDN U23169 ( .A(n18738), .B(n27153), .Z(n18741) );
  NOR U23170 ( .A(n18740), .B(n18739), .Z(n27154) );
  NAND U23171 ( .A(n18741), .B(n27154), .Z(n18742) );
  NANDN U23172 ( .A(n27157), .B(n18742), .Z(n18743) );
  NANDN U23173 ( .A(n27159), .B(n18743), .Z(n18744) );
  AND U23174 ( .A(n27160), .B(n18744), .Z(n18745) );
  OR U23175 ( .A(n27162), .B(n18745), .Z(n18748) );
  NANDN U23176 ( .A(y[3353]), .B(x[3353]), .Z(n18747) );
  ANDN U23177 ( .B(n18747), .A(n18746), .Z(n27164) );
  NAND U23178 ( .A(n18748), .B(n27164), .Z(n18749) );
  NANDN U23179 ( .A(n27167), .B(n18749), .Z(n18752) );
  NANDN U23180 ( .A(y[3354]), .B(x[3354]), .Z(n18751) );
  ANDN U23181 ( .B(n18751), .A(n18750), .Z(n27168) );
  NAND U23182 ( .A(n18752), .B(n27168), .Z(n18753) );
  AND U23183 ( .A(n27172), .B(n18753), .Z(n18755) );
  NAND U23184 ( .A(n18755), .B(n18754), .Z(n18758) );
  NANDN U23185 ( .A(y[3356]), .B(x[3356]), .Z(n18757) );
  ANDN U23186 ( .B(n18757), .A(n18756), .Z(n27174) );
  NAND U23187 ( .A(n18758), .B(n27174), .Z(n18759) );
  NAND U23188 ( .A(n18760), .B(n18759), .Z(n18761) );
  NANDN U23189 ( .A(n18761), .B(n27178), .Z(n18762) );
  AND U23190 ( .A(n27180), .B(n18762), .Z(n18766) );
  NAND U23191 ( .A(n18763), .B(y[3359]), .Z(n18765) );
  ANDN U23192 ( .B(n18765), .A(n18764), .Z(n27183) );
  NANDN U23193 ( .A(n18766), .B(n27183), .Z(n18769) );
  NOR U23194 ( .A(n18768), .B(n18767), .Z(n27184) );
  NAND U23195 ( .A(n18769), .B(n27184), .Z(n18770) );
  NANDN U23196 ( .A(n27187), .B(n18770), .Z(n18771) );
  NANDN U23197 ( .A(n27189), .B(n18771), .Z(n18772) );
  AND U23198 ( .A(n27190), .B(n18772), .Z(n18775) );
  OR U23199 ( .A(n18774), .B(n18773), .Z(n27192) );
  OR U23200 ( .A(n18775), .B(n27192), .Z(n18776) );
  NAND U23201 ( .A(n18777), .B(n18776), .Z(n18778) );
  NANDN U23202 ( .A(n18778), .B(n27195), .Z(n18779) );
  AND U23203 ( .A(n27198), .B(n18779), .Z(n18780) );
  OR U23204 ( .A(n27200), .B(n18780), .Z(n18783) );
  ANDN U23205 ( .B(n18782), .A(n18781), .Z(n27202) );
  NAND U23206 ( .A(n18783), .B(n27202), .Z(n18786) );
  NANDN U23207 ( .A(x[3369]), .B(y[3369]), .Z(n18785) );
  ANDN U23208 ( .B(n18785), .A(n18784), .Z(n27204) );
  NAND U23209 ( .A(n18786), .B(n27204), .Z(n18787) );
  NANDN U23210 ( .A(n27207), .B(n18787), .Z(n18788) );
  AND U23211 ( .A(n27208), .B(n18788), .Z(n18789) );
  OR U23212 ( .A(n27210), .B(n18789), .Z(n18792) );
  NANDN U23213 ( .A(x[3373]), .B(y[3373]), .Z(n18791) );
  ANDN U23214 ( .B(n18791), .A(n18790), .Z(n27212) );
  NAND U23215 ( .A(n18792), .B(n27212), .Z(n18793) );
  NANDN U23216 ( .A(n27215), .B(n18793), .Z(n18794) );
  NANDN U23217 ( .A(n27217), .B(n18794), .Z(n18795) );
  AND U23218 ( .A(n27218), .B(n18795), .Z(n18796) );
  OR U23219 ( .A(n27220), .B(n18796), .Z(n18797) );
  NAND U23220 ( .A(n18797), .B(n27222), .Z(n18798) );
  NAND U23221 ( .A(n18798), .B(n27225), .Z(n18801) );
  NANDN U23222 ( .A(y[3381]), .B(x[3381]), .Z(n18800) );
  ANDN U23223 ( .B(n18800), .A(n18799), .Z(n27226) );
  NAND U23224 ( .A(n18801), .B(n27226), .Z(n18802) );
  NANDN U23225 ( .A(n27228), .B(n18802), .Z(n18803) );
  AND U23226 ( .A(n27230), .B(n18803), .Z(n18804) );
  OR U23227 ( .A(n27232), .B(n18804), .Z(n18807) );
  NANDN U23228 ( .A(y[3384]), .B(x[3384]), .Z(n18806) );
  ANDN U23229 ( .B(n18806), .A(n18805), .Z(n27234) );
  NAND U23230 ( .A(n18807), .B(n27234), .Z(n18808) );
  NANDN U23231 ( .A(n27237), .B(n18808), .Z(n18811) );
  NANDN U23232 ( .A(y[3386]), .B(x[3386]), .Z(n18810) );
  ANDN U23233 ( .B(n18810), .A(n18809), .Z(n27238) );
  NAND U23234 ( .A(n18811), .B(n27238), .Z(n18812) );
  AND U23235 ( .A(n27240), .B(n18812), .Z(n18815) );
  OR U23236 ( .A(n18814), .B(n18813), .Z(n27242) );
  OR U23237 ( .A(n18815), .B(n27242), .Z(n18816) );
  NAND U23238 ( .A(n18817), .B(n18816), .Z(n18818) );
  NANDN U23239 ( .A(n18818), .B(n27245), .Z(n18819) );
  AND U23240 ( .A(n27248), .B(n18819), .Z(n18822) );
  NANDN U23241 ( .A(x[3391]), .B(y[3391]), .Z(n18821) );
  ANDN U23242 ( .B(n18821), .A(n18820), .Z(n27251) );
  NANDN U23243 ( .A(n18822), .B(n27251), .Z(n18825) );
  NOR U23244 ( .A(n18824), .B(n18823), .Z(n27252) );
  NAND U23245 ( .A(n18825), .B(n27252), .Z(n18826) );
  NANDN U23246 ( .A(n27255), .B(n18826), .Z(n18827) );
  NANDN U23247 ( .A(n27257), .B(n18827), .Z(n18828) );
  AND U23248 ( .A(n27258), .B(n18828), .Z(n18829) );
  OR U23249 ( .A(n27260), .B(n18829), .Z(n18832) );
  NANDN U23250 ( .A(x[3398]), .B(y[3398]), .Z(n18831) );
  ANDN U23251 ( .B(n18831), .A(n18830), .Z(n27262) );
  NAND U23252 ( .A(n18832), .B(n27262), .Z(n18833) );
  NANDN U23253 ( .A(n27265), .B(n18833), .Z(n18836) );
  NANDN U23254 ( .A(x[3399]), .B(y[3399]), .Z(n18835) );
  ANDN U23255 ( .B(n18835), .A(n18834), .Z(n27266) );
  NAND U23256 ( .A(n18836), .B(n27266), .Z(n18837) );
  AND U23257 ( .A(n27268), .B(n18837), .Z(n18838) );
  OR U23258 ( .A(n27270), .B(n18838), .Z(n18841) );
  AND U23259 ( .A(n18840), .B(n18839), .Z(n27272) );
  NAND U23260 ( .A(n18841), .B(n27272), .Z(n18844) );
  NANDN U23261 ( .A(x[3403]), .B(y[3403]), .Z(n18843) );
  ANDN U23262 ( .B(n18843), .A(n18842), .Z(n27274) );
  NAND U23263 ( .A(n18844), .B(n27274), .Z(n18845) );
  NANDN U23264 ( .A(n27277), .B(n18845), .Z(n18846) );
  AND U23265 ( .A(n27278), .B(n18846), .Z(n18847) );
  OR U23266 ( .A(n27280), .B(n18847), .Z(n18850) );
  NANDN U23267 ( .A(x[3407]), .B(y[3407]), .Z(n18849) );
  ANDN U23268 ( .B(n18849), .A(n18848), .Z(n27282) );
  NAND U23269 ( .A(n18850), .B(n27282), .Z(n18851) );
  NANDN U23270 ( .A(n27285), .B(n18851), .Z(n18852) );
  NAND U23271 ( .A(n18853), .B(n18852), .Z(n18854) );
  AND U23272 ( .A(n27290), .B(n18854), .Z(n18857) );
  NANDN U23273 ( .A(x[3411]), .B(y[3411]), .Z(n18856) );
  ANDN U23274 ( .B(n18856), .A(n18855), .Z(n27293) );
  NANDN U23275 ( .A(n18857), .B(n27293), .Z(n18860) );
  NANDN U23276 ( .A(y[3413]), .B(x[3413]), .Z(n18859) );
  ANDN U23277 ( .B(n18859), .A(n18858), .Z(n27294) );
  NAND U23278 ( .A(n18860), .B(n27294), .Z(n18861) );
  NANDN U23279 ( .A(n27297), .B(n18861), .Z(n18864) );
  NANDN U23280 ( .A(y[3414]), .B(x[3414]), .Z(n18863) );
  ANDN U23281 ( .B(n18863), .A(n18862), .Z(n27298) );
  NAND U23282 ( .A(n18864), .B(n27298), .Z(n18865) );
  AND U23283 ( .A(n27300), .B(n18865), .Z(n18866) );
  OR U23284 ( .A(n27302), .B(n18866), .Z(n18869) );
  AND U23285 ( .A(n18868), .B(n18867), .Z(n27304) );
  NAND U23286 ( .A(n18869), .B(n27304), .Z(n18872) );
  NANDN U23287 ( .A(y[3418]), .B(x[3418]), .Z(n18871) );
  ANDN U23288 ( .B(n18871), .A(n18870), .Z(n27306) );
  NAND U23289 ( .A(n18872), .B(n27306), .Z(n18873) );
  NANDN U23290 ( .A(n27309), .B(n18873), .Z(n18874) );
  AND U23291 ( .A(n27310), .B(n18874), .Z(n18875) );
  OR U23292 ( .A(n27312), .B(n18875), .Z(n18878) );
  NANDN U23293 ( .A(y[3423]), .B(x[3423]), .Z(n18877) );
  NANDN U23294 ( .A(y[3422]), .B(x[3422]), .Z(n18876) );
  AND U23295 ( .A(n18877), .B(n18876), .Z(n27314) );
  NAND U23296 ( .A(n18878), .B(n27314), .Z(n18879) );
  NANDN U23297 ( .A(n27317), .B(n18879), .Z(n18882) );
  NANDN U23298 ( .A(y[3424]), .B(x[3424]), .Z(n18881) );
  ANDN U23299 ( .B(n18881), .A(n18880), .Z(n27318) );
  NAND U23300 ( .A(n18882), .B(n27318), .Z(n18883) );
  AND U23301 ( .A(n27320), .B(n18883), .Z(n18884) );
  OR U23302 ( .A(n27322), .B(n18884), .Z(n18887) );
  NANDN U23303 ( .A(x[3428]), .B(y[3428]), .Z(n18886) );
  AND U23304 ( .A(n18886), .B(n18885), .Z(n27324) );
  NAND U23305 ( .A(n18887), .B(n27324), .Z(n18888) );
  NANDN U23306 ( .A(n27327), .B(n18888), .Z(n18889) );
  NANDN U23307 ( .A(n27329), .B(n18889), .Z(n18892) );
  OR U23308 ( .A(n18891), .B(n18890), .Z(n27331) );
  ANDN U23309 ( .B(n18892), .A(n27331), .Z(n18893) );
  ANDN U23310 ( .B(n20227), .A(n18893), .Z(n18895) );
  NAND U23311 ( .A(n18895), .B(n18894), .Z(n18896) );
  NANDN U23312 ( .A(n27335), .B(n18896), .Z(n18899) );
  NANDN U23313 ( .A(x[3433]), .B(y[3433]), .Z(n18897) );
  NAND U23314 ( .A(n18898), .B(n18897), .Z(n27337) );
  ANDN U23315 ( .B(n18899), .A(n27337), .Z(n18900) );
  OR U23316 ( .A(n27339), .B(n18900), .Z(n18903) );
  ANDN U23317 ( .B(n18902), .A(n18901), .Z(n27340) );
  NAND U23318 ( .A(n18903), .B(n27340), .Z(n18906) );
  NANDN U23319 ( .A(y[3436]), .B(x[3436]), .Z(n18905) );
  ANDN U23320 ( .B(n18905), .A(n18904), .Z(n27343) );
  NAND U23321 ( .A(n18906), .B(n27343), .Z(n18907) );
  NANDN U23322 ( .A(n27345), .B(n18907), .Z(n18910) );
  NANDN U23323 ( .A(y[3439]), .B(x[3439]), .Z(n18908) );
  NANDN U23324 ( .A(n18909), .B(n18908), .Z(n27347) );
  ANDN U23325 ( .B(n18910), .A(n27347), .Z(n18911) );
  OR U23326 ( .A(n27349), .B(n18911), .Z(n18914) );
  NANDN U23327 ( .A(y[3440]), .B(x[3440]), .Z(n18913) );
  ANDN U23328 ( .B(n18913), .A(n18912), .Z(n27350) );
  NAND U23329 ( .A(n18914), .B(n27350), .Z(n18915) );
  NANDN U23330 ( .A(n27352), .B(n18915), .Z(n18916) );
  NANDN U23331 ( .A(n27355), .B(n18916), .Z(n18919) );
  NAND U23332 ( .A(n18918), .B(n18917), .Z(n27357) );
  ANDN U23333 ( .B(n18919), .A(n27357), .Z(n18922) );
  NANDN U23334 ( .A(y[3444]), .B(x[3444]), .Z(n18921) );
  ANDN U23335 ( .B(n18921), .A(n18920), .Z(n27358) );
  NANDN U23336 ( .A(n18922), .B(n27358), .Z(n18925) );
  NOR U23337 ( .A(n18924), .B(n18923), .Z(n27360) );
  NAND U23338 ( .A(n18925), .B(n27360), .Z(n18926) );
  NANDN U23339 ( .A(n27362), .B(n18926), .Z(n18927) );
  NANDN U23340 ( .A(n27365), .B(n18927), .Z(n18930) );
  NANDN U23341 ( .A(y[3448]), .B(x[3448]), .Z(n18928) );
  NAND U23342 ( .A(n18929), .B(n18928), .Z(n27367) );
  ANDN U23343 ( .B(n18930), .A(n27367), .Z(n18931) );
  OR U23344 ( .A(n27369), .B(n18931), .Z(n18934) );
  NANDN U23345 ( .A(y[3451]), .B(x[3451]), .Z(n18933) );
  ANDN U23346 ( .B(n18933), .A(n18932), .Z(n27370) );
  NAND U23347 ( .A(n18934), .B(n27370), .Z(n18935) );
  NANDN U23348 ( .A(n27372), .B(n18935), .Z(n18938) );
  NANDN U23349 ( .A(y[3452]), .B(x[3452]), .Z(n18937) );
  ANDN U23350 ( .B(n18937), .A(n18936), .Z(n27374) );
  NAND U23351 ( .A(n18938), .B(n27374), .Z(n18941) );
  OR U23352 ( .A(n18940), .B(n18939), .Z(n27377) );
  ANDN U23353 ( .B(n18941), .A(n27377), .Z(n18942) );
  OR U23354 ( .A(n27379), .B(n18942), .Z(n18945) );
  AND U23355 ( .A(n18944), .B(n18943), .Z(n27380) );
  NAND U23356 ( .A(n18945), .B(n27380), .Z(n18948) );
  NANDN U23357 ( .A(y[3456]), .B(x[3456]), .Z(n18947) );
  ANDN U23358 ( .B(n18947), .A(n18946), .Z(n27383) );
  NAND U23359 ( .A(n18948), .B(n27383), .Z(n18949) );
  NANDN U23360 ( .A(n27385), .B(n18949), .Z(n18952) );
  NANDN U23361 ( .A(y[3459]), .B(x[3459]), .Z(n18950) );
  NANDN U23362 ( .A(n18951), .B(n18950), .Z(n27387) );
  ANDN U23363 ( .B(n18952), .A(n27387), .Z(n18953) );
  OR U23364 ( .A(n27389), .B(n18953), .Z(n18956) );
  NANDN U23365 ( .A(y[3460]), .B(x[3460]), .Z(n18955) );
  ANDN U23366 ( .B(n18955), .A(n18954), .Z(n27390) );
  NAND U23367 ( .A(n18956), .B(n27390), .Z(n18957) );
  NANDN U23368 ( .A(n27392), .B(n18957), .Z(n18958) );
  NANDN U23369 ( .A(n27395), .B(n18958), .Z(n18961) );
  NAND U23370 ( .A(n18960), .B(n18959), .Z(n27397) );
  ANDN U23371 ( .B(n18961), .A(n27397), .Z(n18964) );
  NANDN U23372 ( .A(y[3464]), .B(x[3464]), .Z(n18963) );
  ANDN U23373 ( .B(n18963), .A(n18962), .Z(n27398) );
  NANDN U23374 ( .A(n18964), .B(n27398), .Z(n18967) );
  NOR U23375 ( .A(n18966), .B(n18965), .Z(n27400) );
  NAND U23376 ( .A(n18967), .B(n27400), .Z(n18968) );
  NANDN U23377 ( .A(n27402), .B(n18968), .Z(n18969) );
  NANDN U23378 ( .A(n27405), .B(n18969), .Z(n18972) );
  NANDN U23379 ( .A(y[3468]), .B(x[3468]), .Z(n18970) );
  NANDN U23380 ( .A(n18971), .B(n18970), .Z(n27407) );
  ANDN U23381 ( .B(n18972), .A(n27407), .Z(n18973) );
  ANDN U23382 ( .B(n27410), .A(n18973), .Z(n18976) );
  XOR U23383 ( .A(n18974), .B(y[3470]), .Z(n18975) );
  NAND U23384 ( .A(n18976), .B(n18975), .Z(n18977) );
  NANDN U23385 ( .A(n27413), .B(n18977), .Z(n18980) );
  NANDN U23386 ( .A(x[3471]), .B(y[3471]), .Z(n18978) );
  NANDN U23387 ( .A(n18979), .B(n18978), .Z(n27414) );
  ANDN U23388 ( .B(n18980), .A(n27414), .Z(n18981) );
  OR U23389 ( .A(n27417), .B(n18981), .Z(n18982) );
  NANDN U23390 ( .A(n27419), .B(n18982), .Z(n18983) );
  NANDN U23391 ( .A(n27421), .B(n18983), .Z(n18984) );
  NANDN U23392 ( .A(n27423), .B(n18984), .Z(n18988) );
  NAND U23393 ( .A(n18985), .B(x[3476]), .Z(n18986) );
  NANDN U23394 ( .A(n18987), .B(n18986), .Z(n27424) );
  ANDN U23395 ( .B(n18988), .A(n27424), .Z(n18989) );
  ANDN U23396 ( .B(n27427), .A(n18989), .Z(n18991) );
  NAND U23397 ( .A(n18991), .B(n18990), .Z(n18994) );
  NANDN U23398 ( .A(y[3478]), .B(x[3478]), .Z(n18993) );
  ANDN U23399 ( .B(n18993), .A(n18992), .Z(n27430) );
  NAND U23400 ( .A(n18994), .B(n27430), .Z(n18998) );
  NAND U23401 ( .A(n18995), .B(y[3480]), .Z(n18996) );
  NANDN U23402 ( .A(n18997), .B(n18996), .Z(n27432) );
  ANDN U23403 ( .B(n18998), .A(n27432), .Z(n19001) );
  NANDN U23404 ( .A(y[3480]), .B(x[3480]), .Z(n19000) );
  ANDN U23405 ( .B(n19000), .A(n18999), .Z(n27434) );
  NANDN U23406 ( .A(n19001), .B(n27434), .Z(n19002) );
  NANDN U23407 ( .A(n27437), .B(n19002), .Z(n19005) );
  NANDN U23408 ( .A(y[3482]), .B(x[3482]), .Z(n19004) );
  ANDN U23409 ( .B(n19004), .A(n19003), .Z(n27438) );
  NAND U23410 ( .A(n19005), .B(n27438), .Z(n19006) );
  NANDN U23411 ( .A(n27441), .B(n19006), .Z(n19009) );
  NANDN U23412 ( .A(y[3484]), .B(x[3484]), .Z(n19007) );
  NAND U23413 ( .A(n19008), .B(n19007), .Z(n27442) );
  ANDN U23414 ( .B(n19009), .A(n27442), .Z(n19010) );
  OR U23415 ( .A(n27445), .B(n19010), .Z(n19011) );
  NANDN U23416 ( .A(n27447), .B(n19011), .Z(n19012) );
  NANDN U23417 ( .A(n27449), .B(n19012), .Z(n19013) );
  NAND U23418 ( .A(n19013), .B(n27450), .Z(n19014) );
  NAND U23419 ( .A(n19014), .B(n27452), .Z(n19015) );
  AND U23420 ( .A(n27455), .B(n19015), .Z(n19016) );
  NANDN U23421 ( .A(n19016), .B(n27456), .Z(n19017) );
  AND U23422 ( .A(n27459), .B(n19017), .Z(n19020) );
  NOR U23423 ( .A(n19019), .B(n19018), .Z(n27460) );
  NANDN U23424 ( .A(n19020), .B(n27460), .Z(n19021) );
  NANDN U23425 ( .A(n27463), .B(n19021), .Z(n19024) );
  NANDN U23426 ( .A(x[3495]), .B(y[3495]), .Z(n19023) );
  ANDN U23427 ( .B(n19023), .A(n19022), .Z(n27464) );
  NAND U23428 ( .A(n19024), .B(n27464), .Z(n19025) );
  NANDN U23429 ( .A(n27467), .B(n19025), .Z(n19028) );
  NANDN U23430 ( .A(x[3497]), .B(y[3497]), .Z(n19026) );
  NAND U23431 ( .A(n19027), .B(n19026), .Z(n27468) );
  ANDN U23432 ( .B(n19028), .A(n27468), .Z(n19029) );
  OR U23433 ( .A(n27471), .B(n19029), .Z(n19030) );
  NANDN U23434 ( .A(n27473), .B(n19030), .Z(n19031) );
  NANDN U23435 ( .A(n27475), .B(n19031), .Z(n19032) );
  NAND U23436 ( .A(n19033), .B(n19032), .Z(n19034) );
  AND U23437 ( .A(n27480), .B(n19034), .Z(n19035) );
  OR U23438 ( .A(n27483), .B(n19035), .Z(n19036) );
  NANDN U23439 ( .A(n27485), .B(n19036), .Z(n19039) );
  NANDN U23440 ( .A(x[3505]), .B(y[3505]), .Z(n19038) );
  ANDN U23441 ( .B(n19038), .A(n19037), .Z(n27486) );
  NAND U23442 ( .A(n19039), .B(n27486), .Z(n19040) );
  NANDN U23443 ( .A(n27489), .B(n19040), .Z(n19043) );
  OR U23444 ( .A(n19042), .B(n19041), .Z(n27490) );
  ANDN U23445 ( .B(n19043), .A(n27490), .Z(n19046) );
  ANDN U23446 ( .B(n19045), .A(n19044), .Z(n27492) );
  NANDN U23447 ( .A(n19046), .B(n27492), .Z(n19047) );
  NANDN U23448 ( .A(n27495), .B(n19047), .Z(n19050) );
  NANDN U23449 ( .A(y[3510]), .B(x[3510]), .Z(n19049) );
  ANDN U23450 ( .B(n19049), .A(n19048), .Z(n27496) );
  NAND U23451 ( .A(n19050), .B(n27496), .Z(n19051) );
  NANDN U23452 ( .A(n27499), .B(n19051), .Z(n19054) );
  NANDN U23453 ( .A(y[3512]), .B(x[3512]), .Z(n19052) );
  NAND U23454 ( .A(n19053), .B(n19052), .Z(n27500) );
  ANDN U23455 ( .B(n19054), .A(n27500), .Z(n19055) );
  OR U23456 ( .A(n27503), .B(n19055), .Z(n19056) );
  NANDN U23457 ( .A(n27505), .B(n19056), .Z(n19057) );
  NANDN U23458 ( .A(n27507), .B(n19057), .Z(n19060) );
  NANDN U23459 ( .A(y[3516]), .B(x[3516]), .Z(n19059) );
  ANDN U23460 ( .B(n19059), .A(n19058), .Z(n27508) );
  NAND U23461 ( .A(n19060), .B(n27508), .Z(n19064) );
  NAND U23462 ( .A(n19061), .B(y[3518]), .Z(n19062) );
  NANDN U23463 ( .A(n19063), .B(n19062), .Z(n27510) );
  ANDN U23464 ( .B(n19064), .A(n27510), .Z(n19067) );
  NANDN U23465 ( .A(y[3518]), .B(x[3518]), .Z(n19066) );
  ANDN U23466 ( .B(n19066), .A(n19065), .Z(n27512) );
  NANDN U23467 ( .A(n19067), .B(n27512), .Z(n19068) );
  NANDN U23468 ( .A(n27515), .B(n19068), .Z(n19069) );
  NANDN U23469 ( .A(n27517), .B(n19069), .Z(n19070) );
  NANDN U23470 ( .A(n27519), .B(n19070), .Z(n19073) );
  NANDN U23471 ( .A(n19072), .B(n19071), .Z(n27520) );
  ANDN U23472 ( .B(n19073), .A(n27520), .Z(n19074) );
  ANDN U23473 ( .B(n27523), .A(n19074), .Z(n19076) );
  NAND U23474 ( .A(n19076), .B(n19075), .Z(n19079) );
  NANDN U23475 ( .A(y[3524]), .B(x[3524]), .Z(n19078) );
  ANDN U23476 ( .B(n19078), .A(n19077), .Z(n27526) );
  NAND U23477 ( .A(n19079), .B(n27526), .Z(n19083) );
  NAND U23478 ( .A(n19080), .B(y[3526]), .Z(n19081) );
  NANDN U23479 ( .A(n19082), .B(n19081), .Z(n27528) );
  ANDN U23480 ( .B(n19083), .A(n27528), .Z(n19086) );
  NANDN U23481 ( .A(y[3526]), .B(x[3526]), .Z(n19085) );
  ANDN U23482 ( .B(n19085), .A(n19084), .Z(n27530) );
  NANDN U23483 ( .A(n19086), .B(n27530), .Z(n19087) );
  NANDN U23484 ( .A(n27533), .B(n19087), .Z(n19088) );
  NANDN U23485 ( .A(n27535), .B(n19088), .Z(n19089) );
  NANDN U23486 ( .A(n27537), .B(n19089), .Z(n19092) );
  NANDN U23487 ( .A(n19091), .B(n19090), .Z(n27538) );
  ANDN U23488 ( .B(n19092), .A(n27538), .Z(n19093) );
  ANDN U23489 ( .B(n27541), .A(n19093), .Z(n19095) );
  NAND U23490 ( .A(n19095), .B(n19094), .Z(n19098) );
  NANDN U23491 ( .A(y[3532]), .B(x[3532]), .Z(n19097) );
  ANDN U23492 ( .B(n19097), .A(n19096), .Z(n27544) );
  NAND U23493 ( .A(n19098), .B(n27544), .Z(n19102) );
  NAND U23494 ( .A(n19099), .B(y[3534]), .Z(n19100) );
  NANDN U23495 ( .A(n19101), .B(n19100), .Z(n27546) );
  ANDN U23496 ( .B(n19102), .A(n27546), .Z(n19105) );
  NANDN U23497 ( .A(y[3534]), .B(x[3534]), .Z(n19104) );
  ANDN U23498 ( .B(n19104), .A(n19103), .Z(n27548) );
  NANDN U23499 ( .A(n19105), .B(n27548), .Z(n19106) );
  NANDN U23500 ( .A(n27551), .B(n19106), .Z(n19109) );
  NANDN U23501 ( .A(y[3536]), .B(x[3536]), .Z(n19108) );
  ANDN U23502 ( .B(n19108), .A(n19107), .Z(n27552) );
  NAND U23503 ( .A(n19109), .B(n27552), .Z(n19110) );
  NANDN U23504 ( .A(n27555), .B(n19110), .Z(n19113) );
  NANDN U23505 ( .A(y[3538]), .B(x[3538]), .Z(n19111) );
  NANDN U23506 ( .A(n19112), .B(n19111), .Z(n27556) );
  ANDN U23507 ( .B(n19113), .A(n27556), .Z(n19114) );
  OR U23508 ( .A(n27559), .B(n19114), .Z(n19115) );
  NANDN U23509 ( .A(n27561), .B(n19115), .Z(n19116) );
  NAND U23510 ( .A(n19116), .B(n27564), .Z(n19117) );
  ANDN U23511 ( .B(n19118), .A(n19117), .Z(n19121) );
  NANDN U23512 ( .A(y[3542]), .B(x[3542]), .Z(n19120) );
  ANDN U23513 ( .B(n19120), .A(n19119), .Z(n27566) );
  NANDN U23514 ( .A(n19121), .B(n27566), .Z(n19122) );
  NANDN U23515 ( .A(n27568), .B(n19122), .Z(n19125) );
  NANDN U23516 ( .A(y[3544]), .B(x[3544]), .Z(n19124) );
  ANDN U23517 ( .B(n19124), .A(n19123), .Z(n27570) );
  NAND U23518 ( .A(n19125), .B(n27570), .Z(n19126) );
  NANDN U23519 ( .A(n27573), .B(n19126), .Z(n19127) );
  AND U23520 ( .A(n27574), .B(n19127), .Z(n19128) );
  OR U23521 ( .A(n27577), .B(n19128), .Z(n19129) );
  NANDN U23522 ( .A(n27578), .B(n19129), .Z(n19130) );
  NANDN U23523 ( .A(n27581), .B(n19130), .Z(n19133) );
  NANDN U23524 ( .A(y[3550]), .B(x[3550]), .Z(n19132) );
  ANDN U23525 ( .B(n19132), .A(n19131), .Z(n27582) );
  NAND U23526 ( .A(n19133), .B(n27582), .Z(n19134) );
  AND U23527 ( .A(n27584), .B(n19134), .Z(n19137) );
  NANDN U23528 ( .A(y[3552]), .B(x[3552]), .Z(n19136) );
  ANDN U23529 ( .B(n19136), .A(n19135), .Z(n27586) );
  NANDN U23530 ( .A(n19137), .B(n27586), .Z(n19138) );
  NANDN U23531 ( .A(n27588), .B(n19138), .Z(n19141) );
  NANDN U23532 ( .A(y[3554]), .B(x[3554]), .Z(n19140) );
  ANDN U23533 ( .B(n19140), .A(n19139), .Z(n27590) );
  NAND U23534 ( .A(n19141), .B(n27590), .Z(n19142) );
  NANDN U23535 ( .A(n27593), .B(n19142), .Z(n19143) );
  AND U23536 ( .A(n27594), .B(n19143), .Z(n19144) );
  OR U23537 ( .A(n27597), .B(n19144), .Z(n19145) );
  NANDN U23538 ( .A(n27598), .B(n19145), .Z(n19146) );
  NAND U23539 ( .A(n19146), .B(n20225), .Z(n19148) );
  NANDN U23540 ( .A(n19148), .B(n19147), .Z(n19151) );
  NANDN U23541 ( .A(y[3560]), .B(x[3560]), .Z(n19150) );
  ANDN U23542 ( .B(n19150), .A(n19149), .Z(n27602) );
  NAND U23543 ( .A(n19151), .B(n27602), .Z(n19152) );
  NAND U23544 ( .A(n19153), .B(n19152), .Z(n19154) );
  NANDN U23545 ( .A(n19154), .B(n27605), .Z(n19155) );
  AND U23546 ( .A(n27608), .B(n19155), .Z(n19158) );
  NOR U23547 ( .A(n19157), .B(n19156), .Z(n27610) );
  NANDN U23548 ( .A(n19158), .B(n27610), .Z(n19159) );
  NANDN U23549 ( .A(n27613), .B(n19159), .Z(n19162) );
  NOR U23550 ( .A(n19161), .B(n19160), .Z(n27614) );
  NAND U23551 ( .A(n19162), .B(n27614), .Z(n19163) );
  NANDN U23552 ( .A(n27617), .B(n19163), .Z(n19166) );
  NANDN U23553 ( .A(x[3567]), .B(y[3567]), .Z(n19164) );
  NAND U23554 ( .A(n19165), .B(n19164), .Z(n27618) );
  ANDN U23555 ( .B(n19166), .A(n27618), .Z(n19167) );
  OR U23556 ( .A(n27621), .B(n19167), .Z(n19168) );
  NANDN U23557 ( .A(n27623), .B(n19168), .Z(n19169) );
  NANDN U23558 ( .A(n27625), .B(n19169), .Z(n19170) );
  NAND U23559 ( .A(n19171), .B(n19170), .Z(n19172) );
  NANDN U23560 ( .A(n27631), .B(n19172), .Z(n19175) );
  OR U23561 ( .A(n19174), .B(n19173), .Z(n27633) );
  ANDN U23562 ( .B(n19175), .A(n27633), .Z(n19178) );
  ANDN U23563 ( .B(n19177), .A(n19176), .Z(n27634) );
  NANDN U23564 ( .A(n19178), .B(n27634), .Z(n19181) );
  NANDN U23565 ( .A(x[3575]), .B(y[3575]), .Z(n19180) );
  ANDN U23566 ( .B(n19180), .A(n19179), .Z(n27636) );
  NAND U23567 ( .A(n19181), .B(n27636), .Z(n19182) );
  NANDN U23568 ( .A(n27639), .B(n19182), .Z(n19183) );
  NANDN U23569 ( .A(n27640), .B(n19183), .Z(n19184) );
  AND U23570 ( .A(n27642), .B(n19184), .Z(n19185) );
  OR U23571 ( .A(n27645), .B(n19185), .Z(n19188) );
  NANDN U23572 ( .A(y[3580]), .B(x[3580]), .Z(n19187) );
  ANDN U23573 ( .B(n19187), .A(n19186), .Z(n27646) );
  NAND U23574 ( .A(n19188), .B(n27646), .Z(n19189) );
  NANDN U23575 ( .A(n27649), .B(n19189), .Z(n19190) );
  NANDN U23576 ( .A(n27650), .B(n19190), .Z(n19191) );
  AND U23577 ( .A(n19192), .B(n19191), .Z(n19193) );
  OR U23578 ( .A(n27657), .B(n19193), .Z(n19194) );
  NANDN U23579 ( .A(n27658), .B(n19194), .Z(n19197) );
  NOR U23580 ( .A(n19196), .B(n19195), .Z(n27660) );
  NAND U23581 ( .A(n19197), .B(n27660), .Z(n19198) );
  NAND U23582 ( .A(n19199), .B(n19198), .Z(n19200) );
  AND U23583 ( .A(n27666), .B(n19200), .Z(n19201) );
  OR U23584 ( .A(n27669), .B(n19201), .Z(n19202) );
  NANDN U23585 ( .A(n27671), .B(n19202), .Z(n19203) );
  NANDN U23586 ( .A(n27673), .B(n19203), .Z(n19206) );
  NANDN U23587 ( .A(y[3592]), .B(x[3592]), .Z(n19205) );
  ANDN U23588 ( .B(n19205), .A(n19204), .Z(n27674) );
  NAND U23589 ( .A(n19206), .B(n27674), .Z(n19210) );
  NAND U23590 ( .A(n19207), .B(y[3594]), .Z(n19208) );
  NANDN U23591 ( .A(n19209), .B(n19208), .Z(n27676) );
  ANDN U23592 ( .B(n19210), .A(n27676), .Z(n19211) );
  OR U23593 ( .A(n27679), .B(n19211), .Z(n19212) );
  NANDN U23594 ( .A(n27681), .B(n19212), .Z(n19215) );
  NOR U23595 ( .A(n19214), .B(n19213), .Z(n27682) );
  NAND U23596 ( .A(n19215), .B(n27682), .Z(n19216) );
  NAND U23597 ( .A(n19217), .B(n19216), .Z(n19218) );
  AND U23598 ( .A(n27688), .B(n19218), .Z(n19219) );
  ANDN U23599 ( .B(n27692), .A(n19219), .Z(n19221) );
  AND U23600 ( .A(n19221), .B(n19220), .Z(n19224) );
  NANDN U23601 ( .A(y[3600]), .B(x[3600]), .Z(n19223) );
  ANDN U23602 ( .B(n19223), .A(n19222), .Z(n27694) );
  NANDN U23603 ( .A(n19224), .B(n27694), .Z(n19225) );
  NANDN U23604 ( .A(n27696), .B(n19225), .Z(n19226) );
  NANDN U23605 ( .A(n27699), .B(n19226), .Z(n19227) );
  NAND U23606 ( .A(n19228), .B(n19227), .Z(n19231) );
  NANDN U23607 ( .A(y[3604]), .B(x[3604]), .Z(n19230) );
  ANDN U23608 ( .B(n19230), .A(n19229), .Z(n27704) );
  NAND U23609 ( .A(n19231), .B(n27704), .Z(n19232) );
  NAND U23610 ( .A(n19233), .B(n19232), .Z(n19234) );
  NANDN U23611 ( .A(n19234), .B(n27708), .Z(n19235) );
  AND U23612 ( .A(n27710), .B(n19235), .Z(n19238) );
  NOR U23613 ( .A(n19237), .B(n19236), .Z(n27713) );
  NANDN U23614 ( .A(n19238), .B(n27713), .Z(n19241) );
  NANDN U23615 ( .A(y[3609]), .B(x[3609]), .Z(n19240) );
  ANDN U23616 ( .B(n19240), .A(n19239), .Z(n27714) );
  NAND U23617 ( .A(n19241), .B(n27714), .Z(n19244) );
  NANDN U23618 ( .A(x[3609]), .B(y[3609]), .Z(n19243) );
  ANDN U23619 ( .B(n19243), .A(n19242), .Z(n27716) );
  NAND U23620 ( .A(n19244), .B(n27716), .Z(n19245) );
  NANDN U23621 ( .A(n27719), .B(n19245), .Z(n19246) );
  AND U23622 ( .A(n27720), .B(n19246), .Z(n19247) );
  OR U23623 ( .A(n27722), .B(n19247), .Z(n19250) );
  NANDN U23624 ( .A(x[3613]), .B(y[3613]), .Z(n19249) );
  ANDN U23625 ( .B(n19249), .A(n19248), .Z(n27724) );
  NAND U23626 ( .A(n19250), .B(n27724), .Z(n19251) );
  NANDN U23627 ( .A(n27727), .B(n19251), .Z(n19254) );
  NANDN U23628 ( .A(x[3615]), .B(y[3615]), .Z(n19253) );
  ANDN U23629 ( .B(n19253), .A(n19252), .Z(n27728) );
  NAND U23630 ( .A(n19254), .B(n27728), .Z(n19255) );
  AND U23631 ( .A(n27730), .B(n19255), .Z(n19256) );
  OR U23632 ( .A(n27732), .B(n19256), .Z(n19259) );
  NOR U23633 ( .A(n19258), .B(n19257), .Z(n27734) );
  NAND U23634 ( .A(n19259), .B(n27734), .Z(n19260) );
  NAND U23635 ( .A(n19260), .B(n27737), .Z(n19262) );
  NANDN U23636 ( .A(n19262), .B(n19261), .Z(n19263) );
  NANDN U23637 ( .A(n27741), .B(n19263), .Z(n19266) );
  OR U23638 ( .A(n19265), .B(n19264), .Z(n27743) );
  ANDN U23639 ( .B(n19266), .A(n27743), .Z(n19269) );
  ANDN U23640 ( .B(n19268), .A(n19267), .Z(n27744) );
  NANDN U23641 ( .A(n19269), .B(n27744), .Z(n19272) );
  NANDN U23642 ( .A(x[3623]), .B(y[3623]), .Z(n19271) );
  ANDN U23643 ( .B(n19271), .A(n19270), .Z(n27746) );
  NAND U23644 ( .A(n19272), .B(n27746), .Z(n19273) );
  NANDN U23645 ( .A(n27749), .B(n19273), .Z(n19274) );
  NANDN U23646 ( .A(n27750), .B(n19274), .Z(n19275) );
  AND U23647 ( .A(n27752), .B(n19275), .Z(n19276) );
  OR U23648 ( .A(n19277), .B(n19276), .Z(n19280) );
  NANDN U23649 ( .A(y[3628]), .B(x[3628]), .Z(n19279) );
  ANDN U23650 ( .B(n19279), .A(n19278), .Z(n27758) );
  NAND U23651 ( .A(n19280), .B(n27758), .Z(n19283) );
  NOR U23652 ( .A(n19282), .B(n19281), .Z(n27761) );
  NAND U23653 ( .A(n19283), .B(n27761), .Z(n19286) );
  NOR U23654 ( .A(n19285), .B(n19284), .Z(n27762) );
  NAND U23655 ( .A(n19286), .B(n27762), .Z(n19287) );
  NAND U23656 ( .A(n19288), .B(n19287), .Z(n19289) );
  NANDN U23657 ( .A(n19289), .B(n20223), .Z(n19290) );
  AND U23658 ( .A(n27766), .B(n19290), .Z(n19293) );
  NOR U23659 ( .A(n19292), .B(n19291), .Z(n27768) );
  NANDN U23660 ( .A(n19293), .B(n27768), .Z(n19296) );
  NOR U23661 ( .A(n19295), .B(n19294), .Z(n27770) );
  NAND U23662 ( .A(n19296), .B(n27770), .Z(n19299) );
  NOR U23663 ( .A(n19298), .B(n19297), .Z(n27772) );
  NAND U23664 ( .A(n19299), .B(n27772), .Z(n19300) );
  NANDN U23665 ( .A(n27774), .B(n19300), .Z(n19301) );
  AND U23666 ( .A(n27776), .B(n19301), .Z(n19302) );
  OR U23667 ( .A(n27779), .B(n19302), .Z(n19305) );
  NANDN U23668 ( .A(x[3639]), .B(y[3639]), .Z(n19304) );
  ANDN U23669 ( .B(n19304), .A(n19303), .Z(n27780) );
  NAND U23670 ( .A(n19305), .B(n27780), .Z(n19306) );
  NANDN U23671 ( .A(n27783), .B(n19306), .Z(n19307) );
  NANDN U23672 ( .A(n27784), .B(n19307), .Z(n19308) );
  AND U23673 ( .A(n27786), .B(n19308), .Z(n19311) );
  AND U23674 ( .A(n19309), .B(n27789), .Z(n19310) );
  NANDN U23675 ( .A(n19311), .B(n19310), .Z(n19312) );
  NANDN U23676 ( .A(n27793), .B(n19312), .Z(n19315) );
  OR U23677 ( .A(n19314), .B(n19313), .Z(n27795) );
  ANDN U23678 ( .B(n19315), .A(n27795), .Z(n19318) );
  ANDN U23679 ( .B(n19317), .A(n19316), .Z(n27796) );
  NANDN U23680 ( .A(n19318), .B(n27796), .Z(n19321) );
  NANDN U23681 ( .A(x[3647]), .B(y[3647]), .Z(n19320) );
  ANDN U23682 ( .B(n19320), .A(n19319), .Z(n27798) );
  NAND U23683 ( .A(n19321), .B(n27798), .Z(n19322) );
  NANDN U23684 ( .A(n27801), .B(n19322), .Z(n19323) );
  NANDN U23685 ( .A(n27802), .B(n19323), .Z(n19324) );
  AND U23686 ( .A(n27804), .B(n19324), .Z(n19325) );
  ANDN U23687 ( .B(n27807), .A(n19325), .Z(n19327) );
  NAND U23688 ( .A(n19327), .B(n19326), .Z(n19328) );
  AND U23689 ( .A(n27810), .B(n19328), .Z(n19329) );
  ANDN U23690 ( .B(n27814), .A(n19329), .Z(n19330) );
  NAND U23691 ( .A(n19331), .B(n19330), .Z(n19334) );
  NANDN U23692 ( .A(y[3654]), .B(x[3654]), .Z(n19333) );
  ANDN U23693 ( .B(n19333), .A(n19332), .Z(n27816) );
  NAND U23694 ( .A(n19334), .B(n27816), .Z(n19337) );
  NANDN U23695 ( .A(n19336), .B(n19335), .Z(n27818) );
  ANDN U23696 ( .B(n19337), .A(n27818), .Z(n19338) );
  OR U23697 ( .A(n27821), .B(n19338), .Z(n19339) );
  AND U23698 ( .A(n27823), .B(n19339), .Z(n19340) );
  NAND U23699 ( .A(n19341), .B(n19340), .Z(n19342) );
  NANDN U23700 ( .A(n27827), .B(n19342), .Z(n19343) );
  NANDN U23701 ( .A(n27829), .B(n19343), .Z(n19344) );
  ANDN U23702 ( .B(n19344), .A(n27830), .Z(n19345) );
  OR U23703 ( .A(n27833), .B(n19345), .Z(n19346) );
  NANDN U23704 ( .A(n27835), .B(n19346), .Z(n19347) );
  NAND U23705 ( .A(n19347), .B(n27838), .Z(n19350) );
  XOR U23706 ( .A(n19348), .B(y[3664]), .Z(n19349) );
  NANDN U23707 ( .A(n19350), .B(n19349), .Z(n19351) );
  NANDN U23708 ( .A(n27841), .B(n19351), .Z(n19354) );
  NANDN U23709 ( .A(x[3665]), .B(y[3665]), .Z(n19352) );
  NAND U23710 ( .A(n19353), .B(n19352), .Z(n27842) );
  ANDN U23711 ( .B(n19354), .A(n27842), .Z(n19355) );
  OR U23712 ( .A(n27845), .B(n19355), .Z(n19356) );
  NANDN U23713 ( .A(n27847), .B(n19356), .Z(n19359) );
  ANDN U23714 ( .B(n19358), .A(n19357), .Z(n27848) );
  NAND U23715 ( .A(n19359), .B(n27848), .Z(n19360) );
  NANDN U23716 ( .A(n27851), .B(n19360), .Z(n19363) );
  NANDN U23717 ( .A(y[3670]), .B(x[3670]), .Z(n19361) );
  NAND U23718 ( .A(n19362), .B(n19361), .Z(n27852) );
  ANDN U23719 ( .B(n19363), .A(n27852), .Z(n19364) );
  OR U23720 ( .A(n27855), .B(n19364), .Z(n19365) );
  NANDN U23721 ( .A(n27857), .B(n19365), .Z(n19366) );
  NANDN U23722 ( .A(n27859), .B(n19366), .Z(n19369) );
  NANDN U23723 ( .A(y[3674]), .B(x[3674]), .Z(n19368) );
  ANDN U23724 ( .B(n19368), .A(n19367), .Z(n27860) );
  NAND U23725 ( .A(n19369), .B(n27860), .Z(n19373) );
  NAND U23726 ( .A(n19370), .B(y[3676]), .Z(n19371) );
  NANDN U23727 ( .A(n19372), .B(n19371), .Z(n27862) );
  ANDN U23728 ( .B(n19373), .A(n27862), .Z(n19376) );
  NANDN U23729 ( .A(y[3676]), .B(x[3676]), .Z(n19375) );
  ANDN U23730 ( .B(n19375), .A(n19374), .Z(n27864) );
  NANDN U23731 ( .A(n19376), .B(n27864), .Z(n19377) );
  NANDN U23732 ( .A(n27867), .B(n19377), .Z(n19380) );
  NANDN U23733 ( .A(y[3678]), .B(x[3678]), .Z(n19379) );
  ANDN U23734 ( .B(n19379), .A(n19378), .Z(n27868) );
  NAND U23735 ( .A(n19380), .B(n27868), .Z(n19381) );
  NANDN U23736 ( .A(n27871), .B(n19381), .Z(n19384) );
  NANDN U23737 ( .A(y[3680]), .B(x[3680]), .Z(n19382) );
  NAND U23738 ( .A(n19383), .B(n19382), .Z(n27872) );
  ANDN U23739 ( .B(n19384), .A(n27872), .Z(n19385) );
  OR U23740 ( .A(n27875), .B(n19385), .Z(n19386) );
  NANDN U23741 ( .A(n27877), .B(n19386), .Z(n19387) );
  NANDN U23742 ( .A(n27879), .B(n19387), .Z(n19390) );
  NANDN U23743 ( .A(y[3684]), .B(x[3684]), .Z(n19389) );
  ANDN U23744 ( .B(n19389), .A(n19388), .Z(n27880) );
  NAND U23745 ( .A(n19390), .B(n27880), .Z(n19394) );
  NAND U23746 ( .A(n19391), .B(y[3686]), .Z(n19392) );
  NANDN U23747 ( .A(n19393), .B(n19392), .Z(n27882) );
  ANDN U23748 ( .B(n19394), .A(n27882), .Z(n19397) );
  NANDN U23749 ( .A(y[3686]), .B(x[3686]), .Z(n19396) );
  ANDN U23750 ( .B(n19396), .A(n19395), .Z(n27884) );
  NANDN U23751 ( .A(n19397), .B(n27884), .Z(n19398) );
  NANDN U23752 ( .A(n27887), .B(n19398), .Z(n19401) );
  NANDN U23753 ( .A(y[3688]), .B(x[3688]), .Z(n19400) );
  ANDN U23754 ( .B(n19400), .A(n19399), .Z(n27888) );
  NAND U23755 ( .A(n19401), .B(n27888), .Z(n19402) );
  NANDN U23756 ( .A(n27891), .B(n19402), .Z(n19405) );
  NANDN U23757 ( .A(y[3690]), .B(x[3690]), .Z(n19403) );
  NAND U23758 ( .A(n19404), .B(n19403), .Z(n27892) );
  ANDN U23759 ( .B(n19405), .A(n27892), .Z(n19406) );
  OR U23760 ( .A(n27895), .B(n19406), .Z(n19407) );
  NANDN U23761 ( .A(n27897), .B(n19407), .Z(n19408) );
  NANDN U23762 ( .A(n27899), .B(n19408), .Z(n19411) );
  NANDN U23763 ( .A(y[3694]), .B(x[3694]), .Z(n19410) );
  ANDN U23764 ( .B(n19410), .A(n19409), .Z(n27900) );
  NAND U23765 ( .A(n19411), .B(n27900), .Z(n19412) );
  NANDN U23766 ( .A(n27902), .B(n19412), .Z(n19415) );
  NANDN U23767 ( .A(y[3696]), .B(x[3696]), .Z(n19414) );
  ANDN U23768 ( .B(n19414), .A(n19413), .Z(n27904) );
  NAND U23769 ( .A(n19415), .B(n27904), .Z(n19416) );
  NANDN U23770 ( .A(n27907), .B(n19416), .Z(n19417) );
  AND U23771 ( .A(n27908), .B(n19417), .Z(n19420) );
  NOR U23772 ( .A(n27913), .B(n19418), .Z(n19419) );
  NANDN U23773 ( .A(n19420), .B(n19419), .Z(n19423) );
  NANDN U23774 ( .A(y[3700]), .B(x[3700]), .Z(n19422) );
  ANDN U23775 ( .B(n19422), .A(n19421), .Z(n27914) );
  NAND U23776 ( .A(n19423), .B(n27914), .Z(n19427) );
  NAND U23777 ( .A(n19424), .B(y[3702]), .Z(n19425) );
  NANDN U23778 ( .A(n19426), .B(n19425), .Z(n27917) );
  ANDN U23779 ( .B(n19427), .A(n27917), .Z(n19430) );
  NANDN U23780 ( .A(y[3702]), .B(x[3702]), .Z(n19429) );
  ANDN U23781 ( .B(n19429), .A(n19428), .Z(n27918) );
  NANDN U23782 ( .A(n19430), .B(n27918), .Z(n19433) );
  NANDN U23783 ( .A(x[3704]), .B(y[3704]), .Z(n19432) );
  ANDN U23784 ( .B(n19432), .A(n19431), .Z(n27920) );
  NAND U23785 ( .A(n19433), .B(n27920), .Z(n19436) );
  NANDN U23786 ( .A(y[3704]), .B(x[3704]), .Z(n19435) );
  ANDN U23787 ( .B(n19435), .A(n19434), .Z(n27922) );
  NAND U23788 ( .A(n19436), .B(n27922), .Z(n19440) );
  NAND U23789 ( .A(n19437), .B(y[3706]), .Z(n19438) );
  NANDN U23790 ( .A(n19439), .B(n19438), .Z(n27924) );
  ANDN U23791 ( .B(n19440), .A(n27924), .Z(n19443) );
  NANDN U23792 ( .A(y[3706]), .B(x[3706]), .Z(n19442) );
  ANDN U23793 ( .B(n19442), .A(n19441), .Z(n27926) );
  NANDN U23794 ( .A(n19443), .B(n27926), .Z(n19447) );
  NAND U23795 ( .A(n19444), .B(y[3708]), .Z(n19445) );
  NANDN U23796 ( .A(n19446), .B(n19445), .Z(n27929) );
  ANDN U23797 ( .B(n19447), .A(n27929), .Z(n19448) );
  OR U23798 ( .A(n27931), .B(n19448), .Z(n19451) );
  NOR U23799 ( .A(n19450), .B(n19449), .Z(n27932) );
  NAND U23800 ( .A(n19451), .B(n27932), .Z(n19454) );
  NOR U23801 ( .A(n19453), .B(n19452), .Z(n27935) );
  NAND U23802 ( .A(n19454), .B(n27935), .Z(n19455) );
  AND U23803 ( .A(n19456), .B(n19455), .Z(n19459) );
  NANDN U23804 ( .A(y[3712]), .B(x[3712]), .Z(n19458) );
  ANDN U23805 ( .B(n19458), .A(n19457), .Z(n27940) );
  NANDN U23806 ( .A(n19459), .B(n27940), .Z(n19463) );
  NAND U23807 ( .A(n19460), .B(y[3714]), .Z(n19461) );
  NANDN U23808 ( .A(n19462), .B(n19461), .Z(n27942) );
  ANDN U23809 ( .B(n19463), .A(n27942), .Z(n19466) );
  NANDN U23810 ( .A(y[3714]), .B(x[3714]), .Z(n19465) );
  ANDN U23811 ( .B(n19465), .A(n19464), .Z(n27944) );
  NANDN U23812 ( .A(n19466), .B(n27944), .Z(n19467) );
  NANDN U23813 ( .A(n27947), .B(n19467), .Z(n19468) );
  NANDN U23814 ( .A(n27949), .B(n19468), .Z(n19469) );
  AND U23815 ( .A(n27950), .B(n19469), .Z(n19472) );
  NOR U23816 ( .A(n19471), .B(n19470), .Z(n27953) );
  NANDN U23817 ( .A(n19472), .B(n27953), .Z(n19473) );
  AND U23818 ( .A(n19474), .B(n19473), .Z(n19477) );
  NANDN U23819 ( .A(y[3720]), .B(x[3720]), .Z(n19476) );
  ANDN U23820 ( .B(n19476), .A(n19475), .Z(n27958) );
  NANDN U23821 ( .A(n19477), .B(n27958), .Z(n19478) );
  NANDN U23822 ( .A(n27960), .B(n19478), .Z(n19479) );
  NANDN U23823 ( .A(n27963), .B(n19479), .Z(n19482) );
  OR U23824 ( .A(n19481), .B(n19480), .Z(n27965) );
  ANDN U23825 ( .B(n19482), .A(n27965), .Z(n19485) );
  NOR U23826 ( .A(n19484), .B(n19483), .Z(n27966) );
  NANDN U23827 ( .A(n19485), .B(n27966), .Z(n19486) );
  AND U23828 ( .A(n19487), .B(n19486), .Z(n19490) );
  NANDN U23829 ( .A(y[3726]), .B(x[3726]), .Z(n19489) );
  ANDN U23830 ( .B(n19489), .A(n19488), .Z(n27972) );
  NANDN U23831 ( .A(n19490), .B(n27972), .Z(n19491) );
  NANDN U23832 ( .A(n19492), .B(n19491), .Z(n19493) );
  AND U23833 ( .A(n27978), .B(n19493), .Z(n19494) );
  OR U23834 ( .A(n27980), .B(n19494), .Z(n19497) );
  NANDN U23835 ( .A(y[3730]), .B(x[3730]), .Z(n19496) );
  ANDN U23836 ( .B(n19496), .A(n19495), .Z(n27982) );
  NAND U23837 ( .A(n19497), .B(n27982), .Z(n19498) );
  NANDN U23838 ( .A(n27985), .B(n19498), .Z(n19499) );
  AND U23839 ( .A(n27986), .B(n19499), .Z(n19500) );
  OR U23840 ( .A(n27989), .B(n19500), .Z(n19503) );
  NANDN U23841 ( .A(y[3734]), .B(x[3734]), .Z(n19501) );
  NAND U23842 ( .A(n19502), .B(n19501), .Z(n27990) );
  ANDN U23843 ( .B(n19503), .A(n27990), .Z(n19504) );
  OR U23844 ( .A(n27993), .B(n19504), .Z(n19505) );
  NANDN U23845 ( .A(n27995), .B(n19505), .Z(n19506) );
  NANDN U23846 ( .A(n27997), .B(n19506), .Z(n19509) );
  NANDN U23847 ( .A(n19508), .B(n19507), .Z(n27999) );
  ANDN U23848 ( .B(n19509), .A(n27999), .Z(n19512) );
  OR U23849 ( .A(n19510), .B(n20220), .Z(n19511) );
  OR U23850 ( .A(n19512), .B(n19511), .Z(n19513) );
  AND U23851 ( .A(n28002), .B(n19513), .Z(n19514) );
  OR U23852 ( .A(n28005), .B(n19514), .Z(n19517) );
  NANDN U23853 ( .A(y[3742]), .B(x[3742]), .Z(n19516) );
  ANDN U23854 ( .B(n19516), .A(n19515), .Z(n28006) );
  NAND U23855 ( .A(n19517), .B(n28006), .Z(n19518) );
  NANDN U23856 ( .A(n28009), .B(n19518), .Z(n19521) );
  NANDN U23857 ( .A(n19520), .B(n19519), .Z(n28010) );
  ANDN U23858 ( .B(n19521), .A(n28010), .Z(n19524) );
  OR U23859 ( .A(n19522), .B(n20219), .Z(n19523) );
  OR U23860 ( .A(n19524), .B(n19523), .Z(n19525) );
  AND U23861 ( .A(n28014), .B(n19525), .Z(n19526) );
  OR U23862 ( .A(n19527), .B(n19526), .Z(n19530) );
  NANDN U23863 ( .A(y[3748]), .B(x[3748]), .Z(n19529) );
  ANDN U23864 ( .B(n19529), .A(n19528), .Z(n28020) );
  NAND U23865 ( .A(n19530), .B(n28020), .Z(n19533) );
  NOR U23866 ( .A(n19532), .B(n19531), .Z(n28022) );
  NAND U23867 ( .A(n19533), .B(n28022), .Z(n19536) );
  OR U23868 ( .A(n19535), .B(n19534), .Z(n28025) );
  ANDN U23869 ( .B(n19536), .A(n28025), .Z(n19539) );
  NOR U23870 ( .A(n19538), .B(n19537), .Z(n28026) );
  NANDN U23871 ( .A(n19539), .B(n28026), .Z(n19540) );
  AND U23872 ( .A(n28028), .B(n19540), .Z(n19543) );
  NANDN U23873 ( .A(x[3753]), .B(y[3753]), .Z(n19542) );
  ANDN U23874 ( .B(n19542), .A(n19541), .Z(n28031) );
  NANDN U23875 ( .A(n19543), .B(n28031), .Z(n19546) );
  NANDN U23876 ( .A(y[3755]), .B(x[3755]), .Z(n19545) );
  ANDN U23877 ( .B(n19545), .A(n19544), .Z(n28032) );
  NAND U23878 ( .A(n19546), .B(n28032), .Z(n19549) );
  NANDN U23879 ( .A(x[3755]), .B(y[3755]), .Z(n19548) );
  ANDN U23880 ( .B(n19548), .A(n19547), .Z(n28034) );
  NAND U23881 ( .A(n19549), .B(n28034), .Z(n19550) );
  AND U23882 ( .A(n28036), .B(n19550), .Z(n19553) );
  NANDN U23883 ( .A(x[3757]), .B(y[3757]), .Z(n19552) );
  ANDN U23884 ( .B(n19552), .A(n19551), .Z(n28038) );
  NANDN U23885 ( .A(n19553), .B(n28038), .Z(n19554) );
  NANDN U23886 ( .A(n28040), .B(n19554), .Z(n19555) );
  AND U23887 ( .A(n28042), .B(n19555), .Z(n19556) );
  OR U23888 ( .A(n28045), .B(n19556), .Z(n19559) );
  NANDN U23889 ( .A(x[3761]), .B(y[3761]), .Z(n19558) );
  ANDN U23890 ( .B(n19558), .A(n19557), .Z(n28046) );
  NAND U23891 ( .A(n19559), .B(n28046), .Z(n19560) );
  NANDN U23892 ( .A(n28049), .B(n19560), .Z(n19561) );
  NAND U23893 ( .A(n19562), .B(n19561), .Z(n19563) );
  NANDN U23894 ( .A(n28053), .B(n19563), .Z(n19566) );
  OR U23895 ( .A(n19565), .B(n19564), .Z(n28055) );
  ANDN U23896 ( .B(n19566), .A(n28055), .Z(n19569) );
  ANDN U23897 ( .B(n19568), .A(n19567), .Z(n28056) );
  NANDN U23898 ( .A(n19569), .B(n28056), .Z(n19572) );
  NANDN U23899 ( .A(x[3767]), .B(y[3767]), .Z(n19571) );
  ANDN U23900 ( .B(n19571), .A(n19570), .Z(n28058) );
  NAND U23901 ( .A(n19572), .B(n28058), .Z(n19573) );
  NANDN U23902 ( .A(n28060), .B(n19573), .Z(n19574) );
  AND U23903 ( .A(n28062), .B(n19574), .Z(n19577) );
  NOR U23904 ( .A(n19576), .B(n19575), .Z(n28064) );
  NANDN U23905 ( .A(n19577), .B(n28064), .Z(n19578) );
  AND U23906 ( .A(n19579), .B(n19578), .Z(n19582) );
  NANDN U23907 ( .A(y[3772]), .B(x[3772]), .Z(n19581) );
  ANDN U23908 ( .B(n19581), .A(n19580), .Z(n28070) );
  NANDN U23909 ( .A(n19582), .B(n28070), .Z(n19583) );
  NANDN U23910 ( .A(n28072), .B(n19583), .Z(n19584) );
  NANDN U23911 ( .A(n28075), .B(n19584), .Z(n19587) );
  OR U23912 ( .A(n19586), .B(n19585), .Z(n28077) );
  ANDN U23913 ( .B(n19587), .A(n28077), .Z(n19590) );
  NOR U23914 ( .A(n19589), .B(n19588), .Z(n28078) );
  NANDN U23915 ( .A(n19590), .B(n28078), .Z(n19591) );
  AND U23916 ( .A(n19592), .B(n19591), .Z(n19595) );
  NANDN U23917 ( .A(y[3778]), .B(x[3778]), .Z(n19594) );
  ANDN U23918 ( .B(n19594), .A(n19593), .Z(n28084) );
  NANDN U23919 ( .A(n19595), .B(n28084), .Z(n19596) );
  NANDN U23920 ( .A(n28087), .B(n19596), .Z(n19599) );
  NANDN U23921 ( .A(y[3780]), .B(x[3780]), .Z(n19598) );
  ANDN U23922 ( .B(n19598), .A(n19597), .Z(n28088) );
  NAND U23923 ( .A(n19599), .B(n28088), .Z(n19600) );
  AND U23924 ( .A(n28090), .B(n19600), .Z(n19603) );
  NANDN U23925 ( .A(y[3782]), .B(x[3782]), .Z(n19602) );
  ANDN U23926 ( .B(n19602), .A(n19601), .Z(n28092) );
  NANDN U23927 ( .A(n19603), .B(n28092), .Z(n19607) );
  NAND U23928 ( .A(n19604), .B(y[3784]), .Z(n19605) );
  NANDN U23929 ( .A(n19606), .B(n19605), .Z(n28094) );
  ANDN U23930 ( .B(n19607), .A(n28094), .Z(n19610) );
  NANDN U23931 ( .A(y[3784]), .B(x[3784]), .Z(n19609) );
  ANDN U23932 ( .B(n19609), .A(n19608), .Z(n28096) );
  NANDN U23933 ( .A(n19610), .B(n28096), .Z(n19611) );
  NANDN U23934 ( .A(n28099), .B(n19611), .Z(n19614) );
  NANDN U23935 ( .A(y[3786]), .B(x[3786]), .Z(n19613) );
  ANDN U23936 ( .B(n19613), .A(n19612), .Z(n28100) );
  NAND U23937 ( .A(n19614), .B(n28100), .Z(n19615) );
  AND U23938 ( .A(n28102), .B(n19615), .Z(n19618) );
  NANDN U23939 ( .A(y[3788]), .B(x[3788]), .Z(n19616) );
  NAND U23940 ( .A(n19617), .B(n19616), .Z(n28104) );
  OR U23941 ( .A(n19618), .B(n28104), .Z(n19619) );
  NANDN U23942 ( .A(n28107), .B(n19619), .Z(n19622) );
  NANDN U23943 ( .A(y[3790]), .B(x[3790]), .Z(n19620) );
  NANDN U23944 ( .A(n19621), .B(n19620), .Z(n28109) );
  ANDN U23945 ( .B(n19622), .A(n28109), .Z(n19623) );
  OR U23946 ( .A(n28111), .B(n19623), .Z(n19624) );
  NANDN U23947 ( .A(n28113), .B(n19624), .Z(n19625) );
  NANDN U23948 ( .A(n19626), .B(n19625), .Z(n19627) );
  AND U23949 ( .A(n28116), .B(n19627), .Z(n19628) );
  ANDN U23950 ( .B(n28119), .A(n19628), .Z(n19630) );
  AND U23951 ( .A(n19630), .B(n19629), .Z(n19633) );
  NANDN U23952 ( .A(y[3796]), .B(x[3796]), .Z(n19632) );
  ANDN U23953 ( .B(n19632), .A(n19631), .Z(n28122) );
  NANDN U23954 ( .A(n19633), .B(n28122), .Z(n19634) );
  NANDN U23955 ( .A(n28125), .B(n19634), .Z(n19637) );
  NANDN U23956 ( .A(y[3798]), .B(x[3798]), .Z(n19636) );
  ANDN U23957 ( .B(n19636), .A(n19635), .Z(n28126) );
  NAND U23958 ( .A(n19637), .B(n28126), .Z(n19638) );
  AND U23959 ( .A(n28128), .B(n19638), .Z(n19641) );
  NANDN U23960 ( .A(y[3800]), .B(x[3800]), .Z(n19640) );
  ANDN U23961 ( .B(n19640), .A(n19639), .Z(n28130) );
  NANDN U23962 ( .A(n19641), .B(n28130), .Z(n19642) );
  NANDN U23963 ( .A(n28132), .B(n19642), .Z(n19643) );
  AND U23964 ( .A(n28134), .B(n19643), .Z(n19644) );
  OR U23965 ( .A(n28137), .B(n19644), .Z(n19647) );
  NANDN U23966 ( .A(y[3804]), .B(x[3804]), .Z(n19646) );
  ANDN U23967 ( .B(n19646), .A(n19645), .Z(n28138) );
  NAND U23968 ( .A(n19647), .B(n28138), .Z(n19648) );
  NANDN U23969 ( .A(n28141), .B(n19648), .Z(n19651) );
  NANDN U23970 ( .A(y[3806]), .B(x[3806]), .Z(n19650) );
  NANDN U23971 ( .A(y[3807]), .B(x[3807]), .Z(n19649) );
  NAND U23972 ( .A(n19650), .B(n19649), .Z(n28142) );
  ANDN U23973 ( .B(n19651), .A(n28142), .Z(n19652) );
  OR U23974 ( .A(n28144), .B(n19652), .Z(n19653) );
  NAND U23975 ( .A(n19653), .B(n28147), .Z(n19654) );
  NAND U23976 ( .A(n19654), .B(n28148), .Z(n19655) );
  ANDN U23977 ( .B(n19655), .A(n28150), .Z(n19656) );
  OR U23978 ( .A(n28153), .B(n19656), .Z(n19659) );
  OR U23979 ( .A(n19658), .B(n19657), .Z(n28155) );
  ANDN U23980 ( .B(n19659), .A(n28155), .Z(n19660) );
  OR U23981 ( .A(n19661), .B(n19660), .Z(n19664) );
  NANDN U23982 ( .A(y[3814]), .B(x[3814]), .Z(n19663) );
  ANDN U23983 ( .B(n19663), .A(n19662), .Z(n28160) );
  NAND U23984 ( .A(n19664), .B(n28160), .Z(n19665) );
  NANDN U23985 ( .A(n28162), .B(n19665), .Z(n19666) );
  AND U23986 ( .A(n28164), .B(n19666), .Z(n19669) );
  OR U23987 ( .A(n19668), .B(n19667), .Z(n28167) );
  OR U23988 ( .A(n19669), .B(n28167), .Z(n19672) );
  NOR U23989 ( .A(n19671), .B(n19670), .Z(n28168) );
  NAND U23990 ( .A(n19672), .B(n28168), .Z(n19673) );
  AND U23991 ( .A(n28172), .B(n19673), .Z(n19674) );
  NANDN U23992 ( .A(n19675), .B(n19674), .Z(n19676) );
  NANDN U23993 ( .A(n28175), .B(n19676), .Z(n19677) );
  AND U23994 ( .A(n19678), .B(n19677), .Z(n19679) );
  OR U23995 ( .A(n28181), .B(n19679), .Z(n19682) );
  ANDN U23996 ( .B(n28183), .A(n19680), .Z(n19681) );
  NAND U23997 ( .A(n19682), .B(n19681), .Z(n19683) );
  NANDN U23998 ( .A(n28187), .B(n19683), .Z(n19684) );
  NANDN U23999 ( .A(n28188), .B(n19684), .Z(n19685) );
  NANDN U24000 ( .A(n28191), .B(n19685), .Z(n19686) );
  AND U24001 ( .A(n19687), .B(n19686), .Z(n19688) );
  OR U24002 ( .A(n28195), .B(n19688), .Z(n19689) );
  NANDN U24003 ( .A(n28197), .B(n19689), .Z(n19690) );
  NANDN U24004 ( .A(n28199), .B(n19690), .Z(n19691) );
  NAND U24005 ( .A(n19692), .B(n19691), .Z(n19693) );
  NANDN U24006 ( .A(n28205), .B(n19693), .Z(n19696) );
  OR U24007 ( .A(n19695), .B(n19694), .Z(n28207) );
  ANDN U24008 ( .B(n19696), .A(n28207), .Z(n19699) );
  ANDN U24009 ( .B(n19698), .A(n19697), .Z(n28208) );
  NANDN U24010 ( .A(n19699), .B(n28208), .Z(n19702) );
  NANDN U24011 ( .A(x[3835]), .B(y[3835]), .Z(n19701) );
  ANDN U24012 ( .B(n19701), .A(n19700), .Z(n28210) );
  NAND U24013 ( .A(n19702), .B(n28210), .Z(n19703) );
  NANDN U24014 ( .A(n28213), .B(n19703), .Z(n19706) );
  OR U24015 ( .A(n19705), .B(n19704), .Z(n28214) );
  ANDN U24016 ( .B(n19706), .A(n28214), .Z(n19709) );
  ANDN U24017 ( .B(n19708), .A(n19707), .Z(n28216) );
  NANDN U24018 ( .A(n19709), .B(n28216), .Z(n19713) );
  NAND U24019 ( .A(n19710), .B(y[3840]), .Z(n19711) );
  NANDN U24020 ( .A(n19712), .B(n19711), .Z(n28219) );
  ANDN U24021 ( .B(n19713), .A(n28219), .Z(n19716) );
  NANDN U24022 ( .A(y[3840]), .B(x[3840]), .Z(n19715) );
  ANDN U24023 ( .B(n19715), .A(n19714), .Z(n28220) );
  NANDN U24024 ( .A(n19716), .B(n28220), .Z(n19717) );
  NANDN U24025 ( .A(n28222), .B(n19717), .Z(n19718) );
  NANDN U24026 ( .A(n28224), .B(n19718), .Z(n19719) );
  NAND U24027 ( .A(n19719), .B(n28226), .Z(n19720) );
  ANDN U24028 ( .B(n19720), .A(n28228), .Z(n19721) );
  OR U24029 ( .A(n28231), .B(n19721), .Z(n19724) );
  NANDN U24030 ( .A(n19723), .B(n19722), .Z(n28233) );
  ANDN U24031 ( .B(n19724), .A(n28233), .Z(n19725) );
  OR U24032 ( .A(n28235), .B(n19725), .Z(n19726) );
  NANDN U24033 ( .A(n28236), .B(n19726), .Z(n19727) );
  NANDN U24034 ( .A(n28238), .B(n19727), .Z(n19728) );
  AND U24035 ( .A(n28240), .B(n19728), .Z(n19731) );
  NANDN U24036 ( .A(n19729), .B(n28244), .Z(n19730) );
  OR U24037 ( .A(n19731), .B(n19730), .Z(n19732) );
  AND U24038 ( .A(n28246), .B(n19732), .Z(n19733) );
  OR U24039 ( .A(n28248), .B(n19733), .Z(n19736) );
  NANDN U24040 ( .A(y[3854]), .B(x[3854]), .Z(n19735) );
  ANDN U24041 ( .B(n19735), .A(n19734), .Z(n28250) );
  NAND U24042 ( .A(n19736), .B(n28250), .Z(n19737) );
  NANDN U24043 ( .A(n28253), .B(n19737), .Z(n19738) );
  AND U24044 ( .A(n28254), .B(n19738), .Z(n19739) );
  OR U24045 ( .A(n28256), .B(n19739), .Z(n19740) );
  AND U24046 ( .A(n28258), .B(n19740), .Z(n19741) );
  OR U24047 ( .A(n28261), .B(n19741), .Z(n19744) );
  NOR U24048 ( .A(n19743), .B(n19742), .Z(n28262) );
  NAND U24049 ( .A(n19744), .B(n28262), .Z(n19745) );
  NANDN U24050 ( .A(n19746), .B(n19745), .Z(n19747) );
  AND U24051 ( .A(n28268), .B(n19747), .Z(n19748) );
  OR U24052 ( .A(n28270), .B(n19748), .Z(n19749) );
  AND U24053 ( .A(n28272), .B(n19749), .Z(n19750) );
  OR U24054 ( .A(n28275), .B(n19750), .Z(n19753) );
  NANDN U24055 ( .A(y[3866]), .B(x[3866]), .Z(n19752) );
  ANDN U24056 ( .B(n19752), .A(n19751), .Z(n28276) );
  NAND U24057 ( .A(n19753), .B(n28276), .Z(n19754) );
  NANDN U24058 ( .A(n28278), .B(n19754), .Z(n19755) );
  AND U24059 ( .A(n28280), .B(n19755), .Z(n19758) );
  NANDN U24060 ( .A(x[3870]), .B(y[3870]), .Z(n19756) );
  NANDN U24061 ( .A(n19757), .B(n19756), .Z(n28282) );
  OR U24062 ( .A(n19758), .B(n28282), .Z(n19761) );
  NANDN U24063 ( .A(y[3870]), .B(x[3870]), .Z(n19760) );
  ANDN U24064 ( .B(n19760), .A(n19759), .Z(n28284) );
  NAND U24065 ( .A(n19761), .B(n28284), .Z(n19765) );
  NAND U24066 ( .A(n19762), .B(y[3872]), .Z(n19763) );
  NANDN U24067 ( .A(n19764), .B(n19763), .Z(n28287) );
  ANDN U24068 ( .B(n19765), .A(n28287), .Z(n19768) );
  NANDN U24069 ( .A(y[3872]), .B(x[3872]), .Z(n19767) );
  ANDN U24070 ( .B(n19767), .A(n19766), .Z(n28288) );
  NANDN U24071 ( .A(n19768), .B(n28288), .Z(n19769) );
  NANDN U24072 ( .A(n28290), .B(n19769), .Z(n19772) );
  NANDN U24073 ( .A(y[3874]), .B(x[3874]), .Z(n19771) );
  ANDN U24074 ( .B(n19771), .A(n19770), .Z(n28292) );
  NAND U24075 ( .A(n19772), .B(n28292), .Z(n19773) );
  AND U24076 ( .A(n28294), .B(n19773), .Z(n19776) );
  NANDN U24077 ( .A(y[3876]), .B(x[3876]), .Z(n19775) );
  ANDN U24078 ( .B(n19775), .A(n19774), .Z(n28297) );
  NANDN U24079 ( .A(n19776), .B(n28297), .Z(n19777) );
  AND U24080 ( .A(n28298), .B(n19777), .Z(n19780) );
  NANDN U24081 ( .A(y[3878]), .B(x[3878]), .Z(n19779) );
  ANDN U24082 ( .B(n19779), .A(n19778), .Z(n28300) );
  NANDN U24083 ( .A(n19780), .B(n28300), .Z(n19783) );
  NANDN U24084 ( .A(x[3880]), .B(y[3880]), .Z(n19782) );
  ANDN U24085 ( .B(n19782), .A(n19781), .Z(n28302) );
  NAND U24086 ( .A(n19783), .B(n28302), .Z(n19786) );
  NANDN U24087 ( .A(y[3880]), .B(x[3880]), .Z(n19785) );
  ANDN U24088 ( .B(n19785), .A(n19784), .Z(n28305) );
  NAND U24089 ( .A(n19786), .B(n28305), .Z(n19787) );
  AND U24090 ( .A(n28306), .B(n19787), .Z(n19790) );
  NANDN U24091 ( .A(y[3882]), .B(x[3882]), .Z(n19788) );
  NAND U24092 ( .A(n19789), .B(n19788), .Z(n28308) );
  OR U24093 ( .A(n19790), .B(n28308), .Z(n19791) );
  NANDN U24094 ( .A(n28311), .B(n19791), .Z(n19794) );
  NANDN U24095 ( .A(y[3884]), .B(x[3884]), .Z(n19792) );
  NAND U24096 ( .A(n19793), .B(n19792), .Z(n28313) );
  ANDN U24097 ( .B(n19794), .A(n28313), .Z(n19795) );
  OR U24098 ( .A(n28315), .B(n19795), .Z(n19796) );
  NANDN U24099 ( .A(n28316), .B(n19796), .Z(n19797) );
  NANDN U24100 ( .A(n28318), .B(n19797), .Z(n19798) );
  AND U24101 ( .A(n28320), .B(n19798), .Z(n19799) );
  OR U24102 ( .A(n28322), .B(n19799), .Z(n19800) );
  AND U24103 ( .A(n28324), .B(n19800), .Z(n19801) );
  OR U24104 ( .A(n19802), .B(n19801), .Z(n19805) );
  NANDN U24105 ( .A(y[3892]), .B(x[3892]), .Z(n19804) );
  ANDN U24106 ( .B(n19804), .A(n19803), .Z(n28330) );
  NAND U24107 ( .A(n19805), .B(n28330), .Z(n19806) );
  AND U24108 ( .A(n28333), .B(n19806), .Z(n19807) );
  OR U24109 ( .A(n28335), .B(n19807), .Z(n19810) );
  NOR U24110 ( .A(n20210), .B(n19808), .Z(n19809) );
  NAND U24111 ( .A(n19810), .B(n19809), .Z(n19811) );
  NANDN U24112 ( .A(n28339), .B(n19811), .Z(n19812) );
  AND U24113 ( .A(n19813), .B(n19812), .Z(n19814) );
  ANDN U24114 ( .B(n28344), .A(n19814), .Z(n19815) );
  OR U24115 ( .A(n19816), .B(n19815), .Z(n19819) );
  NANDN U24116 ( .A(y[3901]), .B(x[3901]), .Z(n19818) );
  NANDN U24117 ( .A(y[3900]), .B(x[3900]), .Z(n19817) );
  AND U24118 ( .A(n19818), .B(n19817), .Z(n28350) );
  NAND U24119 ( .A(n19819), .B(n28350), .Z(n19820) );
  NANDN U24120 ( .A(n28352), .B(n19820), .Z(n19823) );
  NOR U24121 ( .A(n19822), .B(n19821), .Z(n28354) );
  NAND U24122 ( .A(n19823), .B(n28354), .Z(n19824) );
  NANDN U24123 ( .A(n19825), .B(n19824), .Z(n19826) );
  AND U24124 ( .A(n28360), .B(n19826), .Z(n19827) );
  OR U24125 ( .A(n28362), .B(n19827), .Z(n19830) );
  NOR U24126 ( .A(n19829), .B(n19828), .Z(n28364) );
  NAND U24127 ( .A(n19830), .B(n28364), .Z(n19831) );
  NANDN U24128 ( .A(n19832), .B(n19831), .Z(n19833) );
  AND U24129 ( .A(n28368), .B(n19833), .Z(n19834) );
  ANDN U24130 ( .B(n28371), .A(n19834), .Z(n19836) );
  XNOR U24131 ( .A(x[3910]), .B(y[3910]), .Z(n19835) );
  AND U24132 ( .A(n19836), .B(n19835), .Z(n19837) );
  OR U24133 ( .A(n28375), .B(n19837), .Z(n19838) );
  NANDN U24134 ( .A(n28376), .B(n19838), .Z(n19841) );
  NOR U24135 ( .A(n19840), .B(n19839), .Z(n28378) );
  NAND U24136 ( .A(n19841), .B(n28378), .Z(n19842) );
  AND U24137 ( .A(n19843), .B(n19842), .Z(n19846) );
  NANDN U24138 ( .A(y[3914]), .B(x[3914]), .Z(n19845) );
  ANDN U24139 ( .B(n19845), .A(n19844), .Z(n28382) );
  NANDN U24140 ( .A(n19846), .B(n28382), .Z(n19850) );
  NAND U24141 ( .A(n19847), .B(y[3916]), .Z(n19848) );
  NANDN U24142 ( .A(n19849), .B(n19848), .Z(n28385) );
  ANDN U24143 ( .B(n19850), .A(n28385), .Z(n19851) );
  OR U24144 ( .A(n28387), .B(n19851), .Z(n19852) );
  NANDN U24145 ( .A(n28388), .B(n19852), .Z(n19855) );
  NOR U24146 ( .A(n19854), .B(n19853), .Z(n28390) );
  NAND U24147 ( .A(n19855), .B(n28390), .Z(n19856) );
  AND U24148 ( .A(n19857), .B(n19856), .Z(n19860) );
  NANDN U24149 ( .A(y[3920]), .B(x[3920]), .Z(n19859) );
  ANDN U24150 ( .B(n19859), .A(n19858), .Z(n28394) );
  NANDN U24151 ( .A(n19860), .B(n28394), .Z(n19864) );
  NAND U24152 ( .A(n19861), .B(y[3922]), .Z(n19862) );
  NANDN U24153 ( .A(n19863), .B(n19862), .Z(n28397) );
  ANDN U24154 ( .B(n19864), .A(n28397), .Z(n19867) );
  NANDN U24155 ( .A(y[3922]), .B(x[3922]), .Z(n19866) );
  ANDN U24156 ( .B(n19866), .A(n19865), .Z(n28398) );
  NANDN U24157 ( .A(n19867), .B(n28398), .Z(n19868) );
  NANDN U24158 ( .A(n28400), .B(n19868), .Z(n19869) );
  NANDN U24159 ( .A(n28402), .B(n19869), .Z(n19872) );
  OR U24160 ( .A(n19871), .B(n19870), .Z(n28404) );
  ANDN U24161 ( .B(n19872), .A(n28404), .Z(n19875) );
  NOR U24162 ( .A(n19874), .B(n19873), .Z(n28406) );
  NANDN U24163 ( .A(n19875), .B(n28406), .Z(n19876) );
  AND U24164 ( .A(n19877), .B(n19876), .Z(n19880) );
  NANDN U24165 ( .A(y[3928]), .B(x[3928]), .Z(n19879) );
  ANDN U24166 ( .B(n19879), .A(n19878), .Z(n28412) );
  NANDN U24167 ( .A(n19880), .B(n28412), .Z(n19881) );
  NANDN U24168 ( .A(n28414), .B(n19881), .Z(n19882) );
  NANDN U24169 ( .A(n28416), .B(n19882), .Z(n19883) );
  AND U24170 ( .A(n19884), .B(n19883), .Z(n19885) );
  OR U24171 ( .A(n28421), .B(n19885), .Z(n19888) );
  NANDN U24172 ( .A(n19887), .B(n19886), .Z(n28423) );
  ANDN U24173 ( .B(n19888), .A(n28423), .Z(n19889) );
  OR U24174 ( .A(n28425), .B(n19889), .Z(n19890) );
  NANDN U24175 ( .A(n28426), .B(n19890), .Z(n19891) );
  NANDN U24176 ( .A(n28428), .B(n19891), .Z(n19894) );
  NANDN U24177 ( .A(x[3937]), .B(y[3937]), .Z(n19892) );
  NAND U24178 ( .A(n19893), .B(n19892), .Z(n28430) );
  ANDN U24179 ( .B(n19894), .A(n28430), .Z(n19895) );
  OR U24180 ( .A(n28433), .B(n19895), .Z(n19898) );
  NANDN U24181 ( .A(x[3939]), .B(y[3939]), .Z(n19896) );
  NAND U24182 ( .A(n19897), .B(n19896), .Z(n28435) );
  ANDN U24183 ( .B(n19898), .A(n28435), .Z(n19899) );
  OR U24184 ( .A(n28437), .B(n19899), .Z(n19900) );
  NANDN U24185 ( .A(n28438), .B(n19900), .Z(n19901) );
  NANDN U24186 ( .A(n28441), .B(n19901), .Z(n19904) );
  NANDN U24187 ( .A(x[3943]), .B(y[3943]), .Z(n19902) );
  NANDN U24188 ( .A(n19903), .B(n19902), .Z(n28443) );
  ANDN U24189 ( .B(n19904), .A(n28443), .Z(n19905) );
  OR U24190 ( .A(n28445), .B(n19905), .Z(n19906) );
  AND U24191 ( .A(n19907), .B(n19906), .Z(n19908) );
  OR U24192 ( .A(n28451), .B(n19908), .Z(n19909) );
  NANDN U24193 ( .A(n28452), .B(n19909), .Z(n19912) );
  NOR U24194 ( .A(n19911), .B(n19910), .Z(n28454) );
  NAND U24195 ( .A(n19912), .B(n28454), .Z(n19913) );
  NAND U24196 ( .A(n19914), .B(n19913), .Z(n19918) );
  NAND U24197 ( .A(n19915), .B(x[3950]), .Z(n19917) );
  ANDN U24198 ( .B(n19917), .A(n19916), .Z(n28460) );
  NAND U24199 ( .A(n19918), .B(n28460), .Z(n19919) );
  AND U24200 ( .A(n19920), .B(n19919), .Z(n19921) );
  OR U24201 ( .A(n28466), .B(n19921), .Z(n19924) );
  NOR U24202 ( .A(n28470), .B(n19922), .Z(n19923) );
  NAND U24203 ( .A(n19924), .B(n19923), .Z(n19925) );
  NANDN U24204 ( .A(n28472), .B(n19925), .Z(n19928) );
  OR U24205 ( .A(n19927), .B(n19926), .Z(n28474) );
  ANDN U24206 ( .B(n19928), .A(n28474), .Z(n19929) );
  OR U24207 ( .A(n28477), .B(n19929), .Z(n19931) );
  ANDN U24208 ( .B(n19931), .A(n19930), .Z(n19932) );
  NAND U24209 ( .A(n19932), .B(n28479), .Z(n19933) );
  NANDN U24210 ( .A(n28483), .B(n19933), .Z(n19934) );
  AND U24211 ( .A(n19935), .B(n19934), .Z(n19936) );
  OR U24212 ( .A(n28488), .B(n19936), .Z(n19937) );
  NANDN U24213 ( .A(n28490), .B(n19937), .Z(n19938) );
  NANDN U24214 ( .A(n28493), .B(n19938), .Z(n19941) );
  NANDN U24215 ( .A(n19940), .B(n19939), .Z(n28495) );
  ANDN U24216 ( .B(n19941), .A(n28495), .Z(n19944) );
  NANDN U24217 ( .A(y[3965]), .B(x[3965]), .Z(n19943) );
  ANDN U24218 ( .B(n19943), .A(n19942), .Z(n28496) );
  NANDN U24219 ( .A(n19944), .B(n28496), .Z(n19947) );
  NANDN U24220 ( .A(x[3965]), .B(y[3965]), .Z(n19946) );
  ANDN U24221 ( .B(n19946), .A(n19945), .Z(n28499) );
  NAND U24222 ( .A(n19947), .B(n28499), .Z(n19948) );
  AND U24223 ( .A(n28500), .B(n19948), .Z(n19951) );
  NANDN U24224 ( .A(x[3967]), .B(y[3967]), .Z(n19950) );
  ANDN U24225 ( .B(n19950), .A(n19949), .Z(n28503) );
  NANDN U24226 ( .A(n19951), .B(n28503), .Z(n19954) );
  NOR U24227 ( .A(n19953), .B(n19952), .Z(n28504) );
  NAND U24228 ( .A(n19954), .B(n28504), .Z(n19955) );
  NANDN U24229 ( .A(n19956), .B(n19955), .Z(n19959) );
  NANDN U24230 ( .A(y[3970]), .B(x[3970]), .Z(n19958) );
  ANDN U24231 ( .B(n19958), .A(n19957), .Z(n28510) );
  NAND U24232 ( .A(n19959), .B(n28510), .Z(n19960) );
  NANDN U24233 ( .A(n19961), .B(n19960), .Z(n19962) );
  AND U24234 ( .A(n28516), .B(n19962), .Z(n19965) );
  NANDN U24235 ( .A(x[3973]), .B(y[3973]), .Z(n19964) );
  ANDN U24236 ( .B(n19964), .A(n19963), .Z(n28519) );
  NANDN U24237 ( .A(n19965), .B(n28519), .Z(n19968) );
  NANDN U24238 ( .A(y[3975]), .B(x[3975]), .Z(n19967) );
  ANDN U24239 ( .B(n19967), .A(n19966), .Z(n28520) );
  NAND U24240 ( .A(n19968), .B(n28520), .Z(n19971) );
  NANDN U24241 ( .A(x[3975]), .B(y[3975]), .Z(n19970) );
  ANDN U24242 ( .B(n19970), .A(n19969), .Z(n28522) );
  NAND U24243 ( .A(n19971), .B(n28522), .Z(n19972) );
  AND U24244 ( .A(n28524), .B(n19972), .Z(n19975) );
  NANDN U24245 ( .A(x[3977]), .B(y[3977]), .Z(n19974) );
  ANDN U24246 ( .B(n19974), .A(n19973), .Z(n28527) );
  NANDN U24247 ( .A(n19975), .B(n28527), .Z(n19976) );
  AND U24248 ( .A(n28528), .B(n19976), .Z(n19979) );
  NANDN U24249 ( .A(x[3979]), .B(y[3979]), .Z(n19977) );
  NANDN U24250 ( .A(n19978), .B(n19977), .Z(n28530) );
  OR U24251 ( .A(n19979), .B(n28530), .Z(n19980) );
  NANDN U24252 ( .A(n28533), .B(n19980), .Z(n19981) );
  AND U24253 ( .A(n19982), .B(n19981), .Z(n19983) );
  OR U24254 ( .A(n28539), .B(n19983), .Z(n19984) );
  NANDN U24255 ( .A(n28540), .B(n19984), .Z(n19987) );
  ANDN U24256 ( .B(n19986), .A(n19985), .Z(n28542) );
  NAND U24257 ( .A(n19987), .B(n28542), .Z(n19990) );
  NANDN U24258 ( .A(x[3985]), .B(y[3985]), .Z(n19988) );
  NAND U24259 ( .A(n19989), .B(n19988), .Z(n28544) );
  ANDN U24260 ( .B(n19990), .A(n28544), .Z(n19991) );
  OR U24261 ( .A(n28547), .B(n19991), .Z(n19994) );
  OR U24262 ( .A(n19993), .B(n19992), .Z(n28549) );
  ANDN U24263 ( .B(n19994), .A(n28549), .Z(n19997) );
  ANDN U24264 ( .B(n19996), .A(n19995), .Z(n28550) );
  NANDN U24265 ( .A(n19997), .B(n28550), .Z(n19998) );
  NANDN U24266 ( .A(n28552), .B(n19998), .Z(n20001) );
  NANDN U24267 ( .A(y[3990]), .B(x[3990]), .Z(n20000) );
  ANDN U24268 ( .B(n20000), .A(n19999), .Z(n28554) );
  NAND U24269 ( .A(n20001), .B(n28554), .Z(n20002) );
  AND U24270 ( .A(n28556), .B(n20002), .Z(n20005) );
  NANDN U24271 ( .A(y[3992]), .B(x[3992]), .Z(n20003) );
  NAND U24272 ( .A(n20004), .B(n20003), .Z(n28558) );
  OR U24273 ( .A(n20005), .B(n28558), .Z(n20006) );
  NANDN U24274 ( .A(n28561), .B(n20006), .Z(n20009) );
  NANDN U24275 ( .A(y[3994]), .B(x[3994]), .Z(n20007) );
  NAND U24276 ( .A(n20008), .B(n20007), .Z(n28563) );
  ANDN U24277 ( .B(n20009), .A(n28563), .Z(n20010) );
  OR U24278 ( .A(n28565), .B(n20010), .Z(n20011) );
  NANDN U24279 ( .A(n28566), .B(n20011), .Z(n20012) );
  NANDN U24280 ( .A(n28568), .B(n20012), .Z(n20015) );
  NANDN U24281 ( .A(y[3998]), .B(x[3998]), .Z(n20013) );
  NAND U24282 ( .A(n20014), .B(n20013), .Z(n28570) );
  ANDN U24283 ( .B(n20015), .A(n28570), .Z(n20016) );
  OR U24284 ( .A(n28573), .B(n20016), .Z(n20019) );
  NANDN U24285 ( .A(y[4000]), .B(x[4000]), .Z(n20017) );
  NAND U24286 ( .A(n20018), .B(n20017), .Z(n28575) );
  ANDN U24287 ( .B(n20019), .A(n28575), .Z(n20020) );
  OR U24288 ( .A(n28577), .B(n20020), .Z(n20021) );
  NANDN U24289 ( .A(n28578), .B(n20021), .Z(n20022) );
  NANDN U24290 ( .A(n28581), .B(n20022), .Z(n20023) );
  NAND U24291 ( .A(n20023), .B(n28582), .Z(n20024) );
  AND U24292 ( .A(n28584), .B(n20024), .Z(n20025) );
  NANDN U24293 ( .A(n20025), .B(n28587), .Z(n20026) );
  NAND U24294 ( .A(n20026), .B(n28588), .Z(n20027) );
  NAND U24295 ( .A(n20027), .B(n28590), .Z(n20028) );
  AND U24296 ( .A(n28592), .B(n20028), .Z(n20029) );
  OR U24297 ( .A(n28594), .B(n20029), .Z(n20032) );
  NANDN U24298 ( .A(n20031), .B(n20030), .Z(n28597) );
  ANDN U24299 ( .B(n20032), .A(n28597), .Z(n20033) );
  OR U24300 ( .A(n28599), .B(n20033), .Z(n20034) );
  NANDN U24301 ( .A(n28600), .B(n20034), .Z(n20035) );
  NANDN U24302 ( .A(n28603), .B(n20035), .Z(n20038) );
  NANDN U24303 ( .A(x[4015]), .B(y[4015]), .Z(n20036) );
  NAND U24304 ( .A(n20037), .B(n20036), .Z(n28605) );
  ANDN U24305 ( .B(n20038), .A(n28605), .Z(n20041) );
  NANDN U24306 ( .A(y[4017]), .B(x[4017]), .Z(n20040) );
  ANDN U24307 ( .B(n20040), .A(n20039), .Z(n28606) );
  NANDN U24308 ( .A(n20041), .B(n28606), .Z(n20044) );
  NANDN U24309 ( .A(x[4017]), .B(y[4017]), .Z(n20043) );
  ANDN U24310 ( .B(n20043), .A(n20042), .Z(n28609) );
  NAND U24311 ( .A(n20044), .B(n28609), .Z(n20045) );
  AND U24312 ( .A(n28610), .B(n20045), .Z(n20048) );
  NANDN U24313 ( .A(x[4019]), .B(y[4019]), .Z(n20047) );
  ANDN U24314 ( .B(n20047), .A(n20046), .Z(n28613) );
  NANDN U24315 ( .A(n20048), .B(n28613), .Z(n20051) );
  NANDN U24316 ( .A(y[4021]), .B(x[4021]), .Z(n20050) );
  ANDN U24317 ( .B(n20050), .A(n20049), .Z(n28614) );
  NAND U24318 ( .A(n20051), .B(n28614), .Z(n20052) );
  NANDN U24319 ( .A(n28617), .B(n20052), .Z(n20055) );
  NOR U24320 ( .A(n20054), .B(n20053), .Z(n28618) );
  NAND U24321 ( .A(n20055), .B(n28618), .Z(n20056) );
  NANDN U24322 ( .A(n20057), .B(n20056), .Z(n20058) );
  AND U24323 ( .A(n28624), .B(n20058), .Z(n20059) );
  OR U24324 ( .A(n28627), .B(n20059), .Z(n20060) );
  NANDN U24325 ( .A(n28629), .B(n20060), .Z(n20061) );
  NANDN U24326 ( .A(n20062), .B(n20061), .Z(n20063) );
  AND U24327 ( .A(n28634), .B(n20063), .Z(n20064) );
  OR U24328 ( .A(n28637), .B(n20064), .Z(n20065) );
  NAND U24329 ( .A(n20065), .B(n28638), .Z(n20066) );
  ANDN U24330 ( .B(n20066), .A(n28640), .Z(n20067) );
  NANDN U24331 ( .A(n20067), .B(n28642), .Z(n20070) );
  OR U24332 ( .A(n20069), .B(n20068), .Z(n28645) );
  ANDN U24333 ( .B(n20070), .A(n28645), .Z(n20071) );
  OR U24334 ( .A(n28647), .B(n20071), .Z(n20074) );
  XOR U24335 ( .A(x[4036]), .B(n20075), .Z(n20072) );
  AND U24336 ( .A(n28651), .B(n20072), .Z(n20073) );
  NAND U24337 ( .A(n20074), .B(n20073), .Z(n20078) );
  NAND U24338 ( .A(n20075), .B(x[4036]), .Z(n20077) );
  ANDN U24339 ( .B(n20077), .A(n20076), .Z(n28652) );
  NAND U24340 ( .A(n20078), .B(n28652), .Z(n20079) );
  NAND U24341 ( .A(n20080), .B(n20079), .Z(n20083) );
  NANDN U24342 ( .A(y[4038]), .B(x[4038]), .Z(n20082) );
  ANDN U24343 ( .B(n20082), .A(n20081), .Z(n28658) );
  NAND U24344 ( .A(n20083), .B(n28658), .Z(n20087) );
  NAND U24345 ( .A(n20084), .B(y[4040]), .Z(n20085) );
  NANDN U24346 ( .A(n20086), .B(n20085), .Z(n28660) );
  ANDN U24347 ( .B(n20087), .A(n28660), .Z(n20090) );
  NANDN U24348 ( .A(y[4040]), .B(x[4040]), .Z(n20089) );
  ANDN U24349 ( .B(n20089), .A(n20088), .Z(n28662) );
  NANDN U24350 ( .A(n20090), .B(n28662), .Z(n20091) );
  NANDN U24351 ( .A(n28665), .B(n20091), .Z(n20094) );
  NANDN U24352 ( .A(y[4042]), .B(x[4042]), .Z(n20093) );
  ANDN U24353 ( .B(n20093), .A(n20092), .Z(n28666) );
  NAND U24354 ( .A(n20094), .B(n28666), .Z(n20098) );
  NAND U24355 ( .A(n20095), .B(y[4044]), .Z(n20096) );
  NANDN U24356 ( .A(n20097), .B(n20096), .Z(n28668) );
  ANDN U24357 ( .B(n20098), .A(n28668), .Z(n20101) );
  NANDN U24358 ( .A(y[4044]), .B(x[4044]), .Z(n20100) );
  ANDN U24359 ( .B(n20100), .A(n20099), .Z(n28670) );
  NANDN U24360 ( .A(n20101), .B(n28670), .Z(n20102) );
  AND U24361 ( .A(n28672), .B(n20102), .Z(n20105) );
  NANDN U24362 ( .A(y[4046]), .B(x[4046]), .Z(n20104) );
  ANDN U24363 ( .B(n20104), .A(n20103), .Z(n28675) );
  NANDN U24364 ( .A(n20105), .B(n28675), .Z(n20108) );
  NANDN U24365 ( .A(x[4048]), .B(y[4048]), .Z(n20107) );
  ANDN U24366 ( .B(n20107), .A(n20106), .Z(n28676) );
  NAND U24367 ( .A(n20108), .B(n28676), .Z(n20109) );
  NANDN U24368 ( .A(n28679), .B(n20109), .Z(n20110) );
  AND U24369 ( .A(n28680), .B(n20110), .Z(n20113) );
  NOR U24370 ( .A(n20112), .B(n20111), .Z(n28682) );
  NANDN U24371 ( .A(n20113), .B(n28682), .Z(n20114) );
  AND U24372 ( .A(n20115), .B(n20114), .Z(n20116) );
  OR U24373 ( .A(n28687), .B(n20116), .Z(n20119) );
  NOR U24374 ( .A(n28690), .B(n20117), .Z(n20118) );
  NAND U24375 ( .A(n20119), .B(n20118), .Z(n20122) );
  NANDN U24376 ( .A(y[4054]), .B(x[4054]), .Z(n20121) );
  ANDN U24377 ( .B(n20121), .A(n20120), .Z(n28693) );
  NAND U24378 ( .A(n20122), .B(n28693), .Z(n20123) );
  AND U24379 ( .A(n28694), .B(n20123), .Z(n20126) );
  NANDN U24380 ( .A(y[4056]), .B(x[4056]), .Z(n20125) );
  ANDN U24381 ( .B(n20125), .A(n20124), .Z(n28696) );
  NANDN U24382 ( .A(n20126), .B(n28696), .Z(n20127) );
  AND U24383 ( .A(n28698), .B(n20127), .Z(n20130) );
  NANDN U24384 ( .A(y[4058]), .B(x[4058]), .Z(n20129) );
  ANDN U24385 ( .B(n20129), .A(n20128), .Z(n28701) );
  NANDN U24386 ( .A(n20130), .B(n28701), .Z(n20133) );
  NANDN U24387 ( .A(x[4060]), .B(y[4060]), .Z(n20132) );
  ANDN U24388 ( .B(n20132), .A(n20131), .Z(n28702) );
  NAND U24389 ( .A(n20133), .B(n28702), .Z(n20136) );
  NANDN U24390 ( .A(y[4060]), .B(x[4060]), .Z(n20135) );
  ANDN U24391 ( .B(n20135), .A(n20134), .Z(n28705) );
  NAND U24392 ( .A(n20136), .B(n28705), .Z(n20137) );
  AND U24393 ( .A(n28706), .B(n20137), .Z(n20138) );
  OR U24394 ( .A(n28709), .B(n20138), .Z(n20141) );
  NOR U24395 ( .A(n20140), .B(n20139), .Z(n28710) );
  NAND U24396 ( .A(n20141), .B(n28710), .Z(n20144) );
  NOR U24397 ( .A(n20143), .B(n20142), .Z(n28712) );
  NAND U24398 ( .A(n20144), .B(n28712), .Z(n20145) );
  NAND U24399 ( .A(n20146), .B(n20145), .Z(n20149) );
  NANDN U24400 ( .A(y[4066]), .B(x[4066]), .Z(n20148) );
  ANDN U24401 ( .B(n20148), .A(n20147), .Z(n28719) );
  NAND U24402 ( .A(n20149), .B(n28719), .Z(n20150) );
  AND U24403 ( .A(n28720), .B(n20150), .Z(n20151) );
  OR U24404 ( .A(n28723), .B(n20151), .Z(n20154) );
  NANDN U24405 ( .A(x[4070]), .B(y[4070]), .Z(n20153) );
  ANDN U24406 ( .B(n20153), .A(n20152), .Z(n28724) );
  NAND U24407 ( .A(n20154), .B(n28724), .Z(n20155) );
  NANDN U24408 ( .A(n28726), .B(n20155), .Z(n20156) );
  NANDN U24409 ( .A(n28729), .B(n20156), .Z(n20157) );
  NANDN U24410 ( .A(n28731), .B(n20157), .Z(n20158) );
  AND U24411 ( .A(n20159), .B(n20158), .Z(n20160) );
  OR U24412 ( .A(n28736), .B(n20160), .Z(n20161) );
  NANDN U24413 ( .A(n28738), .B(n20161), .Z(n20162) );
  NANDN U24414 ( .A(n28741), .B(n20162), .Z(n20165) );
  NANDN U24415 ( .A(x[4077]), .B(y[4077]), .Z(n20164) );
  NAND U24416 ( .A(n20164), .B(n20163), .Z(n28743) );
  ANDN U24417 ( .B(n20165), .A(n28743), .Z(n20166) );
  OR U24418 ( .A(n28745), .B(n20166), .Z(n20169) );
  NANDN U24419 ( .A(x[4079]), .B(y[4079]), .Z(n20167) );
  NANDN U24420 ( .A(n20168), .B(n20167), .Z(n28746) );
  ANDN U24421 ( .B(n20169), .A(n28746), .Z(n20170) );
  OR U24422 ( .A(n28749), .B(n20170), .Z(n20173) );
  ANDN U24423 ( .B(n20199), .A(n20171), .Z(n20172) );
  NAND U24424 ( .A(n20173), .B(n20172), .Z(n20174) );
  NANDN U24425 ( .A(n28753), .B(n20174), .Z(n20175) );
  NAND U24426 ( .A(n20176), .B(n20175), .Z(n20177) );
  AND U24427 ( .A(n20178), .B(n20177), .Z(n20179) );
  NAND U24428 ( .A(e), .B(n20179), .Z(n5) );
  ANDN U24429 ( .B(e), .A(n20179), .Z(n28770) );
  OR U24430 ( .A(g), .B(n28770), .Z(n28773) );
  NOR U24431 ( .A(n20181), .B(n20180), .Z(n20185) );
  NANDN U24432 ( .A(n20183), .B(n20182), .Z(n20184) );
  AND U24433 ( .A(n20185), .B(n20184), .Z(n20186) );
  OR U24434 ( .A(n20187), .B(n20186), .Z(n20188) );
  NANDN U24435 ( .A(n20189), .B(n20188), .Z(n20191) );
  NAND U24436 ( .A(n20191), .B(n20190), .Z(n28769) );
  NANDN U24437 ( .A(x[4087]), .B(y[4087]), .Z(n20193) );
  NAND U24438 ( .A(n20193), .B(n20192), .Z(n28765) );
  OR U24439 ( .A(n20195), .B(n20194), .Z(n28759) );
  NOR U24440 ( .A(n20197), .B(n20196), .Z(n28755) );
  ANDN U24441 ( .B(n20199), .A(n20198), .Z(n28751) );
  NOR U24442 ( .A(n20201), .B(n20200), .Z(n28685) );
  NOR U24443 ( .A(n20203), .B(n20202), .Z(n28419) );
  NOR U24444 ( .A(n20205), .B(n20204), .Z(n28393) );
  NOR U24445 ( .A(n20207), .B(n20206), .Z(n28381) );
  ANDN U24446 ( .B(n20209), .A(n20208), .Z(n28367) );
  NOR U24447 ( .A(n20211), .B(n20210), .Z(n28337) );
  ANDN U24448 ( .B(n20213), .A(n20212), .Z(n28193) );
  NOR U24449 ( .A(n20215), .B(n20214), .Z(n28115) );
  AND U24450 ( .A(n20217), .B(n20216), .Z(n28051) );
  NOR U24451 ( .A(n20219), .B(n20218), .Z(n28013) );
  NOR U24452 ( .A(n20221), .B(n20220), .Z(n28001) );
  ANDN U24453 ( .B(n20223), .A(n20222), .Z(n27765) );
  ANDN U24454 ( .B(n20225), .A(n20224), .Z(n27601) );
  AND U24455 ( .A(n20227), .B(n20226), .Z(n27333) );
  AND U24456 ( .A(n20229), .B(n20228), .Z(n27095) );
  ANDN U24457 ( .B(n20231), .A(n20230), .Z(n26995) );
  ANDN U24458 ( .B(n20233), .A(n20232), .Z(n26757) );
  NAND U24459 ( .A(n20234), .B(y[2869]), .Z(n26079) );
  XOR U24460 ( .A(y[2869]), .B(n20234), .Z(n26077) );
  NANDN U24461 ( .A(n20236), .B(n20235), .Z(n25837) );
  NAND U24462 ( .A(n20238), .B(n20237), .Z(n20239) );
  AND U24463 ( .A(n20240), .B(n20239), .Z(n25689) );
  NANDN U24464 ( .A(n20242), .B(n20241), .Z(n25500) );
  ANDN U24465 ( .B(n20244), .A(n20243), .Z(n25380) );
  AND U24466 ( .A(n20246), .B(n20245), .Z(n25210) );
  AND U24467 ( .A(n20248), .B(n20247), .Z(n25030) );
  XNOR U24468 ( .A(x[2438]), .B(y[2438]), .Z(n25028) );
  NANDN U24469 ( .A(n20250), .B(n20249), .Z(n24623) );
  AND U24470 ( .A(n20252), .B(n20251), .Z(n24565) );
  XNOR U24471 ( .A(y[2228]), .B(x[2228]), .Z(n24535) );
  XNOR U24472 ( .A(n20254), .B(n20253), .Z(n24531) );
  AND U24473 ( .A(n20256), .B(n20255), .Z(n24509) );
  XNOR U24474 ( .A(x[2217]), .B(y[2217]), .Z(n24507) );
  AND U24475 ( .A(n20258), .B(n20257), .Z(n24435) );
  XNOR U24476 ( .A(y[2185]), .B(x[2185]), .Z(n24433) );
  NANDN U24477 ( .A(n20260), .B(n20259), .Z(n24230) );
  ANDN U24478 ( .B(n20262), .A(n20261), .Z(n24228) );
  XNOR U24479 ( .A(y[2018]), .B(x[2018]), .Z(n24048) );
  XNOR U24480 ( .A(y[2012]), .B(x[2012]), .Z(n24034) );
  XOR U24481 ( .A(n20263), .B(x[1974]), .Z(n23942) );
  XNOR U24482 ( .A(n20265), .B(n20264), .Z(n23826) );
  NANDN U24483 ( .A(n20267), .B(n20266), .Z(n23708) );
  NAND U24484 ( .A(n20269), .B(n20268), .Z(n23694) );
  XNOR U24485 ( .A(y[1834]), .B(x[1834]), .Z(n23614) );
  NANDN U24486 ( .A(n20271), .B(n20270), .Z(n20273) );
  ANDN U24487 ( .B(n20273), .A(n20272), .Z(n23245) );
  XNOR U24488 ( .A(n20275), .B(n20274), .Z(n23205) );
  AND U24489 ( .A(n20277), .B(n20276), .Z(n23157) );
  AND U24490 ( .A(n20279), .B(n20278), .Z(n23131) );
  XNOR U24491 ( .A(x[1625]), .B(y[1625]), .Z(n23129) );
  NANDN U24492 ( .A(y[1544]), .B(x[1544]), .Z(n20280) );
  AND U24493 ( .A(n20281), .B(n20280), .Z(n22952) );
  XNOR U24494 ( .A(x[1544]), .B(y[1544]), .Z(n22950) );
  NANDN U24495 ( .A(n20283), .B(n20282), .Z(n20285) );
  ANDN U24496 ( .B(n20285), .A(n20284), .Z(n22878) );
  NAND U24497 ( .A(n20288), .B(x[1328]), .Z(n20286) );
  AND U24498 ( .A(n20287), .B(n20286), .Z(n22509) );
  XOR U24499 ( .A(x[1328]), .B(n20288), .Z(n22507) );
  AND U24500 ( .A(n20290), .B(n20289), .Z(n21853) );
  NAND U24501 ( .A(n20292), .B(n20291), .Z(n21827) );
  AND U24502 ( .A(n20294), .B(n20293), .Z(n21713) );
  NANDN U24503 ( .A(n20296), .B(n20295), .Z(n21687) );
  AND U24504 ( .A(n20298), .B(n20297), .Z(n21685) );
  NAND U24505 ( .A(n20300), .B(n20299), .Z(n20301) );
  AND U24506 ( .A(n20302), .B(n20301), .Z(n21150) );
  ANDN U24507 ( .B(n20304), .A(n20303), .Z(n20402) );
  AND U24508 ( .A(n20306), .B(n20305), .Z(n20398) );
  NANDN U24509 ( .A(n20308), .B(n20307), .Z(n20310) );
  ANDN U24510 ( .B(n20310), .A(n20309), .Z(n20312) );
  NAND U24511 ( .A(n20312), .B(n20311), .Z(n20314) );
  NAND U24512 ( .A(n20314), .B(n20313), .Z(n20315) );
  NANDN U24513 ( .A(n20316), .B(n20315), .Z(n20318) );
  ANDN U24514 ( .B(n20318), .A(n20317), .Z(n20320) );
  NANDN U24515 ( .A(n20320), .B(n20319), .Z(n20321) );
  NANDN U24516 ( .A(n20322), .B(n20321), .Z(n20324) );
  NAND U24517 ( .A(n20324), .B(n20323), .Z(n20325) );
  NANDN U24518 ( .A(n20326), .B(n20325), .Z(n20328) );
  NAND U24519 ( .A(n20328), .B(n20327), .Z(n20330) );
  ANDN U24520 ( .B(n20330), .A(n20329), .Z(n20332) );
  NANDN U24521 ( .A(n20332), .B(n20331), .Z(n20333) );
  NANDN U24522 ( .A(n20334), .B(n20333), .Z(n20336) );
  NAND U24523 ( .A(n20336), .B(n20335), .Z(n20337) );
  NANDN U24524 ( .A(n20338), .B(n20337), .Z(n20340) );
  NAND U24525 ( .A(n20340), .B(n20339), .Z(n20342) );
  ANDN U24526 ( .B(n20342), .A(n20341), .Z(n20344) );
  NANDN U24527 ( .A(n20344), .B(n20343), .Z(n20345) );
  NANDN U24528 ( .A(n20346), .B(n20345), .Z(n20348) );
  NAND U24529 ( .A(n20348), .B(n20347), .Z(n20349) );
  NANDN U24530 ( .A(n20350), .B(n20349), .Z(n20352) );
  NAND U24531 ( .A(n20352), .B(n20351), .Z(n20354) );
  ANDN U24532 ( .B(n20354), .A(n20353), .Z(n20356) );
  NANDN U24533 ( .A(n20356), .B(n20355), .Z(n20358) );
  ANDN U24534 ( .B(n20358), .A(n20357), .Z(n20360) );
  ANDN U24535 ( .B(x[312]), .A(y[312]), .Z(n20359) );
  OR U24536 ( .A(n20360), .B(n20359), .Z(n20361) );
  NANDN U24537 ( .A(n20362), .B(n20361), .Z(n20364) );
  NAND U24538 ( .A(n20364), .B(n20363), .Z(n20366) );
  NAND U24539 ( .A(n20366), .B(n20365), .Z(n20368) );
  NAND U24540 ( .A(n20368), .B(n20367), .Z(n20369) );
  AND U24541 ( .A(n20370), .B(n20369), .Z(n20372) );
  NANDN U24542 ( .A(n20372), .B(n20371), .Z(n20374) );
  NAND U24543 ( .A(n20374), .B(n20373), .Z(n20376) );
  NAND U24544 ( .A(n20376), .B(n20375), .Z(n20378) );
  NAND U24545 ( .A(n20378), .B(n20377), .Z(n20380) );
  NAND U24546 ( .A(n20380), .B(n20379), .Z(n20381) );
  AND U24547 ( .A(n20382), .B(n20381), .Z(n20384) );
  NAND U24548 ( .A(n20384), .B(n20383), .Z(n20385) );
  NANDN U24549 ( .A(n20386), .B(n20385), .Z(n20388) );
  ANDN U24550 ( .B(n20388), .A(n20387), .Z(n20389) );
  OR U24551 ( .A(n20390), .B(n20389), .Z(n20392) );
  NAND U24552 ( .A(n20392), .B(n20391), .Z(n20393) );
  AND U24553 ( .A(n20394), .B(n20393), .Z(n20396) );
  NANDN U24554 ( .A(n20396), .B(n20395), .Z(n20397) );
  AND U24555 ( .A(n20398), .B(n20397), .Z(n20399) );
  OR U24556 ( .A(n20400), .B(n20399), .Z(n20401) );
  AND U24557 ( .A(n20402), .B(n20401), .Z(n20403) );
  OR U24558 ( .A(n20404), .B(n20403), .Z(n20406) );
  NAND U24559 ( .A(n20406), .B(n20405), .Z(n20408) );
  NAND U24560 ( .A(n20408), .B(n20407), .Z(n20410) );
  NAND U24561 ( .A(n20410), .B(n20409), .Z(n20412) );
  NAND U24562 ( .A(n20412), .B(n20411), .Z(n20413) );
  AND U24563 ( .A(n20414), .B(n20413), .Z(n20416) );
  NANDN U24564 ( .A(n20416), .B(n20415), .Z(n20418) );
  NAND U24565 ( .A(n20418), .B(n20417), .Z(n20420) );
  NAND U24566 ( .A(n20420), .B(n20419), .Z(n20422) );
  NAND U24567 ( .A(n20422), .B(n20421), .Z(n20424) );
  NAND U24568 ( .A(n20424), .B(n20423), .Z(n20425) );
  AND U24569 ( .A(n20426), .B(n20425), .Z(n20428) );
  NANDN U24570 ( .A(n20428), .B(n20427), .Z(n20430) );
  NAND U24571 ( .A(n20430), .B(n20429), .Z(n20432) );
  NAND U24572 ( .A(n20432), .B(n20431), .Z(n20434) );
  NAND U24573 ( .A(n20434), .B(n20433), .Z(n20436) );
  NAND U24574 ( .A(n20436), .B(n20435), .Z(n20437) );
  AND U24575 ( .A(n20438), .B(n20437), .Z(n20440) );
  NANDN U24576 ( .A(n20440), .B(n20439), .Z(n20442) );
  NAND U24577 ( .A(n20442), .B(n20441), .Z(n20444) );
  NAND U24578 ( .A(n20444), .B(n20443), .Z(n20446) );
  NAND U24579 ( .A(n20446), .B(n20445), .Z(n20448) );
  NAND U24580 ( .A(n20448), .B(n20447), .Z(n20449) );
  AND U24581 ( .A(n20450), .B(n20449), .Z(n20451) );
  OR U24582 ( .A(n20452), .B(n20451), .Z(n20454) );
  NAND U24583 ( .A(n20454), .B(n20453), .Z(n20456) );
  NAND U24584 ( .A(n20456), .B(n20455), .Z(n20458) );
  NAND U24585 ( .A(n20458), .B(n20457), .Z(n20460) );
  NAND U24586 ( .A(n20460), .B(n20459), .Z(n20461) );
  AND U24587 ( .A(n20462), .B(n20461), .Z(n20464) );
  NANDN U24588 ( .A(n20464), .B(n20463), .Z(n20465) );
  AND U24589 ( .A(n20466), .B(n20465), .Z(n20468) );
  NANDN U24590 ( .A(n20468), .B(n20467), .Z(n20470) );
  NAND U24591 ( .A(n20470), .B(n20469), .Z(n20472) );
  NAND U24592 ( .A(n20472), .B(n20471), .Z(n20473) );
  NAND U24593 ( .A(n20474), .B(n20473), .Z(n20475) );
  NANDN U24594 ( .A(n20476), .B(n20475), .Z(n20478) );
  ANDN U24595 ( .B(n20478), .A(n20477), .Z(n20480) );
  NANDN U24596 ( .A(n20480), .B(n20479), .Z(n20482) );
  NAND U24597 ( .A(n20482), .B(n20481), .Z(n20484) );
  NAND U24598 ( .A(n20484), .B(n20483), .Z(n20485) );
  NANDN U24599 ( .A(n20486), .B(n20485), .Z(n20488) );
  NAND U24600 ( .A(n20488), .B(n20487), .Z(n20489) );
  AND U24601 ( .A(n20490), .B(n20489), .Z(n20492) );
  NANDN U24602 ( .A(n20492), .B(n20491), .Z(n20494) );
  NAND U24603 ( .A(n20494), .B(n20493), .Z(n20496) );
  NAND U24604 ( .A(n20496), .B(n20495), .Z(n20497) );
  NANDN U24605 ( .A(n20498), .B(n20497), .Z(n20499) );
  NANDN U24606 ( .A(n20500), .B(n20499), .Z(n20501) );
  AND U24607 ( .A(n20502), .B(n20501), .Z(n20504) );
  NANDN U24608 ( .A(n20504), .B(n20503), .Z(n20506) );
  NAND U24609 ( .A(n20506), .B(n20505), .Z(n20508) );
  NAND U24610 ( .A(n20508), .B(n20507), .Z(n20510) );
  NAND U24611 ( .A(n20510), .B(n20509), .Z(n20512) );
  NAND U24612 ( .A(n20512), .B(n20511), .Z(n20513) );
  AND U24613 ( .A(n20514), .B(n20513), .Z(n20516) );
  NANDN U24614 ( .A(n20516), .B(n20515), .Z(n20518) );
  NAND U24615 ( .A(n20518), .B(n20517), .Z(n20520) );
  NAND U24616 ( .A(n20520), .B(n20519), .Z(n20522) );
  NAND U24617 ( .A(n20522), .B(n20521), .Z(n20524) );
  NAND U24618 ( .A(n20524), .B(n20523), .Z(n20525) );
  AND U24619 ( .A(n20526), .B(n20525), .Z(n20528) );
  NANDN U24620 ( .A(n20528), .B(n20527), .Z(n20530) );
  NAND U24621 ( .A(n20530), .B(n20529), .Z(n20532) );
  NAND U24622 ( .A(n20532), .B(n20531), .Z(n20534) );
  NAND U24623 ( .A(n20534), .B(n20533), .Z(n20536) );
  NAND U24624 ( .A(n20536), .B(n20535), .Z(n20537) );
  AND U24625 ( .A(n20538), .B(n20537), .Z(n20540) );
  NANDN U24626 ( .A(n20540), .B(n20539), .Z(n20542) );
  NAND U24627 ( .A(n20542), .B(n20541), .Z(n20544) );
  NAND U24628 ( .A(n20544), .B(n20543), .Z(n20546) );
  NAND U24629 ( .A(n20546), .B(n20545), .Z(n20548) );
  NAND U24630 ( .A(n20548), .B(n20547), .Z(n20549) );
  AND U24631 ( .A(n20550), .B(n20549), .Z(n20552) );
  NANDN U24632 ( .A(n20552), .B(n20551), .Z(n20554) );
  NAND U24633 ( .A(n20554), .B(n20553), .Z(n20556) );
  NAND U24634 ( .A(n20556), .B(n20555), .Z(n20558) );
  NAND U24635 ( .A(n20558), .B(n20557), .Z(n20560) );
  NAND U24636 ( .A(n20560), .B(n20559), .Z(n20561) );
  AND U24637 ( .A(n20562), .B(n20561), .Z(n20564) );
  NANDN U24638 ( .A(n20564), .B(n20563), .Z(n20566) );
  NAND U24639 ( .A(n20566), .B(n20565), .Z(n20568) );
  NAND U24640 ( .A(n20568), .B(n20567), .Z(n20570) );
  NAND U24641 ( .A(n20570), .B(n20569), .Z(n20572) );
  NAND U24642 ( .A(n20572), .B(n20571), .Z(n20573) );
  AND U24643 ( .A(n20574), .B(n20573), .Z(n20576) );
  NANDN U24644 ( .A(n20576), .B(n20575), .Z(n20578) );
  NAND U24645 ( .A(n20578), .B(n20577), .Z(n20580) );
  NAND U24646 ( .A(n20580), .B(n20579), .Z(n20582) );
  NAND U24647 ( .A(n20582), .B(n20581), .Z(n20584) );
  NAND U24648 ( .A(n20584), .B(n20583), .Z(n20585) );
  AND U24649 ( .A(n20586), .B(n20585), .Z(n20588) );
  NANDN U24650 ( .A(n20588), .B(n20587), .Z(n20589) );
  AND U24651 ( .A(n20590), .B(n20589), .Z(n20592) );
  NANDN U24652 ( .A(n20592), .B(n20591), .Z(n20594) );
  NAND U24653 ( .A(n20594), .B(n20593), .Z(n20596) );
  NAND U24654 ( .A(n20596), .B(n20595), .Z(n20597) );
  NAND U24655 ( .A(n20598), .B(n20597), .Z(n20599) );
  NANDN U24656 ( .A(n20600), .B(n20599), .Z(n20602) );
  ANDN U24657 ( .B(n20602), .A(n20601), .Z(n20604) );
  NANDN U24658 ( .A(n20604), .B(n20603), .Z(n20606) );
  NAND U24659 ( .A(n20606), .B(n20605), .Z(n20608) );
  NAND U24660 ( .A(n20608), .B(n20607), .Z(n20610) );
  NAND U24661 ( .A(n20610), .B(n20609), .Z(n20612) );
  NAND U24662 ( .A(n20612), .B(n20611), .Z(n20613) );
  AND U24663 ( .A(n20614), .B(n20613), .Z(n20616) );
  NANDN U24664 ( .A(n20616), .B(n20615), .Z(n20618) );
  NAND U24665 ( .A(n20618), .B(n20617), .Z(n20620) );
  NAND U24666 ( .A(n20620), .B(n20619), .Z(n20621) );
  NAND U24667 ( .A(n20622), .B(n20621), .Z(n20625) );
  XOR U24668 ( .A(n20622), .B(n20621), .Z(n20623) );
  NAND U24669 ( .A(n20623), .B(y[436]), .Z(n20624) );
  NAND U24670 ( .A(n20625), .B(n20624), .Z(n20626) );
  AND U24671 ( .A(n20627), .B(n20626), .Z(n20629) );
  NANDN U24672 ( .A(n20629), .B(n20628), .Z(n20631) );
  NAND U24673 ( .A(n20631), .B(n20630), .Z(n20633) );
  NAND U24674 ( .A(n20633), .B(n20632), .Z(n20635) );
  NAND U24675 ( .A(n20635), .B(n20634), .Z(n20637) );
  NAND U24676 ( .A(n20637), .B(n20636), .Z(n20638) );
  AND U24677 ( .A(n20639), .B(n20638), .Z(n20641) );
  NANDN U24678 ( .A(n20641), .B(n20640), .Z(n20643) );
  NAND U24679 ( .A(n20643), .B(n20642), .Z(n20645) );
  NAND U24680 ( .A(n20645), .B(n20644), .Z(n20647) );
  NAND U24681 ( .A(n20647), .B(n20646), .Z(n20649) );
  NAND U24682 ( .A(n20649), .B(n20648), .Z(n20650) );
  AND U24683 ( .A(n20651), .B(n20650), .Z(n20653) );
  NANDN U24684 ( .A(n20653), .B(n20652), .Z(n20655) );
  NAND U24685 ( .A(n20655), .B(n20654), .Z(n20657) );
  NAND U24686 ( .A(n20657), .B(n20656), .Z(n20658) );
  NANDN U24687 ( .A(n20659), .B(n20658), .Z(n20661) );
  NAND U24688 ( .A(n20661), .B(n20660), .Z(n20662) );
  AND U24689 ( .A(n20663), .B(n20662), .Z(n20665) );
  NANDN U24690 ( .A(n20665), .B(n20664), .Z(n20667) );
  NAND U24691 ( .A(n20667), .B(n20666), .Z(n20669) );
  NAND U24692 ( .A(n20669), .B(n20668), .Z(n20671) );
  NAND U24693 ( .A(n20671), .B(n20670), .Z(n20673) );
  NAND U24694 ( .A(n20673), .B(n20672), .Z(n20674) );
  AND U24695 ( .A(n20675), .B(n20674), .Z(n20677) );
  NANDN U24696 ( .A(n20677), .B(n20676), .Z(n20679) );
  NAND U24697 ( .A(n20679), .B(n20678), .Z(n20681) );
  NAND U24698 ( .A(n20681), .B(n20680), .Z(n20683) );
  NAND U24699 ( .A(n20683), .B(n20682), .Z(n20685) );
  NAND U24700 ( .A(n20685), .B(n20684), .Z(n20686) );
  AND U24701 ( .A(n20687), .B(n20686), .Z(n20689) );
  NANDN U24702 ( .A(n20689), .B(n20688), .Z(n20691) );
  NAND U24703 ( .A(n20691), .B(n20690), .Z(n20693) );
  NAND U24704 ( .A(n20693), .B(n20692), .Z(n20695) );
  NAND U24705 ( .A(n20695), .B(n20694), .Z(n20697) );
  NAND U24706 ( .A(n20697), .B(n20696), .Z(n20698) );
  AND U24707 ( .A(n20699), .B(n20698), .Z(n20701) );
  NANDN U24708 ( .A(n20701), .B(n20700), .Z(n20703) );
  NAND U24709 ( .A(n20703), .B(n20702), .Z(n20705) );
  NAND U24710 ( .A(n20705), .B(n20704), .Z(n20707) );
  NAND U24711 ( .A(n20707), .B(n20706), .Z(n20709) );
  NAND U24712 ( .A(n20709), .B(n20708), .Z(n20710) );
  AND U24713 ( .A(n20711), .B(n20710), .Z(n20713) );
  NANDN U24714 ( .A(n20713), .B(n20712), .Z(n20714) );
  NANDN U24715 ( .A(n20715), .B(n20714), .Z(n20716) );
  NANDN U24716 ( .A(n20717), .B(n20716), .Z(n20718) );
  NANDN U24717 ( .A(n20719), .B(n20718), .Z(n20721) );
  NAND U24718 ( .A(n20721), .B(n20720), .Z(n20723) );
  ANDN U24719 ( .B(n20723), .A(n20722), .Z(n20725) );
  NANDN U24720 ( .A(n20725), .B(n20724), .Z(n20726) );
  NANDN U24721 ( .A(n20727), .B(n20726), .Z(n20729) );
  NAND U24722 ( .A(n20729), .B(n20728), .Z(n20730) );
  NANDN U24723 ( .A(n20731), .B(n20730), .Z(n20733) );
  NAND U24724 ( .A(n20733), .B(n20732), .Z(n20735) );
  ANDN U24725 ( .B(n20735), .A(n20734), .Z(n20737) );
  NANDN U24726 ( .A(n20737), .B(n20736), .Z(n20738) );
  NANDN U24727 ( .A(n20739), .B(n20738), .Z(n20741) );
  NAND U24728 ( .A(n20741), .B(n20740), .Z(n20742) );
  NANDN U24729 ( .A(n20743), .B(n20742), .Z(n20745) );
  NAND U24730 ( .A(n20745), .B(n20744), .Z(n20747) );
  ANDN U24731 ( .B(n20747), .A(n20746), .Z(n20749) );
  NANDN U24732 ( .A(n20749), .B(n20748), .Z(n20750) );
  NANDN U24733 ( .A(n20751), .B(n20750), .Z(n20753) );
  NAND U24734 ( .A(n20753), .B(n20752), .Z(n20754) );
  NANDN U24735 ( .A(n20755), .B(n20754), .Z(n20757) );
  NAND U24736 ( .A(n20757), .B(n20756), .Z(n20759) );
  ANDN U24737 ( .B(n20759), .A(n20758), .Z(n20761) );
  NANDN U24738 ( .A(n20761), .B(n20760), .Z(n20762) );
  NANDN U24739 ( .A(n20763), .B(n20762), .Z(n20765) );
  NAND U24740 ( .A(n20765), .B(n20764), .Z(n20766) );
  NANDN U24741 ( .A(n20767), .B(n20766), .Z(n20769) );
  NAND U24742 ( .A(n20769), .B(n20768), .Z(n20771) );
  ANDN U24743 ( .B(n20771), .A(n20770), .Z(n20773) );
  NANDN U24744 ( .A(n20773), .B(n20772), .Z(n20774) );
  NANDN U24745 ( .A(n20775), .B(n20774), .Z(n20777) );
  NAND U24746 ( .A(n20777), .B(n20776), .Z(n20779) );
  NAND U24747 ( .A(n20779), .B(n20778), .Z(n20780) );
  NANDN U24748 ( .A(n20781), .B(n20780), .Z(n20783) );
  ANDN U24749 ( .B(n20783), .A(n20782), .Z(n20785) );
  NANDN U24750 ( .A(n20785), .B(n20784), .Z(n20786) );
  NANDN U24751 ( .A(n20787), .B(n20786), .Z(n20789) );
  NAND U24752 ( .A(n20789), .B(n20788), .Z(n20790) );
  NANDN U24753 ( .A(n20791), .B(n20790), .Z(n20793) );
  NAND U24754 ( .A(n20793), .B(n20792), .Z(n20795) );
  ANDN U24755 ( .B(n20795), .A(n20794), .Z(n20797) );
  NANDN U24756 ( .A(n20797), .B(n20796), .Z(n20798) );
  NANDN U24757 ( .A(n20799), .B(n20798), .Z(n20801) );
  NAND U24758 ( .A(n20801), .B(n20800), .Z(n20802) );
  NANDN U24759 ( .A(n20803), .B(n20802), .Z(n20805) );
  NAND U24760 ( .A(n20805), .B(n20804), .Z(n20806) );
  AND U24761 ( .A(n20807), .B(n20806), .Z(n20808) );
  OR U24762 ( .A(n20809), .B(n20808), .Z(n20810) );
  NANDN U24763 ( .A(n20811), .B(n20810), .Z(n20813) );
  NAND U24764 ( .A(n20813), .B(n20812), .Z(n20814) );
  NANDN U24765 ( .A(n20815), .B(n20814), .Z(n20817) );
  NAND U24766 ( .A(n20817), .B(n20816), .Z(n20819) );
  ANDN U24767 ( .B(n20819), .A(n20818), .Z(n20821) );
  NANDN U24768 ( .A(n20821), .B(n20820), .Z(n20822) );
  NANDN U24769 ( .A(n20823), .B(n20822), .Z(n20825) );
  NAND U24770 ( .A(n20825), .B(n20824), .Z(n20826) );
  NANDN U24771 ( .A(n20827), .B(n20826), .Z(n20829) );
  NAND U24772 ( .A(n20829), .B(n20828), .Z(n20831) );
  ANDN U24773 ( .B(n20831), .A(n20830), .Z(n20833) );
  NANDN U24774 ( .A(n20833), .B(n20832), .Z(n20834) );
  NANDN U24775 ( .A(n20835), .B(n20834), .Z(n20837) );
  NAND U24776 ( .A(n20837), .B(n20836), .Z(n20838) );
  NANDN U24777 ( .A(n20839), .B(n20838), .Z(n20841) );
  NAND U24778 ( .A(n20841), .B(n20840), .Z(n20843) );
  ANDN U24779 ( .B(n20843), .A(n20842), .Z(n20845) );
  NANDN U24780 ( .A(n20845), .B(n20844), .Z(n20846) );
  NANDN U24781 ( .A(n20847), .B(n20846), .Z(n20849) );
  NAND U24782 ( .A(n20849), .B(n20848), .Z(n20850) );
  NANDN U24783 ( .A(n20851), .B(n20850), .Z(n20853) );
  NAND U24784 ( .A(n20853), .B(n20852), .Z(n20855) );
  ANDN U24785 ( .B(n20855), .A(n20854), .Z(n20857) );
  NANDN U24786 ( .A(n20857), .B(n20856), .Z(n20858) );
  NANDN U24787 ( .A(n20859), .B(n20858), .Z(n20860) );
  NANDN U24788 ( .A(n20861), .B(n20860), .Z(n20862) );
  NANDN U24789 ( .A(n20863), .B(n20862), .Z(n20865) );
  NAND U24790 ( .A(n20865), .B(n20864), .Z(n20867) );
  ANDN U24791 ( .B(n20867), .A(n20866), .Z(n20869) );
  NANDN U24792 ( .A(n20869), .B(n20868), .Z(n20870) );
  NANDN U24793 ( .A(n20871), .B(n20870), .Z(n20873) );
  NAND U24794 ( .A(n20873), .B(n20872), .Z(n20874) );
  NANDN U24795 ( .A(n20875), .B(n20874), .Z(n20877) );
  NAND U24796 ( .A(n20877), .B(n20876), .Z(n20878) );
  AND U24797 ( .A(n20879), .B(n20878), .Z(n20885) );
  NAND U24798 ( .A(n20881), .B(n20880), .Z(n20883) );
  NAND U24799 ( .A(n20883), .B(n20882), .Z(n20884) );
  NANDN U24800 ( .A(n20885), .B(n20884), .Z(n20886) );
  NANDN U24801 ( .A(n20887), .B(n20886), .Z(n20888) );
  NANDN U24802 ( .A(n20889), .B(n20888), .Z(n20890) );
  AND U24803 ( .A(n20891), .B(n20890), .Z(n20893) );
  NANDN U24804 ( .A(n20893), .B(n20892), .Z(n20895) );
  NAND U24805 ( .A(n20895), .B(n20894), .Z(n20897) );
  NAND U24806 ( .A(n20897), .B(n20896), .Z(n20899) );
  NAND U24807 ( .A(n20899), .B(n20898), .Z(n20901) );
  NAND U24808 ( .A(n20901), .B(n20900), .Z(n20902) );
  AND U24809 ( .A(n20903), .B(n20902), .Z(n20904) );
  OR U24810 ( .A(n20905), .B(n20904), .Z(n20907) );
  NAND U24811 ( .A(n20907), .B(n20906), .Z(n20909) );
  ANDN U24812 ( .B(n20909), .A(n20908), .Z(n20911) );
  NANDN U24813 ( .A(n20911), .B(n20910), .Z(n20913) );
  NAND U24814 ( .A(n20913), .B(n20912), .Z(n20915) );
  NAND U24815 ( .A(n20915), .B(n20914), .Z(n20916) );
  NANDN U24816 ( .A(n20917), .B(n20916), .Z(n20919) );
  NAND U24817 ( .A(n20919), .B(n20918), .Z(n20921) );
  ANDN U24818 ( .B(n20921), .A(n20920), .Z(n20923) );
  NANDN U24819 ( .A(n20923), .B(n20922), .Z(n20924) );
  NANDN U24820 ( .A(n20925), .B(n20924), .Z(n20927) );
  NAND U24821 ( .A(n20927), .B(n20926), .Z(n20928) );
  NANDN U24822 ( .A(n20929), .B(n20928), .Z(n20930) );
  NANDN U24823 ( .A(n20931), .B(n20930), .Z(n20932) );
  AND U24824 ( .A(n20933), .B(n20932), .Z(n20935) );
  NANDN U24825 ( .A(n20935), .B(n20934), .Z(n20936) );
  NANDN U24826 ( .A(n20937), .B(n20936), .Z(n20939) );
  NAND U24827 ( .A(n20939), .B(n20938), .Z(n20940) );
  NANDN U24828 ( .A(n20941), .B(n20940), .Z(n20943) );
  NAND U24829 ( .A(n20943), .B(n20942), .Z(n20945) );
  ANDN U24830 ( .B(n20945), .A(n20944), .Z(n20947) );
  NANDN U24831 ( .A(n20947), .B(n20946), .Z(n20948) );
  NANDN U24832 ( .A(n20949), .B(n20948), .Z(n20951) );
  NAND U24833 ( .A(n20951), .B(n20950), .Z(n20952) );
  NANDN U24834 ( .A(n20953), .B(n20952), .Z(n20954) );
  NANDN U24835 ( .A(n20955), .B(n20954), .Z(n20957) );
  ANDN U24836 ( .B(n20957), .A(n20956), .Z(n20958) );
  OR U24837 ( .A(n20959), .B(n20958), .Z(n20960) );
  NANDN U24838 ( .A(n20961), .B(n20960), .Z(n20963) );
  NAND U24839 ( .A(n20963), .B(n20962), .Z(n20964) );
  NANDN U24840 ( .A(n20965), .B(n20964), .Z(n20967) );
  NAND U24841 ( .A(n20967), .B(n20966), .Z(n20969) );
  ANDN U24842 ( .B(n20969), .A(n20968), .Z(n20971) );
  NANDN U24843 ( .A(n20971), .B(n20970), .Z(n20972) );
  NANDN U24844 ( .A(n20973), .B(n20972), .Z(n20975) );
  NAND U24845 ( .A(n20975), .B(n20974), .Z(n20976) );
  NANDN U24846 ( .A(n20977), .B(n20976), .Z(n20979) );
  NAND U24847 ( .A(n20979), .B(n20978), .Z(n20981) );
  ANDN U24848 ( .B(n20981), .A(n20980), .Z(n20983) );
  NANDN U24849 ( .A(n20983), .B(n20982), .Z(n20984) );
  NANDN U24850 ( .A(n20985), .B(n20984), .Z(n20987) );
  NAND U24851 ( .A(n20987), .B(n20986), .Z(n20988) );
  NANDN U24852 ( .A(n20989), .B(n20988), .Z(n20991) );
  NAND U24853 ( .A(n20991), .B(n20990), .Z(n20993) );
  ANDN U24854 ( .B(n20993), .A(n20992), .Z(n20995) );
  NANDN U24855 ( .A(n20995), .B(n20994), .Z(n20996) );
  NANDN U24856 ( .A(n20997), .B(n20996), .Z(n20999) );
  NAND U24857 ( .A(n20999), .B(n20998), .Z(n21001) );
  NAND U24858 ( .A(n21001), .B(n21000), .Z(n21003) );
  NAND U24859 ( .A(n21003), .B(n21002), .Z(n21005) );
  ANDN U24860 ( .B(n21005), .A(n21004), .Z(n21007) );
  NANDN U24861 ( .A(n21007), .B(n21006), .Z(n21008) );
  NANDN U24862 ( .A(n21009), .B(n21008), .Z(n21011) );
  NAND U24863 ( .A(n21011), .B(n21010), .Z(n21012) );
  NANDN U24864 ( .A(n21013), .B(n21012), .Z(n21014) );
  AND U24865 ( .A(n21015), .B(n21014), .Z(n21016) );
  NANDN U24866 ( .A(n21017), .B(n21016), .Z(n21018) );
  NANDN U24867 ( .A(n21019), .B(n21018), .Z(n21021) );
  NAND U24868 ( .A(n21021), .B(n21020), .Z(n21022) );
  AND U24869 ( .A(n21023), .B(n21022), .Z(n21025) );
  NANDN U24870 ( .A(n21025), .B(n21024), .Z(n21026) );
  NANDN U24871 ( .A(n21027), .B(n21026), .Z(n21029) );
  NAND U24872 ( .A(n21029), .B(n21028), .Z(n21030) );
  NANDN U24873 ( .A(n21031), .B(n21030), .Z(n21033) );
  NAND U24874 ( .A(n21033), .B(n21032), .Z(n21035) );
  ANDN U24875 ( .B(n21035), .A(n21034), .Z(n21037) );
  NANDN U24876 ( .A(n21037), .B(n21036), .Z(n21038) );
  AND U24877 ( .A(n21039), .B(n21038), .Z(n21041) );
  NANDN U24878 ( .A(n21041), .B(n21040), .Z(n21042) );
  NANDN U24879 ( .A(n21043), .B(n21042), .Z(n21045) );
  NAND U24880 ( .A(n21045), .B(n21044), .Z(n21046) );
  NANDN U24881 ( .A(n21047), .B(n21046), .Z(n21048) );
  NANDN U24882 ( .A(n21049), .B(n21048), .Z(n21051) );
  NAND U24883 ( .A(n21051), .B(n21050), .Z(n21052) );
  NANDN U24884 ( .A(n21053), .B(n21052), .Z(n21055) );
  NAND U24885 ( .A(n21055), .B(n21054), .Z(n21057) );
  ANDN U24886 ( .B(n21057), .A(n21056), .Z(n21059) );
  NANDN U24887 ( .A(n21059), .B(n21058), .Z(n21060) );
  NANDN U24888 ( .A(n21061), .B(n21060), .Z(n21063) );
  NAND U24889 ( .A(n21063), .B(n21062), .Z(n21064) );
  NANDN U24890 ( .A(n21065), .B(n21064), .Z(n21067) );
  NAND U24891 ( .A(n21067), .B(n21066), .Z(n21069) );
  ANDN U24892 ( .B(n21069), .A(n21068), .Z(n21071) );
  NANDN U24893 ( .A(n21071), .B(n21070), .Z(n21072) );
  NANDN U24894 ( .A(n21073), .B(n21072), .Z(n21075) );
  NAND U24895 ( .A(n21075), .B(n21074), .Z(n21077) );
  NAND U24896 ( .A(n21077), .B(n21076), .Z(n21078) );
  NANDN U24897 ( .A(n21079), .B(n21078), .Z(n21081) );
  ANDN U24898 ( .B(n21081), .A(n21080), .Z(n21083) );
  NANDN U24899 ( .A(n21083), .B(n21082), .Z(n21084) );
  NANDN U24900 ( .A(n21085), .B(n21084), .Z(n21087) );
  NAND U24901 ( .A(n21087), .B(n21086), .Z(n21088) );
  NANDN U24902 ( .A(n21089), .B(n21088), .Z(n21091) );
  NAND U24903 ( .A(n21091), .B(n21090), .Z(n21093) );
  ANDN U24904 ( .B(n21093), .A(n21092), .Z(n21095) );
  NANDN U24905 ( .A(n21095), .B(n21094), .Z(n21097) );
  NAND U24906 ( .A(n21097), .B(n21096), .Z(n21099) );
  ANDN U24907 ( .B(n21099), .A(n21098), .Z(n21103) );
  ANDN U24908 ( .B(n21101), .A(n21100), .Z(n21102) );
  NANDN U24909 ( .A(n21103), .B(n21102), .Z(n21105) );
  NAND U24910 ( .A(n21105), .B(n21104), .Z(n21107) );
  NANDN U24911 ( .A(n21107), .B(x[675]), .Z(n21110) );
  XOR U24912 ( .A(n21107), .B(n21106), .Z(n21108) );
  NANDN U24913 ( .A(y[675]), .B(n21108), .Z(n21109) );
  AND U24914 ( .A(n21110), .B(n21109), .Z(n21113) );
  OR U24915 ( .A(n21113), .B(y[676]), .Z(n21111) );
  AND U24916 ( .A(n21112), .B(n21111), .Z(n21116) );
  XOR U24917 ( .A(y[676]), .B(n21113), .Z(n21114) );
  NAND U24918 ( .A(n21114), .B(x[676]), .Z(n21115) );
  NAND U24919 ( .A(n21116), .B(n21115), .Z(n21118) );
  NAND U24920 ( .A(n21118), .B(n21117), .Z(n21120) );
  NAND U24921 ( .A(n21120), .B(n21119), .Z(n21121) );
  AND U24922 ( .A(n21122), .B(n21121), .Z(n21124) );
  NANDN U24923 ( .A(n21124), .B(n21123), .Z(n21126) );
  NAND U24924 ( .A(n21126), .B(n21125), .Z(n21128) );
  NAND U24925 ( .A(n21128), .B(n21127), .Z(n21130) );
  NAND U24926 ( .A(n21130), .B(n21129), .Z(n21132) );
  NAND U24927 ( .A(n21132), .B(n21131), .Z(n21133) );
  AND U24928 ( .A(n21134), .B(n21133), .Z(n21136) );
  NANDN U24929 ( .A(n21136), .B(n21135), .Z(n21138) );
  NAND U24930 ( .A(n21138), .B(n21137), .Z(n21140) );
  NAND U24931 ( .A(n21140), .B(n21139), .Z(n21142) );
  NAND U24932 ( .A(n21142), .B(n21141), .Z(n21144) );
  NAND U24933 ( .A(n21144), .B(n21143), .Z(n21146) );
  ANDN U24934 ( .B(n21146), .A(n21145), .Z(n21148) );
  NANDN U24935 ( .A(n21148), .B(n21147), .Z(n21149) );
  NANDN U24936 ( .A(n21150), .B(n21149), .Z(n21152) );
  NAND U24937 ( .A(n21152), .B(n21151), .Z(n21153) );
  NANDN U24938 ( .A(n21154), .B(n21153), .Z(n21155) );
  NANDN U24939 ( .A(n21156), .B(n21155), .Z(n21158) );
  NAND U24940 ( .A(n21158), .B(n21157), .Z(n21159) );
  NANDN U24941 ( .A(n21160), .B(n21159), .Z(n21162) );
  NAND U24942 ( .A(n21162), .B(n21161), .Z(n21164) );
  ANDN U24943 ( .B(n21164), .A(n21163), .Z(n21166) );
  NANDN U24944 ( .A(n21166), .B(n21165), .Z(n21167) );
  NANDN U24945 ( .A(n21168), .B(n21167), .Z(n21170) );
  NAND U24946 ( .A(n21170), .B(n21169), .Z(n21171) );
  NANDN U24947 ( .A(n21172), .B(n21171), .Z(n21174) );
  NAND U24948 ( .A(n21174), .B(n21173), .Z(n21176) );
  ANDN U24949 ( .B(n21176), .A(n21175), .Z(n21178) );
  NANDN U24950 ( .A(n21178), .B(n21177), .Z(n21179) );
  NANDN U24951 ( .A(n21180), .B(n21179), .Z(n21182) );
  NAND U24952 ( .A(n21182), .B(n21181), .Z(n21184) );
  NAND U24953 ( .A(n21184), .B(n21183), .Z(n21185) );
  NANDN U24954 ( .A(n21186), .B(n21185), .Z(n21188) );
  ANDN U24955 ( .B(n21188), .A(n21187), .Z(n21190) );
  NANDN U24956 ( .A(n21190), .B(n21189), .Z(n21191) );
  NANDN U24957 ( .A(n21192), .B(n21191), .Z(n21194) );
  NAND U24958 ( .A(n21194), .B(n21193), .Z(n21195) );
  NANDN U24959 ( .A(n21196), .B(n21195), .Z(n21198) );
  NAND U24960 ( .A(n21198), .B(n21197), .Z(n21200) );
  ANDN U24961 ( .B(n21200), .A(n21199), .Z(n21202) );
  NANDN U24962 ( .A(n21202), .B(n21201), .Z(n21203) );
  NANDN U24963 ( .A(n21204), .B(n21203), .Z(n21206) );
  NAND U24964 ( .A(n21206), .B(n21205), .Z(n21207) );
  NANDN U24965 ( .A(n21208), .B(n21207), .Z(n21210) );
  NAND U24966 ( .A(n21210), .B(n21209), .Z(n21212) );
  ANDN U24967 ( .B(n21212), .A(n21211), .Z(n21214) );
  NANDN U24968 ( .A(n21214), .B(n21213), .Z(n21215) );
  NANDN U24969 ( .A(n21216), .B(n21215), .Z(n21218) );
  NAND U24970 ( .A(n21218), .B(n21217), .Z(n21219) );
  NANDN U24971 ( .A(n21220), .B(n21219), .Z(n21222) );
  NAND U24972 ( .A(n21222), .B(n21221), .Z(n21223) );
  AND U24973 ( .A(n21224), .B(n21223), .Z(n21225) );
  OR U24974 ( .A(n21226), .B(n21225), .Z(n21227) );
  NANDN U24975 ( .A(n21228), .B(n21227), .Z(n21230) );
  NAND U24976 ( .A(n21230), .B(n21229), .Z(n21231) );
  NANDN U24977 ( .A(n21232), .B(n21231), .Z(n21234) );
  NAND U24978 ( .A(n21234), .B(n21233), .Z(n21235) );
  AND U24979 ( .A(n21236), .B(n21235), .Z(n21238) );
  NANDN U24980 ( .A(n21238), .B(n21237), .Z(n21240) );
  NAND U24981 ( .A(n21240), .B(n21239), .Z(n21242) );
  NAND U24982 ( .A(n21242), .B(n21241), .Z(n21244) );
  NAND U24983 ( .A(n21244), .B(n21243), .Z(n21246) );
  NAND U24984 ( .A(n21246), .B(n21245), .Z(n21247) );
  AND U24985 ( .A(n21248), .B(n21247), .Z(n21250) );
  NANDN U24986 ( .A(n21250), .B(n21249), .Z(n21252) );
  NAND U24987 ( .A(n21252), .B(n21251), .Z(n21254) );
  NAND U24988 ( .A(n21254), .B(n21253), .Z(n21256) );
  ANDN U24989 ( .B(n21256), .A(n21255), .Z(n21258) );
  NAND U24990 ( .A(n21258), .B(n21257), .Z(n21259) );
  NANDN U24991 ( .A(n21260), .B(n21259), .Z(n21262) );
  ANDN U24992 ( .B(n21262), .A(n21261), .Z(n21266) );
  NANDN U24993 ( .A(n21264), .B(n21263), .Z(n21265) );
  AND U24994 ( .A(n21266), .B(n21265), .Z(n21268) );
  NANDN U24995 ( .A(n21268), .B(n21267), .Z(n21270) );
  NAND U24996 ( .A(n21270), .B(n21269), .Z(n21272) );
  NAND U24997 ( .A(n21272), .B(n21271), .Z(n21274) );
  NAND U24998 ( .A(n21274), .B(n21273), .Z(n21276) );
  NAND U24999 ( .A(n21276), .B(n21275), .Z(n21277) );
  AND U25000 ( .A(n21278), .B(n21277), .Z(n21280) );
  NANDN U25001 ( .A(n21280), .B(n21279), .Z(n21282) );
  NAND U25002 ( .A(n21282), .B(n21281), .Z(n21284) );
  NAND U25003 ( .A(n21284), .B(n21283), .Z(n21286) );
  NAND U25004 ( .A(n21286), .B(n21285), .Z(n21288) );
  NAND U25005 ( .A(n21288), .B(n21287), .Z(n21290) );
  ANDN U25006 ( .B(n21290), .A(n21289), .Z(n21292) );
  NANDN U25007 ( .A(n21292), .B(n21291), .Z(n21294) );
  NAND U25008 ( .A(n21294), .B(n21293), .Z(n21296) );
  NAND U25009 ( .A(n21296), .B(n21295), .Z(n21298) );
  NAND U25010 ( .A(n21298), .B(n21297), .Z(n21300) );
  NAND U25011 ( .A(n21300), .B(n21299), .Z(n21301) );
  AND U25012 ( .A(n21302), .B(n21301), .Z(n21304) );
  NANDN U25013 ( .A(n21304), .B(n21303), .Z(n21306) );
  ANDN U25014 ( .B(n21306), .A(n21305), .Z(n21307) );
  OR U25015 ( .A(n21308), .B(n21307), .Z(n21310) );
  NAND U25016 ( .A(n21310), .B(n21309), .Z(n21311) );
  AND U25017 ( .A(n21312), .B(n21311), .Z(n21314) );
  NANDN U25018 ( .A(n21314), .B(n21313), .Z(n21316) );
  NAND U25019 ( .A(n21316), .B(n21315), .Z(n21318) );
  NAND U25020 ( .A(n21318), .B(n21317), .Z(n21320) );
  NAND U25021 ( .A(n21320), .B(n21319), .Z(n21322) );
  NAND U25022 ( .A(n21322), .B(n21321), .Z(n21323) );
  AND U25023 ( .A(n21324), .B(n21323), .Z(n21326) );
  NANDN U25024 ( .A(n21326), .B(n21325), .Z(n21328) );
  NAND U25025 ( .A(n21328), .B(n21327), .Z(n21330) );
  NAND U25026 ( .A(n21330), .B(n21329), .Z(n21332) );
  NAND U25027 ( .A(n21332), .B(n21331), .Z(n21334) );
  NAND U25028 ( .A(n21334), .B(n21333), .Z(n21335) );
  AND U25029 ( .A(n21336), .B(n21335), .Z(n21338) );
  NANDN U25030 ( .A(n21338), .B(n21337), .Z(n21340) );
  NAND U25031 ( .A(n21340), .B(n21339), .Z(n21342) );
  NAND U25032 ( .A(n21342), .B(n21341), .Z(n21344) );
  NAND U25033 ( .A(n21344), .B(n21343), .Z(n21346) );
  NAND U25034 ( .A(n21346), .B(n21345), .Z(n21347) );
  AND U25035 ( .A(n21348), .B(n21347), .Z(n21350) );
  NANDN U25036 ( .A(n21350), .B(n21349), .Z(n21352) );
  NAND U25037 ( .A(n21352), .B(n21351), .Z(n21354) );
  NAND U25038 ( .A(n21354), .B(n21353), .Z(n21356) );
  NAND U25039 ( .A(n21356), .B(n21355), .Z(n21358) );
  NAND U25040 ( .A(n21358), .B(n21357), .Z(n21359) );
  AND U25041 ( .A(n21360), .B(n21359), .Z(n21361) );
  OR U25042 ( .A(n21362), .B(n21361), .Z(n21363) );
  NANDN U25043 ( .A(n21364), .B(n21363), .Z(n21366) );
  NAND U25044 ( .A(n21366), .B(n21365), .Z(n21368) );
  NAND U25045 ( .A(n21368), .B(n21367), .Z(n21369) );
  NANDN U25046 ( .A(n21370), .B(n21369), .Z(n21372) );
  NAND U25047 ( .A(n21372), .B(n21371), .Z(n21373) );
  NANDN U25048 ( .A(n21374), .B(n21373), .Z(n21376) );
  NAND U25049 ( .A(n21376), .B(n21375), .Z(n21378) );
  ANDN U25050 ( .B(n21378), .A(n21377), .Z(n21380) );
  NANDN U25051 ( .A(n21380), .B(n21379), .Z(n21381) );
  NANDN U25052 ( .A(n21382), .B(n21381), .Z(n21384) );
  NAND U25053 ( .A(n21384), .B(n21383), .Z(n21385) );
  NANDN U25054 ( .A(n21386), .B(n21385), .Z(n21388) );
  NAND U25055 ( .A(n21388), .B(n21387), .Z(n21390) );
  ANDN U25056 ( .B(n21390), .A(n21389), .Z(n21392) );
  NANDN U25057 ( .A(n21392), .B(n21391), .Z(n21393) );
  NANDN U25058 ( .A(n21394), .B(n21393), .Z(n21396) );
  NAND U25059 ( .A(n21396), .B(n21395), .Z(n21398) );
  NAND U25060 ( .A(n21398), .B(n21397), .Z(n21399) );
  NANDN U25061 ( .A(n21400), .B(n21399), .Z(n21402) );
  ANDN U25062 ( .B(n21402), .A(n21401), .Z(n21404) );
  NANDN U25063 ( .A(n21404), .B(n21403), .Z(n21405) );
  NANDN U25064 ( .A(n21406), .B(n21405), .Z(n21408) );
  NAND U25065 ( .A(n21408), .B(n21407), .Z(n21409) );
  NANDN U25066 ( .A(n21410), .B(n21409), .Z(n21412) );
  NAND U25067 ( .A(n21412), .B(n21411), .Z(n21414) );
  ANDN U25068 ( .B(n21414), .A(n21413), .Z(n21416) );
  NANDN U25069 ( .A(n21416), .B(n21415), .Z(n21417) );
  NANDN U25070 ( .A(n21418), .B(n21417), .Z(n21420) );
  NAND U25071 ( .A(n21420), .B(n21419), .Z(n21421) );
  NANDN U25072 ( .A(n21422), .B(n21421), .Z(n21424) );
  NAND U25073 ( .A(n21424), .B(n21423), .Z(n21426) );
  ANDN U25074 ( .B(n21426), .A(n21425), .Z(n21428) );
  NANDN U25075 ( .A(n21428), .B(n21427), .Z(n21429) );
  NANDN U25076 ( .A(n21430), .B(n21429), .Z(n21431) );
  NANDN U25077 ( .A(n21432), .B(n21431), .Z(n21433) );
  NANDN U25078 ( .A(n21434), .B(n21433), .Z(n21436) );
  NAND U25079 ( .A(n21436), .B(n21435), .Z(n21438) );
  ANDN U25080 ( .B(n21438), .A(n21437), .Z(n21440) );
  NANDN U25081 ( .A(n21440), .B(n21439), .Z(n21441) );
  NANDN U25082 ( .A(n21442), .B(n21441), .Z(n21444) );
  NAND U25083 ( .A(n21444), .B(n21443), .Z(n21445) );
  NANDN U25084 ( .A(n21446), .B(n21445), .Z(n21447) );
  NANDN U25085 ( .A(n21448), .B(n21447), .Z(n21449) );
  AND U25086 ( .A(n21450), .B(n21449), .Z(n21452) );
  NANDN U25087 ( .A(n21452), .B(n21451), .Z(n21454) );
  NAND U25088 ( .A(n21454), .B(n21453), .Z(n21456) );
  NAND U25089 ( .A(n21456), .B(n21455), .Z(n21458) );
  NAND U25090 ( .A(n21458), .B(n21457), .Z(n21460) );
  NAND U25091 ( .A(n21460), .B(n21459), .Z(n21461) );
  AND U25092 ( .A(n21462), .B(n21461), .Z(n21466) );
  AND U25093 ( .A(n21464), .B(n21463), .Z(n21465) );
  NANDN U25094 ( .A(n21466), .B(n21465), .Z(n21468) );
  ANDN U25095 ( .B(n21468), .A(n21467), .Z(n21469) );
  ANDN U25096 ( .B(n21470), .A(n21469), .Z(n21472) );
  NAND U25097 ( .A(n21472), .B(n21471), .Z(n21474) );
  NAND U25098 ( .A(n21474), .B(n21473), .Z(n21475) );
  AND U25099 ( .A(n21476), .B(n21475), .Z(n21477) );
  OR U25100 ( .A(n21478), .B(n21477), .Z(n21479) );
  NANDN U25101 ( .A(n21480), .B(n21479), .Z(n21481) );
  NANDN U25102 ( .A(n21482), .B(n21481), .Z(n21483) );
  NANDN U25103 ( .A(n21484), .B(n21483), .Z(n21485) );
  NANDN U25104 ( .A(n21486), .B(n21485), .Z(n21488) );
  NAND U25105 ( .A(n21488), .B(n21487), .Z(n21489) );
  NANDN U25106 ( .A(n21490), .B(n21489), .Z(n21492) );
  NAND U25107 ( .A(n21492), .B(n21491), .Z(n21493) );
  AND U25108 ( .A(n21494), .B(n21493), .Z(n21496) );
  NANDN U25109 ( .A(n21496), .B(n21495), .Z(n21497) );
  NANDN U25110 ( .A(n21498), .B(n21497), .Z(n21500) );
  NAND U25111 ( .A(n21500), .B(n21499), .Z(n21501) );
  NANDN U25112 ( .A(n21502), .B(n21501), .Z(n21504) );
  NAND U25113 ( .A(n21504), .B(n21503), .Z(n21505) );
  AND U25114 ( .A(n21506), .B(n21505), .Z(n21508) );
  NANDN U25115 ( .A(n21508), .B(n21507), .Z(n21509) );
  NANDN U25116 ( .A(n21510), .B(n21509), .Z(n21512) );
  NAND U25117 ( .A(n21512), .B(n21511), .Z(n21513) );
  NANDN U25118 ( .A(n21514), .B(n21513), .Z(n21516) );
  NAND U25119 ( .A(n21516), .B(n21515), .Z(n21518) );
  ANDN U25120 ( .B(n21518), .A(n21517), .Z(n21522) );
  ANDN U25121 ( .B(n21520), .A(n21519), .Z(n21521) );
  NANDN U25122 ( .A(n21522), .B(n21521), .Z(n21524) );
  NAND U25123 ( .A(n21524), .B(n21523), .Z(n21525) );
  OR U25124 ( .A(n21525), .B(x[883]), .Z(n21528) );
  XOR U25125 ( .A(n21525), .B(x[883]), .Z(n21526) );
  NAND U25126 ( .A(y[883]), .B(n21526), .Z(n21527) );
  NAND U25127 ( .A(n21528), .B(n21527), .Z(n21529) );
  AND U25128 ( .A(n21530), .B(n21529), .Z(n21532) );
  NANDN U25129 ( .A(n21532), .B(n21531), .Z(n21533) );
  NANDN U25130 ( .A(n21534), .B(n21533), .Z(n21536) );
  NAND U25131 ( .A(n21536), .B(n21535), .Z(n21538) );
  NAND U25132 ( .A(n21538), .B(n21537), .Z(n21540) );
  NAND U25133 ( .A(n21540), .B(n21539), .Z(n21542) );
  ANDN U25134 ( .B(n21542), .A(n21541), .Z(n21544) );
  NANDN U25135 ( .A(n21544), .B(n21543), .Z(n21545) );
  NANDN U25136 ( .A(n21546), .B(n21545), .Z(n21548) );
  NAND U25137 ( .A(n21548), .B(n21547), .Z(n21549) );
  NANDN U25138 ( .A(n21550), .B(n21549), .Z(n21551) );
  AND U25139 ( .A(n21552), .B(n21551), .Z(n21554) );
  NAND U25140 ( .A(n21554), .B(n21553), .Z(n21556) );
  NAND U25141 ( .A(n21556), .B(n21555), .Z(n21558) );
  NAND U25142 ( .A(n21558), .B(n21557), .Z(n21560) );
  ANDN U25143 ( .B(n21560), .A(n21559), .Z(n21562) );
  NANDN U25144 ( .A(n21562), .B(n21561), .Z(n21563) );
  NANDN U25145 ( .A(n21564), .B(n21563), .Z(n21566) );
  NAND U25146 ( .A(n21566), .B(n21565), .Z(n21568) );
  NAND U25147 ( .A(n21568), .B(n21567), .Z(n21570) );
  NAND U25148 ( .A(n21570), .B(n21569), .Z(n21571) );
  AND U25149 ( .A(n21572), .B(n21571), .Z(n21574) );
  NANDN U25150 ( .A(n21574), .B(n21573), .Z(n21576) );
  NAND U25151 ( .A(n21576), .B(n21575), .Z(n21578) );
  NAND U25152 ( .A(n21578), .B(n21577), .Z(n21580) );
  NAND U25153 ( .A(n21580), .B(n21579), .Z(n21581) );
  AND U25154 ( .A(n21582), .B(n21581), .Z(n21584) );
  NAND U25155 ( .A(n21584), .B(n21583), .Z(n21586) );
  NAND U25156 ( .A(n21586), .B(n21585), .Z(n21588) );
  NANDN U25157 ( .A(n21588), .B(y[907]), .Z(n21591) );
  XOR U25158 ( .A(n21588), .B(n21587), .Z(n21589) );
  NANDN U25159 ( .A(x[907]), .B(n21589), .Z(n21590) );
  AND U25160 ( .A(n21591), .B(n21590), .Z(n21594) );
  NANDN U25161 ( .A(n21594), .B(n21595), .Z(n21592) );
  AND U25162 ( .A(n21593), .B(n21592), .Z(n21598) );
  XNOR U25163 ( .A(n21595), .B(n21594), .Z(n21596) );
  NAND U25164 ( .A(n21596), .B(y[908]), .Z(n21597) );
  NAND U25165 ( .A(n21598), .B(n21597), .Z(n21600) );
  NAND U25166 ( .A(n21600), .B(n21599), .Z(n21602) );
  NAND U25167 ( .A(n21602), .B(n21601), .Z(n21603) );
  AND U25168 ( .A(n21604), .B(n21603), .Z(n21606) );
  NANDN U25169 ( .A(n21606), .B(n21605), .Z(n21608) );
  NAND U25170 ( .A(n21608), .B(n21607), .Z(n21610) );
  NAND U25171 ( .A(n21610), .B(n21609), .Z(n21612) );
  NAND U25172 ( .A(n21612), .B(n21611), .Z(n21614) );
  NAND U25173 ( .A(n21614), .B(n21613), .Z(n21615) );
  AND U25174 ( .A(n21616), .B(n21615), .Z(n21618) );
  NANDN U25175 ( .A(n21618), .B(n21617), .Z(n21620) );
  NAND U25176 ( .A(n21620), .B(n21619), .Z(n21622) );
  NAND U25177 ( .A(n21622), .B(n21621), .Z(n21624) );
  NAND U25178 ( .A(n21624), .B(n21623), .Z(n21625) );
  NANDN U25179 ( .A(n21626), .B(n21625), .Z(n21628) );
  ANDN U25180 ( .B(n21628), .A(n21627), .Z(n21630) );
  NANDN U25181 ( .A(n21630), .B(n21629), .Z(n21632) );
  NAND U25182 ( .A(n21632), .B(n21631), .Z(n21634) );
  NAND U25183 ( .A(n21634), .B(n21633), .Z(n21636) );
  NAND U25184 ( .A(n21636), .B(n21635), .Z(n21638) );
  NAND U25185 ( .A(n21638), .B(n21637), .Z(n21639) );
  AND U25186 ( .A(n21640), .B(n21639), .Z(n21642) );
  NANDN U25187 ( .A(n21642), .B(n21641), .Z(n21644) );
  NAND U25188 ( .A(n21644), .B(n21643), .Z(n21646) );
  NAND U25189 ( .A(n21646), .B(n21645), .Z(n21648) );
  NANDN U25190 ( .A(n21648), .B(n21647), .Z(n21650) );
  NAND U25191 ( .A(n21650), .B(n21649), .Z(n21652) );
  NANDN U25192 ( .A(n21652), .B(y[931]), .Z(n21655) );
  XOR U25193 ( .A(n21652), .B(n21651), .Z(n21653) );
  NANDN U25194 ( .A(x[931]), .B(n21653), .Z(n21654) );
  AND U25195 ( .A(n21655), .B(n21654), .Z(n21658) );
  OR U25196 ( .A(n21658), .B(x[932]), .Z(n21656) );
  AND U25197 ( .A(n21657), .B(n21656), .Z(n21661) );
  XOR U25198 ( .A(x[932]), .B(n21658), .Z(n21659) );
  NAND U25199 ( .A(n21659), .B(y[932]), .Z(n21660) );
  NAND U25200 ( .A(n21661), .B(n21660), .Z(n21663) );
  NAND U25201 ( .A(n21663), .B(n21662), .Z(n21665) );
  NAND U25202 ( .A(n21665), .B(n21664), .Z(n21666) );
  AND U25203 ( .A(n21667), .B(n21666), .Z(n21669) );
  NANDN U25204 ( .A(n21669), .B(n21668), .Z(n21671) );
  NAND U25205 ( .A(n21671), .B(n21670), .Z(n21673) );
  NAND U25206 ( .A(n21673), .B(n21672), .Z(n21675) );
  NAND U25207 ( .A(n21675), .B(n21674), .Z(n21677) );
  NAND U25208 ( .A(n21677), .B(n21676), .Z(n21678) );
  AND U25209 ( .A(n21679), .B(n21678), .Z(n21683) );
  ANDN U25210 ( .B(n21681), .A(n21680), .Z(n21682) );
  NANDN U25211 ( .A(n21683), .B(n21682), .Z(n21684) );
  AND U25212 ( .A(n21685), .B(n21684), .Z(n21686) );
  ANDN U25213 ( .B(n21687), .A(n21686), .Z(n21689) );
  NAND U25214 ( .A(n21689), .B(n21688), .Z(n21690) );
  NANDN U25215 ( .A(n21691), .B(n21690), .Z(n21693) );
  NAND U25216 ( .A(n21693), .B(n21692), .Z(n21694) );
  AND U25217 ( .A(n21695), .B(n21694), .Z(n21697) );
  NANDN U25218 ( .A(n21697), .B(n21696), .Z(n21699) );
  NAND U25219 ( .A(n21699), .B(n21698), .Z(n21701) );
  NAND U25220 ( .A(n21701), .B(n21700), .Z(n21703) );
  NAND U25221 ( .A(n21703), .B(n21702), .Z(n21705) );
  NAND U25222 ( .A(n21705), .B(n21704), .Z(n21706) );
  AND U25223 ( .A(n21707), .B(n21706), .Z(n21711) );
  ANDN U25224 ( .B(n21709), .A(n21708), .Z(n21710) );
  NANDN U25225 ( .A(n21711), .B(n21710), .Z(n21712) );
  AND U25226 ( .A(n21713), .B(n21712), .Z(n21717) );
  ANDN U25227 ( .B(n21715), .A(n21714), .Z(n21716) );
  NANDN U25228 ( .A(n21717), .B(n21716), .Z(n21719) );
  ANDN U25229 ( .B(n21719), .A(n21718), .Z(n21721) );
  NANDN U25230 ( .A(n21721), .B(n21720), .Z(n21723) );
  ANDN U25231 ( .B(n21723), .A(n21722), .Z(n21724) );
  OR U25232 ( .A(n21725), .B(n21724), .Z(n21726) );
  NANDN U25233 ( .A(n21727), .B(n21726), .Z(n21729) );
  NAND U25234 ( .A(n21729), .B(n21728), .Z(n21730) );
  NANDN U25235 ( .A(n21731), .B(n21730), .Z(n21733) );
  NAND U25236 ( .A(n21733), .B(n21732), .Z(n21735) );
  ANDN U25237 ( .B(n21735), .A(n21734), .Z(n21737) );
  NANDN U25238 ( .A(n21737), .B(n21736), .Z(n21739) );
  NAND U25239 ( .A(n21739), .B(n21738), .Z(n21741) );
  NAND U25240 ( .A(n21741), .B(n21740), .Z(n21742) );
  NANDN U25241 ( .A(n21743), .B(n21742), .Z(n21745) );
  NAND U25242 ( .A(n21745), .B(n21744), .Z(n21747) );
  ANDN U25243 ( .B(n21747), .A(n21746), .Z(n21749) );
  NANDN U25244 ( .A(n21749), .B(n21748), .Z(n21751) );
  NAND U25245 ( .A(n21751), .B(n21750), .Z(n21753) );
  NAND U25246 ( .A(n21753), .B(n21752), .Z(n21754) );
  NANDN U25247 ( .A(n21755), .B(n21754), .Z(n21757) );
  NAND U25248 ( .A(n21757), .B(n21756), .Z(n21759) );
  ANDN U25249 ( .B(n21759), .A(n21758), .Z(n21761) );
  NANDN U25250 ( .A(n21761), .B(n21760), .Z(n21762) );
  NANDN U25251 ( .A(n21763), .B(n21762), .Z(n21765) );
  NAND U25252 ( .A(n21765), .B(n21764), .Z(n21767) );
  NAND U25253 ( .A(n21767), .B(n21766), .Z(n21769) );
  NAND U25254 ( .A(n21769), .B(n21768), .Z(n21771) );
  ANDN U25255 ( .B(n21771), .A(n21770), .Z(n21773) );
  NANDN U25256 ( .A(n21773), .B(n21772), .Z(n21774) );
  NANDN U25257 ( .A(n21775), .B(n21774), .Z(n21777) );
  NAND U25258 ( .A(n21777), .B(n21776), .Z(n21779) );
  NAND U25259 ( .A(n21779), .B(n21778), .Z(n21781) );
  NAND U25260 ( .A(n21781), .B(n21780), .Z(n21783) );
  ANDN U25261 ( .B(n21783), .A(n21782), .Z(n21785) );
  NANDN U25262 ( .A(n21785), .B(n21784), .Z(n21786) );
  NANDN U25263 ( .A(n21787), .B(n21786), .Z(n21789) );
  NAND U25264 ( .A(n21789), .B(n21788), .Z(n21790) );
  NANDN U25265 ( .A(n21791), .B(n21790), .Z(n21792) );
  AND U25266 ( .A(n21793), .B(n21792), .Z(n21795) );
  NAND U25267 ( .A(n21795), .B(n21794), .Z(n21797) );
  NAND U25268 ( .A(n21797), .B(n21796), .Z(n21798) );
  AND U25269 ( .A(n21799), .B(n21798), .Z(n21800) );
  NANDN U25270 ( .A(n21801), .B(n21800), .Z(n21802) );
  NANDN U25271 ( .A(n21803), .B(n21802), .Z(n21805) );
  NAND U25272 ( .A(n21805), .B(n21804), .Z(n21806) );
  AND U25273 ( .A(n21807), .B(n21806), .Z(n21809) );
  NANDN U25274 ( .A(n21809), .B(n21808), .Z(n21811) );
  NAND U25275 ( .A(n21811), .B(n21810), .Z(n21813) );
  NAND U25276 ( .A(n21813), .B(n21812), .Z(n21815) );
  NAND U25277 ( .A(n21815), .B(n21814), .Z(n21817) );
  NAND U25278 ( .A(n21817), .B(n21816), .Z(n21818) );
  AND U25279 ( .A(n21819), .B(n21818), .Z(n21823) );
  AND U25280 ( .A(n21821), .B(n21820), .Z(n21822) );
  NANDN U25281 ( .A(n21823), .B(n21822), .Z(n21825) );
  ANDN U25282 ( .B(n21825), .A(n21824), .Z(n21826) );
  ANDN U25283 ( .B(n21827), .A(n21826), .Z(n21829) );
  NAND U25284 ( .A(n21829), .B(n21828), .Z(n21831) );
  NAND U25285 ( .A(n21831), .B(n21830), .Z(n21833) );
  NAND U25286 ( .A(n21833), .B(n21832), .Z(n21834) );
  AND U25287 ( .A(n21835), .B(n21834), .Z(n21837) );
  NANDN U25288 ( .A(n21837), .B(n21836), .Z(n21839) );
  NAND U25289 ( .A(n21839), .B(n21838), .Z(n21841) );
  NAND U25290 ( .A(n21841), .B(n21840), .Z(n21843) );
  NAND U25291 ( .A(n21843), .B(n21842), .Z(n21845) );
  NAND U25292 ( .A(n21845), .B(n21844), .Z(n21846) );
  AND U25293 ( .A(n21847), .B(n21846), .Z(n21851) );
  AND U25294 ( .A(n21849), .B(n21848), .Z(n21850) );
  NANDN U25295 ( .A(n21851), .B(n21850), .Z(n21852) );
  AND U25296 ( .A(n21853), .B(n21852), .Z(n21854) );
  ANDN U25297 ( .B(n21855), .A(n21854), .Z(n21857) );
  NAND U25298 ( .A(n21857), .B(n21856), .Z(n21859) );
  ANDN U25299 ( .B(n21859), .A(n21858), .Z(n21861) );
  NANDN U25300 ( .A(n21861), .B(n21860), .Z(n21863) );
  NAND U25301 ( .A(n21863), .B(n21862), .Z(n21865) );
  NAND U25302 ( .A(n21865), .B(n21864), .Z(n21866) );
  NANDN U25303 ( .A(n21867), .B(n21866), .Z(n21869) );
  NAND U25304 ( .A(n21869), .B(n21868), .Z(n21870) );
  AND U25305 ( .A(n21871), .B(n21870), .Z(n21873) );
  NANDN U25306 ( .A(n21873), .B(n21872), .Z(n21875) );
  NAND U25307 ( .A(n21875), .B(n21874), .Z(n21877) );
  NAND U25308 ( .A(n21877), .B(n21876), .Z(n21878) );
  NANDN U25309 ( .A(n21879), .B(n21878), .Z(n21881) );
  NAND U25310 ( .A(n21881), .B(n21880), .Z(n21882) );
  AND U25311 ( .A(n21883), .B(n21882), .Z(n21885) );
  NANDN U25312 ( .A(n21885), .B(n21884), .Z(n21887) );
  NAND U25313 ( .A(n21887), .B(n21886), .Z(n21889) );
  NAND U25314 ( .A(n21889), .B(n21888), .Z(n21890) );
  NANDN U25315 ( .A(n21891), .B(n21890), .Z(n21893) );
  NAND U25316 ( .A(n21893), .B(n21892), .Z(n21895) );
  ANDN U25317 ( .B(n21895), .A(n21894), .Z(n21896) );
  OR U25318 ( .A(n21897), .B(n21896), .Z(n21899) );
  NAND U25319 ( .A(n21899), .B(n21898), .Z(n21901) );
  NAND U25320 ( .A(n21901), .B(n21900), .Z(n21903) );
  NAND U25321 ( .A(n21903), .B(n21902), .Z(n21905) );
  NAND U25322 ( .A(n21905), .B(n21904), .Z(n21907) );
  ANDN U25323 ( .B(n21907), .A(n21906), .Z(n21909) );
  NANDN U25324 ( .A(n21909), .B(n21908), .Z(n21910) );
  NANDN U25325 ( .A(n21911), .B(n21910), .Z(n21913) );
  NAND U25326 ( .A(n21913), .B(n21912), .Z(n21915) );
  NAND U25327 ( .A(n21915), .B(n21914), .Z(n21917) );
  NAND U25328 ( .A(n21917), .B(n21916), .Z(n21918) );
  AND U25329 ( .A(n21919), .B(n21918), .Z(n21921) );
  NANDN U25330 ( .A(n21921), .B(n21920), .Z(n21922) );
  NANDN U25331 ( .A(n21923), .B(n21922), .Z(n21925) );
  NAND U25332 ( .A(n21925), .B(n21924), .Z(n21926) );
  NANDN U25333 ( .A(n21927), .B(n21926), .Z(n21928) );
  NANDN U25334 ( .A(n21929), .B(n21928), .Z(n21930) );
  NANDN U25335 ( .A(n21931), .B(n21930), .Z(n21933) );
  NAND U25336 ( .A(n21933), .B(n21932), .Z(n21935) );
  NAND U25337 ( .A(n21935), .B(n21934), .Z(n21936) );
  AND U25338 ( .A(n21937), .B(n21936), .Z(n21939) );
  NANDN U25339 ( .A(n21939), .B(n21938), .Z(n21940) );
  NANDN U25340 ( .A(n21941), .B(n21940), .Z(n21942) );
  NANDN U25341 ( .A(n21943), .B(n21942), .Z(n21945) );
  NAND U25342 ( .A(n21945), .B(n21944), .Z(n21947) );
  NAND U25343 ( .A(n21947), .B(n21946), .Z(n21948) );
  AND U25344 ( .A(n21949), .B(n21948), .Z(n21950) );
  OR U25345 ( .A(n21951), .B(n21950), .Z(n21952) );
  NANDN U25346 ( .A(n21953), .B(n21952), .Z(n21955) );
  ANDN U25347 ( .B(n21955), .A(n21954), .Z(n21957) );
  NANDN U25348 ( .A(n21957), .B(n21956), .Z(n21958) );
  AND U25349 ( .A(n21959), .B(n21958), .Z(n21960) );
  OR U25350 ( .A(n21961), .B(n21960), .Z(n21963) );
  NAND U25351 ( .A(n21963), .B(n21962), .Z(n21965) );
  NAND U25352 ( .A(n21965), .B(n21964), .Z(n21967) );
  NAND U25353 ( .A(n21967), .B(n21966), .Z(n21969) );
  NAND U25354 ( .A(n21969), .B(n21968), .Z(n21970) );
  AND U25355 ( .A(n21971), .B(n21970), .Z(n21973) );
  NANDN U25356 ( .A(n21973), .B(n21972), .Z(n21975) );
  NAND U25357 ( .A(n21975), .B(n21974), .Z(n21976) );
  NANDN U25358 ( .A(n21977), .B(n21976), .Z(n21978) );
  NANDN U25359 ( .A(n21979), .B(n21978), .Z(n21981) );
  NAND U25360 ( .A(n21981), .B(n21980), .Z(n21983) );
  NAND U25361 ( .A(n21983), .B(n21982), .Z(n21984) );
  NANDN U25362 ( .A(n21985), .B(n21984), .Z(n21987) );
  NAND U25363 ( .A(n21987), .B(n21986), .Z(n21988) );
  AND U25364 ( .A(n21989), .B(n21988), .Z(n21991) );
  NANDN U25365 ( .A(n21991), .B(n21990), .Z(n21992) );
  NANDN U25366 ( .A(n21993), .B(n21992), .Z(n21995) );
  NAND U25367 ( .A(n21995), .B(n21994), .Z(n21996) );
  NANDN U25368 ( .A(n21997), .B(n21996), .Z(n21999) );
  NAND U25369 ( .A(n21999), .B(n21998), .Z(n22001) );
  ANDN U25370 ( .B(n22001), .A(n22000), .Z(n22003) );
  NANDN U25371 ( .A(n22003), .B(n22002), .Z(n22004) );
  NANDN U25372 ( .A(n22005), .B(n22004), .Z(n22006) );
  NANDN U25373 ( .A(n22007), .B(n22006), .Z(n22008) );
  NANDN U25374 ( .A(n22009), .B(n22008), .Z(n22011) );
  NAND U25375 ( .A(n22011), .B(n22010), .Z(n22012) );
  AND U25376 ( .A(n22013), .B(n22012), .Z(n22015) );
  NANDN U25377 ( .A(n22015), .B(n22014), .Z(n22017) );
  NAND U25378 ( .A(n22017), .B(n22016), .Z(n22019) );
  NAND U25379 ( .A(n22019), .B(n22018), .Z(n22021) );
  NAND U25380 ( .A(n22021), .B(n22020), .Z(n22023) );
  NAND U25381 ( .A(n22023), .B(n22022), .Z(n22025) );
  ANDN U25382 ( .B(n22025), .A(n22024), .Z(n22026) );
  OR U25383 ( .A(n22027), .B(n22026), .Z(n22029) );
  NAND U25384 ( .A(n22029), .B(n22028), .Z(n22031) );
  NAND U25385 ( .A(n22031), .B(n22030), .Z(n22033) );
  NAND U25386 ( .A(n22033), .B(n22032), .Z(n22035) );
  NAND U25387 ( .A(n22035), .B(n22034), .Z(n22037) );
  ANDN U25388 ( .B(n22037), .A(n22036), .Z(n22038) );
  OR U25389 ( .A(n22039), .B(n22038), .Z(n22041) );
  NAND U25390 ( .A(n22041), .B(n22040), .Z(n22043) );
  NAND U25391 ( .A(n22043), .B(n22042), .Z(n22045) );
  NAND U25392 ( .A(n22045), .B(n22044), .Z(n22047) );
  NAND U25393 ( .A(n22047), .B(n22046), .Z(n22048) );
  AND U25394 ( .A(n22049), .B(n22048), .Z(n22051) );
  NAND U25395 ( .A(n22051), .B(n22050), .Z(n22052) );
  NANDN U25396 ( .A(n22053), .B(n22052), .Z(n22055) );
  NAND U25397 ( .A(n22055), .B(n22054), .Z(n22056) );
  NANDN U25398 ( .A(n22057), .B(n22056), .Z(n22058) );
  NANDN U25399 ( .A(n22059), .B(n22058), .Z(n22061) );
  ANDN U25400 ( .B(n22061), .A(n22060), .Z(n22063) );
  NANDN U25401 ( .A(n22063), .B(n22062), .Z(n22064) );
  NANDN U25402 ( .A(n22065), .B(n22064), .Z(n22067) );
  NAND U25403 ( .A(n22067), .B(n22066), .Z(n22068) );
  NANDN U25404 ( .A(n22069), .B(n22068), .Z(n22071) );
  NAND U25405 ( .A(n22071), .B(n22070), .Z(n22073) );
  ANDN U25406 ( .B(n22073), .A(n22072), .Z(n22075) );
  NANDN U25407 ( .A(n22075), .B(n22074), .Z(n22076) );
  NANDN U25408 ( .A(n22077), .B(n22076), .Z(n22079) );
  NAND U25409 ( .A(n22079), .B(n22078), .Z(n22081) );
  NAND U25410 ( .A(n22081), .B(n22080), .Z(n22083) );
  NAND U25411 ( .A(n22083), .B(n22082), .Z(n22085) );
  ANDN U25412 ( .B(n22085), .A(n22084), .Z(n22087) );
  NANDN U25413 ( .A(n22087), .B(n22086), .Z(n22088) );
  NANDN U25414 ( .A(n22089), .B(n22088), .Z(n22091) );
  NAND U25415 ( .A(n22091), .B(n22090), .Z(n22092) );
  NANDN U25416 ( .A(n22093), .B(n22092), .Z(n22095) );
  NAND U25417 ( .A(n22095), .B(n22094), .Z(n22097) );
  ANDN U25418 ( .B(n22097), .A(n22096), .Z(n22099) );
  NANDN U25419 ( .A(n22099), .B(n22098), .Z(n22101) );
  ANDN U25420 ( .B(n22101), .A(n22100), .Z(n22103) );
  NANDN U25421 ( .A(n22103), .B(n22102), .Z(n22105) );
  NAND U25422 ( .A(n22105), .B(n22104), .Z(n22107) );
  NAND U25423 ( .A(n22107), .B(n22106), .Z(n22109) );
  NAND U25424 ( .A(n22109), .B(n22108), .Z(n22111) );
  NAND U25425 ( .A(n22111), .B(n22110), .Z(n22112) );
  AND U25426 ( .A(n22113), .B(n22112), .Z(n22115) );
  NANDN U25427 ( .A(n22115), .B(n22114), .Z(n22116) );
  NANDN U25428 ( .A(n22117), .B(n22116), .Z(n22119) );
  NAND U25429 ( .A(n22119), .B(n22118), .Z(n22121) );
  NAND U25430 ( .A(n22121), .B(n22120), .Z(n22123) );
  NAND U25431 ( .A(n22123), .B(n22122), .Z(n22124) );
  AND U25432 ( .A(n22125), .B(n22124), .Z(n22127) );
  NANDN U25433 ( .A(n22127), .B(n22126), .Z(n22129) );
  NAND U25434 ( .A(n22129), .B(n22128), .Z(n22131) );
  NAND U25435 ( .A(n22131), .B(n22130), .Z(n22132) );
  NANDN U25436 ( .A(n22133), .B(n22132), .Z(n22134) );
  NANDN U25437 ( .A(n22135), .B(n22134), .Z(n22137) );
  ANDN U25438 ( .B(n22137), .A(n22136), .Z(n22138) );
  OR U25439 ( .A(n22139), .B(n22138), .Z(n22140) );
  NANDN U25440 ( .A(n22141), .B(n22140), .Z(n22143) );
  NAND U25441 ( .A(n22143), .B(n22142), .Z(n22144) );
  NANDN U25442 ( .A(n22145), .B(n22144), .Z(n22147) );
  NAND U25443 ( .A(n22147), .B(n22146), .Z(n22149) );
  ANDN U25444 ( .B(n22149), .A(n22148), .Z(n22151) );
  NANDN U25445 ( .A(n22151), .B(n22150), .Z(n22152) );
  NANDN U25446 ( .A(n22153), .B(n22152), .Z(n22154) );
  NANDN U25447 ( .A(n22155), .B(n22154), .Z(n22156) );
  NANDN U25448 ( .A(n22157), .B(n22156), .Z(n22159) );
  NAND U25449 ( .A(n22159), .B(n22158), .Z(n22161) );
  ANDN U25450 ( .B(n22161), .A(n22160), .Z(n22163) );
  NANDN U25451 ( .A(n22163), .B(n22162), .Z(n22164) );
  NANDN U25452 ( .A(n22165), .B(n22164), .Z(n22167) );
  NAND U25453 ( .A(n22167), .B(n22166), .Z(n22168) );
  NANDN U25454 ( .A(n22169), .B(n22168), .Z(n22171) );
  NAND U25455 ( .A(n22171), .B(n22170), .Z(n22173) );
  ANDN U25456 ( .B(n22173), .A(n22172), .Z(n22177) );
  ANDN U25457 ( .B(n22175), .A(n22174), .Z(n22176) );
  NANDN U25458 ( .A(n22177), .B(n22176), .Z(n22179) );
  ANDN U25459 ( .B(n22179), .A(n22178), .Z(n22181) );
  NANDN U25460 ( .A(n22181), .B(n22180), .Z(n22182) );
  NANDN U25461 ( .A(n22183), .B(n22182), .Z(n22185) );
  NAND U25462 ( .A(n22185), .B(n22184), .Z(n22186) );
  NANDN U25463 ( .A(n22187), .B(n22186), .Z(n22189) );
  NAND U25464 ( .A(n22189), .B(n22188), .Z(n22191) );
  ANDN U25465 ( .B(n22191), .A(n22190), .Z(n22193) );
  NANDN U25466 ( .A(n22193), .B(n22192), .Z(n22194) );
  NANDN U25467 ( .A(n22195), .B(n22194), .Z(n22197) );
  NAND U25468 ( .A(n22197), .B(n22196), .Z(n22199) );
  NAND U25469 ( .A(n22199), .B(n22198), .Z(n22201) );
  NAND U25470 ( .A(n22201), .B(n22200), .Z(n22202) );
  AND U25471 ( .A(n22203), .B(n22202), .Z(n22205) );
  NANDN U25472 ( .A(n22205), .B(n22204), .Z(n22206) );
  NANDN U25473 ( .A(n22207), .B(n22206), .Z(n22209) );
  NAND U25474 ( .A(n22209), .B(n22208), .Z(n22210) );
  NANDN U25475 ( .A(n22211), .B(n22210), .Z(n22212) );
  NANDN U25476 ( .A(n22213), .B(n22212), .Z(n22215) );
  NAND U25477 ( .A(n22215), .B(n22214), .Z(n22216) );
  NANDN U25478 ( .A(n22217), .B(n22216), .Z(n22219) );
  NAND U25479 ( .A(n22219), .B(n22218), .Z(n22221) );
  ANDN U25480 ( .B(n22221), .A(n22220), .Z(n22223) );
  NANDN U25481 ( .A(n22223), .B(n22222), .Z(n22224) );
  AND U25482 ( .A(n22225), .B(n22224), .Z(n22227) );
  NANDN U25483 ( .A(n22227), .B(n22226), .Z(n22228) );
  NANDN U25484 ( .A(n22229), .B(n22228), .Z(n22231) );
  NAND U25485 ( .A(n22231), .B(n22230), .Z(n22233) );
  ANDN U25486 ( .B(n22233), .A(n22232), .Z(n22235) );
  NANDN U25487 ( .A(n22235), .B(n22234), .Z(n22237) );
  NAND U25488 ( .A(n22237), .B(n22236), .Z(n22238) );
  AND U25489 ( .A(n22239), .B(n22238), .Z(n22241) );
  NANDN U25490 ( .A(n22241), .B(n22240), .Z(n22242) );
  NANDN U25491 ( .A(n22243), .B(n22242), .Z(n22245) );
  NAND U25492 ( .A(n22245), .B(n22244), .Z(n22247) );
  NAND U25493 ( .A(n22247), .B(n22246), .Z(n22249) );
  NAND U25494 ( .A(n22249), .B(n22248), .Z(n22250) );
  AND U25495 ( .A(n22251), .B(n22250), .Z(n22253) );
  NANDN U25496 ( .A(n22253), .B(n22252), .Z(n22254) );
  AND U25497 ( .A(n22255), .B(n22254), .Z(n22257) );
  NANDN U25498 ( .A(n22257), .B(n22256), .Z(n22258) );
  NANDN U25499 ( .A(n22259), .B(n22258), .Z(n22261) );
  ANDN U25500 ( .B(n22261), .A(n22260), .Z(n22263) );
  NANDN U25501 ( .A(n22263), .B(n22262), .Z(n22264) );
  NANDN U25502 ( .A(n22265), .B(n22264), .Z(n22267) );
  NAND U25503 ( .A(n22267), .B(n22266), .Z(n22269) );
  NAND U25504 ( .A(n22269), .B(n22268), .Z(n22270) );
  AND U25505 ( .A(n22271), .B(n22270), .Z(n22273) );
  NANDN U25506 ( .A(n22273), .B(n22272), .Z(n22274) );
  NANDN U25507 ( .A(n22275), .B(n22274), .Z(n22277) );
  NAND U25508 ( .A(n22277), .B(n22276), .Z(n22278) );
  NANDN U25509 ( .A(n22279), .B(n22278), .Z(n22281) );
  NAND U25510 ( .A(n22281), .B(n22280), .Z(n22282) );
  AND U25511 ( .A(n22283), .B(n22282), .Z(n22285) );
  NANDN U25512 ( .A(n22285), .B(n22284), .Z(n22287) );
  ANDN U25513 ( .B(n22287), .A(n22286), .Z(n22289) );
  NANDN U25514 ( .A(n22289), .B(n22288), .Z(n22290) );
  NANDN U25515 ( .A(n22291), .B(n22290), .Z(n22293) );
  NAND U25516 ( .A(n22293), .B(n22292), .Z(n22295) );
  NAND U25517 ( .A(n22295), .B(n22294), .Z(n22297) );
  NAND U25518 ( .A(n22297), .B(n22296), .Z(n22299) );
  NAND U25519 ( .A(n22299), .B(n22298), .Z(n22303) );
  NAND U25520 ( .A(n22301), .B(n22300), .Z(n22302) );
  AND U25521 ( .A(n22303), .B(n22302), .Z(n22305) );
  NAND U25522 ( .A(n22305), .B(n22304), .Z(n22306) );
  NANDN U25523 ( .A(n22307), .B(n22306), .Z(n22309) );
  ANDN U25524 ( .B(n22309), .A(n22308), .Z(n22310) );
  OR U25525 ( .A(n22311), .B(n22310), .Z(n22312) );
  NANDN U25526 ( .A(n22313), .B(n22312), .Z(n22315) );
  NAND U25527 ( .A(n22315), .B(n22314), .Z(n22316) );
  NANDN U25528 ( .A(n22317), .B(n22316), .Z(n22319) );
  NAND U25529 ( .A(n22319), .B(n22318), .Z(n22320) );
  AND U25530 ( .A(n22321), .B(n22320), .Z(n22322) );
  OR U25531 ( .A(n22323), .B(n22322), .Z(n22324) );
  NANDN U25532 ( .A(n22325), .B(n22324), .Z(n22326) );
  NANDN U25533 ( .A(n22327), .B(n22326), .Z(n22328) );
  NANDN U25534 ( .A(n22329), .B(n22328), .Z(n22331) );
  NAND U25535 ( .A(n22331), .B(n22330), .Z(n22333) );
  ANDN U25536 ( .B(n22333), .A(n22332), .Z(n22335) );
  NANDN U25537 ( .A(n22335), .B(n22334), .Z(n22336) );
  NANDN U25538 ( .A(n22337), .B(n22336), .Z(n22339) );
  NAND U25539 ( .A(n22339), .B(n22338), .Z(n22340) );
  NANDN U25540 ( .A(n22341), .B(n22340), .Z(n22343) );
  NAND U25541 ( .A(n22343), .B(n22342), .Z(n22344) );
  AND U25542 ( .A(n22345), .B(n22344), .Z(n22347) );
  NANDN U25543 ( .A(n22347), .B(n22346), .Z(n22349) );
  NAND U25544 ( .A(n22349), .B(n22348), .Z(n22351) );
  NAND U25545 ( .A(n22351), .B(n22350), .Z(n22353) );
  ANDN U25546 ( .B(n22353), .A(n22352), .Z(n22354) );
  OR U25547 ( .A(n22355), .B(n22354), .Z(n22356) );
  NANDN U25548 ( .A(n22357), .B(n22356), .Z(n22358) );
  NANDN U25549 ( .A(n22359), .B(n22358), .Z(n22360) );
  NANDN U25550 ( .A(n22361), .B(n22360), .Z(n22363) );
  NAND U25551 ( .A(n22363), .B(n22362), .Z(n22365) );
  ANDN U25552 ( .B(n22365), .A(n22364), .Z(n22367) );
  NANDN U25553 ( .A(n22367), .B(n22366), .Z(n22368) );
  NANDN U25554 ( .A(n22369), .B(n22368), .Z(n22370) );
  NANDN U25555 ( .A(n22371), .B(n22370), .Z(n22373) );
  NAND U25556 ( .A(n22373), .B(n22372), .Z(n22375) );
  NAND U25557 ( .A(n22375), .B(n22374), .Z(n22377) );
  NAND U25558 ( .A(n22377), .B(n22376), .Z(n22379) );
  ANDN U25559 ( .B(n22379), .A(n22378), .Z(n22381) );
  NANDN U25560 ( .A(n22381), .B(n22380), .Z(n22383) );
  ANDN U25561 ( .B(n22383), .A(n22382), .Z(n22384) );
  OR U25562 ( .A(n22385), .B(n22384), .Z(n22386) );
  NANDN U25563 ( .A(n22387), .B(n22386), .Z(n22389) );
  ANDN U25564 ( .B(n22389), .A(n22388), .Z(n22391) );
  NANDN U25565 ( .A(n22391), .B(n22390), .Z(n22393) );
  ANDN U25566 ( .B(n22393), .A(n22392), .Z(n22395) );
  NANDN U25567 ( .A(n22395), .B(n22394), .Z(n22397) );
  ANDN U25568 ( .B(n22397), .A(n22396), .Z(n22398) );
  OR U25569 ( .A(n22399), .B(n22398), .Z(n22401) );
  ANDN U25570 ( .B(n22401), .A(n22400), .Z(n22402) );
  OR U25571 ( .A(n22403), .B(n22402), .Z(n22405) );
  NAND U25572 ( .A(n22405), .B(n22404), .Z(n22406) );
  NANDN U25573 ( .A(n22407), .B(n22406), .Z(n22409) );
  ANDN U25574 ( .B(n22409), .A(n22408), .Z(n22411) );
  NANDN U25575 ( .A(n22411), .B(n22410), .Z(n22412) );
  NANDN U25576 ( .A(n22413), .B(n22412), .Z(n22415) );
  NAND U25577 ( .A(n22415), .B(n22414), .Z(n22416) );
  NANDN U25578 ( .A(n22417), .B(n22416), .Z(n22418) );
  NANDN U25579 ( .A(n22419), .B(n22418), .Z(n22420) );
  NANDN U25580 ( .A(n22421), .B(n22420), .Z(n22423) );
  ANDN U25581 ( .B(n22423), .A(n22422), .Z(n22425) );
  NANDN U25582 ( .A(n22425), .B(n22424), .Z(n22427) );
  NAND U25583 ( .A(n22427), .B(n22426), .Z(n22429) );
  NAND U25584 ( .A(n22429), .B(n22428), .Z(n22431) );
  NAND U25585 ( .A(n22431), .B(n22430), .Z(n22433) );
  NAND U25586 ( .A(n22433), .B(n22432), .Z(n22435) );
  ANDN U25587 ( .B(n22435), .A(n22434), .Z(n22437) );
  NANDN U25588 ( .A(n22437), .B(n22436), .Z(n22438) );
  AND U25589 ( .A(n22439), .B(n22438), .Z(n22441) );
  NANDN U25590 ( .A(n22441), .B(n22440), .Z(n22442) );
  AND U25591 ( .A(n22443), .B(n22442), .Z(n22445) );
  NANDN U25592 ( .A(n22445), .B(n22444), .Z(n22447) );
  NAND U25593 ( .A(n22447), .B(n22446), .Z(n22448) );
  NANDN U25594 ( .A(n22449), .B(n22448), .Z(n22451) );
  NAND U25595 ( .A(n22451), .B(n22450), .Z(n22453) );
  ANDN U25596 ( .B(n22453), .A(n22452), .Z(n22454) );
  OR U25597 ( .A(n22455), .B(n22454), .Z(n22457) );
  NAND U25598 ( .A(n22457), .B(n22456), .Z(n22458) );
  NANDN U25599 ( .A(n22459), .B(n22458), .Z(n22461) );
  ANDN U25600 ( .B(n22461), .A(n22460), .Z(n22463) );
  NANDN U25601 ( .A(n22463), .B(n22462), .Z(n22464) );
  AND U25602 ( .A(n22465), .B(n22464), .Z(n22467) );
  NANDN U25603 ( .A(n22467), .B(n22466), .Z(n22469) );
  NAND U25604 ( .A(n22469), .B(n22468), .Z(n22471) );
  NAND U25605 ( .A(n22471), .B(n22470), .Z(n22473) );
  NAND U25606 ( .A(n22473), .B(n22472), .Z(n22474) );
  AND U25607 ( .A(n22475), .B(n22474), .Z(n22477) );
  NANDN U25608 ( .A(n22477), .B(n22476), .Z(n22478) );
  NANDN U25609 ( .A(n22479), .B(n22478), .Z(n22481) );
  NAND U25610 ( .A(n22481), .B(n22480), .Z(n22483) );
  NAND U25611 ( .A(n22483), .B(n22482), .Z(n22485) );
  NAND U25612 ( .A(n22485), .B(n22484), .Z(n22487) );
  NAND U25613 ( .A(n22487), .B(n22486), .Z(n22488) );
  NANDN U25614 ( .A(n22489), .B(n22488), .Z(n22491) );
  NAND U25615 ( .A(n22491), .B(n22490), .Z(n22493) );
  ANDN U25616 ( .B(n22493), .A(n22492), .Z(n22495) );
  NOR U25617 ( .A(n22495), .B(n22494), .Z(n22497) );
  NANDN U25618 ( .A(n22497), .B(n22496), .Z(n22498) );
  NANDN U25619 ( .A(n22499), .B(n22498), .Z(n22501) );
  NAND U25620 ( .A(n22501), .B(n22500), .Z(n22503) );
  NAND U25621 ( .A(n22503), .B(n22502), .Z(n22505) );
  ANDN U25622 ( .B(n22505), .A(n22504), .Z(n22506) );
  NAND U25623 ( .A(n22507), .B(n22506), .Z(n22508) );
  NAND U25624 ( .A(n22509), .B(n22508), .Z(n22510) );
  NANDN U25625 ( .A(n22511), .B(n22510), .Z(n22513) );
  NAND U25626 ( .A(n22513), .B(n22512), .Z(n22515) );
  ANDN U25627 ( .B(n22515), .A(n22514), .Z(n22517) );
  NANDN U25628 ( .A(n22517), .B(n22516), .Z(n22519) );
  ANDN U25629 ( .B(n22519), .A(n22518), .Z(n22521) );
  NANDN U25630 ( .A(n22521), .B(n22520), .Z(n22523) );
  ANDN U25631 ( .B(n22523), .A(n22522), .Z(n22525) );
  NANDN U25632 ( .A(n22525), .B(n22524), .Z(n22527) );
  ANDN U25633 ( .B(n22527), .A(n22526), .Z(n22529) );
  NANDN U25634 ( .A(n22529), .B(n22528), .Z(n22531) );
  NAND U25635 ( .A(n22531), .B(n22530), .Z(n22532) );
  NANDN U25636 ( .A(n22533), .B(n22532), .Z(n22537) );
  NANDN U25637 ( .A(n22535), .B(n22534), .Z(n22536) );
  AND U25638 ( .A(n22537), .B(n22536), .Z(n22539) );
  NAND U25639 ( .A(n22539), .B(n22538), .Z(n22540) );
  NANDN U25640 ( .A(n22541), .B(n22540), .Z(n22542) );
  NANDN U25641 ( .A(n22543), .B(n22542), .Z(n22545) );
  NAND U25642 ( .A(n22545), .B(n22544), .Z(n22546) );
  NANDN U25643 ( .A(n22547), .B(n22546), .Z(n22549) );
  NAND U25644 ( .A(n22549), .B(n22548), .Z(n22550) );
  AND U25645 ( .A(n22551), .B(n22550), .Z(n22553) );
  NANDN U25646 ( .A(n22553), .B(n22552), .Z(n22555) );
  ANDN U25647 ( .B(n22555), .A(n22554), .Z(n22556) );
  OR U25648 ( .A(n22557), .B(n22556), .Z(n22558) );
  NANDN U25649 ( .A(n22559), .B(n22558), .Z(n22561) );
  NAND U25650 ( .A(n22561), .B(n22560), .Z(n22562) );
  NANDN U25651 ( .A(n22563), .B(n22562), .Z(n22565) );
  NAND U25652 ( .A(n22565), .B(n22564), .Z(n22567) );
  ANDN U25653 ( .B(n22567), .A(n22566), .Z(n22569) );
  NANDN U25654 ( .A(n22569), .B(n22568), .Z(n22571) );
  ANDN U25655 ( .B(n22571), .A(n22570), .Z(n22573) );
  NANDN U25656 ( .A(n22573), .B(n22572), .Z(n22574) );
  NANDN U25657 ( .A(n22575), .B(n22574), .Z(n22577) );
  NAND U25658 ( .A(n22577), .B(n22576), .Z(n22579) );
  NAND U25659 ( .A(n22579), .B(n22578), .Z(n22581) );
  NAND U25660 ( .A(n22581), .B(n22580), .Z(n22582) );
  AND U25661 ( .A(n22583), .B(n22582), .Z(n22585) );
  NANDN U25662 ( .A(n22585), .B(n22584), .Z(n22587) );
  NAND U25663 ( .A(n22587), .B(n22586), .Z(n22589) );
  NAND U25664 ( .A(n22589), .B(n22588), .Z(n22591) );
  NAND U25665 ( .A(n22591), .B(n22590), .Z(n22592) );
  NANDN U25666 ( .A(n22593), .B(n22592), .Z(n22595) );
  NAND U25667 ( .A(n22595), .B(n22594), .Z(n22596) );
  NANDN U25668 ( .A(n22597), .B(n22596), .Z(n22599) );
  NAND U25669 ( .A(n22599), .B(n22598), .Z(n22601) );
  ANDN U25670 ( .B(n22601), .A(n22600), .Z(n22602) );
  OR U25671 ( .A(n22603), .B(n22602), .Z(n22604) );
  NANDN U25672 ( .A(n22605), .B(n22604), .Z(n22606) );
  NANDN U25673 ( .A(n22607), .B(n22606), .Z(n22609) );
  ANDN U25674 ( .B(n22609), .A(n22608), .Z(n22611) );
  NANDN U25675 ( .A(n22611), .B(n22610), .Z(n22612) );
  NANDN U25676 ( .A(n22613), .B(n22612), .Z(n22615) );
  NAND U25677 ( .A(n22615), .B(n22614), .Z(n22617) );
  NAND U25678 ( .A(n22617), .B(n22616), .Z(n22618) );
  AND U25679 ( .A(n22619), .B(n22618), .Z(n22620) );
  OR U25680 ( .A(n22621), .B(n22620), .Z(n22622) );
  NANDN U25681 ( .A(n22623), .B(n22622), .Z(n22625) );
  ANDN U25682 ( .B(n22625), .A(n22624), .Z(n22626) );
  OR U25683 ( .A(n22627), .B(n22626), .Z(n22628) );
  NANDN U25684 ( .A(n22629), .B(n22628), .Z(n22630) );
  NANDN U25685 ( .A(n22631), .B(n22630), .Z(n22632) );
  NANDN U25686 ( .A(n22633), .B(n22632), .Z(n22635) );
  NAND U25687 ( .A(n22635), .B(n22634), .Z(n22637) );
  NAND U25688 ( .A(n22637), .B(n22636), .Z(n22639) );
  NAND U25689 ( .A(n22639), .B(n22638), .Z(n22640) );
  NANDN U25690 ( .A(n22641), .B(n22640), .Z(n22643) );
  ANDN U25691 ( .B(n22643), .A(n22642), .Z(n22645) );
  NANDN U25692 ( .A(n22645), .B(n22644), .Z(n22647) );
  NAND U25693 ( .A(n22647), .B(n22646), .Z(n22648) );
  NANDN U25694 ( .A(n22649), .B(n22648), .Z(n22651) );
  NAND U25695 ( .A(n22651), .B(n22650), .Z(n22653) );
  ANDN U25696 ( .B(n22653), .A(n22652), .Z(n22655) );
  NANDN U25697 ( .A(n22655), .B(n22654), .Z(n22656) );
  NANDN U25698 ( .A(n22657), .B(n22656), .Z(n22659) );
  NAND U25699 ( .A(n22659), .B(n22658), .Z(n22660) );
  NANDN U25700 ( .A(n22661), .B(n22660), .Z(n22663) );
  NAND U25701 ( .A(n22663), .B(n22662), .Z(n22664) );
  AND U25702 ( .A(n22665), .B(n22664), .Z(n22667) );
  NANDN U25703 ( .A(n22667), .B(n22666), .Z(n22668) );
  NANDN U25704 ( .A(n22669), .B(n22668), .Z(n22670) );
  NANDN U25705 ( .A(n22671), .B(n22670), .Z(n22672) );
  NANDN U25706 ( .A(n22673), .B(n22672), .Z(n22674) );
  NANDN U25707 ( .A(n22675), .B(n22674), .Z(n22676) );
  AND U25708 ( .A(n22677), .B(n22676), .Z(n22679) );
  NANDN U25709 ( .A(n22679), .B(n22678), .Z(n22681) );
  NAND U25710 ( .A(n22681), .B(n22680), .Z(n22683) );
  NAND U25711 ( .A(n22683), .B(n22682), .Z(n22684) );
  NANDN U25712 ( .A(n22685), .B(n22684), .Z(n22686) );
  NANDN U25713 ( .A(n22687), .B(n22686), .Z(n22689) );
  NAND U25714 ( .A(n22689), .B(n22688), .Z(n22691) );
  NAND U25715 ( .A(n22691), .B(n22690), .Z(n22692) );
  AND U25716 ( .A(n22693), .B(n22692), .Z(n22695) );
  NANDN U25717 ( .A(n22695), .B(n22694), .Z(n22697) );
  ANDN U25718 ( .B(n22697), .A(n22696), .Z(n22699) );
  OR U25719 ( .A(n22699), .B(n22698), .Z(n22701) );
  ANDN U25720 ( .B(n22701), .A(n22700), .Z(n22703) );
  OR U25721 ( .A(n22703), .B(n22702), .Z(n22704) );
  AND U25722 ( .A(n22705), .B(n22704), .Z(n22707) );
  NANDN U25723 ( .A(n22707), .B(n22706), .Z(n22709) );
  NAND U25724 ( .A(n22709), .B(n22708), .Z(n22711) );
  NAND U25725 ( .A(n22711), .B(n22710), .Z(n22713) );
  NAND U25726 ( .A(n22713), .B(n22712), .Z(n22714) );
  NANDN U25727 ( .A(n22715), .B(n22714), .Z(n22717) );
  NAND U25728 ( .A(n22717), .B(n22716), .Z(n22719) );
  NAND U25729 ( .A(n22719), .B(n22718), .Z(n22720) );
  NANDN U25730 ( .A(n22721), .B(n22720), .Z(n22723) );
  ANDN U25731 ( .B(n22723), .A(n22722), .Z(n22724) );
  OR U25732 ( .A(n22725), .B(n22724), .Z(n22726) );
  NANDN U25733 ( .A(n22727), .B(n22726), .Z(n22728) );
  NANDN U25734 ( .A(n22729), .B(n22728), .Z(n22731) );
  NAND U25735 ( .A(n22731), .B(n22730), .Z(n22732) );
  NANDN U25736 ( .A(n22733), .B(n22732), .Z(n22735) );
  NAND U25737 ( .A(n22735), .B(n22734), .Z(n22736) );
  NANDN U25738 ( .A(n22737), .B(n22736), .Z(n22739) );
  NAND U25739 ( .A(n22739), .B(n22738), .Z(n22740) );
  AND U25740 ( .A(n22741), .B(n22740), .Z(n22743) );
  OR U25741 ( .A(n22743), .B(n22742), .Z(n22745) );
  ANDN U25742 ( .B(n22745), .A(n22744), .Z(n22747) );
  NANDN U25743 ( .A(n22747), .B(n22746), .Z(n22749) );
  NAND U25744 ( .A(n22749), .B(n22748), .Z(n22751) );
  ANDN U25745 ( .B(n22751), .A(n22750), .Z(n22753) );
  NANDN U25746 ( .A(n22753), .B(n22752), .Z(n22754) );
  NANDN U25747 ( .A(n22755), .B(n22754), .Z(n22757) );
  NAND U25748 ( .A(n22757), .B(n22756), .Z(n22758) );
  NANDN U25749 ( .A(n22759), .B(n22758), .Z(n22761) );
  NAND U25750 ( .A(n22761), .B(n22760), .Z(n22762) );
  AND U25751 ( .A(n22763), .B(n22762), .Z(n22765) );
  NANDN U25752 ( .A(n22765), .B(n22764), .Z(n22767) );
  NAND U25753 ( .A(n22767), .B(n22766), .Z(n22769) );
  NAND U25754 ( .A(n22769), .B(n22768), .Z(n22773) );
  NAND U25755 ( .A(n22771), .B(n22770), .Z(n22772) );
  AND U25756 ( .A(n22773), .B(n22772), .Z(n22774) );
  NANDN U25757 ( .A(n22775), .B(n22774), .Z(n22776) );
  NANDN U25758 ( .A(n22777), .B(n22776), .Z(n22779) );
  NAND U25759 ( .A(n22779), .B(n22778), .Z(n22780) );
  AND U25760 ( .A(n22781), .B(n22780), .Z(n22783) );
  NANDN U25761 ( .A(n22783), .B(n22782), .Z(n22785) );
  ANDN U25762 ( .B(n22785), .A(n22784), .Z(n22787) );
  NANDN U25763 ( .A(n22787), .B(n22786), .Z(n22788) );
  NANDN U25764 ( .A(n22789), .B(n22788), .Z(n22791) );
  NAND U25765 ( .A(n22791), .B(n22790), .Z(n22792) );
  NANDN U25766 ( .A(n22793), .B(n22792), .Z(n22795) );
  AND U25767 ( .A(n22795), .B(n22794), .Z(n22796) );
  NANDN U25768 ( .A(n22796), .B(n22797), .Z(n22800) );
  XNOR U25769 ( .A(n22797), .B(n22796), .Z(n22798) );
  NAND U25770 ( .A(n22798), .B(y[1472]), .Z(n22799) );
  NAND U25771 ( .A(n22800), .B(n22799), .Z(n22801) );
  AND U25772 ( .A(n22802), .B(n22801), .Z(n22804) );
  NANDN U25773 ( .A(n22804), .B(n22803), .Z(n22805) );
  NANDN U25774 ( .A(n22806), .B(n22805), .Z(n22807) );
  AND U25775 ( .A(n22808), .B(n22807), .Z(n22809) );
  OR U25776 ( .A(n22810), .B(n22809), .Z(n22811) );
  NANDN U25777 ( .A(n22812), .B(n22811), .Z(n22814) );
  NAND U25778 ( .A(n22814), .B(n22813), .Z(n22815) );
  NANDN U25779 ( .A(n22816), .B(n22815), .Z(n22817) );
  NANDN U25780 ( .A(n22818), .B(n22817), .Z(n22820) );
  NAND U25781 ( .A(n22820), .B(n22819), .Z(n22822) );
  ANDN U25782 ( .B(n22822), .A(n22821), .Z(n22824) );
  NANDN U25783 ( .A(n22824), .B(n22823), .Z(n22826) );
  NAND U25784 ( .A(n22826), .B(n22825), .Z(n22828) );
  NAND U25785 ( .A(n22828), .B(n22827), .Z(n22830) );
  NAND U25786 ( .A(n22830), .B(n22829), .Z(n22832) );
  NAND U25787 ( .A(n22832), .B(n22831), .Z(n22834) );
  ANDN U25788 ( .B(n22834), .A(n22833), .Z(n22835) );
  OR U25789 ( .A(n22836), .B(n22835), .Z(n22837) );
  NANDN U25790 ( .A(n22838), .B(n22837), .Z(n22839) );
  NANDN U25791 ( .A(n22840), .B(n22839), .Z(n22841) );
  NANDN U25792 ( .A(n22842), .B(n22841), .Z(n22844) );
  NAND U25793 ( .A(n22844), .B(n22843), .Z(n22846) );
  ANDN U25794 ( .B(n22846), .A(n22845), .Z(n22848) );
  NANDN U25795 ( .A(n22848), .B(n22847), .Z(n22850) );
  ANDN U25796 ( .B(n22850), .A(n22849), .Z(n22851) );
  ANDN U25797 ( .B(n22852), .A(n22851), .Z(n22854) );
  NANDN U25798 ( .A(n22854), .B(n22853), .Z(n22856) );
  NAND U25799 ( .A(n22856), .B(n22855), .Z(n22858) );
  NAND U25800 ( .A(n22858), .B(n22857), .Z(n22859) );
  NANDN U25801 ( .A(n22860), .B(n22859), .Z(n22862) );
  NAND U25802 ( .A(n22862), .B(n22861), .Z(n22864) );
  ANDN U25803 ( .B(n22864), .A(n22863), .Z(n22865) );
  OR U25804 ( .A(n22866), .B(n22865), .Z(n22868) );
  NAND U25805 ( .A(n22868), .B(n22867), .Z(n22869) );
  AND U25806 ( .A(n22870), .B(n22869), .Z(n22872) );
  NANDN U25807 ( .A(n22872), .B(n22871), .Z(n22874) );
  NAND U25808 ( .A(n22874), .B(n22873), .Z(n22876) );
  NAND U25809 ( .A(n22876), .B(n22875), .Z(n22877) );
  NAND U25810 ( .A(n22878), .B(n22877), .Z(n22879) );
  NANDN U25811 ( .A(n22880), .B(n22879), .Z(n22881) );
  NANDN U25812 ( .A(n22882), .B(n22881), .Z(n22883) );
  NANDN U25813 ( .A(n22884), .B(n22883), .Z(n22885) );
  AND U25814 ( .A(n22886), .B(n22885), .Z(n22888) );
  NANDN U25815 ( .A(n22888), .B(n22887), .Z(n22889) );
  AND U25816 ( .A(n22890), .B(n22889), .Z(n22892) );
  NANDN U25817 ( .A(n22892), .B(n22891), .Z(n22893) );
  AND U25818 ( .A(n22894), .B(n22893), .Z(n22895) );
  OR U25819 ( .A(n22896), .B(n22895), .Z(n22897) );
  NANDN U25820 ( .A(n22898), .B(n22897), .Z(n22900) );
  NAND U25821 ( .A(n22900), .B(n22899), .Z(n22901) );
  NANDN U25822 ( .A(n22902), .B(n22901), .Z(n22903) );
  NANDN U25823 ( .A(n22904), .B(n22903), .Z(n22905) );
  AND U25824 ( .A(n22906), .B(n22905), .Z(n22908) );
  NANDN U25825 ( .A(n22908), .B(n22907), .Z(n22909) );
  AND U25826 ( .A(n22910), .B(n22909), .Z(n22912) );
  NANDN U25827 ( .A(n22912), .B(n22911), .Z(n22913) );
  AND U25828 ( .A(n22914), .B(n22913), .Z(n22916) );
  NANDN U25829 ( .A(n22916), .B(n22915), .Z(n22918) );
  NAND U25830 ( .A(n22918), .B(n22917), .Z(n22920) );
  NAND U25831 ( .A(n22920), .B(n22919), .Z(n22921) );
  NANDN U25832 ( .A(n22922), .B(n22921), .Z(n22924) );
  NAND U25833 ( .A(n22924), .B(n22923), .Z(n22925) );
  NANDN U25834 ( .A(n22926), .B(n22925), .Z(n22928) );
  NAND U25835 ( .A(n22928), .B(n22927), .Z(n22929) );
  AND U25836 ( .A(n22930), .B(n22929), .Z(n22931) );
  ANDN U25837 ( .B(n22932), .A(n22931), .Z(n22934) );
  NANDN U25838 ( .A(n22934), .B(n22933), .Z(n22935) );
  AND U25839 ( .A(n22936), .B(n22935), .Z(n22938) );
  NANDN U25840 ( .A(n22938), .B(n22937), .Z(n22940) );
  NAND U25841 ( .A(n22940), .B(n22939), .Z(n22942) );
  NAND U25842 ( .A(n22942), .B(n22941), .Z(n22943) );
  NANDN U25843 ( .A(n22944), .B(n22943), .Z(n22946) );
  ANDN U25844 ( .B(n22946), .A(n22945), .Z(n22948) );
  NOR U25845 ( .A(n22948), .B(n22947), .Z(n22949) );
  NAND U25846 ( .A(n22950), .B(n22949), .Z(n22951) );
  NAND U25847 ( .A(n22952), .B(n22951), .Z(n22953) );
  NANDN U25848 ( .A(n22954), .B(n22953), .Z(n22956) );
  NAND U25849 ( .A(n22956), .B(n22955), .Z(n22958) );
  ANDN U25850 ( .B(n22958), .A(n22957), .Z(n22960) );
  NANDN U25851 ( .A(n22960), .B(n22959), .Z(n22962) );
  ANDN U25852 ( .B(n22962), .A(n22961), .Z(n22964) );
  NANDN U25853 ( .A(n22964), .B(n22963), .Z(n22966) );
  NAND U25854 ( .A(n22966), .B(n22965), .Z(n22968) );
  NAND U25855 ( .A(n22968), .B(n22967), .Z(n22970) );
  NAND U25856 ( .A(n22970), .B(n22969), .Z(n22972) );
  ANDN U25857 ( .B(n22972), .A(n22971), .Z(n22973) );
  OR U25858 ( .A(n22974), .B(n22973), .Z(n22975) );
  NANDN U25859 ( .A(n22976), .B(n22975), .Z(n22978) );
  NAND U25860 ( .A(n22978), .B(n22977), .Z(n22979) );
  AND U25861 ( .A(n22980), .B(n22979), .Z(n22982) );
  NANDN U25862 ( .A(n22982), .B(n22981), .Z(n22983) );
  NANDN U25863 ( .A(n22984), .B(n22983), .Z(n22986) );
  NAND U25864 ( .A(n22986), .B(n22985), .Z(n22987) );
  NANDN U25865 ( .A(n22988), .B(n22987), .Z(n22990) );
  NAND U25866 ( .A(n22990), .B(n22989), .Z(n22992) );
  NAND U25867 ( .A(n22992), .B(n22991), .Z(n22994) );
  NAND U25868 ( .A(n22994), .B(n22993), .Z(n22996) );
  NAND U25869 ( .A(n22996), .B(n22995), .Z(n22998) );
  ANDN U25870 ( .B(n22998), .A(n22997), .Z(n23000) );
  NANDN U25871 ( .A(n23000), .B(n22999), .Z(n23002) );
  NAND U25872 ( .A(n23002), .B(n23001), .Z(n23004) );
  NAND U25873 ( .A(n23004), .B(n23003), .Z(n23005) );
  NANDN U25874 ( .A(n23006), .B(n23005), .Z(n23008) );
  NAND U25875 ( .A(n23008), .B(n23007), .Z(n23009) );
  AND U25876 ( .A(n23010), .B(n23009), .Z(n23012) );
  NANDN U25877 ( .A(n23012), .B(n23011), .Z(n23013) );
  AND U25878 ( .A(n23014), .B(n23013), .Z(n23016) );
  NANDN U25879 ( .A(n23016), .B(n23015), .Z(n23017) );
  AND U25880 ( .A(n23018), .B(n23017), .Z(n23020) );
  NANDN U25881 ( .A(n23020), .B(n23019), .Z(n23021) );
  AND U25882 ( .A(n23022), .B(n23021), .Z(n23024) );
  NANDN U25883 ( .A(n23024), .B(n23023), .Z(n23026) );
  ANDN U25884 ( .B(n23026), .A(n23025), .Z(n23027) );
  OR U25885 ( .A(n23028), .B(n23027), .Z(n23030) );
  NAND U25886 ( .A(n23030), .B(n23029), .Z(n23031) );
  NANDN U25887 ( .A(n23032), .B(n23031), .Z(n23033) );
  NANDN U25888 ( .A(n23034), .B(n23033), .Z(n23036) );
  NAND U25889 ( .A(n23036), .B(n23035), .Z(n23038) );
  ANDN U25890 ( .B(n23038), .A(n23037), .Z(n23040) );
  NANDN U25891 ( .A(n23040), .B(n23039), .Z(n23041) );
  NANDN U25892 ( .A(n23042), .B(n23041), .Z(n23044) );
  NAND U25893 ( .A(n23044), .B(n23043), .Z(n23045) );
  NANDN U25894 ( .A(n23046), .B(n23045), .Z(n23048) );
  NAND U25895 ( .A(n23048), .B(n23047), .Z(n23050) );
  NAND U25896 ( .A(n23050), .B(n23049), .Z(n23052) );
  NAND U25897 ( .A(n23052), .B(n23051), .Z(n23054) );
  NAND U25898 ( .A(n23054), .B(n23053), .Z(n23056) );
  ANDN U25899 ( .B(n23056), .A(n23055), .Z(n23058) );
  NANDN U25900 ( .A(n23058), .B(n23057), .Z(n23060) );
  ANDN U25901 ( .B(n23060), .A(n23059), .Z(n23062) );
  OR U25902 ( .A(n23062), .B(n23061), .Z(n23064) );
  ANDN U25903 ( .B(n23064), .A(n23063), .Z(n23066) );
  NANDN U25904 ( .A(n23066), .B(n23065), .Z(n23068) );
  NAND U25905 ( .A(n23068), .B(n23067), .Z(n23070) );
  NAND U25906 ( .A(n23070), .B(n23069), .Z(n23072) );
  NAND U25907 ( .A(n23072), .B(n23071), .Z(n23074) );
  NAND U25908 ( .A(n23074), .B(n23073), .Z(n23075) );
  AND U25909 ( .A(n23076), .B(n23075), .Z(n23078) );
  NANDN U25910 ( .A(n23078), .B(n23077), .Z(n23080) );
  NAND U25911 ( .A(n23080), .B(n23079), .Z(n23082) );
  NAND U25912 ( .A(n23082), .B(n23081), .Z(n23083) );
  NANDN U25913 ( .A(n23084), .B(n23083), .Z(n23086) );
  NAND U25914 ( .A(n23086), .B(n23085), .Z(n23088) );
  ANDN U25915 ( .B(n23088), .A(n23087), .Z(n23090) );
  NANDN U25916 ( .A(n23090), .B(n23089), .Z(n23092) );
  NAND U25917 ( .A(n23092), .B(n23091), .Z(n23094) );
  NAND U25918 ( .A(n23094), .B(n23093), .Z(n23095) );
  NANDN U25919 ( .A(n23096), .B(n23095), .Z(n23098) );
  ANDN U25920 ( .B(n23098), .A(n23097), .Z(n23100) );
  NANDN U25921 ( .A(n23100), .B(n23099), .Z(n23102) );
  NAND U25922 ( .A(n23102), .B(n23101), .Z(n23104) );
  NAND U25923 ( .A(n23104), .B(n23103), .Z(n23105) );
  NANDN U25924 ( .A(n23106), .B(n23105), .Z(n23108) );
  NAND U25925 ( .A(n23108), .B(n23107), .Z(n23110) );
  ANDN U25926 ( .B(n23110), .A(n23109), .Z(n23112) );
  NANDN U25927 ( .A(n23112), .B(n23111), .Z(n23113) );
  NANDN U25928 ( .A(n23114), .B(n23113), .Z(n23116) );
  NAND U25929 ( .A(n23116), .B(n23115), .Z(n23117) );
  NANDN U25930 ( .A(n23118), .B(n23117), .Z(n23120) );
  NAND U25931 ( .A(n23120), .B(n23119), .Z(n23121) );
  NANDN U25932 ( .A(n23122), .B(n23121), .Z(n23123) );
  NANDN U25933 ( .A(n23123), .B(x[1624]), .Z(n23127) );
  XNOR U25934 ( .A(n23123), .B(x[1624]), .Z(n23124) );
  NAND U25935 ( .A(n23125), .B(n23124), .Z(n23126) );
  NAND U25936 ( .A(n23127), .B(n23126), .Z(n23128) );
  NAND U25937 ( .A(n23129), .B(n23128), .Z(n23130) );
  NAND U25938 ( .A(n23131), .B(n23130), .Z(n23132) );
  AND U25939 ( .A(n23133), .B(n23132), .Z(n23134) );
  NANDN U25940 ( .A(n23135), .B(n23134), .Z(n23137) );
  NAND U25941 ( .A(n23137), .B(n23136), .Z(n23139) );
  NAND U25942 ( .A(n23139), .B(n23138), .Z(n23140) );
  NANDN U25943 ( .A(n23141), .B(n23140), .Z(n23142) );
  AND U25944 ( .A(n23143), .B(n23142), .Z(n23145) );
  NANDN U25945 ( .A(n23145), .B(n23144), .Z(n23147) );
  NAND U25946 ( .A(n23147), .B(n23146), .Z(n23149) );
  NAND U25947 ( .A(n23149), .B(n23148), .Z(n23150) );
  NANDN U25948 ( .A(n23151), .B(n23150), .Z(n23152) );
  AND U25949 ( .A(n23153), .B(n23152), .Z(n23155) );
  NAND U25950 ( .A(n23155), .B(n23154), .Z(n23156) );
  NAND U25951 ( .A(n23157), .B(n23156), .Z(n23159) );
  ANDN U25952 ( .B(n23159), .A(n23158), .Z(n23160) );
  NANDN U25953 ( .A(n23161), .B(n23160), .Z(n23163) );
  NAND U25954 ( .A(n23163), .B(n23162), .Z(n23165) );
  ANDN U25955 ( .B(n23165), .A(n23164), .Z(n23167) );
  NANDN U25956 ( .A(n23167), .B(n23166), .Z(n23168) );
  AND U25957 ( .A(n23169), .B(n23168), .Z(n23170) );
  OR U25958 ( .A(n23171), .B(n23170), .Z(n23172) );
  NANDN U25959 ( .A(n23173), .B(n23172), .Z(n23175) );
  NAND U25960 ( .A(n23175), .B(n23174), .Z(n23177) );
  NAND U25961 ( .A(n23177), .B(n23176), .Z(n23178) );
  AND U25962 ( .A(n23179), .B(n23178), .Z(n23181) );
  NANDN U25963 ( .A(n23181), .B(n23180), .Z(n23183) );
  NAND U25964 ( .A(n23183), .B(n23182), .Z(n23185) );
  NAND U25965 ( .A(n23185), .B(n23184), .Z(n23186) );
  NANDN U25966 ( .A(n23187), .B(n23186), .Z(n23189) );
  NAND U25967 ( .A(n23189), .B(n23188), .Z(n23191) );
  ANDN U25968 ( .B(n23191), .A(n23190), .Z(n23193) );
  NANDN U25969 ( .A(n23193), .B(n23192), .Z(n23195) );
  NAND U25970 ( .A(n23195), .B(n23194), .Z(n23197) );
  NAND U25971 ( .A(n23197), .B(n23196), .Z(n23198) );
  NANDN U25972 ( .A(n23199), .B(n23198), .Z(n23200) );
  NANDN U25973 ( .A(n23201), .B(n23200), .Z(n23203) );
  NAND U25974 ( .A(n23203), .B(n23202), .Z(n23204) );
  NAND U25975 ( .A(n23205), .B(n23204), .Z(n23206) );
  NAND U25976 ( .A(n23207), .B(n23206), .Z(n23209) );
  NANDN U25977 ( .A(n23209), .B(n23208), .Z(n23210) );
  AND U25978 ( .A(n23211), .B(n23210), .Z(n23212) );
  NANDN U25979 ( .A(n23213), .B(n23212), .Z(n23215) );
  NAND U25980 ( .A(n23215), .B(n23214), .Z(n23217) );
  ANDN U25981 ( .B(n23217), .A(n23216), .Z(n23218) );
  OR U25982 ( .A(n23219), .B(n23218), .Z(n23220) );
  NANDN U25983 ( .A(n23221), .B(n23220), .Z(n23223) );
  NAND U25984 ( .A(n23223), .B(n23222), .Z(n23225) );
  NAND U25985 ( .A(n23225), .B(n23224), .Z(n23226) );
  NANDN U25986 ( .A(n23227), .B(n23226), .Z(n23229) );
  ANDN U25987 ( .B(n23229), .A(n23228), .Z(n23231) );
  NANDN U25988 ( .A(n23231), .B(n23230), .Z(n23232) );
  AND U25989 ( .A(n23233), .B(n23232), .Z(n23235) );
  NANDN U25990 ( .A(n23235), .B(n23234), .Z(n23236) );
  NANDN U25991 ( .A(n23237), .B(n23236), .Z(n23239) );
  NAND U25992 ( .A(n23239), .B(n23238), .Z(n23241) );
  NAND U25993 ( .A(n23241), .B(n23240), .Z(n23243) );
  NAND U25994 ( .A(n23243), .B(n23242), .Z(n23244) );
  AND U25995 ( .A(n23245), .B(n23244), .Z(n23247) );
  NANDN U25996 ( .A(n23247), .B(n23246), .Z(n23249) );
  NAND U25997 ( .A(n23249), .B(n23248), .Z(n23251) );
  NAND U25998 ( .A(n23251), .B(n23250), .Z(n23253) );
  NAND U25999 ( .A(n23253), .B(n23252), .Z(n23255) );
  NAND U26000 ( .A(n23255), .B(n23254), .Z(n23257) );
  ANDN U26001 ( .B(n23257), .A(n23256), .Z(n23259) );
  NANDN U26002 ( .A(n23259), .B(n23258), .Z(n23260) );
  AND U26003 ( .A(n23261), .B(n23260), .Z(n23263) );
  NANDN U26004 ( .A(n23263), .B(n23262), .Z(n23264) );
  NANDN U26005 ( .A(n23265), .B(n23264), .Z(n23267) );
  ANDN U26006 ( .B(n23267), .A(n23266), .Z(n23268) );
  OR U26007 ( .A(n23269), .B(n23268), .Z(n23270) );
  NANDN U26008 ( .A(n23271), .B(n23270), .Z(n23273) );
  NAND U26009 ( .A(n23273), .B(n23272), .Z(n23275) );
  NAND U26010 ( .A(n23275), .B(n23274), .Z(n23277) );
  NAND U26011 ( .A(n23277), .B(n23276), .Z(n23279) );
  ANDN U26012 ( .B(n23279), .A(n23278), .Z(n23281) );
  NANDN U26013 ( .A(n23281), .B(n23280), .Z(n23282) );
  NAND U26014 ( .A(n23283), .B(n23282), .Z(n23285) );
  NAND U26015 ( .A(n23285), .B(n23284), .Z(n23286) );
  NANDN U26016 ( .A(n23287), .B(n23286), .Z(n23289) );
  NAND U26017 ( .A(n23289), .B(n23288), .Z(n23291) );
  ANDN U26018 ( .B(n23291), .A(n23290), .Z(n23293) );
  NANDN U26019 ( .A(n23293), .B(n23292), .Z(n23295) );
  NAND U26020 ( .A(n23295), .B(n23294), .Z(n23297) );
  NAND U26021 ( .A(n23297), .B(n23296), .Z(n23298) );
  AND U26022 ( .A(n23299), .B(n23298), .Z(n23301) );
  NANDN U26023 ( .A(n23301), .B(n23300), .Z(n23303) );
  ANDN U26024 ( .B(n23303), .A(n23302), .Z(n23305) );
  NANDN U26025 ( .A(n23305), .B(n23304), .Z(n23307) );
  NAND U26026 ( .A(n23307), .B(n23306), .Z(n23308) );
  NANDN U26027 ( .A(n23309), .B(n23308), .Z(n23311) );
  NAND U26028 ( .A(n23311), .B(n23310), .Z(n23312) );
  AND U26029 ( .A(n23313), .B(n23312), .Z(n23317) );
  ANDN U26030 ( .B(n23315), .A(n23314), .Z(n23316) );
  NANDN U26031 ( .A(n23317), .B(n23316), .Z(n23319) );
  NAND U26032 ( .A(n23319), .B(n23318), .Z(n23321) );
  NAND U26033 ( .A(n23321), .B(n23320), .Z(n23322) );
  NANDN U26034 ( .A(n23323), .B(n23322), .Z(n23325) );
  ANDN U26035 ( .B(n23325), .A(n23324), .Z(n23326) );
  OR U26036 ( .A(n23327), .B(n23326), .Z(n23328) );
  NANDN U26037 ( .A(n23329), .B(n23328), .Z(n23331) );
  NAND U26038 ( .A(n23331), .B(n23330), .Z(n23332) );
  NANDN U26039 ( .A(n23333), .B(n23332), .Z(n23335) );
  NAND U26040 ( .A(n23335), .B(n23334), .Z(n23336) );
  AND U26041 ( .A(n23337), .B(n23336), .Z(n23339) );
  OR U26042 ( .A(n23339), .B(n23338), .Z(n23341) );
  ANDN U26043 ( .B(n23341), .A(n23340), .Z(n23343) );
  NANDN U26044 ( .A(n23343), .B(n23342), .Z(n23345) );
  NAND U26045 ( .A(n23345), .B(n23344), .Z(n23347) );
  NAND U26046 ( .A(n23347), .B(n23346), .Z(n23348) );
  NANDN U26047 ( .A(n23349), .B(n23348), .Z(n23351) );
  NAND U26048 ( .A(n23351), .B(n23350), .Z(n23353) );
  ANDN U26049 ( .B(n23353), .A(n23352), .Z(n23355) );
  NANDN U26050 ( .A(n23355), .B(n23354), .Z(n23357) );
  ANDN U26051 ( .B(n23357), .A(n23356), .Z(n23359) );
  NANDN U26052 ( .A(n23359), .B(n23358), .Z(n23361) );
  NAND U26053 ( .A(n23361), .B(n23360), .Z(n23362) );
  AND U26054 ( .A(n23363), .B(n23362), .Z(n23365) );
  NANDN U26055 ( .A(n23365), .B(n23364), .Z(n23367) );
  NAND U26056 ( .A(n23367), .B(n23366), .Z(n23369) );
  NAND U26057 ( .A(n23369), .B(n23368), .Z(n23371) );
  NAND U26058 ( .A(n23371), .B(n23370), .Z(n23373) );
  NAND U26059 ( .A(n23373), .B(n23372), .Z(n23374) );
  AND U26060 ( .A(n23375), .B(n23374), .Z(n23377) );
  NANDN U26061 ( .A(n23377), .B(n23376), .Z(n23378) );
  AND U26062 ( .A(n23379), .B(n23378), .Z(n23381) );
  NANDN U26063 ( .A(n23381), .B(n23380), .Z(n23383) );
  NAND U26064 ( .A(n23383), .B(n23382), .Z(n23385) );
  ANDN U26065 ( .B(n23385), .A(n23384), .Z(n23387) );
  NANDN U26066 ( .A(n23387), .B(n23386), .Z(n23389) );
  ANDN U26067 ( .B(n23389), .A(n23388), .Z(n23391) );
  NANDN U26068 ( .A(n23391), .B(n23390), .Z(n23393) );
  NAND U26069 ( .A(n23393), .B(n23392), .Z(n23394) );
  AND U26070 ( .A(n23395), .B(n23394), .Z(n23397) );
  NANDN U26071 ( .A(n23397), .B(n23396), .Z(n23399) );
  NAND U26072 ( .A(n23399), .B(n23398), .Z(n23401) );
  NAND U26073 ( .A(n23401), .B(n23400), .Z(n23403) );
  NAND U26074 ( .A(n23403), .B(n23402), .Z(n23404) );
  NANDN U26075 ( .A(n23405), .B(n23404), .Z(n23407) );
  NAND U26076 ( .A(n23407), .B(n23406), .Z(n23408) );
  NANDN U26077 ( .A(n23409), .B(n23408), .Z(n23411) );
  NAND U26078 ( .A(n23411), .B(n23410), .Z(n23412) );
  AND U26079 ( .A(n23413), .B(n23412), .Z(n23414) );
  OR U26080 ( .A(n23415), .B(n23414), .Z(n23416) );
  NANDN U26081 ( .A(n23417), .B(n23416), .Z(n23419) );
  NAND U26082 ( .A(n23419), .B(n23418), .Z(n23420) );
  NANDN U26083 ( .A(n23421), .B(n23420), .Z(n23423) );
  NAND U26084 ( .A(n23423), .B(n23422), .Z(n23424) );
  AND U26085 ( .A(n23425), .B(n23424), .Z(n23427) );
  NANDN U26086 ( .A(n23427), .B(n23426), .Z(n23428) );
  NANDN U26087 ( .A(n23429), .B(n23428), .Z(n23431) );
  NAND U26088 ( .A(n23431), .B(n23430), .Z(n23433) );
  NAND U26089 ( .A(n23433), .B(n23432), .Z(n23435) );
  NAND U26090 ( .A(n23435), .B(n23434), .Z(n23437) );
  ANDN U26091 ( .B(n23437), .A(n23436), .Z(n23439) );
  NANDN U26092 ( .A(n23439), .B(n23438), .Z(n23441) );
  ANDN U26093 ( .B(n23441), .A(n23440), .Z(n23443) );
  NANDN U26094 ( .A(n23443), .B(n23442), .Z(n23444) );
  NANDN U26095 ( .A(n23445), .B(n23444), .Z(n23447) );
  NAND U26096 ( .A(n23447), .B(n23446), .Z(n23448) );
  NANDN U26097 ( .A(n23449), .B(n23448), .Z(n23451) );
  NAND U26098 ( .A(n23451), .B(n23450), .Z(n23452) );
  AND U26099 ( .A(n23453), .B(n23452), .Z(n23455) );
  NANDN U26100 ( .A(n23455), .B(n23454), .Z(n23457) );
  NAND U26101 ( .A(n23457), .B(n23456), .Z(n23458) );
  NANDN U26102 ( .A(n23459), .B(n23458), .Z(n23460) );
  NANDN U26103 ( .A(n23461), .B(n23460), .Z(n23462) );
  NANDN U26104 ( .A(n23463), .B(n23462), .Z(n23465) );
  ANDN U26105 ( .B(n23465), .A(n23464), .Z(n23467) );
  NANDN U26106 ( .A(n23467), .B(n23466), .Z(n23469) );
  NAND U26107 ( .A(n23469), .B(n23468), .Z(n23471) );
  NAND U26108 ( .A(n23471), .B(n23470), .Z(n23475) );
  NANDN U26109 ( .A(n23473), .B(n23472), .Z(n23474) );
  AND U26110 ( .A(n23475), .B(n23474), .Z(n23477) );
  NAND U26111 ( .A(n23477), .B(n23476), .Z(n23478) );
  NANDN U26112 ( .A(n23479), .B(n23478), .Z(n23481) );
  NAND U26113 ( .A(n23481), .B(n23480), .Z(n23483) );
  NAND U26114 ( .A(n23483), .B(n23482), .Z(n23484) );
  NANDN U26115 ( .A(n23485), .B(n23484), .Z(n23487) );
  NAND U26116 ( .A(n23487), .B(n23486), .Z(n23488) );
  AND U26117 ( .A(n23489), .B(n23488), .Z(n23490) );
  OR U26118 ( .A(n23491), .B(n23490), .Z(n23492) );
  NANDN U26119 ( .A(n23493), .B(n23492), .Z(n23494) );
  NANDN U26120 ( .A(n23495), .B(n23494), .Z(n23497) );
  NAND U26121 ( .A(n23497), .B(n23496), .Z(n23498) );
  NANDN U26122 ( .A(n23499), .B(n23498), .Z(n23501) );
  ANDN U26123 ( .B(n23501), .A(n23500), .Z(n23503) );
  NANDN U26124 ( .A(n23503), .B(n23502), .Z(n23505) );
  NAND U26125 ( .A(n23505), .B(n23504), .Z(n23507) );
  NAND U26126 ( .A(n23507), .B(n23506), .Z(n23508) );
  NANDN U26127 ( .A(n23509), .B(n23508), .Z(n23510) );
  AND U26128 ( .A(n23511), .B(n23510), .Z(n23513) );
  NAND U26129 ( .A(n23513), .B(n23512), .Z(n23514) );
  NANDN U26130 ( .A(n23515), .B(n23514), .Z(n23517) );
  NAND U26131 ( .A(n23517), .B(n23516), .Z(n23518) );
  AND U26132 ( .A(n23519), .B(n23518), .Z(n23521) );
  NANDN U26133 ( .A(n23521), .B(n23520), .Z(n23523) );
  NAND U26134 ( .A(n23523), .B(n23522), .Z(n23525) );
  NAND U26135 ( .A(n23525), .B(n23524), .Z(n23526) );
  NANDN U26136 ( .A(n23527), .B(n23526), .Z(n23529) );
  NAND U26137 ( .A(n23529), .B(n23528), .Z(n23531) );
  ANDN U26138 ( .B(n23531), .A(n23530), .Z(n23533) );
  NANDN U26139 ( .A(n23533), .B(n23532), .Z(n23534) );
  NANDN U26140 ( .A(n23535), .B(n23534), .Z(n23537) );
  NAND U26141 ( .A(n23537), .B(n23536), .Z(n23539) );
  NAND U26142 ( .A(n23539), .B(n23538), .Z(n23541) );
  NAND U26143 ( .A(n23541), .B(n23540), .Z(n23543) );
  ANDN U26144 ( .B(n23543), .A(n23542), .Z(n23545) );
  NANDN U26145 ( .A(n23545), .B(n23544), .Z(n23547) );
  NAND U26146 ( .A(n23547), .B(n23546), .Z(n23549) );
  NAND U26147 ( .A(n23549), .B(n23548), .Z(n23550) );
  NANDN U26148 ( .A(n23551), .B(n23550), .Z(n23552) );
  NANDN U26149 ( .A(n23553), .B(n23552), .Z(n23555) );
  NAND U26150 ( .A(n23555), .B(n23554), .Z(n23557) );
  ANDN U26151 ( .B(n23557), .A(n23556), .Z(n23558) );
  NANDN U26152 ( .A(n23559), .B(n23558), .Z(n23563) );
  ANDN U26153 ( .B(n23561), .A(n23560), .Z(n23562) );
  NAND U26154 ( .A(n23563), .B(n23562), .Z(n23564) );
  NANDN U26155 ( .A(n23565), .B(n23564), .Z(n23567) );
  NAND U26156 ( .A(n23567), .B(n23566), .Z(n23568) );
  AND U26157 ( .A(n23569), .B(n23568), .Z(n23571) );
  NANDN U26158 ( .A(n23571), .B(n23570), .Z(n23572) );
  AND U26159 ( .A(n23573), .B(n23572), .Z(n23575) );
  NANDN U26160 ( .A(n23575), .B(n23574), .Z(n23576) );
  NANDN U26161 ( .A(n23577), .B(n23576), .Z(n23578) );
  NANDN U26162 ( .A(n23579), .B(n23578), .Z(n23580) );
  NANDN U26163 ( .A(n23581), .B(n23580), .Z(n23583) );
  NAND U26164 ( .A(n23583), .B(n23582), .Z(n23585) );
  ANDN U26165 ( .B(n23585), .A(n23584), .Z(n23586) );
  NANDN U26166 ( .A(n23587), .B(n23586), .Z(n23588) );
  AND U26167 ( .A(n23589), .B(n23588), .Z(n23591) );
  NAND U26168 ( .A(n23591), .B(n23590), .Z(n23592) );
  NANDN U26169 ( .A(n23593), .B(n23592), .Z(n23595) );
  NANDN U26170 ( .A(n23595), .B(n23594), .Z(n23596) );
  NANDN U26171 ( .A(n23597), .B(n23596), .Z(n23599) );
  ANDN U26172 ( .B(n23599), .A(n23598), .Z(n23601) );
  NANDN U26173 ( .A(n23601), .B(n23600), .Z(n23602) );
  NANDN U26174 ( .A(n23603), .B(n23602), .Z(n23605) );
  NAND U26175 ( .A(n23605), .B(n23604), .Z(n23606) );
  NANDN U26176 ( .A(n23607), .B(n23606), .Z(n23608) );
  NANDN U26177 ( .A(n23608), .B(y[1833]), .Z(n23612) );
  XNOR U26178 ( .A(n23608), .B(y[1833]), .Z(n23609) );
  NAND U26179 ( .A(n23610), .B(n23609), .Z(n23611) );
  NAND U26180 ( .A(n23612), .B(n23611), .Z(n23613) );
  NAND U26181 ( .A(n23614), .B(n23613), .Z(n23615) );
  NAND U26182 ( .A(n23616), .B(n23615), .Z(n23618) );
  ANDN U26183 ( .B(n23618), .A(n23617), .Z(n23620) );
  NANDN U26184 ( .A(n23620), .B(n23619), .Z(n23621) );
  NANDN U26185 ( .A(n23622), .B(n23621), .Z(n23624) );
  NAND U26186 ( .A(n23624), .B(n23623), .Z(n23626) );
  NAND U26187 ( .A(n23626), .B(n23625), .Z(n23628) );
  NAND U26188 ( .A(n23628), .B(n23627), .Z(n23629) );
  AND U26189 ( .A(n23630), .B(n23629), .Z(n23631) );
  NANDN U26190 ( .A(n23632), .B(n23631), .Z(n23634) );
  NAND U26191 ( .A(n23634), .B(n23633), .Z(n23636) );
  ANDN U26192 ( .B(n23636), .A(n23635), .Z(n23638) );
  NAND U26193 ( .A(n23638), .B(n23637), .Z(n23640) );
  NAND U26194 ( .A(n23640), .B(n23639), .Z(n23642) );
  NAND U26195 ( .A(n23642), .B(n23641), .Z(n23643) );
  NANDN U26196 ( .A(n23644), .B(n23643), .Z(n23646) );
  NAND U26197 ( .A(n23646), .B(n23645), .Z(n23648) );
  NAND U26198 ( .A(n23648), .B(n23647), .Z(n23649) );
  NANDN U26199 ( .A(n23650), .B(n23649), .Z(n23652) );
  NAND U26200 ( .A(n23652), .B(n23651), .Z(n23654) );
  ANDN U26201 ( .B(n23654), .A(n23653), .Z(n23656) );
  NANDN U26202 ( .A(n23656), .B(n23655), .Z(n23657) );
  AND U26203 ( .A(n23658), .B(n23657), .Z(n23659) );
  OR U26204 ( .A(n23660), .B(n23659), .Z(n23661) );
  NANDN U26205 ( .A(n23662), .B(n23661), .Z(n23664) );
  NAND U26206 ( .A(n23664), .B(n23663), .Z(n23665) );
  NANDN U26207 ( .A(n23666), .B(n23665), .Z(n23668) );
  NAND U26208 ( .A(n23668), .B(n23667), .Z(n23669) );
  AND U26209 ( .A(n23670), .B(n23669), .Z(n23672) );
  NANDN U26210 ( .A(n23672), .B(n23671), .Z(n23673) );
  NANDN U26211 ( .A(n23674), .B(n23673), .Z(n23675) );
  NANDN U26212 ( .A(n23676), .B(n23675), .Z(n23677) );
  NANDN U26213 ( .A(n23678), .B(n23677), .Z(n23680) );
  NAND U26214 ( .A(n23680), .B(n23679), .Z(n23682) );
  ANDN U26215 ( .B(n23682), .A(n23681), .Z(n23684) );
  NANDN U26216 ( .A(n23684), .B(n23683), .Z(n23686) );
  ANDN U26217 ( .B(n23686), .A(n23685), .Z(n23687) );
  OR U26218 ( .A(n23688), .B(n23687), .Z(n23689) );
  AND U26219 ( .A(n23690), .B(n23689), .Z(n23691) );
  NANDN U26220 ( .A(n23692), .B(n23691), .Z(n23693) );
  NANDN U26221 ( .A(n23694), .B(n23693), .Z(n23696) );
  ANDN U26222 ( .B(n23696), .A(n23695), .Z(n23698) );
  NAND U26223 ( .A(n23698), .B(n23697), .Z(n23700) );
  NAND U26224 ( .A(n23700), .B(n23699), .Z(n23702) );
  NAND U26225 ( .A(n23702), .B(n23701), .Z(n23704) );
  NAND U26226 ( .A(n23704), .B(n23703), .Z(n23706) );
  ANDN U26227 ( .B(n23706), .A(n23705), .Z(n23707) );
  NAND U26228 ( .A(n23708), .B(n23707), .Z(n23710) );
  NAND U26229 ( .A(n23710), .B(n23709), .Z(n23711) );
  NANDN U26230 ( .A(n23712), .B(n23711), .Z(n23713) );
  NANDN U26231 ( .A(n23714), .B(n23713), .Z(n23716) );
  ANDN U26232 ( .B(n23716), .A(n23715), .Z(n23718) );
  NANDN U26233 ( .A(n23718), .B(n23717), .Z(n23720) );
  NAND U26234 ( .A(n23720), .B(n23719), .Z(n23721) );
  NANDN U26235 ( .A(n23722), .B(n23721), .Z(n23723) );
  NANDN U26236 ( .A(n23724), .B(n23723), .Z(n23726) );
  NAND U26237 ( .A(n23726), .B(n23725), .Z(n23727) );
  NANDN U26238 ( .A(n23728), .B(n23727), .Z(n23730) );
  NAND U26239 ( .A(n23730), .B(n23729), .Z(n23732) );
  NAND U26240 ( .A(n23732), .B(n23731), .Z(n23733) );
  AND U26241 ( .A(n23734), .B(n23733), .Z(n23736) );
  NANDN U26242 ( .A(n23736), .B(n23735), .Z(n23738) );
  NAND U26243 ( .A(n23738), .B(n23737), .Z(n23740) );
  NAND U26244 ( .A(n23740), .B(n23739), .Z(n23741) );
  NANDN U26245 ( .A(n23742), .B(n23741), .Z(n23744) );
  NAND U26246 ( .A(n23744), .B(n23743), .Z(n23745) );
  AND U26247 ( .A(n23746), .B(n23745), .Z(n23748) );
  NANDN U26248 ( .A(n23748), .B(n23747), .Z(n23749) );
  NANDN U26249 ( .A(n23750), .B(n23749), .Z(n23752) );
  NAND U26250 ( .A(n23752), .B(n23751), .Z(n23753) );
  AND U26251 ( .A(n23754), .B(n23753), .Z(n23756) );
  OR U26252 ( .A(n23756), .B(n23755), .Z(n23758) );
  ANDN U26253 ( .B(n23758), .A(n23757), .Z(n23760) );
  NANDN U26254 ( .A(n23760), .B(n23759), .Z(n23762) );
  NAND U26255 ( .A(n23762), .B(n23761), .Z(n23764) );
  NAND U26256 ( .A(n23764), .B(n23763), .Z(n23765) );
  NANDN U26257 ( .A(n23766), .B(n23765), .Z(n23767) );
  NANDN U26258 ( .A(n23768), .B(n23767), .Z(n23770) );
  ANDN U26259 ( .B(n23770), .A(n23769), .Z(n23772) );
  OR U26260 ( .A(n23772), .B(n23771), .Z(n23773) );
  AND U26261 ( .A(n23774), .B(n23773), .Z(n23776) );
  NANDN U26262 ( .A(n23776), .B(n23775), .Z(n23778) );
  NAND U26263 ( .A(n23778), .B(n23777), .Z(n23780) );
  NAND U26264 ( .A(n23780), .B(n23779), .Z(n23781) );
  AND U26265 ( .A(n23782), .B(n23781), .Z(n23783) );
  OR U26266 ( .A(n23783), .B(x[1907]), .Z(n23786) );
  XOR U26267 ( .A(x[1907]), .B(n23783), .Z(n23784) );
  NAND U26268 ( .A(y[1907]), .B(n23784), .Z(n23785) );
  NAND U26269 ( .A(n23786), .B(n23785), .Z(n23788) );
  ANDN U26270 ( .B(n23788), .A(n23787), .Z(n23790) );
  NANDN U26271 ( .A(n23790), .B(n23789), .Z(n23791) );
  NANDN U26272 ( .A(n23792), .B(n23791), .Z(n23794) );
  NAND U26273 ( .A(n23794), .B(n23793), .Z(n23795) );
  NANDN U26274 ( .A(n23796), .B(n23795), .Z(n23798) );
  NAND U26275 ( .A(n23798), .B(n23797), .Z(n23799) );
  AND U26276 ( .A(n23800), .B(n23799), .Z(n23802) );
  NANDN U26277 ( .A(n23802), .B(n23801), .Z(n23803) );
  NANDN U26278 ( .A(n23804), .B(n23803), .Z(n23806) );
  NAND U26279 ( .A(n23806), .B(n23805), .Z(n23807) );
  NANDN U26280 ( .A(n23808), .B(n23807), .Z(n23810) );
  ANDN U26281 ( .B(n23810), .A(n23809), .Z(n23812) );
  NAND U26282 ( .A(n23812), .B(n23811), .Z(n23813) );
  NANDN U26283 ( .A(n23814), .B(n23813), .Z(n23816) );
  NAND U26284 ( .A(n23816), .B(n23815), .Z(n23817) );
  AND U26285 ( .A(n23818), .B(n23817), .Z(n23819) );
  OR U26286 ( .A(n23820), .B(n23819), .Z(n23821) );
  NANDN U26287 ( .A(n23822), .B(n23821), .Z(n23824) );
  NAND U26288 ( .A(n23824), .B(n23823), .Z(n23825) );
  NAND U26289 ( .A(n23826), .B(n23825), .Z(n23827) );
  NAND U26290 ( .A(n23828), .B(n23827), .Z(n23830) );
  NANDN U26291 ( .A(n23830), .B(n23829), .Z(n23831) );
  AND U26292 ( .A(n23832), .B(n23831), .Z(n23834) );
  NAND U26293 ( .A(n23834), .B(n23833), .Z(n23836) );
  NAND U26294 ( .A(n23836), .B(n23835), .Z(n23837) );
  AND U26295 ( .A(n23838), .B(n23837), .Z(n23840) );
  NANDN U26296 ( .A(n23840), .B(n23839), .Z(n23842) );
  ANDN U26297 ( .B(n23842), .A(n23841), .Z(n23844) );
  NANDN U26298 ( .A(n23844), .B(n23843), .Z(n23845) );
  NANDN U26299 ( .A(n23846), .B(n23845), .Z(n23848) );
  NAND U26300 ( .A(n23848), .B(n23847), .Z(n23849) );
  AND U26301 ( .A(n23850), .B(n23849), .Z(n23851) );
  OR U26302 ( .A(n23852), .B(n23851), .Z(n23853) );
  AND U26303 ( .A(n23854), .B(n23853), .Z(n23856) );
  NANDN U26304 ( .A(n23856), .B(n23855), .Z(n23858) );
  NAND U26305 ( .A(n23858), .B(n23857), .Z(n23860) );
  NAND U26306 ( .A(n23860), .B(n23859), .Z(n23862) );
  NAND U26307 ( .A(n23862), .B(n23861), .Z(n23864) );
  NAND U26308 ( .A(n23864), .B(n23863), .Z(n23865) );
  AND U26309 ( .A(n23866), .B(n23865), .Z(n23868) );
  NANDN U26310 ( .A(n23868), .B(n23867), .Z(n23869) );
  AND U26311 ( .A(n23870), .B(n23869), .Z(n23872) );
  NANDN U26312 ( .A(n23872), .B(n23871), .Z(n23873) );
  AND U26313 ( .A(n23874), .B(n23873), .Z(n23876) );
  NANDN U26314 ( .A(n23876), .B(n23875), .Z(n23877) );
  NANDN U26315 ( .A(n23878), .B(n23877), .Z(n23880) );
  NAND U26316 ( .A(n23880), .B(n23879), .Z(n23882) );
  NAND U26317 ( .A(n23882), .B(n23881), .Z(n23884) );
  NAND U26318 ( .A(n23884), .B(n23883), .Z(n23888) );
  NANDN U26319 ( .A(n23886), .B(n23885), .Z(n23887) );
  NANDN U26320 ( .A(n23888), .B(n23887), .Z(n23889) );
  AND U26321 ( .A(n23890), .B(n23889), .Z(n23892) );
  NANDN U26322 ( .A(n23892), .B(n23891), .Z(n23893) );
  NANDN U26323 ( .A(n23894), .B(n23893), .Z(n23896) );
  NAND U26324 ( .A(n23896), .B(n23895), .Z(n23898) );
  NAND U26325 ( .A(n23898), .B(n23897), .Z(n23900) );
  NAND U26326 ( .A(n23900), .B(n23899), .Z(n23902) );
  NAND U26327 ( .A(n23902), .B(n23901), .Z(n23903) );
  OR U26328 ( .A(n23904), .B(n23903), .Z(n23905) );
  NANDN U26329 ( .A(n23906), .B(n23905), .Z(n23907) );
  NANDN U26330 ( .A(n23908), .B(n23907), .Z(n23909) );
  ANDN U26331 ( .B(n23910), .A(n23909), .Z(n23912) );
  NAND U26332 ( .A(n23912), .B(n23911), .Z(n23914) );
  ANDN U26333 ( .B(n23914), .A(n23913), .Z(n23916) );
  NANDN U26334 ( .A(n23916), .B(n23915), .Z(n23917) );
  NANDN U26335 ( .A(n23918), .B(n23917), .Z(n23920) );
  NAND U26336 ( .A(n23920), .B(n23919), .Z(n23921) );
  NANDN U26337 ( .A(n23922), .B(n23921), .Z(n23924) );
  NAND U26338 ( .A(n23924), .B(n23923), .Z(n23926) );
  ANDN U26339 ( .B(n23926), .A(n23925), .Z(n23928) );
  NANDN U26340 ( .A(n23928), .B(n23927), .Z(n23930) );
  NAND U26341 ( .A(n23930), .B(n23929), .Z(n23932) );
  ANDN U26342 ( .B(n23932), .A(n23931), .Z(n23933) );
  OR U26343 ( .A(n23934), .B(n23933), .Z(n23935) );
  NANDN U26344 ( .A(n23936), .B(n23935), .Z(n23938) );
  NAND U26345 ( .A(n23938), .B(n23937), .Z(n23939) );
  NANDN U26346 ( .A(n23940), .B(n23939), .Z(n23941) );
  NAND U26347 ( .A(n23942), .B(n23941), .Z(n23943) );
  NAND U26348 ( .A(n23944), .B(n23943), .Z(n23946) );
  NANDN U26349 ( .A(n23946), .B(n23945), .Z(n23947) );
  AND U26350 ( .A(n23948), .B(n23947), .Z(n23949) );
  OR U26351 ( .A(n23950), .B(n23949), .Z(n23952) );
  NAND U26352 ( .A(n23952), .B(n23951), .Z(n23953) );
  AND U26353 ( .A(n23954), .B(n23953), .Z(n23956) );
  NANDN U26354 ( .A(n23956), .B(n23955), .Z(n23957) );
  NANDN U26355 ( .A(n23958), .B(n23957), .Z(n23960) );
  NAND U26356 ( .A(n23960), .B(n23959), .Z(n23961) );
  NANDN U26357 ( .A(n23962), .B(n23961), .Z(n23963) );
  NANDN U26358 ( .A(n23964), .B(n23963), .Z(n23965) );
  AND U26359 ( .A(n23966), .B(n23965), .Z(n23968) );
  NANDN U26360 ( .A(n23968), .B(n23967), .Z(n23970) );
  ANDN U26361 ( .B(n23970), .A(n23969), .Z(n23972) );
  NANDN U26362 ( .A(n23972), .B(n23971), .Z(n23974) );
  NAND U26363 ( .A(n23974), .B(n23973), .Z(n23975) );
  AND U26364 ( .A(n23976), .B(n23975), .Z(n23977) );
  OR U26365 ( .A(n23978), .B(n23977), .Z(n23979) );
  AND U26366 ( .A(n23980), .B(n23979), .Z(n23984) );
  ANDN U26367 ( .B(n23982), .A(n23981), .Z(n23983) );
  NANDN U26368 ( .A(n23984), .B(n23983), .Z(n23986) );
  NAND U26369 ( .A(n23986), .B(n23985), .Z(n23988) );
  NAND U26370 ( .A(n23988), .B(n23987), .Z(n23989) );
  NANDN U26371 ( .A(n23990), .B(n23989), .Z(n23991) );
  AND U26372 ( .A(n23992), .B(n23991), .Z(n23994) );
  NANDN U26373 ( .A(n23994), .B(n23993), .Z(n23995) );
  NANDN U26374 ( .A(n23996), .B(n23995), .Z(n23997) );
  NANDN U26375 ( .A(n23998), .B(n23997), .Z(n24000) );
  NAND U26376 ( .A(n24000), .B(n23999), .Z(n24002) );
  NAND U26377 ( .A(n24002), .B(n24001), .Z(n24003) );
  AND U26378 ( .A(n24004), .B(n24003), .Z(n24006) );
  NANDN U26379 ( .A(n24006), .B(n24005), .Z(n24007) );
  NANDN U26380 ( .A(n24008), .B(n24007), .Z(n24009) );
  NANDN U26381 ( .A(n24010), .B(n24009), .Z(n24011) );
  NANDN U26382 ( .A(n24012), .B(n24011), .Z(n24014) );
  NAND U26383 ( .A(n24014), .B(n24013), .Z(n24016) );
  ANDN U26384 ( .B(n24016), .A(n24015), .Z(n24017) );
  OR U26385 ( .A(n24018), .B(n24017), .Z(n24019) );
  AND U26386 ( .A(n24020), .B(n24019), .Z(n24022) );
  NANDN U26387 ( .A(n24022), .B(n24021), .Z(n24024) );
  NAND U26388 ( .A(n24024), .B(n24023), .Z(n24026) );
  NAND U26389 ( .A(n24026), .B(n24025), .Z(n24028) );
  NAND U26390 ( .A(n24028), .B(n24027), .Z(n24030) );
  NAND U26391 ( .A(n24030), .B(n24029), .Z(n24032) );
  ANDN U26392 ( .B(n24032), .A(n24031), .Z(n24033) );
  NAND U26393 ( .A(n24034), .B(n24033), .Z(n24035) );
  NAND U26394 ( .A(n24036), .B(n24035), .Z(n24038) );
  ANDN U26395 ( .B(n24038), .A(n24037), .Z(n24040) );
  NANDN U26396 ( .A(n24040), .B(n24039), .Z(n24042) );
  ANDN U26397 ( .B(n24042), .A(n24041), .Z(n24044) );
  NANDN U26398 ( .A(n24044), .B(n24043), .Z(n24045) );
  AND U26399 ( .A(n24046), .B(n24045), .Z(n24047) );
  NAND U26400 ( .A(n24048), .B(n24047), .Z(n24049) );
  NAND U26401 ( .A(n24050), .B(n24049), .Z(n24052) );
  ANDN U26402 ( .B(n24052), .A(n24051), .Z(n24053) );
  OR U26403 ( .A(n24054), .B(n24053), .Z(n24056) );
  ANDN U26404 ( .B(n24056), .A(n24055), .Z(n24057) );
  ANDN U26405 ( .B(n24058), .A(n24057), .Z(n24060) );
  NANDN U26406 ( .A(n24060), .B(n24059), .Z(n24061) );
  NANDN U26407 ( .A(n24062), .B(n24061), .Z(n24064) );
  NAND U26408 ( .A(n24064), .B(n24063), .Z(n24065) );
  NANDN U26409 ( .A(n24066), .B(n24065), .Z(n24068) );
  NAND U26410 ( .A(n24068), .B(n24067), .Z(n24069) );
  AND U26411 ( .A(n24070), .B(n24069), .Z(n24072) );
  OR U26412 ( .A(n24072), .B(n24071), .Z(n24073) );
  AND U26413 ( .A(n24074), .B(n24073), .Z(n24076) );
  NANDN U26414 ( .A(n24076), .B(n24075), .Z(n24078) );
  NAND U26415 ( .A(n24078), .B(n24077), .Z(n24080) );
  ANDN U26416 ( .B(n24080), .A(n24079), .Z(n24081) );
  OR U26417 ( .A(n24082), .B(n24081), .Z(n24084) );
  NAND U26418 ( .A(n24084), .B(n24083), .Z(n24086) );
  NAND U26419 ( .A(n24086), .B(n24085), .Z(n24088) );
  ANDN U26420 ( .B(n24088), .A(n24087), .Z(n24090) );
  NANDN U26421 ( .A(n24090), .B(n24089), .Z(n24091) );
  NANDN U26422 ( .A(n24092), .B(n24091), .Z(n24094) );
  NAND U26423 ( .A(n24094), .B(n24093), .Z(n24096) );
  NAND U26424 ( .A(n24096), .B(n24095), .Z(n24098) );
  NAND U26425 ( .A(n24098), .B(n24097), .Z(n24100) );
  ANDN U26426 ( .B(n24100), .A(n24099), .Z(n24102) );
  NANDN U26427 ( .A(n24102), .B(n24101), .Z(n24104) );
  NAND U26428 ( .A(n24104), .B(n24103), .Z(n24106) );
  NAND U26429 ( .A(n24106), .B(n24105), .Z(n24108) );
  NAND U26430 ( .A(n24108), .B(n24107), .Z(n24110) );
  NAND U26431 ( .A(n24110), .B(n24109), .Z(n24111) );
  AND U26432 ( .A(n24112), .B(n24111), .Z(n24114) );
  NANDN U26433 ( .A(n24114), .B(n24113), .Z(n24116) );
  NAND U26434 ( .A(n24116), .B(n24115), .Z(n24118) );
  NAND U26435 ( .A(n24118), .B(n24117), .Z(n24119) );
  NANDN U26436 ( .A(n24120), .B(n24119), .Z(n24122) );
  NAND U26437 ( .A(n24122), .B(n24121), .Z(n24124) );
  ANDN U26438 ( .B(n24124), .A(n24123), .Z(n24126) );
  NANDN U26439 ( .A(n24126), .B(n24125), .Z(n24127) );
  AND U26440 ( .A(n24128), .B(n24127), .Z(n24130) );
  NANDN U26441 ( .A(n24130), .B(n24129), .Z(n24131) );
  NANDN U26442 ( .A(n24132), .B(n24131), .Z(n24134) );
  NAND U26443 ( .A(n24134), .B(n24133), .Z(n24136) );
  ANDN U26444 ( .B(n24136), .A(n24135), .Z(n24137) );
  NANDN U26445 ( .A(n24138), .B(n24137), .Z(n24139) );
  NANDN U26446 ( .A(n24140), .B(n24139), .Z(n24142) );
  ANDN U26447 ( .B(n24142), .A(n24141), .Z(n24144) );
  NANDN U26448 ( .A(n24144), .B(n24143), .Z(n24146) );
  NAND U26449 ( .A(n24146), .B(n24145), .Z(n24147) );
  NANDN U26450 ( .A(n24148), .B(n24147), .Z(n24150) );
  NAND U26451 ( .A(n24150), .B(n24149), .Z(n24152) );
  NAND U26452 ( .A(n24152), .B(n24151), .Z(n24153) );
  AND U26453 ( .A(n24154), .B(n24153), .Z(n24156) );
  NANDN U26454 ( .A(n24156), .B(n24155), .Z(n24157) );
  NANDN U26455 ( .A(n24158), .B(n24157), .Z(n24160) );
  NAND U26456 ( .A(n24160), .B(n24159), .Z(n24161) );
  NANDN U26457 ( .A(n24162), .B(n24161), .Z(n24164) );
  NAND U26458 ( .A(n24164), .B(n24163), .Z(n24165) );
  NANDN U26459 ( .A(n24166), .B(n24165), .Z(n24167) );
  NANDN U26460 ( .A(n24168), .B(n24167), .Z(n24170) );
  NAND U26461 ( .A(n24170), .B(n24169), .Z(n24171) );
  AND U26462 ( .A(n24172), .B(n24171), .Z(n24174) );
  NANDN U26463 ( .A(n24174), .B(n24173), .Z(n24175) );
  NANDN U26464 ( .A(n24176), .B(n24175), .Z(n24178) );
  NAND U26465 ( .A(n24178), .B(n24177), .Z(n24180) );
  NANDN U26466 ( .A(n24180), .B(n24179), .Z(n24182) );
  ANDN U26467 ( .B(n24182), .A(n24181), .Z(n24184) );
  NANDN U26468 ( .A(n24184), .B(n24183), .Z(n24186) );
  NAND U26469 ( .A(n24186), .B(n24185), .Z(n24188) );
  NAND U26470 ( .A(n24188), .B(n24187), .Z(n24190) );
  NAND U26471 ( .A(n24190), .B(n24189), .Z(n24192) );
  ANDN U26472 ( .B(n24192), .A(n24191), .Z(n24194) );
  NANDN U26473 ( .A(n24194), .B(n24193), .Z(n24196) );
  NAND U26474 ( .A(n24196), .B(n24195), .Z(n24197) );
  AND U26475 ( .A(n24198), .B(n24197), .Z(n24199) );
  OR U26476 ( .A(n24200), .B(n24199), .Z(n24201) );
  NANDN U26477 ( .A(n24202), .B(n24201), .Z(n24204) );
  NAND U26478 ( .A(n24204), .B(n24203), .Z(n24206) );
  NAND U26479 ( .A(n24206), .B(n24205), .Z(n24208) );
  NAND U26480 ( .A(n24208), .B(n24207), .Z(n24210) );
  ANDN U26481 ( .B(n24210), .A(n24209), .Z(n24212) );
  OR U26482 ( .A(n24212), .B(n24211), .Z(n24213) );
  AND U26483 ( .A(n24214), .B(n24213), .Z(n24216) );
  NANDN U26484 ( .A(n24216), .B(n24215), .Z(n24217) );
  NANDN U26485 ( .A(n24218), .B(n24217), .Z(n24220) );
  NAND U26486 ( .A(n24220), .B(n24219), .Z(n24221) );
  NANDN U26487 ( .A(n24222), .B(n24221), .Z(n24224) );
  NAND U26488 ( .A(n24224), .B(n24223), .Z(n24226) );
  NAND U26489 ( .A(n24226), .B(n24225), .Z(n24227) );
  NAND U26490 ( .A(n24228), .B(n24227), .Z(n24229) );
  NANDN U26491 ( .A(n24230), .B(n24229), .Z(n24231) );
  AND U26492 ( .A(n24232), .B(n24231), .Z(n24234) );
  NANDN U26493 ( .A(n24234), .B(n24233), .Z(n24235) );
  NANDN U26494 ( .A(n24236), .B(n24235), .Z(n24238) );
  NAND U26495 ( .A(n24238), .B(n24237), .Z(n24239) );
  NANDN U26496 ( .A(n24240), .B(n24239), .Z(n24242) );
  NAND U26497 ( .A(n24242), .B(n24241), .Z(n24244) );
  ANDN U26498 ( .B(n24244), .A(n24243), .Z(n24246) );
  NANDN U26499 ( .A(n24246), .B(n24245), .Z(n24247) );
  NANDN U26500 ( .A(n24248), .B(n24247), .Z(n24250) );
  NAND U26501 ( .A(n24250), .B(n24249), .Z(n24252) );
  NAND U26502 ( .A(n24252), .B(n24251), .Z(n24254) );
  ANDN U26503 ( .B(n24254), .A(n24253), .Z(n24256) );
  NANDN U26504 ( .A(n24256), .B(n24255), .Z(n24258) );
  NAND U26505 ( .A(n24258), .B(n24257), .Z(n24259) );
  NANDN U26506 ( .A(n24260), .B(n24259), .Z(n24262) );
  NAND U26507 ( .A(n24262), .B(n24261), .Z(n24263) );
  AND U26508 ( .A(n24264), .B(n24263), .Z(n24266) );
  NANDN U26509 ( .A(n24266), .B(n24265), .Z(n24268) );
  ANDN U26510 ( .B(n24268), .A(n24267), .Z(n24270) );
  NANDN U26511 ( .A(n24270), .B(n24269), .Z(n24272) );
  NAND U26512 ( .A(n24272), .B(n24271), .Z(n24274) );
  NAND U26513 ( .A(n24274), .B(n24273), .Z(n24275) );
  NAND U26514 ( .A(n24276), .B(n24275), .Z(n24279) );
  XOR U26515 ( .A(n24276), .B(n24275), .Z(n24277) );
  NAND U26516 ( .A(n24277), .B(y[2117]), .Z(n24278) );
  NAND U26517 ( .A(n24279), .B(n24278), .Z(n24280) );
  AND U26518 ( .A(n24281), .B(n24280), .Z(n24283) );
  NANDN U26519 ( .A(n24283), .B(n24282), .Z(n24284) );
  AND U26520 ( .A(n24285), .B(n24284), .Z(n24286) );
  OR U26521 ( .A(n24287), .B(n24286), .Z(n24289) );
  NAND U26522 ( .A(n24289), .B(n24288), .Z(n24291) );
  ANDN U26523 ( .B(n24291), .A(n24290), .Z(n24293) );
  NANDN U26524 ( .A(n24293), .B(n24292), .Z(n24295) );
  NAND U26525 ( .A(n24295), .B(n24294), .Z(n24297) );
  NAND U26526 ( .A(n24297), .B(n24296), .Z(n24299) );
  NAND U26527 ( .A(n24299), .B(n24298), .Z(n24301) );
  AND U26528 ( .A(n24301), .B(n24300), .Z(n24303) );
  NANDN U26529 ( .A(n24303), .B(n24302), .Z(n24304) );
  NANDN U26530 ( .A(n24305), .B(n24304), .Z(n24307) );
  NAND U26531 ( .A(n24307), .B(n24306), .Z(n24309) );
  NAND U26532 ( .A(n24309), .B(n24308), .Z(n24311) );
  NAND U26533 ( .A(n24311), .B(n24310), .Z(n24313) );
  ANDN U26534 ( .B(n24313), .A(n24312), .Z(n24315) );
  NANDN U26535 ( .A(n24315), .B(n24314), .Z(n24316) );
  NAND U26536 ( .A(n24317), .B(n24316), .Z(n24319) );
  NAND U26537 ( .A(n24319), .B(n24318), .Z(n24321) );
  NAND U26538 ( .A(n24321), .B(n24320), .Z(n24323) );
  ANDN U26539 ( .B(n24323), .A(n24322), .Z(n24324) );
  ANDN U26540 ( .B(n24325), .A(n24324), .Z(n24327) );
  NANDN U26541 ( .A(n24327), .B(n24326), .Z(n24328) );
  NANDN U26542 ( .A(n24329), .B(n24328), .Z(n24331) );
  NAND U26543 ( .A(n24331), .B(n24330), .Z(n24332) );
  AND U26544 ( .A(n24333), .B(n24332), .Z(n24335) );
  NANDN U26545 ( .A(n24335), .B(n24334), .Z(n24337) );
  NAND U26546 ( .A(n24337), .B(n24336), .Z(n24339) );
  NAND U26547 ( .A(n24339), .B(n24338), .Z(n24340) );
  AND U26548 ( .A(n24341), .B(n24340), .Z(n24343) );
  NANDN U26549 ( .A(n24343), .B(n24342), .Z(n24345) );
  NAND U26550 ( .A(n24345), .B(n24344), .Z(n24347) );
  NAND U26551 ( .A(n24347), .B(n24346), .Z(n24349) );
  NAND U26552 ( .A(n24349), .B(n24348), .Z(n24350) );
  NANDN U26553 ( .A(n24351), .B(n24350), .Z(n24353) );
  NAND U26554 ( .A(n24353), .B(n24352), .Z(n24354) );
  AND U26555 ( .A(n24355), .B(n24354), .Z(n24356) );
  ANDN U26556 ( .B(n24357), .A(n24356), .Z(n24358) );
  OR U26557 ( .A(n24359), .B(n24358), .Z(n24360) );
  NANDN U26558 ( .A(n24361), .B(n24360), .Z(n24362) );
  NANDN U26559 ( .A(n24363), .B(n24362), .Z(n24364) );
  NAND U26560 ( .A(n24365), .B(n24364), .Z(n24367) );
  NANDN U26561 ( .A(n24367), .B(n24366), .Z(n24369) );
  NAND U26562 ( .A(n24369), .B(n24368), .Z(n24371) );
  NAND U26563 ( .A(n24371), .B(n24370), .Z(n24373) );
  NAND U26564 ( .A(n24373), .B(n24372), .Z(n24375) );
  NAND U26565 ( .A(n24375), .B(n24374), .Z(n24376) );
  AND U26566 ( .A(n24377), .B(n24376), .Z(n24379) );
  NANDN U26567 ( .A(n24379), .B(n24378), .Z(n24380) );
  NANDN U26568 ( .A(n24381), .B(n24380), .Z(n24383) );
  NAND U26569 ( .A(n24383), .B(n24382), .Z(n24385) );
  NAND U26570 ( .A(n24385), .B(n24384), .Z(n24387) );
  NAND U26571 ( .A(n24387), .B(n24386), .Z(n24389) );
  NAND U26572 ( .A(n24389), .B(n24388), .Z(n24391) );
  ANDN U26573 ( .B(n24391), .A(n24390), .Z(n24392) );
  OR U26574 ( .A(n24393), .B(n24392), .Z(n24395) );
  NAND U26575 ( .A(n24395), .B(n24394), .Z(n24396) );
  AND U26576 ( .A(n24397), .B(n24396), .Z(n24398) );
  OR U26577 ( .A(n24399), .B(n24398), .Z(n24400) );
  NANDN U26578 ( .A(n24401), .B(n24400), .Z(n24402) );
  NANDN U26579 ( .A(n24403), .B(n24402), .Z(n24405) );
  NAND U26580 ( .A(n24405), .B(n24404), .Z(n24407) );
  ANDN U26581 ( .B(n24407), .A(n24406), .Z(n24409) );
  NANDN U26582 ( .A(n24409), .B(n24408), .Z(n24410) );
  NANDN U26583 ( .A(n24411), .B(n24410), .Z(n24412) );
  NANDN U26584 ( .A(n24413), .B(n24412), .Z(n24415) );
  NAND U26585 ( .A(n24415), .B(n24414), .Z(n24416) );
  AND U26586 ( .A(n24417), .B(n24416), .Z(n24419) );
  NANDN U26587 ( .A(n24419), .B(n24418), .Z(n24421) );
  ANDN U26588 ( .B(n24421), .A(n24420), .Z(n24423) );
  OR U26589 ( .A(n24423), .B(n24422), .Z(n24424) );
  NANDN U26590 ( .A(n24425), .B(n24424), .Z(n24427) );
  ANDN U26591 ( .B(n24427), .A(n24426), .Z(n24429) );
  NANDN U26592 ( .A(n24429), .B(n24428), .Z(n24430) );
  AND U26593 ( .A(n24431), .B(n24430), .Z(n24432) );
  NAND U26594 ( .A(n24433), .B(n24432), .Z(n24434) );
  NAND U26595 ( .A(n24435), .B(n24434), .Z(n24436) );
  NANDN U26596 ( .A(n24437), .B(n24436), .Z(n24439) );
  NAND U26597 ( .A(n24439), .B(n24438), .Z(n24440) );
  AND U26598 ( .A(n24441), .B(n24440), .Z(n24443) );
  NANDN U26599 ( .A(n24443), .B(n24442), .Z(n24445) );
  ANDN U26600 ( .B(n24445), .A(n24444), .Z(n24447) );
  NANDN U26601 ( .A(n24447), .B(n24446), .Z(n24448) );
  NANDN U26602 ( .A(n24449), .B(n24448), .Z(n24451) );
  NAND U26603 ( .A(n24451), .B(n24450), .Z(n24453) );
  NAND U26604 ( .A(n24453), .B(n24452), .Z(n24455) );
  NAND U26605 ( .A(n24455), .B(n24454), .Z(n24456) );
  NANDN U26606 ( .A(n24457), .B(n24456), .Z(n24458) );
  NANDN U26607 ( .A(n24459), .B(n24458), .Z(n24461) );
  NAND U26608 ( .A(n24461), .B(n24460), .Z(n24463) );
  ANDN U26609 ( .B(n24463), .A(n24462), .Z(n24464) );
  OR U26610 ( .A(n24465), .B(n24464), .Z(n24467) );
  ANDN U26611 ( .B(n24467), .A(n24466), .Z(n24471) );
  AND U26612 ( .A(n24469), .B(n24468), .Z(n24470) );
  NANDN U26613 ( .A(n24471), .B(n24470), .Z(n24472) );
  AND U26614 ( .A(n24473), .B(n24472), .Z(n24475) );
  NANDN U26615 ( .A(n24475), .B(n24474), .Z(n24477) );
  ANDN U26616 ( .B(n24477), .A(n24476), .Z(n24479) );
  NANDN U26617 ( .A(n24479), .B(n24478), .Z(n24481) );
  ANDN U26618 ( .B(n24481), .A(n24480), .Z(n24483) );
  NANDN U26619 ( .A(n24483), .B(n24482), .Z(n24484) );
  NANDN U26620 ( .A(n24485), .B(n24484), .Z(n24487) );
  NAND U26621 ( .A(n24487), .B(n24486), .Z(n24489) );
  ANDN U26622 ( .B(n24489), .A(n24488), .Z(n24491) );
  OR U26623 ( .A(n24491), .B(n24490), .Z(n24492) );
  NANDN U26624 ( .A(n24493), .B(n24492), .Z(n24494) );
  NANDN U26625 ( .A(n24495), .B(n24494), .Z(n24497) );
  ANDN U26626 ( .B(n24497), .A(n24496), .Z(n24499) );
  NANDN U26627 ( .A(n24499), .B(n24498), .Z(n24501) );
  ANDN U26628 ( .B(n24501), .A(n24500), .Z(n24503) );
  NANDN U26629 ( .A(n24503), .B(n24502), .Z(n24504) );
  AND U26630 ( .A(n24505), .B(n24504), .Z(n24506) );
  NAND U26631 ( .A(n24507), .B(n24506), .Z(n24508) );
  NAND U26632 ( .A(n24509), .B(n24508), .Z(n24511) );
  ANDN U26633 ( .B(n24511), .A(n24510), .Z(n24513) );
  NANDN U26634 ( .A(n24513), .B(n24512), .Z(n24515) );
  NAND U26635 ( .A(n24515), .B(n24514), .Z(n24517) );
  NAND U26636 ( .A(n24517), .B(n24516), .Z(n24519) );
  NAND U26637 ( .A(n24519), .B(n24518), .Z(n24520) );
  NANDN U26638 ( .A(n24521), .B(n24520), .Z(n24523) );
  NAND U26639 ( .A(n24523), .B(n24522), .Z(n24525) );
  AND U26640 ( .A(n24525), .B(n24524), .Z(n24527) );
  NAND U26641 ( .A(n24527), .B(n24526), .Z(n24529) );
  NAND U26642 ( .A(n24529), .B(n24528), .Z(n24530) );
  NAND U26643 ( .A(n24531), .B(n24530), .Z(n24532) );
  NAND U26644 ( .A(n24533), .B(n24532), .Z(n24534) );
  NAND U26645 ( .A(n24535), .B(n24534), .Z(n24536) );
  NAND U26646 ( .A(n24537), .B(n24536), .Z(n24538) );
  AND U26647 ( .A(n24539), .B(n24538), .Z(n24541) );
  NANDN U26648 ( .A(n24541), .B(n24540), .Z(n24543) );
  NAND U26649 ( .A(n24543), .B(n24542), .Z(n24545) );
  NAND U26650 ( .A(n24545), .B(n24544), .Z(n24546) );
  AND U26651 ( .A(n24547), .B(n24546), .Z(n24548) );
  OR U26652 ( .A(n24549), .B(n24548), .Z(n24551) );
  NAND U26653 ( .A(n24551), .B(n24550), .Z(n24553) );
  ANDN U26654 ( .B(n24553), .A(n24552), .Z(n24555) );
  NANDN U26655 ( .A(n24555), .B(n24554), .Z(n24556) );
  AND U26656 ( .A(n24557), .B(n24556), .Z(n24559) );
  OR U26657 ( .A(n24559), .B(n24558), .Z(n24560) );
  AND U26658 ( .A(n24561), .B(n24560), .Z(n24563) );
  NANDN U26659 ( .A(n24563), .B(n24562), .Z(n24564) );
  AND U26660 ( .A(n24565), .B(n24564), .Z(n24567) );
  NANDN U26661 ( .A(n24567), .B(n24566), .Z(n24568) );
  NANDN U26662 ( .A(n24569), .B(n24568), .Z(n24571) );
  NAND U26663 ( .A(n24571), .B(n24570), .Z(n24572) );
  AND U26664 ( .A(n24573), .B(n24572), .Z(n24575) );
  NANDN U26665 ( .A(n24575), .B(n24574), .Z(n24577) );
  NAND U26666 ( .A(n24577), .B(n24576), .Z(n24578) );
  AND U26667 ( .A(n24579), .B(n24578), .Z(n24581) );
  NANDN U26668 ( .A(n24581), .B(n24580), .Z(n24583) );
  NAND U26669 ( .A(n24583), .B(n24582), .Z(n24585) );
  NAND U26670 ( .A(n24585), .B(n24584), .Z(n24587) );
  ANDN U26671 ( .B(n24587), .A(n24586), .Z(n24589) );
  NANDN U26672 ( .A(n24589), .B(n24588), .Z(n24590) );
  AND U26673 ( .A(n24591), .B(n24590), .Z(n24593) );
  NANDN U26674 ( .A(n24593), .B(n24592), .Z(n24594) );
  NANDN U26675 ( .A(n24595), .B(n24594), .Z(n24597) );
  NAND U26676 ( .A(n24597), .B(n24596), .Z(n24599) );
  ANDN U26677 ( .B(n24599), .A(n24598), .Z(n24601) );
  NANDN U26678 ( .A(n24601), .B(n24600), .Z(n24602) );
  NANDN U26679 ( .A(n24603), .B(n24602), .Z(n24605) );
  NAND U26680 ( .A(n24605), .B(n24604), .Z(n24607) );
  ANDN U26681 ( .B(n24607), .A(n24606), .Z(n24609) );
  NANDN U26682 ( .A(n24609), .B(n24608), .Z(n24611) );
  NAND U26683 ( .A(n24611), .B(n24610), .Z(n24613) );
  ANDN U26684 ( .B(n24613), .A(n24612), .Z(n24615) );
  NANDN U26685 ( .A(n24615), .B(n24614), .Z(n24617) );
  NAND U26686 ( .A(n24617), .B(n24616), .Z(n24619) );
  NAND U26687 ( .A(n24619), .B(n24618), .Z(n24620) );
  AND U26688 ( .A(n24621), .B(n24620), .Z(n24622) );
  OR U26689 ( .A(n24623), .B(n24622), .Z(n24625) );
  NAND U26690 ( .A(n24625), .B(n24624), .Z(n24627) );
  NAND U26691 ( .A(n24627), .B(n24626), .Z(n24629) );
  ANDN U26692 ( .B(n24629), .A(n24628), .Z(n24630) );
  OR U26693 ( .A(n24631), .B(n24630), .Z(n24632) );
  NANDN U26694 ( .A(n24633), .B(n24632), .Z(n24635) );
  NAND U26695 ( .A(n24635), .B(n24634), .Z(n24637) );
  ANDN U26696 ( .B(n24637), .A(n24636), .Z(n24639) );
  NANDN U26697 ( .A(n24639), .B(n24638), .Z(n24640) );
  NANDN U26698 ( .A(n24641), .B(n24640), .Z(n24643) );
  NAND U26699 ( .A(n24643), .B(n24642), .Z(n24644) );
  NANDN U26700 ( .A(n24645), .B(n24644), .Z(n24647) );
  NAND U26701 ( .A(n24647), .B(n24646), .Z(n24648) );
  AND U26702 ( .A(n24649), .B(n24648), .Z(n24651) );
  NANDN U26703 ( .A(n24651), .B(n24650), .Z(n24653) );
  ANDN U26704 ( .B(n24653), .A(n24652), .Z(n24655) );
  NANDN U26705 ( .A(n24655), .B(n24654), .Z(n24656) );
  NANDN U26706 ( .A(n24657), .B(n24656), .Z(n24659) );
  NAND U26707 ( .A(n24659), .B(n24658), .Z(n24661) );
  NANDN U26708 ( .A(n24661), .B(n24660), .Z(n24662) );
  NANDN U26709 ( .A(n24663), .B(n24662), .Z(n24665) );
  NAND U26710 ( .A(n24665), .B(n24664), .Z(n24666) );
  AND U26711 ( .A(n24667), .B(n24666), .Z(n24669) );
  NANDN U26712 ( .A(n24669), .B(n24668), .Z(n24671) );
  NAND U26713 ( .A(n24671), .B(n24670), .Z(n24673) );
  NAND U26714 ( .A(n24673), .B(n24672), .Z(n24674) );
  AND U26715 ( .A(n24675), .B(n24674), .Z(n24677) );
  NANDN U26716 ( .A(n24677), .B(n24676), .Z(n24678) );
  NANDN U26717 ( .A(n24679), .B(n24678), .Z(n24681) );
  NAND U26718 ( .A(n24681), .B(n24680), .Z(n24683) );
  ANDN U26719 ( .B(n24683), .A(n24682), .Z(n24685) );
  NANDN U26720 ( .A(n24685), .B(n24684), .Z(n24687) );
  NAND U26721 ( .A(n24687), .B(n24686), .Z(n24689) );
  NAND U26722 ( .A(n24689), .B(n24688), .Z(n24690) );
  AND U26723 ( .A(n24691), .B(n24690), .Z(n24692) );
  OR U26724 ( .A(n24693), .B(n24692), .Z(n24695) );
  NAND U26725 ( .A(n24695), .B(n24694), .Z(n24696) );
  AND U26726 ( .A(n24697), .B(n24696), .Z(n24699) );
  NANDN U26727 ( .A(n24699), .B(n24698), .Z(n24700) );
  AND U26728 ( .A(n24701), .B(n24700), .Z(n24703) );
  NANDN U26729 ( .A(n24703), .B(n24702), .Z(n24704) );
  AND U26730 ( .A(n24705), .B(n24704), .Z(n24707) );
  NANDN U26731 ( .A(n24707), .B(n24706), .Z(n24709) );
  NAND U26732 ( .A(n24709), .B(n24708), .Z(n24711) );
  NAND U26733 ( .A(n24711), .B(n24710), .Z(n24712) );
  AND U26734 ( .A(n24713), .B(n24712), .Z(n24714) );
  NANDN U26735 ( .A(n24715), .B(n24714), .Z(n24717) );
  NAND U26736 ( .A(n24717), .B(n24716), .Z(n24718) );
  AND U26737 ( .A(n24719), .B(n24718), .Z(n24720) );
  NANDN U26738 ( .A(n24721), .B(n24720), .Z(n24723) );
  NAND U26739 ( .A(n24723), .B(n24722), .Z(n24725) );
  ANDN U26740 ( .B(n24725), .A(n24724), .Z(n24727) );
  NANDN U26741 ( .A(n24727), .B(n24726), .Z(n24728) );
  AND U26742 ( .A(n24729), .B(n24728), .Z(n24731) );
  NANDN U26743 ( .A(n24731), .B(n24730), .Z(n24732) );
  AND U26744 ( .A(n24733), .B(n24732), .Z(n24734) );
  OR U26745 ( .A(n24735), .B(n24734), .Z(n24737) );
  NAND U26746 ( .A(n24737), .B(n24736), .Z(n24739) );
  ANDN U26747 ( .B(n24739), .A(n24738), .Z(n24741) );
  NANDN U26748 ( .A(n24741), .B(n24740), .Z(n24742) );
  NANDN U26749 ( .A(n24743), .B(n24742), .Z(n24745) );
  NAND U26750 ( .A(n24745), .B(n24744), .Z(n24746) );
  NANDN U26751 ( .A(n24747), .B(n24746), .Z(n24748) );
  NANDN U26752 ( .A(n24749), .B(n24748), .Z(n24751) );
  NAND U26753 ( .A(n24751), .B(n24750), .Z(n24753) );
  ANDN U26754 ( .B(n24753), .A(n24752), .Z(n24754) );
  OR U26755 ( .A(n24755), .B(n24754), .Z(n24757) );
  NAND U26756 ( .A(n24757), .B(n24756), .Z(n24759) );
  ANDN U26757 ( .B(n24759), .A(n24758), .Z(n24761) );
  NANDN U26758 ( .A(n24761), .B(n24760), .Z(n24762) );
  NANDN U26759 ( .A(n24763), .B(n24762), .Z(n24765) );
  NAND U26760 ( .A(n24765), .B(n24764), .Z(n24766) );
  NAND U26761 ( .A(n24767), .B(n24766), .Z(n24770) );
  XOR U26762 ( .A(n24767), .B(n24766), .Z(n24768) );
  NAND U26763 ( .A(n24768), .B(x[2328]), .Z(n24769) );
  NAND U26764 ( .A(n24770), .B(n24769), .Z(n24771) );
  AND U26765 ( .A(n24772), .B(n24771), .Z(n24774) );
  NANDN U26766 ( .A(n24774), .B(n24773), .Z(n24776) );
  NAND U26767 ( .A(n24776), .B(n24775), .Z(n24778) );
  ANDN U26768 ( .B(n24778), .A(n24777), .Z(n24780) );
  NANDN U26769 ( .A(n24780), .B(n24779), .Z(n24781) );
  AND U26770 ( .A(n24782), .B(n24781), .Z(n24784) );
  NANDN U26771 ( .A(n24784), .B(n24783), .Z(n24785) );
  NANDN U26772 ( .A(n24786), .B(n24785), .Z(n24788) );
  NAND U26773 ( .A(n24788), .B(n24787), .Z(n24789) );
  AND U26774 ( .A(n24790), .B(n24789), .Z(n24792) );
  NANDN U26775 ( .A(n24792), .B(n24791), .Z(n24793) );
  NANDN U26776 ( .A(n24794), .B(n24793), .Z(n24796) );
  NAND U26777 ( .A(n24796), .B(n24795), .Z(n24797) );
  AND U26778 ( .A(n24798), .B(n24797), .Z(n24800) );
  NANDN U26779 ( .A(n24800), .B(n24799), .Z(n24801) );
  NANDN U26780 ( .A(n24802), .B(n24801), .Z(n24804) );
  NAND U26781 ( .A(n24804), .B(n24803), .Z(n24805) );
  AND U26782 ( .A(n24806), .B(n24805), .Z(n24808) );
  NANDN U26783 ( .A(n24808), .B(n24807), .Z(n24809) );
  NANDN U26784 ( .A(n24810), .B(n24809), .Z(n24812) );
  NAND U26785 ( .A(n24812), .B(n24811), .Z(n24814) );
  NAND U26786 ( .A(n24814), .B(n24813), .Z(n24816) );
  NAND U26787 ( .A(n24816), .B(n24815), .Z(n24817) );
  AND U26788 ( .A(n24818), .B(n24817), .Z(n24820) );
  NANDN U26789 ( .A(n24820), .B(n24819), .Z(n24821) );
  NANDN U26790 ( .A(n24822), .B(n24821), .Z(n24823) );
  NANDN U26791 ( .A(n24824), .B(n24823), .Z(n24825) );
  AND U26792 ( .A(n24826), .B(n24825), .Z(n24828) );
  NANDN U26793 ( .A(n24828), .B(n24827), .Z(n24830) );
  NAND U26794 ( .A(n24830), .B(n24829), .Z(n24832) );
  NAND U26795 ( .A(n24832), .B(n24831), .Z(n24834) );
  NAND U26796 ( .A(n24834), .B(n24833), .Z(n24836) );
  ANDN U26797 ( .B(n24836), .A(n24835), .Z(n24838) );
  NANDN U26798 ( .A(n24838), .B(n24837), .Z(n24839) );
  AND U26799 ( .A(n24840), .B(n24839), .Z(n24842) );
  NANDN U26800 ( .A(n24842), .B(n24841), .Z(n24843) );
  NANDN U26801 ( .A(n24844), .B(n24843), .Z(n24846) );
  NAND U26802 ( .A(n24846), .B(n24845), .Z(n24848) );
  NAND U26803 ( .A(n24848), .B(n24847), .Z(n24850) );
  ANDN U26804 ( .B(n24850), .A(n24849), .Z(n24851) );
  NANDN U26805 ( .A(n24852), .B(n24851), .Z(n24854) );
  NAND U26806 ( .A(n24854), .B(n24853), .Z(n24856) );
  ANDN U26807 ( .B(n24856), .A(n24855), .Z(n24858) );
  OR U26808 ( .A(n24858), .B(n24857), .Z(n24860) );
  ANDN U26809 ( .B(n24860), .A(n24859), .Z(n24862) );
  NANDN U26810 ( .A(n24862), .B(n24861), .Z(n24863) );
  AND U26811 ( .A(n24864), .B(n24863), .Z(n24866) );
  NANDN U26812 ( .A(n24866), .B(n24865), .Z(n24868) );
  NAND U26813 ( .A(n24868), .B(n24867), .Z(n24870) );
  NAND U26814 ( .A(n24870), .B(n24869), .Z(n24871) );
  AND U26815 ( .A(n24872), .B(n24871), .Z(n24874) );
  NANDN U26816 ( .A(n24874), .B(n24873), .Z(n24876) );
  ANDN U26817 ( .B(n24876), .A(n24875), .Z(n24877) );
  NANDN U26818 ( .A(n24878), .B(n24877), .Z(n24880) );
  NAND U26819 ( .A(n24880), .B(n24879), .Z(n24882) );
  ANDN U26820 ( .B(n24882), .A(n24881), .Z(n24884) );
  NANDN U26821 ( .A(n24884), .B(n24883), .Z(n24886) );
  NAND U26822 ( .A(n24886), .B(n24885), .Z(n24888) );
  NAND U26823 ( .A(n24888), .B(n24887), .Z(n24890) );
  NAND U26824 ( .A(n24890), .B(n24889), .Z(n24892) );
  ANDN U26825 ( .B(n24892), .A(n24891), .Z(n24894) );
  NANDN U26826 ( .A(n24894), .B(n24893), .Z(n24896) );
  NAND U26827 ( .A(n24896), .B(n24895), .Z(n24897) );
  NANDN U26828 ( .A(n24898), .B(n24897), .Z(n24899) );
  NANDN U26829 ( .A(n24900), .B(n24899), .Z(n24902) );
  NAND U26830 ( .A(n24902), .B(n24901), .Z(n24904) );
  NAND U26831 ( .A(n24904), .B(n24903), .Z(n24906) );
  ANDN U26832 ( .B(n24906), .A(n24905), .Z(n24908) );
  OR U26833 ( .A(n24908), .B(n24907), .Z(n24910) );
  ANDN U26834 ( .B(n24910), .A(n24909), .Z(n24912) );
  NANDN U26835 ( .A(n24912), .B(n24911), .Z(n24913) );
  AND U26836 ( .A(n24914), .B(n24913), .Z(n24920) );
  NANDN U26837 ( .A(n24916), .B(n24915), .Z(n24918) );
  ANDN U26838 ( .B(n24918), .A(n24917), .Z(n24919) );
  NANDN U26839 ( .A(n24920), .B(n24919), .Z(n24922) );
  NAND U26840 ( .A(n24922), .B(n24921), .Z(n24924) );
  NAND U26841 ( .A(n24924), .B(n24923), .Z(n24926) );
  ANDN U26842 ( .B(n24926), .A(n24925), .Z(n24928) );
  NANDN U26843 ( .A(n24928), .B(n24927), .Z(n24930) );
  NAND U26844 ( .A(n24930), .B(n24929), .Z(n24932) );
  NAND U26845 ( .A(n24932), .B(n24931), .Z(n24933) );
  AND U26846 ( .A(n24934), .B(n24933), .Z(n24936) );
  NANDN U26847 ( .A(n24936), .B(n24935), .Z(n24938) );
  ANDN U26848 ( .B(n24938), .A(n24937), .Z(n24940) );
  NANDN U26849 ( .A(n24940), .B(n24939), .Z(n24941) );
  NANDN U26850 ( .A(n24942), .B(n24941), .Z(n24944) );
  NAND U26851 ( .A(n24944), .B(n24943), .Z(n24945) );
  AND U26852 ( .A(n24946), .B(n24945), .Z(n24948) );
  NANDN U26853 ( .A(n24948), .B(n24947), .Z(n24949) );
  NANDN U26854 ( .A(n24950), .B(n24949), .Z(n24952) );
  NAND U26855 ( .A(n24952), .B(n24951), .Z(n24954) );
  ANDN U26856 ( .B(n24954), .A(n24953), .Z(n24956) );
  NAND U26857 ( .A(n24956), .B(n24955), .Z(n24958) );
  NAND U26858 ( .A(n24958), .B(n24957), .Z(n24960) );
  NAND U26859 ( .A(n24960), .B(n24959), .Z(n24962) );
  ANDN U26860 ( .B(n24962), .A(n24961), .Z(n24964) );
  NANDN U26861 ( .A(n24964), .B(n24963), .Z(n24965) );
  AND U26862 ( .A(n24966), .B(n24965), .Z(n24968) );
  NANDN U26863 ( .A(n24968), .B(n24967), .Z(n24969) );
  AND U26864 ( .A(n24970), .B(n24969), .Z(n24972) );
  NANDN U26865 ( .A(n24972), .B(n24971), .Z(n24974) );
  NAND U26866 ( .A(n24974), .B(n24973), .Z(n24975) );
  AND U26867 ( .A(n24976), .B(n24975), .Z(n24978) );
  NANDN U26868 ( .A(n24978), .B(n24977), .Z(n24980) );
  ANDN U26869 ( .B(n24980), .A(n24979), .Z(n24981) );
  OR U26870 ( .A(n24982), .B(n24981), .Z(n24983) );
  NANDN U26871 ( .A(n24984), .B(n24983), .Z(n24986) );
  NAND U26872 ( .A(n24986), .B(n24985), .Z(n24988) );
  ANDN U26873 ( .B(n24988), .A(n24987), .Z(n24990) );
  NANDN U26874 ( .A(n24990), .B(n24989), .Z(n24991) );
  NANDN U26875 ( .A(n24992), .B(n24991), .Z(n24994) );
  NAND U26876 ( .A(n24994), .B(n24993), .Z(n24996) );
  ANDN U26877 ( .B(n24996), .A(n24995), .Z(n24998) );
  NAND U26878 ( .A(n24998), .B(n24997), .Z(n25000) );
  NAND U26879 ( .A(n25000), .B(n24999), .Z(n25002) );
  AND U26880 ( .A(n25002), .B(n25001), .Z(n25004) );
  NANDN U26881 ( .A(n25004), .B(n25003), .Z(n25006) );
  NAND U26882 ( .A(n25006), .B(n25005), .Z(n25007) );
  AND U26883 ( .A(n25008), .B(n25007), .Z(n25010) );
  NANDN U26884 ( .A(n25010), .B(n25009), .Z(n25012) );
  NAND U26885 ( .A(n25012), .B(n25011), .Z(n25014) );
  NAND U26886 ( .A(n25014), .B(n25013), .Z(n25016) );
  NANDN U26887 ( .A(n25016), .B(n25015), .Z(n25018) );
  ANDN U26888 ( .B(n25018), .A(n25017), .Z(n25020) );
  NANDN U26889 ( .A(n25020), .B(n25019), .Z(n25022) );
  ANDN U26890 ( .B(n25022), .A(n25021), .Z(n25024) );
  NANDN U26891 ( .A(n25024), .B(n25023), .Z(n25026) );
  ANDN U26892 ( .B(n25026), .A(n25025), .Z(n25027) );
  NAND U26893 ( .A(n25028), .B(n25027), .Z(n25029) );
  NAND U26894 ( .A(n25030), .B(n25029), .Z(n25031) );
  NANDN U26895 ( .A(n25032), .B(n25031), .Z(n25034) );
  NAND U26896 ( .A(n25034), .B(n25033), .Z(n25035) );
  AND U26897 ( .A(n25036), .B(n25035), .Z(n25038) );
  NANDN U26898 ( .A(n25038), .B(n25037), .Z(n25039) );
  NANDN U26899 ( .A(n25040), .B(n25039), .Z(n25042) );
  NAND U26900 ( .A(n25042), .B(n25041), .Z(n25044) );
  NAND U26901 ( .A(n25044), .B(n25043), .Z(n25046) );
  NAND U26902 ( .A(n25046), .B(n25045), .Z(n25048) );
  NAND U26903 ( .A(n25048), .B(n25047), .Z(n25050) );
  ANDN U26904 ( .B(n25050), .A(n25049), .Z(n25051) );
  NANDN U26905 ( .A(n25052), .B(n25051), .Z(n25054) );
  NAND U26906 ( .A(n25054), .B(n25053), .Z(n25056) );
  ANDN U26907 ( .B(n25056), .A(n25055), .Z(n25058) );
  NANDN U26908 ( .A(n25058), .B(n25057), .Z(n25059) );
  NANDN U26909 ( .A(n25060), .B(n25059), .Z(n25062) );
  NAND U26910 ( .A(n25062), .B(n25061), .Z(n25063) );
  NAND U26911 ( .A(n25064), .B(n25063), .Z(n25066) );
  NAND U26912 ( .A(n25066), .B(n25065), .Z(n25068) );
  ANDN U26913 ( .B(n25068), .A(n25067), .Z(n25070) );
  NANDN U26914 ( .A(n25070), .B(n25069), .Z(n25072) );
  NAND U26915 ( .A(n25072), .B(n25071), .Z(n25074) );
  NAND U26916 ( .A(n25074), .B(n25073), .Z(n25075) );
  AND U26917 ( .A(n25076), .B(n25075), .Z(n25078) );
  NANDN U26918 ( .A(n25078), .B(n25077), .Z(n25079) );
  NANDN U26919 ( .A(n25080), .B(n25079), .Z(n25081) );
  NANDN U26920 ( .A(n25082), .B(n25081), .Z(n25084) );
  ANDN U26921 ( .B(n25084), .A(n25083), .Z(n25086) );
  NANDN U26922 ( .A(n25086), .B(n25085), .Z(n25088) );
  NAND U26923 ( .A(n25088), .B(n25087), .Z(n25090) );
  NAND U26924 ( .A(n25090), .B(n25089), .Z(n25091) );
  AND U26925 ( .A(n25092), .B(n25091), .Z(n25094) );
  NANDN U26926 ( .A(n25094), .B(n25093), .Z(n25095) );
  AND U26927 ( .A(n25096), .B(n25095), .Z(n25098) );
  NANDN U26928 ( .A(n25098), .B(n25097), .Z(n25100) );
  NAND U26929 ( .A(n25100), .B(n25099), .Z(n25102) );
  NAND U26930 ( .A(n25102), .B(n25101), .Z(n25103) );
  AND U26931 ( .A(n25104), .B(n25103), .Z(n25106) );
  NANDN U26932 ( .A(n25106), .B(n25105), .Z(n25108) );
  NAND U26933 ( .A(n25108), .B(n25107), .Z(n25110) );
  NAND U26934 ( .A(n25110), .B(n25109), .Z(n25111) );
  AND U26935 ( .A(n25112), .B(n25111), .Z(n25114) );
  NANDN U26936 ( .A(n25114), .B(n25113), .Z(n25115) );
  NANDN U26937 ( .A(n25116), .B(n25115), .Z(n25118) );
  NAND U26938 ( .A(n25118), .B(n25117), .Z(n25119) );
  AND U26939 ( .A(n25120), .B(n25119), .Z(n25122) );
  NANDN U26940 ( .A(n25122), .B(n25121), .Z(n25124) );
  NAND U26941 ( .A(n25124), .B(n25123), .Z(n25126) );
  NAND U26942 ( .A(n25126), .B(n25125), .Z(n25127) );
  AND U26943 ( .A(n25128), .B(n25127), .Z(n25130) );
  NANDN U26944 ( .A(n25130), .B(n25129), .Z(n25132) );
  NAND U26945 ( .A(n25132), .B(n25131), .Z(n25134) );
  NAND U26946 ( .A(n25134), .B(n25133), .Z(n25135) );
  AND U26947 ( .A(n25136), .B(n25135), .Z(n25138) );
  NANDN U26948 ( .A(n25138), .B(n25137), .Z(n25139) );
  NANDN U26949 ( .A(n25140), .B(n25139), .Z(n25142) );
  NAND U26950 ( .A(n25142), .B(n25141), .Z(n25144) );
  NAND U26951 ( .A(n25144), .B(n25143), .Z(n25146) );
  NAND U26952 ( .A(n25146), .B(n25145), .Z(n25147) );
  AND U26953 ( .A(n25148), .B(n25147), .Z(n25150) );
  NANDN U26954 ( .A(n25150), .B(n25149), .Z(n25152) );
  ANDN U26955 ( .B(n25152), .A(n25151), .Z(n25154) );
  NANDN U26956 ( .A(n25154), .B(n25153), .Z(n25156) );
  NAND U26957 ( .A(n25156), .B(n25155), .Z(n25158) );
  NAND U26958 ( .A(n25158), .B(n25157), .Z(n25159) );
  AND U26959 ( .A(n25160), .B(n25159), .Z(n25162) );
  NAND U26960 ( .A(n25162), .B(n25161), .Z(n25163) );
  NANDN U26961 ( .A(n25164), .B(n25163), .Z(n25166) );
  NAND U26962 ( .A(n25166), .B(n25165), .Z(n25167) );
  AND U26963 ( .A(n25168), .B(n25167), .Z(n25170) );
  NANDN U26964 ( .A(n25170), .B(n25169), .Z(n25171) );
  NANDN U26965 ( .A(n25172), .B(n25171), .Z(n25174) );
  NAND U26966 ( .A(n25174), .B(n25173), .Z(n25176) );
  NAND U26967 ( .A(n25176), .B(n25175), .Z(n25178) );
  NAND U26968 ( .A(n25178), .B(n25177), .Z(n25179) );
  NANDN U26969 ( .A(n25180), .B(n25179), .Z(n25182) );
  ANDN U26970 ( .B(n25182), .A(n25181), .Z(n25184) );
  OR U26971 ( .A(n25184), .B(n25183), .Z(n25186) );
  NAND U26972 ( .A(n25186), .B(n25185), .Z(n25187) );
  AND U26973 ( .A(n25188), .B(n25187), .Z(n25190) );
  NANDN U26974 ( .A(n25190), .B(n25189), .Z(n25191) );
  NANDN U26975 ( .A(n25192), .B(n25191), .Z(n25194) );
  NAND U26976 ( .A(n25194), .B(n25193), .Z(n25195) );
  NANDN U26977 ( .A(n25196), .B(n25195), .Z(n25198) );
  NAND U26978 ( .A(n25198), .B(n25197), .Z(n25199) );
  NANDN U26979 ( .A(n25200), .B(n25199), .Z(n25201) );
  NANDN U26980 ( .A(n25202), .B(n25201), .Z(n25204) );
  NAND U26981 ( .A(n25204), .B(n25203), .Z(n25205) );
  AND U26982 ( .A(n25206), .B(n25205), .Z(n25208) );
  NANDN U26983 ( .A(n25208), .B(n25207), .Z(n25209) );
  NAND U26984 ( .A(n25210), .B(n25209), .Z(n25211) );
  NANDN U26985 ( .A(n25212), .B(n25211), .Z(n25213) );
  AND U26986 ( .A(n25214), .B(n25213), .Z(n25216) );
  NAND U26987 ( .A(n25216), .B(n25215), .Z(n25217) );
  AND U26988 ( .A(n25218), .B(n25217), .Z(n25220) );
  NANDN U26989 ( .A(n25220), .B(n25219), .Z(n25221) );
  AND U26990 ( .A(n25222), .B(n25221), .Z(n25224) );
  NANDN U26991 ( .A(n25224), .B(n25223), .Z(n25226) );
  NAND U26992 ( .A(n25226), .B(n25225), .Z(n25228) );
  NAND U26993 ( .A(n25228), .B(n25227), .Z(n25229) );
  NANDN U26994 ( .A(n25230), .B(n25229), .Z(n25232) );
  NAND U26995 ( .A(n25232), .B(n25231), .Z(n25233) );
  AND U26996 ( .A(n25234), .B(n25233), .Z(n25236) );
  NANDN U26997 ( .A(n25236), .B(n25235), .Z(n25238) );
  NAND U26998 ( .A(n25238), .B(n25237), .Z(n25240) );
  NAND U26999 ( .A(n25240), .B(n25239), .Z(n25242) );
  NAND U27000 ( .A(n25242), .B(n25241), .Z(n25244) );
  NAND U27001 ( .A(n25244), .B(n25243), .Z(n25245) );
  AND U27002 ( .A(n25246), .B(n25245), .Z(n25248) );
  NANDN U27003 ( .A(n25248), .B(n25247), .Z(n25250) );
  ANDN U27004 ( .B(n25250), .A(n25249), .Z(n25252) );
  NANDN U27005 ( .A(n25252), .B(n25251), .Z(n25253) );
  AND U27006 ( .A(n25254), .B(n25253), .Z(n25256) );
  NANDN U27007 ( .A(n25256), .B(n25255), .Z(n25258) );
  ANDN U27008 ( .B(n25258), .A(n25257), .Z(n25260) );
  NANDN U27009 ( .A(n25260), .B(n25259), .Z(n25262) );
  ANDN U27010 ( .B(n25262), .A(n25261), .Z(n25264) );
  NANDN U27011 ( .A(n25264), .B(n25263), .Z(n25266) );
  ANDN U27012 ( .B(n25266), .A(n25265), .Z(n25268) );
  NANDN U27013 ( .A(n25268), .B(n25267), .Z(n25270) );
  ANDN U27014 ( .B(n25270), .A(n25269), .Z(n25272) );
  NANDN U27015 ( .A(n25272), .B(n25271), .Z(n25273) );
  NANDN U27016 ( .A(n25274), .B(n25273), .Z(n25276) );
  NAND U27017 ( .A(n25276), .B(n25275), .Z(n25277) );
  NANDN U27018 ( .A(n25278), .B(n25277), .Z(n25280) );
  NAND U27019 ( .A(n25280), .B(n25279), .Z(n25281) );
  AND U27020 ( .A(n25282), .B(n25281), .Z(n25284) );
  NANDN U27021 ( .A(n25284), .B(n25283), .Z(n25286) );
  ANDN U27022 ( .B(n25286), .A(n25285), .Z(n25288) );
  NANDN U27023 ( .A(n25288), .B(n25287), .Z(n25289) );
  AND U27024 ( .A(n25290), .B(n25289), .Z(n25292) );
  NANDN U27025 ( .A(n25292), .B(n25291), .Z(n25294) );
  ANDN U27026 ( .B(n25294), .A(n25293), .Z(n25296) );
  NANDN U27027 ( .A(n25296), .B(n25295), .Z(n25297) );
  AND U27028 ( .A(n25298), .B(n25297), .Z(n25300) );
  NANDN U27029 ( .A(n25300), .B(n25299), .Z(n25302) );
  ANDN U27030 ( .B(n25302), .A(n25301), .Z(n25304) );
  NANDN U27031 ( .A(n25304), .B(n25303), .Z(n25305) );
  NANDN U27032 ( .A(n25306), .B(n25305), .Z(n25308) );
  NAND U27033 ( .A(n25308), .B(n25307), .Z(n25310) );
  NAND U27034 ( .A(n25310), .B(n25309), .Z(n25312) );
  NAND U27035 ( .A(n25312), .B(n25311), .Z(n25314) );
  ANDN U27036 ( .B(n25314), .A(n25313), .Z(n25316) );
  NANDN U27037 ( .A(n25316), .B(n25315), .Z(n25318) );
  NAND U27038 ( .A(n25318), .B(n25317), .Z(n25320) );
  NAND U27039 ( .A(n25320), .B(n25319), .Z(n25321) );
  AND U27040 ( .A(n25322), .B(n25321), .Z(n25324) );
  NANDN U27041 ( .A(n25324), .B(n25323), .Z(n25326) );
  NAND U27042 ( .A(n25326), .B(n25325), .Z(n25328) );
  NAND U27043 ( .A(n25328), .B(n25327), .Z(n25330) );
  ANDN U27044 ( .B(n25330), .A(n25329), .Z(n25332) );
  NANDN U27045 ( .A(n25332), .B(n25331), .Z(n25333) );
  NANDN U27046 ( .A(n25334), .B(n25333), .Z(n25336) );
  NAND U27047 ( .A(n25336), .B(n25335), .Z(n25337) );
  NANDN U27048 ( .A(n25338), .B(n25337), .Z(n25340) );
  NAND U27049 ( .A(n25340), .B(n25339), .Z(n25342) );
  NAND U27050 ( .A(n25342), .B(n25341), .Z(n25343) );
  AND U27051 ( .A(n25344), .B(n25343), .Z(n25348) );
  ANDN U27052 ( .B(n25346), .A(n25345), .Z(n25347) );
  NANDN U27053 ( .A(n25348), .B(n25347), .Z(n25349) );
  NANDN U27054 ( .A(n25350), .B(n25349), .Z(n25352) );
  NAND U27055 ( .A(n25352), .B(n25351), .Z(n25354) );
  ANDN U27056 ( .B(n25354), .A(n25353), .Z(n25355) );
  AND U27057 ( .A(n25356), .B(n25355), .Z(n25358) );
  NANDN U27058 ( .A(n25358), .B(n25357), .Z(n25359) );
  NANDN U27059 ( .A(n25360), .B(n25359), .Z(n25361) );
  NANDN U27060 ( .A(n25362), .B(n25361), .Z(n25364) );
  ANDN U27061 ( .B(n25364), .A(n25363), .Z(n25366) );
  NANDN U27062 ( .A(n25366), .B(n25365), .Z(n25368) );
  NAND U27063 ( .A(n25368), .B(n25367), .Z(n25370) );
  NAND U27064 ( .A(n25370), .B(n25369), .Z(n25371) );
  NANDN U27065 ( .A(n25372), .B(n25371), .Z(n25374) );
  ANDN U27066 ( .B(n25374), .A(n25373), .Z(n25376) );
  NANDN U27067 ( .A(n25376), .B(n25375), .Z(n25378) );
  NAND U27068 ( .A(n25378), .B(n25377), .Z(n25379) );
  AND U27069 ( .A(n25380), .B(n25379), .Z(n25382) );
  NANDN U27070 ( .A(n25382), .B(n25381), .Z(n25384) );
  NAND U27071 ( .A(n25384), .B(n25383), .Z(n25386) );
  NAND U27072 ( .A(n25386), .B(n25385), .Z(n25388) );
  NAND U27073 ( .A(n25388), .B(n25387), .Z(n25390) );
  ANDN U27074 ( .B(n25390), .A(n25389), .Z(n25392) );
  NANDN U27075 ( .A(n25392), .B(n25391), .Z(n25393) );
  NANDN U27076 ( .A(n25394), .B(n25393), .Z(n25396) );
  NAND U27077 ( .A(n25396), .B(n25395), .Z(n25398) );
  NAND U27078 ( .A(n25398), .B(n25397), .Z(n25400) );
  NAND U27079 ( .A(n25400), .B(n25399), .Z(n25401) );
  AND U27080 ( .A(n25402), .B(n25401), .Z(n25404) );
  NANDN U27081 ( .A(n25404), .B(n25403), .Z(n25405) );
  NANDN U27082 ( .A(n25406), .B(n25405), .Z(n25408) );
  NAND U27083 ( .A(n25408), .B(n25407), .Z(n25410) );
  ANDN U27084 ( .B(n25410), .A(n25409), .Z(n25412) );
  NANDN U27085 ( .A(n25412), .B(n25411), .Z(n25413) );
  NANDN U27086 ( .A(n25414), .B(n25413), .Z(n25416) );
  NAND U27087 ( .A(n25416), .B(n25415), .Z(n25417) );
  NANDN U27088 ( .A(n25418), .B(n25417), .Z(n25420) );
  NAND U27089 ( .A(n25420), .B(n25419), .Z(n25422) );
  ANDN U27090 ( .B(n25422), .A(n25421), .Z(n25424) );
  NANDN U27091 ( .A(n25424), .B(n25423), .Z(n25426) );
  ANDN U27092 ( .B(n25426), .A(n25425), .Z(n25428) );
  NANDN U27093 ( .A(n25428), .B(n25427), .Z(n25430) );
  ANDN U27094 ( .B(n25430), .A(n25429), .Z(n25432) );
  NANDN U27095 ( .A(n25432), .B(n25431), .Z(n25434) );
  ANDN U27096 ( .B(n25434), .A(n25433), .Z(n25436) );
  OR U27097 ( .A(n25436), .B(n25435), .Z(n25437) );
  AND U27098 ( .A(n25438), .B(n25437), .Z(n25440) );
  NANDN U27099 ( .A(n25440), .B(n25439), .Z(n25442) );
  ANDN U27100 ( .B(n25442), .A(n25441), .Z(n25444) );
  NANDN U27101 ( .A(n25444), .B(n25443), .Z(n25446) );
  NAND U27102 ( .A(n25446), .B(n25445), .Z(n25448) );
  ANDN U27103 ( .B(n25448), .A(n25447), .Z(n25450) );
  NANDN U27104 ( .A(n25450), .B(n25449), .Z(n25452) );
  ANDN U27105 ( .B(n25452), .A(n25451), .Z(n25453) );
  AND U27106 ( .A(n25454), .B(n25453), .Z(n25456) );
  OR U27107 ( .A(n25456), .B(n25455), .Z(n25457) );
  OR U27108 ( .A(n25457), .B(y[2621]), .Z(n25460) );
  XOR U27109 ( .A(n25457), .B(y[2621]), .Z(n25458) );
  NAND U27110 ( .A(n25458), .B(x[2621]), .Z(n25459) );
  NAND U27111 ( .A(n25460), .B(n25459), .Z(n25461) );
  AND U27112 ( .A(n25462), .B(n25461), .Z(n25463) );
  OR U27113 ( .A(n25464), .B(n25463), .Z(n25465) );
  AND U27114 ( .A(n25466), .B(n25465), .Z(n25468) );
  NANDN U27115 ( .A(n25468), .B(n25467), .Z(n25470) );
  ANDN U27116 ( .B(n25470), .A(n25469), .Z(n25471) );
  OR U27117 ( .A(n25472), .B(n25471), .Z(n25473) );
  NANDN U27118 ( .A(n25474), .B(n25473), .Z(n25476) );
  NAND U27119 ( .A(n25476), .B(n25475), .Z(n25477) );
  AND U27120 ( .A(n25478), .B(n25477), .Z(n25480) );
  NANDN U27121 ( .A(n25480), .B(n25479), .Z(n25482) );
  ANDN U27122 ( .B(n25482), .A(n25481), .Z(n25484) );
  NANDN U27123 ( .A(n25484), .B(n25483), .Z(n25485) );
  NANDN U27124 ( .A(n25486), .B(n25485), .Z(n25488) );
  NAND U27125 ( .A(n25488), .B(n25487), .Z(n25489) );
  AND U27126 ( .A(n25490), .B(n25489), .Z(n25492) );
  NANDN U27127 ( .A(n25492), .B(n25491), .Z(n25494) );
  NAND U27128 ( .A(n25494), .B(n25493), .Z(n25496) );
  NAND U27129 ( .A(n25496), .B(n25495), .Z(n25497) );
  AND U27130 ( .A(n25498), .B(n25497), .Z(n25499) );
  NAND U27131 ( .A(n25500), .B(n25499), .Z(n25502) );
  NAND U27132 ( .A(n25502), .B(n25501), .Z(n25504) );
  ANDN U27133 ( .B(n25504), .A(n25503), .Z(n25506) );
  OR U27134 ( .A(n25506), .B(n25505), .Z(n25508) );
  NAND U27135 ( .A(n25508), .B(n25507), .Z(n25509) );
  AND U27136 ( .A(n25510), .B(n25509), .Z(n25512) );
  NANDN U27137 ( .A(n25512), .B(n25511), .Z(n25513) );
  NANDN U27138 ( .A(n25514), .B(n25513), .Z(n25516) );
  NAND U27139 ( .A(n25516), .B(n25515), .Z(n25518) );
  NAND U27140 ( .A(n25518), .B(n25517), .Z(n25520) );
  NAND U27141 ( .A(n25520), .B(n25519), .Z(n25521) );
  AND U27142 ( .A(n25522), .B(n25521), .Z(n25524) );
  NANDN U27143 ( .A(n25524), .B(n25523), .Z(n25525) );
  AND U27144 ( .A(n25526), .B(n25525), .Z(n25527) );
  OR U27145 ( .A(n25528), .B(n25527), .Z(n25529) );
  NANDN U27146 ( .A(n25530), .B(n25529), .Z(n25532) );
  NAND U27147 ( .A(n25532), .B(n25531), .Z(n25533) );
  NANDN U27148 ( .A(n25534), .B(n25533), .Z(n25535) );
  NANDN U27149 ( .A(n25536), .B(n25535), .Z(n25538) );
  NAND U27150 ( .A(n25538), .B(n25537), .Z(n25539) );
  AND U27151 ( .A(n25540), .B(n25539), .Z(n25542) );
  NANDN U27152 ( .A(n25542), .B(n25541), .Z(n25543) );
  NANDN U27153 ( .A(n25544), .B(n25543), .Z(n25546) );
  NAND U27154 ( .A(n25546), .B(n25545), .Z(n25547) );
  AND U27155 ( .A(n25548), .B(n25547), .Z(n25550) );
  NANDN U27156 ( .A(n25550), .B(n25549), .Z(n25552) );
  NAND U27157 ( .A(n25552), .B(n25551), .Z(n25554) );
  NAND U27158 ( .A(n25554), .B(n25553), .Z(n25555) );
  AND U27159 ( .A(n25556), .B(n25555), .Z(n25558) );
  NANDN U27160 ( .A(n25558), .B(n25557), .Z(n25560) );
  NAND U27161 ( .A(n25560), .B(n25559), .Z(n25562) );
  NAND U27162 ( .A(n25562), .B(n25561), .Z(n25564) );
  ANDN U27163 ( .B(n25564), .A(n25563), .Z(n25566) );
  NANDN U27164 ( .A(n25566), .B(n25565), .Z(n25568) );
  NAND U27165 ( .A(n25568), .B(n25567), .Z(n25570) );
  NAND U27166 ( .A(n25570), .B(n25569), .Z(n25571) );
  AND U27167 ( .A(n25572), .B(n25571), .Z(n25574) );
  NANDN U27168 ( .A(n25574), .B(n25573), .Z(n25575) );
  NANDN U27169 ( .A(n25576), .B(n25575), .Z(n25578) );
  NAND U27170 ( .A(n25578), .B(n25577), .Z(n25580) );
  ANDN U27171 ( .B(n25580), .A(n25579), .Z(n25582) );
  OR U27172 ( .A(n25582), .B(n25581), .Z(n25584) );
  NAND U27173 ( .A(n25584), .B(n25583), .Z(n25586) );
  ANDN U27174 ( .B(n25586), .A(n25585), .Z(n25588) );
  NANDN U27175 ( .A(n25588), .B(n25587), .Z(n25590) );
  NAND U27176 ( .A(n25590), .B(n25589), .Z(n25592) );
  NAND U27177 ( .A(n25592), .B(n25591), .Z(n25593) );
  NANDN U27178 ( .A(n25594), .B(n25593), .Z(n25596) );
  ANDN U27179 ( .B(n25596), .A(n25595), .Z(n25598) );
  NANDN U27180 ( .A(n25598), .B(n25597), .Z(n25599) );
  AND U27181 ( .A(n25600), .B(n25599), .Z(n25602) );
  NANDN U27182 ( .A(n25602), .B(n25601), .Z(n25604) );
  ANDN U27183 ( .B(n25604), .A(n25603), .Z(n25605) );
  OR U27184 ( .A(n25606), .B(n25605), .Z(n25608) );
  NAND U27185 ( .A(n25608), .B(n25607), .Z(n25609) );
  NANDN U27186 ( .A(n25610), .B(n25609), .Z(n25611) );
  NANDN U27187 ( .A(n25611), .B(y[2686]), .Z(n25614) );
  XNOR U27188 ( .A(n25611), .B(y[2686]), .Z(n25612) );
  NANDN U27189 ( .A(x[2686]), .B(n25612), .Z(n25613) );
  NAND U27190 ( .A(n25614), .B(n25613), .Z(n25617) );
  NANDN U27191 ( .A(n25617), .B(n25618), .Z(n25615) );
  AND U27192 ( .A(n25616), .B(n25615), .Z(n25621) );
  XNOR U27193 ( .A(n25618), .B(n25617), .Z(n25619) );
  NAND U27194 ( .A(n25619), .B(x[2687]), .Z(n25620) );
  NAND U27195 ( .A(n25621), .B(n25620), .Z(n25622) );
  AND U27196 ( .A(n25623), .B(n25622), .Z(n25625) );
  NANDN U27197 ( .A(n25625), .B(n25624), .Z(n25627) );
  NAND U27198 ( .A(n25627), .B(n25626), .Z(n25629) );
  NAND U27199 ( .A(n25629), .B(n25628), .Z(n25631) );
  NAND U27200 ( .A(n25631), .B(n25630), .Z(n25633) );
  NAND U27201 ( .A(n25633), .B(n25632), .Z(n25639) );
  NANDN U27202 ( .A(n25635), .B(n25634), .Z(n25636) );
  AND U27203 ( .A(n25637), .B(n25636), .Z(n25638) );
  NAND U27204 ( .A(n25639), .B(n25638), .Z(n25641) );
  NAND U27205 ( .A(n25641), .B(n25640), .Z(n25642) );
  NANDN U27206 ( .A(n25643), .B(n25642), .Z(n25644) );
  NANDN U27207 ( .A(n25645), .B(n25644), .Z(n25646) );
  AND U27208 ( .A(n25647), .B(n25646), .Z(n25649) );
  NANDN U27209 ( .A(n25649), .B(n25648), .Z(n25651) );
  ANDN U27210 ( .B(n25651), .A(n25650), .Z(n25653) );
  NANDN U27211 ( .A(n25653), .B(n25652), .Z(n25655) );
  NAND U27212 ( .A(n25655), .B(n25654), .Z(n25657) );
  NAND U27213 ( .A(n25657), .B(n25656), .Z(n25659) );
  ANDN U27214 ( .B(n25659), .A(n25658), .Z(n25663) );
  ANDN U27215 ( .B(n25661), .A(n25660), .Z(n25662) );
  NANDN U27216 ( .A(n25663), .B(n25662), .Z(n25665) );
  NAND U27217 ( .A(n25665), .B(n25664), .Z(n25667) );
  ANDN U27218 ( .B(n25667), .A(n25666), .Z(n25669) );
  NANDN U27219 ( .A(n25669), .B(n25668), .Z(n25670) );
  NANDN U27220 ( .A(n25671), .B(n25670), .Z(n25673) );
  NAND U27221 ( .A(n25673), .B(n25672), .Z(n25675) );
  NANDN U27222 ( .A(n25675), .B(n25674), .Z(n25676) );
  NANDN U27223 ( .A(n25677), .B(n25676), .Z(n25679) );
  NAND U27224 ( .A(n25679), .B(n25678), .Z(n25680) );
  NANDN U27225 ( .A(n25681), .B(n25680), .Z(n25682) );
  NANDN U27226 ( .A(n25683), .B(n25682), .Z(n25684) );
  AND U27227 ( .A(n25685), .B(n25684), .Z(n25687) );
  NANDN U27228 ( .A(n25687), .B(n25686), .Z(n25688) );
  AND U27229 ( .A(n25689), .B(n25688), .Z(n25691) );
  NANDN U27230 ( .A(n25691), .B(n25690), .Z(n25693) );
  NAND U27231 ( .A(n25693), .B(n25692), .Z(n25695) );
  NAND U27232 ( .A(n25695), .B(n25694), .Z(n25696) );
  NANDN U27233 ( .A(n25697), .B(n25696), .Z(n25699) );
  ANDN U27234 ( .B(n25699), .A(n25698), .Z(n25700) );
  OR U27235 ( .A(n25701), .B(n25700), .Z(n25702) );
  NANDN U27236 ( .A(n25703), .B(n25702), .Z(n25704) );
  NANDN U27237 ( .A(n25705), .B(n25704), .Z(n25707) );
  NAND U27238 ( .A(n25707), .B(n25706), .Z(n25708) );
  AND U27239 ( .A(n25709), .B(n25708), .Z(n25711) );
  NANDN U27240 ( .A(n25711), .B(n25710), .Z(n25713) );
  ANDN U27241 ( .B(n25713), .A(n25712), .Z(n25715) );
  NANDN U27242 ( .A(n25715), .B(n25714), .Z(n25717) );
  ANDN U27243 ( .B(n25717), .A(n25716), .Z(n25719) );
  NANDN U27244 ( .A(n25719), .B(n25718), .Z(n25720) );
  AND U27245 ( .A(n25721), .B(n25720), .Z(n25723) );
  NANDN U27246 ( .A(n25723), .B(n25722), .Z(n25725) );
  ANDN U27247 ( .B(n25725), .A(n25724), .Z(n25727) );
  OR U27248 ( .A(n25727), .B(n25726), .Z(n25728) );
  AND U27249 ( .A(n25729), .B(n25728), .Z(n25731) );
  NANDN U27250 ( .A(n25731), .B(n25730), .Z(n25733) );
  ANDN U27251 ( .B(n25733), .A(n25732), .Z(n25734) );
  OR U27252 ( .A(n25735), .B(n25734), .Z(n25736) );
  NANDN U27253 ( .A(n25737), .B(n25736), .Z(n25739) );
  NAND U27254 ( .A(n25739), .B(n25738), .Z(n25740) );
  NANDN U27255 ( .A(n25741), .B(n25740), .Z(n25742) );
  NANDN U27256 ( .A(n25743), .B(n25742), .Z(n25745) );
  ANDN U27257 ( .B(n25745), .A(n25744), .Z(n25747) );
  NANDN U27258 ( .A(n25747), .B(n25746), .Z(n25749) );
  NAND U27259 ( .A(n25749), .B(n25748), .Z(n25751) );
  NAND U27260 ( .A(n25751), .B(n25750), .Z(n25752) );
  NANDN U27261 ( .A(n25753), .B(n25752), .Z(n25755) );
  NAND U27262 ( .A(n25755), .B(n25754), .Z(n25756) );
  AND U27263 ( .A(n25757), .B(n25756), .Z(n25759) );
  NANDN U27264 ( .A(n25759), .B(n25758), .Z(n25761) );
  NAND U27265 ( .A(n25761), .B(n25760), .Z(n25763) );
  NAND U27266 ( .A(n25763), .B(n25762), .Z(n25764) );
  NAND U27267 ( .A(n25765), .B(n25764), .Z(n25767) );
  NAND U27268 ( .A(n25767), .B(n25766), .Z(n25769) );
  ANDN U27269 ( .B(n25769), .A(n25768), .Z(n25770) );
  OR U27270 ( .A(n25771), .B(n25770), .Z(n25772) );
  NANDN U27271 ( .A(n25773), .B(n25772), .Z(n25774) );
  NANDN U27272 ( .A(n25775), .B(n25774), .Z(n25777) );
  NAND U27273 ( .A(n25777), .B(n25776), .Z(n25779) );
  NAND U27274 ( .A(n25779), .B(n25778), .Z(n25781) );
  NAND U27275 ( .A(n25781), .B(n25780), .Z(n25782) );
  AND U27276 ( .A(n25783), .B(n25782), .Z(n25785) );
  NANDN U27277 ( .A(n25785), .B(n25784), .Z(n25786) );
  NANDN U27278 ( .A(n25787), .B(n25786), .Z(n25788) );
  NANDN U27279 ( .A(n25789), .B(n25788), .Z(n25790) );
  AND U27280 ( .A(n25791), .B(n25790), .Z(n25793) );
  NANDN U27281 ( .A(n25793), .B(n25792), .Z(n25794) );
  NANDN U27282 ( .A(n25795), .B(n25794), .Z(n25797) );
  NAND U27283 ( .A(n25797), .B(n25796), .Z(n25799) );
  ANDN U27284 ( .B(n25799), .A(n25798), .Z(n25801) );
  NANDN U27285 ( .A(n25801), .B(n25800), .Z(n25802) );
  AND U27286 ( .A(n25803), .B(n25802), .Z(n25805) );
  NANDN U27287 ( .A(n25805), .B(n25804), .Z(n25806) );
  NANDN U27288 ( .A(n25807), .B(n25806), .Z(n25808) );
  AND U27289 ( .A(n25809), .B(n25808), .Z(n25811) );
  NANDN U27290 ( .A(n25811), .B(n25810), .Z(n25813) );
  ANDN U27291 ( .B(n25813), .A(n25812), .Z(n25814) );
  OR U27292 ( .A(n25815), .B(n25814), .Z(n25816) );
  NANDN U27293 ( .A(n25817), .B(n25816), .Z(n25818) );
  NANDN U27294 ( .A(n25819), .B(n25818), .Z(n25820) );
  AND U27295 ( .A(n25821), .B(n25820), .Z(n25823) );
  NANDN U27296 ( .A(n25823), .B(n25822), .Z(n25824) );
  NANDN U27297 ( .A(n25825), .B(n25824), .Z(n25826) );
  AND U27298 ( .A(n25827), .B(n25826), .Z(n25829) );
  NANDN U27299 ( .A(n25829), .B(n25828), .Z(n25830) );
  AND U27300 ( .A(n25831), .B(n25830), .Z(n25833) );
  NANDN U27301 ( .A(n25833), .B(n25832), .Z(n25834) );
  AND U27302 ( .A(n25835), .B(n25834), .Z(n25836) );
  ANDN U27303 ( .B(n25837), .A(n25836), .Z(n25839) );
  NAND U27304 ( .A(n25839), .B(n25838), .Z(n25840) );
  AND U27305 ( .A(n25841), .B(n25840), .Z(n25843) );
  NANDN U27306 ( .A(n25843), .B(n25842), .Z(n25845) );
  NAND U27307 ( .A(n25845), .B(n25844), .Z(n25847) );
  NAND U27308 ( .A(n25847), .B(n25846), .Z(n25848) );
  AND U27309 ( .A(n25849), .B(n25848), .Z(n25851) );
  NANDN U27310 ( .A(n25851), .B(n25850), .Z(n25853) );
  ANDN U27311 ( .B(n25853), .A(n25852), .Z(n25855) );
  NANDN U27312 ( .A(n25855), .B(n25854), .Z(n25857) );
  NAND U27313 ( .A(n25857), .B(n25856), .Z(n25858) );
  NANDN U27314 ( .A(n25859), .B(n25858), .Z(n25861) );
  NANDN U27315 ( .A(n25861), .B(y[2788]), .Z(n25864) );
  XOR U27316 ( .A(n25861), .B(n25860), .Z(n25862) );
  NANDN U27317 ( .A(x[2788]), .B(n25862), .Z(n25863) );
  NAND U27318 ( .A(n25864), .B(n25863), .Z(n25865) );
  NANDN U27319 ( .A(n25866), .B(n25865), .Z(n25867) );
  NANDN U27320 ( .A(n25868), .B(n25867), .Z(n25870) );
  NAND U27321 ( .A(n25870), .B(n25869), .Z(n25871) );
  NANDN U27322 ( .A(n25872), .B(n25871), .Z(n25874) );
  NAND U27323 ( .A(n25874), .B(n25873), .Z(n25875) );
  AND U27324 ( .A(n25876), .B(n25875), .Z(n25878) );
  NANDN U27325 ( .A(n25878), .B(n25877), .Z(n25880) );
  ANDN U27326 ( .B(n25880), .A(n25879), .Z(n25882) );
  OR U27327 ( .A(n25882), .B(n25881), .Z(n25883) );
  AND U27328 ( .A(n25884), .B(n25883), .Z(n25886) );
  NANDN U27329 ( .A(n25886), .B(n25885), .Z(n25888) );
  ANDN U27330 ( .B(n25888), .A(n25887), .Z(n25890) );
  OR U27331 ( .A(n25890), .B(n25889), .Z(n25891) );
  AND U27332 ( .A(n25892), .B(n25891), .Z(n25894) );
  NANDN U27333 ( .A(n25894), .B(n25893), .Z(n25895) );
  AND U27334 ( .A(n25896), .B(n25895), .Z(n25898) );
  NANDN U27335 ( .A(n25898), .B(n25897), .Z(n25899) );
  NANDN U27336 ( .A(n25900), .B(n25899), .Z(n25902) );
  NAND U27337 ( .A(n25902), .B(n25901), .Z(n25904) );
  NAND U27338 ( .A(n25904), .B(n25903), .Z(n25905) );
  NANDN U27339 ( .A(n25906), .B(n25905), .Z(n25907) );
  NANDN U27340 ( .A(n25908), .B(n25907), .Z(n25910) );
  ANDN U27341 ( .B(n25910), .A(n25909), .Z(n25912) );
  NANDN U27342 ( .A(n25912), .B(n25911), .Z(n25914) );
  NAND U27343 ( .A(n25914), .B(n25913), .Z(n25915) );
  AND U27344 ( .A(n25916), .B(n25915), .Z(n25918) );
  NANDN U27345 ( .A(n25918), .B(n25917), .Z(n25920) );
  ANDN U27346 ( .B(n25920), .A(n25919), .Z(n25922) );
  NANDN U27347 ( .A(n25922), .B(n25921), .Z(n25924) );
  NAND U27348 ( .A(n25924), .B(n25923), .Z(n25925) );
  NANDN U27349 ( .A(n25926), .B(n25925), .Z(n25927) );
  NANDN U27350 ( .A(n25927), .B(y[2815]), .Z(n25931) );
  XNOR U27351 ( .A(n25927), .B(y[2815]), .Z(n25928) );
  NAND U27352 ( .A(n25929), .B(n25928), .Z(n25930) );
  AND U27353 ( .A(n25931), .B(n25930), .Z(n25934) );
  OR U27354 ( .A(n25934), .B(x[2816]), .Z(n25932) );
  AND U27355 ( .A(n25933), .B(n25932), .Z(n25937) );
  XOR U27356 ( .A(n25934), .B(x[2816]), .Z(n25935) );
  NAND U27357 ( .A(n25935), .B(y[2816]), .Z(n25936) );
  NAND U27358 ( .A(n25937), .B(n25936), .Z(n25941) );
  NAND U27359 ( .A(n25939), .B(n25938), .Z(n25940) );
  AND U27360 ( .A(n25941), .B(n25940), .Z(n25942) );
  NANDN U27361 ( .A(n25943), .B(n25942), .Z(n25945) );
  ANDN U27362 ( .B(n25945), .A(n25944), .Z(n25947) );
  NANDN U27363 ( .A(n25947), .B(n25946), .Z(n25949) );
  NAND U27364 ( .A(n25949), .B(n25948), .Z(n25951) );
  NAND U27365 ( .A(n25951), .B(n25950), .Z(n25952) );
  AND U27366 ( .A(n25953), .B(n25952), .Z(n25955) );
  NANDN U27367 ( .A(n25955), .B(n25954), .Z(n25957) );
  ANDN U27368 ( .B(n25957), .A(n25956), .Z(n25959) );
  NANDN U27369 ( .A(n25959), .B(n25958), .Z(n25961) );
  NAND U27370 ( .A(n25961), .B(n25960), .Z(n25963) );
  NAND U27371 ( .A(n25963), .B(n25962), .Z(n25965) );
  NAND U27372 ( .A(n25965), .B(n25964), .Z(n25967) );
  NAND U27373 ( .A(n25967), .B(n25966), .Z(n25969) );
  ANDN U27374 ( .B(n25969), .A(n25968), .Z(n25971) );
  NAND U27375 ( .A(n25971), .B(n25970), .Z(n25972) );
  AND U27376 ( .A(n25973), .B(n25972), .Z(n25975) );
  NAND U27377 ( .A(n25975), .B(n25974), .Z(n25976) );
  AND U27378 ( .A(n25977), .B(n25976), .Z(n25978) );
  NANDN U27379 ( .A(n25979), .B(n25978), .Z(n25981) );
  NAND U27380 ( .A(n25981), .B(n25980), .Z(n25985) );
  NAND U27381 ( .A(n25983), .B(n25982), .Z(n25984) );
  NANDN U27382 ( .A(n25985), .B(n25984), .Z(n25986) );
  AND U27383 ( .A(n25987), .B(n25986), .Z(n25989) );
  NANDN U27384 ( .A(n25989), .B(n25988), .Z(n25991) );
  ANDN U27385 ( .B(n25991), .A(n25990), .Z(n25993) );
  NANDN U27386 ( .A(n25993), .B(n25992), .Z(n25995) );
  ANDN U27387 ( .B(n25995), .A(n25994), .Z(n25997) );
  NANDN U27388 ( .A(n25997), .B(n25996), .Z(n25998) );
  AND U27389 ( .A(n25999), .B(n25998), .Z(n26001) );
  NANDN U27390 ( .A(n26001), .B(n26000), .Z(n26003) );
  ANDN U27391 ( .B(n26003), .A(n26002), .Z(n26005) );
  NANDN U27392 ( .A(n26005), .B(n26004), .Z(n26006) );
  AND U27393 ( .A(n26007), .B(n26006), .Z(n26009) );
  NANDN U27394 ( .A(n26009), .B(n26008), .Z(n26011) );
  ANDN U27395 ( .B(n26011), .A(n26010), .Z(n26013) );
  NANDN U27396 ( .A(n26013), .B(n26012), .Z(n26015) );
  ANDN U27397 ( .B(n26015), .A(n26014), .Z(n26017) );
  NANDN U27398 ( .A(n26017), .B(n26016), .Z(n26018) );
  AND U27399 ( .A(n26019), .B(n26018), .Z(n26021) );
  NANDN U27400 ( .A(n26021), .B(n26020), .Z(n26022) );
  NANDN U27401 ( .A(n26023), .B(n26022), .Z(n26024) );
  AND U27402 ( .A(n26025), .B(n26024), .Z(n26027) );
  NANDN U27403 ( .A(n26027), .B(n26026), .Z(n26029) );
  ANDN U27404 ( .B(n26029), .A(n26028), .Z(n26030) );
  OR U27405 ( .A(n26031), .B(n26030), .Z(n26032) );
  NANDN U27406 ( .A(n26033), .B(n26032), .Z(n26035) );
  NAND U27407 ( .A(n26035), .B(n26034), .Z(n26037) );
  NAND U27408 ( .A(n26037), .B(n26036), .Z(n26039) );
  NAND U27409 ( .A(n26039), .B(n26038), .Z(n26041) );
  ANDN U27410 ( .B(n26041), .A(n26040), .Z(n26043) );
  NANDN U27411 ( .A(n26043), .B(n26042), .Z(n26045) );
  NAND U27412 ( .A(n26045), .B(n26044), .Z(n26047) );
  NAND U27413 ( .A(n26047), .B(n26046), .Z(n26049) );
  ANDN U27414 ( .B(n26049), .A(n26048), .Z(n26051) );
  NAND U27415 ( .A(n26051), .B(n26050), .Z(n26053) );
  NAND U27416 ( .A(n26053), .B(n26052), .Z(n26055) );
  ANDN U27417 ( .B(n26055), .A(n26054), .Z(n26057) );
  NANDN U27418 ( .A(n26057), .B(n26056), .Z(n26059) );
  NAND U27419 ( .A(n26059), .B(n26058), .Z(n26061) );
  NAND U27420 ( .A(n26061), .B(n26060), .Z(n26062) );
  AND U27421 ( .A(n26063), .B(n26062), .Z(n26065) );
  NANDN U27422 ( .A(n26065), .B(n26064), .Z(n26067) );
  NAND U27423 ( .A(n26067), .B(n26066), .Z(n26069) );
  NAND U27424 ( .A(n26069), .B(n26068), .Z(n26070) );
  NANDN U27425 ( .A(n26071), .B(n26070), .Z(n26073) );
  NAND U27426 ( .A(n26073), .B(n26072), .Z(n26075) );
  ANDN U27427 ( .B(n26075), .A(n26074), .Z(n26076) );
  NAND U27428 ( .A(n26077), .B(n26076), .Z(n26078) );
  NAND U27429 ( .A(n26079), .B(n26078), .Z(n26081) );
  ANDN U27430 ( .B(n26081), .A(n26080), .Z(n26083) );
  OR U27431 ( .A(n26083), .B(n26082), .Z(n26084) );
  NANDN U27432 ( .A(n26085), .B(n26084), .Z(n26087) );
  NAND U27433 ( .A(n26087), .B(n26086), .Z(n26089) );
  NAND U27434 ( .A(n26089), .B(n26088), .Z(n26090) );
  NANDN U27435 ( .A(n26091), .B(n26090), .Z(n26092) );
  NANDN U27436 ( .A(n26093), .B(n26092), .Z(n26095) );
  ANDN U27437 ( .B(n26095), .A(n26094), .Z(n26097) );
  NANDN U27438 ( .A(n26097), .B(n26096), .Z(n26099) );
  NAND U27439 ( .A(n26099), .B(n26098), .Z(n26101) );
  NAND U27440 ( .A(n26101), .B(n26100), .Z(n26102) );
  AND U27441 ( .A(n26103), .B(n26102), .Z(n26105) );
  NANDN U27442 ( .A(n26105), .B(n26104), .Z(n26106) );
  NANDN U27443 ( .A(n26107), .B(n26106), .Z(n26109) );
  NAND U27444 ( .A(n26109), .B(n26108), .Z(n26111) );
  ANDN U27445 ( .B(n26111), .A(n26110), .Z(n26113) );
  OR U27446 ( .A(n26113), .B(n26112), .Z(n26115) );
  NAND U27447 ( .A(n26115), .B(n26114), .Z(n26117) );
  ANDN U27448 ( .B(n26117), .A(n26116), .Z(n26119) );
  NANDN U27449 ( .A(n26119), .B(n26118), .Z(n26121) );
  NAND U27450 ( .A(n26121), .B(n26120), .Z(n26123) );
  NAND U27451 ( .A(n26123), .B(n26122), .Z(n26125) );
  NAND U27452 ( .A(n26125), .B(n26124), .Z(n26127) );
  ANDN U27453 ( .B(n26127), .A(n26126), .Z(n26129) );
  NANDN U27454 ( .A(n26129), .B(n26128), .Z(n26130) );
  AND U27455 ( .A(n26131), .B(n26130), .Z(n26133) );
  NANDN U27456 ( .A(n26133), .B(n26132), .Z(n26135) );
  ANDN U27457 ( .B(n26135), .A(n26134), .Z(n26137) );
  NANDN U27458 ( .A(n26137), .B(n26136), .Z(n26138) );
  AND U27459 ( .A(n26139), .B(n26138), .Z(n26141) );
  NANDN U27460 ( .A(n26141), .B(n26140), .Z(n26143) );
  ANDN U27461 ( .B(n26143), .A(n26142), .Z(n26145) );
  OR U27462 ( .A(n26145), .B(n26144), .Z(n26146) );
  AND U27463 ( .A(n26147), .B(n26146), .Z(n26149) );
  NANDN U27464 ( .A(n26149), .B(n26148), .Z(n26151) );
  ANDN U27465 ( .B(n26151), .A(n26150), .Z(n26153) );
  NANDN U27466 ( .A(n26153), .B(n26152), .Z(n26155) );
  NAND U27467 ( .A(n26155), .B(n26154), .Z(n26157) );
  NAND U27468 ( .A(n26157), .B(n26156), .Z(n26159) );
  NAND U27469 ( .A(n26159), .B(n26158), .Z(n26161) );
  NAND U27470 ( .A(n26161), .B(n26160), .Z(n26163) );
  ANDN U27471 ( .B(n26163), .A(n26162), .Z(n26165) );
  NANDN U27472 ( .A(n26165), .B(n26164), .Z(n26166) );
  NANDN U27473 ( .A(n26167), .B(n26166), .Z(n26169) );
  NAND U27474 ( .A(n26169), .B(n26168), .Z(n26171) );
  NAND U27475 ( .A(n26171), .B(n26170), .Z(n26173) );
  NAND U27476 ( .A(n26173), .B(n26172), .Z(n26174) );
  AND U27477 ( .A(n26175), .B(n26174), .Z(n26177) );
  NANDN U27478 ( .A(n26177), .B(n26176), .Z(n26179) );
  ANDN U27479 ( .B(n26179), .A(n26178), .Z(n26181) );
  NANDN U27480 ( .A(n26181), .B(n26180), .Z(n26183) );
  AND U27481 ( .A(n26183), .B(n26182), .Z(n26187) );
  ANDN U27482 ( .B(n26185), .A(n26184), .Z(n26186) );
  NANDN U27483 ( .A(n26187), .B(n26186), .Z(n26188) );
  NANDN U27484 ( .A(n26189), .B(n26188), .Z(n26191) );
  NAND U27485 ( .A(n26191), .B(n26190), .Z(n26192) );
  AND U27486 ( .A(n26193), .B(n26192), .Z(n26195) );
  NANDN U27487 ( .A(n26195), .B(n26194), .Z(n26196) );
  NANDN U27488 ( .A(n26197), .B(n26196), .Z(n26199) );
  NAND U27489 ( .A(n26199), .B(n26198), .Z(n26200) );
  NANDN U27490 ( .A(n26201), .B(n26200), .Z(n26202) );
  NANDN U27491 ( .A(n26203), .B(n26202), .Z(n26205) );
  ANDN U27492 ( .B(n26205), .A(n26204), .Z(n26207) );
  NANDN U27493 ( .A(n26207), .B(n26206), .Z(n26208) );
  AND U27494 ( .A(n26209), .B(n26208), .Z(n26211) );
  NANDN U27495 ( .A(n26211), .B(n26210), .Z(n26213) );
  ANDN U27496 ( .B(n26213), .A(n26212), .Z(n26215) );
  OR U27497 ( .A(n26215), .B(n26214), .Z(n26216) );
  AND U27498 ( .A(n26217), .B(n26216), .Z(n26219) );
  NANDN U27499 ( .A(n26219), .B(n26218), .Z(n26221) );
  ANDN U27500 ( .B(n26221), .A(n26220), .Z(n26223) );
  NANDN U27501 ( .A(n26223), .B(n26222), .Z(n26224) );
  NANDN U27502 ( .A(n26225), .B(n26224), .Z(n26227) );
  NAND U27503 ( .A(n26227), .B(n26226), .Z(n26229) );
  NAND U27504 ( .A(n26229), .B(n26228), .Z(n26231) );
  NAND U27505 ( .A(n26231), .B(n26230), .Z(n26233) );
  ANDN U27506 ( .B(n26233), .A(n26232), .Z(n26235) );
  NANDN U27507 ( .A(n26235), .B(n26234), .Z(n26237) );
  NAND U27508 ( .A(n26237), .B(n26236), .Z(n26239) );
  NAND U27509 ( .A(n26239), .B(n26238), .Z(n26241) );
  ANDN U27510 ( .B(n26241), .A(n26240), .Z(n26242) );
  OR U27511 ( .A(n26243), .B(n26242), .Z(n26245) );
  NAND U27512 ( .A(n26245), .B(n26244), .Z(n26246) );
  AND U27513 ( .A(n26247), .B(n26246), .Z(n26249) );
  NANDN U27514 ( .A(n26249), .B(n26248), .Z(n26250) );
  NANDN U27515 ( .A(n26251), .B(n26250), .Z(n26253) );
  NAND U27516 ( .A(n26253), .B(n26252), .Z(n26255) );
  NAND U27517 ( .A(n26255), .B(n26254), .Z(n26257) );
  NAND U27518 ( .A(n26257), .B(n26256), .Z(n26259) );
  ANDN U27519 ( .B(n26259), .A(n26258), .Z(n26261) );
  NANDN U27520 ( .A(n26261), .B(n26260), .Z(n26263) );
  ANDN U27521 ( .B(n26263), .A(n26262), .Z(n26265) );
  NANDN U27522 ( .A(n26265), .B(n26264), .Z(n26267) );
  ANDN U27523 ( .B(n26267), .A(n26266), .Z(n26269) );
  NANDN U27524 ( .A(n26269), .B(n26268), .Z(n26271) );
  NAND U27525 ( .A(n26271), .B(n26270), .Z(n26272) );
  NANDN U27526 ( .A(n26273), .B(n26272), .Z(n26275) );
  NAND U27527 ( .A(n26275), .B(n26274), .Z(n26276) );
  AND U27528 ( .A(n26277), .B(n26276), .Z(n26279) );
  NANDN U27529 ( .A(n26279), .B(n26278), .Z(n26281) );
  ANDN U27530 ( .B(n26281), .A(n26280), .Z(n26283) );
  OR U27531 ( .A(n26283), .B(n26282), .Z(n26284) );
  AND U27532 ( .A(n26285), .B(n26284), .Z(n26287) );
  NANDN U27533 ( .A(n26287), .B(n26286), .Z(n26289) );
  ANDN U27534 ( .B(n26289), .A(n26288), .Z(n26291) );
  NANDN U27535 ( .A(n26291), .B(n26290), .Z(n26292) );
  NANDN U27536 ( .A(n26293), .B(n26292), .Z(n26295) );
  NAND U27537 ( .A(n26295), .B(n26294), .Z(n26297) );
  NAND U27538 ( .A(n26297), .B(n26296), .Z(n26298) );
  NANDN U27539 ( .A(n26299), .B(n26298), .Z(n26300) );
  NANDN U27540 ( .A(n26301), .B(n26300), .Z(n26302) );
  AND U27541 ( .A(n26303), .B(n26302), .Z(n26305) );
  NANDN U27542 ( .A(n26305), .B(n26304), .Z(n26307) );
  NAND U27543 ( .A(n26307), .B(n26306), .Z(n26309) );
  NAND U27544 ( .A(n26309), .B(n26308), .Z(n26311) );
  ANDN U27545 ( .B(n26311), .A(n26310), .Z(n26313) );
  NANDN U27546 ( .A(n26313), .B(n26312), .Z(n26315) );
  NAND U27547 ( .A(n26315), .B(n26314), .Z(n26317) );
  NAND U27548 ( .A(n26317), .B(n26316), .Z(n26318) );
  AND U27549 ( .A(n26319), .B(n26318), .Z(n26321) );
  NANDN U27550 ( .A(n26321), .B(n26320), .Z(n26323) );
  NAND U27551 ( .A(n26323), .B(n26322), .Z(n26325) );
  NAND U27552 ( .A(n26325), .B(n26324), .Z(n26327) );
  ANDN U27553 ( .B(n26327), .A(n26326), .Z(n26328) );
  OR U27554 ( .A(n26329), .B(n26328), .Z(n26331) );
  NAND U27555 ( .A(n26331), .B(n26330), .Z(n26333) );
  NAND U27556 ( .A(n26333), .B(n26332), .Z(n26335) );
  ANDN U27557 ( .B(n26335), .A(n26334), .Z(n26337) );
  NANDN U27558 ( .A(n26337), .B(n26336), .Z(n26339) );
  NAND U27559 ( .A(n26339), .B(n26338), .Z(n26340) );
  AND U27560 ( .A(n26341), .B(n26340), .Z(n26343) );
  NANDN U27561 ( .A(n26343), .B(n26342), .Z(n26344) );
  NANDN U27562 ( .A(n26345), .B(n26344), .Z(n26346) );
  NANDN U27563 ( .A(n26347), .B(n26346), .Z(n26349) );
  NAND U27564 ( .A(n26349), .B(n26348), .Z(n26351) );
  NAND U27565 ( .A(n26351), .B(n26350), .Z(n26353) );
  NAND U27566 ( .A(n26353), .B(n26352), .Z(n26354) );
  AND U27567 ( .A(n26355), .B(n26354), .Z(n26357) );
  NANDN U27568 ( .A(n26357), .B(n26356), .Z(n26359) );
  NAND U27569 ( .A(n26359), .B(n26358), .Z(n26361) );
  NAND U27570 ( .A(n26361), .B(n26360), .Z(n26363) );
  ANDN U27571 ( .B(n26363), .A(n26362), .Z(n26364) );
  OR U27572 ( .A(n26365), .B(n26364), .Z(n26367) );
  NAND U27573 ( .A(n26367), .B(n26366), .Z(n26369) );
  NAND U27574 ( .A(n26369), .B(n26368), .Z(n26371) );
  ANDN U27575 ( .B(n26371), .A(n26370), .Z(n26373) );
  NANDN U27576 ( .A(n26373), .B(n26372), .Z(n26375) );
  NAND U27577 ( .A(n26375), .B(n26374), .Z(n26376) );
  AND U27578 ( .A(n26377), .B(n26376), .Z(n26379) );
  NANDN U27579 ( .A(n26379), .B(n26378), .Z(n26380) );
  NANDN U27580 ( .A(n26381), .B(n26380), .Z(n26382) );
  NANDN U27581 ( .A(n26383), .B(n26382), .Z(n26385) );
  NAND U27582 ( .A(n26385), .B(n26384), .Z(n26387) );
  NAND U27583 ( .A(n26387), .B(n26386), .Z(n26389) );
  NAND U27584 ( .A(n26389), .B(n26388), .Z(n26390) );
  AND U27585 ( .A(n26391), .B(n26390), .Z(n26393) );
  NANDN U27586 ( .A(n26393), .B(n26392), .Z(n26395) );
  NAND U27587 ( .A(n26395), .B(n26394), .Z(n26397) );
  NAND U27588 ( .A(n26397), .B(n26396), .Z(n26399) );
  ANDN U27589 ( .B(n26399), .A(n26398), .Z(n26400) );
  OR U27590 ( .A(n26401), .B(n26400), .Z(n26403) );
  NAND U27591 ( .A(n26403), .B(n26402), .Z(n26405) );
  NAND U27592 ( .A(n26405), .B(n26404), .Z(n26407) );
  ANDN U27593 ( .B(n26407), .A(n26406), .Z(n26409) );
  NANDN U27594 ( .A(n26409), .B(n26408), .Z(n26411) );
  NAND U27595 ( .A(n26411), .B(n26410), .Z(n26412) );
  AND U27596 ( .A(n26413), .B(n26412), .Z(n26415) );
  NANDN U27597 ( .A(n26415), .B(n26414), .Z(n26416) );
  NANDN U27598 ( .A(n26417), .B(n26416), .Z(n26418) );
  NANDN U27599 ( .A(n26419), .B(n26418), .Z(n26421) );
  NAND U27600 ( .A(n26421), .B(n26420), .Z(n26423) );
  NAND U27601 ( .A(n26423), .B(n26422), .Z(n26425) );
  NAND U27602 ( .A(n26425), .B(n26424), .Z(n26426) );
  AND U27603 ( .A(n26427), .B(n26426), .Z(n26429) );
  NANDN U27604 ( .A(n26429), .B(n26428), .Z(n26431) );
  NAND U27605 ( .A(n26431), .B(n26430), .Z(n26433) );
  NAND U27606 ( .A(n26433), .B(n26432), .Z(n26435) );
  ANDN U27607 ( .B(n26435), .A(n26434), .Z(n26436) );
  OR U27608 ( .A(n26437), .B(n26436), .Z(n26439) );
  NAND U27609 ( .A(n26439), .B(n26438), .Z(n26441) );
  NAND U27610 ( .A(n26441), .B(n26440), .Z(n26443) );
  ANDN U27611 ( .B(n26443), .A(n26442), .Z(n26445) );
  NANDN U27612 ( .A(n26445), .B(n26444), .Z(n26447) );
  NAND U27613 ( .A(n26447), .B(n26446), .Z(n26448) );
  AND U27614 ( .A(n26449), .B(n26448), .Z(n26451) );
  NANDN U27615 ( .A(n26451), .B(n26450), .Z(n26452) );
  NANDN U27616 ( .A(n26453), .B(n26452), .Z(n26455) );
  NAND U27617 ( .A(n26455), .B(n26454), .Z(n26457) );
  NAND U27618 ( .A(n26457), .B(n26456), .Z(n26459) );
  NAND U27619 ( .A(n26459), .B(n26458), .Z(n26460) );
  NANDN U27620 ( .A(n26461), .B(n26460), .Z(n26463) );
  ANDN U27621 ( .B(n26463), .A(n26462), .Z(n26465) );
  NANDN U27622 ( .A(n26465), .B(n26464), .Z(n26467) );
  NAND U27623 ( .A(n26467), .B(n26466), .Z(n26469) );
  NAND U27624 ( .A(n26469), .B(n26468), .Z(n26471) );
  ANDN U27625 ( .B(n26471), .A(n26470), .Z(n26473) );
  NANDN U27626 ( .A(n26473), .B(n26472), .Z(n26475) );
  NAND U27627 ( .A(n26475), .B(n26474), .Z(n26477) );
  NAND U27628 ( .A(n26477), .B(n26476), .Z(n26479) );
  ANDN U27629 ( .B(n26479), .A(n26478), .Z(n26481) );
  NANDN U27630 ( .A(n26481), .B(n26480), .Z(n26483) );
  NAND U27631 ( .A(n26483), .B(n26482), .Z(n26484) );
  AND U27632 ( .A(n26485), .B(n26484), .Z(n26487) );
  NANDN U27633 ( .A(n26487), .B(n26486), .Z(n26488) );
  NANDN U27634 ( .A(n26489), .B(n26488), .Z(n26490) );
  NANDN U27635 ( .A(n26491), .B(n26490), .Z(n26493) );
  NAND U27636 ( .A(n26493), .B(n26492), .Z(n26495) );
  NAND U27637 ( .A(n26495), .B(n26494), .Z(n26497) );
  NAND U27638 ( .A(n26497), .B(n26496), .Z(n26498) );
  AND U27639 ( .A(n26499), .B(n26498), .Z(n26501) );
  NANDN U27640 ( .A(n26501), .B(n26500), .Z(n26502) );
  NANDN U27641 ( .A(n26503), .B(n26502), .Z(n26504) );
  NANDN U27642 ( .A(n26505), .B(n26504), .Z(n26507) );
  ANDN U27643 ( .B(n26507), .A(n26506), .Z(n26508) );
  OR U27644 ( .A(n26509), .B(n26508), .Z(n26511) );
  NAND U27645 ( .A(n26511), .B(n26510), .Z(n26513) );
  NAND U27646 ( .A(n26513), .B(n26512), .Z(n26515) );
  ANDN U27647 ( .B(n26515), .A(n26514), .Z(n26517) );
  NANDN U27648 ( .A(n26517), .B(n26516), .Z(n26519) );
  NAND U27649 ( .A(n26519), .B(n26518), .Z(n26520) );
  AND U27650 ( .A(n26521), .B(n26520), .Z(n26523) );
  NANDN U27651 ( .A(n26523), .B(n26522), .Z(n26524) );
  NANDN U27652 ( .A(n26525), .B(n26524), .Z(n26526) );
  NANDN U27653 ( .A(n26527), .B(n26526), .Z(n26529) );
  NAND U27654 ( .A(n26529), .B(n26528), .Z(n26531) );
  NAND U27655 ( .A(n26531), .B(n26530), .Z(n26533) );
  NAND U27656 ( .A(n26533), .B(n26532), .Z(n26534) );
  AND U27657 ( .A(n26535), .B(n26534), .Z(n26537) );
  NANDN U27658 ( .A(n26537), .B(n26536), .Z(n26539) );
  NAND U27659 ( .A(n26539), .B(n26538), .Z(n26541) );
  NAND U27660 ( .A(n26541), .B(n26540), .Z(n26542) );
  AND U27661 ( .A(n26543), .B(n26542), .Z(n26544) );
  NANDN U27662 ( .A(n26545), .B(n26544), .Z(n26547) );
  NAND U27663 ( .A(n26547), .B(n26546), .Z(n26548) );
  AND U27664 ( .A(n26549), .B(n26548), .Z(n26551) );
  NANDN U27665 ( .A(n26551), .B(n26550), .Z(n26553) );
  ANDN U27666 ( .B(n26553), .A(n26552), .Z(n26555) );
  OR U27667 ( .A(n26555), .B(n26554), .Z(n26556) );
  AND U27668 ( .A(n26557), .B(n26556), .Z(n26559) );
  NANDN U27669 ( .A(n26559), .B(n26558), .Z(n26560) );
  AND U27670 ( .A(n26561), .B(n26560), .Z(n26563) );
  NANDN U27671 ( .A(n26563), .B(n26562), .Z(n26564) );
  NANDN U27672 ( .A(n26565), .B(n26564), .Z(n26567) );
  NAND U27673 ( .A(n26567), .B(n26566), .Z(n26569) );
  NAND U27674 ( .A(n26569), .B(n26568), .Z(n26570) );
  NANDN U27675 ( .A(n26571), .B(n26570), .Z(n26572) );
  NANDN U27676 ( .A(n26573), .B(n26572), .Z(n26574) );
  AND U27677 ( .A(n26575), .B(n26574), .Z(n26577) );
  NANDN U27678 ( .A(n26577), .B(n26576), .Z(n26579) );
  NAND U27679 ( .A(n26579), .B(n26578), .Z(n26581) );
  NAND U27680 ( .A(n26581), .B(n26580), .Z(n26584) );
  NANDN U27681 ( .A(y[3068]), .B(n26584), .Z(n26582) );
  AND U27682 ( .A(n26583), .B(n26582), .Z(n26587) );
  XNOR U27683 ( .A(n26584), .B(y[3068]), .Z(n26585) );
  NAND U27684 ( .A(n26585), .B(x[3068]), .Z(n26586) );
  NAND U27685 ( .A(n26587), .B(n26586), .Z(n26589) );
  ANDN U27686 ( .B(n26589), .A(n26588), .Z(n26591) );
  NANDN U27687 ( .A(n26591), .B(n26590), .Z(n26592) );
  NANDN U27688 ( .A(n26593), .B(n26592), .Z(n26595) );
  ANDN U27689 ( .B(n26595), .A(n26594), .Z(n26596) );
  OR U27690 ( .A(n26597), .B(n26596), .Z(n26598) );
  NANDN U27691 ( .A(n26599), .B(n26598), .Z(n26600) );
  NANDN U27692 ( .A(n26601), .B(n26600), .Z(n26603) );
  NAND U27693 ( .A(n26603), .B(n26602), .Z(n26605) );
  ANDN U27694 ( .B(n26605), .A(n26604), .Z(n26607) );
  NANDN U27695 ( .A(n26607), .B(n26606), .Z(n26608) );
  NANDN U27696 ( .A(n26609), .B(n26608), .Z(n26610) );
  NANDN U27697 ( .A(n26611), .B(n26610), .Z(n26613) );
  NAND U27698 ( .A(n26613), .B(n26612), .Z(n26615) );
  ANDN U27699 ( .B(n26615), .A(n26614), .Z(n26616) );
  OR U27700 ( .A(n26617), .B(n26616), .Z(n26618) );
  NANDN U27701 ( .A(n26619), .B(n26618), .Z(n26620) );
  NANDN U27702 ( .A(n26621), .B(n26620), .Z(n26623) );
  NAND U27703 ( .A(n26623), .B(n26622), .Z(n26625) );
  ANDN U27704 ( .B(n26625), .A(n26624), .Z(n26626) );
  OR U27705 ( .A(n26627), .B(n26626), .Z(n26628) );
  NANDN U27706 ( .A(n26629), .B(n26628), .Z(n26631) );
  NAND U27707 ( .A(n26631), .B(n26630), .Z(n26633) );
  ANDN U27708 ( .B(n26633), .A(n26632), .Z(n26635) );
  NAND U27709 ( .A(n26635), .B(n26634), .Z(n26637) );
  NAND U27710 ( .A(n26637), .B(n26636), .Z(n26638) );
  AND U27711 ( .A(n26639), .B(n26638), .Z(n26641) );
  NAND U27712 ( .A(n26641), .B(n26640), .Z(n26642) );
  NANDN U27713 ( .A(n26643), .B(n26642), .Z(n26645) );
  ANDN U27714 ( .B(n26645), .A(n26644), .Z(n26647) );
  NANDN U27715 ( .A(n26647), .B(n26646), .Z(n26648) );
  NANDN U27716 ( .A(n26649), .B(n26648), .Z(n26651) );
  NAND U27717 ( .A(n26651), .B(n26650), .Z(n26652) );
  NANDN U27718 ( .A(n26653), .B(n26652), .Z(n26655) );
  ANDN U27719 ( .B(n26655), .A(n26654), .Z(n26657) );
  NANDN U27720 ( .A(n26657), .B(n26656), .Z(n26658) );
  NANDN U27721 ( .A(n26659), .B(n26658), .Z(n26661) );
  NAND U27722 ( .A(n26661), .B(n26660), .Z(n26662) );
  NANDN U27723 ( .A(n26663), .B(n26662), .Z(n26665) );
  ANDN U27724 ( .B(n26665), .A(n26664), .Z(n26666) );
  OR U27725 ( .A(n26667), .B(n26666), .Z(n26668) );
  NANDN U27726 ( .A(n26669), .B(n26668), .Z(n26671) );
  NAND U27727 ( .A(n26671), .B(n26670), .Z(n26673) );
  NAND U27728 ( .A(n26673), .B(n26672), .Z(n26675) );
  ANDN U27729 ( .B(n26675), .A(n26674), .Z(n26676) );
  OR U27730 ( .A(n26677), .B(n26676), .Z(n26678) );
  NANDN U27731 ( .A(n26679), .B(n26678), .Z(n26681) );
  NAND U27732 ( .A(n26681), .B(n26680), .Z(n26682) );
  NANDN U27733 ( .A(n26683), .B(n26682), .Z(n26685) );
  ANDN U27734 ( .B(n26685), .A(n26684), .Z(n26686) );
  OR U27735 ( .A(n26687), .B(n26686), .Z(n26689) );
  NAND U27736 ( .A(n26689), .B(n26688), .Z(n26691) );
  NAND U27737 ( .A(n26691), .B(n26690), .Z(n26692) );
  NANDN U27738 ( .A(n26693), .B(n26692), .Z(n26695) );
  ANDN U27739 ( .B(n26695), .A(n26694), .Z(n26697) );
  NANDN U27740 ( .A(n26697), .B(n26696), .Z(n26698) );
  NANDN U27741 ( .A(n26699), .B(n26698), .Z(n26701) );
  NAND U27742 ( .A(n26701), .B(n26700), .Z(n26702) );
  NANDN U27743 ( .A(n26703), .B(n26702), .Z(n26705) );
  ANDN U27744 ( .B(n26705), .A(n26704), .Z(n26706) );
  OR U27745 ( .A(n26707), .B(n26706), .Z(n26708) );
  NANDN U27746 ( .A(n26709), .B(n26708), .Z(n26711) );
  NAND U27747 ( .A(n26711), .B(n26710), .Z(n26712) );
  NANDN U27748 ( .A(n26713), .B(n26712), .Z(n26715) );
  NAND U27749 ( .A(n26715), .B(n26714), .Z(n26717) );
  ANDN U27750 ( .B(n26717), .A(n26716), .Z(n26719) );
  NANDN U27751 ( .A(n26719), .B(n26718), .Z(n26721) );
  ANDN U27752 ( .B(n26721), .A(n26720), .Z(n26723) );
  NANDN U27753 ( .A(n26723), .B(n26722), .Z(n26725) );
  ANDN U27754 ( .B(n26725), .A(n26724), .Z(n26727) );
  NANDN U27755 ( .A(n26727), .B(n26726), .Z(n26729) );
  ANDN U27756 ( .B(n26729), .A(n26728), .Z(n26731) );
  NANDN U27757 ( .A(n26731), .B(n26730), .Z(n26733) );
  NAND U27758 ( .A(n26733), .B(n26732), .Z(n26734) );
  NANDN U27759 ( .A(n26735), .B(n26734), .Z(n26737) );
  NAND U27760 ( .A(n26737), .B(n26736), .Z(n26739) );
  ANDN U27761 ( .B(n26739), .A(n26738), .Z(n26741) );
  NANDN U27762 ( .A(n26741), .B(n26740), .Z(n26742) );
  NANDN U27763 ( .A(n26743), .B(n26742), .Z(n26745) );
  NAND U27764 ( .A(n26745), .B(n26744), .Z(n26747) );
  NAND U27765 ( .A(n26747), .B(n26746), .Z(n26748) );
  NANDN U27766 ( .A(n26749), .B(n26748), .Z(n26751) );
  NAND U27767 ( .A(n26751), .B(n26750), .Z(n26753) );
  ANDN U27768 ( .B(n26753), .A(n26752), .Z(n26755) );
  NANDN U27769 ( .A(n26755), .B(n26754), .Z(n26756) );
  AND U27770 ( .A(n26757), .B(n26756), .Z(n26759) );
  NANDN U27771 ( .A(n26759), .B(n26758), .Z(n26761) );
  NAND U27772 ( .A(n26761), .B(n26760), .Z(n26763) );
  NAND U27773 ( .A(n26763), .B(n26762), .Z(n26764) );
  NANDN U27774 ( .A(n26765), .B(n26764), .Z(n26767) );
  ANDN U27775 ( .B(n26767), .A(n26766), .Z(n26769) );
  NANDN U27776 ( .A(n26769), .B(n26768), .Z(n26771) );
  NAND U27777 ( .A(n26771), .B(n26770), .Z(n26773) );
  NAND U27778 ( .A(n26773), .B(n26772), .Z(n26774) );
  NANDN U27779 ( .A(n26775), .B(n26774), .Z(n26777) );
  ANDN U27780 ( .B(n26777), .A(n26776), .Z(n26779) );
  NANDN U27781 ( .A(n26779), .B(n26778), .Z(n26780) );
  NANDN U27782 ( .A(n26781), .B(n26780), .Z(n26783) );
  NAND U27783 ( .A(n26783), .B(n26782), .Z(n26784) );
  NANDN U27784 ( .A(n26785), .B(n26784), .Z(n26786) );
  AND U27785 ( .A(n26787), .B(n26786), .Z(n26789) );
  NANDN U27786 ( .A(n26789), .B(n26788), .Z(n26790) );
  NANDN U27787 ( .A(n26791), .B(n26790), .Z(n26793) );
  NAND U27788 ( .A(n26793), .B(n26792), .Z(n26795) );
  NAND U27789 ( .A(n26795), .B(n26794), .Z(n26797) );
  ANDN U27790 ( .B(n26797), .A(n26796), .Z(n26799) );
  NANDN U27791 ( .A(n26799), .B(n26798), .Z(n26803) );
  ANDN U27792 ( .B(n26801), .A(n26800), .Z(n26802) );
  NAND U27793 ( .A(n26803), .B(n26802), .Z(n26804) );
  NANDN U27794 ( .A(n26805), .B(n26804), .Z(n26806) );
  NANDN U27795 ( .A(n26807), .B(n26806), .Z(n26808) );
  NANDN U27796 ( .A(n26809), .B(n26808), .Z(n26811) );
  NAND U27797 ( .A(n26811), .B(n26810), .Z(n26812) );
  NANDN U27798 ( .A(n26813), .B(n26812), .Z(n26814) );
  AND U27799 ( .A(n26815), .B(n26814), .Z(n26817) );
  NANDN U27800 ( .A(n26817), .B(n26816), .Z(n26818) );
  NANDN U27801 ( .A(n26819), .B(n26818), .Z(n26821) );
  NAND U27802 ( .A(n26821), .B(n26820), .Z(n26823) );
  NAND U27803 ( .A(n26823), .B(n26822), .Z(n26825) );
  ANDN U27804 ( .B(n26825), .A(n26824), .Z(n26827) );
  NANDN U27805 ( .A(n26827), .B(n26826), .Z(n26828) );
  NANDN U27806 ( .A(n26829), .B(n26828), .Z(n26831) );
  NAND U27807 ( .A(n26831), .B(n26830), .Z(n26832) );
  NANDN U27808 ( .A(n26833), .B(n26832), .Z(n26835) );
  ANDN U27809 ( .B(n26835), .A(n26834), .Z(n26837) );
  NANDN U27810 ( .A(n26837), .B(n26836), .Z(n26839) );
  NAND U27811 ( .A(n26839), .B(n26838), .Z(n26841) );
  NAND U27812 ( .A(n26841), .B(n26840), .Z(n26842) );
  NANDN U27813 ( .A(n26843), .B(n26842), .Z(n26845) );
  ANDN U27814 ( .B(n26845), .A(n26844), .Z(n26847) );
  NANDN U27815 ( .A(n26847), .B(n26846), .Z(n26848) );
  NANDN U27816 ( .A(n26849), .B(n26848), .Z(n26851) );
  NAND U27817 ( .A(n26851), .B(n26850), .Z(n26852) );
  NANDN U27818 ( .A(n26853), .B(n26852), .Z(n26854) );
  AND U27819 ( .A(n26855), .B(n26854), .Z(n26857) );
  NANDN U27820 ( .A(n26857), .B(n26856), .Z(n26858) );
  NANDN U27821 ( .A(n26859), .B(n26858), .Z(n26861) );
  NAND U27822 ( .A(n26861), .B(n26860), .Z(n26863) );
  NAND U27823 ( .A(n26863), .B(n26862), .Z(n26865) );
  ANDN U27824 ( .B(n26865), .A(n26864), .Z(n26867) );
  NANDN U27825 ( .A(n26867), .B(n26866), .Z(n26868) );
  NANDN U27826 ( .A(n26869), .B(n26868), .Z(n26871) );
  NAND U27827 ( .A(n26871), .B(n26870), .Z(n26872) );
  NANDN U27828 ( .A(n26873), .B(n26872), .Z(n26875) );
  ANDN U27829 ( .B(n26875), .A(n26874), .Z(n26877) );
  NANDN U27830 ( .A(n26877), .B(n26876), .Z(n26879) );
  NAND U27831 ( .A(n26879), .B(n26878), .Z(n26881) );
  NAND U27832 ( .A(n26881), .B(n26880), .Z(n26882) );
  NANDN U27833 ( .A(n26883), .B(n26882), .Z(n26885) );
  ANDN U27834 ( .B(n26885), .A(n26884), .Z(n26887) );
  NANDN U27835 ( .A(n26887), .B(n26886), .Z(n26888) );
  NANDN U27836 ( .A(n26889), .B(n26888), .Z(n26891) );
  NAND U27837 ( .A(n26891), .B(n26890), .Z(n26892) );
  NANDN U27838 ( .A(n26893), .B(n26892), .Z(n26894) );
  AND U27839 ( .A(n26895), .B(n26894), .Z(n26897) );
  NANDN U27840 ( .A(n26897), .B(n26896), .Z(n26898) );
  NANDN U27841 ( .A(n26899), .B(n26898), .Z(n26901) );
  NAND U27842 ( .A(n26901), .B(n26900), .Z(n26903) );
  NAND U27843 ( .A(n26903), .B(n26902), .Z(n26905) );
  ANDN U27844 ( .B(n26905), .A(n26904), .Z(n26907) );
  NANDN U27845 ( .A(n26907), .B(n26906), .Z(n26908) );
  NANDN U27846 ( .A(n26909), .B(n26908), .Z(n26911) );
  NAND U27847 ( .A(n26911), .B(n26910), .Z(n26912) );
  NANDN U27848 ( .A(n26913), .B(n26912), .Z(n26915) );
  ANDN U27849 ( .B(n26915), .A(n26914), .Z(n26917) );
  NANDN U27850 ( .A(n26917), .B(n26916), .Z(n26919) );
  NAND U27851 ( .A(n26919), .B(n26918), .Z(n26921) );
  NAND U27852 ( .A(n26921), .B(n26920), .Z(n26922) );
  NANDN U27853 ( .A(n26923), .B(n26922), .Z(n26925) );
  ANDN U27854 ( .B(n26925), .A(n26924), .Z(n26927) );
  NANDN U27855 ( .A(n26927), .B(n26926), .Z(n26928) );
  NANDN U27856 ( .A(n26929), .B(n26928), .Z(n26931) );
  NAND U27857 ( .A(n26931), .B(n26930), .Z(n26932) );
  NANDN U27858 ( .A(n26933), .B(n26932), .Z(n26934) );
  AND U27859 ( .A(n26935), .B(n26934), .Z(n26937) );
  NANDN U27860 ( .A(n26937), .B(n26936), .Z(n26938) );
  NANDN U27861 ( .A(n26939), .B(n26938), .Z(n26941) );
  NAND U27862 ( .A(n26941), .B(n26940), .Z(n26943) );
  NAND U27863 ( .A(n26943), .B(n26942), .Z(n26945) );
  ANDN U27864 ( .B(n26945), .A(n26944), .Z(n26947) );
  NANDN U27865 ( .A(n26947), .B(n26946), .Z(n26948) );
  NANDN U27866 ( .A(n26949), .B(n26948), .Z(n26951) );
  NAND U27867 ( .A(n26951), .B(n26950), .Z(n26952) );
  NANDN U27868 ( .A(n26953), .B(n26952), .Z(n26955) );
  ANDN U27869 ( .B(n26955), .A(n26954), .Z(n26957) );
  NANDN U27870 ( .A(n26957), .B(n26956), .Z(n26959) );
  NAND U27871 ( .A(n26959), .B(n26958), .Z(n26961) );
  NAND U27872 ( .A(n26961), .B(n26960), .Z(n26962) );
  NANDN U27873 ( .A(n26963), .B(n26962), .Z(n26965) );
  ANDN U27874 ( .B(n26965), .A(n26964), .Z(n26967) );
  NANDN U27875 ( .A(n26967), .B(n26966), .Z(n26968) );
  NANDN U27876 ( .A(n26969), .B(n26968), .Z(n26971) );
  NAND U27877 ( .A(n26971), .B(n26970), .Z(n26973) );
  ANDN U27878 ( .B(n26973), .A(n26972), .Z(n26975) );
  NANDN U27879 ( .A(n26975), .B(n26974), .Z(n26976) );
  NANDN U27880 ( .A(n26977), .B(n26976), .Z(n26979) );
  NAND U27881 ( .A(n26979), .B(n26978), .Z(n26980) );
  NANDN U27882 ( .A(n26981), .B(n26980), .Z(n26983) );
  ANDN U27883 ( .B(n26983), .A(n26982), .Z(n26985) );
  NANDN U27884 ( .A(n26985), .B(n26984), .Z(n26986) );
  AND U27885 ( .A(n26987), .B(n26986), .Z(n26989) );
  NANDN U27886 ( .A(n26989), .B(n26988), .Z(n26990) );
  AND U27887 ( .A(n26991), .B(n26990), .Z(n26993) );
  NANDN U27888 ( .A(n26993), .B(n26992), .Z(n26994) );
  AND U27889 ( .A(n26995), .B(n26994), .Z(n26997) );
  NANDN U27890 ( .A(n26997), .B(n26996), .Z(n26999) );
  NAND U27891 ( .A(n26999), .B(n26998), .Z(n27001) );
  NAND U27892 ( .A(n27001), .B(n27000), .Z(n27002) );
  NANDN U27893 ( .A(n27003), .B(n27002), .Z(n27004) );
  AND U27894 ( .A(n27005), .B(n27004), .Z(n27007) );
  NANDN U27895 ( .A(n27007), .B(n27006), .Z(n27008) );
  NANDN U27896 ( .A(n27009), .B(n27008), .Z(n27011) );
  NAND U27897 ( .A(n27011), .B(n27010), .Z(n27013) );
  NAND U27898 ( .A(n27013), .B(n27012), .Z(n27015) );
  ANDN U27899 ( .B(n27015), .A(n27014), .Z(n27017) );
  NANDN U27900 ( .A(n27017), .B(n27016), .Z(n27018) );
  NANDN U27901 ( .A(n27019), .B(n27018), .Z(n27021) );
  NAND U27902 ( .A(n27021), .B(n27020), .Z(n27022) );
  NANDN U27903 ( .A(n27023), .B(n27022), .Z(n27024) );
  AND U27904 ( .A(n27025), .B(n27024), .Z(n27027) );
  NANDN U27905 ( .A(n27027), .B(n27026), .Z(n27028) );
  NANDN U27906 ( .A(n27029), .B(n27028), .Z(n27031) );
  NAND U27907 ( .A(n27031), .B(n27030), .Z(n27032) );
  NANDN U27908 ( .A(n27033), .B(n27032), .Z(n27035) );
  ANDN U27909 ( .B(n27035), .A(n27034), .Z(n27037) );
  NANDN U27910 ( .A(n27037), .B(n27036), .Z(n27038) );
  NANDN U27911 ( .A(n27039), .B(n27038), .Z(n27041) );
  NAND U27912 ( .A(n27041), .B(n27040), .Z(n27042) );
  NANDN U27913 ( .A(n27043), .B(n27042), .Z(n27045) );
  ANDN U27914 ( .B(n27045), .A(n27044), .Z(n27047) );
  NANDN U27915 ( .A(n27047), .B(n27046), .Z(n27049) );
  NAND U27916 ( .A(n27049), .B(n27048), .Z(n27051) );
  NAND U27917 ( .A(n27051), .B(n27050), .Z(n27052) );
  NANDN U27918 ( .A(n27053), .B(n27052), .Z(n27055) );
  ANDN U27919 ( .B(n27055), .A(n27054), .Z(n27057) );
  NANDN U27920 ( .A(n27057), .B(n27056), .Z(n27058) );
  NANDN U27921 ( .A(n27059), .B(n27058), .Z(n27061) );
  NAND U27922 ( .A(n27061), .B(n27060), .Z(n27062) );
  NANDN U27923 ( .A(n27063), .B(n27062), .Z(n27065) );
  ANDN U27924 ( .B(n27065), .A(n27064), .Z(n27067) );
  NANDN U27925 ( .A(n27067), .B(n27066), .Z(n27068) );
  NANDN U27926 ( .A(n27069), .B(n27068), .Z(n27071) );
  NAND U27927 ( .A(n27071), .B(n27070), .Z(n27073) );
  NAND U27928 ( .A(n27073), .B(n27072), .Z(n27075) );
  ANDN U27929 ( .B(n27075), .A(n27074), .Z(n27077) );
  NANDN U27930 ( .A(n27077), .B(n27076), .Z(n27078) );
  NANDN U27931 ( .A(n27079), .B(n27078), .Z(n27081) );
  NAND U27932 ( .A(n27081), .B(n27080), .Z(n27082) );
  NANDN U27933 ( .A(n27083), .B(n27082), .Z(n27084) );
  AND U27934 ( .A(n27085), .B(n27084), .Z(n27087) );
  NANDN U27935 ( .A(n27087), .B(n27086), .Z(n27088) );
  NANDN U27936 ( .A(n27089), .B(n27088), .Z(n27091) );
  NAND U27937 ( .A(n27091), .B(n27090), .Z(n27092) );
  NANDN U27938 ( .A(n27093), .B(n27092), .Z(n27094) );
  AND U27939 ( .A(n27095), .B(n27094), .Z(n27096) );
  OR U27940 ( .A(n27097), .B(n27096), .Z(n27098) );
  NANDN U27941 ( .A(n27099), .B(n27098), .Z(n27101) );
  NAND U27942 ( .A(n27101), .B(n27100), .Z(n27103) );
  NAND U27943 ( .A(n27103), .B(n27102), .Z(n27105) );
  ANDN U27944 ( .B(n27105), .A(n27104), .Z(n27109) );
  ANDN U27945 ( .B(n27107), .A(n27106), .Z(n27108) );
  NANDN U27946 ( .A(n27109), .B(n27108), .Z(n27111) );
  NAND U27947 ( .A(n27111), .B(n27110), .Z(n27112) );
  AND U27948 ( .A(n27113), .B(n27112), .Z(n27115) );
  NANDN U27949 ( .A(n27115), .B(n27114), .Z(n27116) );
  NANDN U27950 ( .A(n27117), .B(n27116), .Z(n27119) );
  NAND U27951 ( .A(n27119), .B(n27118), .Z(n27120) );
  NANDN U27952 ( .A(n27121), .B(n27120), .Z(n27123) );
  ANDN U27953 ( .B(n27123), .A(n27122), .Z(n27125) );
  NANDN U27954 ( .A(n27125), .B(n27124), .Z(n27127) );
  ANDN U27955 ( .B(n27127), .A(n27126), .Z(n27129) );
  NANDN U27956 ( .A(n27129), .B(n27128), .Z(n27131) );
  ANDN U27957 ( .B(n27131), .A(n27130), .Z(n27132) );
  OR U27958 ( .A(n27133), .B(n27132), .Z(n27134) );
  NANDN U27959 ( .A(n27135), .B(n27134), .Z(n27136) );
  NANDN U27960 ( .A(n27137), .B(n27136), .Z(n27139) );
  NANDN U27961 ( .A(n27139), .B(n27138), .Z(n27141) );
  NAND U27962 ( .A(n27141), .B(n27140), .Z(n27142) );
  AND U27963 ( .A(n27143), .B(n27142), .Z(n27145) );
  NANDN U27964 ( .A(n27145), .B(n27144), .Z(n27146) );
  NANDN U27965 ( .A(n27147), .B(n27146), .Z(n27148) );
  NANDN U27966 ( .A(n27149), .B(n27148), .Z(n27151) );
  NAND U27967 ( .A(n27151), .B(n27150), .Z(n27152) );
  AND U27968 ( .A(n27153), .B(n27152), .Z(n27155) );
  NANDN U27969 ( .A(n27155), .B(n27154), .Z(n27156) );
  NANDN U27970 ( .A(n27157), .B(n27156), .Z(n27158) );
  NANDN U27971 ( .A(n27159), .B(n27158), .Z(n27161) );
  NAND U27972 ( .A(n27161), .B(n27160), .Z(n27163) );
  ANDN U27973 ( .B(n27163), .A(n27162), .Z(n27165) );
  NANDN U27974 ( .A(n27165), .B(n27164), .Z(n27166) );
  NANDN U27975 ( .A(n27167), .B(n27166), .Z(n27169) );
  NAND U27976 ( .A(n27169), .B(n27168), .Z(n27171) );
  ANDN U27977 ( .B(n27171), .A(n27170), .Z(n27173) );
  NAND U27978 ( .A(n27173), .B(n27172), .Z(n27175) );
  NAND U27979 ( .A(n27175), .B(n27174), .Z(n27177) );
  ANDN U27980 ( .B(n27177), .A(n27176), .Z(n27179) );
  NAND U27981 ( .A(n27179), .B(n27178), .Z(n27181) );
  NAND U27982 ( .A(n27181), .B(n27180), .Z(n27182) );
  AND U27983 ( .A(n27183), .B(n27182), .Z(n27185) );
  NANDN U27984 ( .A(n27185), .B(n27184), .Z(n27186) );
  NANDN U27985 ( .A(n27187), .B(n27186), .Z(n27188) );
  NANDN U27986 ( .A(n27189), .B(n27188), .Z(n27191) );
  NAND U27987 ( .A(n27191), .B(n27190), .Z(n27193) );
  ANDN U27988 ( .B(n27193), .A(n27192), .Z(n27197) );
  ANDN U27989 ( .B(n27195), .A(n27194), .Z(n27196) );
  NANDN U27990 ( .A(n27197), .B(n27196), .Z(n27199) );
  NAND U27991 ( .A(n27199), .B(n27198), .Z(n27201) );
  ANDN U27992 ( .B(n27201), .A(n27200), .Z(n27203) );
  NANDN U27993 ( .A(n27203), .B(n27202), .Z(n27205) );
  NAND U27994 ( .A(n27205), .B(n27204), .Z(n27206) );
  NANDN U27995 ( .A(n27207), .B(n27206), .Z(n27209) );
  NAND U27996 ( .A(n27209), .B(n27208), .Z(n27211) );
  ANDN U27997 ( .B(n27211), .A(n27210), .Z(n27213) );
  NANDN U27998 ( .A(n27213), .B(n27212), .Z(n27214) );
  NANDN U27999 ( .A(n27215), .B(n27214), .Z(n27216) );
  NANDN U28000 ( .A(n27217), .B(n27216), .Z(n27219) );
  NAND U28001 ( .A(n27219), .B(n27218), .Z(n27221) );
  ANDN U28002 ( .B(n27221), .A(n27220), .Z(n27223) );
  NANDN U28003 ( .A(n27223), .B(n27222), .Z(n27224) );
  AND U28004 ( .A(n27225), .B(n27224), .Z(n27227) );
  NANDN U28005 ( .A(n27227), .B(n27226), .Z(n27229) );
  ANDN U28006 ( .B(n27229), .A(n27228), .Z(n27231) );
  NANDN U28007 ( .A(n27231), .B(n27230), .Z(n27233) );
  ANDN U28008 ( .B(n27233), .A(n27232), .Z(n27235) );
  NANDN U28009 ( .A(n27235), .B(n27234), .Z(n27236) );
  NANDN U28010 ( .A(n27237), .B(n27236), .Z(n27239) );
  NAND U28011 ( .A(n27239), .B(n27238), .Z(n27241) );
  NAND U28012 ( .A(n27241), .B(n27240), .Z(n27243) );
  ANDN U28013 ( .B(n27243), .A(n27242), .Z(n27247) );
  ANDN U28014 ( .B(n27245), .A(n27244), .Z(n27246) );
  NANDN U28015 ( .A(n27247), .B(n27246), .Z(n27249) );
  NAND U28016 ( .A(n27249), .B(n27248), .Z(n27250) );
  AND U28017 ( .A(n27251), .B(n27250), .Z(n27253) );
  NANDN U28018 ( .A(n27253), .B(n27252), .Z(n27254) );
  NANDN U28019 ( .A(n27255), .B(n27254), .Z(n27256) );
  NANDN U28020 ( .A(n27257), .B(n27256), .Z(n27259) );
  NAND U28021 ( .A(n27259), .B(n27258), .Z(n27261) );
  ANDN U28022 ( .B(n27261), .A(n27260), .Z(n27263) );
  NANDN U28023 ( .A(n27263), .B(n27262), .Z(n27264) );
  NANDN U28024 ( .A(n27265), .B(n27264), .Z(n27267) );
  NAND U28025 ( .A(n27267), .B(n27266), .Z(n27269) );
  NAND U28026 ( .A(n27269), .B(n27268), .Z(n27271) );
  ANDN U28027 ( .B(n27271), .A(n27270), .Z(n27273) );
  NANDN U28028 ( .A(n27273), .B(n27272), .Z(n27275) );
  NAND U28029 ( .A(n27275), .B(n27274), .Z(n27276) );
  NANDN U28030 ( .A(n27277), .B(n27276), .Z(n27279) );
  NAND U28031 ( .A(n27279), .B(n27278), .Z(n27281) );
  ANDN U28032 ( .B(n27281), .A(n27280), .Z(n27283) );
  NANDN U28033 ( .A(n27283), .B(n27282), .Z(n27284) );
  NANDN U28034 ( .A(n27285), .B(n27284), .Z(n27287) );
  NAND U28035 ( .A(n27287), .B(n27286), .Z(n27289) );
  NANDN U28036 ( .A(n27289), .B(n27288), .Z(n27291) );
  NAND U28037 ( .A(n27291), .B(n27290), .Z(n27292) );
  AND U28038 ( .A(n27293), .B(n27292), .Z(n27295) );
  NANDN U28039 ( .A(n27295), .B(n27294), .Z(n27296) );
  NANDN U28040 ( .A(n27297), .B(n27296), .Z(n27299) );
  NAND U28041 ( .A(n27299), .B(n27298), .Z(n27301) );
  NAND U28042 ( .A(n27301), .B(n27300), .Z(n27303) );
  ANDN U28043 ( .B(n27303), .A(n27302), .Z(n27305) );
  NANDN U28044 ( .A(n27305), .B(n27304), .Z(n27307) );
  NAND U28045 ( .A(n27307), .B(n27306), .Z(n27308) );
  NANDN U28046 ( .A(n27309), .B(n27308), .Z(n27311) );
  NAND U28047 ( .A(n27311), .B(n27310), .Z(n27313) );
  ANDN U28048 ( .B(n27313), .A(n27312), .Z(n27315) );
  NANDN U28049 ( .A(n27315), .B(n27314), .Z(n27316) );
  NANDN U28050 ( .A(n27317), .B(n27316), .Z(n27319) );
  NAND U28051 ( .A(n27319), .B(n27318), .Z(n27321) );
  NAND U28052 ( .A(n27321), .B(n27320), .Z(n27323) );
  ANDN U28053 ( .B(n27323), .A(n27322), .Z(n27325) );
  NANDN U28054 ( .A(n27325), .B(n27324), .Z(n27326) );
  NANDN U28055 ( .A(n27327), .B(n27326), .Z(n27328) );
  NANDN U28056 ( .A(n27329), .B(n27328), .Z(n27330) );
  NANDN U28057 ( .A(n27331), .B(n27330), .Z(n27332) );
  AND U28058 ( .A(n27333), .B(n27332), .Z(n27334) );
  OR U28059 ( .A(n27335), .B(n27334), .Z(n27336) );
  NANDN U28060 ( .A(n27337), .B(n27336), .Z(n27338) );
  NANDN U28061 ( .A(n27339), .B(n27338), .Z(n27341) );
  NAND U28062 ( .A(n27341), .B(n27340), .Z(n27342) );
  AND U28063 ( .A(n27343), .B(n27342), .Z(n27344) );
  OR U28064 ( .A(n27345), .B(n27344), .Z(n27346) );
  NANDN U28065 ( .A(n27347), .B(n27346), .Z(n27348) );
  NANDN U28066 ( .A(n27349), .B(n27348), .Z(n27351) );
  NAND U28067 ( .A(n27351), .B(n27350), .Z(n27353) );
  ANDN U28068 ( .B(n27353), .A(n27352), .Z(n27354) );
  OR U28069 ( .A(n27355), .B(n27354), .Z(n27356) );
  NANDN U28070 ( .A(n27357), .B(n27356), .Z(n27359) );
  NAND U28071 ( .A(n27359), .B(n27358), .Z(n27361) );
  NAND U28072 ( .A(n27361), .B(n27360), .Z(n27363) );
  ANDN U28073 ( .B(n27363), .A(n27362), .Z(n27364) );
  OR U28074 ( .A(n27365), .B(n27364), .Z(n27366) );
  NANDN U28075 ( .A(n27367), .B(n27366), .Z(n27368) );
  NANDN U28076 ( .A(n27369), .B(n27368), .Z(n27371) );
  NAND U28077 ( .A(n27371), .B(n27370), .Z(n27373) );
  ANDN U28078 ( .B(n27373), .A(n27372), .Z(n27375) );
  NANDN U28079 ( .A(n27375), .B(n27374), .Z(n27376) );
  NANDN U28080 ( .A(n27377), .B(n27376), .Z(n27378) );
  NANDN U28081 ( .A(n27379), .B(n27378), .Z(n27381) );
  NAND U28082 ( .A(n27381), .B(n27380), .Z(n27382) );
  AND U28083 ( .A(n27383), .B(n27382), .Z(n27384) );
  OR U28084 ( .A(n27385), .B(n27384), .Z(n27386) );
  NANDN U28085 ( .A(n27387), .B(n27386), .Z(n27388) );
  NANDN U28086 ( .A(n27389), .B(n27388), .Z(n27391) );
  NAND U28087 ( .A(n27391), .B(n27390), .Z(n27393) );
  ANDN U28088 ( .B(n27393), .A(n27392), .Z(n27394) );
  OR U28089 ( .A(n27395), .B(n27394), .Z(n27396) );
  NANDN U28090 ( .A(n27397), .B(n27396), .Z(n27399) );
  NAND U28091 ( .A(n27399), .B(n27398), .Z(n27401) );
  NAND U28092 ( .A(n27401), .B(n27400), .Z(n27403) );
  ANDN U28093 ( .B(n27403), .A(n27402), .Z(n27404) );
  OR U28094 ( .A(n27405), .B(n27404), .Z(n27406) );
  NANDN U28095 ( .A(n27407), .B(n27406), .Z(n27409) );
  NAND U28096 ( .A(n27409), .B(n27408), .Z(n27411) );
  NANDN U28097 ( .A(n27411), .B(n27410), .Z(n27412) );
  NANDN U28098 ( .A(n27413), .B(n27412), .Z(n27415) );
  ANDN U28099 ( .B(n27415), .A(n27414), .Z(n27416) );
  OR U28100 ( .A(n27417), .B(n27416), .Z(n27418) );
  NANDN U28101 ( .A(n27419), .B(n27418), .Z(n27420) );
  NANDN U28102 ( .A(n27421), .B(n27420), .Z(n27422) );
  NANDN U28103 ( .A(n27423), .B(n27422), .Z(n27425) );
  ANDN U28104 ( .B(n27425), .A(n27424), .Z(n27429) );
  ANDN U28105 ( .B(n27427), .A(n27426), .Z(n27428) );
  NANDN U28106 ( .A(n27429), .B(n27428), .Z(n27431) );
  NAND U28107 ( .A(n27431), .B(n27430), .Z(n27433) );
  ANDN U28108 ( .B(n27433), .A(n27432), .Z(n27435) );
  NANDN U28109 ( .A(n27435), .B(n27434), .Z(n27436) );
  NANDN U28110 ( .A(n27437), .B(n27436), .Z(n27439) );
  NAND U28111 ( .A(n27439), .B(n27438), .Z(n27440) );
  NANDN U28112 ( .A(n27441), .B(n27440), .Z(n27443) );
  ANDN U28113 ( .B(n27443), .A(n27442), .Z(n27444) );
  OR U28114 ( .A(n27445), .B(n27444), .Z(n27446) );
  NANDN U28115 ( .A(n27447), .B(n27446), .Z(n27448) );
  NANDN U28116 ( .A(n27449), .B(n27448), .Z(n27451) );
  NAND U28117 ( .A(n27451), .B(n27450), .Z(n27453) );
  NAND U28118 ( .A(n27453), .B(n27452), .Z(n27454) );
  AND U28119 ( .A(n27455), .B(n27454), .Z(n27457) );
  NANDN U28120 ( .A(n27457), .B(n27456), .Z(n27458) );
  AND U28121 ( .A(n27459), .B(n27458), .Z(n27461) );
  NANDN U28122 ( .A(n27461), .B(n27460), .Z(n27462) );
  NANDN U28123 ( .A(n27463), .B(n27462), .Z(n27465) );
  NAND U28124 ( .A(n27465), .B(n27464), .Z(n27466) );
  NANDN U28125 ( .A(n27467), .B(n27466), .Z(n27469) );
  ANDN U28126 ( .B(n27469), .A(n27468), .Z(n27470) );
  OR U28127 ( .A(n27471), .B(n27470), .Z(n27472) );
  NANDN U28128 ( .A(n27473), .B(n27472), .Z(n27474) );
  NANDN U28129 ( .A(n27475), .B(n27474), .Z(n27477) );
  AND U28130 ( .A(n27477), .B(n27476), .Z(n27479) );
  NAND U28131 ( .A(n27479), .B(n27478), .Z(n27481) );
  NAND U28132 ( .A(n27481), .B(n27480), .Z(n27482) );
  NANDN U28133 ( .A(n27483), .B(n27482), .Z(n27484) );
  NANDN U28134 ( .A(n27485), .B(n27484), .Z(n27487) );
  NAND U28135 ( .A(n27487), .B(n27486), .Z(n27488) );
  NANDN U28136 ( .A(n27489), .B(n27488), .Z(n27491) );
  ANDN U28137 ( .B(n27491), .A(n27490), .Z(n27493) );
  NANDN U28138 ( .A(n27493), .B(n27492), .Z(n27494) );
  NANDN U28139 ( .A(n27495), .B(n27494), .Z(n27497) );
  NAND U28140 ( .A(n27497), .B(n27496), .Z(n27498) );
  NANDN U28141 ( .A(n27499), .B(n27498), .Z(n27501) );
  ANDN U28142 ( .B(n27501), .A(n27500), .Z(n27502) );
  OR U28143 ( .A(n27503), .B(n27502), .Z(n27504) );
  NANDN U28144 ( .A(n27505), .B(n27504), .Z(n27506) );
  NANDN U28145 ( .A(n27507), .B(n27506), .Z(n27509) );
  NAND U28146 ( .A(n27509), .B(n27508), .Z(n27511) );
  ANDN U28147 ( .B(n27511), .A(n27510), .Z(n27513) );
  NANDN U28148 ( .A(n27513), .B(n27512), .Z(n27514) );
  NANDN U28149 ( .A(n27515), .B(n27514), .Z(n27516) );
  NANDN U28150 ( .A(n27517), .B(n27516), .Z(n27518) );
  NANDN U28151 ( .A(n27519), .B(n27518), .Z(n27521) );
  ANDN U28152 ( .B(n27521), .A(n27520), .Z(n27525) );
  ANDN U28153 ( .B(n27523), .A(n27522), .Z(n27524) );
  NANDN U28154 ( .A(n27525), .B(n27524), .Z(n27527) );
  NAND U28155 ( .A(n27527), .B(n27526), .Z(n27529) );
  ANDN U28156 ( .B(n27529), .A(n27528), .Z(n27531) );
  NANDN U28157 ( .A(n27531), .B(n27530), .Z(n27532) );
  NANDN U28158 ( .A(n27533), .B(n27532), .Z(n27534) );
  NANDN U28159 ( .A(n27535), .B(n27534), .Z(n27536) );
  NANDN U28160 ( .A(n27537), .B(n27536), .Z(n27539) );
  ANDN U28161 ( .B(n27539), .A(n27538), .Z(n27543) );
  ANDN U28162 ( .B(n27541), .A(n27540), .Z(n27542) );
  NANDN U28163 ( .A(n27543), .B(n27542), .Z(n27545) );
  NAND U28164 ( .A(n27545), .B(n27544), .Z(n27547) );
  ANDN U28165 ( .B(n27547), .A(n27546), .Z(n27549) );
  NANDN U28166 ( .A(n27549), .B(n27548), .Z(n27550) );
  NANDN U28167 ( .A(n27551), .B(n27550), .Z(n27553) );
  NAND U28168 ( .A(n27553), .B(n27552), .Z(n27554) );
  NANDN U28169 ( .A(n27555), .B(n27554), .Z(n27557) );
  ANDN U28170 ( .B(n27557), .A(n27556), .Z(n27558) );
  OR U28171 ( .A(n27559), .B(n27558), .Z(n27560) );
  NANDN U28172 ( .A(n27561), .B(n27560), .Z(n27563) );
  NAND U28173 ( .A(n27563), .B(n27562), .Z(n27565) );
  NANDN U28174 ( .A(n27565), .B(n27564), .Z(n27567) );
  NAND U28175 ( .A(n27567), .B(n27566), .Z(n27569) );
  ANDN U28176 ( .B(n27569), .A(n27568), .Z(n27571) );
  NANDN U28177 ( .A(n27571), .B(n27570), .Z(n27572) );
  NANDN U28178 ( .A(n27573), .B(n27572), .Z(n27575) );
  NAND U28179 ( .A(n27575), .B(n27574), .Z(n27576) );
  NANDN U28180 ( .A(n27577), .B(n27576), .Z(n27579) );
  ANDN U28181 ( .B(n27579), .A(n27578), .Z(n27580) );
  OR U28182 ( .A(n27581), .B(n27580), .Z(n27583) );
  NAND U28183 ( .A(n27583), .B(n27582), .Z(n27585) );
  NAND U28184 ( .A(n27585), .B(n27584), .Z(n27587) );
  NAND U28185 ( .A(n27587), .B(n27586), .Z(n27589) );
  ANDN U28186 ( .B(n27589), .A(n27588), .Z(n27591) );
  NANDN U28187 ( .A(n27591), .B(n27590), .Z(n27592) );
  NANDN U28188 ( .A(n27593), .B(n27592), .Z(n27595) );
  NAND U28189 ( .A(n27595), .B(n27594), .Z(n27596) );
  NANDN U28190 ( .A(n27597), .B(n27596), .Z(n27599) );
  ANDN U28191 ( .B(n27599), .A(n27598), .Z(n27600) );
  ANDN U28192 ( .B(n27601), .A(n27600), .Z(n27603) );
  NANDN U28193 ( .A(n27603), .B(n27602), .Z(n27607) );
  ANDN U28194 ( .B(n27605), .A(n27604), .Z(n27606) );
  NAND U28195 ( .A(n27607), .B(n27606), .Z(n27609) );
  NAND U28196 ( .A(n27609), .B(n27608), .Z(n27611) );
  NAND U28197 ( .A(n27611), .B(n27610), .Z(n27612) );
  NANDN U28198 ( .A(n27613), .B(n27612), .Z(n27615) );
  NAND U28199 ( .A(n27615), .B(n27614), .Z(n27616) );
  NANDN U28200 ( .A(n27617), .B(n27616), .Z(n27619) );
  ANDN U28201 ( .B(n27619), .A(n27618), .Z(n27620) );
  OR U28202 ( .A(n27621), .B(n27620), .Z(n27622) );
  NANDN U28203 ( .A(n27623), .B(n27622), .Z(n27624) );
  NANDN U28204 ( .A(n27625), .B(n27624), .Z(n27627) );
  AND U28205 ( .A(n27627), .B(n27626), .Z(n27629) );
  NAND U28206 ( .A(n27629), .B(n27628), .Z(n27630) );
  NANDN U28207 ( .A(n27631), .B(n27630), .Z(n27632) );
  NANDN U28208 ( .A(n27633), .B(n27632), .Z(n27635) );
  NAND U28209 ( .A(n27635), .B(n27634), .Z(n27637) );
  NAND U28210 ( .A(n27637), .B(n27636), .Z(n27638) );
  NANDN U28211 ( .A(n27639), .B(n27638), .Z(n27641) );
  ANDN U28212 ( .B(n27641), .A(n27640), .Z(n27643) );
  NANDN U28213 ( .A(n27643), .B(n27642), .Z(n27644) );
  NANDN U28214 ( .A(n27645), .B(n27644), .Z(n27647) );
  NAND U28215 ( .A(n27647), .B(n27646), .Z(n27648) );
  NANDN U28216 ( .A(n27649), .B(n27648), .Z(n27651) );
  ANDN U28217 ( .B(n27651), .A(n27650), .Z(n27655) );
  NOR U28218 ( .A(n27653), .B(n27652), .Z(n27654) );
  NANDN U28219 ( .A(n27655), .B(n27654), .Z(n27656) );
  NANDN U28220 ( .A(n27657), .B(n27656), .Z(n27659) );
  ANDN U28221 ( .B(n27659), .A(n27658), .Z(n27661) );
  NANDN U28222 ( .A(n27661), .B(n27660), .Z(n27665) );
  NOR U28223 ( .A(n27663), .B(n27662), .Z(n27664) );
  NAND U28224 ( .A(n27665), .B(n27664), .Z(n27667) );
  NAND U28225 ( .A(n27667), .B(n27666), .Z(n27668) );
  NANDN U28226 ( .A(n27669), .B(n27668), .Z(n27670) );
  NANDN U28227 ( .A(n27671), .B(n27670), .Z(n27672) );
  NANDN U28228 ( .A(n27673), .B(n27672), .Z(n27675) );
  NAND U28229 ( .A(n27675), .B(n27674), .Z(n27677) );
  ANDN U28230 ( .B(n27677), .A(n27676), .Z(n27678) );
  OR U28231 ( .A(n27679), .B(n27678), .Z(n27680) );
  NANDN U28232 ( .A(n27681), .B(n27680), .Z(n27683) );
  NAND U28233 ( .A(n27683), .B(n27682), .Z(n27685) );
  ANDN U28234 ( .B(n27685), .A(n27684), .Z(n27686) );
  NANDN U28235 ( .A(n27687), .B(n27686), .Z(n27689) );
  NAND U28236 ( .A(n27689), .B(n27688), .Z(n27691) );
  ANDN U28237 ( .B(n27691), .A(n27690), .Z(n27693) );
  NAND U28238 ( .A(n27693), .B(n27692), .Z(n27695) );
  NAND U28239 ( .A(n27695), .B(n27694), .Z(n27697) );
  ANDN U28240 ( .B(n27697), .A(n27696), .Z(n27698) );
  OR U28241 ( .A(n27699), .B(n27698), .Z(n27703) );
  NOR U28242 ( .A(n27701), .B(n27700), .Z(n27702) );
  NAND U28243 ( .A(n27703), .B(n27702), .Z(n27705) );
  NAND U28244 ( .A(n27705), .B(n27704), .Z(n27706) );
  AND U28245 ( .A(n27707), .B(n27706), .Z(n27709) );
  NAND U28246 ( .A(n27709), .B(n27708), .Z(n27711) );
  NAND U28247 ( .A(n27711), .B(n27710), .Z(n27712) );
  AND U28248 ( .A(n27713), .B(n27712), .Z(n27715) );
  NANDN U28249 ( .A(n27715), .B(n27714), .Z(n27717) );
  NAND U28250 ( .A(n27717), .B(n27716), .Z(n27718) );
  NANDN U28251 ( .A(n27719), .B(n27718), .Z(n27721) );
  NAND U28252 ( .A(n27721), .B(n27720), .Z(n27723) );
  ANDN U28253 ( .B(n27723), .A(n27722), .Z(n27725) );
  NANDN U28254 ( .A(n27725), .B(n27724), .Z(n27726) );
  NANDN U28255 ( .A(n27727), .B(n27726), .Z(n27729) );
  NAND U28256 ( .A(n27729), .B(n27728), .Z(n27731) );
  NAND U28257 ( .A(n27731), .B(n27730), .Z(n27733) );
  ANDN U28258 ( .B(n27733), .A(n27732), .Z(n27735) );
  NANDN U28259 ( .A(n27735), .B(n27734), .Z(n27739) );
  AND U28260 ( .A(n27737), .B(n27736), .Z(n27738) );
  NAND U28261 ( .A(n27739), .B(n27738), .Z(n27740) );
  NANDN U28262 ( .A(n27741), .B(n27740), .Z(n27742) );
  NANDN U28263 ( .A(n27743), .B(n27742), .Z(n27745) );
  NAND U28264 ( .A(n27745), .B(n27744), .Z(n27747) );
  NAND U28265 ( .A(n27747), .B(n27746), .Z(n27748) );
  NANDN U28266 ( .A(n27749), .B(n27748), .Z(n27751) );
  ANDN U28267 ( .B(n27751), .A(n27750), .Z(n27753) );
  NANDN U28268 ( .A(n27753), .B(n27752), .Z(n27757) );
  NOR U28269 ( .A(n27755), .B(n27754), .Z(n27756) );
  NAND U28270 ( .A(n27757), .B(n27756), .Z(n27759) );
  NAND U28271 ( .A(n27759), .B(n27758), .Z(n27760) );
  AND U28272 ( .A(n27761), .B(n27760), .Z(n27763) );
  NANDN U28273 ( .A(n27763), .B(n27762), .Z(n27764) );
  AND U28274 ( .A(n27765), .B(n27764), .Z(n27767) );
  NANDN U28275 ( .A(n27767), .B(n27766), .Z(n27769) );
  NAND U28276 ( .A(n27769), .B(n27768), .Z(n27771) );
  NAND U28277 ( .A(n27771), .B(n27770), .Z(n27773) );
  NAND U28278 ( .A(n27773), .B(n27772), .Z(n27775) );
  ANDN U28279 ( .B(n27775), .A(n27774), .Z(n27777) );
  NANDN U28280 ( .A(n27777), .B(n27776), .Z(n27778) );
  NANDN U28281 ( .A(n27779), .B(n27778), .Z(n27781) );
  NAND U28282 ( .A(n27781), .B(n27780), .Z(n27782) );
  NANDN U28283 ( .A(n27783), .B(n27782), .Z(n27785) );
  ANDN U28284 ( .B(n27785), .A(n27784), .Z(n27787) );
  NANDN U28285 ( .A(n27787), .B(n27786), .Z(n27791) );
  AND U28286 ( .A(n27789), .B(n27788), .Z(n27790) );
  NAND U28287 ( .A(n27791), .B(n27790), .Z(n27792) );
  NANDN U28288 ( .A(n27793), .B(n27792), .Z(n27794) );
  NANDN U28289 ( .A(n27795), .B(n27794), .Z(n27797) );
  NAND U28290 ( .A(n27797), .B(n27796), .Z(n27799) );
  NAND U28291 ( .A(n27799), .B(n27798), .Z(n27800) );
  NANDN U28292 ( .A(n27801), .B(n27800), .Z(n27803) );
  ANDN U28293 ( .B(n27803), .A(n27802), .Z(n27805) );
  NANDN U28294 ( .A(n27805), .B(n27804), .Z(n27809) );
  ANDN U28295 ( .B(n27807), .A(n27806), .Z(n27808) );
  NAND U28296 ( .A(n27809), .B(n27808), .Z(n27811) );
  NAND U28297 ( .A(n27811), .B(n27810), .Z(n27813) );
  ANDN U28298 ( .B(n27813), .A(n27812), .Z(n27815) );
  NAND U28299 ( .A(n27815), .B(n27814), .Z(n27817) );
  NAND U28300 ( .A(n27817), .B(n27816), .Z(n27819) );
  ANDN U28301 ( .B(n27819), .A(n27818), .Z(n27820) );
  OR U28302 ( .A(n27821), .B(n27820), .Z(n27825) );
  ANDN U28303 ( .B(n27823), .A(n27822), .Z(n27824) );
  NAND U28304 ( .A(n27825), .B(n27824), .Z(n27826) );
  NANDN U28305 ( .A(n27827), .B(n27826), .Z(n27828) );
  NANDN U28306 ( .A(n27829), .B(n27828), .Z(n27831) );
  ANDN U28307 ( .B(n27831), .A(n27830), .Z(n27832) );
  OR U28308 ( .A(n27833), .B(n27832), .Z(n27834) );
  NANDN U28309 ( .A(n27835), .B(n27834), .Z(n27837) );
  NAND U28310 ( .A(n27837), .B(n27836), .Z(n27839) );
  NANDN U28311 ( .A(n27839), .B(n27838), .Z(n27840) );
  NANDN U28312 ( .A(n27841), .B(n27840), .Z(n27843) );
  ANDN U28313 ( .B(n27843), .A(n27842), .Z(n27844) );
  OR U28314 ( .A(n27845), .B(n27844), .Z(n27846) );
  NANDN U28315 ( .A(n27847), .B(n27846), .Z(n27849) );
  NAND U28316 ( .A(n27849), .B(n27848), .Z(n27850) );
  NANDN U28317 ( .A(n27851), .B(n27850), .Z(n27853) );
  ANDN U28318 ( .B(n27853), .A(n27852), .Z(n27854) );
  OR U28319 ( .A(n27855), .B(n27854), .Z(n27856) );
  NANDN U28320 ( .A(n27857), .B(n27856), .Z(n27858) );
  NANDN U28321 ( .A(n27859), .B(n27858), .Z(n27861) );
  NAND U28322 ( .A(n27861), .B(n27860), .Z(n27863) );
  ANDN U28323 ( .B(n27863), .A(n27862), .Z(n27865) );
  NANDN U28324 ( .A(n27865), .B(n27864), .Z(n27866) );
  NANDN U28325 ( .A(n27867), .B(n27866), .Z(n27869) );
  NAND U28326 ( .A(n27869), .B(n27868), .Z(n27870) );
  NANDN U28327 ( .A(n27871), .B(n27870), .Z(n27873) );
  ANDN U28328 ( .B(n27873), .A(n27872), .Z(n27874) );
  OR U28329 ( .A(n27875), .B(n27874), .Z(n27876) );
  NANDN U28330 ( .A(n27877), .B(n27876), .Z(n27878) );
  NANDN U28331 ( .A(n27879), .B(n27878), .Z(n27881) );
  NAND U28332 ( .A(n27881), .B(n27880), .Z(n27883) );
  ANDN U28333 ( .B(n27883), .A(n27882), .Z(n27885) );
  NANDN U28334 ( .A(n27885), .B(n27884), .Z(n27886) );
  NANDN U28335 ( .A(n27887), .B(n27886), .Z(n27889) );
  NAND U28336 ( .A(n27889), .B(n27888), .Z(n27890) );
  NANDN U28337 ( .A(n27891), .B(n27890), .Z(n27893) );
  ANDN U28338 ( .B(n27893), .A(n27892), .Z(n27894) );
  OR U28339 ( .A(n27895), .B(n27894), .Z(n27896) );
  NANDN U28340 ( .A(n27897), .B(n27896), .Z(n27898) );
  NANDN U28341 ( .A(n27899), .B(n27898), .Z(n27901) );
  NAND U28342 ( .A(n27901), .B(n27900), .Z(n27903) );
  ANDN U28343 ( .B(n27903), .A(n27902), .Z(n27905) );
  NANDN U28344 ( .A(n27905), .B(n27904), .Z(n27906) );
  NANDN U28345 ( .A(n27907), .B(n27906), .Z(n27909) );
  NAND U28346 ( .A(n27909), .B(n27908), .Z(n27910) );
  AND U28347 ( .A(n27911), .B(n27910), .Z(n27912) );
  NANDN U28348 ( .A(n27913), .B(n27912), .Z(n27915) );
  NAND U28349 ( .A(n27915), .B(n27914), .Z(n27916) );
  NANDN U28350 ( .A(n27917), .B(n27916), .Z(n27919) );
  NAND U28351 ( .A(n27919), .B(n27918), .Z(n27921) );
  NAND U28352 ( .A(n27921), .B(n27920), .Z(n27923) );
  NAND U28353 ( .A(n27923), .B(n27922), .Z(n27925) );
  ANDN U28354 ( .B(n27925), .A(n27924), .Z(n27927) );
  NANDN U28355 ( .A(n27927), .B(n27926), .Z(n27928) );
  NANDN U28356 ( .A(n27929), .B(n27928), .Z(n27930) );
  NANDN U28357 ( .A(n27931), .B(n27930), .Z(n27933) );
  NAND U28358 ( .A(n27933), .B(n27932), .Z(n27934) );
  AND U28359 ( .A(n27935), .B(n27934), .Z(n27939) );
  NOR U28360 ( .A(n27937), .B(n27936), .Z(n27938) );
  NANDN U28361 ( .A(n27939), .B(n27938), .Z(n27941) );
  NAND U28362 ( .A(n27941), .B(n27940), .Z(n27943) );
  ANDN U28363 ( .B(n27943), .A(n27942), .Z(n27945) );
  NANDN U28364 ( .A(n27945), .B(n27944), .Z(n27946) );
  NANDN U28365 ( .A(n27947), .B(n27946), .Z(n27948) );
  NANDN U28366 ( .A(n27949), .B(n27948), .Z(n27951) );
  NAND U28367 ( .A(n27951), .B(n27950), .Z(n27952) );
  AND U28368 ( .A(n27953), .B(n27952), .Z(n27957) );
  NOR U28369 ( .A(n27955), .B(n27954), .Z(n27956) );
  NANDN U28370 ( .A(n27957), .B(n27956), .Z(n27959) );
  NAND U28371 ( .A(n27959), .B(n27958), .Z(n27961) );
  ANDN U28372 ( .B(n27961), .A(n27960), .Z(n27962) );
  OR U28373 ( .A(n27963), .B(n27962), .Z(n27964) );
  NANDN U28374 ( .A(n27965), .B(n27964), .Z(n27967) );
  NAND U28375 ( .A(n27967), .B(n27966), .Z(n27969) );
  ANDN U28376 ( .B(n27969), .A(n27968), .Z(n27970) );
  NANDN U28377 ( .A(n27971), .B(n27970), .Z(n27973) );
  NAND U28378 ( .A(n27973), .B(n27972), .Z(n27974) );
  AND U28379 ( .A(n27975), .B(n27974), .Z(n27976) );
  NANDN U28380 ( .A(n27977), .B(n27976), .Z(n27979) );
  NAND U28381 ( .A(n27979), .B(n27978), .Z(n27981) );
  ANDN U28382 ( .B(n27981), .A(n27980), .Z(n27983) );
  NANDN U28383 ( .A(n27983), .B(n27982), .Z(n27984) );
  NANDN U28384 ( .A(n27985), .B(n27984), .Z(n27987) );
  NAND U28385 ( .A(n27987), .B(n27986), .Z(n27988) );
  NANDN U28386 ( .A(n27989), .B(n27988), .Z(n27991) );
  ANDN U28387 ( .B(n27991), .A(n27990), .Z(n27992) );
  OR U28388 ( .A(n27993), .B(n27992), .Z(n27994) );
  NANDN U28389 ( .A(n27995), .B(n27994), .Z(n27996) );
  NANDN U28390 ( .A(n27997), .B(n27996), .Z(n27998) );
  NANDN U28391 ( .A(n27999), .B(n27998), .Z(n28000) );
  AND U28392 ( .A(n28001), .B(n28000), .Z(n28003) );
  NANDN U28393 ( .A(n28003), .B(n28002), .Z(n28004) );
  NANDN U28394 ( .A(n28005), .B(n28004), .Z(n28007) );
  NAND U28395 ( .A(n28007), .B(n28006), .Z(n28008) );
  NANDN U28396 ( .A(n28009), .B(n28008), .Z(n28011) );
  ANDN U28397 ( .B(n28011), .A(n28010), .Z(n28012) );
  ANDN U28398 ( .B(n28013), .A(n28012), .Z(n28015) );
  NANDN U28399 ( .A(n28015), .B(n28014), .Z(n28019) );
  ANDN U28400 ( .B(n28017), .A(n28016), .Z(n28018) );
  NAND U28401 ( .A(n28019), .B(n28018), .Z(n28021) );
  NAND U28402 ( .A(n28021), .B(n28020), .Z(n28023) );
  NAND U28403 ( .A(n28023), .B(n28022), .Z(n28024) );
  NANDN U28404 ( .A(n28025), .B(n28024), .Z(n28027) );
  NAND U28405 ( .A(n28027), .B(n28026), .Z(n28029) );
  NAND U28406 ( .A(n28029), .B(n28028), .Z(n28030) );
  AND U28407 ( .A(n28031), .B(n28030), .Z(n28033) );
  NANDN U28408 ( .A(n28033), .B(n28032), .Z(n28035) );
  NAND U28409 ( .A(n28035), .B(n28034), .Z(n28037) );
  NAND U28410 ( .A(n28037), .B(n28036), .Z(n28039) );
  NAND U28411 ( .A(n28039), .B(n28038), .Z(n28041) );
  ANDN U28412 ( .B(n28041), .A(n28040), .Z(n28043) );
  NANDN U28413 ( .A(n28043), .B(n28042), .Z(n28044) );
  NANDN U28414 ( .A(n28045), .B(n28044), .Z(n28047) );
  NAND U28415 ( .A(n28047), .B(n28046), .Z(n28048) );
  NANDN U28416 ( .A(n28049), .B(n28048), .Z(n28050) );
  AND U28417 ( .A(n28051), .B(n28050), .Z(n28052) );
  OR U28418 ( .A(n28053), .B(n28052), .Z(n28054) );
  NANDN U28419 ( .A(n28055), .B(n28054), .Z(n28057) );
  NAND U28420 ( .A(n28057), .B(n28056), .Z(n28059) );
  NAND U28421 ( .A(n28059), .B(n28058), .Z(n28061) );
  ANDN U28422 ( .B(n28061), .A(n28060), .Z(n28063) );
  NANDN U28423 ( .A(n28063), .B(n28062), .Z(n28065) );
  NAND U28424 ( .A(n28065), .B(n28064), .Z(n28067) );
  NAND U28425 ( .A(n28067), .B(n28066), .Z(n28069) );
  NANDN U28426 ( .A(n28069), .B(n28068), .Z(n28071) );
  NAND U28427 ( .A(n28071), .B(n28070), .Z(n28073) );
  ANDN U28428 ( .B(n28073), .A(n28072), .Z(n28074) );
  OR U28429 ( .A(n28075), .B(n28074), .Z(n28076) );
  NANDN U28430 ( .A(n28077), .B(n28076), .Z(n28079) );
  NAND U28431 ( .A(n28079), .B(n28078), .Z(n28080) );
  AND U28432 ( .A(n28081), .B(n28080), .Z(n28082) );
  NANDN U28433 ( .A(n28083), .B(n28082), .Z(n28085) );
  NAND U28434 ( .A(n28085), .B(n28084), .Z(n28086) );
  NANDN U28435 ( .A(n28087), .B(n28086), .Z(n28089) );
  NAND U28436 ( .A(n28089), .B(n28088), .Z(n28091) );
  NAND U28437 ( .A(n28091), .B(n28090), .Z(n28093) );
  NAND U28438 ( .A(n28093), .B(n28092), .Z(n28095) );
  ANDN U28439 ( .B(n28095), .A(n28094), .Z(n28097) );
  NANDN U28440 ( .A(n28097), .B(n28096), .Z(n28098) );
  NANDN U28441 ( .A(n28099), .B(n28098), .Z(n28101) );
  NAND U28442 ( .A(n28101), .B(n28100), .Z(n28103) );
  NAND U28443 ( .A(n28103), .B(n28102), .Z(n28105) );
  ANDN U28444 ( .B(n28105), .A(n28104), .Z(n28106) );
  OR U28445 ( .A(n28107), .B(n28106), .Z(n28108) );
  NANDN U28446 ( .A(n28109), .B(n28108), .Z(n28110) );
  NANDN U28447 ( .A(n28111), .B(n28110), .Z(n28112) );
  NANDN U28448 ( .A(n28113), .B(n28112), .Z(n28114) );
  AND U28449 ( .A(n28115), .B(n28114), .Z(n28117) );
  NANDN U28450 ( .A(n28117), .B(n28116), .Z(n28121) );
  ANDN U28451 ( .B(n28119), .A(n28118), .Z(n28120) );
  NAND U28452 ( .A(n28121), .B(n28120), .Z(n28123) );
  NAND U28453 ( .A(n28123), .B(n28122), .Z(n28124) );
  NANDN U28454 ( .A(n28125), .B(n28124), .Z(n28127) );
  NAND U28455 ( .A(n28127), .B(n28126), .Z(n28129) );
  NAND U28456 ( .A(n28129), .B(n28128), .Z(n28131) );
  NAND U28457 ( .A(n28131), .B(n28130), .Z(n28133) );
  ANDN U28458 ( .B(n28133), .A(n28132), .Z(n28135) );
  NANDN U28459 ( .A(n28135), .B(n28134), .Z(n28136) );
  NANDN U28460 ( .A(n28137), .B(n28136), .Z(n28139) );
  NAND U28461 ( .A(n28139), .B(n28138), .Z(n28140) );
  NANDN U28462 ( .A(n28141), .B(n28140), .Z(n28143) );
  ANDN U28463 ( .B(n28143), .A(n28142), .Z(n28145) );
  OR U28464 ( .A(n28145), .B(n28144), .Z(n28146) );
  AND U28465 ( .A(n28147), .B(n28146), .Z(n28149) );
  NANDN U28466 ( .A(n28149), .B(n28148), .Z(n28151) );
  ANDN U28467 ( .B(n28151), .A(n28150), .Z(n28152) );
  OR U28468 ( .A(n28153), .B(n28152), .Z(n28154) );
  NANDN U28469 ( .A(n28155), .B(n28154), .Z(n28157) );
  NAND U28470 ( .A(n28157), .B(n28156), .Z(n28159) );
  NANDN U28471 ( .A(n28159), .B(n28158), .Z(n28161) );
  NAND U28472 ( .A(n28161), .B(n28160), .Z(n28163) );
  ANDN U28473 ( .B(n28163), .A(n28162), .Z(n28165) );
  NANDN U28474 ( .A(n28165), .B(n28164), .Z(n28166) );
  NANDN U28475 ( .A(n28167), .B(n28166), .Z(n28169) );
  NAND U28476 ( .A(n28169), .B(n28168), .Z(n28171) );
  ANDN U28477 ( .B(n28171), .A(n28170), .Z(n28173) );
  NAND U28478 ( .A(n28173), .B(n28172), .Z(n28174) );
  NANDN U28479 ( .A(n28175), .B(n28174), .Z(n28177) );
  ANDN U28480 ( .B(n28177), .A(n28176), .Z(n28179) );
  ANDN U28481 ( .B(n28179), .A(n28178), .Z(n28180) );
  OR U28482 ( .A(n28181), .B(n28180), .Z(n28185) );
  ANDN U28483 ( .B(n28183), .A(n28182), .Z(n28184) );
  NAND U28484 ( .A(n28185), .B(n28184), .Z(n28186) );
  NANDN U28485 ( .A(n28187), .B(n28186), .Z(n28189) );
  ANDN U28486 ( .B(n28189), .A(n28188), .Z(n28190) );
  OR U28487 ( .A(n28191), .B(n28190), .Z(n28192) );
  AND U28488 ( .A(n28193), .B(n28192), .Z(n28194) );
  OR U28489 ( .A(n28195), .B(n28194), .Z(n28196) );
  NANDN U28490 ( .A(n28197), .B(n28196), .Z(n28198) );
  NANDN U28491 ( .A(n28199), .B(n28198), .Z(n28201) );
  AND U28492 ( .A(n28201), .B(n28200), .Z(n28203) );
  NAND U28493 ( .A(n28203), .B(n28202), .Z(n28204) );
  NANDN U28494 ( .A(n28205), .B(n28204), .Z(n28206) );
  NANDN U28495 ( .A(n28207), .B(n28206), .Z(n28209) );
  NAND U28496 ( .A(n28209), .B(n28208), .Z(n28211) );
  NAND U28497 ( .A(n28211), .B(n28210), .Z(n28212) );
  NANDN U28498 ( .A(n28213), .B(n28212), .Z(n28215) );
  ANDN U28499 ( .B(n28215), .A(n28214), .Z(n28217) );
  NANDN U28500 ( .A(n28217), .B(n28216), .Z(n28218) );
  NANDN U28501 ( .A(n28219), .B(n28218), .Z(n28221) );
  NAND U28502 ( .A(n28221), .B(n28220), .Z(n28223) );
  ANDN U28503 ( .B(n28223), .A(n28222), .Z(n28225) );
  OR U28504 ( .A(n28225), .B(n28224), .Z(n28227) );
  NAND U28505 ( .A(n28227), .B(n28226), .Z(n28229) );
  ANDN U28506 ( .B(n28229), .A(n28228), .Z(n28230) );
  OR U28507 ( .A(n28231), .B(n28230), .Z(n28232) );
  NANDN U28508 ( .A(n28233), .B(n28232), .Z(n28234) );
  NANDN U28509 ( .A(n28235), .B(n28234), .Z(n28237) );
  ANDN U28510 ( .B(n28237), .A(n28236), .Z(n28239) );
  OR U28511 ( .A(n28239), .B(n28238), .Z(n28241) );
  NAND U28512 ( .A(n28241), .B(n28240), .Z(n28243) );
  ANDN U28513 ( .B(n28243), .A(n28242), .Z(n28245) );
  AND U28514 ( .A(n28245), .B(n28244), .Z(n28247) );
  NANDN U28515 ( .A(n28247), .B(n28246), .Z(n28249) );
  ANDN U28516 ( .B(n28249), .A(n28248), .Z(n28251) );
  NANDN U28517 ( .A(n28251), .B(n28250), .Z(n28252) );
  NANDN U28518 ( .A(n28253), .B(n28252), .Z(n28255) );
  NAND U28519 ( .A(n28255), .B(n28254), .Z(n28257) );
  ANDN U28520 ( .B(n28257), .A(n28256), .Z(n28259) );
  NANDN U28521 ( .A(n28259), .B(n28258), .Z(n28260) );
  NANDN U28522 ( .A(n28261), .B(n28260), .Z(n28263) );
  NAND U28523 ( .A(n28263), .B(n28262), .Z(n28265) );
  ANDN U28524 ( .B(n28265), .A(n28264), .Z(n28266) );
  NANDN U28525 ( .A(n28267), .B(n28266), .Z(n28269) );
  NAND U28526 ( .A(n28269), .B(n28268), .Z(n28271) );
  ANDN U28527 ( .B(n28271), .A(n28270), .Z(n28273) );
  NANDN U28528 ( .A(n28273), .B(n28272), .Z(n28274) );
  NANDN U28529 ( .A(n28275), .B(n28274), .Z(n28277) );
  NAND U28530 ( .A(n28277), .B(n28276), .Z(n28279) );
  ANDN U28531 ( .B(n28279), .A(n28278), .Z(n28281) );
  NANDN U28532 ( .A(n28281), .B(n28280), .Z(n28283) );
  ANDN U28533 ( .B(n28283), .A(n28282), .Z(n28285) );
  NANDN U28534 ( .A(n28285), .B(n28284), .Z(n28286) );
  NANDN U28535 ( .A(n28287), .B(n28286), .Z(n28289) );
  NAND U28536 ( .A(n28289), .B(n28288), .Z(n28291) );
  ANDN U28537 ( .B(n28291), .A(n28290), .Z(n28293) );
  NANDN U28538 ( .A(n28293), .B(n28292), .Z(n28295) );
  NAND U28539 ( .A(n28295), .B(n28294), .Z(n28296) );
  AND U28540 ( .A(n28297), .B(n28296), .Z(n28299) );
  NANDN U28541 ( .A(n28299), .B(n28298), .Z(n28301) );
  NAND U28542 ( .A(n28301), .B(n28300), .Z(n28303) );
  NAND U28543 ( .A(n28303), .B(n28302), .Z(n28304) );
  AND U28544 ( .A(n28305), .B(n28304), .Z(n28307) );
  NANDN U28545 ( .A(n28307), .B(n28306), .Z(n28309) );
  ANDN U28546 ( .B(n28309), .A(n28308), .Z(n28310) );
  OR U28547 ( .A(n28311), .B(n28310), .Z(n28312) );
  NANDN U28548 ( .A(n28313), .B(n28312), .Z(n28314) );
  NANDN U28549 ( .A(n28315), .B(n28314), .Z(n28317) );
  ANDN U28550 ( .B(n28317), .A(n28316), .Z(n28319) );
  OR U28551 ( .A(n28319), .B(n28318), .Z(n28321) );
  NAND U28552 ( .A(n28321), .B(n28320), .Z(n28323) );
  ANDN U28553 ( .B(n28323), .A(n28322), .Z(n28325) );
  NANDN U28554 ( .A(n28325), .B(n28324), .Z(n28329) );
  NOR U28555 ( .A(n28327), .B(n28326), .Z(n28328) );
  NAND U28556 ( .A(n28329), .B(n28328), .Z(n28331) );
  NAND U28557 ( .A(n28331), .B(n28330), .Z(n28332) );
  AND U28558 ( .A(n28333), .B(n28332), .Z(n28334) );
  OR U28559 ( .A(n28335), .B(n28334), .Z(n28336) );
  AND U28560 ( .A(n28337), .B(n28336), .Z(n28338) );
  OR U28561 ( .A(n28339), .B(n28338), .Z(n28343) );
  NOR U28562 ( .A(n28341), .B(n28340), .Z(n28342) );
  NAND U28563 ( .A(n28343), .B(n28342), .Z(n28345) );
  NAND U28564 ( .A(n28345), .B(n28344), .Z(n28346) );
  AND U28565 ( .A(n28347), .B(n28346), .Z(n28349) );
  NAND U28566 ( .A(n28349), .B(n28348), .Z(n28351) );
  NAND U28567 ( .A(n28351), .B(n28350), .Z(n28353) );
  ANDN U28568 ( .B(n28353), .A(n28352), .Z(n28355) );
  NANDN U28569 ( .A(n28355), .B(n28354), .Z(n28359) );
  AND U28570 ( .A(n28357), .B(n28356), .Z(n28358) );
  NAND U28571 ( .A(n28359), .B(n28358), .Z(n28361) );
  NAND U28572 ( .A(n28361), .B(n28360), .Z(n28363) );
  ANDN U28573 ( .B(n28363), .A(n28362), .Z(n28365) );
  NANDN U28574 ( .A(n28365), .B(n28364), .Z(n28366) );
  AND U28575 ( .A(n28367), .B(n28366), .Z(n28369) );
  NANDN U28576 ( .A(n28369), .B(n28368), .Z(n28373) );
  ANDN U28577 ( .B(n28371), .A(n28370), .Z(n28372) );
  NAND U28578 ( .A(n28373), .B(n28372), .Z(n28374) );
  NANDN U28579 ( .A(n28375), .B(n28374), .Z(n28377) );
  ANDN U28580 ( .B(n28377), .A(n28376), .Z(n28379) );
  NANDN U28581 ( .A(n28379), .B(n28378), .Z(n28380) );
  AND U28582 ( .A(n28381), .B(n28380), .Z(n28383) );
  NANDN U28583 ( .A(n28383), .B(n28382), .Z(n28384) );
  NANDN U28584 ( .A(n28385), .B(n28384), .Z(n28386) );
  NANDN U28585 ( .A(n28387), .B(n28386), .Z(n28389) );
  ANDN U28586 ( .B(n28389), .A(n28388), .Z(n28391) );
  NANDN U28587 ( .A(n28391), .B(n28390), .Z(n28392) );
  AND U28588 ( .A(n28393), .B(n28392), .Z(n28395) );
  NANDN U28589 ( .A(n28395), .B(n28394), .Z(n28396) );
  NANDN U28590 ( .A(n28397), .B(n28396), .Z(n28399) );
  NAND U28591 ( .A(n28399), .B(n28398), .Z(n28401) );
  ANDN U28592 ( .B(n28401), .A(n28400), .Z(n28403) );
  OR U28593 ( .A(n28403), .B(n28402), .Z(n28405) );
  ANDN U28594 ( .B(n28405), .A(n28404), .Z(n28407) );
  NANDN U28595 ( .A(n28407), .B(n28406), .Z(n28411) );
  NOR U28596 ( .A(n28409), .B(n28408), .Z(n28410) );
  NAND U28597 ( .A(n28411), .B(n28410), .Z(n28413) );
  NAND U28598 ( .A(n28413), .B(n28412), .Z(n28415) );
  ANDN U28599 ( .B(n28415), .A(n28414), .Z(n28417) );
  OR U28600 ( .A(n28417), .B(n28416), .Z(n28418) );
  AND U28601 ( .A(n28419), .B(n28418), .Z(n28420) );
  OR U28602 ( .A(n28421), .B(n28420), .Z(n28422) );
  NANDN U28603 ( .A(n28423), .B(n28422), .Z(n28424) );
  NANDN U28604 ( .A(n28425), .B(n28424), .Z(n28427) );
  ANDN U28605 ( .B(n28427), .A(n28426), .Z(n28429) );
  OR U28606 ( .A(n28429), .B(n28428), .Z(n28431) );
  ANDN U28607 ( .B(n28431), .A(n28430), .Z(n28432) );
  OR U28608 ( .A(n28433), .B(n28432), .Z(n28434) );
  NANDN U28609 ( .A(n28435), .B(n28434), .Z(n28436) );
  NANDN U28610 ( .A(n28437), .B(n28436), .Z(n28439) );
  ANDN U28611 ( .B(n28439), .A(n28438), .Z(n28440) );
  OR U28612 ( .A(n28441), .B(n28440), .Z(n28442) );
  NANDN U28613 ( .A(n28443), .B(n28442), .Z(n28444) );
  NANDN U28614 ( .A(n28445), .B(n28444), .Z(n28446) );
  AND U28615 ( .A(n28447), .B(n28446), .Z(n28449) );
  NAND U28616 ( .A(n28449), .B(n28448), .Z(n28450) );
  NANDN U28617 ( .A(n28451), .B(n28450), .Z(n28453) );
  ANDN U28618 ( .B(n28453), .A(n28452), .Z(n28455) );
  NANDN U28619 ( .A(n28455), .B(n28454), .Z(n28459) );
  ANDN U28620 ( .B(n28457), .A(n28456), .Z(n28458) );
  NAND U28621 ( .A(n28459), .B(n28458), .Z(n28461) );
  NAND U28622 ( .A(n28461), .B(n28460), .Z(n28463) );
  ANDN U28623 ( .B(n28463), .A(n28462), .Z(n28464) );
  AND U28624 ( .A(n28465), .B(n28464), .Z(n28467) );
  OR U28625 ( .A(n28467), .B(n28466), .Z(n28469) );
  ANDN U28626 ( .B(n28469), .A(n28468), .Z(n28471) );
  ANDN U28627 ( .B(n28471), .A(n28470), .Z(n28473) );
  OR U28628 ( .A(n28473), .B(n28472), .Z(n28475) );
  ANDN U28629 ( .B(n28475), .A(n28474), .Z(n28476) );
  OR U28630 ( .A(n28477), .B(n28476), .Z(n28481) );
  AND U28631 ( .A(n28479), .B(n28478), .Z(n28480) );
  NAND U28632 ( .A(n28481), .B(n28480), .Z(n28482) );
  NANDN U28633 ( .A(n28483), .B(n28482), .Z(n28485) );
  ANDN U28634 ( .B(n28485), .A(n28484), .Z(n28487) );
  ANDN U28635 ( .B(n28487), .A(n28486), .Z(n28489) );
  OR U28636 ( .A(n28489), .B(n28488), .Z(n28491) );
  ANDN U28637 ( .B(n28491), .A(n28490), .Z(n28492) );
  OR U28638 ( .A(n28493), .B(n28492), .Z(n28494) );
  NANDN U28639 ( .A(n28495), .B(n28494), .Z(n28497) );
  NAND U28640 ( .A(n28497), .B(n28496), .Z(n28498) );
  AND U28641 ( .A(n28499), .B(n28498), .Z(n28501) );
  NANDN U28642 ( .A(n28501), .B(n28500), .Z(n28502) );
  AND U28643 ( .A(n28503), .B(n28502), .Z(n28505) );
  NANDN U28644 ( .A(n28505), .B(n28504), .Z(n28509) );
  NOR U28645 ( .A(n28507), .B(n28506), .Z(n28508) );
  NAND U28646 ( .A(n28509), .B(n28508), .Z(n28511) );
  NAND U28647 ( .A(n28511), .B(n28510), .Z(n28512) );
  AND U28648 ( .A(n28513), .B(n28512), .Z(n28515) );
  ANDN U28649 ( .B(n28515), .A(n28514), .Z(n28517) );
  NANDN U28650 ( .A(n28517), .B(n28516), .Z(n28518) );
  AND U28651 ( .A(n28519), .B(n28518), .Z(n28521) );
  NANDN U28652 ( .A(n28521), .B(n28520), .Z(n28523) );
  NAND U28653 ( .A(n28523), .B(n28522), .Z(n28525) );
  NAND U28654 ( .A(n28525), .B(n28524), .Z(n28526) );
  AND U28655 ( .A(n28527), .B(n28526), .Z(n28529) );
  NANDN U28656 ( .A(n28529), .B(n28528), .Z(n28531) );
  ANDN U28657 ( .B(n28531), .A(n28530), .Z(n28532) );
  OR U28658 ( .A(n28533), .B(n28532), .Z(n28537) );
  AND U28659 ( .A(n28535), .B(n28534), .Z(n28536) );
  NAND U28660 ( .A(n28537), .B(n28536), .Z(n28538) );
  NANDN U28661 ( .A(n28539), .B(n28538), .Z(n28541) );
  ANDN U28662 ( .B(n28541), .A(n28540), .Z(n28543) );
  NANDN U28663 ( .A(n28543), .B(n28542), .Z(n28545) );
  ANDN U28664 ( .B(n28545), .A(n28544), .Z(n28546) );
  OR U28665 ( .A(n28547), .B(n28546), .Z(n28548) );
  NANDN U28666 ( .A(n28549), .B(n28548), .Z(n28551) );
  NAND U28667 ( .A(n28551), .B(n28550), .Z(n28553) );
  ANDN U28668 ( .B(n28553), .A(n28552), .Z(n28555) );
  NANDN U28669 ( .A(n28555), .B(n28554), .Z(n28557) );
  NAND U28670 ( .A(n28557), .B(n28556), .Z(n28559) );
  ANDN U28671 ( .B(n28559), .A(n28558), .Z(n28560) );
  OR U28672 ( .A(n28561), .B(n28560), .Z(n28562) );
  NANDN U28673 ( .A(n28563), .B(n28562), .Z(n28564) );
  NANDN U28674 ( .A(n28565), .B(n28564), .Z(n28567) );
  ANDN U28675 ( .B(n28567), .A(n28566), .Z(n28569) );
  OR U28676 ( .A(n28569), .B(n28568), .Z(n28571) );
  ANDN U28677 ( .B(n28571), .A(n28570), .Z(n28572) );
  OR U28678 ( .A(n28573), .B(n28572), .Z(n28574) );
  NANDN U28679 ( .A(n28575), .B(n28574), .Z(n28576) );
  NANDN U28680 ( .A(n28577), .B(n28576), .Z(n28579) );
  ANDN U28681 ( .B(n28579), .A(n28578), .Z(n28580) );
  OR U28682 ( .A(n28581), .B(n28580), .Z(n28583) );
  NAND U28683 ( .A(n28583), .B(n28582), .Z(n28585) );
  NAND U28684 ( .A(n28585), .B(n28584), .Z(n28586) );
  AND U28685 ( .A(n28587), .B(n28586), .Z(n28589) );
  NANDN U28686 ( .A(n28589), .B(n28588), .Z(n28591) );
  NAND U28687 ( .A(n28591), .B(n28590), .Z(n28593) );
  NAND U28688 ( .A(n28593), .B(n28592), .Z(n28595) );
  ANDN U28689 ( .B(n28595), .A(n28594), .Z(n28596) );
  OR U28690 ( .A(n28597), .B(n28596), .Z(n28598) );
  NANDN U28691 ( .A(n28599), .B(n28598), .Z(n28601) );
  ANDN U28692 ( .B(n28601), .A(n28600), .Z(n28602) );
  OR U28693 ( .A(n28603), .B(n28602), .Z(n28604) );
  NANDN U28694 ( .A(n28605), .B(n28604), .Z(n28607) );
  NAND U28695 ( .A(n28607), .B(n28606), .Z(n28608) );
  AND U28696 ( .A(n28609), .B(n28608), .Z(n28611) );
  NANDN U28697 ( .A(n28611), .B(n28610), .Z(n28612) );
  AND U28698 ( .A(n28613), .B(n28612), .Z(n28615) );
  NANDN U28699 ( .A(n28615), .B(n28614), .Z(n28616) );
  NANDN U28700 ( .A(n28617), .B(n28616), .Z(n28619) );
  NAND U28701 ( .A(n28619), .B(n28618), .Z(n28621) );
  ANDN U28702 ( .B(n28621), .A(n28620), .Z(n28622) );
  AND U28703 ( .A(n28623), .B(n28622), .Z(n28625) );
  NANDN U28704 ( .A(n28625), .B(n28624), .Z(n28626) );
  NANDN U28705 ( .A(n28627), .B(n28626), .Z(n28628) );
  NANDN U28706 ( .A(n28629), .B(n28628), .Z(n28631) );
  ANDN U28707 ( .B(n28631), .A(n28630), .Z(n28633) );
  AND U28708 ( .A(n28633), .B(n28632), .Z(n28635) );
  NANDN U28709 ( .A(n28635), .B(n28634), .Z(n28636) );
  NANDN U28710 ( .A(n28637), .B(n28636), .Z(n28639) );
  NAND U28711 ( .A(n28639), .B(n28638), .Z(n28641) );
  ANDN U28712 ( .B(n28641), .A(n28640), .Z(n28643) );
  NANDN U28713 ( .A(n28643), .B(n28642), .Z(n28644) );
  NANDN U28714 ( .A(n28645), .B(n28644), .Z(n28646) );
  NANDN U28715 ( .A(n28647), .B(n28646), .Z(n28649) );
  ANDN U28716 ( .B(n28649), .A(n28648), .Z(n28650) );
  AND U28717 ( .A(n28651), .B(n28650), .Z(n28653) );
  NANDN U28718 ( .A(n28653), .B(n28652), .Z(n28655) );
  ANDN U28719 ( .B(n28655), .A(n28654), .Z(n28656) );
  AND U28720 ( .A(n28657), .B(n28656), .Z(n28659) );
  NANDN U28721 ( .A(n28659), .B(n28658), .Z(n28661) );
  ANDN U28722 ( .B(n28661), .A(n28660), .Z(n28663) );
  NANDN U28723 ( .A(n28663), .B(n28662), .Z(n28664) );
  NANDN U28724 ( .A(n28665), .B(n28664), .Z(n28667) );
  NAND U28725 ( .A(n28667), .B(n28666), .Z(n28669) );
  ANDN U28726 ( .B(n28669), .A(n28668), .Z(n28671) );
  NANDN U28727 ( .A(n28671), .B(n28670), .Z(n28673) );
  NAND U28728 ( .A(n28673), .B(n28672), .Z(n28674) );
  AND U28729 ( .A(n28675), .B(n28674), .Z(n28677) );
  NANDN U28730 ( .A(n28677), .B(n28676), .Z(n28678) );
  NANDN U28731 ( .A(n28679), .B(n28678), .Z(n28681) );
  NAND U28732 ( .A(n28681), .B(n28680), .Z(n28683) );
  NAND U28733 ( .A(n28683), .B(n28682), .Z(n28684) );
  NAND U28734 ( .A(n28685), .B(n28684), .Z(n28686) );
  NANDN U28735 ( .A(n28687), .B(n28686), .Z(n28688) );
  AND U28736 ( .A(n28689), .B(n28688), .Z(n28691) );
  ANDN U28737 ( .B(n28691), .A(n28690), .Z(n28692) );
  ANDN U28738 ( .B(n28693), .A(n28692), .Z(n28695) );
  NANDN U28739 ( .A(n28695), .B(n28694), .Z(n28697) );
  NAND U28740 ( .A(n28697), .B(n28696), .Z(n28699) );
  NAND U28741 ( .A(n28699), .B(n28698), .Z(n28700) );
  AND U28742 ( .A(n28701), .B(n28700), .Z(n28703) );
  NANDN U28743 ( .A(n28703), .B(n28702), .Z(n28704) );
  AND U28744 ( .A(n28705), .B(n28704), .Z(n28707) );
  NANDN U28745 ( .A(n28707), .B(n28706), .Z(n28708) );
  NANDN U28746 ( .A(n28709), .B(n28708), .Z(n28711) );
  NAND U28747 ( .A(n28711), .B(n28710), .Z(n28713) );
  NAND U28748 ( .A(n28713), .B(n28712), .Z(n28715) );
  ANDN U28749 ( .B(n28715), .A(n28714), .Z(n28717) );
  NAND U28750 ( .A(n28717), .B(n28716), .Z(n28718) );
  AND U28751 ( .A(n28719), .B(n28718), .Z(n28721) );
  NANDN U28752 ( .A(n28721), .B(n28720), .Z(n28722) );
  NANDN U28753 ( .A(n28723), .B(n28722), .Z(n28725) );
  NAND U28754 ( .A(n28725), .B(n28724), .Z(n28727) );
  ANDN U28755 ( .B(n28727), .A(n28726), .Z(n28728) );
  OR U28756 ( .A(n28729), .B(n28728), .Z(n28730) );
  NANDN U28757 ( .A(n28731), .B(n28730), .Z(n28732) );
  AND U28758 ( .A(n28733), .B(n28732), .Z(n28735) );
  ANDN U28759 ( .B(n28735), .A(n28734), .Z(n28737) );
  OR U28760 ( .A(n28737), .B(n28736), .Z(n28739) );
  ANDN U28761 ( .B(n28739), .A(n28738), .Z(n28740) );
  OR U28762 ( .A(n28741), .B(n28740), .Z(n28742) );
  NANDN U28763 ( .A(n28743), .B(n28742), .Z(n28744) );
  NANDN U28764 ( .A(n28745), .B(n28744), .Z(n28747) );
  ANDN U28765 ( .B(n28747), .A(n28746), .Z(n28748) );
  OR U28766 ( .A(n28749), .B(n28748), .Z(n28750) );
  NAND U28767 ( .A(n28751), .B(n28750), .Z(n28752) );
  NANDN U28768 ( .A(n28753), .B(n28752), .Z(n28754) );
  NAND U28769 ( .A(n28755), .B(n28754), .Z(n28757) );
  ANDN U28770 ( .B(n28757), .A(n28756), .Z(n28758) );
  OR U28771 ( .A(n28759), .B(n28758), .Z(n28763) );
  AND U28772 ( .A(n28761), .B(n28760), .Z(n28762) );
  NAND U28773 ( .A(n28763), .B(n28762), .Z(n28764) );
  NANDN U28774 ( .A(n28765), .B(n28764), .Z(n28767) );
  ANDN U28775 ( .B(n28767), .A(n28766), .Z(n28768) );
  OR U28776 ( .A(n28769), .B(n28768), .Z(n28771) );
  NAND U28777 ( .A(n28771), .B(n28770), .Z(n28772) );
  AND U28778 ( .A(n28773), .B(n28772), .Z(n4) );
endmodule

