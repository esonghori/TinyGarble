
module sum_N256_CC1 ( clk, rst, a, b, c );
  input [255:0] a;
  input [255:0] b;
  output [255:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018;

  XNOR U2 ( .A(a[2]), .B(n1014), .Z(n78) );
  XNOR U3 ( .A(a[5]), .B(n1005), .Z(n45) );
  XNOR U4 ( .A(a[8]), .B(n996), .Z(n12) );
  XNOR U5 ( .A(a[11]), .B(n987), .Z(n644) );
  XNOR U6 ( .A(a[14]), .B(n978), .Z(n521) );
  XNOR U7 ( .A(a[17]), .B(n969), .Z(n398) );
  XNOR U8 ( .A(a[20]), .B(n960), .Z(n274) );
  XNOR U9 ( .A(a[23]), .B(n951), .Z(n151) );
  XNOR U10 ( .A(a[26]), .B(n942), .Z(n82) );
  XNOR U11 ( .A(a[29]), .B(n933), .Z(n79) );
  XNOR U12 ( .A(a[32]), .B(n924), .Z(n75) );
  XNOR U13 ( .A(a[35]), .B(n915), .Z(n72) );
  XNOR U14 ( .A(a[38]), .B(n906), .Z(n69) );
  XNOR U15 ( .A(a[41]), .B(n897), .Z(n65) );
  XNOR U16 ( .A(a[44]), .B(n888), .Z(n62) );
  XNOR U17 ( .A(a[47]), .B(n879), .Z(n59) );
  XNOR U18 ( .A(a[50]), .B(n870), .Z(n55) );
  XNOR U19 ( .A(a[53]), .B(n861), .Z(n52) );
  XNOR U20 ( .A(a[56]), .B(n852), .Z(n49) );
  XNOR U21 ( .A(a[59]), .B(n843), .Z(n46) );
  XNOR U22 ( .A(a[62]), .B(n834), .Z(n42) );
  XNOR U23 ( .A(a[65]), .B(n825), .Z(n39) );
  XNOR U24 ( .A(a[68]), .B(n816), .Z(n36) );
  XNOR U25 ( .A(a[71]), .B(n807), .Z(n32) );
  XNOR U26 ( .A(a[74]), .B(n798), .Z(n29) );
  XNOR U27 ( .A(a[77]), .B(n789), .Z(n26) );
  XNOR U28 ( .A(a[80]), .B(n780), .Z(n22) );
  XNOR U29 ( .A(a[83]), .B(n771), .Z(n19) );
  XNOR U30 ( .A(a[86]), .B(n762), .Z(n16) );
  XNOR U31 ( .A(a[89]), .B(n753), .Z(n13) );
  XNOR U32 ( .A(a[92]), .B(n744), .Z(n9) );
  XNOR U33 ( .A(a[95]), .B(n735), .Z(n6) );
  XNOR U34 ( .A(a[98]), .B(n726), .Z(n3) );
  XNOR U35 ( .A(a[101]), .B(n715), .Z(n717) );
  XNOR U36 ( .A(a[104]), .B(n703), .Z(n705) );
  XNOR U37 ( .A(a[107]), .B(n691), .Z(n693) );
  XNOR U38 ( .A(a[110]), .B(n678), .Z(n680) );
  XNOR U39 ( .A(a[113]), .B(n666), .Z(n668) );
  XNOR U40 ( .A(a[116]), .B(n654), .Z(n656) );
  XNOR U41 ( .A(a[119]), .B(n641), .Z(n643) );
  XNOR U42 ( .A(a[122]), .B(n629), .Z(n631) );
  XNOR U43 ( .A(a[125]), .B(n617), .Z(n619) );
  XNOR U44 ( .A(a[128]), .B(n605), .Z(n607) );
  XNOR U45 ( .A(a[131]), .B(n592), .Z(n594) );
  XNOR U46 ( .A(a[134]), .B(n580), .Z(n582) );
  XNOR U47 ( .A(a[137]), .B(n568), .Z(n570) );
  XNOR U48 ( .A(a[140]), .B(n555), .Z(n557) );
  XNOR U49 ( .A(a[143]), .B(n543), .Z(n545) );
  XNOR U50 ( .A(a[146]), .B(n531), .Z(n533) );
  XNOR U51 ( .A(a[149]), .B(n518), .Z(n520) );
  XNOR U52 ( .A(a[152]), .B(n506), .Z(n508) );
  XNOR U53 ( .A(a[155]), .B(n494), .Z(n496) );
  XNOR U54 ( .A(a[158]), .B(n482), .Z(n484) );
  XNOR U55 ( .A(a[161]), .B(n469), .Z(n471) );
  XNOR U56 ( .A(a[164]), .B(n457), .Z(n459) );
  XNOR U57 ( .A(a[167]), .B(n445), .Z(n447) );
  XNOR U58 ( .A(a[170]), .B(n432), .Z(n434) );
  XNOR U59 ( .A(a[173]), .B(n420), .Z(n422) );
  XNOR U60 ( .A(a[176]), .B(n408), .Z(n410) );
  XNOR U61 ( .A(a[179]), .B(n395), .Z(n397) );
  XNOR U62 ( .A(a[182]), .B(n383), .Z(n385) );
  XNOR U63 ( .A(a[185]), .B(n371), .Z(n373) );
  XNOR U64 ( .A(a[188]), .B(n359), .Z(n361) );
  XNOR U65 ( .A(a[191]), .B(n346), .Z(n348) );
  XNOR U66 ( .A(a[194]), .B(n334), .Z(n336) );
  XNOR U67 ( .A(a[197]), .B(n322), .Z(n324) );
  XNOR U68 ( .A(a[200]), .B(n308), .Z(n310) );
  XNOR U69 ( .A(a[203]), .B(n296), .Z(n298) );
  XNOR U70 ( .A(a[206]), .B(n284), .Z(n286) );
  XNOR U71 ( .A(a[209]), .B(n271), .Z(n273) );
  XNOR U72 ( .A(a[212]), .B(n259), .Z(n261) );
  XNOR U73 ( .A(a[215]), .B(n247), .Z(n249) );
  XNOR U74 ( .A(a[218]), .B(n235), .Z(n237) );
  XNOR U75 ( .A(a[221]), .B(n222), .Z(n224) );
  XNOR U76 ( .A(a[224]), .B(n210), .Z(n212) );
  XNOR U77 ( .A(a[227]), .B(n198), .Z(n200) );
  XNOR U78 ( .A(a[230]), .B(n185), .Z(n187) );
  XNOR U79 ( .A(a[233]), .B(n173), .Z(n175) );
  XNOR U80 ( .A(a[236]), .B(n161), .Z(n163) );
  XNOR U81 ( .A(a[239]), .B(n148), .Z(n150) );
  XNOR U82 ( .A(a[242]), .B(n136), .Z(n138) );
  XNOR U83 ( .A(a[245]), .B(n124), .Z(n126) );
  XNOR U84 ( .A(a[248]), .B(n112), .Z(n114) );
  XNOR U85 ( .A(a[251]), .B(n99), .Z(n101) );
  XNOR U86 ( .A(a[3]), .B(n1011), .Z(n67) );
  XNOR U87 ( .A(a[6]), .B(n1002), .Z(n34) );
  XNOR U88 ( .A(a[9]), .B(n993), .Z(n1) );
  XNOR U89 ( .A(a[12]), .B(n984), .Z(n603) );
  XNOR U90 ( .A(a[15]), .B(n975), .Z(n480) );
  XNOR U91 ( .A(a[18]), .B(n966), .Z(n357) );
  XNOR U92 ( .A(a[21]), .B(n957), .Z(n233) );
  XNOR U93 ( .A(a[24]), .B(n948), .Z(n110) );
  XNOR U94 ( .A(a[27]), .B(n939), .Z(n81) );
  XNOR U95 ( .A(a[30]), .B(n930), .Z(n77) );
  XNOR U96 ( .A(a[33]), .B(n921), .Z(n74) );
  XNOR U97 ( .A(a[36]), .B(n912), .Z(n71) );
  XNOR U98 ( .A(a[39]), .B(n903), .Z(n68) );
  XNOR U99 ( .A(a[42]), .B(n894), .Z(n64) );
  XNOR U100 ( .A(a[45]), .B(n885), .Z(n61) );
  XNOR U101 ( .A(a[48]), .B(n876), .Z(n58) );
  XNOR U102 ( .A(a[51]), .B(n867), .Z(n54) );
  XNOR U103 ( .A(a[54]), .B(n858), .Z(n51) );
  XNOR U104 ( .A(a[57]), .B(n849), .Z(n48) );
  XNOR U105 ( .A(a[60]), .B(n840), .Z(n44) );
  XNOR U106 ( .A(a[63]), .B(n831), .Z(n41) );
  XNOR U107 ( .A(a[66]), .B(n822), .Z(n38) );
  XNOR U108 ( .A(a[69]), .B(n813), .Z(n35) );
  XNOR U109 ( .A(a[72]), .B(n804), .Z(n31) );
  XNOR U110 ( .A(a[75]), .B(n795), .Z(n28) );
  XNOR U111 ( .A(a[78]), .B(n786), .Z(n25) );
  XNOR U112 ( .A(a[81]), .B(n777), .Z(n21) );
  XNOR U113 ( .A(a[84]), .B(n768), .Z(n18) );
  XNOR U114 ( .A(a[87]), .B(n759), .Z(n15) );
  XNOR U115 ( .A(a[90]), .B(n750), .Z(n11) );
  XNOR U116 ( .A(a[93]), .B(n741), .Z(n8) );
  XNOR U117 ( .A(a[96]), .B(n732), .Z(n5) );
  XNOR U118 ( .A(a[99]), .B(n723), .Z(n2) );
  XNOR U119 ( .A(a[102]), .B(n711), .Z(n713) );
  XNOR U120 ( .A(a[105]), .B(n699), .Z(n701) );
  XNOR U121 ( .A(a[108]), .B(n687), .Z(n689) );
  XNOR U122 ( .A(a[111]), .B(n674), .Z(n676) );
  XNOR U123 ( .A(a[114]), .B(n662), .Z(n664) );
  XNOR U124 ( .A(a[117]), .B(n650), .Z(n652) );
  XNOR U125 ( .A(a[120]), .B(n637), .Z(n639) );
  XNOR U126 ( .A(a[123]), .B(n625), .Z(n627) );
  XNOR U127 ( .A(a[126]), .B(n613), .Z(n615) );
  XNOR U128 ( .A(a[129]), .B(n600), .Z(n602) );
  XNOR U129 ( .A(a[132]), .B(n588), .Z(n590) );
  XNOR U130 ( .A(a[135]), .B(n576), .Z(n578) );
  XNOR U131 ( .A(a[138]), .B(n564), .Z(n566) );
  XNOR U132 ( .A(a[141]), .B(n551), .Z(n553) );
  XNOR U133 ( .A(a[144]), .B(n539), .Z(n541) );
  XNOR U134 ( .A(a[147]), .B(n527), .Z(n529) );
  XNOR U135 ( .A(a[150]), .B(n514), .Z(n516) );
  XNOR U136 ( .A(a[153]), .B(n502), .Z(n504) );
  XNOR U137 ( .A(a[156]), .B(n490), .Z(n492) );
  XNOR U138 ( .A(a[159]), .B(n477), .Z(n479) );
  XNOR U139 ( .A(a[162]), .B(n465), .Z(n467) );
  XNOR U140 ( .A(a[165]), .B(n453), .Z(n455) );
  XNOR U141 ( .A(a[168]), .B(n441), .Z(n443) );
  XNOR U142 ( .A(a[171]), .B(n428), .Z(n430) );
  XNOR U143 ( .A(a[174]), .B(n416), .Z(n418) );
  XNOR U144 ( .A(a[177]), .B(n404), .Z(n406) );
  XNOR U145 ( .A(a[180]), .B(n391), .Z(n393) );
  XNOR U146 ( .A(a[183]), .B(n379), .Z(n381) );
  XNOR U147 ( .A(a[186]), .B(n367), .Z(n369) );
  XNOR U148 ( .A(a[189]), .B(n354), .Z(n356) );
  XNOR U149 ( .A(a[192]), .B(n342), .Z(n344) );
  XNOR U150 ( .A(a[195]), .B(n330), .Z(n332) );
  XNOR U151 ( .A(a[198]), .B(n318), .Z(n320) );
  XNOR U152 ( .A(a[201]), .B(n304), .Z(n306) );
  XNOR U153 ( .A(a[204]), .B(n292), .Z(n294) );
  XNOR U154 ( .A(a[207]), .B(n280), .Z(n282) );
  XNOR U155 ( .A(a[210]), .B(n267), .Z(n269) );
  XNOR U156 ( .A(a[213]), .B(n255), .Z(n257) );
  XNOR U157 ( .A(a[216]), .B(n243), .Z(n245) );
  XNOR U158 ( .A(a[219]), .B(n230), .Z(n232) );
  XNOR U159 ( .A(a[222]), .B(n218), .Z(n220) );
  XNOR U160 ( .A(a[225]), .B(n206), .Z(n208) );
  XNOR U161 ( .A(a[228]), .B(n194), .Z(n196) );
  XNOR U162 ( .A(a[231]), .B(n181), .Z(n183) );
  XNOR U163 ( .A(a[234]), .B(n169), .Z(n171) );
  XNOR U164 ( .A(a[237]), .B(n157), .Z(n159) );
  XNOR U165 ( .A(a[240]), .B(n144), .Z(n146) );
  XNOR U166 ( .A(a[243]), .B(n132), .Z(n134) );
  XNOR U167 ( .A(a[246]), .B(n120), .Z(n122) );
  XNOR U168 ( .A(a[249]), .B(n107), .Z(n109) );
  XNOR U169 ( .A(a[252]), .B(n95), .Z(n97) );
  XNOR U170 ( .A(a[4]), .B(n1008), .Z(n56) );
  XNOR U171 ( .A(a[7]), .B(n999), .Z(n23) );
  XNOR U172 ( .A(a[10]), .B(n990), .Z(n685) );
  XNOR U173 ( .A(a[13]), .B(n981), .Z(n562) );
  XNOR U174 ( .A(a[16]), .B(n972), .Z(n439) );
  XNOR U175 ( .A(a[19]), .B(n963), .Z(n316) );
  XNOR U176 ( .A(a[22]), .B(n954), .Z(n192) );
  XNOR U177 ( .A(a[25]), .B(n945), .Z(n83) );
  XNOR U178 ( .A(a[28]), .B(n936), .Z(n80) );
  XNOR U179 ( .A(a[31]), .B(n927), .Z(n76) );
  XNOR U180 ( .A(a[34]), .B(n918), .Z(n73) );
  XNOR U181 ( .A(a[37]), .B(n909), .Z(n70) );
  XNOR U182 ( .A(a[40]), .B(n900), .Z(n66) );
  XNOR U183 ( .A(a[43]), .B(n891), .Z(n63) );
  XNOR U184 ( .A(a[46]), .B(n882), .Z(n60) );
  XNOR U185 ( .A(a[49]), .B(n873), .Z(n57) );
  XNOR U186 ( .A(a[52]), .B(n864), .Z(n53) );
  XNOR U187 ( .A(a[55]), .B(n855), .Z(n50) );
  XNOR U188 ( .A(a[58]), .B(n846), .Z(n47) );
  XNOR U189 ( .A(a[61]), .B(n837), .Z(n43) );
  XNOR U190 ( .A(a[64]), .B(n828), .Z(n40) );
  XNOR U191 ( .A(a[67]), .B(n819), .Z(n37) );
  XNOR U192 ( .A(a[70]), .B(n810), .Z(n33) );
  XNOR U193 ( .A(a[73]), .B(n801), .Z(n30) );
  XNOR U194 ( .A(a[76]), .B(n792), .Z(n27) );
  XNOR U195 ( .A(a[79]), .B(n783), .Z(n24) );
  XNOR U196 ( .A(a[82]), .B(n774), .Z(n20) );
  XNOR U197 ( .A(a[85]), .B(n765), .Z(n17) );
  XNOR U198 ( .A(a[88]), .B(n756), .Z(n14) );
  XNOR U199 ( .A(a[91]), .B(n747), .Z(n10) );
  XNOR U200 ( .A(a[94]), .B(n738), .Z(n7) );
  XNOR U201 ( .A(a[97]), .B(n729), .Z(n4) );
  XNOR U202 ( .A(a[100]), .B(n719), .Z(n721) );
  XNOR U203 ( .A(a[103]), .B(n707), .Z(n709) );
  XNOR U204 ( .A(a[106]), .B(n695), .Z(n697) );
  XNOR U205 ( .A(a[109]), .B(n682), .Z(n684) );
  XNOR U206 ( .A(a[112]), .B(n670), .Z(n672) );
  XNOR U207 ( .A(a[115]), .B(n658), .Z(n660) );
  XNOR U208 ( .A(a[118]), .B(n646), .Z(n648) );
  XNOR U209 ( .A(a[121]), .B(n633), .Z(n635) );
  XNOR U210 ( .A(a[124]), .B(n621), .Z(n623) );
  XNOR U211 ( .A(a[127]), .B(n609), .Z(n611) );
  XNOR U212 ( .A(a[130]), .B(n596), .Z(n598) );
  XNOR U213 ( .A(a[133]), .B(n584), .Z(n586) );
  XNOR U214 ( .A(a[136]), .B(n572), .Z(n574) );
  XNOR U215 ( .A(a[139]), .B(n559), .Z(n561) );
  XNOR U216 ( .A(a[142]), .B(n547), .Z(n549) );
  XNOR U217 ( .A(a[145]), .B(n535), .Z(n537) );
  XNOR U218 ( .A(a[148]), .B(n523), .Z(n525) );
  XNOR U219 ( .A(a[151]), .B(n510), .Z(n512) );
  XNOR U220 ( .A(a[154]), .B(n498), .Z(n500) );
  XNOR U221 ( .A(a[157]), .B(n486), .Z(n488) );
  XNOR U222 ( .A(a[160]), .B(n473), .Z(n475) );
  XNOR U223 ( .A(a[163]), .B(n461), .Z(n463) );
  XNOR U224 ( .A(a[166]), .B(n449), .Z(n451) );
  XNOR U225 ( .A(a[169]), .B(n436), .Z(n438) );
  XNOR U226 ( .A(a[172]), .B(n424), .Z(n426) );
  XNOR U227 ( .A(a[175]), .B(n412), .Z(n414) );
  XNOR U228 ( .A(a[178]), .B(n400), .Z(n402) );
  XNOR U229 ( .A(a[181]), .B(n387), .Z(n389) );
  XNOR U230 ( .A(a[184]), .B(n375), .Z(n377) );
  XNOR U231 ( .A(a[187]), .B(n363), .Z(n365) );
  XNOR U232 ( .A(a[190]), .B(n350), .Z(n352) );
  XNOR U233 ( .A(a[193]), .B(n338), .Z(n340) );
  XNOR U234 ( .A(a[196]), .B(n326), .Z(n328) );
  XNOR U235 ( .A(a[199]), .B(n312), .Z(n314) );
  XNOR U236 ( .A(a[202]), .B(n300), .Z(n302) );
  XNOR U237 ( .A(a[205]), .B(n288), .Z(n290) );
  XNOR U238 ( .A(a[208]), .B(n276), .Z(n278) );
  XNOR U239 ( .A(a[211]), .B(n263), .Z(n265) );
  XNOR U240 ( .A(a[214]), .B(n251), .Z(n253) );
  XNOR U241 ( .A(a[217]), .B(n239), .Z(n241) );
  XNOR U242 ( .A(a[220]), .B(n226), .Z(n228) );
  XNOR U243 ( .A(a[223]), .B(n214), .Z(n216) );
  XNOR U244 ( .A(a[226]), .B(n202), .Z(n204) );
  XNOR U245 ( .A(a[229]), .B(n189), .Z(n191) );
  XNOR U246 ( .A(a[232]), .B(n177), .Z(n179) );
  XNOR U247 ( .A(a[235]), .B(n165), .Z(n167) );
  XNOR U248 ( .A(a[238]), .B(n153), .Z(n155) );
  XNOR U249 ( .A(a[241]), .B(n140), .Z(n142) );
  XNOR U250 ( .A(a[244]), .B(n128), .Z(n130) );
  XNOR U251 ( .A(a[247]), .B(n116), .Z(n118) );
  XNOR U252 ( .A(a[250]), .B(n103), .Z(n105) );
  XNOR U253 ( .A(a[253]), .B(n91), .Z(n93) );
  XNOR U254 ( .A(b[9]), .B(n1), .Z(c[9]) );
  XNOR U255 ( .A(b[99]), .B(n2), .Z(c[99]) );
  XNOR U256 ( .A(b[98]), .B(n3), .Z(c[98]) );
  XNOR U257 ( .A(b[97]), .B(n4), .Z(c[97]) );
  XNOR U258 ( .A(b[96]), .B(n5), .Z(c[96]) );
  XNOR U259 ( .A(b[95]), .B(n6), .Z(c[95]) );
  XNOR U260 ( .A(b[94]), .B(n7), .Z(c[94]) );
  XNOR U261 ( .A(b[93]), .B(n8), .Z(c[93]) );
  XNOR U262 ( .A(b[92]), .B(n9), .Z(c[92]) );
  XNOR U263 ( .A(b[91]), .B(n10), .Z(c[91]) );
  XNOR U264 ( .A(b[90]), .B(n11), .Z(c[90]) );
  XNOR U265 ( .A(b[8]), .B(n12), .Z(c[8]) );
  XNOR U266 ( .A(b[89]), .B(n13), .Z(c[89]) );
  XNOR U267 ( .A(b[88]), .B(n14), .Z(c[88]) );
  XNOR U268 ( .A(b[87]), .B(n15), .Z(c[87]) );
  XNOR U269 ( .A(b[86]), .B(n16), .Z(c[86]) );
  XNOR U270 ( .A(b[85]), .B(n17), .Z(c[85]) );
  XNOR U271 ( .A(b[84]), .B(n18), .Z(c[84]) );
  XNOR U272 ( .A(b[83]), .B(n19), .Z(c[83]) );
  XNOR U273 ( .A(b[82]), .B(n20), .Z(c[82]) );
  XNOR U274 ( .A(b[81]), .B(n21), .Z(c[81]) );
  XNOR U275 ( .A(b[80]), .B(n22), .Z(c[80]) );
  XNOR U276 ( .A(b[7]), .B(n23), .Z(c[7]) );
  XNOR U277 ( .A(b[79]), .B(n24), .Z(c[79]) );
  XNOR U278 ( .A(b[78]), .B(n25), .Z(c[78]) );
  XNOR U279 ( .A(b[77]), .B(n26), .Z(c[77]) );
  XNOR U280 ( .A(b[76]), .B(n27), .Z(c[76]) );
  XNOR U281 ( .A(b[75]), .B(n28), .Z(c[75]) );
  XNOR U282 ( .A(b[74]), .B(n29), .Z(c[74]) );
  XNOR U283 ( .A(b[73]), .B(n30), .Z(c[73]) );
  XNOR U284 ( .A(b[72]), .B(n31), .Z(c[72]) );
  XNOR U285 ( .A(b[71]), .B(n32), .Z(c[71]) );
  XNOR U286 ( .A(b[70]), .B(n33), .Z(c[70]) );
  XNOR U287 ( .A(b[6]), .B(n34), .Z(c[6]) );
  XNOR U288 ( .A(b[69]), .B(n35), .Z(c[69]) );
  XNOR U289 ( .A(b[68]), .B(n36), .Z(c[68]) );
  XNOR U290 ( .A(b[67]), .B(n37), .Z(c[67]) );
  XNOR U291 ( .A(b[66]), .B(n38), .Z(c[66]) );
  XNOR U292 ( .A(b[65]), .B(n39), .Z(c[65]) );
  XNOR U293 ( .A(b[64]), .B(n40), .Z(c[64]) );
  XNOR U294 ( .A(b[63]), .B(n41), .Z(c[63]) );
  XNOR U295 ( .A(b[62]), .B(n42), .Z(c[62]) );
  XNOR U296 ( .A(b[61]), .B(n43), .Z(c[61]) );
  XNOR U297 ( .A(b[60]), .B(n44), .Z(c[60]) );
  XNOR U298 ( .A(b[5]), .B(n45), .Z(c[5]) );
  XNOR U299 ( .A(b[59]), .B(n46), .Z(c[59]) );
  XNOR U300 ( .A(b[58]), .B(n47), .Z(c[58]) );
  XNOR U301 ( .A(b[57]), .B(n48), .Z(c[57]) );
  XNOR U302 ( .A(b[56]), .B(n49), .Z(c[56]) );
  XNOR U303 ( .A(b[55]), .B(n50), .Z(c[55]) );
  XNOR U304 ( .A(b[54]), .B(n51), .Z(c[54]) );
  XNOR U305 ( .A(b[53]), .B(n52), .Z(c[53]) );
  XNOR U306 ( .A(b[52]), .B(n53), .Z(c[52]) );
  XNOR U307 ( .A(b[51]), .B(n54), .Z(c[51]) );
  XNOR U308 ( .A(b[50]), .B(n55), .Z(c[50]) );
  XNOR U309 ( .A(b[4]), .B(n56), .Z(c[4]) );
  XNOR U310 ( .A(b[49]), .B(n57), .Z(c[49]) );
  XNOR U311 ( .A(b[48]), .B(n58), .Z(c[48]) );
  XNOR U312 ( .A(b[47]), .B(n59), .Z(c[47]) );
  XNOR U313 ( .A(b[46]), .B(n60), .Z(c[46]) );
  XNOR U314 ( .A(b[45]), .B(n61), .Z(c[45]) );
  XNOR U315 ( .A(b[44]), .B(n62), .Z(c[44]) );
  XNOR U316 ( .A(b[43]), .B(n63), .Z(c[43]) );
  XNOR U317 ( .A(b[42]), .B(n64), .Z(c[42]) );
  XNOR U318 ( .A(b[41]), .B(n65), .Z(c[41]) );
  XNOR U319 ( .A(b[40]), .B(n66), .Z(c[40]) );
  XNOR U320 ( .A(b[3]), .B(n67), .Z(c[3]) );
  XNOR U321 ( .A(b[39]), .B(n68), .Z(c[39]) );
  XNOR U322 ( .A(b[38]), .B(n69), .Z(c[38]) );
  XNOR U323 ( .A(b[37]), .B(n70), .Z(c[37]) );
  XNOR U324 ( .A(b[36]), .B(n71), .Z(c[36]) );
  XNOR U325 ( .A(b[35]), .B(n72), .Z(c[35]) );
  XNOR U326 ( .A(b[34]), .B(n73), .Z(c[34]) );
  XNOR U327 ( .A(b[33]), .B(n74), .Z(c[33]) );
  XNOR U328 ( .A(b[32]), .B(n75), .Z(c[32]) );
  XNOR U329 ( .A(b[31]), .B(n76), .Z(c[31]) );
  XNOR U330 ( .A(b[30]), .B(n77), .Z(c[30]) );
  XNOR U331 ( .A(b[2]), .B(n78), .Z(c[2]) );
  XNOR U332 ( .A(b[29]), .B(n79), .Z(c[29]) );
  XNOR U333 ( .A(b[28]), .B(n80), .Z(c[28]) );
  XNOR U334 ( .A(b[27]), .B(n81), .Z(c[27]) );
  XNOR U335 ( .A(b[26]), .B(n82), .Z(c[26]) );
  XNOR U336 ( .A(b[25]), .B(n83), .Z(c[25]) );
  XOR U337 ( .A(n84), .B(n85), .Z(c[255]) );
  XOR U338 ( .A(n86), .B(n87), .Z(n85) );
  ANDN U339 ( .B(n88), .A(n89), .Z(n86) );
  XOR U340 ( .A(b[254]), .B(n87), .Z(n88) );
  XOR U341 ( .A(b[255]), .B(a[255]), .Z(n84) );
  XNOR U342 ( .A(b[254]), .B(n89), .Z(c[254]) );
  XNOR U343 ( .A(a[254]), .B(n87), .Z(n89) );
  XOR U344 ( .A(n90), .B(n91), .Z(n87) );
  ANDN U345 ( .B(n92), .A(n93), .Z(n90) );
  XOR U346 ( .A(b[253]), .B(n91), .Z(n92) );
  XNOR U347 ( .A(b[253]), .B(n93), .Z(c[253]) );
  XOR U348 ( .A(n94), .B(n95), .Z(n91) );
  ANDN U349 ( .B(n96), .A(n97), .Z(n94) );
  XOR U350 ( .A(b[252]), .B(n95), .Z(n96) );
  XNOR U351 ( .A(b[252]), .B(n97), .Z(c[252]) );
  XOR U352 ( .A(n98), .B(n99), .Z(n95) );
  ANDN U353 ( .B(n100), .A(n101), .Z(n98) );
  XOR U354 ( .A(b[251]), .B(n99), .Z(n100) );
  XNOR U355 ( .A(b[251]), .B(n101), .Z(c[251]) );
  XOR U356 ( .A(n102), .B(n103), .Z(n99) );
  ANDN U357 ( .B(n104), .A(n105), .Z(n102) );
  XOR U358 ( .A(b[250]), .B(n103), .Z(n104) );
  XNOR U359 ( .A(b[250]), .B(n105), .Z(c[250]) );
  XOR U360 ( .A(n106), .B(n107), .Z(n103) );
  ANDN U361 ( .B(n108), .A(n109), .Z(n106) );
  XOR U362 ( .A(b[249]), .B(n107), .Z(n108) );
  XNOR U363 ( .A(b[24]), .B(n110), .Z(c[24]) );
  XNOR U364 ( .A(b[249]), .B(n109), .Z(c[249]) );
  XOR U365 ( .A(n111), .B(n112), .Z(n107) );
  ANDN U366 ( .B(n113), .A(n114), .Z(n111) );
  XOR U367 ( .A(b[248]), .B(n112), .Z(n113) );
  XNOR U368 ( .A(b[248]), .B(n114), .Z(c[248]) );
  XOR U369 ( .A(n115), .B(n116), .Z(n112) );
  ANDN U370 ( .B(n117), .A(n118), .Z(n115) );
  XOR U371 ( .A(b[247]), .B(n116), .Z(n117) );
  XNOR U372 ( .A(b[247]), .B(n118), .Z(c[247]) );
  XOR U373 ( .A(n119), .B(n120), .Z(n116) );
  ANDN U374 ( .B(n121), .A(n122), .Z(n119) );
  XOR U375 ( .A(b[246]), .B(n120), .Z(n121) );
  XNOR U376 ( .A(b[246]), .B(n122), .Z(c[246]) );
  XOR U377 ( .A(n123), .B(n124), .Z(n120) );
  ANDN U378 ( .B(n125), .A(n126), .Z(n123) );
  XOR U379 ( .A(b[245]), .B(n124), .Z(n125) );
  XNOR U380 ( .A(b[245]), .B(n126), .Z(c[245]) );
  XOR U381 ( .A(n127), .B(n128), .Z(n124) );
  ANDN U382 ( .B(n129), .A(n130), .Z(n127) );
  XOR U383 ( .A(b[244]), .B(n128), .Z(n129) );
  XNOR U384 ( .A(b[244]), .B(n130), .Z(c[244]) );
  XOR U385 ( .A(n131), .B(n132), .Z(n128) );
  ANDN U386 ( .B(n133), .A(n134), .Z(n131) );
  XOR U387 ( .A(b[243]), .B(n132), .Z(n133) );
  XNOR U388 ( .A(b[243]), .B(n134), .Z(c[243]) );
  XOR U389 ( .A(n135), .B(n136), .Z(n132) );
  ANDN U390 ( .B(n137), .A(n138), .Z(n135) );
  XOR U391 ( .A(b[242]), .B(n136), .Z(n137) );
  XNOR U392 ( .A(b[242]), .B(n138), .Z(c[242]) );
  XOR U393 ( .A(n139), .B(n140), .Z(n136) );
  ANDN U394 ( .B(n141), .A(n142), .Z(n139) );
  XOR U395 ( .A(b[241]), .B(n140), .Z(n141) );
  XNOR U396 ( .A(b[241]), .B(n142), .Z(c[241]) );
  XOR U397 ( .A(n143), .B(n144), .Z(n140) );
  ANDN U398 ( .B(n145), .A(n146), .Z(n143) );
  XOR U399 ( .A(b[240]), .B(n144), .Z(n145) );
  XNOR U400 ( .A(b[240]), .B(n146), .Z(c[240]) );
  XOR U401 ( .A(n147), .B(n148), .Z(n144) );
  ANDN U402 ( .B(n149), .A(n150), .Z(n147) );
  XOR U403 ( .A(b[239]), .B(n148), .Z(n149) );
  XNOR U404 ( .A(b[23]), .B(n151), .Z(c[23]) );
  XNOR U405 ( .A(b[239]), .B(n150), .Z(c[239]) );
  XOR U406 ( .A(n152), .B(n153), .Z(n148) );
  ANDN U407 ( .B(n154), .A(n155), .Z(n152) );
  XOR U408 ( .A(b[238]), .B(n153), .Z(n154) );
  XNOR U409 ( .A(b[238]), .B(n155), .Z(c[238]) );
  XOR U410 ( .A(n156), .B(n157), .Z(n153) );
  ANDN U411 ( .B(n158), .A(n159), .Z(n156) );
  XOR U412 ( .A(b[237]), .B(n157), .Z(n158) );
  XNOR U413 ( .A(b[237]), .B(n159), .Z(c[237]) );
  XOR U414 ( .A(n160), .B(n161), .Z(n157) );
  ANDN U415 ( .B(n162), .A(n163), .Z(n160) );
  XOR U416 ( .A(b[236]), .B(n161), .Z(n162) );
  XNOR U417 ( .A(b[236]), .B(n163), .Z(c[236]) );
  XOR U418 ( .A(n164), .B(n165), .Z(n161) );
  ANDN U419 ( .B(n166), .A(n167), .Z(n164) );
  XOR U420 ( .A(b[235]), .B(n165), .Z(n166) );
  XNOR U421 ( .A(b[235]), .B(n167), .Z(c[235]) );
  XOR U422 ( .A(n168), .B(n169), .Z(n165) );
  ANDN U423 ( .B(n170), .A(n171), .Z(n168) );
  XOR U424 ( .A(b[234]), .B(n169), .Z(n170) );
  XNOR U425 ( .A(b[234]), .B(n171), .Z(c[234]) );
  XOR U426 ( .A(n172), .B(n173), .Z(n169) );
  ANDN U427 ( .B(n174), .A(n175), .Z(n172) );
  XOR U428 ( .A(b[233]), .B(n173), .Z(n174) );
  XNOR U429 ( .A(b[233]), .B(n175), .Z(c[233]) );
  XOR U430 ( .A(n176), .B(n177), .Z(n173) );
  ANDN U431 ( .B(n178), .A(n179), .Z(n176) );
  XOR U432 ( .A(b[232]), .B(n177), .Z(n178) );
  XNOR U433 ( .A(b[232]), .B(n179), .Z(c[232]) );
  XOR U434 ( .A(n180), .B(n181), .Z(n177) );
  ANDN U435 ( .B(n182), .A(n183), .Z(n180) );
  XOR U436 ( .A(b[231]), .B(n181), .Z(n182) );
  XNOR U437 ( .A(b[231]), .B(n183), .Z(c[231]) );
  XOR U438 ( .A(n184), .B(n185), .Z(n181) );
  ANDN U439 ( .B(n186), .A(n187), .Z(n184) );
  XOR U440 ( .A(b[230]), .B(n185), .Z(n186) );
  XNOR U441 ( .A(b[230]), .B(n187), .Z(c[230]) );
  XOR U442 ( .A(n188), .B(n189), .Z(n185) );
  ANDN U443 ( .B(n190), .A(n191), .Z(n188) );
  XOR U444 ( .A(b[229]), .B(n189), .Z(n190) );
  XNOR U445 ( .A(b[22]), .B(n192), .Z(c[22]) );
  XNOR U446 ( .A(b[229]), .B(n191), .Z(c[229]) );
  XOR U447 ( .A(n193), .B(n194), .Z(n189) );
  ANDN U448 ( .B(n195), .A(n196), .Z(n193) );
  XOR U449 ( .A(b[228]), .B(n194), .Z(n195) );
  XNOR U450 ( .A(b[228]), .B(n196), .Z(c[228]) );
  XOR U451 ( .A(n197), .B(n198), .Z(n194) );
  ANDN U452 ( .B(n199), .A(n200), .Z(n197) );
  XOR U453 ( .A(b[227]), .B(n198), .Z(n199) );
  XNOR U454 ( .A(b[227]), .B(n200), .Z(c[227]) );
  XOR U455 ( .A(n201), .B(n202), .Z(n198) );
  ANDN U456 ( .B(n203), .A(n204), .Z(n201) );
  XOR U457 ( .A(b[226]), .B(n202), .Z(n203) );
  XNOR U458 ( .A(b[226]), .B(n204), .Z(c[226]) );
  XOR U459 ( .A(n205), .B(n206), .Z(n202) );
  ANDN U460 ( .B(n207), .A(n208), .Z(n205) );
  XOR U461 ( .A(b[225]), .B(n206), .Z(n207) );
  XNOR U462 ( .A(b[225]), .B(n208), .Z(c[225]) );
  XOR U463 ( .A(n209), .B(n210), .Z(n206) );
  ANDN U464 ( .B(n211), .A(n212), .Z(n209) );
  XOR U465 ( .A(b[224]), .B(n210), .Z(n211) );
  XNOR U466 ( .A(b[224]), .B(n212), .Z(c[224]) );
  XOR U467 ( .A(n213), .B(n214), .Z(n210) );
  ANDN U468 ( .B(n215), .A(n216), .Z(n213) );
  XOR U469 ( .A(b[223]), .B(n214), .Z(n215) );
  XNOR U470 ( .A(b[223]), .B(n216), .Z(c[223]) );
  XOR U471 ( .A(n217), .B(n218), .Z(n214) );
  ANDN U472 ( .B(n219), .A(n220), .Z(n217) );
  XOR U473 ( .A(b[222]), .B(n218), .Z(n219) );
  XNOR U474 ( .A(b[222]), .B(n220), .Z(c[222]) );
  XOR U475 ( .A(n221), .B(n222), .Z(n218) );
  ANDN U476 ( .B(n223), .A(n224), .Z(n221) );
  XOR U477 ( .A(b[221]), .B(n222), .Z(n223) );
  XNOR U478 ( .A(b[221]), .B(n224), .Z(c[221]) );
  XOR U479 ( .A(n225), .B(n226), .Z(n222) );
  ANDN U480 ( .B(n227), .A(n228), .Z(n225) );
  XOR U481 ( .A(b[220]), .B(n226), .Z(n227) );
  XNOR U482 ( .A(b[220]), .B(n228), .Z(c[220]) );
  XOR U483 ( .A(n229), .B(n230), .Z(n226) );
  ANDN U484 ( .B(n231), .A(n232), .Z(n229) );
  XOR U485 ( .A(b[219]), .B(n230), .Z(n231) );
  XNOR U486 ( .A(b[21]), .B(n233), .Z(c[21]) );
  XNOR U487 ( .A(b[219]), .B(n232), .Z(c[219]) );
  XOR U488 ( .A(n234), .B(n235), .Z(n230) );
  ANDN U489 ( .B(n236), .A(n237), .Z(n234) );
  XOR U490 ( .A(b[218]), .B(n235), .Z(n236) );
  XNOR U491 ( .A(b[218]), .B(n237), .Z(c[218]) );
  XOR U492 ( .A(n238), .B(n239), .Z(n235) );
  ANDN U493 ( .B(n240), .A(n241), .Z(n238) );
  XOR U494 ( .A(b[217]), .B(n239), .Z(n240) );
  XNOR U495 ( .A(b[217]), .B(n241), .Z(c[217]) );
  XOR U496 ( .A(n242), .B(n243), .Z(n239) );
  ANDN U497 ( .B(n244), .A(n245), .Z(n242) );
  XOR U498 ( .A(b[216]), .B(n243), .Z(n244) );
  XNOR U499 ( .A(b[216]), .B(n245), .Z(c[216]) );
  XOR U500 ( .A(n246), .B(n247), .Z(n243) );
  ANDN U501 ( .B(n248), .A(n249), .Z(n246) );
  XOR U502 ( .A(b[215]), .B(n247), .Z(n248) );
  XNOR U503 ( .A(b[215]), .B(n249), .Z(c[215]) );
  XOR U504 ( .A(n250), .B(n251), .Z(n247) );
  ANDN U505 ( .B(n252), .A(n253), .Z(n250) );
  XOR U506 ( .A(b[214]), .B(n251), .Z(n252) );
  XNOR U507 ( .A(b[214]), .B(n253), .Z(c[214]) );
  XOR U508 ( .A(n254), .B(n255), .Z(n251) );
  ANDN U509 ( .B(n256), .A(n257), .Z(n254) );
  XOR U510 ( .A(b[213]), .B(n255), .Z(n256) );
  XNOR U511 ( .A(b[213]), .B(n257), .Z(c[213]) );
  XOR U512 ( .A(n258), .B(n259), .Z(n255) );
  ANDN U513 ( .B(n260), .A(n261), .Z(n258) );
  XOR U514 ( .A(b[212]), .B(n259), .Z(n260) );
  XNOR U515 ( .A(b[212]), .B(n261), .Z(c[212]) );
  XOR U516 ( .A(n262), .B(n263), .Z(n259) );
  ANDN U517 ( .B(n264), .A(n265), .Z(n262) );
  XOR U518 ( .A(b[211]), .B(n263), .Z(n264) );
  XNOR U519 ( .A(b[211]), .B(n265), .Z(c[211]) );
  XOR U520 ( .A(n266), .B(n267), .Z(n263) );
  ANDN U521 ( .B(n268), .A(n269), .Z(n266) );
  XOR U522 ( .A(b[210]), .B(n267), .Z(n268) );
  XNOR U523 ( .A(b[210]), .B(n269), .Z(c[210]) );
  XOR U524 ( .A(n270), .B(n271), .Z(n267) );
  ANDN U525 ( .B(n272), .A(n273), .Z(n270) );
  XOR U526 ( .A(b[209]), .B(n271), .Z(n272) );
  XNOR U527 ( .A(b[20]), .B(n274), .Z(c[20]) );
  XNOR U528 ( .A(b[209]), .B(n273), .Z(c[209]) );
  XOR U529 ( .A(n275), .B(n276), .Z(n271) );
  ANDN U530 ( .B(n277), .A(n278), .Z(n275) );
  XOR U531 ( .A(b[208]), .B(n276), .Z(n277) );
  XNOR U532 ( .A(b[208]), .B(n278), .Z(c[208]) );
  XOR U533 ( .A(n279), .B(n280), .Z(n276) );
  ANDN U534 ( .B(n281), .A(n282), .Z(n279) );
  XOR U535 ( .A(b[207]), .B(n280), .Z(n281) );
  XNOR U536 ( .A(b[207]), .B(n282), .Z(c[207]) );
  XOR U537 ( .A(n283), .B(n284), .Z(n280) );
  ANDN U538 ( .B(n285), .A(n286), .Z(n283) );
  XOR U539 ( .A(b[206]), .B(n284), .Z(n285) );
  XNOR U540 ( .A(b[206]), .B(n286), .Z(c[206]) );
  XOR U541 ( .A(n287), .B(n288), .Z(n284) );
  ANDN U542 ( .B(n289), .A(n290), .Z(n287) );
  XOR U543 ( .A(b[205]), .B(n288), .Z(n289) );
  XNOR U544 ( .A(b[205]), .B(n290), .Z(c[205]) );
  XOR U545 ( .A(n291), .B(n292), .Z(n288) );
  ANDN U546 ( .B(n293), .A(n294), .Z(n291) );
  XOR U547 ( .A(b[204]), .B(n292), .Z(n293) );
  XNOR U548 ( .A(b[204]), .B(n294), .Z(c[204]) );
  XOR U549 ( .A(n295), .B(n296), .Z(n292) );
  ANDN U550 ( .B(n297), .A(n298), .Z(n295) );
  XOR U551 ( .A(b[203]), .B(n296), .Z(n297) );
  XNOR U552 ( .A(b[203]), .B(n298), .Z(c[203]) );
  XOR U553 ( .A(n299), .B(n300), .Z(n296) );
  ANDN U554 ( .B(n301), .A(n302), .Z(n299) );
  XOR U555 ( .A(b[202]), .B(n300), .Z(n301) );
  XNOR U556 ( .A(b[202]), .B(n302), .Z(c[202]) );
  XOR U557 ( .A(n303), .B(n304), .Z(n300) );
  ANDN U558 ( .B(n305), .A(n306), .Z(n303) );
  XOR U559 ( .A(b[201]), .B(n304), .Z(n305) );
  XNOR U560 ( .A(b[201]), .B(n306), .Z(c[201]) );
  XOR U561 ( .A(n307), .B(n308), .Z(n304) );
  ANDN U562 ( .B(n309), .A(n310), .Z(n307) );
  XOR U563 ( .A(b[200]), .B(n308), .Z(n309) );
  XNOR U564 ( .A(b[200]), .B(n310), .Z(c[200]) );
  XOR U565 ( .A(n311), .B(n312), .Z(n308) );
  ANDN U566 ( .B(n313), .A(n314), .Z(n311) );
  XOR U567 ( .A(b[199]), .B(n312), .Z(n313) );
  XNOR U568 ( .A(b[1]), .B(n315), .Z(c[1]) );
  XNOR U569 ( .A(b[19]), .B(n316), .Z(c[19]) );
  XNOR U570 ( .A(b[199]), .B(n314), .Z(c[199]) );
  XOR U571 ( .A(n317), .B(n318), .Z(n312) );
  ANDN U572 ( .B(n319), .A(n320), .Z(n317) );
  XOR U573 ( .A(b[198]), .B(n318), .Z(n319) );
  XNOR U574 ( .A(b[198]), .B(n320), .Z(c[198]) );
  XOR U575 ( .A(n321), .B(n322), .Z(n318) );
  ANDN U576 ( .B(n323), .A(n324), .Z(n321) );
  XOR U577 ( .A(b[197]), .B(n322), .Z(n323) );
  XNOR U578 ( .A(b[197]), .B(n324), .Z(c[197]) );
  XOR U579 ( .A(n325), .B(n326), .Z(n322) );
  ANDN U580 ( .B(n327), .A(n328), .Z(n325) );
  XOR U581 ( .A(b[196]), .B(n326), .Z(n327) );
  XNOR U582 ( .A(b[196]), .B(n328), .Z(c[196]) );
  XOR U583 ( .A(n329), .B(n330), .Z(n326) );
  ANDN U584 ( .B(n331), .A(n332), .Z(n329) );
  XOR U585 ( .A(b[195]), .B(n330), .Z(n331) );
  XNOR U586 ( .A(b[195]), .B(n332), .Z(c[195]) );
  XOR U587 ( .A(n333), .B(n334), .Z(n330) );
  ANDN U588 ( .B(n335), .A(n336), .Z(n333) );
  XOR U589 ( .A(b[194]), .B(n334), .Z(n335) );
  XNOR U590 ( .A(b[194]), .B(n336), .Z(c[194]) );
  XOR U591 ( .A(n337), .B(n338), .Z(n334) );
  ANDN U592 ( .B(n339), .A(n340), .Z(n337) );
  XOR U593 ( .A(b[193]), .B(n338), .Z(n339) );
  XNOR U594 ( .A(b[193]), .B(n340), .Z(c[193]) );
  XOR U595 ( .A(n341), .B(n342), .Z(n338) );
  ANDN U596 ( .B(n343), .A(n344), .Z(n341) );
  XOR U597 ( .A(b[192]), .B(n342), .Z(n343) );
  XNOR U598 ( .A(b[192]), .B(n344), .Z(c[192]) );
  XOR U599 ( .A(n345), .B(n346), .Z(n342) );
  ANDN U600 ( .B(n347), .A(n348), .Z(n345) );
  XOR U601 ( .A(b[191]), .B(n346), .Z(n347) );
  XNOR U602 ( .A(b[191]), .B(n348), .Z(c[191]) );
  XOR U603 ( .A(n349), .B(n350), .Z(n346) );
  ANDN U604 ( .B(n351), .A(n352), .Z(n349) );
  XOR U605 ( .A(b[190]), .B(n350), .Z(n351) );
  XNOR U606 ( .A(b[190]), .B(n352), .Z(c[190]) );
  XOR U607 ( .A(n353), .B(n354), .Z(n350) );
  ANDN U608 ( .B(n355), .A(n356), .Z(n353) );
  XOR U609 ( .A(b[189]), .B(n354), .Z(n355) );
  XNOR U610 ( .A(b[18]), .B(n357), .Z(c[18]) );
  XNOR U611 ( .A(b[189]), .B(n356), .Z(c[189]) );
  XOR U612 ( .A(n358), .B(n359), .Z(n354) );
  ANDN U613 ( .B(n360), .A(n361), .Z(n358) );
  XOR U614 ( .A(b[188]), .B(n359), .Z(n360) );
  XNOR U615 ( .A(b[188]), .B(n361), .Z(c[188]) );
  XOR U616 ( .A(n362), .B(n363), .Z(n359) );
  ANDN U617 ( .B(n364), .A(n365), .Z(n362) );
  XOR U618 ( .A(b[187]), .B(n363), .Z(n364) );
  XNOR U619 ( .A(b[187]), .B(n365), .Z(c[187]) );
  XOR U620 ( .A(n366), .B(n367), .Z(n363) );
  ANDN U621 ( .B(n368), .A(n369), .Z(n366) );
  XOR U622 ( .A(b[186]), .B(n367), .Z(n368) );
  XNOR U623 ( .A(b[186]), .B(n369), .Z(c[186]) );
  XOR U624 ( .A(n370), .B(n371), .Z(n367) );
  ANDN U625 ( .B(n372), .A(n373), .Z(n370) );
  XOR U626 ( .A(b[185]), .B(n371), .Z(n372) );
  XNOR U627 ( .A(b[185]), .B(n373), .Z(c[185]) );
  XOR U628 ( .A(n374), .B(n375), .Z(n371) );
  ANDN U629 ( .B(n376), .A(n377), .Z(n374) );
  XOR U630 ( .A(b[184]), .B(n375), .Z(n376) );
  XNOR U631 ( .A(b[184]), .B(n377), .Z(c[184]) );
  XOR U632 ( .A(n378), .B(n379), .Z(n375) );
  ANDN U633 ( .B(n380), .A(n381), .Z(n378) );
  XOR U634 ( .A(b[183]), .B(n379), .Z(n380) );
  XNOR U635 ( .A(b[183]), .B(n381), .Z(c[183]) );
  XOR U636 ( .A(n382), .B(n383), .Z(n379) );
  ANDN U637 ( .B(n384), .A(n385), .Z(n382) );
  XOR U638 ( .A(b[182]), .B(n383), .Z(n384) );
  XNOR U639 ( .A(b[182]), .B(n385), .Z(c[182]) );
  XOR U640 ( .A(n386), .B(n387), .Z(n383) );
  ANDN U641 ( .B(n388), .A(n389), .Z(n386) );
  XOR U642 ( .A(b[181]), .B(n387), .Z(n388) );
  XNOR U643 ( .A(b[181]), .B(n389), .Z(c[181]) );
  XOR U644 ( .A(n390), .B(n391), .Z(n387) );
  ANDN U645 ( .B(n392), .A(n393), .Z(n390) );
  XOR U646 ( .A(b[180]), .B(n391), .Z(n392) );
  XNOR U647 ( .A(b[180]), .B(n393), .Z(c[180]) );
  XOR U648 ( .A(n394), .B(n395), .Z(n391) );
  ANDN U649 ( .B(n396), .A(n397), .Z(n394) );
  XOR U650 ( .A(b[179]), .B(n395), .Z(n396) );
  XNOR U651 ( .A(b[17]), .B(n398), .Z(c[17]) );
  XNOR U652 ( .A(b[179]), .B(n397), .Z(c[179]) );
  XOR U653 ( .A(n399), .B(n400), .Z(n395) );
  ANDN U654 ( .B(n401), .A(n402), .Z(n399) );
  XOR U655 ( .A(b[178]), .B(n400), .Z(n401) );
  XNOR U656 ( .A(b[178]), .B(n402), .Z(c[178]) );
  XOR U657 ( .A(n403), .B(n404), .Z(n400) );
  ANDN U658 ( .B(n405), .A(n406), .Z(n403) );
  XOR U659 ( .A(b[177]), .B(n404), .Z(n405) );
  XNOR U660 ( .A(b[177]), .B(n406), .Z(c[177]) );
  XOR U661 ( .A(n407), .B(n408), .Z(n404) );
  ANDN U662 ( .B(n409), .A(n410), .Z(n407) );
  XOR U663 ( .A(b[176]), .B(n408), .Z(n409) );
  XNOR U664 ( .A(b[176]), .B(n410), .Z(c[176]) );
  XOR U665 ( .A(n411), .B(n412), .Z(n408) );
  ANDN U666 ( .B(n413), .A(n414), .Z(n411) );
  XOR U667 ( .A(b[175]), .B(n412), .Z(n413) );
  XNOR U668 ( .A(b[175]), .B(n414), .Z(c[175]) );
  XOR U669 ( .A(n415), .B(n416), .Z(n412) );
  ANDN U670 ( .B(n417), .A(n418), .Z(n415) );
  XOR U671 ( .A(b[174]), .B(n416), .Z(n417) );
  XNOR U672 ( .A(b[174]), .B(n418), .Z(c[174]) );
  XOR U673 ( .A(n419), .B(n420), .Z(n416) );
  ANDN U674 ( .B(n421), .A(n422), .Z(n419) );
  XOR U675 ( .A(b[173]), .B(n420), .Z(n421) );
  XNOR U676 ( .A(b[173]), .B(n422), .Z(c[173]) );
  XOR U677 ( .A(n423), .B(n424), .Z(n420) );
  ANDN U678 ( .B(n425), .A(n426), .Z(n423) );
  XOR U679 ( .A(b[172]), .B(n424), .Z(n425) );
  XNOR U680 ( .A(b[172]), .B(n426), .Z(c[172]) );
  XOR U681 ( .A(n427), .B(n428), .Z(n424) );
  ANDN U682 ( .B(n429), .A(n430), .Z(n427) );
  XOR U683 ( .A(b[171]), .B(n428), .Z(n429) );
  XNOR U684 ( .A(b[171]), .B(n430), .Z(c[171]) );
  XOR U685 ( .A(n431), .B(n432), .Z(n428) );
  ANDN U686 ( .B(n433), .A(n434), .Z(n431) );
  XOR U687 ( .A(b[170]), .B(n432), .Z(n433) );
  XNOR U688 ( .A(b[170]), .B(n434), .Z(c[170]) );
  XOR U689 ( .A(n435), .B(n436), .Z(n432) );
  ANDN U690 ( .B(n437), .A(n438), .Z(n435) );
  XOR U691 ( .A(b[169]), .B(n436), .Z(n437) );
  XNOR U692 ( .A(b[16]), .B(n439), .Z(c[16]) );
  XNOR U693 ( .A(b[169]), .B(n438), .Z(c[169]) );
  XOR U694 ( .A(n440), .B(n441), .Z(n436) );
  ANDN U695 ( .B(n442), .A(n443), .Z(n440) );
  XOR U696 ( .A(b[168]), .B(n441), .Z(n442) );
  XNOR U697 ( .A(b[168]), .B(n443), .Z(c[168]) );
  XOR U698 ( .A(n444), .B(n445), .Z(n441) );
  ANDN U699 ( .B(n446), .A(n447), .Z(n444) );
  XOR U700 ( .A(b[167]), .B(n445), .Z(n446) );
  XNOR U701 ( .A(b[167]), .B(n447), .Z(c[167]) );
  XOR U702 ( .A(n448), .B(n449), .Z(n445) );
  ANDN U703 ( .B(n450), .A(n451), .Z(n448) );
  XOR U704 ( .A(b[166]), .B(n449), .Z(n450) );
  XNOR U705 ( .A(b[166]), .B(n451), .Z(c[166]) );
  XOR U706 ( .A(n452), .B(n453), .Z(n449) );
  ANDN U707 ( .B(n454), .A(n455), .Z(n452) );
  XOR U708 ( .A(b[165]), .B(n453), .Z(n454) );
  XNOR U709 ( .A(b[165]), .B(n455), .Z(c[165]) );
  XOR U710 ( .A(n456), .B(n457), .Z(n453) );
  ANDN U711 ( .B(n458), .A(n459), .Z(n456) );
  XOR U712 ( .A(b[164]), .B(n457), .Z(n458) );
  XNOR U713 ( .A(b[164]), .B(n459), .Z(c[164]) );
  XOR U714 ( .A(n460), .B(n461), .Z(n457) );
  ANDN U715 ( .B(n462), .A(n463), .Z(n460) );
  XOR U716 ( .A(b[163]), .B(n461), .Z(n462) );
  XNOR U717 ( .A(b[163]), .B(n463), .Z(c[163]) );
  XOR U718 ( .A(n464), .B(n465), .Z(n461) );
  ANDN U719 ( .B(n466), .A(n467), .Z(n464) );
  XOR U720 ( .A(b[162]), .B(n465), .Z(n466) );
  XNOR U721 ( .A(b[162]), .B(n467), .Z(c[162]) );
  XOR U722 ( .A(n468), .B(n469), .Z(n465) );
  ANDN U723 ( .B(n470), .A(n471), .Z(n468) );
  XOR U724 ( .A(b[161]), .B(n469), .Z(n470) );
  XNOR U725 ( .A(b[161]), .B(n471), .Z(c[161]) );
  XOR U726 ( .A(n472), .B(n473), .Z(n469) );
  ANDN U727 ( .B(n474), .A(n475), .Z(n472) );
  XOR U728 ( .A(b[160]), .B(n473), .Z(n474) );
  XNOR U729 ( .A(b[160]), .B(n475), .Z(c[160]) );
  XOR U730 ( .A(n476), .B(n477), .Z(n473) );
  ANDN U731 ( .B(n478), .A(n479), .Z(n476) );
  XOR U732 ( .A(b[159]), .B(n477), .Z(n478) );
  XNOR U733 ( .A(b[15]), .B(n480), .Z(c[15]) );
  XNOR U734 ( .A(b[159]), .B(n479), .Z(c[159]) );
  XOR U735 ( .A(n481), .B(n482), .Z(n477) );
  ANDN U736 ( .B(n483), .A(n484), .Z(n481) );
  XOR U737 ( .A(b[158]), .B(n482), .Z(n483) );
  XNOR U738 ( .A(b[158]), .B(n484), .Z(c[158]) );
  XOR U739 ( .A(n485), .B(n486), .Z(n482) );
  ANDN U740 ( .B(n487), .A(n488), .Z(n485) );
  XOR U741 ( .A(b[157]), .B(n486), .Z(n487) );
  XNOR U742 ( .A(b[157]), .B(n488), .Z(c[157]) );
  XOR U743 ( .A(n489), .B(n490), .Z(n486) );
  ANDN U744 ( .B(n491), .A(n492), .Z(n489) );
  XOR U745 ( .A(b[156]), .B(n490), .Z(n491) );
  XNOR U746 ( .A(b[156]), .B(n492), .Z(c[156]) );
  XOR U747 ( .A(n493), .B(n494), .Z(n490) );
  ANDN U748 ( .B(n495), .A(n496), .Z(n493) );
  XOR U749 ( .A(b[155]), .B(n494), .Z(n495) );
  XNOR U750 ( .A(b[155]), .B(n496), .Z(c[155]) );
  XOR U751 ( .A(n497), .B(n498), .Z(n494) );
  ANDN U752 ( .B(n499), .A(n500), .Z(n497) );
  XOR U753 ( .A(b[154]), .B(n498), .Z(n499) );
  XNOR U754 ( .A(b[154]), .B(n500), .Z(c[154]) );
  XOR U755 ( .A(n501), .B(n502), .Z(n498) );
  ANDN U756 ( .B(n503), .A(n504), .Z(n501) );
  XOR U757 ( .A(b[153]), .B(n502), .Z(n503) );
  XNOR U758 ( .A(b[153]), .B(n504), .Z(c[153]) );
  XOR U759 ( .A(n505), .B(n506), .Z(n502) );
  ANDN U760 ( .B(n507), .A(n508), .Z(n505) );
  XOR U761 ( .A(b[152]), .B(n506), .Z(n507) );
  XNOR U762 ( .A(b[152]), .B(n508), .Z(c[152]) );
  XOR U763 ( .A(n509), .B(n510), .Z(n506) );
  ANDN U764 ( .B(n511), .A(n512), .Z(n509) );
  XOR U765 ( .A(b[151]), .B(n510), .Z(n511) );
  XNOR U766 ( .A(b[151]), .B(n512), .Z(c[151]) );
  XOR U767 ( .A(n513), .B(n514), .Z(n510) );
  ANDN U768 ( .B(n515), .A(n516), .Z(n513) );
  XOR U769 ( .A(b[150]), .B(n514), .Z(n515) );
  XNOR U770 ( .A(b[150]), .B(n516), .Z(c[150]) );
  XOR U771 ( .A(n517), .B(n518), .Z(n514) );
  ANDN U772 ( .B(n519), .A(n520), .Z(n517) );
  XOR U773 ( .A(b[149]), .B(n518), .Z(n519) );
  XNOR U774 ( .A(b[14]), .B(n521), .Z(c[14]) );
  XNOR U775 ( .A(b[149]), .B(n520), .Z(c[149]) );
  XOR U776 ( .A(n522), .B(n523), .Z(n518) );
  ANDN U777 ( .B(n524), .A(n525), .Z(n522) );
  XOR U778 ( .A(b[148]), .B(n523), .Z(n524) );
  XNOR U779 ( .A(b[148]), .B(n525), .Z(c[148]) );
  XOR U780 ( .A(n526), .B(n527), .Z(n523) );
  ANDN U781 ( .B(n528), .A(n529), .Z(n526) );
  XOR U782 ( .A(b[147]), .B(n527), .Z(n528) );
  XNOR U783 ( .A(b[147]), .B(n529), .Z(c[147]) );
  XOR U784 ( .A(n530), .B(n531), .Z(n527) );
  ANDN U785 ( .B(n532), .A(n533), .Z(n530) );
  XOR U786 ( .A(b[146]), .B(n531), .Z(n532) );
  XNOR U787 ( .A(b[146]), .B(n533), .Z(c[146]) );
  XOR U788 ( .A(n534), .B(n535), .Z(n531) );
  ANDN U789 ( .B(n536), .A(n537), .Z(n534) );
  XOR U790 ( .A(b[145]), .B(n535), .Z(n536) );
  XNOR U791 ( .A(b[145]), .B(n537), .Z(c[145]) );
  XOR U792 ( .A(n538), .B(n539), .Z(n535) );
  ANDN U793 ( .B(n540), .A(n541), .Z(n538) );
  XOR U794 ( .A(b[144]), .B(n539), .Z(n540) );
  XNOR U795 ( .A(b[144]), .B(n541), .Z(c[144]) );
  XOR U796 ( .A(n542), .B(n543), .Z(n539) );
  ANDN U797 ( .B(n544), .A(n545), .Z(n542) );
  XOR U798 ( .A(b[143]), .B(n543), .Z(n544) );
  XNOR U799 ( .A(b[143]), .B(n545), .Z(c[143]) );
  XOR U800 ( .A(n546), .B(n547), .Z(n543) );
  ANDN U801 ( .B(n548), .A(n549), .Z(n546) );
  XOR U802 ( .A(b[142]), .B(n547), .Z(n548) );
  XNOR U803 ( .A(b[142]), .B(n549), .Z(c[142]) );
  XOR U804 ( .A(n550), .B(n551), .Z(n547) );
  ANDN U805 ( .B(n552), .A(n553), .Z(n550) );
  XOR U806 ( .A(b[141]), .B(n551), .Z(n552) );
  XNOR U807 ( .A(b[141]), .B(n553), .Z(c[141]) );
  XOR U808 ( .A(n554), .B(n555), .Z(n551) );
  ANDN U809 ( .B(n556), .A(n557), .Z(n554) );
  XOR U810 ( .A(b[140]), .B(n555), .Z(n556) );
  XNOR U811 ( .A(b[140]), .B(n557), .Z(c[140]) );
  XOR U812 ( .A(n558), .B(n559), .Z(n555) );
  ANDN U813 ( .B(n560), .A(n561), .Z(n558) );
  XOR U814 ( .A(b[139]), .B(n559), .Z(n560) );
  XNOR U815 ( .A(b[13]), .B(n562), .Z(c[13]) );
  XNOR U816 ( .A(b[139]), .B(n561), .Z(c[139]) );
  XOR U817 ( .A(n563), .B(n564), .Z(n559) );
  ANDN U818 ( .B(n565), .A(n566), .Z(n563) );
  XOR U819 ( .A(b[138]), .B(n564), .Z(n565) );
  XNOR U820 ( .A(b[138]), .B(n566), .Z(c[138]) );
  XOR U821 ( .A(n567), .B(n568), .Z(n564) );
  ANDN U822 ( .B(n569), .A(n570), .Z(n567) );
  XOR U823 ( .A(b[137]), .B(n568), .Z(n569) );
  XNOR U824 ( .A(b[137]), .B(n570), .Z(c[137]) );
  XOR U825 ( .A(n571), .B(n572), .Z(n568) );
  ANDN U826 ( .B(n573), .A(n574), .Z(n571) );
  XOR U827 ( .A(b[136]), .B(n572), .Z(n573) );
  XNOR U828 ( .A(b[136]), .B(n574), .Z(c[136]) );
  XOR U829 ( .A(n575), .B(n576), .Z(n572) );
  ANDN U830 ( .B(n577), .A(n578), .Z(n575) );
  XOR U831 ( .A(b[135]), .B(n576), .Z(n577) );
  XNOR U832 ( .A(b[135]), .B(n578), .Z(c[135]) );
  XOR U833 ( .A(n579), .B(n580), .Z(n576) );
  ANDN U834 ( .B(n581), .A(n582), .Z(n579) );
  XOR U835 ( .A(b[134]), .B(n580), .Z(n581) );
  XNOR U836 ( .A(b[134]), .B(n582), .Z(c[134]) );
  XOR U837 ( .A(n583), .B(n584), .Z(n580) );
  ANDN U838 ( .B(n585), .A(n586), .Z(n583) );
  XOR U839 ( .A(b[133]), .B(n584), .Z(n585) );
  XNOR U840 ( .A(b[133]), .B(n586), .Z(c[133]) );
  XOR U841 ( .A(n587), .B(n588), .Z(n584) );
  ANDN U842 ( .B(n589), .A(n590), .Z(n587) );
  XOR U843 ( .A(b[132]), .B(n588), .Z(n589) );
  XNOR U844 ( .A(b[132]), .B(n590), .Z(c[132]) );
  XOR U845 ( .A(n591), .B(n592), .Z(n588) );
  ANDN U846 ( .B(n593), .A(n594), .Z(n591) );
  XOR U847 ( .A(b[131]), .B(n592), .Z(n593) );
  XNOR U848 ( .A(b[131]), .B(n594), .Z(c[131]) );
  XOR U849 ( .A(n595), .B(n596), .Z(n592) );
  ANDN U850 ( .B(n597), .A(n598), .Z(n595) );
  XOR U851 ( .A(b[130]), .B(n596), .Z(n597) );
  XNOR U852 ( .A(b[130]), .B(n598), .Z(c[130]) );
  XOR U853 ( .A(n599), .B(n600), .Z(n596) );
  ANDN U854 ( .B(n601), .A(n602), .Z(n599) );
  XOR U855 ( .A(b[129]), .B(n600), .Z(n601) );
  XNOR U856 ( .A(b[12]), .B(n603), .Z(c[12]) );
  XNOR U857 ( .A(b[129]), .B(n602), .Z(c[129]) );
  XOR U858 ( .A(n604), .B(n605), .Z(n600) );
  ANDN U859 ( .B(n606), .A(n607), .Z(n604) );
  XOR U860 ( .A(b[128]), .B(n605), .Z(n606) );
  XNOR U861 ( .A(b[128]), .B(n607), .Z(c[128]) );
  XOR U862 ( .A(n608), .B(n609), .Z(n605) );
  ANDN U863 ( .B(n610), .A(n611), .Z(n608) );
  XOR U864 ( .A(b[127]), .B(n609), .Z(n610) );
  XNOR U865 ( .A(b[127]), .B(n611), .Z(c[127]) );
  XOR U866 ( .A(n612), .B(n613), .Z(n609) );
  ANDN U867 ( .B(n614), .A(n615), .Z(n612) );
  XOR U868 ( .A(b[126]), .B(n613), .Z(n614) );
  XNOR U869 ( .A(b[126]), .B(n615), .Z(c[126]) );
  XOR U870 ( .A(n616), .B(n617), .Z(n613) );
  ANDN U871 ( .B(n618), .A(n619), .Z(n616) );
  XOR U872 ( .A(b[125]), .B(n617), .Z(n618) );
  XNOR U873 ( .A(b[125]), .B(n619), .Z(c[125]) );
  XOR U874 ( .A(n620), .B(n621), .Z(n617) );
  ANDN U875 ( .B(n622), .A(n623), .Z(n620) );
  XOR U876 ( .A(b[124]), .B(n621), .Z(n622) );
  XNOR U877 ( .A(b[124]), .B(n623), .Z(c[124]) );
  XOR U878 ( .A(n624), .B(n625), .Z(n621) );
  ANDN U879 ( .B(n626), .A(n627), .Z(n624) );
  XOR U880 ( .A(b[123]), .B(n625), .Z(n626) );
  XNOR U881 ( .A(b[123]), .B(n627), .Z(c[123]) );
  XOR U882 ( .A(n628), .B(n629), .Z(n625) );
  ANDN U883 ( .B(n630), .A(n631), .Z(n628) );
  XOR U884 ( .A(b[122]), .B(n629), .Z(n630) );
  XNOR U885 ( .A(b[122]), .B(n631), .Z(c[122]) );
  XOR U886 ( .A(n632), .B(n633), .Z(n629) );
  ANDN U887 ( .B(n634), .A(n635), .Z(n632) );
  XOR U888 ( .A(b[121]), .B(n633), .Z(n634) );
  XNOR U889 ( .A(b[121]), .B(n635), .Z(c[121]) );
  XOR U890 ( .A(n636), .B(n637), .Z(n633) );
  ANDN U891 ( .B(n638), .A(n639), .Z(n636) );
  XOR U892 ( .A(b[120]), .B(n637), .Z(n638) );
  XNOR U893 ( .A(b[120]), .B(n639), .Z(c[120]) );
  XOR U894 ( .A(n640), .B(n641), .Z(n637) );
  ANDN U895 ( .B(n642), .A(n643), .Z(n640) );
  XOR U896 ( .A(b[119]), .B(n641), .Z(n642) );
  XNOR U897 ( .A(b[11]), .B(n644), .Z(c[11]) );
  XNOR U898 ( .A(b[119]), .B(n643), .Z(c[119]) );
  XOR U899 ( .A(n645), .B(n646), .Z(n641) );
  ANDN U900 ( .B(n647), .A(n648), .Z(n645) );
  XOR U901 ( .A(b[118]), .B(n646), .Z(n647) );
  XNOR U902 ( .A(b[118]), .B(n648), .Z(c[118]) );
  XOR U903 ( .A(n649), .B(n650), .Z(n646) );
  ANDN U904 ( .B(n651), .A(n652), .Z(n649) );
  XOR U905 ( .A(b[117]), .B(n650), .Z(n651) );
  XNOR U906 ( .A(b[117]), .B(n652), .Z(c[117]) );
  XOR U907 ( .A(n653), .B(n654), .Z(n650) );
  ANDN U908 ( .B(n655), .A(n656), .Z(n653) );
  XOR U909 ( .A(b[116]), .B(n654), .Z(n655) );
  XNOR U910 ( .A(b[116]), .B(n656), .Z(c[116]) );
  XOR U911 ( .A(n657), .B(n658), .Z(n654) );
  ANDN U912 ( .B(n659), .A(n660), .Z(n657) );
  XOR U913 ( .A(b[115]), .B(n658), .Z(n659) );
  XNOR U914 ( .A(b[115]), .B(n660), .Z(c[115]) );
  XOR U915 ( .A(n661), .B(n662), .Z(n658) );
  ANDN U916 ( .B(n663), .A(n664), .Z(n661) );
  XOR U917 ( .A(b[114]), .B(n662), .Z(n663) );
  XNOR U918 ( .A(b[114]), .B(n664), .Z(c[114]) );
  XOR U919 ( .A(n665), .B(n666), .Z(n662) );
  ANDN U920 ( .B(n667), .A(n668), .Z(n665) );
  XOR U921 ( .A(b[113]), .B(n666), .Z(n667) );
  XNOR U922 ( .A(b[113]), .B(n668), .Z(c[113]) );
  XOR U923 ( .A(n669), .B(n670), .Z(n666) );
  ANDN U924 ( .B(n671), .A(n672), .Z(n669) );
  XOR U925 ( .A(b[112]), .B(n670), .Z(n671) );
  XNOR U926 ( .A(b[112]), .B(n672), .Z(c[112]) );
  XOR U927 ( .A(n673), .B(n674), .Z(n670) );
  ANDN U928 ( .B(n675), .A(n676), .Z(n673) );
  XOR U929 ( .A(b[111]), .B(n674), .Z(n675) );
  XNOR U930 ( .A(b[111]), .B(n676), .Z(c[111]) );
  XOR U931 ( .A(n677), .B(n678), .Z(n674) );
  ANDN U932 ( .B(n679), .A(n680), .Z(n677) );
  XOR U933 ( .A(b[110]), .B(n678), .Z(n679) );
  XNOR U934 ( .A(b[110]), .B(n680), .Z(c[110]) );
  XOR U935 ( .A(n681), .B(n682), .Z(n678) );
  ANDN U936 ( .B(n683), .A(n684), .Z(n681) );
  XOR U937 ( .A(b[109]), .B(n682), .Z(n683) );
  XNOR U938 ( .A(b[10]), .B(n685), .Z(c[10]) );
  XNOR U939 ( .A(b[109]), .B(n684), .Z(c[109]) );
  XOR U940 ( .A(n686), .B(n687), .Z(n682) );
  ANDN U941 ( .B(n688), .A(n689), .Z(n686) );
  XOR U942 ( .A(b[108]), .B(n687), .Z(n688) );
  XNOR U943 ( .A(b[108]), .B(n689), .Z(c[108]) );
  XOR U944 ( .A(n690), .B(n691), .Z(n687) );
  ANDN U945 ( .B(n692), .A(n693), .Z(n690) );
  XOR U946 ( .A(b[107]), .B(n691), .Z(n692) );
  XNOR U947 ( .A(b[107]), .B(n693), .Z(c[107]) );
  XOR U948 ( .A(n694), .B(n695), .Z(n691) );
  ANDN U949 ( .B(n696), .A(n697), .Z(n694) );
  XOR U950 ( .A(b[106]), .B(n695), .Z(n696) );
  XNOR U951 ( .A(b[106]), .B(n697), .Z(c[106]) );
  XOR U952 ( .A(n698), .B(n699), .Z(n695) );
  ANDN U953 ( .B(n700), .A(n701), .Z(n698) );
  XOR U954 ( .A(b[105]), .B(n699), .Z(n700) );
  XNOR U955 ( .A(b[105]), .B(n701), .Z(c[105]) );
  XOR U956 ( .A(n702), .B(n703), .Z(n699) );
  ANDN U957 ( .B(n704), .A(n705), .Z(n702) );
  XOR U958 ( .A(b[104]), .B(n703), .Z(n704) );
  XNOR U959 ( .A(b[104]), .B(n705), .Z(c[104]) );
  XOR U960 ( .A(n706), .B(n707), .Z(n703) );
  ANDN U961 ( .B(n708), .A(n709), .Z(n706) );
  XOR U962 ( .A(b[103]), .B(n707), .Z(n708) );
  XNOR U963 ( .A(b[103]), .B(n709), .Z(c[103]) );
  XOR U964 ( .A(n710), .B(n711), .Z(n707) );
  ANDN U965 ( .B(n712), .A(n713), .Z(n710) );
  XOR U966 ( .A(b[102]), .B(n711), .Z(n712) );
  XNOR U967 ( .A(b[102]), .B(n713), .Z(c[102]) );
  XOR U968 ( .A(n714), .B(n715), .Z(n711) );
  ANDN U969 ( .B(n716), .A(n717), .Z(n714) );
  XOR U970 ( .A(b[101]), .B(n715), .Z(n716) );
  XNOR U971 ( .A(b[101]), .B(n717), .Z(c[101]) );
  XOR U972 ( .A(n718), .B(n719), .Z(n715) );
  ANDN U973 ( .B(n720), .A(n721), .Z(n718) );
  XOR U974 ( .A(b[100]), .B(n719), .Z(n720) );
  XNOR U975 ( .A(b[100]), .B(n721), .Z(c[100]) );
  XOR U976 ( .A(n722), .B(n723), .Z(n719) );
  ANDN U977 ( .B(n724), .A(n2), .Z(n722) );
  XOR U978 ( .A(b[99]), .B(n723), .Z(n724) );
  XOR U979 ( .A(n725), .B(n726), .Z(n723) );
  ANDN U980 ( .B(n727), .A(n3), .Z(n725) );
  XOR U981 ( .A(b[98]), .B(n726), .Z(n727) );
  XOR U982 ( .A(n728), .B(n729), .Z(n726) );
  ANDN U983 ( .B(n730), .A(n4), .Z(n728) );
  XOR U984 ( .A(b[97]), .B(n729), .Z(n730) );
  XOR U985 ( .A(n731), .B(n732), .Z(n729) );
  ANDN U986 ( .B(n733), .A(n5), .Z(n731) );
  XOR U987 ( .A(b[96]), .B(n732), .Z(n733) );
  XOR U988 ( .A(n734), .B(n735), .Z(n732) );
  ANDN U989 ( .B(n736), .A(n6), .Z(n734) );
  XOR U990 ( .A(b[95]), .B(n735), .Z(n736) );
  XOR U991 ( .A(n737), .B(n738), .Z(n735) );
  ANDN U992 ( .B(n739), .A(n7), .Z(n737) );
  XOR U993 ( .A(b[94]), .B(n738), .Z(n739) );
  XOR U994 ( .A(n740), .B(n741), .Z(n738) );
  ANDN U995 ( .B(n742), .A(n8), .Z(n740) );
  XOR U996 ( .A(b[93]), .B(n741), .Z(n742) );
  XOR U997 ( .A(n743), .B(n744), .Z(n741) );
  ANDN U998 ( .B(n745), .A(n9), .Z(n743) );
  XOR U999 ( .A(b[92]), .B(n744), .Z(n745) );
  XOR U1000 ( .A(n746), .B(n747), .Z(n744) );
  ANDN U1001 ( .B(n748), .A(n10), .Z(n746) );
  XOR U1002 ( .A(b[91]), .B(n747), .Z(n748) );
  XOR U1003 ( .A(n749), .B(n750), .Z(n747) );
  ANDN U1004 ( .B(n751), .A(n11), .Z(n749) );
  XOR U1005 ( .A(b[90]), .B(n750), .Z(n751) );
  XOR U1006 ( .A(n752), .B(n753), .Z(n750) );
  ANDN U1007 ( .B(n754), .A(n13), .Z(n752) );
  XOR U1008 ( .A(b[89]), .B(n753), .Z(n754) );
  XOR U1009 ( .A(n755), .B(n756), .Z(n753) );
  ANDN U1010 ( .B(n757), .A(n14), .Z(n755) );
  XOR U1011 ( .A(b[88]), .B(n756), .Z(n757) );
  XOR U1012 ( .A(n758), .B(n759), .Z(n756) );
  ANDN U1013 ( .B(n760), .A(n15), .Z(n758) );
  XOR U1014 ( .A(b[87]), .B(n759), .Z(n760) );
  XOR U1015 ( .A(n761), .B(n762), .Z(n759) );
  ANDN U1016 ( .B(n763), .A(n16), .Z(n761) );
  XOR U1017 ( .A(b[86]), .B(n762), .Z(n763) );
  XOR U1018 ( .A(n764), .B(n765), .Z(n762) );
  ANDN U1019 ( .B(n766), .A(n17), .Z(n764) );
  XOR U1020 ( .A(b[85]), .B(n765), .Z(n766) );
  XOR U1021 ( .A(n767), .B(n768), .Z(n765) );
  ANDN U1022 ( .B(n769), .A(n18), .Z(n767) );
  XOR U1023 ( .A(b[84]), .B(n768), .Z(n769) );
  XOR U1024 ( .A(n770), .B(n771), .Z(n768) );
  ANDN U1025 ( .B(n772), .A(n19), .Z(n770) );
  XOR U1026 ( .A(b[83]), .B(n771), .Z(n772) );
  XOR U1027 ( .A(n773), .B(n774), .Z(n771) );
  ANDN U1028 ( .B(n775), .A(n20), .Z(n773) );
  XOR U1029 ( .A(b[82]), .B(n774), .Z(n775) );
  XOR U1030 ( .A(n776), .B(n777), .Z(n774) );
  ANDN U1031 ( .B(n778), .A(n21), .Z(n776) );
  XOR U1032 ( .A(b[81]), .B(n777), .Z(n778) );
  XOR U1033 ( .A(n779), .B(n780), .Z(n777) );
  ANDN U1034 ( .B(n781), .A(n22), .Z(n779) );
  XOR U1035 ( .A(b[80]), .B(n780), .Z(n781) );
  XOR U1036 ( .A(n782), .B(n783), .Z(n780) );
  ANDN U1037 ( .B(n784), .A(n24), .Z(n782) );
  XOR U1038 ( .A(b[79]), .B(n783), .Z(n784) );
  XOR U1039 ( .A(n785), .B(n786), .Z(n783) );
  ANDN U1040 ( .B(n787), .A(n25), .Z(n785) );
  XOR U1041 ( .A(b[78]), .B(n786), .Z(n787) );
  XOR U1042 ( .A(n788), .B(n789), .Z(n786) );
  ANDN U1043 ( .B(n790), .A(n26), .Z(n788) );
  XOR U1044 ( .A(b[77]), .B(n789), .Z(n790) );
  XOR U1045 ( .A(n791), .B(n792), .Z(n789) );
  ANDN U1046 ( .B(n793), .A(n27), .Z(n791) );
  XOR U1047 ( .A(b[76]), .B(n792), .Z(n793) );
  XOR U1048 ( .A(n794), .B(n795), .Z(n792) );
  ANDN U1049 ( .B(n796), .A(n28), .Z(n794) );
  XOR U1050 ( .A(b[75]), .B(n795), .Z(n796) );
  XOR U1051 ( .A(n797), .B(n798), .Z(n795) );
  ANDN U1052 ( .B(n799), .A(n29), .Z(n797) );
  XOR U1053 ( .A(b[74]), .B(n798), .Z(n799) );
  XOR U1054 ( .A(n800), .B(n801), .Z(n798) );
  ANDN U1055 ( .B(n802), .A(n30), .Z(n800) );
  XOR U1056 ( .A(b[73]), .B(n801), .Z(n802) );
  XOR U1057 ( .A(n803), .B(n804), .Z(n801) );
  ANDN U1058 ( .B(n805), .A(n31), .Z(n803) );
  XOR U1059 ( .A(b[72]), .B(n804), .Z(n805) );
  XOR U1060 ( .A(n806), .B(n807), .Z(n804) );
  ANDN U1061 ( .B(n808), .A(n32), .Z(n806) );
  XOR U1062 ( .A(b[71]), .B(n807), .Z(n808) );
  XOR U1063 ( .A(n809), .B(n810), .Z(n807) );
  ANDN U1064 ( .B(n811), .A(n33), .Z(n809) );
  XOR U1065 ( .A(b[70]), .B(n810), .Z(n811) );
  XOR U1066 ( .A(n812), .B(n813), .Z(n810) );
  ANDN U1067 ( .B(n814), .A(n35), .Z(n812) );
  XOR U1068 ( .A(b[69]), .B(n813), .Z(n814) );
  XOR U1069 ( .A(n815), .B(n816), .Z(n813) );
  ANDN U1070 ( .B(n817), .A(n36), .Z(n815) );
  XOR U1071 ( .A(b[68]), .B(n816), .Z(n817) );
  XOR U1072 ( .A(n818), .B(n819), .Z(n816) );
  ANDN U1073 ( .B(n820), .A(n37), .Z(n818) );
  XOR U1074 ( .A(b[67]), .B(n819), .Z(n820) );
  XOR U1075 ( .A(n821), .B(n822), .Z(n819) );
  ANDN U1076 ( .B(n823), .A(n38), .Z(n821) );
  XOR U1077 ( .A(b[66]), .B(n822), .Z(n823) );
  XOR U1078 ( .A(n824), .B(n825), .Z(n822) );
  ANDN U1079 ( .B(n826), .A(n39), .Z(n824) );
  XOR U1080 ( .A(b[65]), .B(n825), .Z(n826) );
  XOR U1081 ( .A(n827), .B(n828), .Z(n825) );
  ANDN U1082 ( .B(n829), .A(n40), .Z(n827) );
  XOR U1083 ( .A(b[64]), .B(n828), .Z(n829) );
  XOR U1084 ( .A(n830), .B(n831), .Z(n828) );
  ANDN U1085 ( .B(n832), .A(n41), .Z(n830) );
  XOR U1086 ( .A(b[63]), .B(n831), .Z(n832) );
  XOR U1087 ( .A(n833), .B(n834), .Z(n831) );
  ANDN U1088 ( .B(n835), .A(n42), .Z(n833) );
  XOR U1089 ( .A(b[62]), .B(n834), .Z(n835) );
  XOR U1090 ( .A(n836), .B(n837), .Z(n834) );
  ANDN U1091 ( .B(n838), .A(n43), .Z(n836) );
  XOR U1092 ( .A(b[61]), .B(n837), .Z(n838) );
  XOR U1093 ( .A(n839), .B(n840), .Z(n837) );
  ANDN U1094 ( .B(n841), .A(n44), .Z(n839) );
  XOR U1095 ( .A(b[60]), .B(n840), .Z(n841) );
  XOR U1096 ( .A(n842), .B(n843), .Z(n840) );
  ANDN U1097 ( .B(n844), .A(n46), .Z(n842) );
  XOR U1098 ( .A(b[59]), .B(n843), .Z(n844) );
  XOR U1099 ( .A(n845), .B(n846), .Z(n843) );
  ANDN U1100 ( .B(n847), .A(n47), .Z(n845) );
  XOR U1101 ( .A(b[58]), .B(n846), .Z(n847) );
  XOR U1102 ( .A(n848), .B(n849), .Z(n846) );
  ANDN U1103 ( .B(n850), .A(n48), .Z(n848) );
  XOR U1104 ( .A(b[57]), .B(n849), .Z(n850) );
  XOR U1105 ( .A(n851), .B(n852), .Z(n849) );
  ANDN U1106 ( .B(n853), .A(n49), .Z(n851) );
  XOR U1107 ( .A(b[56]), .B(n852), .Z(n853) );
  XOR U1108 ( .A(n854), .B(n855), .Z(n852) );
  ANDN U1109 ( .B(n856), .A(n50), .Z(n854) );
  XOR U1110 ( .A(b[55]), .B(n855), .Z(n856) );
  XOR U1111 ( .A(n857), .B(n858), .Z(n855) );
  ANDN U1112 ( .B(n859), .A(n51), .Z(n857) );
  XOR U1113 ( .A(b[54]), .B(n858), .Z(n859) );
  XOR U1114 ( .A(n860), .B(n861), .Z(n858) );
  ANDN U1115 ( .B(n862), .A(n52), .Z(n860) );
  XOR U1116 ( .A(b[53]), .B(n861), .Z(n862) );
  XOR U1117 ( .A(n863), .B(n864), .Z(n861) );
  ANDN U1118 ( .B(n865), .A(n53), .Z(n863) );
  XOR U1119 ( .A(b[52]), .B(n864), .Z(n865) );
  XOR U1120 ( .A(n866), .B(n867), .Z(n864) );
  ANDN U1121 ( .B(n868), .A(n54), .Z(n866) );
  XOR U1122 ( .A(b[51]), .B(n867), .Z(n868) );
  XOR U1123 ( .A(n869), .B(n870), .Z(n867) );
  ANDN U1124 ( .B(n871), .A(n55), .Z(n869) );
  XOR U1125 ( .A(b[50]), .B(n870), .Z(n871) );
  XOR U1126 ( .A(n872), .B(n873), .Z(n870) );
  ANDN U1127 ( .B(n874), .A(n57), .Z(n872) );
  XOR U1128 ( .A(b[49]), .B(n873), .Z(n874) );
  XOR U1129 ( .A(n875), .B(n876), .Z(n873) );
  ANDN U1130 ( .B(n877), .A(n58), .Z(n875) );
  XOR U1131 ( .A(b[48]), .B(n876), .Z(n877) );
  XOR U1132 ( .A(n878), .B(n879), .Z(n876) );
  ANDN U1133 ( .B(n880), .A(n59), .Z(n878) );
  XOR U1134 ( .A(b[47]), .B(n879), .Z(n880) );
  XOR U1135 ( .A(n881), .B(n882), .Z(n879) );
  ANDN U1136 ( .B(n883), .A(n60), .Z(n881) );
  XOR U1137 ( .A(b[46]), .B(n882), .Z(n883) );
  XOR U1138 ( .A(n884), .B(n885), .Z(n882) );
  ANDN U1139 ( .B(n886), .A(n61), .Z(n884) );
  XOR U1140 ( .A(b[45]), .B(n885), .Z(n886) );
  XOR U1141 ( .A(n887), .B(n888), .Z(n885) );
  ANDN U1142 ( .B(n889), .A(n62), .Z(n887) );
  XOR U1143 ( .A(b[44]), .B(n888), .Z(n889) );
  XOR U1144 ( .A(n890), .B(n891), .Z(n888) );
  ANDN U1145 ( .B(n892), .A(n63), .Z(n890) );
  XOR U1146 ( .A(b[43]), .B(n891), .Z(n892) );
  XOR U1147 ( .A(n893), .B(n894), .Z(n891) );
  ANDN U1148 ( .B(n895), .A(n64), .Z(n893) );
  XOR U1149 ( .A(b[42]), .B(n894), .Z(n895) );
  XOR U1150 ( .A(n896), .B(n897), .Z(n894) );
  ANDN U1151 ( .B(n898), .A(n65), .Z(n896) );
  XOR U1152 ( .A(b[41]), .B(n897), .Z(n898) );
  XOR U1153 ( .A(n899), .B(n900), .Z(n897) );
  ANDN U1154 ( .B(n901), .A(n66), .Z(n899) );
  XOR U1155 ( .A(b[40]), .B(n900), .Z(n901) );
  XOR U1156 ( .A(n902), .B(n903), .Z(n900) );
  ANDN U1157 ( .B(n904), .A(n68), .Z(n902) );
  XOR U1158 ( .A(b[39]), .B(n903), .Z(n904) );
  XOR U1159 ( .A(n905), .B(n906), .Z(n903) );
  ANDN U1160 ( .B(n907), .A(n69), .Z(n905) );
  XOR U1161 ( .A(b[38]), .B(n906), .Z(n907) );
  XOR U1162 ( .A(n908), .B(n909), .Z(n906) );
  ANDN U1163 ( .B(n910), .A(n70), .Z(n908) );
  XOR U1164 ( .A(b[37]), .B(n909), .Z(n910) );
  XOR U1165 ( .A(n911), .B(n912), .Z(n909) );
  ANDN U1166 ( .B(n913), .A(n71), .Z(n911) );
  XOR U1167 ( .A(b[36]), .B(n912), .Z(n913) );
  XOR U1168 ( .A(n914), .B(n915), .Z(n912) );
  ANDN U1169 ( .B(n916), .A(n72), .Z(n914) );
  XOR U1170 ( .A(b[35]), .B(n915), .Z(n916) );
  XOR U1171 ( .A(n917), .B(n918), .Z(n915) );
  ANDN U1172 ( .B(n919), .A(n73), .Z(n917) );
  XOR U1173 ( .A(b[34]), .B(n918), .Z(n919) );
  XOR U1174 ( .A(n920), .B(n921), .Z(n918) );
  ANDN U1175 ( .B(n922), .A(n74), .Z(n920) );
  XOR U1176 ( .A(b[33]), .B(n921), .Z(n922) );
  XOR U1177 ( .A(n923), .B(n924), .Z(n921) );
  ANDN U1178 ( .B(n925), .A(n75), .Z(n923) );
  XOR U1179 ( .A(b[32]), .B(n924), .Z(n925) );
  XOR U1180 ( .A(n926), .B(n927), .Z(n924) );
  ANDN U1181 ( .B(n928), .A(n76), .Z(n926) );
  XOR U1182 ( .A(b[31]), .B(n927), .Z(n928) );
  XOR U1183 ( .A(n929), .B(n930), .Z(n927) );
  ANDN U1184 ( .B(n931), .A(n77), .Z(n929) );
  XOR U1185 ( .A(b[30]), .B(n930), .Z(n931) );
  XOR U1186 ( .A(n932), .B(n933), .Z(n930) );
  ANDN U1187 ( .B(n934), .A(n79), .Z(n932) );
  XOR U1188 ( .A(b[29]), .B(n933), .Z(n934) );
  XOR U1189 ( .A(n935), .B(n936), .Z(n933) );
  ANDN U1190 ( .B(n937), .A(n80), .Z(n935) );
  XOR U1191 ( .A(b[28]), .B(n936), .Z(n937) );
  XOR U1192 ( .A(n938), .B(n939), .Z(n936) );
  ANDN U1193 ( .B(n940), .A(n81), .Z(n938) );
  XOR U1194 ( .A(b[27]), .B(n939), .Z(n940) );
  XOR U1195 ( .A(n941), .B(n942), .Z(n939) );
  ANDN U1196 ( .B(n943), .A(n82), .Z(n941) );
  XOR U1197 ( .A(b[26]), .B(n942), .Z(n943) );
  XOR U1198 ( .A(n944), .B(n945), .Z(n942) );
  ANDN U1199 ( .B(n946), .A(n83), .Z(n944) );
  XOR U1200 ( .A(b[25]), .B(n945), .Z(n946) );
  XOR U1201 ( .A(n947), .B(n948), .Z(n945) );
  ANDN U1202 ( .B(n949), .A(n110), .Z(n947) );
  XOR U1203 ( .A(b[24]), .B(n948), .Z(n949) );
  XOR U1204 ( .A(n950), .B(n951), .Z(n948) );
  ANDN U1205 ( .B(n952), .A(n151), .Z(n950) );
  XOR U1206 ( .A(b[23]), .B(n951), .Z(n952) );
  XOR U1207 ( .A(n953), .B(n954), .Z(n951) );
  ANDN U1208 ( .B(n955), .A(n192), .Z(n953) );
  XOR U1209 ( .A(b[22]), .B(n954), .Z(n955) );
  XOR U1210 ( .A(n956), .B(n957), .Z(n954) );
  ANDN U1211 ( .B(n958), .A(n233), .Z(n956) );
  XOR U1212 ( .A(b[21]), .B(n957), .Z(n958) );
  XOR U1213 ( .A(n959), .B(n960), .Z(n957) );
  ANDN U1214 ( .B(n961), .A(n274), .Z(n959) );
  XOR U1215 ( .A(b[20]), .B(n960), .Z(n961) );
  XOR U1216 ( .A(n962), .B(n963), .Z(n960) );
  ANDN U1217 ( .B(n964), .A(n316), .Z(n962) );
  XOR U1218 ( .A(b[19]), .B(n963), .Z(n964) );
  XOR U1219 ( .A(n965), .B(n966), .Z(n963) );
  ANDN U1220 ( .B(n967), .A(n357), .Z(n965) );
  XOR U1221 ( .A(b[18]), .B(n966), .Z(n967) );
  XOR U1222 ( .A(n968), .B(n969), .Z(n966) );
  ANDN U1223 ( .B(n970), .A(n398), .Z(n968) );
  XOR U1224 ( .A(b[17]), .B(n969), .Z(n970) );
  XOR U1225 ( .A(n971), .B(n972), .Z(n969) );
  ANDN U1226 ( .B(n973), .A(n439), .Z(n971) );
  XOR U1227 ( .A(b[16]), .B(n972), .Z(n973) );
  XOR U1228 ( .A(n974), .B(n975), .Z(n972) );
  ANDN U1229 ( .B(n976), .A(n480), .Z(n974) );
  XOR U1230 ( .A(b[15]), .B(n975), .Z(n976) );
  XOR U1231 ( .A(n977), .B(n978), .Z(n975) );
  ANDN U1232 ( .B(n979), .A(n521), .Z(n977) );
  XOR U1233 ( .A(b[14]), .B(n978), .Z(n979) );
  XOR U1234 ( .A(n980), .B(n981), .Z(n978) );
  ANDN U1235 ( .B(n982), .A(n562), .Z(n980) );
  XOR U1236 ( .A(b[13]), .B(n981), .Z(n982) );
  XOR U1237 ( .A(n983), .B(n984), .Z(n981) );
  ANDN U1238 ( .B(n985), .A(n603), .Z(n983) );
  XOR U1239 ( .A(b[12]), .B(n984), .Z(n985) );
  XOR U1240 ( .A(n986), .B(n987), .Z(n984) );
  ANDN U1241 ( .B(n988), .A(n644), .Z(n986) );
  XOR U1242 ( .A(b[11]), .B(n987), .Z(n988) );
  XOR U1243 ( .A(n989), .B(n990), .Z(n987) );
  ANDN U1244 ( .B(n991), .A(n685), .Z(n989) );
  XOR U1245 ( .A(b[10]), .B(n990), .Z(n991) );
  XOR U1246 ( .A(n992), .B(n993), .Z(n990) );
  ANDN U1247 ( .B(n994), .A(n1), .Z(n992) );
  XOR U1248 ( .A(b[9]), .B(n993), .Z(n994) );
  XOR U1249 ( .A(n995), .B(n996), .Z(n993) );
  ANDN U1250 ( .B(n997), .A(n12), .Z(n995) );
  XOR U1251 ( .A(b[8]), .B(n996), .Z(n997) );
  XOR U1252 ( .A(n998), .B(n999), .Z(n996) );
  ANDN U1253 ( .B(n1000), .A(n23), .Z(n998) );
  XOR U1254 ( .A(b[7]), .B(n999), .Z(n1000) );
  XOR U1255 ( .A(n1001), .B(n1002), .Z(n999) );
  ANDN U1256 ( .B(n1003), .A(n34), .Z(n1001) );
  XOR U1257 ( .A(b[6]), .B(n1002), .Z(n1003) );
  XOR U1258 ( .A(n1004), .B(n1005), .Z(n1002) );
  ANDN U1259 ( .B(n1006), .A(n45), .Z(n1004) );
  XOR U1260 ( .A(b[5]), .B(n1005), .Z(n1006) );
  XOR U1261 ( .A(n1007), .B(n1008), .Z(n1005) );
  ANDN U1262 ( .B(n1009), .A(n56), .Z(n1007) );
  XOR U1263 ( .A(b[4]), .B(n1008), .Z(n1009) );
  XOR U1264 ( .A(n1010), .B(n1011), .Z(n1008) );
  ANDN U1265 ( .B(n1012), .A(n67), .Z(n1010) );
  XOR U1266 ( .A(b[3]), .B(n1011), .Z(n1012) );
  XOR U1267 ( .A(n1013), .B(n1014), .Z(n1011) );
  ANDN U1268 ( .B(n1015), .A(n78), .Z(n1013) );
  XOR U1269 ( .A(b[2]), .B(n1014), .Z(n1015) );
  XNOR U1270 ( .A(n1016), .B(n1017), .Z(n1014) );
  NANDN U1271 ( .A(n315), .B(n1018), .Z(n1017) );
  XOR U1272 ( .A(b[1]), .B(n1016), .Z(n1018) );
  XNOR U1273 ( .A(a[1]), .B(n1016), .Z(n315) );
  AND U1274 ( .A(b[0]), .B(a[0]), .Z(n1016) );
  XOR U1275 ( .A(b[0]), .B(a[0]), .Z(c[0]) );
endmodule

