
module sum ( a, b, c );
  input [127:0] a;
  input [127:0] b;
  output [128:0] c;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112;

  IV U2 ( .A(n977), .Z(n2) );
  IV U3 ( .A(b[3]), .Z(n3) );
  NOR U4 ( .A(n2), .B(n3), .Z(n4) );
  XOR U5 ( .A(n977), .B(n3), .Z(n5) );
  IV U6 ( .A(a[3]), .Z(n6) );
  NOR U7 ( .A(n5), .B(n6), .Z(n7) );
  NOR U8 ( .A(n4), .B(n7), .Z(n8) );
  IV U9 ( .A(n8), .Z(n999) );
  IV U10 ( .A(n1043), .Z(n9) );
  IV U11 ( .A(b[6]), .Z(n10) );
  NOR U12 ( .A(n9), .B(n10), .Z(n11) );
  XOR U13 ( .A(n1043), .B(n10), .Z(n12) );
  IV U14 ( .A(a[6]), .Z(n13) );
  NOR U15 ( .A(n12), .B(n13), .Z(n14) );
  NOR U16 ( .A(n11), .B(n14), .Z(n15) );
  IV U17 ( .A(n15), .Z(n1065) );
  IV U18 ( .A(n1109), .Z(n16) );
  IV U19 ( .A(a[9]), .Z(n17) );
  NOR U20 ( .A(n16), .B(n17), .Z(n18) );
  XOR U21 ( .A(n1109), .B(n17), .Z(n19) );
  IV U22 ( .A(b[9]), .Z(n20) );
  NOR U23 ( .A(n19), .B(n20), .Z(n21) );
  NOR U24 ( .A(n18), .B(n21), .Z(n22) );
  IV U25 ( .A(n22), .Z(n834) );
  IV U26 ( .A(n916), .Z(n23) );
  IV U27 ( .A(b[12]), .Z(n24) );
  NOR U28 ( .A(n23), .B(n24), .Z(n25) );
  XOR U29 ( .A(n916), .B(n24), .Z(n26) );
  IV U30 ( .A(a[12]), .Z(n27) );
  NOR U31 ( .A(n26), .B(n27), .Z(n28) );
  NOR U32 ( .A(n25), .B(n28), .Z(n29) );
  IV U33 ( .A(n29), .Z(n918) );
  IV U34 ( .A(n922), .Z(n30) );
  IV U35 ( .A(b[15]), .Z(n31) );
  NOR U36 ( .A(n30), .B(n31), .Z(n32) );
  XOR U37 ( .A(n922), .B(n31), .Z(n33) );
  IV U38 ( .A(a[15]), .Z(n34) );
  NOR U39 ( .A(n33), .B(n34), .Z(n35) );
  NOR U40 ( .A(n32), .B(n35), .Z(n36) );
  IV U41 ( .A(n36), .Z(n924) );
  IV U42 ( .A(n928), .Z(n37) );
  IV U43 ( .A(b[18]), .Z(n38) );
  NOR U44 ( .A(n37), .B(n38), .Z(n39) );
  XOR U45 ( .A(n928), .B(n38), .Z(n40) );
  IV U46 ( .A(a[18]), .Z(n41) );
  NOR U47 ( .A(n40), .B(n41), .Z(n42) );
  NOR U48 ( .A(n39), .B(n42), .Z(n43) );
  IV U49 ( .A(n43), .Z(n930) );
  IV U50 ( .A(n936), .Z(n44) );
  IV U51 ( .A(b[21]), .Z(n45) );
  NOR U52 ( .A(n44), .B(n45), .Z(n46) );
  XOR U53 ( .A(n936), .B(n45), .Z(n47) );
  IV U54 ( .A(a[21]), .Z(n48) );
  NOR U55 ( .A(n47), .B(n48), .Z(n49) );
  NOR U56 ( .A(n46), .B(n49), .Z(n50) );
  IV U57 ( .A(n50), .Z(n938) );
  IV U58 ( .A(n942), .Z(n51) );
  IV U59 ( .A(b[24]), .Z(n52) );
  NOR U60 ( .A(n51), .B(n52), .Z(n53) );
  XOR U61 ( .A(n942), .B(n52), .Z(n54) );
  IV U62 ( .A(a[24]), .Z(n55) );
  NOR U63 ( .A(n54), .B(n55), .Z(n56) );
  NOR U64 ( .A(n53), .B(n56), .Z(n57) );
  IV U65 ( .A(n57), .Z(n944) );
  IV U66 ( .A(n948), .Z(n58) );
  IV U67 ( .A(b[27]), .Z(n59) );
  NOR U68 ( .A(n58), .B(n59), .Z(n60) );
  XOR U69 ( .A(n948), .B(n59), .Z(n61) );
  IV U70 ( .A(a[27]), .Z(n62) );
  NOR U71 ( .A(n61), .B(n62), .Z(n63) );
  NOR U72 ( .A(n60), .B(n63), .Z(n64) );
  IV U73 ( .A(n64), .Z(n950) );
  IV U74 ( .A(n957), .Z(n65) );
  IV U75 ( .A(b[30]), .Z(n66) );
  NOR U76 ( .A(n65), .B(n66), .Z(n67) );
  XOR U77 ( .A(n957), .B(n66), .Z(n68) );
  IV U78 ( .A(a[30]), .Z(n69) );
  NOR U79 ( .A(n68), .B(n69), .Z(n70) );
  NOR U80 ( .A(n67), .B(n70), .Z(n71) );
  IV U81 ( .A(n71), .Z(n959) );
  IV U82 ( .A(n963), .Z(n72) );
  IV U83 ( .A(b[33]), .Z(n73) );
  NOR U84 ( .A(n72), .B(n73), .Z(n74) );
  XOR U85 ( .A(n963), .B(n73), .Z(n75) );
  IV U86 ( .A(a[33]), .Z(n76) );
  NOR U87 ( .A(n75), .B(n76), .Z(n77) );
  NOR U88 ( .A(n74), .B(n77), .Z(n78) );
  IV U89 ( .A(n78), .Z(n965) );
  IV U90 ( .A(n969), .Z(n79) );
  IV U91 ( .A(b[36]), .Z(n80) );
  NOR U92 ( .A(n79), .B(n80), .Z(n81) );
  XOR U93 ( .A(n969), .B(n80), .Z(n82) );
  IV U94 ( .A(a[36]), .Z(n83) );
  NOR U95 ( .A(n82), .B(n83), .Z(n84) );
  NOR U96 ( .A(n81), .B(n84), .Z(n85) );
  IV U97 ( .A(n85), .Z(n971) );
  IV U98 ( .A(n975), .Z(n86) );
  IV U99 ( .A(b[39]), .Z(n87) );
  NOR U100 ( .A(n86), .B(n87), .Z(n88) );
  XOR U101 ( .A(n975), .B(n87), .Z(n89) );
  IV U102 ( .A(a[39]), .Z(n90) );
  NOR U103 ( .A(n89), .B(n90), .Z(n91) );
  NOR U104 ( .A(n88), .B(n91), .Z(n92) );
  IV U105 ( .A(n92), .Z(n979) );
  IV U106 ( .A(n983), .Z(n93) );
  IV U107 ( .A(b[42]), .Z(n94) );
  NOR U108 ( .A(n93), .B(n94), .Z(n95) );
  XOR U109 ( .A(n983), .B(n94), .Z(n96) );
  IV U110 ( .A(a[42]), .Z(n97) );
  NOR U111 ( .A(n96), .B(n97), .Z(n98) );
  NOR U112 ( .A(n95), .B(n98), .Z(n99) );
  IV U113 ( .A(n99), .Z(n985) );
  IV U114 ( .A(n989), .Z(n100) );
  IV U115 ( .A(b[45]), .Z(n101) );
  NOR U116 ( .A(n100), .B(n101), .Z(n102) );
  XOR U117 ( .A(n989), .B(n101), .Z(n103) );
  IV U118 ( .A(a[45]), .Z(n104) );
  NOR U119 ( .A(n103), .B(n104), .Z(n105) );
  NOR U120 ( .A(n102), .B(n105), .Z(n106) );
  IV U121 ( .A(n106), .Z(n991) );
  IV U122 ( .A(n995), .Z(n107) );
  IV U123 ( .A(b[48]), .Z(n108) );
  NOR U124 ( .A(n107), .B(n108), .Z(n109) );
  XOR U125 ( .A(n995), .B(n108), .Z(n110) );
  IV U126 ( .A(a[48]), .Z(n111) );
  NOR U127 ( .A(n110), .B(n111), .Z(n112) );
  NOR U128 ( .A(n109), .B(n112), .Z(n113) );
  IV U129 ( .A(n113), .Z(n997) );
  IV U130 ( .A(n1003), .Z(n114) );
  IV U131 ( .A(b[51]), .Z(n115) );
  NOR U132 ( .A(n114), .B(n115), .Z(n116) );
  XOR U133 ( .A(n1003), .B(n115), .Z(n117) );
  IV U134 ( .A(a[51]), .Z(n118) );
  NOR U135 ( .A(n117), .B(n118), .Z(n119) );
  NOR U136 ( .A(n116), .B(n119), .Z(n120) );
  IV U137 ( .A(n120), .Z(n1005) );
  IV U138 ( .A(n1009), .Z(n121) );
  IV U139 ( .A(b[54]), .Z(n122) );
  NOR U140 ( .A(n121), .B(n122), .Z(n123) );
  XOR U141 ( .A(n1009), .B(n122), .Z(n124) );
  IV U142 ( .A(a[54]), .Z(n125) );
  NOR U143 ( .A(n124), .B(n125), .Z(n126) );
  NOR U144 ( .A(n123), .B(n126), .Z(n127) );
  IV U145 ( .A(n127), .Z(n1011) );
  IV U146 ( .A(n1015), .Z(n128) );
  IV U147 ( .A(b[57]), .Z(n129) );
  NOR U148 ( .A(n128), .B(n129), .Z(n130) );
  XOR U149 ( .A(n1015), .B(n129), .Z(n131) );
  IV U150 ( .A(a[57]), .Z(n132) );
  NOR U151 ( .A(n131), .B(n132), .Z(n133) );
  NOR U152 ( .A(n130), .B(n133), .Z(n134) );
  IV U153 ( .A(n134), .Z(n1017) );
  IV U154 ( .A(n1023), .Z(n135) );
  IV U155 ( .A(b[60]), .Z(n136) );
  NOR U156 ( .A(n135), .B(n136), .Z(n137) );
  XOR U157 ( .A(n1023), .B(n136), .Z(n138) );
  IV U158 ( .A(a[60]), .Z(n139) );
  NOR U159 ( .A(n138), .B(n139), .Z(n140) );
  NOR U160 ( .A(n137), .B(n140), .Z(n141) );
  IV U161 ( .A(n141), .Z(n1025) );
  IV U162 ( .A(n1029), .Z(n142) );
  IV U163 ( .A(b[63]), .Z(n143) );
  NOR U164 ( .A(n142), .B(n143), .Z(n144) );
  XOR U165 ( .A(n1029), .B(n143), .Z(n145) );
  IV U166 ( .A(a[63]), .Z(n146) );
  NOR U167 ( .A(n145), .B(n146), .Z(n147) );
  NOR U168 ( .A(n144), .B(n147), .Z(n148) );
  IV U169 ( .A(n148), .Z(n1031) );
  IV U170 ( .A(n1035), .Z(n149) );
  IV U171 ( .A(b[66]), .Z(n150) );
  NOR U172 ( .A(n149), .B(n150), .Z(n151) );
  XOR U173 ( .A(n1035), .B(n150), .Z(n152) );
  IV U174 ( .A(a[66]), .Z(n153) );
  NOR U175 ( .A(n152), .B(n153), .Z(n154) );
  NOR U176 ( .A(n151), .B(n154), .Z(n155) );
  IV U177 ( .A(n155), .Z(n1037) );
  IV U178 ( .A(n1041), .Z(n156) );
  IV U179 ( .A(b[69]), .Z(n157) );
  NOR U180 ( .A(n156), .B(n157), .Z(n158) );
  XOR U181 ( .A(n1041), .B(n157), .Z(n159) );
  IV U182 ( .A(a[69]), .Z(n160) );
  NOR U183 ( .A(n159), .B(n160), .Z(n161) );
  NOR U184 ( .A(n158), .B(n161), .Z(n162) );
  IV U185 ( .A(n162), .Z(n1045) );
  IV U186 ( .A(n1049), .Z(n163) );
  IV U187 ( .A(b[72]), .Z(n164) );
  NOR U188 ( .A(n163), .B(n164), .Z(n165) );
  XOR U189 ( .A(n1049), .B(n164), .Z(n166) );
  IV U190 ( .A(a[72]), .Z(n167) );
  NOR U191 ( .A(n166), .B(n167), .Z(n168) );
  NOR U192 ( .A(n165), .B(n168), .Z(n169) );
  IV U193 ( .A(n169), .Z(n1051) );
  IV U194 ( .A(n1055), .Z(n170) );
  IV U195 ( .A(b[75]), .Z(n171) );
  NOR U196 ( .A(n170), .B(n171), .Z(n172) );
  XOR U197 ( .A(n1055), .B(n171), .Z(n173) );
  IV U198 ( .A(a[75]), .Z(n174) );
  NOR U199 ( .A(n173), .B(n174), .Z(n175) );
  NOR U200 ( .A(n172), .B(n175), .Z(n176) );
  IV U201 ( .A(n176), .Z(n1057) );
  IV U202 ( .A(n1061), .Z(n177) );
  IV U203 ( .A(b[78]), .Z(n178) );
  NOR U204 ( .A(n177), .B(n178), .Z(n179) );
  XOR U205 ( .A(n1061), .B(n178), .Z(n180) );
  IV U206 ( .A(a[78]), .Z(n181) );
  NOR U207 ( .A(n180), .B(n181), .Z(n182) );
  NOR U208 ( .A(n179), .B(n182), .Z(n183) );
  IV U209 ( .A(n183), .Z(n1063) );
  IV U210 ( .A(n1069), .Z(n184) );
  IV U211 ( .A(b[81]), .Z(n185) );
  NOR U212 ( .A(n184), .B(n185), .Z(n186) );
  XOR U213 ( .A(n1069), .B(n185), .Z(n187) );
  IV U214 ( .A(a[81]), .Z(n188) );
  NOR U215 ( .A(n187), .B(n188), .Z(n189) );
  NOR U216 ( .A(n186), .B(n189), .Z(n190) );
  IV U217 ( .A(n190), .Z(n1071) );
  IV U218 ( .A(n1075), .Z(n191) );
  IV U219 ( .A(b[84]), .Z(n192) );
  NOR U220 ( .A(n191), .B(n192), .Z(n193) );
  XOR U221 ( .A(n1075), .B(n192), .Z(n194) );
  IV U222 ( .A(a[84]), .Z(n195) );
  NOR U223 ( .A(n194), .B(n195), .Z(n196) );
  NOR U224 ( .A(n193), .B(n196), .Z(n197) );
  IV U225 ( .A(n197), .Z(n1077) );
  IV U226 ( .A(n1081), .Z(n198) );
  IV U227 ( .A(b[87]), .Z(n199) );
  NOR U228 ( .A(n198), .B(n199), .Z(n200) );
  XOR U229 ( .A(n1081), .B(n199), .Z(n201) );
  IV U230 ( .A(a[87]), .Z(n202) );
  NOR U231 ( .A(n201), .B(n202), .Z(n203) );
  NOR U232 ( .A(n200), .B(n203), .Z(n204) );
  IV U233 ( .A(n204), .Z(n1083) );
  IV U234 ( .A(n1089), .Z(n205) );
  IV U235 ( .A(b[90]), .Z(n206) );
  NOR U236 ( .A(n205), .B(n206), .Z(n207) );
  XOR U237 ( .A(n1089), .B(n206), .Z(n208) );
  IV U238 ( .A(a[90]), .Z(n209) );
  NOR U239 ( .A(n208), .B(n209), .Z(n210) );
  NOR U240 ( .A(n207), .B(n210), .Z(n211) );
  IV U241 ( .A(n211), .Z(n1091) );
  IV U242 ( .A(n1095), .Z(n212) );
  IV U243 ( .A(b[93]), .Z(n213) );
  NOR U244 ( .A(n212), .B(n213), .Z(n214) );
  XOR U245 ( .A(n1095), .B(n213), .Z(n215) );
  IV U246 ( .A(a[93]), .Z(n216) );
  NOR U247 ( .A(n215), .B(n216), .Z(n217) );
  NOR U248 ( .A(n214), .B(n217), .Z(n218) );
  IV U249 ( .A(n218), .Z(n1097) );
  IV U250 ( .A(n1101), .Z(n219) );
  IV U251 ( .A(b[96]), .Z(n220) );
  NOR U252 ( .A(n219), .B(n220), .Z(n221) );
  XOR U253 ( .A(n1101), .B(n220), .Z(n222) );
  IV U254 ( .A(a[96]), .Z(n223) );
  NOR U255 ( .A(n222), .B(n223), .Z(n224) );
  NOR U256 ( .A(n221), .B(n224), .Z(n225) );
  IV U257 ( .A(n225), .Z(n1103) );
  IV U258 ( .A(n1107), .Z(n226) );
  IV U259 ( .A(a[99]), .Z(n227) );
  NOR U260 ( .A(n226), .B(n227), .Z(n228) );
  XOR U261 ( .A(n1107), .B(n227), .Z(n229) );
  IV U262 ( .A(b[99]), .Z(n230) );
  NOR U263 ( .A(n229), .B(n230), .Z(n231) );
  NOR U264 ( .A(n228), .B(n231), .Z(n232) );
  IV U265 ( .A(n232), .Z(n816) );
  IV U266 ( .A(n820), .Z(n233) );
  IV U267 ( .A(b[102]), .Z(n234) );
  NOR U268 ( .A(n233), .B(n234), .Z(n235) );
  XOR U269 ( .A(n820), .B(n234), .Z(n236) );
  IV U270 ( .A(a[102]), .Z(n237) );
  NOR U271 ( .A(n236), .B(n237), .Z(n238) );
  NOR U272 ( .A(n235), .B(n238), .Z(n239) );
  IV U273 ( .A(n239), .Z(n822) );
  IV U274 ( .A(n826), .Z(n240) );
  IV U275 ( .A(b[105]), .Z(n241) );
  NOR U276 ( .A(n240), .B(n241), .Z(n242) );
  XOR U277 ( .A(n826), .B(n241), .Z(n243) );
  IV U278 ( .A(a[105]), .Z(n244) );
  NOR U279 ( .A(n243), .B(n244), .Z(n245) );
  NOR U280 ( .A(n242), .B(n245), .Z(n246) );
  IV U281 ( .A(n246), .Z(n828) );
  IV U282 ( .A(n832), .Z(n247) );
  IV U283 ( .A(b[108]), .Z(n248) );
  NOR U284 ( .A(n247), .B(n248), .Z(n249) );
  XOR U285 ( .A(n832), .B(n248), .Z(n250) );
  IV U286 ( .A(a[108]), .Z(n251) );
  NOR U287 ( .A(n250), .B(n251), .Z(n252) );
  NOR U288 ( .A(n249), .B(n252), .Z(n253) );
  IV U289 ( .A(n253), .Z(n836) );
  IV U290 ( .A(n840), .Z(n254) );
  IV U291 ( .A(b[111]), .Z(n255) );
  NOR U292 ( .A(n254), .B(n255), .Z(n256) );
  XOR U293 ( .A(n840), .B(n255), .Z(n257) );
  IV U294 ( .A(a[111]), .Z(n258) );
  NOR U295 ( .A(n257), .B(n258), .Z(n259) );
  NOR U296 ( .A(n256), .B(n259), .Z(n260) );
  IV U297 ( .A(n260), .Z(n842) );
  IV U298 ( .A(n846), .Z(n261) );
  IV U299 ( .A(b[114]), .Z(n262) );
  NOR U300 ( .A(n261), .B(n262), .Z(n263) );
  XOR U301 ( .A(n846), .B(n262), .Z(n264) );
  IV U302 ( .A(a[114]), .Z(n265) );
  NOR U303 ( .A(n264), .B(n265), .Z(n266) );
  NOR U304 ( .A(n263), .B(n266), .Z(n267) );
  IV U305 ( .A(n267), .Z(n848) );
  IV U306 ( .A(n999), .Z(n268) );
  IV U307 ( .A(b[4]), .Z(n269) );
  NOR U308 ( .A(n268), .B(n269), .Z(n270) );
  XOR U309 ( .A(n999), .B(n269), .Z(n271) );
  IV U310 ( .A(a[4]), .Z(n272) );
  NOR U311 ( .A(n271), .B(n272), .Z(n273) );
  NOR U312 ( .A(n270), .B(n273), .Z(n274) );
  IV U313 ( .A(n274), .Z(n1021) );
  IV U314 ( .A(n1065), .Z(n275) );
  IV U315 ( .A(b[7]), .Z(n276) );
  NOR U316 ( .A(n275), .B(n276), .Z(n277) );
  XOR U317 ( .A(n1065), .B(n276), .Z(n278) );
  IV U318 ( .A(a[7]), .Z(n279) );
  NOR U319 ( .A(n278), .B(n279), .Z(n280) );
  NOR U320 ( .A(n277), .B(n280), .Z(n281) );
  IV U321 ( .A(n281), .Z(n1087) );
  IV U322 ( .A(n834), .Z(n282) );
  IV U323 ( .A(b[10]), .Z(n283) );
  NOR U324 ( .A(n282), .B(n283), .Z(n284) );
  XOR U325 ( .A(n834), .B(n283), .Z(n285) );
  IV U326 ( .A(a[10]), .Z(n286) );
  NOR U327 ( .A(n285), .B(n286), .Z(n287) );
  NOR U328 ( .A(n284), .B(n287), .Z(n288) );
  IV U329 ( .A(n288), .Z(n865) );
  IV U330 ( .A(n918), .Z(n289) );
  IV U331 ( .A(b[13]), .Z(n290) );
  NOR U332 ( .A(n289), .B(n290), .Z(n291) );
  XOR U333 ( .A(n918), .B(n290), .Z(n292) );
  IV U334 ( .A(a[13]), .Z(n293) );
  NOR U335 ( .A(n292), .B(n293), .Z(n294) );
  NOR U336 ( .A(n291), .B(n294), .Z(n295) );
  IV U337 ( .A(n295), .Z(n920) );
  IV U338 ( .A(n924), .Z(n296) );
  IV U339 ( .A(b[16]), .Z(n297) );
  NOR U340 ( .A(n296), .B(n297), .Z(n298) );
  XOR U341 ( .A(n924), .B(n297), .Z(n299) );
  IV U342 ( .A(a[16]), .Z(n300) );
  NOR U343 ( .A(n299), .B(n300), .Z(n301) );
  NOR U344 ( .A(n298), .B(n301), .Z(n302) );
  IV U345 ( .A(n302), .Z(n926) );
  IV U346 ( .A(n930), .Z(n303) );
  IV U347 ( .A(b[19]), .Z(n304) );
  NOR U348 ( .A(n303), .B(n304), .Z(n305) );
  XOR U349 ( .A(n930), .B(n304), .Z(n306) );
  IV U350 ( .A(a[19]), .Z(n307) );
  NOR U351 ( .A(n306), .B(n307), .Z(n308) );
  NOR U352 ( .A(n305), .B(n308), .Z(n309) );
  IV U353 ( .A(n309), .Z(n934) );
  IV U354 ( .A(n938), .Z(n310) );
  IV U355 ( .A(b[22]), .Z(n311) );
  NOR U356 ( .A(n310), .B(n311), .Z(n312) );
  XOR U357 ( .A(n938), .B(n311), .Z(n313) );
  IV U358 ( .A(a[22]), .Z(n314) );
  NOR U359 ( .A(n313), .B(n314), .Z(n315) );
  NOR U360 ( .A(n312), .B(n315), .Z(n316) );
  IV U361 ( .A(n316), .Z(n940) );
  IV U362 ( .A(n944), .Z(n317) );
  IV U363 ( .A(b[25]), .Z(n318) );
  NOR U364 ( .A(n317), .B(n318), .Z(n319) );
  XOR U365 ( .A(n944), .B(n318), .Z(n320) );
  IV U366 ( .A(a[25]), .Z(n321) );
  NOR U367 ( .A(n320), .B(n321), .Z(n322) );
  NOR U368 ( .A(n319), .B(n322), .Z(n323) );
  IV U369 ( .A(n323), .Z(n946) );
  IV U370 ( .A(n950), .Z(n324) );
  IV U371 ( .A(b[28]), .Z(n325) );
  NOR U372 ( .A(n324), .B(n325), .Z(n326) );
  XOR U373 ( .A(n950), .B(n325), .Z(n327) );
  IV U374 ( .A(a[28]), .Z(n328) );
  NOR U375 ( .A(n327), .B(n328), .Z(n329) );
  NOR U376 ( .A(n326), .B(n329), .Z(n330) );
  IV U377 ( .A(n330), .Z(n952) );
  IV U378 ( .A(n959), .Z(n331) );
  IV U379 ( .A(b[31]), .Z(n332) );
  NOR U380 ( .A(n331), .B(n332), .Z(n333) );
  XOR U381 ( .A(n959), .B(n332), .Z(n334) );
  IV U382 ( .A(a[31]), .Z(n335) );
  NOR U383 ( .A(n334), .B(n335), .Z(n336) );
  NOR U384 ( .A(n333), .B(n336), .Z(n337) );
  IV U385 ( .A(n337), .Z(n961) );
  IV U386 ( .A(n965), .Z(n338) );
  IV U387 ( .A(b[34]), .Z(n339) );
  NOR U388 ( .A(n338), .B(n339), .Z(n340) );
  XOR U389 ( .A(n965), .B(n339), .Z(n341) );
  IV U390 ( .A(a[34]), .Z(n342) );
  NOR U391 ( .A(n341), .B(n342), .Z(n343) );
  NOR U392 ( .A(n340), .B(n343), .Z(n344) );
  IV U393 ( .A(n344), .Z(n967) );
  IV U394 ( .A(n971), .Z(n345) );
  IV U395 ( .A(b[37]), .Z(n346) );
  NOR U396 ( .A(n345), .B(n346), .Z(n347) );
  XOR U397 ( .A(n971), .B(n346), .Z(n348) );
  IV U398 ( .A(a[37]), .Z(n349) );
  NOR U399 ( .A(n348), .B(n349), .Z(n350) );
  NOR U400 ( .A(n347), .B(n350), .Z(n351) );
  IV U401 ( .A(n351), .Z(n973) );
  IV U402 ( .A(n979), .Z(n352) );
  IV U403 ( .A(b[40]), .Z(n353) );
  NOR U404 ( .A(n352), .B(n353), .Z(n354) );
  XOR U405 ( .A(n979), .B(n353), .Z(n355) );
  IV U406 ( .A(a[40]), .Z(n356) );
  NOR U407 ( .A(n355), .B(n356), .Z(n357) );
  NOR U408 ( .A(n354), .B(n357), .Z(n358) );
  IV U409 ( .A(n358), .Z(n981) );
  IV U410 ( .A(n985), .Z(n359) );
  IV U411 ( .A(b[43]), .Z(n360) );
  NOR U412 ( .A(n359), .B(n360), .Z(n361) );
  XOR U413 ( .A(n985), .B(n360), .Z(n362) );
  IV U414 ( .A(a[43]), .Z(n363) );
  NOR U415 ( .A(n362), .B(n363), .Z(n364) );
  NOR U416 ( .A(n361), .B(n364), .Z(n365) );
  IV U417 ( .A(n365), .Z(n987) );
  IV U418 ( .A(n991), .Z(n366) );
  IV U419 ( .A(b[46]), .Z(n367) );
  NOR U420 ( .A(n366), .B(n367), .Z(n368) );
  XOR U421 ( .A(n991), .B(n367), .Z(n369) );
  IV U422 ( .A(a[46]), .Z(n370) );
  NOR U423 ( .A(n369), .B(n370), .Z(n371) );
  NOR U424 ( .A(n368), .B(n371), .Z(n372) );
  IV U425 ( .A(n372), .Z(n993) );
  IV U426 ( .A(n997), .Z(n373) );
  IV U427 ( .A(b[49]), .Z(n374) );
  NOR U428 ( .A(n373), .B(n374), .Z(n375) );
  XOR U429 ( .A(n997), .B(n374), .Z(n376) );
  IV U430 ( .A(a[49]), .Z(n377) );
  NOR U431 ( .A(n376), .B(n377), .Z(n378) );
  NOR U432 ( .A(n375), .B(n378), .Z(n379) );
  IV U433 ( .A(n379), .Z(n1001) );
  IV U434 ( .A(n1005), .Z(n380) );
  IV U435 ( .A(b[52]), .Z(n381) );
  NOR U436 ( .A(n380), .B(n381), .Z(n382) );
  XOR U437 ( .A(n1005), .B(n381), .Z(n383) );
  IV U438 ( .A(a[52]), .Z(n384) );
  NOR U439 ( .A(n383), .B(n384), .Z(n385) );
  NOR U440 ( .A(n382), .B(n385), .Z(n386) );
  IV U441 ( .A(n386), .Z(n1007) );
  IV U442 ( .A(n1011), .Z(n387) );
  IV U443 ( .A(b[55]), .Z(n388) );
  NOR U444 ( .A(n387), .B(n388), .Z(n389) );
  XOR U445 ( .A(n1011), .B(n388), .Z(n390) );
  IV U446 ( .A(a[55]), .Z(n391) );
  NOR U447 ( .A(n390), .B(n391), .Z(n392) );
  NOR U448 ( .A(n389), .B(n392), .Z(n393) );
  IV U449 ( .A(n393), .Z(n1013) );
  IV U450 ( .A(n1017), .Z(n394) );
  IV U451 ( .A(b[58]), .Z(n395) );
  NOR U452 ( .A(n394), .B(n395), .Z(n396) );
  XOR U453 ( .A(n1017), .B(n395), .Z(n397) );
  IV U454 ( .A(a[58]), .Z(n398) );
  NOR U455 ( .A(n397), .B(n398), .Z(n399) );
  NOR U456 ( .A(n396), .B(n399), .Z(n400) );
  IV U457 ( .A(n400), .Z(n1019) );
  IV U458 ( .A(n1025), .Z(n401) );
  IV U459 ( .A(b[61]), .Z(n402) );
  NOR U460 ( .A(n401), .B(n402), .Z(n403) );
  XOR U461 ( .A(n1025), .B(n402), .Z(n404) );
  IV U462 ( .A(a[61]), .Z(n405) );
  NOR U463 ( .A(n404), .B(n405), .Z(n406) );
  NOR U464 ( .A(n403), .B(n406), .Z(n407) );
  IV U465 ( .A(n407), .Z(n1027) );
  IV U466 ( .A(n1031), .Z(n408) );
  IV U467 ( .A(b[64]), .Z(n409) );
  NOR U468 ( .A(n408), .B(n409), .Z(n410) );
  XOR U469 ( .A(n1031), .B(n409), .Z(n411) );
  IV U470 ( .A(a[64]), .Z(n412) );
  NOR U471 ( .A(n411), .B(n412), .Z(n413) );
  NOR U472 ( .A(n410), .B(n413), .Z(n414) );
  IV U473 ( .A(n414), .Z(n1033) );
  IV U474 ( .A(n1037), .Z(n415) );
  IV U475 ( .A(b[67]), .Z(n416) );
  NOR U476 ( .A(n415), .B(n416), .Z(n417) );
  XOR U477 ( .A(n1037), .B(n416), .Z(n418) );
  IV U478 ( .A(a[67]), .Z(n419) );
  NOR U479 ( .A(n418), .B(n419), .Z(n420) );
  NOR U480 ( .A(n417), .B(n420), .Z(n421) );
  IV U481 ( .A(n421), .Z(n1039) );
  IV U482 ( .A(n1045), .Z(n422) );
  IV U483 ( .A(b[70]), .Z(n423) );
  NOR U484 ( .A(n422), .B(n423), .Z(n424) );
  XOR U485 ( .A(n1045), .B(n423), .Z(n425) );
  IV U486 ( .A(a[70]), .Z(n426) );
  NOR U487 ( .A(n425), .B(n426), .Z(n427) );
  NOR U488 ( .A(n424), .B(n427), .Z(n428) );
  IV U489 ( .A(n428), .Z(n1047) );
  IV U490 ( .A(n1051), .Z(n429) );
  IV U491 ( .A(b[73]), .Z(n430) );
  NOR U492 ( .A(n429), .B(n430), .Z(n431) );
  XOR U493 ( .A(n1051), .B(n430), .Z(n432) );
  IV U494 ( .A(a[73]), .Z(n433) );
  NOR U495 ( .A(n432), .B(n433), .Z(n434) );
  NOR U496 ( .A(n431), .B(n434), .Z(n435) );
  IV U497 ( .A(n435), .Z(n1053) );
  IV U498 ( .A(n1057), .Z(n436) );
  IV U499 ( .A(b[76]), .Z(n437) );
  NOR U500 ( .A(n436), .B(n437), .Z(n438) );
  XOR U501 ( .A(n1057), .B(n437), .Z(n439) );
  IV U502 ( .A(a[76]), .Z(n440) );
  NOR U503 ( .A(n439), .B(n440), .Z(n441) );
  NOR U504 ( .A(n438), .B(n441), .Z(n442) );
  IV U505 ( .A(n442), .Z(n1059) );
  IV U506 ( .A(n1063), .Z(n443) );
  IV U507 ( .A(b[79]), .Z(n444) );
  NOR U508 ( .A(n443), .B(n444), .Z(n445) );
  XOR U509 ( .A(n1063), .B(n444), .Z(n446) );
  IV U510 ( .A(a[79]), .Z(n447) );
  NOR U511 ( .A(n446), .B(n447), .Z(n448) );
  NOR U512 ( .A(n445), .B(n448), .Z(n449) );
  IV U513 ( .A(n449), .Z(n1067) );
  IV U514 ( .A(n1071), .Z(n450) );
  IV U515 ( .A(b[82]), .Z(n451) );
  NOR U516 ( .A(n450), .B(n451), .Z(n452) );
  XOR U517 ( .A(n1071), .B(n451), .Z(n453) );
  IV U518 ( .A(a[82]), .Z(n454) );
  NOR U519 ( .A(n453), .B(n454), .Z(n455) );
  NOR U520 ( .A(n452), .B(n455), .Z(n456) );
  IV U521 ( .A(n456), .Z(n1073) );
  IV U522 ( .A(n1077), .Z(n457) );
  IV U523 ( .A(b[85]), .Z(n458) );
  NOR U524 ( .A(n457), .B(n458), .Z(n459) );
  XOR U525 ( .A(n1077), .B(n458), .Z(n460) );
  IV U526 ( .A(a[85]), .Z(n461) );
  NOR U527 ( .A(n460), .B(n461), .Z(n462) );
  NOR U528 ( .A(n459), .B(n462), .Z(n463) );
  IV U529 ( .A(n463), .Z(n1079) );
  IV U530 ( .A(n1083), .Z(n464) );
  IV U531 ( .A(b[88]), .Z(n465) );
  NOR U532 ( .A(n464), .B(n465), .Z(n466) );
  XOR U533 ( .A(n1083), .B(n465), .Z(n467) );
  IV U534 ( .A(a[88]), .Z(n468) );
  NOR U535 ( .A(n467), .B(n468), .Z(n469) );
  NOR U536 ( .A(n466), .B(n469), .Z(n470) );
  IV U537 ( .A(n470), .Z(n1085) );
  IV U538 ( .A(n1091), .Z(n471) );
  IV U539 ( .A(b[91]), .Z(n472) );
  NOR U540 ( .A(n471), .B(n472), .Z(n473) );
  XOR U541 ( .A(n1091), .B(n472), .Z(n474) );
  IV U542 ( .A(a[91]), .Z(n475) );
  NOR U543 ( .A(n474), .B(n475), .Z(n476) );
  NOR U544 ( .A(n473), .B(n476), .Z(n477) );
  IV U545 ( .A(n477), .Z(n1093) );
  IV U546 ( .A(n1097), .Z(n478) );
  IV U547 ( .A(b[94]), .Z(n479) );
  NOR U548 ( .A(n478), .B(n479), .Z(n480) );
  XOR U549 ( .A(n1097), .B(n479), .Z(n481) );
  IV U550 ( .A(a[94]), .Z(n482) );
  NOR U551 ( .A(n481), .B(n482), .Z(n483) );
  NOR U552 ( .A(n480), .B(n483), .Z(n484) );
  IV U553 ( .A(n484), .Z(n1099) );
  IV U554 ( .A(n1103), .Z(n485) );
  IV U555 ( .A(b[97]), .Z(n486) );
  NOR U556 ( .A(n485), .B(n486), .Z(n487) );
  XOR U557 ( .A(n1103), .B(n486), .Z(n488) );
  IV U558 ( .A(a[97]), .Z(n489) );
  NOR U559 ( .A(n488), .B(n489), .Z(n490) );
  NOR U560 ( .A(n487), .B(n490), .Z(n491) );
  IV U561 ( .A(n491), .Z(n1105) );
  IV U562 ( .A(n816), .Z(n492) );
  IV U563 ( .A(b[100]), .Z(n493) );
  NOR U564 ( .A(n492), .B(n493), .Z(n494) );
  XOR U565 ( .A(n816), .B(n493), .Z(n495) );
  IV U566 ( .A(a[100]), .Z(n496) );
  NOR U567 ( .A(n495), .B(n496), .Z(n497) );
  NOR U568 ( .A(n494), .B(n497), .Z(n498) );
  IV U569 ( .A(n498), .Z(n818) );
  IV U570 ( .A(n822), .Z(n499) );
  IV U571 ( .A(b[103]), .Z(n500) );
  NOR U572 ( .A(n499), .B(n500), .Z(n501) );
  XOR U573 ( .A(n822), .B(n500), .Z(n502) );
  IV U574 ( .A(a[103]), .Z(n503) );
  NOR U575 ( .A(n502), .B(n503), .Z(n504) );
  NOR U576 ( .A(n501), .B(n504), .Z(n505) );
  IV U577 ( .A(n505), .Z(n824) );
  IV U578 ( .A(n828), .Z(n506) );
  IV U579 ( .A(b[106]), .Z(n507) );
  NOR U580 ( .A(n506), .B(n507), .Z(n508) );
  XOR U581 ( .A(n828), .B(n507), .Z(n509) );
  IV U582 ( .A(a[106]), .Z(n510) );
  NOR U583 ( .A(n509), .B(n510), .Z(n511) );
  NOR U584 ( .A(n508), .B(n511), .Z(n512) );
  IV U585 ( .A(n512), .Z(n830) );
  IV U586 ( .A(n836), .Z(n513) );
  IV U587 ( .A(b[109]), .Z(n514) );
  NOR U588 ( .A(n513), .B(n514), .Z(n515) );
  XOR U589 ( .A(n836), .B(n514), .Z(n516) );
  IV U590 ( .A(a[109]), .Z(n517) );
  NOR U591 ( .A(n516), .B(n517), .Z(n518) );
  NOR U592 ( .A(n515), .B(n518), .Z(n519) );
  IV U593 ( .A(n519), .Z(n838) );
  IV U594 ( .A(n842), .Z(n520) );
  IV U595 ( .A(b[112]), .Z(n521) );
  NOR U596 ( .A(n520), .B(n521), .Z(n522) );
  XOR U597 ( .A(n842), .B(n521), .Z(n523) );
  IV U598 ( .A(a[112]), .Z(n524) );
  NOR U599 ( .A(n523), .B(n524), .Z(n525) );
  NOR U600 ( .A(n522), .B(n525), .Z(n526) );
  IV U601 ( .A(n526), .Z(n844) );
  IV U602 ( .A(n848), .Z(n527) );
  IV U603 ( .A(b[115]), .Z(n528) );
  NOR U604 ( .A(n527), .B(n528), .Z(n529) );
  XOR U605 ( .A(n848), .B(n528), .Z(n530) );
  IV U606 ( .A(a[115]), .Z(n531) );
  NOR U607 ( .A(n530), .B(n531), .Z(n532) );
  NOR U608 ( .A(n529), .B(n532), .Z(n533) );
  IV U609 ( .A(n533), .Z(n850) );
  IV U610 ( .A(n1021), .Z(n534) );
  IV U611 ( .A(b[5]), .Z(n535) );
  NOR U612 ( .A(n534), .B(n535), .Z(n536) );
  XOR U613 ( .A(n1021), .B(n535), .Z(n537) );
  IV U614 ( .A(a[5]), .Z(n538) );
  NOR U615 ( .A(n537), .B(n538), .Z(n539) );
  NOR U616 ( .A(n536), .B(n539), .Z(n540) );
  IV U617 ( .A(n540), .Z(n1043) );
  IV U618 ( .A(n1087), .Z(n541) );
  IV U619 ( .A(b[8]), .Z(n542) );
  NOR U620 ( .A(n541), .B(n542), .Z(n543) );
  XOR U621 ( .A(n1087), .B(n542), .Z(n544) );
  IV U622 ( .A(a[8]), .Z(n545) );
  NOR U623 ( .A(n544), .B(n545), .Z(n546) );
  NOR U624 ( .A(n543), .B(n546), .Z(n547) );
  IV U625 ( .A(n547), .Z(n1109) );
  IV U626 ( .A(n865), .Z(n548) );
  IV U627 ( .A(b[11]), .Z(n549) );
  NOR U628 ( .A(n548), .B(n549), .Z(n550) );
  XOR U629 ( .A(n865), .B(n549), .Z(n551) );
  IV U630 ( .A(a[11]), .Z(n552) );
  NOR U631 ( .A(n551), .B(n552), .Z(n553) );
  NOR U632 ( .A(n550), .B(n553), .Z(n554) );
  IV U633 ( .A(n554), .Z(n916) );
  IV U634 ( .A(n920), .Z(n555) );
  IV U635 ( .A(b[14]), .Z(n556) );
  NOR U636 ( .A(n555), .B(n556), .Z(n557) );
  XOR U637 ( .A(n920), .B(n556), .Z(n558) );
  IV U638 ( .A(a[14]), .Z(n559) );
  NOR U639 ( .A(n558), .B(n559), .Z(n560) );
  NOR U640 ( .A(n557), .B(n560), .Z(n561) );
  IV U641 ( .A(n561), .Z(n922) );
  IV U642 ( .A(n926), .Z(n562) );
  IV U643 ( .A(b[17]), .Z(n563) );
  NOR U644 ( .A(n562), .B(n563), .Z(n564) );
  XOR U645 ( .A(n926), .B(n563), .Z(n565) );
  IV U646 ( .A(a[17]), .Z(n566) );
  NOR U647 ( .A(n565), .B(n566), .Z(n567) );
  NOR U648 ( .A(n564), .B(n567), .Z(n568) );
  IV U649 ( .A(n568), .Z(n928) );
  IV U650 ( .A(n934), .Z(n569) );
  IV U651 ( .A(b[20]), .Z(n570) );
  NOR U652 ( .A(n569), .B(n570), .Z(n571) );
  XOR U653 ( .A(n934), .B(n570), .Z(n572) );
  IV U654 ( .A(a[20]), .Z(n573) );
  NOR U655 ( .A(n572), .B(n573), .Z(n574) );
  NOR U656 ( .A(n571), .B(n574), .Z(n575) );
  IV U657 ( .A(n575), .Z(n936) );
  IV U658 ( .A(n940), .Z(n576) );
  IV U659 ( .A(b[23]), .Z(n577) );
  NOR U660 ( .A(n576), .B(n577), .Z(n578) );
  XOR U661 ( .A(n940), .B(n577), .Z(n579) );
  IV U662 ( .A(a[23]), .Z(n580) );
  NOR U663 ( .A(n579), .B(n580), .Z(n581) );
  NOR U664 ( .A(n578), .B(n581), .Z(n582) );
  IV U665 ( .A(n582), .Z(n942) );
  IV U666 ( .A(n946), .Z(n583) );
  IV U667 ( .A(b[26]), .Z(n584) );
  NOR U668 ( .A(n583), .B(n584), .Z(n585) );
  XOR U669 ( .A(n946), .B(n584), .Z(n586) );
  IV U670 ( .A(a[26]), .Z(n587) );
  NOR U671 ( .A(n586), .B(n587), .Z(n588) );
  NOR U672 ( .A(n585), .B(n588), .Z(n589) );
  IV U673 ( .A(n589), .Z(n948) );
  IV U674 ( .A(n952), .Z(n590) );
  IV U675 ( .A(b[29]), .Z(n591) );
  NOR U676 ( .A(n590), .B(n591), .Z(n592) );
  XOR U677 ( .A(n952), .B(n591), .Z(n593) );
  IV U678 ( .A(a[29]), .Z(n594) );
  NOR U679 ( .A(n593), .B(n594), .Z(n595) );
  NOR U680 ( .A(n592), .B(n595), .Z(n596) );
  IV U681 ( .A(n596), .Z(n957) );
  IV U682 ( .A(n961), .Z(n597) );
  IV U683 ( .A(b[32]), .Z(n598) );
  NOR U684 ( .A(n597), .B(n598), .Z(n599) );
  XOR U685 ( .A(n961), .B(n598), .Z(n600) );
  IV U686 ( .A(a[32]), .Z(n601) );
  NOR U687 ( .A(n600), .B(n601), .Z(n602) );
  NOR U688 ( .A(n599), .B(n602), .Z(n603) );
  IV U689 ( .A(n603), .Z(n963) );
  IV U690 ( .A(n967), .Z(n604) );
  IV U691 ( .A(b[35]), .Z(n605) );
  NOR U692 ( .A(n604), .B(n605), .Z(n606) );
  XOR U693 ( .A(n967), .B(n605), .Z(n607) );
  IV U694 ( .A(a[35]), .Z(n608) );
  NOR U695 ( .A(n607), .B(n608), .Z(n609) );
  NOR U696 ( .A(n606), .B(n609), .Z(n610) );
  IV U697 ( .A(n610), .Z(n969) );
  IV U698 ( .A(n973), .Z(n611) );
  IV U699 ( .A(b[38]), .Z(n612) );
  NOR U700 ( .A(n611), .B(n612), .Z(n613) );
  XOR U701 ( .A(n973), .B(n612), .Z(n614) );
  IV U702 ( .A(a[38]), .Z(n615) );
  NOR U703 ( .A(n614), .B(n615), .Z(n616) );
  NOR U704 ( .A(n613), .B(n616), .Z(n617) );
  IV U705 ( .A(n617), .Z(n975) );
  IV U706 ( .A(n981), .Z(n618) );
  IV U707 ( .A(b[41]), .Z(n619) );
  NOR U708 ( .A(n618), .B(n619), .Z(n620) );
  XOR U709 ( .A(n981), .B(n619), .Z(n621) );
  IV U710 ( .A(a[41]), .Z(n622) );
  NOR U711 ( .A(n621), .B(n622), .Z(n623) );
  NOR U712 ( .A(n620), .B(n623), .Z(n624) );
  IV U713 ( .A(n624), .Z(n983) );
  IV U714 ( .A(n987), .Z(n625) );
  IV U715 ( .A(b[44]), .Z(n626) );
  NOR U716 ( .A(n625), .B(n626), .Z(n627) );
  XOR U717 ( .A(n987), .B(n626), .Z(n628) );
  IV U718 ( .A(a[44]), .Z(n629) );
  NOR U719 ( .A(n628), .B(n629), .Z(n630) );
  NOR U720 ( .A(n627), .B(n630), .Z(n631) );
  IV U721 ( .A(n631), .Z(n989) );
  IV U722 ( .A(n993), .Z(n632) );
  IV U723 ( .A(b[47]), .Z(n633) );
  NOR U724 ( .A(n632), .B(n633), .Z(n634) );
  XOR U725 ( .A(n993), .B(n633), .Z(n635) );
  IV U726 ( .A(a[47]), .Z(n636) );
  NOR U727 ( .A(n635), .B(n636), .Z(n637) );
  NOR U728 ( .A(n634), .B(n637), .Z(n638) );
  IV U729 ( .A(n638), .Z(n995) );
  IV U730 ( .A(n1001), .Z(n639) );
  IV U731 ( .A(b[50]), .Z(n640) );
  NOR U732 ( .A(n639), .B(n640), .Z(n641) );
  XOR U733 ( .A(n1001), .B(n640), .Z(n642) );
  IV U734 ( .A(a[50]), .Z(n643) );
  NOR U735 ( .A(n642), .B(n643), .Z(n644) );
  NOR U736 ( .A(n641), .B(n644), .Z(n645) );
  IV U737 ( .A(n645), .Z(n1003) );
  IV U738 ( .A(n1007), .Z(n646) );
  IV U739 ( .A(b[53]), .Z(n647) );
  NOR U740 ( .A(n646), .B(n647), .Z(n648) );
  XOR U741 ( .A(n1007), .B(n647), .Z(n649) );
  IV U742 ( .A(a[53]), .Z(n650) );
  NOR U743 ( .A(n649), .B(n650), .Z(n651) );
  NOR U744 ( .A(n648), .B(n651), .Z(n652) );
  IV U745 ( .A(n652), .Z(n1009) );
  IV U746 ( .A(n1013), .Z(n653) );
  IV U747 ( .A(b[56]), .Z(n654) );
  NOR U748 ( .A(n653), .B(n654), .Z(n655) );
  XOR U749 ( .A(n1013), .B(n654), .Z(n656) );
  IV U750 ( .A(a[56]), .Z(n657) );
  NOR U751 ( .A(n656), .B(n657), .Z(n658) );
  NOR U752 ( .A(n655), .B(n658), .Z(n659) );
  IV U753 ( .A(n659), .Z(n1015) );
  IV U754 ( .A(n1019), .Z(n660) );
  IV U755 ( .A(b[59]), .Z(n661) );
  NOR U756 ( .A(n660), .B(n661), .Z(n662) );
  XOR U757 ( .A(n1019), .B(n661), .Z(n663) );
  IV U758 ( .A(a[59]), .Z(n664) );
  NOR U759 ( .A(n663), .B(n664), .Z(n665) );
  NOR U760 ( .A(n662), .B(n665), .Z(n666) );
  IV U761 ( .A(n666), .Z(n1023) );
  IV U762 ( .A(n1027), .Z(n667) );
  IV U763 ( .A(b[62]), .Z(n668) );
  NOR U764 ( .A(n667), .B(n668), .Z(n669) );
  XOR U765 ( .A(n1027), .B(n668), .Z(n670) );
  IV U766 ( .A(a[62]), .Z(n671) );
  NOR U767 ( .A(n670), .B(n671), .Z(n672) );
  NOR U768 ( .A(n669), .B(n672), .Z(n673) );
  IV U769 ( .A(n673), .Z(n1029) );
  IV U770 ( .A(n1033), .Z(n674) );
  IV U771 ( .A(b[65]), .Z(n675) );
  NOR U772 ( .A(n674), .B(n675), .Z(n676) );
  XOR U773 ( .A(n1033), .B(n675), .Z(n677) );
  IV U774 ( .A(a[65]), .Z(n678) );
  NOR U775 ( .A(n677), .B(n678), .Z(n679) );
  NOR U776 ( .A(n676), .B(n679), .Z(n680) );
  IV U777 ( .A(n680), .Z(n1035) );
  IV U778 ( .A(n1039), .Z(n681) );
  IV U779 ( .A(b[68]), .Z(n682) );
  NOR U780 ( .A(n681), .B(n682), .Z(n683) );
  XOR U781 ( .A(n1039), .B(n682), .Z(n684) );
  IV U782 ( .A(a[68]), .Z(n685) );
  NOR U783 ( .A(n684), .B(n685), .Z(n686) );
  NOR U784 ( .A(n683), .B(n686), .Z(n687) );
  IV U785 ( .A(n687), .Z(n1041) );
  IV U786 ( .A(n1047), .Z(n688) );
  IV U787 ( .A(b[71]), .Z(n689) );
  NOR U788 ( .A(n688), .B(n689), .Z(n690) );
  XOR U789 ( .A(n1047), .B(n689), .Z(n691) );
  IV U790 ( .A(a[71]), .Z(n692) );
  NOR U791 ( .A(n691), .B(n692), .Z(n693) );
  NOR U792 ( .A(n690), .B(n693), .Z(n694) );
  IV U793 ( .A(n694), .Z(n1049) );
  IV U794 ( .A(n1053), .Z(n695) );
  IV U795 ( .A(b[74]), .Z(n696) );
  NOR U796 ( .A(n695), .B(n696), .Z(n697) );
  XOR U797 ( .A(n1053), .B(n696), .Z(n698) );
  IV U798 ( .A(a[74]), .Z(n699) );
  NOR U799 ( .A(n698), .B(n699), .Z(n700) );
  NOR U800 ( .A(n697), .B(n700), .Z(n701) );
  IV U801 ( .A(n701), .Z(n1055) );
  IV U802 ( .A(n1059), .Z(n702) );
  IV U803 ( .A(b[77]), .Z(n703) );
  NOR U804 ( .A(n702), .B(n703), .Z(n704) );
  XOR U805 ( .A(n1059), .B(n703), .Z(n705) );
  IV U806 ( .A(a[77]), .Z(n706) );
  NOR U807 ( .A(n705), .B(n706), .Z(n707) );
  NOR U808 ( .A(n704), .B(n707), .Z(n708) );
  IV U809 ( .A(n708), .Z(n1061) );
  IV U810 ( .A(n1067), .Z(n709) );
  IV U811 ( .A(b[80]), .Z(n710) );
  NOR U812 ( .A(n709), .B(n710), .Z(n711) );
  XOR U813 ( .A(n1067), .B(n710), .Z(n712) );
  IV U814 ( .A(a[80]), .Z(n713) );
  NOR U815 ( .A(n712), .B(n713), .Z(n714) );
  NOR U816 ( .A(n711), .B(n714), .Z(n715) );
  IV U817 ( .A(n715), .Z(n1069) );
  IV U818 ( .A(n1073), .Z(n716) );
  IV U819 ( .A(b[83]), .Z(n717) );
  NOR U820 ( .A(n716), .B(n717), .Z(n718) );
  XOR U821 ( .A(n1073), .B(n717), .Z(n719) );
  IV U822 ( .A(a[83]), .Z(n720) );
  NOR U823 ( .A(n719), .B(n720), .Z(n721) );
  NOR U824 ( .A(n718), .B(n721), .Z(n722) );
  IV U825 ( .A(n722), .Z(n1075) );
  IV U826 ( .A(n1079), .Z(n723) );
  IV U827 ( .A(b[86]), .Z(n724) );
  NOR U828 ( .A(n723), .B(n724), .Z(n725) );
  XOR U829 ( .A(n1079), .B(n724), .Z(n726) );
  IV U830 ( .A(a[86]), .Z(n727) );
  NOR U831 ( .A(n726), .B(n727), .Z(n728) );
  NOR U832 ( .A(n725), .B(n728), .Z(n729) );
  IV U833 ( .A(n729), .Z(n1081) );
  IV U834 ( .A(n1085), .Z(n730) );
  IV U835 ( .A(b[89]), .Z(n731) );
  NOR U836 ( .A(n730), .B(n731), .Z(n732) );
  XOR U837 ( .A(n1085), .B(n731), .Z(n733) );
  IV U838 ( .A(a[89]), .Z(n734) );
  NOR U839 ( .A(n733), .B(n734), .Z(n735) );
  NOR U840 ( .A(n732), .B(n735), .Z(n736) );
  IV U841 ( .A(n736), .Z(n1089) );
  IV U842 ( .A(n1093), .Z(n737) );
  IV U843 ( .A(b[92]), .Z(n738) );
  NOR U844 ( .A(n737), .B(n738), .Z(n739) );
  XOR U845 ( .A(n1093), .B(n738), .Z(n740) );
  IV U846 ( .A(a[92]), .Z(n741) );
  NOR U847 ( .A(n740), .B(n741), .Z(n742) );
  NOR U848 ( .A(n739), .B(n742), .Z(n743) );
  IV U849 ( .A(n743), .Z(n1095) );
  IV U850 ( .A(n1099), .Z(n744) );
  IV U851 ( .A(b[95]), .Z(n745) );
  NOR U852 ( .A(n744), .B(n745), .Z(n746) );
  XOR U853 ( .A(n1099), .B(n745), .Z(n747) );
  IV U854 ( .A(a[95]), .Z(n748) );
  NOR U855 ( .A(n747), .B(n748), .Z(n749) );
  NOR U856 ( .A(n746), .B(n749), .Z(n750) );
  IV U857 ( .A(n750), .Z(n1101) );
  IV U858 ( .A(n1105), .Z(n751) );
  IV U859 ( .A(b[98]), .Z(n752) );
  NOR U860 ( .A(n751), .B(n752), .Z(n753) );
  XOR U861 ( .A(n1105), .B(n752), .Z(n754) );
  IV U862 ( .A(a[98]), .Z(n755) );
  NOR U863 ( .A(n754), .B(n755), .Z(n756) );
  NOR U864 ( .A(n753), .B(n756), .Z(n757) );
  IV U865 ( .A(n757), .Z(n1107) );
  IV U866 ( .A(n818), .Z(n758) );
  IV U867 ( .A(b[101]), .Z(n759) );
  NOR U868 ( .A(n758), .B(n759), .Z(n760) );
  XOR U869 ( .A(n818), .B(n759), .Z(n761) );
  IV U870 ( .A(a[101]), .Z(n762) );
  NOR U871 ( .A(n761), .B(n762), .Z(n763) );
  NOR U872 ( .A(n760), .B(n763), .Z(n764) );
  IV U873 ( .A(n764), .Z(n820) );
  IV U874 ( .A(n824), .Z(n765) );
  IV U875 ( .A(b[104]), .Z(n766) );
  NOR U876 ( .A(n765), .B(n766), .Z(n767) );
  XOR U877 ( .A(n824), .B(n766), .Z(n768) );
  IV U878 ( .A(a[104]), .Z(n769) );
  NOR U879 ( .A(n768), .B(n769), .Z(n770) );
  NOR U880 ( .A(n767), .B(n770), .Z(n771) );
  IV U881 ( .A(n771), .Z(n826) );
  IV U882 ( .A(n830), .Z(n772) );
  IV U883 ( .A(b[107]), .Z(n773) );
  NOR U884 ( .A(n772), .B(n773), .Z(n774) );
  XOR U885 ( .A(n830), .B(n773), .Z(n775) );
  IV U886 ( .A(a[107]), .Z(n776) );
  NOR U887 ( .A(n775), .B(n776), .Z(n777) );
  NOR U888 ( .A(n774), .B(n777), .Z(n778) );
  IV U889 ( .A(n778), .Z(n832) );
  IV U890 ( .A(n838), .Z(n779) );
  IV U891 ( .A(b[110]), .Z(n780) );
  NOR U892 ( .A(n779), .B(n780), .Z(n781) );
  XOR U893 ( .A(n838), .B(n780), .Z(n782) );
  IV U894 ( .A(a[110]), .Z(n783) );
  NOR U895 ( .A(n782), .B(n783), .Z(n784) );
  NOR U896 ( .A(n781), .B(n784), .Z(n785) );
  IV U897 ( .A(n785), .Z(n840) );
  IV U898 ( .A(n844), .Z(n786) );
  IV U899 ( .A(b[113]), .Z(n787) );
  NOR U900 ( .A(n786), .B(n787), .Z(n788) );
  XOR U901 ( .A(n844), .B(n787), .Z(n789) );
  IV U902 ( .A(a[113]), .Z(n790) );
  NOR U903 ( .A(n789), .B(n790), .Z(n791) );
  NOR U904 ( .A(n788), .B(n791), .Z(n792) );
  IV U905 ( .A(n792), .Z(n846) );
  IV U906 ( .A(b[116]), .Z(n793) );
  IV U907 ( .A(a[116]), .Z(n794) );
  IV U908 ( .A(n850), .Z(n795) );
  NOR U909 ( .A(n795), .B(n793), .Z(n796) );
  XOR U910 ( .A(n850), .B(n793), .Z(n797) );
  NOR U911 ( .A(n797), .B(n794), .Z(n798) );
  NOR U912 ( .A(n796), .B(n798), .Z(n799) );
  IV U913 ( .A(n799), .Z(n852) );
  IV U914 ( .A(a[127]), .Z(n800) );
  NOR U915 ( .A(a[127]), .B(n1112), .Z(n801) );
  NOR U916 ( .A(n1111), .B(n800), .Z(n802) );
  NOR U917 ( .A(b[127]), .B(n802), .Z(n803) );
  NOR U918 ( .A(n801), .B(n803), .Z(c[128]) );
  XOR U919 ( .A(a[0]), .B(b[0]), .Z(c[0]) );
  IV U920 ( .A(a[1]), .Z(n804) );
  IV U921 ( .A(b[1]), .Z(n805) );
  NOR U922 ( .A(n804), .B(n805), .Z(n810) );
  XOR U923 ( .A(a[1]), .B(n805), .Z(n933) );
  IV U924 ( .A(a[0]), .Z(n807) );
  IV U925 ( .A(b[0]), .Z(n806) );
  NOR U926 ( .A(n807), .B(n806), .Z(n808) );
  IV U927 ( .A(n808), .Z(n932) );
  NOR U928 ( .A(n933), .B(n932), .Z(n809) );
  NOR U929 ( .A(n810), .B(n809), .Z(n954) );
  IV U930 ( .A(n954), .Z(n811) );
  NOR U931 ( .A(a[2]), .B(n811), .Z(n814) );
  IV U932 ( .A(a[2]), .Z(n956) );
  NOR U933 ( .A(n954), .B(n956), .Z(n812) );
  NOR U934 ( .A(b[2]), .B(n812), .Z(n813) );
  NOR U935 ( .A(n814), .B(n813), .Z(n977) );
  XOR U936 ( .A(b[100]), .B(n816), .Z(n815) );
  XOR U937 ( .A(a[100]), .B(n815), .Z(c[100]) );
  XOR U938 ( .A(b[101]), .B(n818), .Z(n817) );
  XOR U939 ( .A(a[101]), .B(n817), .Z(c[101]) );
  XOR U940 ( .A(b[102]), .B(n820), .Z(n819) );
  XOR U941 ( .A(a[102]), .B(n819), .Z(c[102]) );
  XOR U942 ( .A(b[103]), .B(n822), .Z(n821) );
  XOR U943 ( .A(a[103]), .B(n821), .Z(c[103]) );
  XOR U944 ( .A(b[104]), .B(n824), .Z(n823) );
  XOR U945 ( .A(a[104]), .B(n823), .Z(c[104]) );
  XOR U946 ( .A(b[105]), .B(n826), .Z(n825) );
  XOR U947 ( .A(a[105]), .B(n825), .Z(c[105]) );
  XOR U948 ( .A(b[106]), .B(n828), .Z(n827) );
  XOR U949 ( .A(a[106]), .B(n827), .Z(c[106]) );
  XOR U950 ( .A(b[107]), .B(n830), .Z(n829) );
  XOR U951 ( .A(a[107]), .B(n829), .Z(c[107]) );
  XOR U952 ( .A(b[108]), .B(n832), .Z(n831) );
  XOR U953 ( .A(a[108]), .B(n831), .Z(c[108]) );
  XOR U954 ( .A(b[109]), .B(n836), .Z(n833) );
  XOR U955 ( .A(a[109]), .B(n833), .Z(c[109]) );
  XOR U956 ( .A(b[10]), .B(n834), .Z(n835) );
  XOR U957 ( .A(a[10]), .B(n835), .Z(c[10]) );
  XOR U958 ( .A(b[110]), .B(n838), .Z(n837) );
  XOR U959 ( .A(a[110]), .B(n837), .Z(c[110]) );
  XOR U960 ( .A(b[111]), .B(n840), .Z(n839) );
  XOR U961 ( .A(a[111]), .B(n839), .Z(c[111]) );
  XOR U962 ( .A(b[112]), .B(n842), .Z(n841) );
  XOR U963 ( .A(a[112]), .B(n841), .Z(c[112]) );
  XOR U964 ( .A(b[113]), .B(n844), .Z(n843) );
  XOR U965 ( .A(a[113]), .B(n843), .Z(c[113]) );
  XOR U966 ( .A(b[114]), .B(n846), .Z(n845) );
  XOR U967 ( .A(a[114]), .B(n845), .Z(c[114]) );
  XOR U968 ( .A(b[115]), .B(n848), .Z(n847) );
  XOR U969 ( .A(a[115]), .B(n847), .Z(c[115]) );
  XOR U970 ( .A(b[116]), .B(n850), .Z(n849) );
  XOR U971 ( .A(a[116]), .B(n849), .Z(c[116]) );
  XOR U972 ( .A(b[117]), .B(n852), .Z(n851) );
  XOR U973 ( .A(a[117]), .B(n851), .Z(c[117]) );
  IV U974 ( .A(a[118]), .Z(n859) );
  IV U975 ( .A(n852), .Z(n855) );
  XOR U976 ( .A(b[117]), .B(n855), .Z(n854) );
  IV U977 ( .A(a[117]), .Z(n853) );
  NOR U978 ( .A(n854), .B(n853), .Z(n858) );
  IV U979 ( .A(b[117]), .Z(n856) );
  NOR U980 ( .A(n856), .B(n855), .Z(n857) );
  NOR U981 ( .A(n858), .B(n857), .Z(n861) );
  XOR U982 ( .A(b[118]), .B(n861), .Z(n860) );
  XOR U983 ( .A(n859), .B(n860), .Z(c[118]) );
  IV U984 ( .A(a[119]), .Z(n867) );
  NOR U985 ( .A(n860), .B(n859), .Z(n864) );
  IV U986 ( .A(b[118]), .Z(n862) );
  NOR U987 ( .A(n862), .B(n861), .Z(n863) );
  NOR U988 ( .A(n864), .B(n863), .Z(n869) );
  XOR U989 ( .A(b[119]), .B(n869), .Z(n868) );
  XOR U990 ( .A(n867), .B(n868), .Z(c[119]) );
  XOR U991 ( .A(b[11]), .B(n865), .Z(n866) );
  XOR U992 ( .A(a[11]), .B(n866), .Z(c[11]) );
  IV U993 ( .A(a[120]), .Z(n873) );
  NOR U994 ( .A(n868), .B(n867), .Z(n872) );
  IV U995 ( .A(b[119]), .Z(n870) );
  NOR U996 ( .A(n870), .B(n869), .Z(n871) );
  NOR U997 ( .A(n872), .B(n871), .Z(n875) );
  XOR U998 ( .A(b[120]), .B(n875), .Z(n874) );
  XOR U999 ( .A(n873), .B(n874), .Z(c[120]) );
  IV U1000 ( .A(a[121]), .Z(n879) );
  NOR U1001 ( .A(n874), .B(n873), .Z(n878) );
  IV U1002 ( .A(b[120]), .Z(n876) );
  NOR U1003 ( .A(n876), .B(n875), .Z(n877) );
  NOR U1004 ( .A(n878), .B(n877), .Z(n881) );
  XOR U1005 ( .A(b[121]), .B(n881), .Z(n880) );
  XOR U1006 ( .A(n879), .B(n880), .Z(c[121]) );
  IV U1007 ( .A(a[122]), .Z(n885) );
  NOR U1008 ( .A(n880), .B(n879), .Z(n884) );
  IV U1009 ( .A(b[121]), .Z(n882) );
  NOR U1010 ( .A(n882), .B(n881), .Z(n883) );
  NOR U1011 ( .A(n884), .B(n883), .Z(n887) );
  XOR U1012 ( .A(b[122]), .B(n887), .Z(n886) );
  XOR U1013 ( .A(n885), .B(n886), .Z(c[122]) );
  IV U1014 ( .A(a[123]), .Z(n891) );
  NOR U1015 ( .A(n886), .B(n885), .Z(n890) );
  IV U1016 ( .A(b[122]), .Z(n888) );
  NOR U1017 ( .A(n888), .B(n887), .Z(n889) );
  NOR U1018 ( .A(n890), .B(n889), .Z(n893) );
  XOR U1019 ( .A(b[123]), .B(n893), .Z(n892) );
  XOR U1020 ( .A(n891), .B(n892), .Z(c[123]) );
  IV U1021 ( .A(a[124]), .Z(n897) );
  NOR U1022 ( .A(n892), .B(n891), .Z(n896) );
  IV U1023 ( .A(b[123]), .Z(n894) );
  NOR U1024 ( .A(n894), .B(n893), .Z(n895) );
  NOR U1025 ( .A(n896), .B(n895), .Z(n899) );
  XOR U1026 ( .A(b[124]), .B(n899), .Z(n898) );
  XOR U1027 ( .A(n897), .B(n898), .Z(c[124]) );
  IV U1028 ( .A(a[125]), .Z(n903) );
  NOR U1029 ( .A(n898), .B(n897), .Z(n902) );
  IV U1030 ( .A(b[124]), .Z(n900) );
  NOR U1031 ( .A(n900), .B(n899), .Z(n901) );
  NOR U1032 ( .A(n902), .B(n901), .Z(n905) );
  XOR U1033 ( .A(b[125]), .B(n905), .Z(n904) );
  XOR U1034 ( .A(n903), .B(n904), .Z(c[125]) );
  IV U1035 ( .A(a[126]), .Z(n909) );
  NOR U1036 ( .A(n904), .B(n903), .Z(n908) );
  IV U1037 ( .A(b[125]), .Z(n906) );
  NOR U1038 ( .A(n906), .B(n905), .Z(n907) );
  NOR U1039 ( .A(n908), .B(n907), .Z(n911) );
  XOR U1040 ( .A(b[126]), .B(n911), .Z(n910) );
  XOR U1041 ( .A(n909), .B(n910), .Z(c[126]) );
  NOR U1042 ( .A(n910), .B(n909), .Z(n914) );
  IV U1043 ( .A(b[126]), .Z(n912) );
  NOR U1044 ( .A(n912), .B(n911), .Z(n913) );
  NOR U1045 ( .A(n914), .B(n913), .Z(n1111) );
  IV U1046 ( .A(n1111), .Z(n1112) );
  XOR U1047 ( .A(a[127]), .B(n1112), .Z(n915) );
  XOR U1048 ( .A(b[127]), .B(n915), .Z(c[127]) );
  XOR U1049 ( .A(b[12]), .B(n916), .Z(n917) );
  XOR U1050 ( .A(a[12]), .B(n917), .Z(c[12]) );
  XOR U1051 ( .A(b[13]), .B(n918), .Z(n919) );
  XOR U1052 ( .A(a[13]), .B(n919), .Z(c[13]) );
  XOR U1053 ( .A(b[14]), .B(n920), .Z(n921) );
  XOR U1054 ( .A(a[14]), .B(n921), .Z(c[14]) );
  XOR U1055 ( .A(b[15]), .B(n922), .Z(n923) );
  XOR U1056 ( .A(a[15]), .B(n923), .Z(c[15]) );
  XOR U1057 ( .A(b[16]), .B(n924), .Z(n925) );
  XOR U1058 ( .A(a[16]), .B(n925), .Z(c[16]) );
  XOR U1059 ( .A(b[17]), .B(n926), .Z(n927) );
  XOR U1060 ( .A(a[17]), .B(n927), .Z(c[17]) );
  XOR U1061 ( .A(b[18]), .B(n928), .Z(n929) );
  XOR U1062 ( .A(a[18]), .B(n929), .Z(c[18]) );
  XOR U1063 ( .A(b[19]), .B(n930), .Z(n931) );
  XOR U1064 ( .A(a[19]), .B(n931), .Z(c[19]) );
  XOR U1065 ( .A(n933), .B(n932), .Z(c[1]) );
  XOR U1066 ( .A(b[20]), .B(n934), .Z(n935) );
  XOR U1067 ( .A(a[20]), .B(n935), .Z(c[20]) );
  XOR U1068 ( .A(b[21]), .B(n936), .Z(n937) );
  XOR U1069 ( .A(a[21]), .B(n937), .Z(c[21]) );
  XOR U1070 ( .A(b[22]), .B(n938), .Z(n939) );
  XOR U1071 ( .A(a[22]), .B(n939), .Z(c[22]) );
  XOR U1072 ( .A(b[23]), .B(n940), .Z(n941) );
  XOR U1073 ( .A(a[23]), .B(n941), .Z(c[23]) );
  XOR U1074 ( .A(b[24]), .B(n942), .Z(n943) );
  XOR U1075 ( .A(a[24]), .B(n943), .Z(c[24]) );
  XOR U1076 ( .A(b[25]), .B(n944), .Z(n945) );
  XOR U1077 ( .A(a[25]), .B(n945), .Z(c[25]) );
  XOR U1078 ( .A(b[26]), .B(n946), .Z(n947) );
  XOR U1079 ( .A(a[26]), .B(n947), .Z(c[26]) );
  XOR U1080 ( .A(b[27]), .B(n948), .Z(n949) );
  XOR U1081 ( .A(a[27]), .B(n949), .Z(c[27]) );
  XOR U1082 ( .A(b[28]), .B(n950), .Z(n951) );
  XOR U1083 ( .A(a[28]), .B(n951), .Z(c[28]) );
  XOR U1084 ( .A(b[29]), .B(n952), .Z(n953) );
  XOR U1085 ( .A(a[29]), .B(n953), .Z(c[29]) );
  XOR U1086 ( .A(b[2]), .B(n954), .Z(n955) );
  XOR U1087 ( .A(n956), .B(n955), .Z(c[2]) );
  XOR U1088 ( .A(b[30]), .B(n957), .Z(n958) );
  XOR U1089 ( .A(a[30]), .B(n958), .Z(c[30]) );
  XOR U1090 ( .A(b[31]), .B(n959), .Z(n960) );
  XOR U1091 ( .A(a[31]), .B(n960), .Z(c[31]) );
  XOR U1092 ( .A(b[32]), .B(n961), .Z(n962) );
  XOR U1093 ( .A(a[32]), .B(n962), .Z(c[32]) );
  XOR U1094 ( .A(b[33]), .B(n963), .Z(n964) );
  XOR U1095 ( .A(a[33]), .B(n964), .Z(c[33]) );
  XOR U1096 ( .A(b[34]), .B(n965), .Z(n966) );
  XOR U1097 ( .A(a[34]), .B(n966), .Z(c[34]) );
  XOR U1098 ( .A(b[35]), .B(n967), .Z(n968) );
  XOR U1099 ( .A(a[35]), .B(n968), .Z(c[35]) );
  XOR U1100 ( .A(b[36]), .B(n969), .Z(n970) );
  XOR U1101 ( .A(a[36]), .B(n970), .Z(c[36]) );
  XOR U1102 ( .A(b[37]), .B(n971), .Z(n972) );
  XOR U1103 ( .A(a[37]), .B(n972), .Z(c[37]) );
  XOR U1104 ( .A(b[38]), .B(n973), .Z(n974) );
  XOR U1105 ( .A(a[38]), .B(n974), .Z(c[38]) );
  XOR U1106 ( .A(b[39]), .B(n975), .Z(n976) );
  XOR U1107 ( .A(a[39]), .B(n976), .Z(c[39]) );
  XOR U1108 ( .A(b[3]), .B(n977), .Z(n978) );
  XOR U1109 ( .A(a[3]), .B(n978), .Z(c[3]) );
  XOR U1110 ( .A(b[40]), .B(n979), .Z(n980) );
  XOR U1111 ( .A(a[40]), .B(n980), .Z(c[40]) );
  XOR U1112 ( .A(b[41]), .B(n981), .Z(n982) );
  XOR U1113 ( .A(a[41]), .B(n982), .Z(c[41]) );
  XOR U1114 ( .A(b[42]), .B(n983), .Z(n984) );
  XOR U1115 ( .A(a[42]), .B(n984), .Z(c[42]) );
  XOR U1116 ( .A(b[43]), .B(n985), .Z(n986) );
  XOR U1117 ( .A(a[43]), .B(n986), .Z(c[43]) );
  XOR U1118 ( .A(b[44]), .B(n987), .Z(n988) );
  XOR U1119 ( .A(a[44]), .B(n988), .Z(c[44]) );
  XOR U1120 ( .A(b[45]), .B(n989), .Z(n990) );
  XOR U1121 ( .A(a[45]), .B(n990), .Z(c[45]) );
  XOR U1122 ( .A(b[46]), .B(n991), .Z(n992) );
  XOR U1123 ( .A(a[46]), .B(n992), .Z(c[46]) );
  XOR U1124 ( .A(b[47]), .B(n993), .Z(n994) );
  XOR U1125 ( .A(a[47]), .B(n994), .Z(c[47]) );
  XOR U1126 ( .A(b[48]), .B(n995), .Z(n996) );
  XOR U1127 ( .A(a[48]), .B(n996), .Z(c[48]) );
  XOR U1128 ( .A(b[49]), .B(n997), .Z(n998) );
  XOR U1129 ( .A(a[49]), .B(n998), .Z(c[49]) );
  XOR U1130 ( .A(b[4]), .B(n999), .Z(n1000) );
  XOR U1131 ( .A(a[4]), .B(n1000), .Z(c[4]) );
  XOR U1132 ( .A(b[50]), .B(n1001), .Z(n1002) );
  XOR U1133 ( .A(a[50]), .B(n1002), .Z(c[50]) );
  XOR U1134 ( .A(b[51]), .B(n1003), .Z(n1004) );
  XOR U1135 ( .A(a[51]), .B(n1004), .Z(c[51]) );
  XOR U1136 ( .A(b[52]), .B(n1005), .Z(n1006) );
  XOR U1137 ( .A(a[52]), .B(n1006), .Z(c[52]) );
  XOR U1138 ( .A(b[53]), .B(n1007), .Z(n1008) );
  XOR U1139 ( .A(a[53]), .B(n1008), .Z(c[53]) );
  XOR U1140 ( .A(b[54]), .B(n1009), .Z(n1010) );
  XOR U1141 ( .A(a[54]), .B(n1010), .Z(c[54]) );
  XOR U1142 ( .A(b[55]), .B(n1011), .Z(n1012) );
  XOR U1143 ( .A(a[55]), .B(n1012), .Z(c[55]) );
  XOR U1144 ( .A(b[56]), .B(n1013), .Z(n1014) );
  XOR U1145 ( .A(a[56]), .B(n1014), .Z(c[56]) );
  XOR U1146 ( .A(b[57]), .B(n1015), .Z(n1016) );
  XOR U1147 ( .A(a[57]), .B(n1016), .Z(c[57]) );
  XOR U1148 ( .A(b[58]), .B(n1017), .Z(n1018) );
  XOR U1149 ( .A(a[58]), .B(n1018), .Z(c[58]) );
  XOR U1150 ( .A(b[59]), .B(n1019), .Z(n1020) );
  XOR U1151 ( .A(a[59]), .B(n1020), .Z(c[59]) );
  XOR U1152 ( .A(b[5]), .B(n1021), .Z(n1022) );
  XOR U1153 ( .A(a[5]), .B(n1022), .Z(c[5]) );
  XOR U1154 ( .A(b[60]), .B(n1023), .Z(n1024) );
  XOR U1155 ( .A(a[60]), .B(n1024), .Z(c[60]) );
  XOR U1156 ( .A(b[61]), .B(n1025), .Z(n1026) );
  XOR U1157 ( .A(a[61]), .B(n1026), .Z(c[61]) );
  XOR U1158 ( .A(b[62]), .B(n1027), .Z(n1028) );
  XOR U1159 ( .A(a[62]), .B(n1028), .Z(c[62]) );
  XOR U1160 ( .A(b[63]), .B(n1029), .Z(n1030) );
  XOR U1161 ( .A(a[63]), .B(n1030), .Z(c[63]) );
  XOR U1162 ( .A(b[64]), .B(n1031), .Z(n1032) );
  XOR U1163 ( .A(a[64]), .B(n1032), .Z(c[64]) );
  XOR U1164 ( .A(b[65]), .B(n1033), .Z(n1034) );
  XOR U1165 ( .A(a[65]), .B(n1034), .Z(c[65]) );
  XOR U1166 ( .A(b[66]), .B(n1035), .Z(n1036) );
  XOR U1167 ( .A(a[66]), .B(n1036), .Z(c[66]) );
  XOR U1168 ( .A(b[67]), .B(n1037), .Z(n1038) );
  XOR U1169 ( .A(a[67]), .B(n1038), .Z(c[67]) );
  XOR U1170 ( .A(b[68]), .B(n1039), .Z(n1040) );
  XOR U1171 ( .A(a[68]), .B(n1040), .Z(c[68]) );
  XOR U1172 ( .A(b[69]), .B(n1041), .Z(n1042) );
  XOR U1173 ( .A(a[69]), .B(n1042), .Z(c[69]) );
  XOR U1174 ( .A(b[6]), .B(n1043), .Z(n1044) );
  XOR U1175 ( .A(a[6]), .B(n1044), .Z(c[6]) );
  XOR U1176 ( .A(b[70]), .B(n1045), .Z(n1046) );
  XOR U1177 ( .A(a[70]), .B(n1046), .Z(c[70]) );
  XOR U1178 ( .A(b[71]), .B(n1047), .Z(n1048) );
  XOR U1179 ( .A(a[71]), .B(n1048), .Z(c[71]) );
  XOR U1180 ( .A(b[72]), .B(n1049), .Z(n1050) );
  XOR U1181 ( .A(a[72]), .B(n1050), .Z(c[72]) );
  XOR U1182 ( .A(b[73]), .B(n1051), .Z(n1052) );
  XOR U1183 ( .A(a[73]), .B(n1052), .Z(c[73]) );
  XOR U1184 ( .A(b[74]), .B(n1053), .Z(n1054) );
  XOR U1185 ( .A(a[74]), .B(n1054), .Z(c[74]) );
  XOR U1186 ( .A(b[75]), .B(n1055), .Z(n1056) );
  XOR U1187 ( .A(a[75]), .B(n1056), .Z(c[75]) );
  XOR U1188 ( .A(b[76]), .B(n1057), .Z(n1058) );
  XOR U1189 ( .A(a[76]), .B(n1058), .Z(c[76]) );
  XOR U1190 ( .A(b[77]), .B(n1059), .Z(n1060) );
  XOR U1191 ( .A(a[77]), .B(n1060), .Z(c[77]) );
  XOR U1192 ( .A(b[78]), .B(n1061), .Z(n1062) );
  XOR U1193 ( .A(a[78]), .B(n1062), .Z(c[78]) );
  XOR U1194 ( .A(b[79]), .B(n1063), .Z(n1064) );
  XOR U1195 ( .A(a[79]), .B(n1064), .Z(c[79]) );
  XOR U1196 ( .A(b[7]), .B(n1065), .Z(n1066) );
  XOR U1197 ( .A(a[7]), .B(n1066), .Z(c[7]) );
  XOR U1198 ( .A(b[80]), .B(n1067), .Z(n1068) );
  XOR U1199 ( .A(a[80]), .B(n1068), .Z(c[80]) );
  XOR U1200 ( .A(b[81]), .B(n1069), .Z(n1070) );
  XOR U1201 ( .A(a[81]), .B(n1070), .Z(c[81]) );
  XOR U1202 ( .A(b[82]), .B(n1071), .Z(n1072) );
  XOR U1203 ( .A(a[82]), .B(n1072), .Z(c[82]) );
  XOR U1204 ( .A(b[83]), .B(n1073), .Z(n1074) );
  XOR U1205 ( .A(a[83]), .B(n1074), .Z(c[83]) );
  XOR U1206 ( .A(b[84]), .B(n1075), .Z(n1076) );
  XOR U1207 ( .A(a[84]), .B(n1076), .Z(c[84]) );
  XOR U1208 ( .A(b[85]), .B(n1077), .Z(n1078) );
  XOR U1209 ( .A(a[85]), .B(n1078), .Z(c[85]) );
  XOR U1210 ( .A(b[86]), .B(n1079), .Z(n1080) );
  XOR U1211 ( .A(a[86]), .B(n1080), .Z(c[86]) );
  XOR U1212 ( .A(b[87]), .B(n1081), .Z(n1082) );
  XOR U1213 ( .A(a[87]), .B(n1082), .Z(c[87]) );
  XOR U1214 ( .A(b[88]), .B(n1083), .Z(n1084) );
  XOR U1215 ( .A(a[88]), .B(n1084), .Z(c[88]) );
  XOR U1216 ( .A(b[89]), .B(n1085), .Z(n1086) );
  XOR U1217 ( .A(a[89]), .B(n1086), .Z(c[89]) );
  XOR U1218 ( .A(b[8]), .B(n1087), .Z(n1088) );
  XOR U1219 ( .A(a[8]), .B(n1088), .Z(c[8]) );
  XOR U1220 ( .A(b[90]), .B(n1089), .Z(n1090) );
  XOR U1221 ( .A(a[90]), .B(n1090), .Z(c[90]) );
  XOR U1222 ( .A(b[91]), .B(n1091), .Z(n1092) );
  XOR U1223 ( .A(a[91]), .B(n1092), .Z(c[91]) );
  XOR U1224 ( .A(b[92]), .B(n1093), .Z(n1094) );
  XOR U1225 ( .A(a[92]), .B(n1094), .Z(c[92]) );
  XOR U1226 ( .A(b[93]), .B(n1095), .Z(n1096) );
  XOR U1227 ( .A(a[93]), .B(n1096), .Z(c[93]) );
  XOR U1228 ( .A(b[94]), .B(n1097), .Z(n1098) );
  XOR U1229 ( .A(a[94]), .B(n1098), .Z(c[94]) );
  XOR U1230 ( .A(b[95]), .B(n1099), .Z(n1100) );
  XOR U1231 ( .A(a[95]), .B(n1100), .Z(c[95]) );
  XOR U1232 ( .A(b[96]), .B(n1101), .Z(n1102) );
  XOR U1233 ( .A(a[96]), .B(n1102), .Z(c[96]) );
  XOR U1234 ( .A(b[97]), .B(n1103), .Z(n1104) );
  XOR U1235 ( .A(a[97]), .B(n1104), .Z(c[97]) );
  XOR U1236 ( .A(b[98]), .B(n1105), .Z(n1106) );
  XOR U1237 ( .A(a[98]), .B(n1106), .Z(c[98]) );
  XOR U1238 ( .A(a[99]), .B(n1107), .Z(n1108) );
  XOR U1239 ( .A(b[99]), .B(n1108), .Z(c[99]) );
  XOR U1240 ( .A(a[9]), .B(n1109), .Z(n1110) );
  XOR U1241 ( .A(b[9]), .B(n1110), .Z(c[9]) );
endmodule

