
module sum ( a, b, c );
  input [1023:0] a;
  input [1023:0] b;
  output [1024:0] c;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143;

  IV U2 ( .A(a[0]), .Z(n1003) );
  IV U3 ( .A(b[0]), .Z(n1002) );
  XOR U4 ( .A(n1003), .B(n1002), .Z(c[0]) );
  IV U5 ( .A(b[999]), .Z(n3998) );
  IV U6 ( .A(a[999]), .Z(n2) );
  NOR U7 ( .A(n3998), .B(n2), .Z(n4000) );
  IV U8 ( .A(a[998]), .Z(n3995) );
  IV U9 ( .A(b[998]), .Z(n3) );
  NOR U10 ( .A(n3995), .B(n3), .Z(n3997) );
  IV U11 ( .A(a[997]), .Z(n3992) );
  IV U12 ( .A(b[997]), .Z(n4) );
  NOR U13 ( .A(n3992), .B(n4), .Z(n3994) );
  IV U14 ( .A(a[996]), .Z(n3989) );
  IV U15 ( .A(b[996]), .Z(n5) );
  NOR U16 ( .A(n3989), .B(n5), .Z(n3991) );
  IV U17 ( .A(a[995]), .Z(n3986) );
  IV U18 ( .A(b[995]), .Z(n6) );
  NOR U19 ( .A(n3986), .B(n6), .Z(n3988) );
  IV U20 ( .A(a[994]), .Z(n3983) );
  IV U21 ( .A(b[994]), .Z(n7) );
  NOR U22 ( .A(n3983), .B(n7), .Z(n3985) );
  IV U23 ( .A(a[993]), .Z(n3980) );
  IV U24 ( .A(b[993]), .Z(n8) );
  NOR U25 ( .A(n3980), .B(n8), .Z(n3982) );
  IV U26 ( .A(a[992]), .Z(n3977) );
  IV U27 ( .A(b[992]), .Z(n9) );
  NOR U28 ( .A(n3977), .B(n9), .Z(n3979) );
  IV U29 ( .A(a[991]), .Z(n3974) );
  IV U30 ( .A(b[991]), .Z(n10) );
  NOR U31 ( .A(n3974), .B(n10), .Z(n3976) );
  IV U32 ( .A(a[990]), .Z(n3971) );
  IV U33 ( .A(b[990]), .Z(n11) );
  NOR U34 ( .A(n3971), .B(n11), .Z(n3973) );
  IV U35 ( .A(a[989]), .Z(n3968) );
  IV U36 ( .A(b[989]), .Z(n12) );
  NOR U37 ( .A(n3968), .B(n12), .Z(n3970) );
  IV U38 ( .A(a[988]), .Z(n3965) );
  IV U39 ( .A(b[988]), .Z(n13) );
  NOR U40 ( .A(n3965), .B(n13), .Z(n3967) );
  IV U41 ( .A(a[987]), .Z(n3962) );
  IV U42 ( .A(b[987]), .Z(n14) );
  NOR U43 ( .A(n3962), .B(n14), .Z(n3964) );
  IV U44 ( .A(a[986]), .Z(n3959) );
  IV U45 ( .A(b[986]), .Z(n15) );
  NOR U46 ( .A(n3959), .B(n15), .Z(n3961) );
  IV U47 ( .A(a[985]), .Z(n3956) );
  IV U48 ( .A(b[985]), .Z(n16) );
  NOR U49 ( .A(n3956), .B(n16), .Z(n3958) );
  IV U50 ( .A(a[984]), .Z(n3953) );
  IV U51 ( .A(b[984]), .Z(n17) );
  NOR U52 ( .A(n3953), .B(n17), .Z(n3955) );
  IV U53 ( .A(a[983]), .Z(n3950) );
  IV U54 ( .A(b[983]), .Z(n18) );
  NOR U55 ( .A(n3950), .B(n18), .Z(n3952) );
  IV U56 ( .A(a[982]), .Z(n3947) );
  IV U57 ( .A(b[982]), .Z(n19) );
  NOR U58 ( .A(n3947), .B(n19), .Z(n3949) );
  IV U59 ( .A(a[981]), .Z(n3944) );
  IV U60 ( .A(b[981]), .Z(n20) );
  NOR U61 ( .A(n3944), .B(n20), .Z(n3946) );
  IV U62 ( .A(a[980]), .Z(n3941) );
  IV U63 ( .A(b[980]), .Z(n21) );
  NOR U64 ( .A(n3941), .B(n21), .Z(n3943) );
  IV U65 ( .A(a[979]), .Z(n3938) );
  IV U66 ( .A(b[979]), .Z(n22) );
  NOR U67 ( .A(n3938), .B(n22), .Z(n3940) );
  IV U68 ( .A(a[978]), .Z(n3935) );
  IV U69 ( .A(b[978]), .Z(n23) );
  NOR U70 ( .A(n3935), .B(n23), .Z(n3937) );
  IV U71 ( .A(a[977]), .Z(n3932) );
  IV U72 ( .A(b[977]), .Z(n24) );
  NOR U73 ( .A(n3932), .B(n24), .Z(n3934) );
  IV U74 ( .A(a[976]), .Z(n3929) );
  IV U75 ( .A(b[976]), .Z(n25) );
  NOR U76 ( .A(n3929), .B(n25), .Z(n3931) );
  IV U77 ( .A(a[975]), .Z(n3926) );
  IV U78 ( .A(b[975]), .Z(n26) );
  NOR U79 ( .A(n3926), .B(n26), .Z(n3928) );
  IV U80 ( .A(a[974]), .Z(n3923) );
  IV U81 ( .A(b[974]), .Z(n27) );
  NOR U82 ( .A(n3923), .B(n27), .Z(n3925) );
  IV U83 ( .A(a[973]), .Z(n3920) );
  IV U84 ( .A(b[973]), .Z(n28) );
  NOR U85 ( .A(n3920), .B(n28), .Z(n3922) );
  IV U86 ( .A(a[972]), .Z(n3917) );
  IV U87 ( .A(b[972]), .Z(n29) );
  NOR U88 ( .A(n3917), .B(n29), .Z(n3919) );
  IV U89 ( .A(a[971]), .Z(n3914) );
  IV U90 ( .A(b[971]), .Z(n30) );
  NOR U91 ( .A(n3914), .B(n30), .Z(n3916) );
  IV U92 ( .A(a[970]), .Z(n3911) );
  IV U93 ( .A(b[970]), .Z(n31) );
  NOR U94 ( .A(n3911), .B(n31), .Z(n3913) );
  IV U95 ( .A(a[969]), .Z(n3908) );
  IV U96 ( .A(b[969]), .Z(n32) );
  NOR U97 ( .A(n3908), .B(n32), .Z(n3910) );
  IV U98 ( .A(a[968]), .Z(n3905) );
  IV U99 ( .A(b[968]), .Z(n33) );
  NOR U100 ( .A(n3905), .B(n33), .Z(n3907) );
  IV U101 ( .A(a[967]), .Z(n3902) );
  IV U102 ( .A(b[967]), .Z(n34) );
  NOR U103 ( .A(n3902), .B(n34), .Z(n3904) );
  IV U104 ( .A(a[966]), .Z(n3899) );
  IV U105 ( .A(b[966]), .Z(n35) );
  NOR U106 ( .A(n3899), .B(n35), .Z(n3901) );
  IV U107 ( .A(a[965]), .Z(n3896) );
  IV U108 ( .A(b[965]), .Z(n36) );
  NOR U109 ( .A(n3896), .B(n36), .Z(n3898) );
  IV U110 ( .A(a[964]), .Z(n3893) );
  IV U111 ( .A(b[964]), .Z(n37) );
  NOR U112 ( .A(n3893), .B(n37), .Z(n3895) );
  IV U113 ( .A(a[963]), .Z(n3890) );
  IV U114 ( .A(b[963]), .Z(n38) );
  NOR U115 ( .A(n3890), .B(n38), .Z(n3892) );
  IV U116 ( .A(a[962]), .Z(n3887) );
  IV U117 ( .A(b[962]), .Z(n39) );
  NOR U118 ( .A(n3887), .B(n39), .Z(n3889) );
  IV U119 ( .A(a[961]), .Z(n3884) );
  IV U120 ( .A(b[961]), .Z(n40) );
  NOR U121 ( .A(n3884), .B(n40), .Z(n3886) );
  IV U122 ( .A(a[960]), .Z(n3881) );
  IV U123 ( .A(b[960]), .Z(n41) );
  NOR U124 ( .A(n3881), .B(n41), .Z(n3883) );
  IV U125 ( .A(a[959]), .Z(n3878) );
  IV U126 ( .A(b[959]), .Z(n42) );
  NOR U127 ( .A(n3878), .B(n42), .Z(n3880) );
  IV U128 ( .A(a[958]), .Z(n3875) );
  IV U129 ( .A(b[958]), .Z(n43) );
  NOR U130 ( .A(n3875), .B(n43), .Z(n3877) );
  IV U131 ( .A(a[957]), .Z(n3872) );
  IV U132 ( .A(b[957]), .Z(n44) );
  NOR U133 ( .A(n3872), .B(n44), .Z(n3874) );
  IV U134 ( .A(a[956]), .Z(n3869) );
  IV U135 ( .A(b[956]), .Z(n45) );
  NOR U136 ( .A(n3869), .B(n45), .Z(n3871) );
  IV U137 ( .A(a[955]), .Z(n3866) );
  IV U138 ( .A(b[955]), .Z(n46) );
  NOR U139 ( .A(n3866), .B(n46), .Z(n3868) );
  IV U140 ( .A(a[954]), .Z(n3863) );
  IV U141 ( .A(b[954]), .Z(n47) );
  NOR U142 ( .A(n3863), .B(n47), .Z(n3865) );
  IV U143 ( .A(a[953]), .Z(n3860) );
  IV U144 ( .A(b[953]), .Z(n48) );
  NOR U145 ( .A(n3860), .B(n48), .Z(n3862) );
  IV U146 ( .A(a[952]), .Z(n3857) );
  IV U147 ( .A(b[952]), .Z(n49) );
  NOR U148 ( .A(n3857), .B(n49), .Z(n3859) );
  IV U149 ( .A(a[951]), .Z(n3854) );
  IV U150 ( .A(b[951]), .Z(n50) );
  NOR U151 ( .A(n3854), .B(n50), .Z(n3856) );
  IV U152 ( .A(a[950]), .Z(n3851) );
  IV U153 ( .A(b[950]), .Z(n51) );
  NOR U154 ( .A(n3851), .B(n51), .Z(n3853) );
  IV U155 ( .A(a[949]), .Z(n3848) );
  IV U156 ( .A(b[949]), .Z(n52) );
  NOR U157 ( .A(n3848), .B(n52), .Z(n3850) );
  IV U158 ( .A(a[948]), .Z(n3845) );
  IV U159 ( .A(b[948]), .Z(n53) );
  NOR U160 ( .A(n3845), .B(n53), .Z(n3847) );
  IV U161 ( .A(a[947]), .Z(n3842) );
  IV U162 ( .A(b[947]), .Z(n54) );
  NOR U163 ( .A(n3842), .B(n54), .Z(n3844) );
  IV U164 ( .A(a[946]), .Z(n3839) );
  IV U165 ( .A(b[946]), .Z(n55) );
  NOR U166 ( .A(n3839), .B(n55), .Z(n3841) );
  IV U167 ( .A(a[945]), .Z(n3836) );
  IV U168 ( .A(b[945]), .Z(n56) );
  NOR U169 ( .A(n3836), .B(n56), .Z(n3838) );
  IV U170 ( .A(a[944]), .Z(n3833) );
  IV U171 ( .A(b[944]), .Z(n57) );
  NOR U172 ( .A(n3833), .B(n57), .Z(n3835) );
  IV U173 ( .A(a[943]), .Z(n3830) );
  IV U174 ( .A(b[943]), .Z(n58) );
  NOR U175 ( .A(n3830), .B(n58), .Z(n3832) );
  IV U176 ( .A(a[942]), .Z(n3827) );
  IV U177 ( .A(b[942]), .Z(n59) );
  NOR U178 ( .A(n3827), .B(n59), .Z(n3829) );
  IV U179 ( .A(a[941]), .Z(n3824) );
  IV U180 ( .A(b[941]), .Z(n60) );
  NOR U181 ( .A(n3824), .B(n60), .Z(n3826) );
  IV U182 ( .A(a[940]), .Z(n3821) );
  IV U183 ( .A(b[940]), .Z(n61) );
  NOR U184 ( .A(n3821), .B(n61), .Z(n3823) );
  IV U185 ( .A(a[939]), .Z(n3818) );
  IV U186 ( .A(b[939]), .Z(n62) );
  NOR U187 ( .A(n3818), .B(n62), .Z(n3820) );
  IV U188 ( .A(a[938]), .Z(n3815) );
  IV U189 ( .A(b[938]), .Z(n63) );
  NOR U190 ( .A(n3815), .B(n63), .Z(n3817) );
  IV U191 ( .A(a[937]), .Z(n3812) );
  IV U192 ( .A(b[937]), .Z(n64) );
  NOR U193 ( .A(n3812), .B(n64), .Z(n3814) );
  IV U194 ( .A(a[936]), .Z(n3809) );
  IV U195 ( .A(b[936]), .Z(n65) );
  NOR U196 ( .A(n3809), .B(n65), .Z(n3811) );
  IV U197 ( .A(a[935]), .Z(n3806) );
  IV U198 ( .A(b[935]), .Z(n66) );
  NOR U199 ( .A(n3806), .B(n66), .Z(n3808) );
  IV U200 ( .A(a[934]), .Z(n3803) );
  IV U201 ( .A(b[934]), .Z(n67) );
  NOR U202 ( .A(n3803), .B(n67), .Z(n3805) );
  IV U203 ( .A(a[933]), .Z(n3800) );
  IV U204 ( .A(b[933]), .Z(n68) );
  NOR U205 ( .A(n3800), .B(n68), .Z(n3802) );
  IV U206 ( .A(a[932]), .Z(n3797) );
  IV U207 ( .A(b[932]), .Z(n69) );
  NOR U208 ( .A(n3797), .B(n69), .Z(n3799) );
  IV U209 ( .A(a[931]), .Z(n3794) );
  IV U210 ( .A(b[931]), .Z(n70) );
  NOR U211 ( .A(n3794), .B(n70), .Z(n3796) );
  IV U212 ( .A(a[930]), .Z(n3791) );
  IV U213 ( .A(b[930]), .Z(n71) );
  NOR U214 ( .A(n3791), .B(n71), .Z(n3793) );
  IV U215 ( .A(a[929]), .Z(n3788) );
  IV U216 ( .A(b[929]), .Z(n72) );
  NOR U217 ( .A(n3788), .B(n72), .Z(n3790) );
  IV U218 ( .A(a[928]), .Z(n3785) );
  IV U219 ( .A(b[928]), .Z(n73) );
  NOR U220 ( .A(n3785), .B(n73), .Z(n3787) );
  IV U221 ( .A(a[927]), .Z(n3782) );
  IV U222 ( .A(b[927]), .Z(n74) );
  NOR U223 ( .A(n3782), .B(n74), .Z(n3784) );
  IV U224 ( .A(a[926]), .Z(n3779) );
  IV U225 ( .A(b[926]), .Z(n75) );
  NOR U226 ( .A(n3779), .B(n75), .Z(n3781) );
  IV U227 ( .A(a[925]), .Z(n3776) );
  IV U228 ( .A(b[925]), .Z(n76) );
  NOR U229 ( .A(n3776), .B(n76), .Z(n3778) );
  IV U230 ( .A(a[924]), .Z(n3773) );
  IV U231 ( .A(b[924]), .Z(n77) );
  NOR U232 ( .A(n3773), .B(n77), .Z(n3775) );
  IV U233 ( .A(a[923]), .Z(n3770) );
  IV U234 ( .A(b[923]), .Z(n78) );
  NOR U235 ( .A(n3770), .B(n78), .Z(n3772) );
  IV U236 ( .A(a[922]), .Z(n3767) );
  IV U237 ( .A(b[922]), .Z(n79) );
  NOR U238 ( .A(n3767), .B(n79), .Z(n3769) );
  IV U239 ( .A(a[921]), .Z(n3764) );
  IV U240 ( .A(b[921]), .Z(n80) );
  NOR U241 ( .A(n3764), .B(n80), .Z(n3766) );
  IV U242 ( .A(a[920]), .Z(n3761) );
  IV U243 ( .A(b[920]), .Z(n81) );
  NOR U244 ( .A(n3761), .B(n81), .Z(n3763) );
  IV U245 ( .A(a[919]), .Z(n3758) );
  IV U246 ( .A(b[919]), .Z(n82) );
  NOR U247 ( .A(n3758), .B(n82), .Z(n3760) );
  IV U248 ( .A(a[918]), .Z(n3755) );
  IV U249 ( .A(b[918]), .Z(n83) );
  NOR U250 ( .A(n3755), .B(n83), .Z(n3757) );
  IV U251 ( .A(a[917]), .Z(n3752) );
  IV U252 ( .A(b[917]), .Z(n84) );
  NOR U253 ( .A(n3752), .B(n84), .Z(n3754) );
  IV U254 ( .A(a[916]), .Z(n3749) );
  IV U255 ( .A(b[916]), .Z(n85) );
  NOR U256 ( .A(n3749), .B(n85), .Z(n3751) );
  IV U257 ( .A(a[915]), .Z(n3746) );
  IV U258 ( .A(b[915]), .Z(n86) );
  NOR U259 ( .A(n3746), .B(n86), .Z(n3748) );
  IV U260 ( .A(a[914]), .Z(n3743) );
  IV U261 ( .A(b[914]), .Z(n87) );
  NOR U262 ( .A(n3743), .B(n87), .Z(n3745) );
  IV U263 ( .A(a[913]), .Z(n3740) );
  IV U264 ( .A(b[913]), .Z(n88) );
  NOR U265 ( .A(n3740), .B(n88), .Z(n3742) );
  IV U266 ( .A(a[912]), .Z(n3737) );
  IV U267 ( .A(b[912]), .Z(n89) );
  NOR U268 ( .A(n3737), .B(n89), .Z(n3739) );
  IV U269 ( .A(a[911]), .Z(n3734) );
  IV U270 ( .A(b[911]), .Z(n90) );
  NOR U271 ( .A(n3734), .B(n90), .Z(n3736) );
  IV U272 ( .A(a[910]), .Z(n3731) );
  IV U273 ( .A(b[910]), .Z(n91) );
  NOR U274 ( .A(n3731), .B(n91), .Z(n3733) );
  IV U275 ( .A(a[909]), .Z(n3728) );
  IV U276 ( .A(b[909]), .Z(n92) );
  NOR U277 ( .A(n3728), .B(n92), .Z(n3730) );
  IV U278 ( .A(a[908]), .Z(n3725) );
  IV U279 ( .A(b[908]), .Z(n93) );
  NOR U280 ( .A(n3725), .B(n93), .Z(n3727) );
  IV U281 ( .A(a[907]), .Z(n3722) );
  IV U282 ( .A(b[907]), .Z(n94) );
  NOR U283 ( .A(n3722), .B(n94), .Z(n3724) );
  IV U284 ( .A(a[906]), .Z(n3719) );
  IV U285 ( .A(b[906]), .Z(n95) );
  NOR U286 ( .A(n3719), .B(n95), .Z(n3721) );
  IV U287 ( .A(a[905]), .Z(n3716) );
  IV U288 ( .A(b[905]), .Z(n96) );
  NOR U289 ( .A(n3716), .B(n96), .Z(n3718) );
  IV U290 ( .A(a[904]), .Z(n3713) );
  IV U291 ( .A(b[904]), .Z(n97) );
  NOR U292 ( .A(n3713), .B(n97), .Z(n3715) );
  IV U293 ( .A(a[903]), .Z(n3710) );
  IV U294 ( .A(b[903]), .Z(n98) );
  NOR U295 ( .A(n3710), .B(n98), .Z(n3712) );
  IV U296 ( .A(a[902]), .Z(n3707) );
  IV U297 ( .A(b[902]), .Z(n99) );
  NOR U298 ( .A(n3707), .B(n99), .Z(n3709) );
  IV U299 ( .A(a[901]), .Z(n3704) );
  IV U300 ( .A(b[901]), .Z(n100) );
  NOR U301 ( .A(n3704), .B(n100), .Z(n3706) );
  IV U302 ( .A(a[900]), .Z(n3701) );
  IV U303 ( .A(b[900]), .Z(n101) );
  NOR U304 ( .A(n3701), .B(n101), .Z(n3703) );
  IV U305 ( .A(a[899]), .Z(n3698) );
  IV U306 ( .A(b[899]), .Z(n102) );
  NOR U307 ( .A(n3698), .B(n102), .Z(n3700) );
  IV U308 ( .A(a[898]), .Z(n3695) );
  IV U309 ( .A(b[898]), .Z(n103) );
  NOR U310 ( .A(n3695), .B(n103), .Z(n3697) );
  IV U311 ( .A(a[897]), .Z(n3692) );
  IV U312 ( .A(b[897]), .Z(n104) );
  NOR U313 ( .A(n3692), .B(n104), .Z(n3694) );
  IV U314 ( .A(a[896]), .Z(n3689) );
  IV U315 ( .A(b[896]), .Z(n105) );
  NOR U316 ( .A(n3689), .B(n105), .Z(n3691) );
  IV U317 ( .A(a[895]), .Z(n3686) );
  IV U318 ( .A(b[895]), .Z(n106) );
  NOR U319 ( .A(n3686), .B(n106), .Z(n3688) );
  IV U320 ( .A(a[894]), .Z(n3683) );
  IV U321 ( .A(b[894]), .Z(n107) );
  NOR U322 ( .A(n3683), .B(n107), .Z(n3685) );
  IV U323 ( .A(a[893]), .Z(n3680) );
  IV U324 ( .A(b[893]), .Z(n108) );
  NOR U325 ( .A(n3680), .B(n108), .Z(n3682) );
  IV U326 ( .A(a[892]), .Z(n3677) );
  IV U327 ( .A(b[892]), .Z(n109) );
  NOR U328 ( .A(n3677), .B(n109), .Z(n3679) );
  IV U329 ( .A(a[891]), .Z(n3674) );
  IV U330 ( .A(b[891]), .Z(n110) );
  NOR U331 ( .A(n3674), .B(n110), .Z(n3676) );
  IV U332 ( .A(a[890]), .Z(n3671) );
  IV U333 ( .A(b[890]), .Z(n111) );
  NOR U334 ( .A(n3671), .B(n111), .Z(n3673) );
  IV U335 ( .A(a[889]), .Z(n3668) );
  IV U336 ( .A(b[889]), .Z(n112) );
  NOR U337 ( .A(n3668), .B(n112), .Z(n3670) );
  IV U338 ( .A(a[888]), .Z(n3665) );
  IV U339 ( .A(b[888]), .Z(n113) );
  NOR U340 ( .A(n3665), .B(n113), .Z(n3667) );
  IV U341 ( .A(a[887]), .Z(n3662) );
  IV U342 ( .A(b[887]), .Z(n114) );
  NOR U343 ( .A(n3662), .B(n114), .Z(n3664) );
  IV U344 ( .A(a[886]), .Z(n3659) );
  IV U345 ( .A(b[886]), .Z(n115) );
  NOR U346 ( .A(n3659), .B(n115), .Z(n3661) );
  IV U347 ( .A(a[885]), .Z(n3656) );
  IV U348 ( .A(b[885]), .Z(n116) );
  NOR U349 ( .A(n3656), .B(n116), .Z(n3658) );
  IV U350 ( .A(a[884]), .Z(n3653) );
  IV U351 ( .A(b[884]), .Z(n117) );
  NOR U352 ( .A(n3653), .B(n117), .Z(n3655) );
  IV U353 ( .A(a[883]), .Z(n3650) );
  IV U354 ( .A(b[883]), .Z(n118) );
  NOR U355 ( .A(n3650), .B(n118), .Z(n3652) );
  IV U356 ( .A(a[882]), .Z(n3647) );
  IV U357 ( .A(b[882]), .Z(n119) );
  NOR U358 ( .A(n3647), .B(n119), .Z(n3649) );
  IV U359 ( .A(a[881]), .Z(n3644) );
  IV U360 ( .A(b[881]), .Z(n120) );
  NOR U361 ( .A(n3644), .B(n120), .Z(n3646) );
  IV U362 ( .A(a[880]), .Z(n3641) );
  IV U363 ( .A(b[880]), .Z(n121) );
  NOR U364 ( .A(n3641), .B(n121), .Z(n3643) );
  IV U365 ( .A(a[879]), .Z(n3638) );
  IV U366 ( .A(b[879]), .Z(n122) );
  NOR U367 ( .A(n3638), .B(n122), .Z(n3640) );
  IV U368 ( .A(a[878]), .Z(n3635) );
  IV U369 ( .A(b[878]), .Z(n123) );
  NOR U370 ( .A(n3635), .B(n123), .Z(n3637) );
  IV U371 ( .A(a[877]), .Z(n3632) );
  IV U372 ( .A(b[877]), .Z(n124) );
  NOR U373 ( .A(n3632), .B(n124), .Z(n3634) );
  IV U374 ( .A(a[876]), .Z(n3629) );
  IV U375 ( .A(b[876]), .Z(n125) );
  NOR U376 ( .A(n3629), .B(n125), .Z(n3631) );
  IV U377 ( .A(a[875]), .Z(n3626) );
  IV U378 ( .A(b[875]), .Z(n126) );
  NOR U379 ( .A(n3626), .B(n126), .Z(n3628) );
  IV U380 ( .A(a[874]), .Z(n3623) );
  IV U381 ( .A(b[874]), .Z(n127) );
  NOR U382 ( .A(n3623), .B(n127), .Z(n3625) );
  IV U383 ( .A(a[873]), .Z(n3620) );
  IV U384 ( .A(b[873]), .Z(n128) );
  NOR U385 ( .A(n3620), .B(n128), .Z(n3622) );
  IV U386 ( .A(a[872]), .Z(n3617) );
  IV U387 ( .A(b[872]), .Z(n129) );
  NOR U388 ( .A(n3617), .B(n129), .Z(n3619) );
  IV U389 ( .A(a[871]), .Z(n3614) );
  IV U390 ( .A(b[871]), .Z(n130) );
  NOR U391 ( .A(n3614), .B(n130), .Z(n3616) );
  IV U392 ( .A(a[870]), .Z(n3611) );
  IV U393 ( .A(b[870]), .Z(n131) );
  NOR U394 ( .A(n3611), .B(n131), .Z(n3613) );
  IV U395 ( .A(a[869]), .Z(n3608) );
  IV U396 ( .A(b[869]), .Z(n132) );
  NOR U397 ( .A(n3608), .B(n132), .Z(n3610) );
  IV U398 ( .A(a[868]), .Z(n3605) );
  IV U399 ( .A(b[868]), .Z(n133) );
  NOR U400 ( .A(n3605), .B(n133), .Z(n3607) );
  IV U401 ( .A(a[867]), .Z(n3602) );
  IV U402 ( .A(b[867]), .Z(n134) );
  NOR U403 ( .A(n3602), .B(n134), .Z(n3604) );
  IV U404 ( .A(a[866]), .Z(n3599) );
  IV U405 ( .A(b[866]), .Z(n135) );
  NOR U406 ( .A(n3599), .B(n135), .Z(n3601) );
  IV U407 ( .A(a[865]), .Z(n3596) );
  IV U408 ( .A(b[865]), .Z(n136) );
  NOR U409 ( .A(n3596), .B(n136), .Z(n3598) );
  IV U410 ( .A(a[864]), .Z(n3593) );
  IV U411 ( .A(b[864]), .Z(n137) );
  NOR U412 ( .A(n3593), .B(n137), .Z(n3595) );
  IV U413 ( .A(a[863]), .Z(n3590) );
  IV U414 ( .A(b[863]), .Z(n138) );
  NOR U415 ( .A(n3590), .B(n138), .Z(n3592) );
  IV U416 ( .A(a[862]), .Z(n3587) );
  IV U417 ( .A(b[862]), .Z(n139) );
  NOR U418 ( .A(n3587), .B(n139), .Z(n3589) );
  IV U419 ( .A(a[861]), .Z(n3584) );
  IV U420 ( .A(b[861]), .Z(n140) );
  NOR U421 ( .A(n3584), .B(n140), .Z(n3586) );
  IV U422 ( .A(a[860]), .Z(n3581) );
  IV U423 ( .A(b[860]), .Z(n141) );
  NOR U424 ( .A(n3581), .B(n141), .Z(n3583) );
  IV U425 ( .A(a[859]), .Z(n3578) );
  IV U426 ( .A(b[859]), .Z(n142) );
  NOR U427 ( .A(n3578), .B(n142), .Z(n3580) );
  IV U428 ( .A(a[858]), .Z(n3575) );
  IV U429 ( .A(b[858]), .Z(n143) );
  NOR U430 ( .A(n3575), .B(n143), .Z(n3577) );
  IV U431 ( .A(a[857]), .Z(n3572) );
  IV U432 ( .A(b[857]), .Z(n144) );
  NOR U433 ( .A(n3572), .B(n144), .Z(n3574) );
  IV U434 ( .A(a[856]), .Z(n3569) );
  IV U435 ( .A(b[856]), .Z(n145) );
  NOR U436 ( .A(n3569), .B(n145), .Z(n3571) );
  IV U437 ( .A(a[855]), .Z(n3566) );
  IV U438 ( .A(b[855]), .Z(n146) );
  NOR U439 ( .A(n3566), .B(n146), .Z(n3568) );
  IV U440 ( .A(a[854]), .Z(n3563) );
  IV U441 ( .A(b[854]), .Z(n147) );
  NOR U442 ( .A(n3563), .B(n147), .Z(n3565) );
  IV U443 ( .A(a[853]), .Z(n3560) );
  IV U444 ( .A(b[853]), .Z(n148) );
  NOR U445 ( .A(n3560), .B(n148), .Z(n3562) );
  IV U446 ( .A(a[852]), .Z(n3557) );
  IV U447 ( .A(b[852]), .Z(n149) );
  NOR U448 ( .A(n3557), .B(n149), .Z(n3559) );
  IV U449 ( .A(a[851]), .Z(n3554) );
  IV U450 ( .A(b[851]), .Z(n150) );
  NOR U451 ( .A(n3554), .B(n150), .Z(n3556) );
  IV U452 ( .A(a[850]), .Z(n3551) );
  IV U453 ( .A(b[850]), .Z(n151) );
  NOR U454 ( .A(n3551), .B(n151), .Z(n3553) );
  IV U455 ( .A(a[849]), .Z(n3548) );
  IV U456 ( .A(b[849]), .Z(n152) );
  NOR U457 ( .A(n3548), .B(n152), .Z(n3550) );
  IV U458 ( .A(a[848]), .Z(n3545) );
  IV U459 ( .A(b[848]), .Z(n153) );
  NOR U460 ( .A(n3545), .B(n153), .Z(n3547) );
  IV U461 ( .A(a[847]), .Z(n3542) );
  IV U462 ( .A(b[847]), .Z(n154) );
  NOR U463 ( .A(n3542), .B(n154), .Z(n3544) );
  IV U464 ( .A(a[846]), .Z(n3539) );
  IV U465 ( .A(b[846]), .Z(n155) );
  NOR U466 ( .A(n3539), .B(n155), .Z(n3541) );
  IV U467 ( .A(a[845]), .Z(n3536) );
  IV U468 ( .A(b[845]), .Z(n156) );
  NOR U469 ( .A(n3536), .B(n156), .Z(n3538) );
  IV U470 ( .A(a[844]), .Z(n3533) );
  IV U471 ( .A(b[844]), .Z(n157) );
  NOR U472 ( .A(n3533), .B(n157), .Z(n3535) );
  IV U473 ( .A(a[843]), .Z(n3530) );
  IV U474 ( .A(b[843]), .Z(n158) );
  NOR U475 ( .A(n3530), .B(n158), .Z(n3532) );
  IV U476 ( .A(a[842]), .Z(n3527) );
  IV U477 ( .A(b[842]), .Z(n159) );
  NOR U478 ( .A(n3527), .B(n159), .Z(n3529) );
  IV U479 ( .A(a[841]), .Z(n3524) );
  IV U480 ( .A(b[841]), .Z(n160) );
  NOR U481 ( .A(n3524), .B(n160), .Z(n3526) );
  IV U482 ( .A(a[840]), .Z(n3521) );
  IV U483 ( .A(b[840]), .Z(n161) );
  NOR U484 ( .A(n3521), .B(n161), .Z(n3523) );
  IV U485 ( .A(a[839]), .Z(n3518) );
  IV U486 ( .A(b[839]), .Z(n162) );
  NOR U487 ( .A(n3518), .B(n162), .Z(n3520) );
  IV U488 ( .A(a[838]), .Z(n3515) );
  IV U489 ( .A(b[838]), .Z(n163) );
  NOR U490 ( .A(n3515), .B(n163), .Z(n3517) );
  IV U491 ( .A(a[837]), .Z(n3512) );
  IV U492 ( .A(b[837]), .Z(n164) );
  NOR U493 ( .A(n3512), .B(n164), .Z(n3514) );
  IV U494 ( .A(a[836]), .Z(n3509) );
  IV U495 ( .A(b[836]), .Z(n165) );
  NOR U496 ( .A(n3509), .B(n165), .Z(n3511) );
  IV U497 ( .A(a[835]), .Z(n3506) );
  IV U498 ( .A(b[835]), .Z(n166) );
  NOR U499 ( .A(n3506), .B(n166), .Z(n3508) );
  IV U500 ( .A(a[834]), .Z(n3503) );
  IV U501 ( .A(b[834]), .Z(n167) );
  NOR U502 ( .A(n3503), .B(n167), .Z(n3505) );
  IV U503 ( .A(a[833]), .Z(n3500) );
  IV U504 ( .A(b[833]), .Z(n168) );
  NOR U505 ( .A(n3500), .B(n168), .Z(n3502) );
  IV U506 ( .A(a[832]), .Z(n3497) );
  IV U507 ( .A(b[832]), .Z(n169) );
  NOR U508 ( .A(n3497), .B(n169), .Z(n3499) );
  IV U509 ( .A(a[831]), .Z(n3494) );
  IV U510 ( .A(b[831]), .Z(n170) );
  NOR U511 ( .A(n3494), .B(n170), .Z(n3496) );
  IV U512 ( .A(a[830]), .Z(n3491) );
  IV U513 ( .A(b[830]), .Z(n171) );
  NOR U514 ( .A(n3491), .B(n171), .Z(n3493) );
  IV U515 ( .A(a[829]), .Z(n3488) );
  IV U516 ( .A(b[829]), .Z(n172) );
  NOR U517 ( .A(n3488), .B(n172), .Z(n3490) );
  IV U518 ( .A(a[828]), .Z(n3485) );
  IV U519 ( .A(b[828]), .Z(n173) );
  NOR U520 ( .A(n3485), .B(n173), .Z(n3487) );
  IV U521 ( .A(a[827]), .Z(n3482) );
  IV U522 ( .A(b[827]), .Z(n174) );
  NOR U523 ( .A(n3482), .B(n174), .Z(n3484) );
  IV U524 ( .A(a[826]), .Z(n3479) );
  IV U525 ( .A(b[826]), .Z(n175) );
  NOR U526 ( .A(n3479), .B(n175), .Z(n3481) );
  IV U527 ( .A(a[825]), .Z(n3476) );
  IV U528 ( .A(b[825]), .Z(n176) );
  NOR U529 ( .A(n3476), .B(n176), .Z(n3478) );
  IV U530 ( .A(a[824]), .Z(n3473) );
  IV U531 ( .A(b[824]), .Z(n177) );
  NOR U532 ( .A(n3473), .B(n177), .Z(n3475) );
  IV U533 ( .A(a[823]), .Z(n3470) );
  IV U534 ( .A(b[823]), .Z(n178) );
  NOR U535 ( .A(n3470), .B(n178), .Z(n3472) );
  IV U536 ( .A(a[822]), .Z(n3467) );
  IV U537 ( .A(b[822]), .Z(n179) );
  NOR U538 ( .A(n3467), .B(n179), .Z(n3469) );
  IV U539 ( .A(a[821]), .Z(n3464) );
  IV U540 ( .A(b[821]), .Z(n180) );
  NOR U541 ( .A(n3464), .B(n180), .Z(n3466) );
  IV U542 ( .A(a[820]), .Z(n3461) );
  IV U543 ( .A(b[820]), .Z(n181) );
  NOR U544 ( .A(n3461), .B(n181), .Z(n3463) );
  IV U545 ( .A(a[819]), .Z(n3458) );
  IV U546 ( .A(b[819]), .Z(n182) );
  NOR U547 ( .A(n3458), .B(n182), .Z(n3460) );
  IV U548 ( .A(a[818]), .Z(n3455) );
  IV U549 ( .A(b[818]), .Z(n183) );
  NOR U550 ( .A(n3455), .B(n183), .Z(n3457) );
  IV U551 ( .A(a[817]), .Z(n3452) );
  IV U552 ( .A(b[817]), .Z(n184) );
  NOR U553 ( .A(n3452), .B(n184), .Z(n3454) );
  IV U554 ( .A(a[816]), .Z(n3449) );
  IV U555 ( .A(b[816]), .Z(n185) );
  NOR U556 ( .A(n3449), .B(n185), .Z(n3451) );
  IV U557 ( .A(a[815]), .Z(n3446) );
  IV U558 ( .A(b[815]), .Z(n186) );
  NOR U559 ( .A(n3446), .B(n186), .Z(n3448) );
  IV U560 ( .A(a[814]), .Z(n3443) );
  IV U561 ( .A(b[814]), .Z(n187) );
  NOR U562 ( .A(n3443), .B(n187), .Z(n3445) );
  IV U563 ( .A(a[813]), .Z(n3440) );
  IV U564 ( .A(b[813]), .Z(n188) );
  NOR U565 ( .A(n3440), .B(n188), .Z(n3442) );
  IV U566 ( .A(a[812]), .Z(n3437) );
  IV U567 ( .A(b[812]), .Z(n189) );
  NOR U568 ( .A(n3437), .B(n189), .Z(n3439) );
  IV U569 ( .A(a[811]), .Z(n3434) );
  IV U570 ( .A(b[811]), .Z(n190) );
  NOR U571 ( .A(n3434), .B(n190), .Z(n3436) );
  IV U572 ( .A(a[810]), .Z(n3431) );
  IV U573 ( .A(b[810]), .Z(n191) );
  NOR U574 ( .A(n3431), .B(n191), .Z(n3433) );
  IV U575 ( .A(a[809]), .Z(n3428) );
  IV U576 ( .A(b[809]), .Z(n192) );
  NOR U577 ( .A(n3428), .B(n192), .Z(n3430) );
  IV U578 ( .A(a[808]), .Z(n3425) );
  IV U579 ( .A(b[808]), .Z(n193) );
  NOR U580 ( .A(n3425), .B(n193), .Z(n3427) );
  IV U581 ( .A(a[807]), .Z(n3422) );
  IV U582 ( .A(b[807]), .Z(n194) );
  NOR U583 ( .A(n3422), .B(n194), .Z(n3424) );
  IV U584 ( .A(a[806]), .Z(n3419) );
  IV U585 ( .A(b[806]), .Z(n195) );
  NOR U586 ( .A(n3419), .B(n195), .Z(n3421) );
  IV U587 ( .A(a[805]), .Z(n3416) );
  IV U588 ( .A(b[805]), .Z(n196) );
  NOR U589 ( .A(n3416), .B(n196), .Z(n3418) );
  IV U590 ( .A(a[804]), .Z(n3413) );
  IV U591 ( .A(b[804]), .Z(n197) );
  NOR U592 ( .A(n3413), .B(n197), .Z(n3415) );
  IV U593 ( .A(a[803]), .Z(n3410) );
  IV U594 ( .A(b[803]), .Z(n198) );
  NOR U595 ( .A(n3410), .B(n198), .Z(n3412) );
  IV U596 ( .A(a[802]), .Z(n3407) );
  IV U597 ( .A(b[802]), .Z(n199) );
  NOR U598 ( .A(n3407), .B(n199), .Z(n3409) );
  IV U599 ( .A(a[801]), .Z(n3404) );
  IV U600 ( .A(b[801]), .Z(n200) );
  NOR U601 ( .A(n3404), .B(n200), .Z(n3406) );
  IV U602 ( .A(a[800]), .Z(n3401) );
  IV U603 ( .A(b[800]), .Z(n201) );
  NOR U604 ( .A(n3401), .B(n201), .Z(n3403) );
  IV U605 ( .A(a[799]), .Z(n3398) );
  IV U606 ( .A(b[799]), .Z(n202) );
  NOR U607 ( .A(n3398), .B(n202), .Z(n3400) );
  IV U608 ( .A(a[798]), .Z(n3395) );
  IV U609 ( .A(b[798]), .Z(n203) );
  NOR U610 ( .A(n3395), .B(n203), .Z(n3397) );
  IV U611 ( .A(a[797]), .Z(n3392) );
  IV U612 ( .A(b[797]), .Z(n204) );
  NOR U613 ( .A(n3392), .B(n204), .Z(n3394) );
  IV U614 ( .A(a[796]), .Z(n3389) );
  IV U615 ( .A(b[796]), .Z(n205) );
  NOR U616 ( .A(n3389), .B(n205), .Z(n3391) );
  IV U617 ( .A(a[795]), .Z(n3386) );
  IV U618 ( .A(b[795]), .Z(n206) );
  NOR U619 ( .A(n3386), .B(n206), .Z(n3388) );
  IV U620 ( .A(a[794]), .Z(n3383) );
  IV U621 ( .A(b[794]), .Z(n207) );
  NOR U622 ( .A(n3383), .B(n207), .Z(n3385) );
  IV U623 ( .A(a[793]), .Z(n3380) );
  IV U624 ( .A(b[793]), .Z(n208) );
  NOR U625 ( .A(n3380), .B(n208), .Z(n3382) );
  IV U626 ( .A(a[792]), .Z(n3377) );
  IV U627 ( .A(b[792]), .Z(n209) );
  NOR U628 ( .A(n3377), .B(n209), .Z(n3379) );
  IV U629 ( .A(a[791]), .Z(n3374) );
  IV U630 ( .A(b[791]), .Z(n210) );
  NOR U631 ( .A(n3374), .B(n210), .Z(n3376) );
  IV U632 ( .A(a[790]), .Z(n3371) );
  IV U633 ( .A(b[790]), .Z(n211) );
  NOR U634 ( .A(n3371), .B(n211), .Z(n3373) );
  IV U635 ( .A(a[789]), .Z(n3368) );
  IV U636 ( .A(b[789]), .Z(n212) );
  NOR U637 ( .A(n3368), .B(n212), .Z(n3370) );
  IV U638 ( .A(a[788]), .Z(n3365) );
  IV U639 ( .A(b[788]), .Z(n213) );
  NOR U640 ( .A(n3365), .B(n213), .Z(n3367) );
  IV U641 ( .A(a[787]), .Z(n3362) );
  IV U642 ( .A(b[787]), .Z(n214) );
  NOR U643 ( .A(n3362), .B(n214), .Z(n3364) );
  IV U644 ( .A(a[786]), .Z(n3359) );
  IV U645 ( .A(b[786]), .Z(n215) );
  NOR U646 ( .A(n3359), .B(n215), .Z(n3361) );
  IV U647 ( .A(a[785]), .Z(n3356) );
  IV U648 ( .A(b[785]), .Z(n216) );
  NOR U649 ( .A(n3356), .B(n216), .Z(n3358) );
  IV U650 ( .A(a[784]), .Z(n3353) );
  IV U651 ( .A(b[784]), .Z(n217) );
  NOR U652 ( .A(n3353), .B(n217), .Z(n3355) );
  IV U653 ( .A(a[783]), .Z(n3350) );
  IV U654 ( .A(b[783]), .Z(n218) );
  NOR U655 ( .A(n3350), .B(n218), .Z(n3352) );
  IV U656 ( .A(a[782]), .Z(n3347) );
  IV U657 ( .A(b[782]), .Z(n219) );
  NOR U658 ( .A(n3347), .B(n219), .Z(n3349) );
  IV U659 ( .A(a[781]), .Z(n3344) );
  IV U660 ( .A(b[781]), .Z(n220) );
  NOR U661 ( .A(n3344), .B(n220), .Z(n3346) );
  IV U662 ( .A(a[780]), .Z(n3341) );
  IV U663 ( .A(b[780]), .Z(n221) );
  NOR U664 ( .A(n3341), .B(n221), .Z(n3343) );
  IV U665 ( .A(a[779]), .Z(n3338) );
  IV U666 ( .A(b[779]), .Z(n222) );
  NOR U667 ( .A(n3338), .B(n222), .Z(n3340) );
  IV U668 ( .A(a[778]), .Z(n3335) );
  IV U669 ( .A(b[778]), .Z(n223) );
  NOR U670 ( .A(n3335), .B(n223), .Z(n3337) );
  IV U671 ( .A(a[777]), .Z(n3332) );
  IV U672 ( .A(b[777]), .Z(n224) );
  NOR U673 ( .A(n3332), .B(n224), .Z(n3334) );
  IV U674 ( .A(a[776]), .Z(n3329) );
  IV U675 ( .A(b[776]), .Z(n225) );
  NOR U676 ( .A(n3329), .B(n225), .Z(n3331) );
  IV U677 ( .A(a[775]), .Z(n3326) );
  IV U678 ( .A(b[775]), .Z(n226) );
  NOR U679 ( .A(n3326), .B(n226), .Z(n3328) );
  IV U680 ( .A(a[774]), .Z(n3323) );
  IV U681 ( .A(b[774]), .Z(n227) );
  NOR U682 ( .A(n3323), .B(n227), .Z(n3325) );
  IV U683 ( .A(a[773]), .Z(n3320) );
  IV U684 ( .A(b[773]), .Z(n228) );
  NOR U685 ( .A(n3320), .B(n228), .Z(n3322) );
  IV U686 ( .A(a[772]), .Z(n3317) );
  IV U687 ( .A(b[772]), .Z(n229) );
  NOR U688 ( .A(n3317), .B(n229), .Z(n3319) );
  IV U689 ( .A(a[771]), .Z(n3314) );
  IV U690 ( .A(b[771]), .Z(n230) );
  NOR U691 ( .A(n3314), .B(n230), .Z(n3316) );
  IV U692 ( .A(a[770]), .Z(n3311) );
  IV U693 ( .A(b[770]), .Z(n231) );
  NOR U694 ( .A(n3311), .B(n231), .Z(n3313) );
  IV U695 ( .A(a[769]), .Z(n3308) );
  IV U696 ( .A(b[769]), .Z(n232) );
  NOR U697 ( .A(n3308), .B(n232), .Z(n3310) );
  IV U698 ( .A(a[768]), .Z(n3305) );
  IV U699 ( .A(b[768]), .Z(n233) );
  NOR U700 ( .A(n3305), .B(n233), .Z(n3307) );
  IV U701 ( .A(a[767]), .Z(n3302) );
  IV U702 ( .A(b[767]), .Z(n234) );
  NOR U703 ( .A(n3302), .B(n234), .Z(n3304) );
  IV U704 ( .A(a[766]), .Z(n3299) );
  IV U705 ( .A(b[766]), .Z(n235) );
  NOR U706 ( .A(n3299), .B(n235), .Z(n3301) );
  IV U707 ( .A(a[765]), .Z(n3296) );
  IV U708 ( .A(b[765]), .Z(n236) );
  NOR U709 ( .A(n3296), .B(n236), .Z(n3298) );
  IV U710 ( .A(a[764]), .Z(n3293) );
  IV U711 ( .A(b[764]), .Z(n237) );
  NOR U712 ( .A(n3293), .B(n237), .Z(n3295) );
  IV U713 ( .A(a[763]), .Z(n3290) );
  IV U714 ( .A(b[763]), .Z(n238) );
  NOR U715 ( .A(n3290), .B(n238), .Z(n3292) );
  IV U716 ( .A(a[762]), .Z(n3287) );
  IV U717 ( .A(b[762]), .Z(n239) );
  NOR U718 ( .A(n3287), .B(n239), .Z(n3289) );
  IV U719 ( .A(a[761]), .Z(n3284) );
  IV U720 ( .A(b[761]), .Z(n240) );
  NOR U721 ( .A(n3284), .B(n240), .Z(n3286) );
  IV U722 ( .A(a[760]), .Z(n3281) );
  IV U723 ( .A(b[760]), .Z(n241) );
  NOR U724 ( .A(n3281), .B(n241), .Z(n3283) );
  IV U725 ( .A(a[759]), .Z(n3278) );
  IV U726 ( .A(b[759]), .Z(n242) );
  NOR U727 ( .A(n3278), .B(n242), .Z(n3280) );
  IV U728 ( .A(a[758]), .Z(n3275) );
  IV U729 ( .A(b[758]), .Z(n243) );
  NOR U730 ( .A(n3275), .B(n243), .Z(n3277) );
  IV U731 ( .A(a[757]), .Z(n3272) );
  IV U732 ( .A(b[757]), .Z(n244) );
  NOR U733 ( .A(n3272), .B(n244), .Z(n3274) );
  IV U734 ( .A(a[756]), .Z(n3269) );
  IV U735 ( .A(b[756]), .Z(n245) );
  NOR U736 ( .A(n3269), .B(n245), .Z(n3271) );
  IV U737 ( .A(a[755]), .Z(n3266) );
  IV U738 ( .A(b[755]), .Z(n246) );
  NOR U739 ( .A(n3266), .B(n246), .Z(n3268) );
  IV U740 ( .A(a[754]), .Z(n3263) );
  IV U741 ( .A(b[754]), .Z(n247) );
  NOR U742 ( .A(n3263), .B(n247), .Z(n3265) );
  IV U743 ( .A(a[753]), .Z(n3260) );
  IV U744 ( .A(b[753]), .Z(n248) );
  NOR U745 ( .A(n3260), .B(n248), .Z(n3262) );
  IV U746 ( .A(a[752]), .Z(n3257) );
  IV U747 ( .A(b[752]), .Z(n249) );
  NOR U748 ( .A(n3257), .B(n249), .Z(n3259) );
  IV U749 ( .A(a[751]), .Z(n3254) );
  IV U750 ( .A(b[751]), .Z(n250) );
  NOR U751 ( .A(n3254), .B(n250), .Z(n3256) );
  IV U752 ( .A(a[750]), .Z(n3251) );
  IV U753 ( .A(b[750]), .Z(n251) );
  NOR U754 ( .A(n3251), .B(n251), .Z(n3253) );
  IV U755 ( .A(a[749]), .Z(n3248) );
  IV U756 ( .A(b[749]), .Z(n252) );
  NOR U757 ( .A(n3248), .B(n252), .Z(n3250) );
  IV U758 ( .A(a[748]), .Z(n3245) );
  IV U759 ( .A(b[748]), .Z(n253) );
  NOR U760 ( .A(n3245), .B(n253), .Z(n3247) );
  IV U761 ( .A(a[747]), .Z(n3242) );
  IV U762 ( .A(b[747]), .Z(n254) );
  NOR U763 ( .A(n3242), .B(n254), .Z(n3244) );
  IV U764 ( .A(a[746]), .Z(n3239) );
  IV U765 ( .A(b[746]), .Z(n255) );
  NOR U766 ( .A(n3239), .B(n255), .Z(n3241) );
  IV U767 ( .A(a[745]), .Z(n3236) );
  IV U768 ( .A(b[745]), .Z(n256) );
  NOR U769 ( .A(n3236), .B(n256), .Z(n3238) );
  IV U770 ( .A(a[744]), .Z(n3233) );
  IV U771 ( .A(b[744]), .Z(n257) );
  NOR U772 ( .A(n3233), .B(n257), .Z(n3235) );
  IV U773 ( .A(a[743]), .Z(n3230) );
  IV U774 ( .A(b[743]), .Z(n258) );
  NOR U775 ( .A(n3230), .B(n258), .Z(n3232) );
  IV U776 ( .A(a[742]), .Z(n3227) );
  IV U777 ( .A(b[742]), .Z(n259) );
  NOR U778 ( .A(n3227), .B(n259), .Z(n3229) );
  IV U779 ( .A(a[741]), .Z(n3224) );
  IV U780 ( .A(b[741]), .Z(n260) );
  NOR U781 ( .A(n3224), .B(n260), .Z(n3226) );
  IV U782 ( .A(a[740]), .Z(n3221) );
  IV U783 ( .A(b[740]), .Z(n261) );
  NOR U784 ( .A(n3221), .B(n261), .Z(n3223) );
  IV U785 ( .A(a[739]), .Z(n3218) );
  IV U786 ( .A(b[739]), .Z(n262) );
  NOR U787 ( .A(n3218), .B(n262), .Z(n3220) );
  IV U788 ( .A(a[738]), .Z(n3215) );
  IV U789 ( .A(b[738]), .Z(n263) );
  NOR U790 ( .A(n3215), .B(n263), .Z(n3217) );
  IV U791 ( .A(a[737]), .Z(n3212) );
  IV U792 ( .A(b[737]), .Z(n264) );
  NOR U793 ( .A(n3212), .B(n264), .Z(n3214) );
  IV U794 ( .A(a[736]), .Z(n3209) );
  IV U795 ( .A(b[736]), .Z(n265) );
  NOR U796 ( .A(n3209), .B(n265), .Z(n3211) );
  IV U797 ( .A(a[735]), .Z(n3206) );
  IV U798 ( .A(b[735]), .Z(n266) );
  NOR U799 ( .A(n3206), .B(n266), .Z(n3208) );
  IV U800 ( .A(a[734]), .Z(n3203) );
  IV U801 ( .A(b[734]), .Z(n267) );
  NOR U802 ( .A(n3203), .B(n267), .Z(n3205) );
  IV U803 ( .A(a[733]), .Z(n3200) );
  IV U804 ( .A(b[733]), .Z(n268) );
  NOR U805 ( .A(n3200), .B(n268), .Z(n3202) );
  IV U806 ( .A(a[732]), .Z(n3197) );
  IV U807 ( .A(b[732]), .Z(n269) );
  NOR U808 ( .A(n3197), .B(n269), .Z(n3199) );
  IV U809 ( .A(a[731]), .Z(n3194) );
  IV U810 ( .A(b[731]), .Z(n270) );
  NOR U811 ( .A(n3194), .B(n270), .Z(n3196) );
  IV U812 ( .A(a[730]), .Z(n3191) );
  IV U813 ( .A(b[730]), .Z(n271) );
  NOR U814 ( .A(n3191), .B(n271), .Z(n3193) );
  IV U815 ( .A(a[729]), .Z(n3188) );
  IV U816 ( .A(b[729]), .Z(n272) );
  NOR U817 ( .A(n3188), .B(n272), .Z(n3190) );
  IV U818 ( .A(a[728]), .Z(n3185) );
  IV U819 ( .A(b[728]), .Z(n273) );
  NOR U820 ( .A(n3185), .B(n273), .Z(n3187) );
  IV U821 ( .A(a[727]), .Z(n3182) );
  IV U822 ( .A(b[727]), .Z(n274) );
  NOR U823 ( .A(n3182), .B(n274), .Z(n3184) );
  IV U824 ( .A(a[726]), .Z(n3179) );
  IV U825 ( .A(b[726]), .Z(n275) );
  NOR U826 ( .A(n3179), .B(n275), .Z(n3181) );
  IV U827 ( .A(a[725]), .Z(n3176) );
  IV U828 ( .A(b[725]), .Z(n276) );
  NOR U829 ( .A(n3176), .B(n276), .Z(n3178) );
  IV U830 ( .A(a[724]), .Z(n3173) );
  IV U831 ( .A(b[724]), .Z(n277) );
  NOR U832 ( .A(n3173), .B(n277), .Z(n3175) );
  IV U833 ( .A(a[723]), .Z(n3170) );
  IV U834 ( .A(b[723]), .Z(n278) );
  NOR U835 ( .A(n3170), .B(n278), .Z(n3172) );
  IV U836 ( .A(a[722]), .Z(n3167) );
  IV U837 ( .A(b[722]), .Z(n279) );
  NOR U838 ( .A(n3167), .B(n279), .Z(n3169) );
  IV U839 ( .A(a[721]), .Z(n3164) );
  IV U840 ( .A(b[721]), .Z(n280) );
  NOR U841 ( .A(n3164), .B(n280), .Z(n3166) );
  IV U842 ( .A(a[720]), .Z(n3161) );
  IV U843 ( .A(b[720]), .Z(n281) );
  NOR U844 ( .A(n3161), .B(n281), .Z(n3163) );
  IV U845 ( .A(a[719]), .Z(n3158) );
  IV U846 ( .A(b[719]), .Z(n282) );
  NOR U847 ( .A(n3158), .B(n282), .Z(n3160) );
  IV U848 ( .A(a[718]), .Z(n3155) );
  IV U849 ( .A(b[718]), .Z(n283) );
  NOR U850 ( .A(n3155), .B(n283), .Z(n3157) );
  IV U851 ( .A(a[717]), .Z(n3152) );
  IV U852 ( .A(b[717]), .Z(n284) );
  NOR U853 ( .A(n3152), .B(n284), .Z(n3154) );
  IV U854 ( .A(a[716]), .Z(n3149) );
  IV U855 ( .A(b[716]), .Z(n285) );
  NOR U856 ( .A(n3149), .B(n285), .Z(n3151) );
  IV U857 ( .A(a[715]), .Z(n3146) );
  IV U858 ( .A(b[715]), .Z(n286) );
  NOR U859 ( .A(n3146), .B(n286), .Z(n3148) );
  IV U860 ( .A(a[714]), .Z(n3143) );
  IV U861 ( .A(b[714]), .Z(n287) );
  NOR U862 ( .A(n3143), .B(n287), .Z(n3145) );
  IV U863 ( .A(a[713]), .Z(n3140) );
  IV U864 ( .A(b[713]), .Z(n288) );
  NOR U865 ( .A(n3140), .B(n288), .Z(n3142) );
  IV U866 ( .A(a[712]), .Z(n3137) );
  IV U867 ( .A(b[712]), .Z(n289) );
  NOR U868 ( .A(n3137), .B(n289), .Z(n3139) );
  IV U869 ( .A(a[711]), .Z(n3134) );
  IV U870 ( .A(b[711]), .Z(n290) );
  NOR U871 ( .A(n3134), .B(n290), .Z(n3136) );
  IV U872 ( .A(a[710]), .Z(n3131) );
  IV U873 ( .A(b[710]), .Z(n291) );
  NOR U874 ( .A(n3131), .B(n291), .Z(n3133) );
  IV U875 ( .A(a[709]), .Z(n3128) );
  IV U876 ( .A(b[709]), .Z(n292) );
  NOR U877 ( .A(n3128), .B(n292), .Z(n3130) );
  IV U878 ( .A(a[708]), .Z(n3125) );
  IV U879 ( .A(b[708]), .Z(n293) );
  NOR U880 ( .A(n3125), .B(n293), .Z(n3127) );
  IV U881 ( .A(a[707]), .Z(n3122) );
  IV U882 ( .A(b[707]), .Z(n294) );
  NOR U883 ( .A(n3122), .B(n294), .Z(n3124) );
  IV U884 ( .A(a[706]), .Z(n3119) );
  IV U885 ( .A(b[706]), .Z(n295) );
  NOR U886 ( .A(n3119), .B(n295), .Z(n3121) );
  IV U887 ( .A(a[705]), .Z(n3116) );
  IV U888 ( .A(b[705]), .Z(n296) );
  NOR U889 ( .A(n3116), .B(n296), .Z(n3118) );
  IV U890 ( .A(a[704]), .Z(n3113) );
  IV U891 ( .A(b[704]), .Z(n297) );
  NOR U892 ( .A(n3113), .B(n297), .Z(n3115) );
  IV U893 ( .A(a[703]), .Z(n3110) );
  IV U894 ( .A(b[703]), .Z(n298) );
  NOR U895 ( .A(n3110), .B(n298), .Z(n3112) );
  IV U896 ( .A(a[702]), .Z(n3107) );
  IV U897 ( .A(b[702]), .Z(n299) );
  NOR U898 ( .A(n3107), .B(n299), .Z(n3109) );
  IV U899 ( .A(a[701]), .Z(n3104) );
  IV U900 ( .A(b[701]), .Z(n300) );
  NOR U901 ( .A(n3104), .B(n300), .Z(n3106) );
  IV U902 ( .A(a[700]), .Z(n3101) );
  IV U903 ( .A(b[700]), .Z(n301) );
  NOR U904 ( .A(n3101), .B(n301), .Z(n3103) );
  IV U905 ( .A(a[699]), .Z(n3098) );
  IV U906 ( .A(b[699]), .Z(n302) );
  NOR U907 ( .A(n3098), .B(n302), .Z(n3100) );
  IV U908 ( .A(a[698]), .Z(n3095) );
  IV U909 ( .A(b[698]), .Z(n303) );
  NOR U910 ( .A(n3095), .B(n303), .Z(n3097) );
  IV U911 ( .A(a[697]), .Z(n3092) );
  IV U912 ( .A(b[697]), .Z(n304) );
  NOR U913 ( .A(n3092), .B(n304), .Z(n3094) );
  IV U914 ( .A(a[696]), .Z(n3089) );
  IV U915 ( .A(b[696]), .Z(n305) );
  NOR U916 ( .A(n3089), .B(n305), .Z(n3091) );
  IV U917 ( .A(a[695]), .Z(n3086) );
  IV U918 ( .A(b[695]), .Z(n306) );
  NOR U919 ( .A(n3086), .B(n306), .Z(n3088) );
  IV U920 ( .A(a[694]), .Z(n3083) );
  IV U921 ( .A(b[694]), .Z(n307) );
  NOR U922 ( .A(n3083), .B(n307), .Z(n3085) );
  IV U923 ( .A(a[693]), .Z(n3080) );
  IV U924 ( .A(b[693]), .Z(n308) );
  NOR U925 ( .A(n3080), .B(n308), .Z(n3082) );
  IV U926 ( .A(a[692]), .Z(n3077) );
  IV U927 ( .A(b[692]), .Z(n309) );
  NOR U928 ( .A(n3077), .B(n309), .Z(n3079) );
  IV U929 ( .A(a[691]), .Z(n3074) );
  IV U930 ( .A(b[691]), .Z(n310) );
  NOR U931 ( .A(n3074), .B(n310), .Z(n3076) );
  IV U932 ( .A(a[690]), .Z(n3071) );
  IV U933 ( .A(b[690]), .Z(n311) );
  NOR U934 ( .A(n3071), .B(n311), .Z(n3073) );
  IV U935 ( .A(a[689]), .Z(n3068) );
  IV U936 ( .A(b[689]), .Z(n312) );
  NOR U937 ( .A(n3068), .B(n312), .Z(n3070) );
  IV U938 ( .A(a[688]), .Z(n3065) );
  IV U939 ( .A(b[688]), .Z(n313) );
  NOR U940 ( .A(n3065), .B(n313), .Z(n3067) );
  IV U941 ( .A(a[687]), .Z(n3062) );
  IV U942 ( .A(b[687]), .Z(n314) );
  NOR U943 ( .A(n3062), .B(n314), .Z(n3064) );
  IV U944 ( .A(a[686]), .Z(n3059) );
  IV U945 ( .A(b[686]), .Z(n315) );
  NOR U946 ( .A(n3059), .B(n315), .Z(n3061) );
  IV U947 ( .A(a[685]), .Z(n3056) );
  IV U948 ( .A(b[685]), .Z(n316) );
  NOR U949 ( .A(n3056), .B(n316), .Z(n3058) );
  IV U950 ( .A(a[684]), .Z(n3053) );
  IV U951 ( .A(b[684]), .Z(n317) );
  NOR U952 ( .A(n3053), .B(n317), .Z(n3055) );
  IV U953 ( .A(a[683]), .Z(n3050) );
  IV U954 ( .A(b[683]), .Z(n318) );
  NOR U955 ( .A(n3050), .B(n318), .Z(n3052) );
  IV U956 ( .A(a[682]), .Z(n3047) );
  IV U957 ( .A(b[682]), .Z(n319) );
  NOR U958 ( .A(n3047), .B(n319), .Z(n3049) );
  IV U959 ( .A(a[681]), .Z(n3044) );
  IV U960 ( .A(b[681]), .Z(n320) );
  NOR U961 ( .A(n3044), .B(n320), .Z(n3046) );
  IV U962 ( .A(a[680]), .Z(n3041) );
  IV U963 ( .A(b[680]), .Z(n321) );
  NOR U964 ( .A(n3041), .B(n321), .Z(n3043) );
  IV U965 ( .A(a[679]), .Z(n3038) );
  IV U966 ( .A(b[679]), .Z(n322) );
  NOR U967 ( .A(n3038), .B(n322), .Z(n3040) );
  IV U968 ( .A(a[678]), .Z(n3035) );
  IV U969 ( .A(b[678]), .Z(n323) );
  NOR U970 ( .A(n3035), .B(n323), .Z(n3037) );
  IV U971 ( .A(a[677]), .Z(n3032) );
  IV U972 ( .A(b[677]), .Z(n324) );
  NOR U973 ( .A(n3032), .B(n324), .Z(n3034) );
  IV U974 ( .A(a[676]), .Z(n3029) );
  IV U975 ( .A(b[676]), .Z(n325) );
  NOR U976 ( .A(n3029), .B(n325), .Z(n3031) );
  IV U977 ( .A(a[675]), .Z(n3026) );
  IV U978 ( .A(b[675]), .Z(n326) );
  NOR U979 ( .A(n3026), .B(n326), .Z(n3028) );
  IV U980 ( .A(a[674]), .Z(n3023) );
  IV U981 ( .A(b[674]), .Z(n327) );
  NOR U982 ( .A(n3023), .B(n327), .Z(n3025) );
  IV U983 ( .A(a[673]), .Z(n3020) );
  IV U984 ( .A(b[673]), .Z(n328) );
  NOR U985 ( .A(n3020), .B(n328), .Z(n3022) );
  IV U986 ( .A(a[672]), .Z(n3017) );
  IV U987 ( .A(b[672]), .Z(n329) );
  NOR U988 ( .A(n3017), .B(n329), .Z(n3019) );
  IV U989 ( .A(a[671]), .Z(n3014) );
  IV U990 ( .A(b[671]), .Z(n330) );
  NOR U991 ( .A(n3014), .B(n330), .Z(n3016) );
  IV U992 ( .A(a[670]), .Z(n3011) );
  IV U993 ( .A(b[670]), .Z(n331) );
  NOR U994 ( .A(n3011), .B(n331), .Z(n3013) );
  IV U995 ( .A(a[669]), .Z(n3008) );
  IV U996 ( .A(b[669]), .Z(n332) );
  NOR U997 ( .A(n3008), .B(n332), .Z(n3010) );
  IV U998 ( .A(a[668]), .Z(n3005) );
  IV U999 ( .A(b[668]), .Z(n333) );
  NOR U1000 ( .A(n3005), .B(n333), .Z(n3007) );
  IV U1001 ( .A(a[667]), .Z(n3002) );
  IV U1002 ( .A(b[667]), .Z(n334) );
  NOR U1003 ( .A(n3002), .B(n334), .Z(n3004) );
  IV U1004 ( .A(a[666]), .Z(n2999) );
  IV U1005 ( .A(b[666]), .Z(n335) );
  NOR U1006 ( .A(n2999), .B(n335), .Z(n3001) );
  IV U1007 ( .A(a[665]), .Z(n2996) );
  IV U1008 ( .A(b[665]), .Z(n336) );
  NOR U1009 ( .A(n2996), .B(n336), .Z(n2998) );
  IV U1010 ( .A(a[664]), .Z(n2993) );
  IV U1011 ( .A(b[664]), .Z(n337) );
  NOR U1012 ( .A(n2993), .B(n337), .Z(n2995) );
  IV U1013 ( .A(a[663]), .Z(n2990) );
  IV U1014 ( .A(b[663]), .Z(n338) );
  NOR U1015 ( .A(n2990), .B(n338), .Z(n2992) );
  IV U1016 ( .A(a[662]), .Z(n2987) );
  IV U1017 ( .A(b[662]), .Z(n339) );
  NOR U1018 ( .A(n2987), .B(n339), .Z(n2989) );
  IV U1019 ( .A(a[661]), .Z(n2984) );
  IV U1020 ( .A(b[661]), .Z(n340) );
  NOR U1021 ( .A(n2984), .B(n340), .Z(n2986) );
  IV U1022 ( .A(a[660]), .Z(n2981) );
  IV U1023 ( .A(b[660]), .Z(n341) );
  NOR U1024 ( .A(n2981), .B(n341), .Z(n2983) );
  IV U1025 ( .A(a[659]), .Z(n2978) );
  IV U1026 ( .A(b[659]), .Z(n342) );
  NOR U1027 ( .A(n2978), .B(n342), .Z(n2980) );
  IV U1028 ( .A(a[658]), .Z(n2975) );
  IV U1029 ( .A(b[658]), .Z(n343) );
  NOR U1030 ( .A(n2975), .B(n343), .Z(n2977) );
  IV U1031 ( .A(a[657]), .Z(n2972) );
  IV U1032 ( .A(b[657]), .Z(n344) );
  NOR U1033 ( .A(n2972), .B(n344), .Z(n2974) );
  IV U1034 ( .A(a[656]), .Z(n2969) );
  IV U1035 ( .A(b[656]), .Z(n345) );
  NOR U1036 ( .A(n2969), .B(n345), .Z(n2971) );
  IV U1037 ( .A(a[655]), .Z(n2966) );
  IV U1038 ( .A(b[655]), .Z(n346) );
  NOR U1039 ( .A(n2966), .B(n346), .Z(n2968) );
  IV U1040 ( .A(a[654]), .Z(n2963) );
  IV U1041 ( .A(b[654]), .Z(n347) );
  NOR U1042 ( .A(n2963), .B(n347), .Z(n2965) );
  IV U1043 ( .A(a[653]), .Z(n2960) );
  IV U1044 ( .A(b[653]), .Z(n348) );
  NOR U1045 ( .A(n2960), .B(n348), .Z(n2962) );
  IV U1046 ( .A(a[652]), .Z(n2957) );
  IV U1047 ( .A(b[652]), .Z(n349) );
  NOR U1048 ( .A(n2957), .B(n349), .Z(n2959) );
  IV U1049 ( .A(a[651]), .Z(n2954) );
  IV U1050 ( .A(b[651]), .Z(n350) );
  NOR U1051 ( .A(n2954), .B(n350), .Z(n2956) );
  IV U1052 ( .A(a[650]), .Z(n2951) );
  IV U1053 ( .A(b[650]), .Z(n351) );
  NOR U1054 ( .A(n2951), .B(n351), .Z(n2953) );
  IV U1055 ( .A(a[649]), .Z(n2948) );
  IV U1056 ( .A(b[649]), .Z(n352) );
  NOR U1057 ( .A(n2948), .B(n352), .Z(n2950) );
  IV U1058 ( .A(a[648]), .Z(n2945) );
  IV U1059 ( .A(b[648]), .Z(n353) );
  NOR U1060 ( .A(n2945), .B(n353), .Z(n2947) );
  IV U1061 ( .A(a[647]), .Z(n2942) );
  IV U1062 ( .A(b[647]), .Z(n354) );
  NOR U1063 ( .A(n2942), .B(n354), .Z(n2944) );
  IV U1064 ( .A(a[646]), .Z(n2939) );
  IV U1065 ( .A(b[646]), .Z(n355) );
  NOR U1066 ( .A(n2939), .B(n355), .Z(n2941) );
  IV U1067 ( .A(a[645]), .Z(n2936) );
  IV U1068 ( .A(b[645]), .Z(n356) );
  NOR U1069 ( .A(n2936), .B(n356), .Z(n2938) );
  IV U1070 ( .A(a[644]), .Z(n2933) );
  IV U1071 ( .A(b[644]), .Z(n357) );
  NOR U1072 ( .A(n2933), .B(n357), .Z(n2935) );
  IV U1073 ( .A(a[643]), .Z(n2930) );
  IV U1074 ( .A(b[643]), .Z(n358) );
  NOR U1075 ( .A(n2930), .B(n358), .Z(n2932) );
  IV U1076 ( .A(a[642]), .Z(n2927) );
  IV U1077 ( .A(b[642]), .Z(n359) );
  NOR U1078 ( .A(n2927), .B(n359), .Z(n2929) );
  IV U1079 ( .A(a[641]), .Z(n2924) );
  IV U1080 ( .A(b[641]), .Z(n360) );
  NOR U1081 ( .A(n2924), .B(n360), .Z(n2926) );
  IV U1082 ( .A(a[640]), .Z(n2921) );
  IV U1083 ( .A(b[640]), .Z(n361) );
  NOR U1084 ( .A(n2921), .B(n361), .Z(n2923) );
  IV U1085 ( .A(a[639]), .Z(n2918) );
  IV U1086 ( .A(b[639]), .Z(n362) );
  NOR U1087 ( .A(n2918), .B(n362), .Z(n2920) );
  IV U1088 ( .A(a[638]), .Z(n2915) );
  IV U1089 ( .A(b[638]), .Z(n363) );
  NOR U1090 ( .A(n2915), .B(n363), .Z(n2917) );
  IV U1091 ( .A(a[637]), .Z(n2912) );
  IV U1092 ( .A(b[637]), .Z(n364) );
  NOR U1093 ( .A(n2912), .B(n364), .Z(n2914) );
  IV U1094 ( .A(a[636]), .Z(n2909) );
  IV U1095 ( .A(b[636]), .Z(n365) );
  NOR U1096 ( .A(n2909), .B(n365), .Z(n2911) );
  IV U1097 ( .A(a[635]), .Z(n2906) );
  IV U1098 ( .A(b[635]), .Z(n366) );
  NOR U1099 ( .A(n2906), .B(n366), .Z(n2908) );
  IV U1100 ( .A(a[634]), .Z(n2903) );
  IV U1101 ( .A(b[634]), .Z(n367) );
  NOR U1102 ( .A(n2903), .B(n367), .Z(n2905) );
  IV U1103 ( .A(a[633]), .Z(n2900) );
  IV U1104 ( .A(b[633]), .Z(n368) );
  NOR U1105 ( .A(n2900), .B(n368), .Z(n2902) );
  IV U1106 ( .A(a[632]), .Z(n2897) );
  IV U1107 ( .A(b[632]), .Z(n369) );
  NOR U1108 ( .A(n2897), .B(n369), .Z(n2899) );
  IV U1109 ( .A(a[631]), .Z(n2894) );
  IV U1110 ( .A(b[631]), .Z(n370) );
  NOR U1111 ( .A(n2894), .B(n370), .Z(n2896) );
  IV U1112 ( .A(a[630]), .Z(n2891) );
  IV U1113 ( .A(b[630]), .Z(n371) );
  NOR U1114 ( .A(n2891), .B(n371), .Z(n2893) );
  IV U1115 ( .A(a[629]), .Z(n2888) );
  IV U1116 ( .A(b[629]), .Z(n372) );
  NOR U1117 ( .A(n2888), .B(n372), .Z(n2890) );
  IV U1118 ( .A(a[628]), .Z(n2885) );
  IV U1119 ( .A(b[628]), .Z(n373) );
  NOR U1120 ( .A(n2885), .B(n373), .Z(n2887) );
  IV U1121 ( .A(a[627]), .Z(n2882) );
  IV U1122 ( .A(b[627]), .Z(n374) );
  NOR U1123 ( .A(n2882), .B(n374), .Z(n2884) );
  IV U1124 ( .A(a[626]), .Z(n2879) );
  IV U1125 ( .A(b[626]), .Z(n375) );
  NOR U1126 ( .A(n2879), .B(n375), .Z(n2881) );
  IV U1127 ( .A(a[625]), .Z(n2876) );
  IV U1128 ( .A(b[625]), .Z(n376) );
  NOR U1129 ( .A(n2876), .B(n376), .Z(n2878) );
  IV U1130 ( .A(a[624]), .Z(n2873) );
  IV U1131 ( .A(b[624]), .Z(n377) );
  NOR U1132 ( .A(n2873), .B(n377), .Z(n2875) );
  IV U1133 ( .A(a[623]), .Z(n2870) );
  IV U1134 ( .A(b[623]), .Z(n378) );
  NOR U1135 ( .A(n2870), .B(n378), .Z(n2872) );
  IV U1136 ( .A(a[622]), .Z(n2867) );
  IV U1137 ( .A(b[622]), .Z(n379) );
  NOR U1138 ( .A(n2867), .B(n379), .Z(n2869) );
  IV U1139 ( .A(a[621]), .Z(n2864) );
  IV U1140 ( .A(b[621]), .Z(n380) );
  NOR U1141 ( .A(n2864), .B(n380), .Z(n2866) );
  IV U1142 ( .A(a[620]), .Z(n2861) );
  IV U1143 ( .A(b[620]), .Z(n381) );
  NOR U1144 ( .A(n2861), .B(n381), .Z(n2863) );
  IV U1145 ( .A(a[619]), .Z(n2858) );
  IV U1146 ( .A(b[619]), .Z(n382) );
  NOR U1147 ( .A(n2858), .B(n382), .Z(n2860) );
  IV U1148 ( .A(a[618]), .Z(n2855) );
  IV U1149 ( .A(b[618]), .Z(n383) );
  NOR U1150 ( .A(n2855), .B(n383), .Z(n2857) );
  IV U1151 ( .A(a[617]), .Z(n2852) );
  IV U1152 ( .A(b[617]), .Z(n384) );
  NOR U1153 ( .A(n2852), .B(n384), .Z(n2854) );
  IV U1154 ( .A(a[616]), .Z(n2849) );
  IV U1155 ( .A(b[616]), .Z(n385) );
  NOR U1156 ( .A(n2849), .B(n385), .Z(n2851) );
  IV U1157 ( .A(a[615]), .Z(n2846) );
  IV U1158 ( .A(b[615]), .Z(n386) );
  NOR U1159 ( .A(n2846), .B(n386), .Z(n2848) );
  IV U1160 ( .A(a[614]), .Z(n2843) );
  IV U1161 ( .A(b[614]), .Z(n387) );
  NOR U1162 ( .A(n2843), .B(n387), .Z(n2845) );
  IV U1163 ( .A(a[613]), .Z(n2840) );
  IV U1164 ( .A(b[613]), .Z(n388) );
  NOR U1165 ( .A(n2840), .B(n388), .Z(n2842) );
  IV U1166 ( .A(a[612]), .Z(n2837) );
  IV U1167 ( .A(b[612]), .Z(n389) );
  NOR U1168 ( .A(n2837), .B(n389), .Z(n2839) );
  IV U1169 ( .A(a[611]), .Z(n2834) );
  IV U1170 ( .A(b[611]), .Z(n390) );
  NOR U1171 ( .A(n2834), .B(n390), .Z(n2836) );
  IV U1172 ( .A(a[610]), .Z(n2831) );
  IV U1173 ( .A(b[610]), .Z(n391) );
  NOR U1174 ( .A(n2831), .B(n391), .Z(n2833) );
  IV U1175 ( .A(a[609]), .Z(n2828) );
  IV U1176 ( .A(b[609]), .Z(n392) );
  NOR U1177 ( .A(n2828), .B(n392), .Z(n2830) );
  IV U1178 ( .A(a[608]), .Z(n2825) );
  IV U1179 ( .A(b[608]), .Z(n393) );
  NOR U1180 ( .A(n2825), .B(n393), .Z(n2827) );
  IV U1181 ( .A(a[607]), .Z(n2822) );
  IV U1182 ( .A(b[607]), .Z(n394) );
  NOR U1183 ( .A(n2822), .B(n394), .Z(n2824) );
  IV U1184 ( .A(a[606]), .Z(n2819) );
  IV U1185 ( .A(b[606]), .Z(n395) );
  NOR U1186 ( .A(n2819), .B(n395), .Z(n2821) );
  IV U1187 ( .A(a[605]), .Z(n2816) );
  IV U1188 ( .A(b[605]), .Z(n396) );
  NOR U1189 ( .A(n2816), .B(n396), .Z(n2818) );
  IV U1190 ( .A(a[604]), .Z(n2813) );
  IV U1191 ( .A(b[604]), .Z(n397) );
  NOR U1192 ( .A(n2813), .B(n397), .Z(n2815) );
  IV U1193 ( .A(a[603]), .Z(n2810) );
  IV U1194 ( .A(b[603]), .Z(n398) );
  NOR U1195 ( .A(n2810), .B(n398), .Z(n2812) );
  IV U1196 ( .A(a[602]), .Z(n2807) );
  IV U1197 ( .A(b[602]), .Z(n399) );
  NOR U1198 ( .A(n2807), .B(n399), .Z(n2809) );
  IV U1199 ( .A(a[601]), .Z(n2804) );
  IV U1200 ( .A(b[601]), .Z(n400) );
  NOR U1201 ( .A(n2804), .B(n400), .Z(n2806) );
  IV U1202 ( .A(a[600]), .Z(n2801) );
  IV U1203 ( .A(b[600]), .Z(n401) );
  NOR U1204 ( .A(n2801), .B(n401), .Z(n2803) );
  IV U1205 ( .A(a[599]), .Z(n2798) );
  IV U1206 ( .A(b[599]), .Z(n402) );
  NOR U1207 ( .A(n2798), .B(n402), .Z(n2800) );
  IV U1208 ( .A(a[598]), .Z(n2795) );
  IV U1209 ( .A(b[598]), .Z(n403) );
  NOR U1210 ( .A(n2795), .B(n403), .Z(n2797) );
  IV U1211 ( .A(a[597]), .Z(n2792) );
  IV U1212 ( .A(b[597]), .Z(n404) );
  NOR U1213 ( .A(n2792), .B(n404), .Z(n2794) );
  IV U1214 ( .A(a[596]), .Z(n2789) );
  IV U1215 ( .A(b[596]), .Z(n405) );
  NOR U1216 ( .A(n2789), .B(n405), .Z(n2791) );
  IV U1217 ( .A(a[595]), .Z(n2786) );
  IV U1218 ( .A(b[595]), .Z(n406) );
  NOR U1219 ( .A(n2786), .B(n406), .Z(n2788) );
  IV U1220 ( .A(a[594]), .Z(n2783) );
  IV U1221 ( .A(b[594]), .Z(n407) );
  NOR U1222 ( .A(n2783), .B(n407), .Z(n2785) );
  IV U1223 ( .A(a[593]), .Z(n2780) );
  IV U1224 ( .A(b[593]), .Z(n408) );
  NOR U1225 ( .A(n2780), .B(n408), .Z(n2782) );
  IV U1226 ( .A(a[592]), .Z(n2777) );
  IV U1227 ( .A(b[592]), .Z(n409) );
  NOR U1228 ( .A(n2777), .B(n409), .Z(n2779) );
  IV U1229 ( .A(a[591]), .Z(n2774) );
  IV U1230 ( .A(b[591]), .Z(n410) );
  NOR U1231 ( .A(n2774), .B(n410), .Z(n2776) );
  IV U1232 ( .A(a[590]), .Z(n2771) );
  IV U1233 ( .A(b[590]), .Z(n411) );
  NOR U1234 ( .A(n2771), .B(n411), .Z(n2773) );
  IV U1235 ( .A(a[589]), .Z(n2768) );
  IV U1236 ( .A(b[589]), .Z(n412) );
  NOR U1237 ( .A(n2768), .B(n412), .Z(n2770) );
  IV U1238 ( .A(a[588]), .Z(n2765) );
  IV U1239 ( .A(b[588]), .Z(n413) );
  NOR U1240 ( .A(n2765), .B(n413), .Z(n2767) );
  IV U1241 ( .A(a[587]), .Z(n2762) );
  IV U1242 ( .A(b[587]), .Z(n414) );
  NOR U1243 ( .A(n2762), .B(n414), .Z(n2764) );
  IV U1244 ( .A(a[586]), .Z(n2759) );
  IV U1245 ( .A(b[586]), .Z(n415) );
  NOR U1246 ( .A(n2759), .B(n415), .Z(n2761) );
  IV U1247 ( .A(a[585]), .Z(n2756) );
  IV U1248 ( .A(b[585]), .Z(n416) );
  NOR U1249 ( .A(n2756), .B(n416), .Z(n2758) );
  IV U1250 ( .A(a[584]), .Z(n2753) );
  IV U1251 ( .A(b[584]), .Z(n417) );
  NOR U1252 ( .A(n2753), .B(n417), .Z(n2755) );
  IV U1253 ( .A(a[583]), .Z(n2750) );
  IV U1254 ( .A(b[583]), .Z(n418) );
  NOR U1255 ( .A(n2750), .B(n418), .Z(n2752) );
  IV U1256 ( .A(a[582]), .Z(n2747) );
  IV U1257 ( .A(b[582]), .Z(n419) );
  NOR U1258 ( .A(n2747), .B(n419), .Z(n2749) );
  IV U1259 ( .A(a[581]), .Z(n2744) );
  IV U1260 ( .A(b[581]), .Z(n420) );
  NOR U1261 ( .A(n2744), .B(n420), .Z(n2746) );
  IV U1262 ( .A(a[580]), .Z(n2741) );
  IV U1263 ( .A(b[580]), .Z(n421) );
  NOR U1264 ( .A(n2741), .B(n421), .Z(n2743) );
  IV U1265 ( .A(a[579]), .Z(n2738) );
  IV U1266 ( .A(b[579]), .Z(n422) );
  NOR U1267 ( .A(n2738), .B(n422), .Z(n2740) );
  IV U1268 ( .A(a[578]), .Z(n2735) );
  IV U1269 ( .A(b[578]), .Z(n423) );
  NOR U1270 ( .A(n2735), .B(n423), .Z(n2737) );
  IV U1271 ( .A(a[577]), .Z(n2732) );
  IV U1272 ( .A(b[577]), .Z(n424) );
  NOR U1273 ( .A(n2732), .B(n424), .Z(n2734) );
  IV U1274 ( .A(a[576]), .Z(n2729) );
  IV U1275 ( .A(b[576]), .Z(n425) );
  NOR U1276 ( .A(n2729), .B(n425), .Z(n2731) );
  IV U1277 ( .A(a[575]), .Z(n2726) );
  IV U1278 ( .A(b[575]), .Z(n426) );
  NOR U1279 ( .A(n2726), .B(n426), .Z(n2728) );
  IV U1280 ( .A(a[574]), .Z(n2723) );
  IV U1281 ( .A(b[574]), .Z(n427) );
  NOR U1282 ( .A(n2723), .B(n427), .Z(n2725) );
  IV U1283 ( .A(a[573]), .Z(n2720) );
  IV U1284 ( .A(b[573]), .Z(n428) );
  NOR U1285 ( .A(n2720), .B(n428), .Z(n2722) );
  IV U1286 ( .A(a[572]), .Z(n2717) );
  IV U1287 ( .A(b[572]), .Z(n429) );
  NOR U1288 ( .A(n2717), .B(n429), .Z(n2719) );
  IV U1289 ( .A(a[571]), .Z(n2714) );
  IV U1290 ( .A(b[571]), .Z(n430) );
  NOR U1291 ( .A(n2714), .B(n430), .Z(n2716) );
  IV U1292 ( .A(a[570]), .Z(n2711) );
  IV U1293 ( .A(b[570]), .Z(n431) );
  NOR U1294 ( .A(n2711), .B(n431), .Z(n2713) );
  IV U1295 ( .A(a[569]), .Z(n2708) );
  IV U1296 ( .A(b[569]), .Z(n432) );
  NOR U1297 ( .A(n2708), .B(n432), .Z(n2710) );
  IV U1298 ( .A(a[568]), .Z(n2705) );
  IV U1299 ( .A(b[568]), .Z(n433) );
  NOR U1300 ( .A(n2705), .B(n433), .Z(n2707) );
  IV U1301 ( .A(a[567]), .Z(n2702) );
  IV U1302 ( .A(b[567]), .Z(n434) );
  NOR U1303 ( .A(n2702), .B(n434), .Z(n2704) );
  IV U1304 ( .A(a[566]), .Z(n2699) );
  IV U1305 ( .A(b[566]), .Z(n435) );
  NOR U1306 ( .A(n2699), .B(n435), .Z(n2701) );
  IV U1307 ( .A(a[565]), .Z(n2696) );
  IV U1308 ( .A(b[565]), .Z(n436) );
  NOR U1309 ( .A(n2696), .B(n436), .Z(n2698) );
  IV U1310 ( .A(a[564]), .Z(n2693) );
  IV U1311 ( .A(b[564]), .Z(n437) );
  NOR U1312 ( .A(n2693), .B(n437), .Z(n2695) );
  IV U1313 ( .A(a[563]), .Z(n2690) );
  IV U1314 ( .A(b[563]), .Z(n438) );
  NOR U1315 ( .A(n2690), .B(n438), .Z(n2692) );
  IV U1316 ( .A(a[562]), .Z(n2687) );
  IV U1317 ( .A(b[562]), .Z(n439) );
  NOR U1318 ( .A(n2687), .B(n439), .Z(n2689) );
  IV U1319 ( .A(a[561]), .Z(n2684) );
  IV U1320 ( .A(b[561]), .Z(n440) );
  NOR U1321 ( .A(n2684), .B(n440), .Z(n2686) );
  IV U1322 ( .A(a[560]), .Z(n2681) );
  IV U1323 ( .A(b[560]), .Z(n441) );
  NOR U1324 ( .A(n2681), .B(n441), .Z(n2683) );
  IV U1325 ( .A(a[559]), .Z(n2678) );
  IV U1326 ( .A(b[559]), .Z(n442) );
  NOR U1327 ( .A(n2678), .B(n442), .Z(n2680) );
  IV U1328 ( .A(a[558]), .Z(n2675) );
  IV U1329 ( .A(b[558]), .Z(n443) );
  NOR U1330 ( .A(n2675), .B(n443), .Z(n2677) );
  IV U1331 ( .A(a[557]), .Z(n2672) );
  IV U1332 ( .A(b[557]), .Z(n444) );
  NOR U1333 ( .A(n2672), .B(n444), .Z(n2674) );
  IV U1334 ( .A(a[556]), .Z(n2669) );
  IV U1335 ( .A(b[556]), .Z(n445) );
  NOR U1336 ( .A(n2669), .B(n445), .Z(n2671) );
  IV U1337 ( .A(a[555]), .Z(n2666) );
  IV U1338 ( .A(b[555]), .Z(n446) );
  NOR U1339 ( .A(n2666), .B(n446), .Z(n2668) );
  IV U1340 ( .A(a[554]), .Z(n2663) );
  IV U1341 ( .A(b[554]), .Z(n447) );
  NOR U1342 ( .A(n2663), .B(n447), .Z(n2665) );
  IV U1343 ( .A(a[553]), .Z(n2660) );
  IV U1344 ( .A(b[553]), .Z(n448) );
  NOR U1345 ( .A(n2660), .B(n448), .Z(n2662) );
  IV U1346 ( .A(a[552]), .Z(n2657) );
  IV U1347 ( .A(b[552]), .Z(n449) );
  NOR U1348 ( .A(n2657), .B(n449), .Z(n2659) );
  IV U1349 ( .A(a[551]), .Z(n2654) );
  IV U1350 ( .A(b[551]), .Z(n450) );
  NOR U1351 ( .A(n2654), .B(n450), .Z(n2656) );
  IV U1352 ( .A(a[550]), .Z(n2651) );
  IV U1353 ( .A(b[550]), .Z(n451) );
  NOR U1354 ( .A(n2651), .B(n451), .Z(n2653) );
  IV U1355 ( .A(a[549]), .Z(n2648) );
  IV U1356 ( .A(b[549]), .Z(n452) );
  NOR U1357 ( .A(n2648), .B(n452), .Z(n2650) );
  IV U1358 ( .A(a[548]), .Z(n2645) );
  IV U1359 ( .A(b[548]), .Z(n453) );
  NOR U1360 ( .A(n2645), .B(n453), .Z(n2647) );
  IV U1361 ( .A(a[547]), .Z(n2642) );
  IV U1362 ( .A(b[547]), .Z(n454) );
  NOR U1363 ( .A(n2642), .B(n454), .Z(n2644) );
  IV U1364 ( .A(a[546]), .Z(n2639) );
  IV U1365 ( .A(b[546]), .Z(n455) );
  NOR U1366 ( .A(n2639), .B(n455), .Z(n2641) );
  IV U1367 ( .A(a[545]), .Z(n2636) );
  IV U1368 ( .A(b[545]), .Z(n456) );
  NOR U1369 ( .A(n2636), .B(n456), .Z(n2638) );
  IV U1370 ( .A(a[544]), .Z(n2633) );
  IV U1371 ( .A(b[544]), .Z(n457) );
  NOR U1372 ( .A(n2633), .B(n457), .Z(n2635) );
  IV U1373 ( .A(a[543]), .Z(n2630) );
  IV U1374 ( .A(b[543]), .Z(n458) );
  NOR U1375 ( .A(n2630), .B(n458), .Z(n2632) );
  IV U1376 ( .A(a[542]), .Z(n2627) );
  IV U1377 ( .A(b[542]), .Z(n459) );
  NOR U1378 ( .A(n2627), .B(n459), .Z(n2629) );
  IV U1379 ( .A(a[541]), .Z(n2624) );
  IV U1380 ( .A(b[541]), .Z(n460) );
  NOR U1381 ( .A(n2624), .B(n460), .Z(n2626) );
  IV U1382 ( .A(a[540]), .Z(n2621) );
  IV U1383 ( .A(b[540]), .Z(n461) );
  NOR U1384 ( .A(n2621), .B(n461), .Z(n2623) );
  IV U1385 ( .A(a[539]), .Z(n2618) );
  IV U1386 ( .A(b[539]), .Z(n462) );
  NOR U1387 ( .A(n2618), .B(n462), .Z(n2620) );
  IV U1388 ( .A(a[538]), .Z(n2615) );
  IV U1389 ( .A(b[538]), .Z(n463) );
  NOR U1390 ( .A(n2615), .B(n463), .Z(n2617) );
  IV U1391 ( .A(a[537]), .Z(n2612) );
  IV U1392 ( .A(b[537]), .Z(n464) );
  NOR U1393 ( .A(n2612), .B(n464), .Z(n2614) );
  IV U1394 ( .A(a[536]), .Z(n2609) );
  IV U1395 ( .A(b[536]), .Z(n465) );
  NOR U1396 ( .A(n2609), .B(n465), .Z(n2611) );
  IV U1397 ( .A(a[535]), .Z(n2606) );
  IV U1398 ( .A(b[535]), .Z(n466) );
  NOR U1399 ( .A(n2606), .B(n466), .Z(n2608) );
  IV U1400 ( .A(a[534]), .Z(n2603) );
  IV U1401 ( .A(b[534]), .Z(n467) );
  NOR U1402 ( .A(n2603), .B(n467), .Z(n2605) );
  IV U1403 ( .A(a[533]), .Z(n2600) );
  IV U1404 ( .A(b[533]), .Z(n468) );
  NOR U1405 ( .A(n2600), .B(n468), .Z(n2602) );
  IV U1406 ( .A(a[532]), .Z(n2597) );
  IV U1407 ( .A(b[532]), .Z(n469) );
  NOR U1408 ( .A(n2597), .B(n469), .Z(n2599) );
  IV U1409 ( .A(a[531]), .Z(n2594) );
  IV U1410 ( .A(b[531]), .Z(n470) );
  NOR U1411 ( .A(n2594), .B(n470), .Z(n2596) );
  IV U1412 ( .A(a[530]), .Z(n2591) );
  IV U1413 ( .A(b[530]), .Z(n471) );
  NOR U1414 ( .A(n2591), .B(n471), .Z(n2593) );
  IV U1415 ( .A(a[529]), .Z(n2588) );
  IV U1416 ( .A(b[529]), .Z(n472) );
  NOR U1417 ( .A(n2588), .B(n472), .Z(n2590) );
  IV U1418 ( .A(a[528]), .Z(n2585) );
  IV U1419 ( .A(b[528]), .Z(n473) );
  NOR U1420 ( .A(n2585), .B(n473), .Z(n2587) );
  IV U1421 ( .A(a[527]), .Z(n2582) );
  IV U1422 ( .A(b[527]), .Z(n474) );
  NOR U1423 ( .A(n2582), .B(n474), .Z(n2584) );
  IV U1424 ( .A(a[526]), .Z(n2579) );
  IV U1425 ( .A(b[526]), .Z(n475) );
  NOR U1426 ( .A(n2579), .B(n475), .Z(n2581) );
  IV U1427 ( .A(a[525]), .Z(n2576) );
  IV U1428 ( .A(b[525]), .Z(n476) );
  NOR U1429 ( .A(n2576), .B(n476), .Z(n2578) );
  IV U1430 ( .A(a[524]), .Z(n2573) );
  IV U1431 ( .A(b[524]), .Z(n477) );
  NOR U1432 ( .A(n2573), .B(n477), .Z(n2575) );
  IV U1433 ( .A(a[523]), .Z(n2570) );
  IV U1434 ( .A(b[523]), .Z(n478) );
  NOR U1435 ( .A(n2570), .B(n478), .Z(n2572) );
  IV U1436 ( .A(a[522]), .Z(n2567) );
  IV U1437 ( .A(b[522]), .Z(n479) );
  NOR U1438 ( .A(n2567), .B(n479), .Z(n2569) );
  IV U1439 ( .A(a[521]), .Z(n2564) );
  IV U1440 ( .A(b[521]), .Z(n480) );
  NOR U1441 ( .A(n2564), .B(n480), .Z(n2566) );
  IV U1442 ( .A(a[520]), .Z(n2561) );
  IV U1443 ( .A(b[520]), .Z(n481) );
  NOR U1444 ( .A(n2561), .B(n481), .Z(n2563) );
  IV U1445 ( .A(a[519]), .Z(n2558) );
  IV U1446 ( .A(b[519]), .Z(n482) );
  NOR U1447 ( .A(n2558), .B(n482), .Z(n2560) );
  IV U1448 ( .A(a[518]), .Z(n2555) );
  IV U1449 ( .A(b[518]), .Z(n483) );
  NOR U1450 ( .A(n2555), .B(n483), .Z(n2557) );
  IV U1451 ( .A(a[517]), .Z(n2552) );
  IV U1452 ( .A(b[517]), .Z(n484) );
  NOR U1453 ( .A(n2552), .B(n484), .Z(n2554) );
  IV U1454 ( .A(a[516]), .Z(n2549) );
  IV U1455 ( .A(b[516]), .Z(n485) );
  NOR U1456 ( .A(n2549), .B(n485), .Z(n2551) );
  IV U1457 ( .A(a[515]), .Z(n2546) );
  IV U1458 ( .A(b[515]), .Z(n486) );
  NOR U1459 ( .A(n2546), .B(n486), .Z(n2548) );
  IV U1460 ( .A(a[514]), .Z(n2543) );
  IV U1461 ( .A(b[514]), .Z(n487) );
  NOR U1462 ( .A(n2543), .B(n487), .Z(n2545) );
  IV U1463 ( .A(a[513]), .Z(n2540) );
  IV U1464 ( .A(b[513]), .Z(n488) );
  NOR U1465 ( .A(n2540), .B(n488), .Z(n2542) );
  IV U1466 ( .A(a[512]), .Z(n2537) );
  IV U1467 ( .A(b[512]), .Z(n489) );
  NOR U1468 ( .A(n2537), .B(n489), .Z(n2539) );
  IV U1469 ( .A(a[511]), .Z(n2534) );
  IV U1470 ( .A(b[511]), .Z(n490) );
  NOR U1471 ( .A(n2534), .B(n490), .Z(n2536) );
  IV U1472 ( .A(a[510]), .Z(n2531) );
  IV U1473 ( .A(b[510]), .Z(n491) );
  NOR U1474 ( .A(n2531), .B(n491), .Z(n2533) );
  IV U1475 ( .A(a[509]), .Z(n2528) );
  IV U1476 ( .A(b[509]), .Z(n492) );
  NOR U1477 ( .A(n2528), .B(n492), .Z(n2530) );
  IV U1478 ( .A(a[508]), .Z(n2525) );
  IV U1479 ( .A(b[508]), .Z(n493) );
  NOR U1480 ( .A(n2525), .B(n493), .Z(n2527) );
  IV U1481 ( .A(a[507]), .Z(n2522) );
  IV U1482 ( .A(b[507]), .Z(n494) );
  NOR U1483 ( .A(n2522), .B(n494), .Z(n2524) );
  IV U1484 ( .A(a[506]), .Z(n2519) );
  IV U1485 ( .A(b[506]), .Z(n495) );
  NOR U1486 ( .A(n2519), .B(n495), .Z(n2521) );
  IV U1487 ( .A(a[505]), .Z(n2516) );
  IV U1488 ( .A(b[505]), .Z(n496) );
  NOR U1489 ( .A(n2516), .B(n496), .Z(n2518) );
  IV U1490 ( .A(a[504]), .Z(n2513) );
  IV U1491 ( .A(b[504]), .Z(n497) );
  NOR U1492 ( .A(n2513), .B(n497), .Z(n2515) );
  IV U1493 ( .A(a[503]), .Z(n2510) );
  IV U1494 ( .A(b[503]), .Z(n498) );
  NOR U1495 ( .A(n2510), .B(n498), .Z(n2512) );
  IV U1496 ( .A(a[502]), .Z(n2507) );
  IV U1497 ( .A(b[502]), .Z(n499) );
  NOR U1498 ( .A(n2507), .B(n499), .Z(n2509) );
  IV U1499 ( .A(a[501]), .Z(n2504) );
  IV U1500 ( .A(b[501]), .Z(n500) );
  NOR U1501 ( .A(n2504), .B(n500), .Z(n2506) );
  IV U1502 ( .A(a[500]), .Z(n2501) );
  IV U1503 ( .A(b[500]), .Z(n501) );
  NOR U1504 ( .A(n2501), .B(n501), .Z(n2503) );
  IV U1505 ( .A(a[499]), .Z(n2498) );
  IV U1506 ( .A(b[499]), .Z(n502) );
  NOR U1507 ( .A(n2498), .B(n502), .Z(n2500) );
  IV U1508 ( .A(a[498]), .Z(n2495) );
  IV U1509 ( .A(b[498]), .Z(n503) );
  NOR U1510 ( .A(n2495), .B(n503), .Z(n2497) );
  IV U1511 ( .A(a[497]), .Z(n2492) );
  IV U1512 ( .A(b[497]), .Z(n504) );
  NOR U1513 ( .A(n2492), .B(n504), .Z(n2494) );
  IV U1514 ( .A(a[496]), .Z(n2489) );
  IV U1515 ( .A(b[496]), .Z(n505) );
  NOR U1516 ( .A(n2489), .B(n505), .Z(n2491) );
  IV U1517 ( .A(a[495]), .Z(n2486) );
  IV U1518 ( .A(b[495]), .Z(n506) );
  NOR U1519 ( .A(n2486), .B(n506), .Z(n2488) );
  IV U1520 ( .A(a[494]), .Z(n2483) );
  IV U1521 ( .A(b[494]), .Z(n507) );
  NOR U1522 ( .A(n2483), .B(n507), .Z(n2485) );
  IV U1523 ( .A(a[493]), .Z(n2480) );
  IV U1524 ( .A(b[493]), .Z(n508) );
  NOR U1525 ( .A(n2480), .B(n508), .Z(n2482) );
  IV U1526 ( .A(a[492]), .Z(n2477) );
  IV U1527 ( .A(b[492]), .Z(n509) );
  NOR U1528 ( .A(n2477), .B(n509), .Z(n2479) );
  IV U1529 ( .A(a[491]), .Z(n2474) );
  IV U1530 ( .A(b[491]), .Z(n510) );
  NOR U1531 ( .A(n2474), .B(n510), .Z(n2476) );
  IV U1532 ( .A(a[490]), .Z(n2471) );
  IV U1533 ( .A(b[490]), .Z(n511) );
  NOR U1534 ( .A(n2471), .B(n511), .Z(n2473) );
  IV U1535 ( .A(a[489]), .Z(n2468) );
  IV U1536 ( .A(b[489]), .Z(n512) );
  NOR U1537 ( .A(n2468), .B(n512), .Z(n2470) );
  IV U1538 ( .A(a[488]), .Z(n2465) );
  IV U1539 ( .A(b[488]), .Z(n513) );
  NOR U1540 ( .A(n2465), .B(n513), .Z(n2467) );
  IV U1541 ( .A(a[487]), .Z(n2462) );
  IV U1542 ( .A(b[487]), .Z(n514) );
  NOR U1543 ( .A(n2462), .B(n514), .Z(n2464) );
  IV U1544 ( .A(a[486]), .Z(n2459) );
  IV U1545 ( .A(b[486]), .Z(n515) );
  NOR U1546 ( .A(n2459), .B(n515), .Z(n2461) );
  IV U1547 ( .A(a[485]), .Z(n2456) );
  IV U1548 ( .A(b[485]), .Z(n516) );
  NOR U1549 ( .A(n2456), .B(n516), .Z(n2458) );
  IV U1550 ( .A(a[484]), .Z(n2453) );
  IV U1551 ( .A(b[484]), .Z(n517) );
  NOR U1552 ( .A(n2453), .B(n517), .Z(n2455) );
  IV U1553 ( .A(a[483]), .Z(n2450) );
  IV U1554 ( .A(b[483]), .Z(n518) );
  NOR U1555 ( .A(n2450), .B(n518), .Z(n2452) );
  IV U1556 ( .A(a[482]), .Z(n2447) );
  IV U1557 ( .A(b[482]), .Z(n519) );
  NOR U1558 ( .A(n2447), .B(n519), .Z(n2449) );
  IV U1559 ( .A(a[481]), .Z(n2444) );
  IV U1560 ( .A(b[481]), .Z(n520) );
  NOR U1561 ( .A(n2444), .B(n520), .Z(n2446) );
  IV U1562 ( .A(a[480]), .Z(n2441) );
  IV U1563 ( .A(b[480]), .Z(n521) );
  NOR U1564 ( .A(n2441), .B(n521), .Z(n2443) );
  IV U1565 ( .A(a[479]), .Z(n2438) );
  IV U1566 ( .A(b[479]), .Z(n522) );
  NOR U1567 ( .A(n2438), .B(n522), .Z(n2440) );
  IV U1568 ( .A(a[478]), .Z(n2435) );
  IV U1569 ( .A(b[478]), .Z(n523) );
  NOR U1570 ( .A(n2435), .B(n523), .Z(n2437) );
  IV U1571 ( .A(a[477]), .Z(n2432) );
  IV U1572 ( .A(b[477]), .Z(n524) );
  NOR U1573 ( .A(n2432), .B(n524), .Z(n2434) );
  IV U1574 ( .A(a[476]), .Z(n2429) );
  IV U1575 ( .A(b[476]), .Z(n525) );
  NOR U1576 ( .A(n2429), .B(n525), .Z(n2431) );
  IV U1577 ( .A(a[475]), .Z(n2426) );
  IV U1578 ( .A(b[475]), .Z(n526) );
  NOR U1579 ( .A(n2426), .B(n526), .Z(n2428) );
  IV U1580 ( .A(a[474]), .Z(n2423) );
  IV U1581 ( .A(b[474]), .Z(n527) );
  NOR U1582 ( .A(n2423), .B(n527), .Z(n2425) );
  IV U1583 ( .A(a[473]), .Z(n2420) );
  IV U1584 ( .A(b[473]), .Z(n528) );
  NOR U1585 ( .A(n2420), .B(n528), .Z(n2422) );
  IV U1586 ( .A(a[472]), .Z(n2417) );
  IV U1587 ( .A(b[472]), .Z(n529) );
  NOR U1588 ( .A(n2417), .B(n529), .Z(n2419) );
  IV U1589 ( .A(a[471]), .Z(n2414) );
  IV U1590 ( .A(b[471]), .Z(n530) );
  NOR U1591 ( .A(n2414), .B(n530), .Z(n2416) );
  IV U1592 ( .A(a[470]), .Z(n2411) );
  IV U1593 ( .A(b[470]), .Z(n531) );
  NOR U1594 ( .A(n2411), .B(n531), .Z(n2413) );
  IV U1595 ( .A(a[469]), .Z(n2408) );
  IV U1596 ( .A(b[469]), .Z(n532) );
  NOR U1597 ( .A(n2408), .B(n532), .Z(n2410) );
  IV U1598 ( .A(a[468]), .Z(n2405) );
  IV U1599 ( .A(b[468]), .Z(n533) );
  NOR U1600 ( .A(n2405), .B(n533), .Z(n2407) );
  IV U1601 ( .A(a[467]), .Z(n2402) );
  IV U1602 ( .A(b[467]), .Z(n534) );
  NOR U1603 ( .A(n2402), .B(n534), .Z(n2404) );
  IV U1604 ( .A(a[466]), .Z(n2399) );
  IV U1605 ( .A(b[466]), .Z(n535) );
  NOR U1606 ( .A(n2399), .B(n535), .Z(n2401) );
  IV U1607 ( .A(a[465]), .Z(n2396) );
  IV U1608 ( .A(b[465]), .Z(n536) );
  NOR U1609 ( .A(n2396), .B(n536), .Z(n2398) );
  IV U1610 ( .A(a[464]), .Z(n2393) );
  IV U1611 ( .A(b[464]), .Z(n537) );
  NOR U1612 ( .A(n2393), .B(n537), .Z(n2395) );
  IV U1613 ( .A(a[463]), .Z(n2390) );
  IV U1614 ( .A(b[463]), .Z(n538) );
  NOR U1615 ( .A(n2390), .B(n538), .Z(n2392) );
  IV U1616 ( .A(a[462]), .Z(n2387) );
  IV U1617 ( .A(b[462]), .Z(n539) );
  NOR U1618 ( .A(n2387), .B(n539), .Z(n2389) );
  IV U1619 ( .A(a[461]), .Z(n2384) );
  IV U1620 ( .A(b[461]), .Z(n540) );
  NOR U1621 ( .A(n2384), .B(n540), .Z(n2386) );
  IV U1622 ( .A(a[460]), .Z(n2381) );
  IV U1623 ( .A(b[460]), .Z(n541) );
  NOR U1624 ( .A(n2381), .B(n541), .Z(n2383) );
  IV U1625 ( .A(a[459]), .Z(n2378) );
  IV U1626 ( .A(b[459]), .Z(n542) );
  NOR U1627 ( .A(n2378), .B(n542), .Z(n2380) );
  IV U1628 ( .A(a[458]), .Z(n2375) );
  IV U1629 ( .A(b[458]), .Z(n543) );
  NOR U1630 ( .A(n2375), .B(n543), .Z(n2377) );
  IV U1631 ( .A(a[457]), .Z(n2372) );
  IV U1632 ( .A(b[457]), .Z(n544) );
  NOR U1633 ( .A(n2372), .B(n544), .Z(n2374) );
  IV U1634 ( .A(a[456]), .Z(n2369) );
  IV U1635 ( .A(b[456]), .Z(n545) );
  NOR U1636 ( .A(n2369), .B(n545), .Z(n2371) );
  IV U1637 ( .A(a[455]), .Z(n2366) );
  IV U1638 ( .A(b[455]), .Z(n546) );
  NOR U1639 ( .A(n2366), .B(n546), .Z(n2368) );
  IV U1640 ( .A(a[454]), .Z(n2363) );
  IV U1641 ( .A(b[454]), .Z(n547) );
  NOR U1642 ( .A(n2363), .B(n547), .Z(n2365) );
  IV U1643 ( .A(a[453]), .Z(n2360) );
  IV U1644 ( .A(b[453]), .Z(n548) );
  NOR U1645 ( .A(n2360), .B(n548), .Z(n2362) );
  IV U1646 ( .A(a[452]), .Z(n2357) );
  IV U1647 ( .A(b[452]), .Z(n549) );
  NOR U1648 ( .A(n2357), .B(n549), .Z(n2359) );
  IV U1649 ( .A(a[451]), .Z(n2354) );
  IV U1650 ( .A(b[451]), .Z(n550) );
  NOR U1651 ( .A(n2354), .B(n550), .Z(n2356) );
  IV U1652 ( .A(a[450]), .Z(n2351) );
  IV U1653 ( .A(b[450]), .Z(n551) );
  NOR U1654 ( .A(n2351), .B(n551), .Z(n2353) );
  IV U1655 ( .A(a[449]), .Z(n2348) );
  IV U1656 ( .A(b[449]), .Z(n552) );
  NOR U1657 ( .A(n2348), .B(n552), .Z(n2350) );
  IV U1658 ( .A(a[448]), .Z(n2345) );
  IV U1659 ( .A(b[448]), .Z(n553) );
  NOR U1660 ( .A(n2345), .B(n553), .Z(n2347) );
  IV U1661 ( .A(a[447]), .Z(n2342) );
  IV U1662 ( .A(b[447]), .Z(n554) );
  NOR U1663 ( .A(n2342), .B(n554), .Z(n2344) );
  IV U1664 ( .A(a[446]), .Z(n2339) );
  IV U1665 ( .A(b[446]), .Z(n555) );
  NOR U1666 ( .A(n2339), .B(n555), .Z(n2341) );
  IV U1667 ( .A(a[445]), .Z(n2336) );
  IV U1668 ( .A(b[445]), .Z(n556) );
  NOR U1669 ( .A(n2336), .B(n556), .Z(n2338) );
  IV U1670 ( .A(a[444]), .Z(n2333) );
  IV U1671 ( .A(b[444]), .Z(n557) );
  NOR U1672 ( .A(n2333), .B(n557), .Z(n2335) );
  IV U1673 ( .A(a[443]), .Z(n2330) );
  IV U1674 ( .A(b[443]), .Z(n558) );
  NOR U1675 ( .A(n2330), .B(n558), .Z(n2332) );
  IV U1676 ( .A(a[442]), .Z(n2327) );
  IV U1677 ( .A(b[442]), .Z(n559) );
  NOR U1678 ( .A(n2327), .B(n559), .Z(n2329) );
  IV U1679 ( .A(a[441]), .Z(n2324) );
  IV U1680 ( .A(b[441]), .Z(n560) );
  NOR U1681 ( .A(n2324), .B(n560), .Z(n2326) );
  IV U1682 ( .A(a[440]), .Z(n2321) );
  IV U1683 ( .A(b[440]), .Z(n561) );
  NOR U1684 ( .A(n2321), .B(n561), .Z(n2323) );
  IV U1685 ( .A(a[439]), .Z(n2318) );
  IV U1686 ( .A(b[439]), .Z(n562) );
  NOR U1687 ( .A(n2318), .B(n562), .Z(n2320) );
  IV U1688 ( .A(a[438]), .Z(n2315) );
  IV U1689 ( .A(b[438]), .Z(n563) );
  NOR U1690 ( .A(n2315), .B(n563), .Z(n2317) );
  IV U1691 ( .A(a[437]), .Z(n2312) );
  IV U1692 ( .A(b[437]), .Z(n564) );
  NOR U1693 ( .A(n2312), .B(n564), .Z(n2314) );
  IV U1694 ( .A(a[436]), .Z(n2309) );
  IV U1695 ( .A(b[436]), .Z(n565) );
  NOR U1696 ( .A(n2309), .B(n565), .Z(n2311) );
  IV U1697 ( .A(a[435]), .Z(n2306) );
  IV U1698 ( .A(b[435]), .Z(n566) );
  NOR U1699 ( .A(n2306), .B(n566), .Z(n2308) );
  IV U1700 ( .A(a[434]), .Z(n2303) );
  IV U1701 ( .A(b[434]), .Z(n567) );
  NOR U1702 ( .A(n2303), .B(n567), .Z(n2305) );
  IV U1703 ( .A(a[433]), .Z(n2300) );
  IV U1704 ( .A(b[433]), .Z(n568) );
  NOR U1705 ( .A(n2300), .B(n568), .Z(n2302) );
  IV U1706 ( .A(a[432]), .Z(n2297) );
  IV U1707 ( .A(b[432]), .Z(n569) );
  NOR U1708 ( .A(n2297), .B(n569), .Z(n2299) );
  IV U1709 ( .A(a[431]), .Z(n2294) );
  IV U1710 ( .A(b[431]), .Z(n570) );
  NOR U1711 ( .A(n2294), .B(n570), .Z(n2296) );
  IV U1712 ( .A(a[430]), .Z(n2291) );
  IV U1713 ( .A(b[430]), .Z(n571) );
  NOR U1714 ( .A(n2291), .B(n571), .Z(n2293) );
  IV U1715 ( .A(a[429]), .Z(n2288) );
  IV U1716 ( .A(b[429]), .Z(n572) );
  NOR U1717 ( .A(n2288), .B(n572), .Z(n2290) );
  IV U1718 ( .A(a[428]), .Z(n2285) );
  IV U1719 ( .A(b[428]), .Z(n573) );
  NOR U1720 ( .A(n2285), .B(n573), .Z(n2287) );
  IV U1721 ( .A(a[427]), .Z(n2282) );
  IV U1722 ( .A(b[427]), .Z(n574) );
  NOR U1723 ( .A(n2282), .B(n574), .Z(n2284) );
  IV U1724 ( .A(a[426]), .Z(n2279) );
  IV U1725 ( .A(b[426]), .Z(n575) );
  NOR U1726 ( .A(n2279), .B(n575), .Z(n2281) );
  IV U1727 ( .A(a[425]), .Z(n2276) );
  IV U1728 ( .A(b[425]), .Z(n576) );
  NOR U1729 ( .A(n2276), .B(n576), .Z(n2278) );
  IV U1730 ( .A(a[424]), .Z(n2273) );
  IV U1731 ( .A(b[424]), .Z(n577) );
  NOR U1732 ( .A(n2273), .B(n577), .Z(n2275) );
  IV U1733 ( .A(a[423]), .Z(n2270) );
  IV U1734 ( .A(b[423]), .Z(n578) );
  NOR U1735 ( .A(n2270), .B(n578), .Z(n2272) );
  IV U1736 ( .A(a[422]), .Z(n2267) );
  IV U1737 ( .A(b[422]), .Z(n579) );
  NOR U1738 ( .A(n2267), .B(n579), .Z(n2269) );
  IV U1739 ( .A(a[421]), .Z(n2264) );
  IV U1740 ( .A(b[421]), .Z(n580) );
  NOR U1741 ( .A(n2264), .B(n580), .Z(n2266) );
  IV U1742 ( .A(a[420]), .Z(n2261) );
  IV U1743 ( .A(b[420]), .Z(n581) );
  NOR U1744 ( .A(n2261), .B(n581), .Z(n2263) );
  IV U1745 ( .A(a[419]), .Z(n2258) );
  IV U1746 ( .A(b[419]), .Z(n582) );
  NOR U1747 ( .A(n2258), .B(n582), .Z(n2260) );
  IV U1748 ( .A(a[418]), .Z(n2255) );
  IV U1749 ( .A(b[418]), .Z(n583) );
  NOR U1750 ( .A(n2255), .B(n583), .Z(n2257) );
  IV U1751 ( .A(a[417]), .Z(n2252) );
  IV U1752 ( .A(b[417]), .Z(n584) );
  NOR U1753 ( .A(n2252), .B(n584), .Z(n2254) );
  IV U1754 ( .A(a[416]), .Z(n2249) );
  IV U1755 ( .A(b[416]), .Z(n585) );
  NOR U1756 ( .A(n2249), .B(n585), .Z(n2251) );
  IV U1757 ( .A(a[415]), .Z(n2246) );
  IV U1758 ( .A(b[415]), .Z(n586) );
  NOR U1759 ( .A(n2246), .B(n586), .Z(n2248) );
  IV U1760 ( .A(a[414]), .Z(n2243) );
  IV U1761 ( .A(b[414]), .Z(n587) );
  NOR U1762 ( .A(n2243), .B(n587), .Z(n2245) );
  IV U1763 ( .A(a[413]), .Z(n2240) );
  IV U1764 ( .A(b[413]), .Z(n588) );
  NOR U1765 ( .A(n2240), .B(n588), .Z(n2242) );
  IV U1766 ( .A(a[412]), .Z(n2237) );
  IV U1767 ( .A(b[412]), .Z(n589) );
  NOR U1768 ( .A(n2237), .B(n589), .Z(n2239) );
  IV U1769 ( .A(a[411]), .Z(n2234) );
  IV U1770 ( .A(b[411]), .Z(n590) );
  NOR U1771 ( .A(n2234), .B(n590), .Z(n2236) );
  IV U1772 ( .A(a[410]), .Z(n2231) );
  IV U1773 ( .A(b[410]), .Z(n591) );
  NOR U1774 ( .A(n2231), .B(n591), .Z(n2233) );
  IV U1775 ( .A(a[409]), .Z(n2228) );
  IV U1776 ( .A(b[409]), .Z(n592) );
  NOR U1777 ( .A(n2228), .B(n592), .Z(n2230) );
  IV U1778 ( .A(a[408]), .Z(n2225) );
  IV U1779 ( .A(b[408]), .Z(n593) );
  NOR U1780 ( .A(n2225), .B(n593), .Z(n2227) );
  IV U1781 ( .A(a[407]), .Z(n2222) );
  IV U1782 ( .A(b[407]), .Z(n594) );
  NOR U1783 ( .A(n2222), .B(n594), .Z(n2224) );
  IV U1784 ( .A(a[406]), .Z(n2219) );
  IV U1785 ( .A(b[406]), .Z(n595) );
  NOR U1786 ( .A(n2219), .B(n595), .Z(n2221) );
  IV U1787 ( .A(a[405]), .Z(n2216) );
  IV U1788 ( .A(b[405]), .Z(n596) );
  NOR U1789 ( .A(n2216), .B(n596), .Z(n2218) );
  IV U1790 ( .A(a[404]), .Z(n2213) );
  IV U1791 ( .A(b[404]), .Z(n597) );
  NOR U1792 ( .A(n2213), .B(n597), .Z(n2215) );
  IV U1793 ( .A(a[403]), .Z(n2210) );
  IV U1794 ( .A(b[403]), .Z(n598) );
  NOR U1795 ( .A(n2210), .B(n598), .Z(n2212) );
  IV U1796 ( .A(a[402]), .Z(n2207) );
  IV U1797 ( .A(b[402]), .Z(n599) );
  NOR U1798 ( .A(n2207), .B(n599), .Z(n2209) );
  IV U1799 ( .A(a[401]), .Z(n2204) );
  IV U1800 ( .A(b[401]), .Z(n600) );
  NOR U1801 ( .A(n2204), .B(n600), .Z(n2206) );
  IV U1802 ( .A(a[400]), .Z(n2201) );
  IV U1803 ( .A(b[400]), .Z(n601) );
  NOR U1804 ( .A(n2201), .B(n601), .Z(n2203) );
  IV U1805 ( .A(a[399]), .Z(n2198) );
  IV U1806 ( .A(b[399]), .Z(n602) );
  NOR U1807 ( .A(n2198), .B(n602), .Z(n2200) );
  IV U1808 ( .A(a[398]), .Z(n2195) );
  IV U1809 ( .A(b[398]), .Z(n603) );
  NOR U1810 ( .A(n2195), .B(n603), .Z(n2197) );
  IV U1811 ( .A(a[397]), .Z(n2192) );
  IV U1812 ( .A(b[397]), .Z(n604) );
  NOR U1813 ( .A(n2192), .B(n604), .Z(n2194) );
  IV U1814 ( .A(a[396]), .Z(n2189) );
  IV U1815 ( .A(b[396]), .Z(n605) );
  NOR U1816 ( .A(n2189), .B(n605), .Z(n2191) );
  IV U1817 ( .A(a[395]), .Z(n2186) );
  IV U1818 ( .A(b[395]), .Z(n606) );
  NOR U1819 ( .A(n2186), .B(n606), .Z(n2188) );
  IV U1820 ( .A(a[394]), .Z(n2183) );
  IV U1821 ( .A(b[394]), .Z(n607) );
  NOR U1822 ( .A(n2183), .B(n607), .Z(n2185) );
  IV U1823 ( .A(a[393]), .Z(n2180) );
  IV U1824 ( .A(b[393]), .Z(n608) );
  NOR U1825 ( .A(n2180), .B(n608), .Z(n2182) );
  IV U1826 ( .A(a[392]), .Z(n2177) );
  IV U1827 ( .A(b[392]), .Z(n609) );
  NOR U1828 ( .A(n2177), .B(n609), .Z(n2179) );
  IV U1829 ( .A(a[391]), .Z(n2174) );
  IV U1830 ( .A(b[391]), .Z(n610) );
  NOR U1831 ( .A(n2174), .B(n610), .Z(n2176) );
  IV U1832 ( .A(a[390]), .Z(n2171) );
  IV U1833 ( .A(b[390]), .Z(n611) );
  NOR U1834 ( .A(n2171), .B(n611), .Z(n2173) );
  IV U1835 ( .A(a[389]), .Z(n2168) );
  IV U1836 ( .A(b[389]), .Z(n612) );
  NOR U1837 ( .A(n2168), .B(n612), .Z(n2170) );
  IV U1838 ( .A(a[388]), .Z(n2165) );
  IV U1839 ( .A(b[388]), .Z(n613) );
  NOR U1840 ( .A(n2165), .B(n613), .Z(n2167) );
  IV U1841 ( .A(a[387]), .Z(n2162) );
  IV U1842 ( .A(b[387]), .Z(n614) );
  NOR U1843 ( .A(n2162), .B(n614), .Z(n2164) );
  IV U1844 ( .A(a[386]), .Z(n2159) );
  IV U1845 ( .A(b[386]), .Z(n615) );
  NOR U1846 ( .A(n2159), .B(n615), .Z(n2161) );
  IV U1847 ( .A(a[385]), .Z(n2156) );
  IV U1848 ( .A(b[385]), .Z(n616) );
  NOR U1849 ( .A(n2156), .B(n616), .Z(n2158) );
  IV U1850 ( .A(a[384]), .Z(n2153) );
  IV U1851 ( .A(b[384]), .Z(n617) );
  NOR U1852 ( .A(n2153), .B(n617), .Z(n2155) );
  IV U1853 ( .A(a[383]), .Z(n2150) );
  IV U1854 ( .A(b[383]), .Z(n618) );
  NOR U1855 ( .A(n2150), .B(n618), .Z(n2152) );
  IV U1856 ( .A(a[382]), .Z(n2147) );
  IV U1857 ( .A(b[382]), .Z(n619) );
  NOR U1858 ( .A(n2147), .B(n619), .Z(n2149) );
  IV U1859 ( .A(a[381]), .Z(n2144) );
  IV U1860 ( .A(b[381]), .Z(n620) );
  NOR U1861 ( .A(n2144), .B(n620), .Z(n2146) );
  IV U1862 ( .A(a[380]), .Z(n2141) );
  IV U1863 ( .A(b[380]), .Z(n621) );
  NOR U1864 ( .A(n2141), .B(n621), .Z(n2143) );
  IV U1865 ( .A(a[379]), .Z(n2138) );
  IV U1866 ( .A(b[379]), .Z(n622) );
  NOR U1867 ( .A(n2138), .B(n622), .Z(n2140) );
  IV U1868 ( .A(a[378]), .Z(n2135) );
  IV U1869 ( .A(b[378]), .Z(n623) );
  NOR U1870 ( .A(n2135), .B(n623), .Z(n2137) );
  IV U1871 ( .A(a[377]), .Z(n2132) );
  IV U1872 ( .A(b[377]), .Z(n624) );
  NOR U1873 ( .A(n2132), .B(n624), .Z(n2134) );
  IV U1874 ( .A(a[376]), .Z(n2129) );
  IV U1875 ( .A(b[376]), .Z(n625) );
  NOR U1876 ( .A(n2129), .B(n625), .Z(n2131) );
  IV U1877 ( .A(a[375]), .Z(n2126) );
  IV U1878 ( .A(b[375]), .Z(n626) );
  NOR U1879 ( .A(n2126), .B(n626), .Z(n2128) );
  IV U1880 ( .A(a[374]), .Z(n2123) );
  IV U1881 ( .A(b[374]), .Z(n627) );
  NOR U1882 ( .A(n2123), .B(n627), .Z(n2125) );
  IV U1883 ( .A(a[373]), .Z(n2120) );
  IV U1884 ( .A(b[373]), .Z(n628) );
  NOR U1885 ( .A(n2120), .B(n628), .Z(n2122) );
  IV U1886 ( .A(a[372]), .Z(n2117) );
  IV U1887 ( .A(b[372]), .Z(n629) );
  NOR U1888 ( .A(n2117), .B(n629), .Z(n2119) );
  IV U1889 ( .A(a[371]), .Z(n2114) );
  IV U1890 ( .A(b[371]), .Z(n630) );
  NOR U1891 ( .A(n2114), .B(n630), .Z(n2116) );
  IV U1892 ( .A(a[370]), .Z(n2111) );
  IV U1893 ( .A(b[370]), .Z(n631) );
  NOR U1894 ( .A(n2111), .B(n631), .Z(n2113) );
  IV U1895 ( .A(a[369]), .Z(n2108) );
  IV U1896 ( .A(b[369]), .Z(n632) );
  NOR U1897 ( .A(n2108), .B(n632), .Z(n2110) );
  IV U1898 ( .A(a[368]), .Z(n2105) );
  IV U1899 ( .A(b[368]), .Z(n633) );
  NOR U1900 ( .A(n2105), .B(n633), .Z(n2107) );
  IV U1901 ( .A(a[367]), .Z(n2102) );
  IV U1902 ( .A(b[367]), .Z(n634) );
  NOR U1903 ( .A(n2102), .B(n634), .Z(n2104) );
  IV U1904 ( .A(a[366]), .Z(n2099) );
  IV U1905 ( .A(b[366]), .Z(n635) );
  NOR U1906 ( .A(n2099), .B(n635), .Z(n2101) );
  IV U1907 ( .A(a[365]), .Z(n2096) );
  IV U1908 ( .A(b[365]), .Z(n636) );
  NOR U1909 ( .A(n2096), .B(n636), .Z(n2098) );
  IV U1910 ( .A(a[364]), .Z(n2093) );
  IV U1911 ( .A(b[364]), .Z(n637) );
  NOR U1912 ( .A(n2093), .B(n637), .Z(n2095) );
  IV U1913 ( .A(a[363]), .Z(n2090) );
  IV U1914 ( .A(b[363]), .Z(n638) );
  NOR U1915 ( .A(n2090), .B(n638), .Z(n2092) );
  IV U1916 ( .A(a[362]), .Z(n2087) );
  IV U1917 ( .A(b[362]), .Z(n639) );
  NOR U1918 ( .A(n2087), .B(n639), .Z(n2089) );
  IV U1919 ( .A(a[361]), .Z(n2084) );
  IV U1920 ( .A(b[361]), .Z(n640) );
  NOR U1921 ( .A(n2084), .B(n640), .Z(n2086) );
  IV U1922 ( .A(a[360]), .Z(n2081) );
  IV U1923 ( .A(b[360]), .Z(n641) );
  NOR U1924 ( .A(n2081), .B(n641), .Z(n2083) );
  IV U1925 ( .A(a[359]), .Z(n2078) );
  IV U1926 ( .A(b[359]), .Z(n642) );
  NOR U1927 ( .A(n2078), .B(n642), .Z(n2080) );
  IV U1928 ( .A(a[358]), .Z(n2075) );
  IV U1929 ( .A(b[358]), .Z(n643) );
  NOR U1930 ( .A(n2075), .B(n643), .Z(n2077) );
  IV U1931 ( .A(a[357]), .Z(n2072) );
  IV U1932 ( .A(b[357]), .Z(n644) );
  NOR U1933 ( .A(n2072), .B(n644), .Z(n2074) );
  IV U1934 ( .A(a[356]), .Z(n2069) );
  IV U1935 ( .A(b[356]), .Z(n645) );
  NOR U1936 ( .A(n2069), .B(n645), .Z(n2071) );
  IV U1937 ( .A(a[355]), .Z(n2066) );
  IV U1938 ( .A(b[355]), .Z(n646) );
  NOR U1939 ( .A(n2066), .B(n646), .Z(n2068) );
  IV U1940 ( .A(a[354]), .Z(n2063) );
  IV U1941 ( .A(b[354]), .Z(n647) );
  NOR U1942 ( .A(n2063), .B(n647), .Z(n2065) );
  IV U1943 ( .A(a[353]), .Z(n2060) );
  IV U1944 ( .A(b[353]), .Z(n648) );
  NOR U1945 ( .A(n2060), .B(n648), .Z(n2062) );
  IV U1946 ( .A(a[352]), .Z(n2057) );
  IV U1947 ( .A(b[352]), .Z(n649) );
  NOR U1948 ( .A(n2057), .B(n649), .Z(n2059) );
  IV U1949 ( .A(a[351]), .Z(n2054) );
  IV U1950 ( .A(b[351]), .Z(n650) );
  NOR U1951 ( .A(n2054), .B(n650), .Z(n2056) );
  IV U1952 ( .A(a[350]), .Z(n2051) );
  IV U1953 ( .A(b[350]), .Z(n651) );
  NOR U1954 ( .A(n2051), .B(n651), .Z(n2053) );
  IV U1955 ( .A(a[349]), .Z(n2048) );
  IV U1956 ( .A(b[349]), .Z(n652) );
  NOR U1957 ( .A(n2048), .B(n652), .Z(n2050) );
  IV U1958 ( .A(a[348]), .Z(n2045) );
  IV U1959 ( .A(b[348]), .Z(n653) );
  NOR U1960 ( .A(n2045), .B(n653), .Z(n2047) );
  IV U1961 ( .A(a[347]), .Z(n2042) );
  IV U1962 ( .A(b[347]), .Z(n654) );
  NOR U1963 ( .A(n2042), .B(n654), .Z(n2044) );
  IV U1964 ( .A(a[346]), .Z(n2039) );
  IV U1965 ( .A(b[346]), .Z(n655) );
  NOR U1966 ( .A(n2039), .B(n655), .Z(n2041) );
  IV U1967 ( .A(a[345]), .Z(n2036) );
  IV U1968 ( .A(b[345]), .Z(n656) );
  NOR U1969 ( .A(n2036), .B(n656), .Z(n2038) );
  IV U1970 ( .A(a[344]), .Z(n2033) );
  IV U1971 ( .A(b[344]), .Z(n657) );
  NOR U1972 ( .A(n2033), .B(n657), .Z(n2035) );
  IV U1973 ( .A(a[343]), .Z(n2030) );
  IV U1974 ( .A(b[343]), .Z(n658) );
  NOR U1975 ( .A(n2030), .B(n658), .Z(n2032) );
  IV U1976 ( .A(a[342]), .Z(n2027) );
  IV U1977 ( .A(b[342]), .Z(n659) );
  NOR U1978 ( .A(n2027), .B(n659), .Z(n2029) );
  IV U1979 ( .A(a[341]), .Z(n2024) );
  IV U1980 ( .A(b[341]), .Z(n660) );
  NOR U1981 ( .A(n2024), .B(n660), .Z(n2026) );
  IV U1982 ( .A(a[340]), .Z(n2021) );
  IV U1983 ( .A(b[340]), .Z(n661) );
  NOR U1984 ( .A(n2021), .B(n661), .Z(n2023) );
  IV U1985 ( .A(a[339]), .Z(n2018) );
  IV U1986 ( .A(b[339]), .Z(n662) );
  NOR U1987 ( .A(n2018), .B(n662), .Z(n2020) );
  IV U1988 ( .A(a[338]), .Z(n2015) );
  IV U1989 ( .A(b[338]), .Z(n663) );
  NOR U1990 ( .A(n2015), .B(n663), .Z(n2017) );
  IV U1991 ( .A(a[337]), .Z(n2012) );
  IV U1992 ( .A(b[337]), .Z(n664) );
  NOR U1993 ( .A(n2012), .B(n664), .Z(n2014) );
  IV U1994 ( .A(a[336]), .Z(n2009) );
  IV U1995 ( .A(b[336]), .Z(n665) );
  NOR U1996 ( .A(n2009), .B(n665), .Z(n2011) );
  IV U1997 ( .A(a[335]), .Z(n2006) );
  IV U1998 ( .A(b[335]), .Z(n666) );
  NOR U1999 ( .A(n2006), .B(n666), .Z(n2008) );
  IV U2000 ( .A(a[334]), .Z(n2003) );
  IV U2001 ( .A(b[334]), .Z(n667) );
  NOR U2002 ( .A(n2003), .B(n667), .Z(n2005) );
  IV U2003 ( .A(a[333]), .Z(n2000) );
  IV U2004 ( .A(b[333]), .Z(n668) );
  NOR U2005 ( .A(n2000), .B(n668), .Z(n2002) );
  IV U2006 ( .A(a[332]), .Z(n1997) );
  IV U2007 ( .A(b[332]), .Z(n669) );
  NOR U2008 ( .A(n1997), .B(n669), .Z(n1999) );
  IV U2009 ( .A(a[331]), .Z(n1994) );
  IV U2010 ( .A(b[331]), .Z(n670) );
  NOR U2011 ( .A(n1994), .B(n670), .Z(n1996) );
  IV U2012 ( .A(a[330]), .Z(n1991) );
  IV U2013 ( .A(b[330]), .Z(n671) );
  NOR U2014 ( .A(n1991), .B(n671), .Z(n1993) );
  IV U2015 ( .A(a[329]), .Z(n1988) );
  IV U2016 ( .A(b[329]), .Z(n672) );
  NOR U2017 ( .A(n1988), .B(n672), .Z(n1990) );
  IV U2018 ( .A(a[328]), .Z(n1985) );
  IV U2019 ( .A(b[328]), .Z(n673) );
  NOR U2020 ( .A(n1985), .B(n673), .Z(n1987) );
  IV U2021 ( .A(a[327]), .Z(n1982) );
  IV U2022 ( .A(b[327]), .Z(n674) );
  NOR U2023 ( .A(n1982), .B(n674), .Z(n1984) );
  IV U2024 ( .A(a[326]), .Z(n1979) );
  IV U2025 ( .A(b[326]), .Z(n675) );
  NOR U2026 ( .A(n1979), .B(n675), .Z(n1981) );
  IV U2027 ( .A(a[325]), .Z(n1976) );
  IV U2028 ( .A(b[325]), .Z(n676) );
  NOR U2029 ( .A(n1976), .B(n676), .Z(n1978) );
  IV U2030 ( .A(a[324]), .Z(n1973) );
  IV U2031 ( .A(b[324]), .Z(n677) );
  NOR U2032 ( .A(n1973), .B(n677), .Z(n1975) );
  IV U2033 ( .A(a[323]), .Z(n1970) );
  IV U2034 ( .A(b[323]), .Z(n678) );
  NOR U2035 ( .A(n1970), .B(n678), .Z(n1972) );
  IV U2036 ( .A(a[322]), .Z(n1967) );
  IV U2037 ( .A(b[322]), .Z(n679) );
  NOR U2038 ( .A(n1967), .B(n679), .Z(n1969) );
  IV U2039 ( .A(a[321]), .Z(n1964) );
  IV U2040 ( .A(b[321]), .Z(n680) );
  NOR U2041 ( .A(n1964), .B(n680), .Z(n1966) );
  IV U2042 ( .A(a[320]), .Z(n1961) );
  IV U2043 ( .A(b[320]), .Z(n681) );
  NOR U2044 ( .A(n1961), .B(n681), .Z(n1963) );
  IV U2045 ( .A(a[319]), .Z(n1958) );
  IV U2046 ( .A(b[319]), .Z(n682) );
  NOR U2047 ( .A(n1958), .B(n682), .Z(n1960) );
  IV U2048 ( .A(a[318]), .Z(n1955) );
  IV U2049 ( .A(b[318]), .Z(n683) );
  NOR U2050 ( .A(n1955), .B(n683), .Z(n1957) );
  IV U2051 ( .A(a[317]), .Z(n1952) );
  IV U2052 ( .A(b[317]), .Z(n684) );
  NOR U2053 ( .A(n1952), .B(n684), .Z(n1954) );
  IV U2054 ( .A(a[316]), .Z(n1949) );
  IV U2055 ( .A(b[316]), .Z(n685) );
  NOR U2056 ( .A(n1949), .B(n685), .Z(n1951) );
  IV U2057 ( .A(a[315]), .Z(n1946) );
  IV U2058 ( .A(b[315]), .Z(n686) );
  NOR U2059 ( .A(n1946), .B(n686), .Z(n1948) );
  IV U2060 ( .A(a[314]), .Z(n1943) );
  IV U2061 ( .A(b[314]), .Z(n687) );
  NOR U2062 ( .A(n1943), .B(n687), .Z(n1945) );
  IV U2063 ( .A(a[313]), .Z(n1940) );
  IV U2064 ( .A(b[313]), .Z(n688) );
  NOR U2065 ( .A(n1940), .B(n688), .Z(n1942) );
  IV U2066 ( .A(a[312]), .Z(n1937) );
  IV U2067 ( .A(b[312]), .Z(n689) );
  NOR U2068 ( .A(n1937), .B(n689), .Z(n1939) );
  IV U2069 ( .A(a[311]), .Z(n1934) );
  IV U2070 ( .A(b[311]), .Z(n690) );
  NOR U2071 ( .A(n1934), .B(n690), .Z(n1936) );
  IV U2072 ( .A(a[310]), .Z(n1931) );
  IV U2073 ( .A(b[310]), .Z(n691) );
  NOR U2074 ( .A(n1931), .B(n691), .Z(n1933) );
  IV U2075 ( .A(a[309]), .Z(n1928) );
  IV U2076 ( .A(b[309]), .Z(n692) );
  NOR U2077 ( .A(n1928), .B(n692), .Z(n1930) );
  IV U2078 ( .A(a[308]), .Z(n1925) );
  IV U2079 ( .A(b[308]), .Z(n693) );
  NOR U2080 ( .A(n1925), .B(n693), .Z(n1927) );
  IV U2081 ( .A(a[307]), .Z(n1922) );
  IV U2082 ( .A(b[307]), .Z(n694) );
  NOR U2083 ( .A(n1922), .B(n694), .Z(n1924) );
  IV U2084 ( .A(a[306]), .Z(n1919) );
  IV U2085 ( .A(b[306]), .Z(n695) );
  NOR U2086 ( .A(n1919), .B(n695), .Z(n1921) );
  IV U2087 ( .A(a[305]), .Z(n1916) );
  IV U2088 ( .A(b[305]), .Z(n696) );
  NOR U2089 ( .A(n1916), .B(n696), .Z(n1918) );
  IV U2090 ( .A(a[304]), .Z(n1913) );
  IV U2091 ( .A(b[304]), .Z(n697) );
  NOR U2092 ( .A(n1913), .B(n697), .Z(n1915) );
  IV U2093 ( .A(a[303]), .Z(n1910) );
  IV U2094 ( .A(b[303]), .Z(n698) );
  NOR U2095 ( .A(n1910), .B(n698), .Z(n1912) );
  IV U2096 ( .A(a[302]), .Z(n1907) );
  IV U2097 ( .A(b[302]), .Z(n699) );
  NOR U2098 ( .A(n1907), .B(n699), .Z(n1909) );
  IV U2099 ( .A(a[301]), .Z(n1904) );
  IV U2100 ( .A(b[301]), .Z(n700) );
  NOR U2101 ( .A(n1904), .B(n700), .Z(n1906) );
  IV U2102 ( .A(a[300]), .Z(n1901) );
  IV U2103 ( .A(b[300]), .Z(n701) );
  NOR U2104 ( .A(n1901), .B(n701), .Z(n1903) );
  IV U2105 ( .A(a[299]), .Z(n1898) );
  IV U2106 ( .A(b[299]), .Z(n702) );
  NOR U2107 ( .A(n1898), .B(n702), .Z(n1900) );
  IV U2108 ( .A(a[298]), .Z(n1895) );
  IV U2109 ( .A(b[298]), .Z(n703) );
  NOR U2110 ( .A(n1895), .B(n703), .Z(n1897) );
  IV U2111 ( .A(a[297]), .Z(n1892) );
  IV U2112 ( .A(b[297]), .Z(n704) );
  NOR U2113 ( .A(n1892), .B(n704), .Z(n1894) );
  IV U2114 ( .A(a[296]), .Z(n1889) );
  IV U2115 ( .A(b[296]), .Z(n705) );
  NOR U2116 ( .A(n1889), .B(n705), .Z(n1891) );
  IV U2117 ( .A(a[295]), .Z(n1886) );
  IV U2118 ( .A(b[295]), .Z(n706) );
  NOR U2119 ( .A(n1886), .B(n706), .Z(n1888) );
  IV U2120 ( .A(a[294]), .Z(n1883) );
  IV U2121 ( .A(b[294]), .Z(n707) );
  NOR U2122 ( .A(n1883), .B(n707), .Z(n1885) );
  IV U2123 ( .A(a[293]), .Z(n1880) );
  IV U2124 ( .A(b[293]), .Z(n708) );
  NOR U2125 ( .A(n1880), .B(n708), .Z(n1882) );
  IV U2126 ( .A(a[292]), .Z(n1877) );
  IV U2127 ( .A(b[292]), .Z(n709) );
  NOR U2128 ( .A(n1877), .B(n709), .Z(n1879) );
  IV U2129 ( .A(a[291]), .Z(n1874) );
  IV U2130 ( .A(b[291]), .Z(n710) );
  NOR U2131 ( .A(n1874), .B(n710), .Z(n1876) );
  IV U2132 ( .A(a[290]), .Z(n1871) );
  IV U2133 ( .A(b[290]), .Z(n711) );
  NOR U2134 ( .A(n1871), .B(n711), .Z(n1873) );
  IV U2135 ( .A(a[289]), .Z(n1868) );
  IV U2136 ( .A(b[289]), .Z(n712) );
  NOR U2137 ( .A(n1868), .B(n712), .Z(n1870) );
  IV U2138 ( .A(a[288]), .Z(n1865) );
  IV U2139 ( .A(b[288]), .Z(n713) );
  NOR U2140 ( .A(n1865), .B(n713), .Z(n1867) );
  IV U2141 ( .A(a[287]), .Z(n1862) );
  IV U2142 ( .A(b[287]), .Z(n714) );
  NOR U2143 ( .A(n1862), .B(n714), .Z(n1864) );
  IV U2144 ( .A(a[286]), .Z(n1859) );
  IV U2145 ( .A(b[286]), .Z(n715) );
  NOR U2146 ( .A(n1859), .B(n715), .Z(n1861) );
  IV U2147 ( .A(a[285]), .Z(n1856) );
  IV U2148 ( .A(b[285]), .Z(n716) );
  NOR U2149 ( .A(n1856), .B(n716), .Z(n1858) );
  IV U2150 ( .A(a[284]), .Z(n1853) );
  IV U2151 ( .A(b[284]), .Z(n717) );
  NOR U2152 ( .A(n1853), .B(n717), .Z(n1855) );
  IV U2153 ( .A(a[283]), .Z(n1850) );
  IV U2154 ( .A(b[283]), .Z(n718) );
  NOR U2155 ( .A(n1850), .B(n718), .Z(n1852) );
  IV U2156 ( .A(a[282]), .Z(n1847) );
  IV U2157 ( .A(b[282]), .Z(n719) );
  NOR U2158 ( .A(n1847), .B(n719), .Z(n1849) );
  IV U2159 ( .A(a[281]), .Z(n1844) );
  IV U2160 ( .A(b[281]), .Z(n720) );
  NOR U2161 ( .A(n1844), .B(n720), .Z(n1846) );
  IV U2162 ( .A(a[280]), .Z(n1841) );
  IV U2163 ( .A(b[280]), .Z(n721) );
  NOR U2164 ( .A(n1841), .B(n721), .Z(n1843) );
  IV U2165 ( .A(a[279]), .Z(n1838) );
  IV U2166 ( .A(b[279]), .Z(n722) );
  NOR U2167 ( .A(n1838), .B(n722), .Z(n1840) );
  IV U2168 ( .A(a[278]), .Z(n1835) );
  IV U2169 ( .A(b[278]), .Z(n723) );
  NOR U2170 ( .A(n1835), .B(n723), .Z(n1837) );
  IV U2171 ( .A(a[277]), .Z(n1832) );
  IV U2172 ( .A(b[277]), .Z(n724) );
  NOR U2173 ( .A(n1832), .B(n724), .Z(n1834) );
  IV U2174 ( .A(a[276]), .Z(n1829) );
  IV U2175 ( .A(b[276]), .Z(n725) );
  NOR U2176 ( .A(n1829), .B(n725), .Z(n1831) );
  IV U2177 ( .A(a[275]), .Z(n1826) );
  IV U2178 ( .A(b[275]), .Z(n726) );
  NOR U2179 ( .A(n1826), .B(n726), .Z(n1828) );
  IV U2180 ( .A(a[274]), .Z(n1823) );
  IV U2181 ( .A(b[274]), .Z(n727) );
  NOR U2182 ( .A(n1823), .B(n727), .Z(n1825) );
  IV U2183 ( .A(a[273]), .Z(n1820) );
  IV U2184 ( .A(b[273]), .Z(n728) );
  NOR U2185 ( .A(n1820), .B(n728), .Z(n1822) );
  IV U2186 ( .A(a[272]), .Z(n1817) );
  IV U2187 ( .A(b[272]), .Z(n729) );
  NOR U2188 ( .A(n1817), .B(n729), .Z(n1819) );
  IV U2189 ( .A(a[271]), .Z(n1814) );
  IV U2190 ( .A(b[271]), .Z(n730) );
  NOR U2191 ( .A(n1814), .B(n730), .Z(n1816) );
  IV U2192 ( .A(a[270]), .Z(n1811) );
  IV U2193 ( .A(b[270]), .Z(n731) );
  NOR U2194 ( .A(n1811), .B(n731), .Z(n1813) );
  IV U2195 ( .A(a[269]), .Z(n1808) );
  IV U2196 ( .A(b[269]), .Z(n732) );
  NOR U2197 ( .A(n1808), .B(n732), .Z(n1810) );
  IV U2198 ( .A(a[268]), .Z(n1805) );
  IV U2199 ( .A(b[268]), .Z(n733) );
  NOR U2200 ( .A(n1805), .B(n733), .Z(n1807) );
  IV U2201 ( .A(a[267]), .Z(n1802) );
  IV U2202 ( .A(b[267]), .Z(n734) );
  NOR U2203 ( .A(n1802), .B(n734), .Z(n1804) );
  IV U2204 ( .A(a[266]), .Z(n1799) );
  IV U2205 ( .A(b[266]), .Z(n735) );
  NOR U2206 ( .A(n1799), .B(n735), .Z(n1801) );
  IV U2207 ( .A(a[265]), .Z(n1796) );
  IV U2208 ( .A(b[265]), .Z(n736) );
  NOR U2209 ( .A(n1796), .B(n736), .Z(n1798) );
  IV U2210 ( .A(a[264]), .Z(n1793) );
  IV U2211 ( .A(b[264]), .Z(n737) );
  NOR U2212 ( .A(n1793), .B(n737), .Z(n1795) );
  IV U2213 ( .A(a[263]), .Z(n1790) );
  IV U2214 ( .A(b[263]), .Z(n738) );
  NOR U2215 ( .A(n1790), .B(n738), .Z(n1792) );
  IV U2216 ( .A(a[262]), .Z(n1787) );
  IV U2217 ( .A(b[262]), .Z(n739) );
  NOR U2218 ( .A(n1787), .B(n739), .Z(n1789) );
  IV U2219 ( .A(a[261]), .Z(n1784) );
  IV U2220 ( .A(b[261]), .Z(n740) );
  NOR U2221 ( .A(n1784), .B(n740), .Z(n1786) );
  IV U2222 ( .A(a[260]), .Z(n1781) );
  IV U2223 ( .A(b[260]), .Z(n741) );
  NOR U2224 ( .A(n1781), .B(n741), .Z(n1783) );
  IV U2225 ( .A(a[259]), .Z(n1778) );
  IV U2226 ( .A(b[259]), .Z(n742) );
  NOR U2227 ( .A(n1778), .B(n742), .Z(n1780) );
  IV U2228 ( .A(a[258]), .Z(n1775) );
  IV U2229 ( .A(b[258]), .Z(n743) );
  NOR U2230 ( .A(n1775), .B(n743), .Z(n1777) );
  IV U2231 ( .A(a[257]), .Z(n1772) );
  IV U2232 ( .A(b[257]), .Z(n744) );
  NOR U2233 ( .A(n1772), .B(n744), .Z(n1774) );
  IV U2234 ( .A(a[256]), .Z(n1769) );
  IV U2235 ( .A(b[256]), .Z(n745) );
  NOR U2236 ( .A(n1769), .B(n745), .Z(n1771) );
  IV U2237 ( .A(a[255]), .Z(n1766) );
  IV U2238 ( .A(b[255]), .Z(n746) );
  NOR U2239 ( .A(n1766), .B(n746), .Z(n1768) );
  IV U2240 ( .A(a[254]), .Z(n1763) );
  IV U2241 ( .A(b[254]), .Z(n747) );
  NOR U2242 ( .A(n1763), .B(n747), .Z(n1765) );
  IV U2243 ( .A(a[253]), .Z(n1760) );
  IV U2244 ( .A(b[253]), .Z(n748) );
  NOR U2245 ( .A(n1760), .B(n748), .Z(n1762) );
  IV U2246 ( .A(a[252]), .Z(n1757) );
  IV U2247 ( .A(b[252]), .Z(n749) );
  NOR U2248 ( .A(n1757), .B(n749), .Z(n1759) );
  IV U2249 ( .A(a[251]), .Z(n1754) );
  IV U2250 ( .A(b[251]), .Z(n750) );
  NOR U2251 ( .A(n1754), .B(n750), .Z(n1756) );
  IV U2252 ( .A(a[250]), .Z(n1751) );
  IV U2253 ( .A(b[250]), .Z(n751) );
  NOR U2254 ( .A(n1751), .B(n751), .Z(n1753) );
  IV U2255 ( .A(a[249]), .Z(n1748) );
  IV U2256 ( .A(b[249]), .Z(n752) );
  NOR U2257 ( .A(n1748), .B(n752), .Z(n1750) );
  IV U2258 ( .A(a[248]), .Z(n1745) );
  IV U2259 ( .A(b[248]), .Z(n753) );
  NOR U2260 ( .A(n1745), .B(n753), .Z(n1747) );
  IV U2261 ( .A(a[247]), .Z(n1742) );
  IV U2262 ( .A(b[247]), .Z(n754) );
  NOR U2263 ( .A(n1742), .B(n754), .Z(n1744) );
  IV U2264 ( .A(a[246]), .Z(n1739) );
  IV U2265 ( .A(b[246]), .Z(n755) );
  NOR U2266 ( .A(n1739), .B(n755), .Z(n1741) );
  IV U2267 ( .A(a[245]), .Z(n1736) );
  IV U2268 ( .A(b[245]), .Z(n756) );
  NOR U2269 ( .A(n1736), .B(n756), .Z(n1738) );
  IV U2270 ( .A(a[244]), .Z(n1733) );
  IV U2271 ( .A(b[244]), .Z(n757) );
  NOR U2272 ( .A(n1733), .B(n757), .Z(n1735) );
  IV U2273 ( .A(a[243]), .Z(n1730) );
  IV U2274 ( .A(b[243]), .Z(n758) );
  NOR U2275 ( .A(n1730), .B(n758), .Z(n1732) );
  IV U2276 ( .A(a[242]), .Z(n1727) );
  IV U2277 ( .A(b[242]), .Z(n759) );
  NOR U2278 ( .A(n1727), .B(n759), .Z(n1729) );
  IV U2279 ( .A(a[241]), .Z(n1724) );
  IV U2280 ( .A(b[241]), .Z(n760) );
  NOR U2281 ( .A(n1724), .B(n760), .Z(n1726) );
  IV U2282 ( .A(a[240]), .Z(n1721) );
  IV U2283 ( .A(b[240]), .Z(n761) );
  NOR U2284 ( .A(n1721), .B(n761), .Z(n1723) );
  IV U2285 ( .A(a[239]), .Z(n1718) );
  IV U2286 ( .A(b[239]), .Z(n762) );
  NOR U2287 ( .A(n1718), .B(n762), .Z(n1720) );
  IV U2288 ( .A(a[238]), .Z(n1715) );
  IV U2289 ( .A(b[238]), .Z(n763) );
  NOR U2290 ( .A(n1715), .B(n763), .Z(n1717) );
  IV U2291 ( .A(a[237]), .Z(n1712) );
  IV U2292 ( .A(b[237]), .Z(n764) );
  NOR U2293 ( .A(n1712), .B(n764), .Z(n1714) );
  IV U2294 ( .A(a[236]), .Z(n1709) );
  IV U2295 ( .A(b[236]), .Z(n765) );
  NOR U2296 ( .A(n1709), .B(n765), .Z(n1711) );
  IV U2297 ( .A(a[235]), .Z(n1706) );
  IV U2298 ( .A(b[235]), .Z(n766) );
  NOR U2299 ( .A(n1706), .B(n766), .Z(n1708) );
  IV U2300 ( .A(a[234]), .Z(n1703) );
  IV U2301 ( .A(b[234]), .Z(n767) );
  NOR U2302 ( .A(n1703), .B(n767), .Z(n1705) );
  IV U2303 ( .A(a[233]), .Z(n1700) );
  IV U2304 ( .A(b[233]), .Z(n768) );
  NOR U2305 ( .A(n1700), .B(n768), .Z(n1702) );
  IV U2306 ( .A(a[232]), .Z(n1697) );
  IV U2307 ( .A(b[232]), .Z(n769) );
  NOR U2308 ( .A(n1697), .B(n769), .Z(n1699) );
  IV U2309 ( .A(a[231]), .Z(n1694) );
  IV U2310 ( .A(b[231]), .Z(n770) );
  NOR U2311 ( .A(n1694), .B(n770), .Z(n1696) );
  IV U2312 ( .A(a[230]), .Z(n1691) );
  IV U2313 ( .A(b[230]), .Z(n771) );
  NOR U2314 ( .A(n1691), .B(n771), .Z(n1693) );
  IV U2315 ( .A(a[229]), .Z(n1688) );
  IV U2316 ( .A(b[229]), .Z(n772) );
  NOR U2317 ( .A(n1688), .B(n772), .Z(n1690) );
  IV U2318 ( .A(a[228]), .Z(n1685) );
  IV U2319 ( .A(b[228]), .Z(n773) );
  NOR U2320 ( .A(n1685), .B(n773), .Z(n1687) );
  IV U2321 ( .A(a[227]), .Z(n1682) );
  IV U2322 ( .A(b[227]), .Z(n774) );
  NOR U2323 ( .A(n1682), .B(n774), .Z(n1684) );
  IV U2324 ( .A(a[226]), .Z(n1679) );
  IV U2325 ( .A(b[226]), .Z(n775) );
  NOR U2326 ( .A(n1679), .B(n775), .Z(n1681) );
  IV U2327 ( .A(a[225]), .Z(n1676) );
  IV U2328 ( .A(b[225]), .Z(n776) );
  NOR U2329 ( .A(n1676), .B(n776), .Z(n1678) );
  IV U2330 ( .A(a[224]), .Z(n1673) );
  IV U2331 ( .A(b[224]), .Z(n777) );
  NOR U2332 ( .A(n1673), .B(n777), .Z(n1675) );
  IV U2333 ( .A(a[223]), .Z(n1670) );
  IV U2334 ( .A(b[223]), .Z(n778) );
  NOR U2335 ( .A(n1670), .B(n778), .Z(n1672) );
  IV U2336 ( .A(a[222]), .Z(n1667) );
  IV U2337 ( .A(b[222]), .Z(n779) );
  NOR U2338 ( .A(n1667), .B(n779), .Z(n1669) );
  IV U2339 ( .A(a[221]), .Z(n1664) );
  IV U2340 ( .A(b[221]), .Z(n780) );
  NOR U2341 ( .A(n1664), .B(n780), .Z(n1666) );
  IV U2342 ( .A(a[220]), .Z(n1661) );
  IV U2343 ( .A(b[220]), .Z(n781) );
  NOR U2344 ( .A(n1661), .B(n781), .Z(n1663) );
  IV U2345 ( .A(a[219]), .Z(n1658) );
  IV U2346 ( .A(b[219]), .Z(n782) );
  NOR U2347 ( .A(n1658), .B(n782), .Z(n1660) );
  IV U2348 ( .A(a[218]), .Z(n1655) );
  IV U2349 ( .A(b[218]), .Z(n783) );
  NOR U2350 ( .A(n1655), .B(n783), .Z(n1657) );
  IV U2351 ( .A(a[217]), .Z(n1652) );
  IV U2352 ( .A(b[217]), .Z(n784) );
  NOR U2353 ( .A(n1652), .B(n784), .Z(n1654) );
  IV U2354 ( .A(a[216]), .Z(n1649) );
  IV U2355 ( .A(b[216]), .Z(n785) );
  NOR U2356 ( .A(n1649), .B(n785), .Z(n1651) );
  IV U2357 ( .A(a[215]), .Z(n1646) );
  IV U2358 ( .A(b[215]), .Z(n786) );
  NOR U2359 ( .A(n1646), .B(n786), .Z(n1648) );
  IV U2360 ( .A(a[214]), .Z(n1643) );
  IV U2361 ( .A(b[214]), .Z(n787) );
  NOR U2362 ( .A(n1643), .B(n787), .Z(n1645) );
  IV U2363 ( .A(a[213]), .Z(n1640) );
  IV U2364 ( .A(b[213]), .Z(n788) );
  NOR U2365 ( .A(n1640), .B(n788), .Z(n1642) );
  IV U2366 ( .A(a[212]), .Z(n1637) );
  IV U2367 ( .A(b[212]), .Z(n789) );
  NOR U2368 ( .A(n1637), .B(n789), .Z(n1639) );
  IV U2369 ( .A(a[211]), .Z(n1634) );
  IV U2370 ( .A(b[211]), .Z(n790) );
  NOR U2371 ( .A(n1634), .B(n790), .Z(n1636) );
  IV U2372 ( .A(a[210]), .Z(n1631) );
  IV U2373 ( .A(b[210]), .Z(n791) );
  NOR U2374 ( .A(n1631), .B(n791), .Z(n1633) );
  IV U2375 ( .A(a[209]), .Z(n1628) );
  IV U2376 ( .A(b[209]), .Z(n792) );
  NOR U2377 ( .A(n1628), .B(n792), .Z(n1630) );
  IV U2378 ( .A(a[208]), .Z(n1625) );
  IV U2379 ( .A(b[208]), .Z(n793) );
  NOR U2380 ( .A(n1625), .B(n793), .Z(n1627) );
  IV U2381 ( .A(a[207]), .Z(n1622) );
  IV U2382 ( .A(b[207]), .Z(n794) );
  NOR U2383 ( .A(n1622), .B(n794), .Z(n1624) );
  IV U2384 ( .A(a[206]), .Z(n1619) );
  IV U2385 ( .A(b[206]), .Z(n795) );
  NOR U2386 ( .A(n1619), .B(n795), .Z(n1621) );
  IV U2387 ( .A(a[205]), .Z(n1616) );
  IV U2388 ( .A(b[205]), .Z(n796) );
  NOR U2389 ( .A(n1616), .B(n796), .Z(n1618) );
  IV U2390 ( .A(a[204]), .Z(n1613) );
  IV U2391 ( .A(b[204]), .Z(n797) );
  NOR U2392 ( .A(n1613), .B(n797), .Z(n1615) );
  IV U2393 ( .A(a[203]), .Z(n1610) );
  IV U2394 ( .A(b[203]), .Z(n798) );
  NOR U2395 ( .A(n1610), .B(n798), .Z(n1612) );
  IV U2396 ( .A(a[202]), .Z(n1607) );
  IV U2397 ( .A(b[202]), .Z(n799) );
  NOR U2398 ( .A(n1607), .B(n799), .Z(n1609) );
  IV U2399 ( .A(a[201]), .Z(n1604) );
  IV U2400 ( .A(b[201]), .Z(n800) );
  NOR U2401 ( .A(n1604), .B(n800), .Z(n1606) );
  IV U2402 ( .A(a[200]), .Z(n1601) );
  IV U2403 ( .A(b[200]), .Z(n801) );
  NOR U2404 ( .A(n1601), .B(n801), .Z(n1603) );
  IV U2405 ( .A(a[199]), .Z(n1598) );
  IV U2406 ( .A(b[199]), .Z(n802) );
  NOR U2407 ( .A(n1598), .B(n802), .Z(n1600) );
  IV U2408 ( .A(a[198]), .Z(n1595) );
  IV U2409 ( .A(b[198]), .Z(n803) );
  NOR U2410 ( .A(n1595), .B(n803), .Z(n1597) );
  IV U2411 ( .A(a[197]), .Z(n1592) );
  IV U2412 ( .A(b[197]), .Z(n804) );
  NOR U2413 ( .A(n1592), .B(n804), .Z(n1594) );
  IV U2414 ( .A(a[196]), .Z(n1589) );
  IV U2415 ( .A(b[196]), .Z(n805) );
  NOR U2416 ( .A(n1589), .B(n805), .Z(n1591) );
  IV U2417 ( .A(a[195]), .Z(n1586) );
  IV U2418 ( .A(b[195]), .Z(n806) );
  NOR U2419 ( .A(n1586), .B(n806), .Z(n1588) );
  IV U2420 ( .A(a[194]), .Z(n1583) );
  IV U2421 ( .A(b[194]), .Z(n807) );
  NOR U2422 ( .A(n1583), .B(n807), .Z(n1585) );
  IV U2423 ( .A(a[193]), .Z(n1580) );
  IV U2424 ( .A(b[193]), .Z(n808) );
  NOR U2425 ( .A(n1580), .B(n808), .Z(n1582) );
  IV U2426 ( .A(a[192]), .Z(n1577) );
  IV U2427 ( .A(b[192]), .Z(n809) );
  NOR U2428 ( .A(n1577), .B(n809), .Z(n1579) );
  IV U2429 ( .A(a[191]), .Z(n1574) );
  IV U2430 ( .A(b[191]), .Z(n810) );
  NOR U2431 ( .A(n1574), .B(n810), .Z(n1576) );
  IV U2432 ( .A(a[190]), .Z(n1571) );
  IV U2433 ( .A(b[190]), .Z(n811) );
  NOR U2434 ( .A(n1571), .B(n811), .Z(n1573) );
  IV U2435 ( .A(a[189]), .Z(n1568) );
  IV U2436 ( .A(b[189]), .Z(n812) );
  NOR U2437 ( .A(n1568), .B(n812), .Z(n1570) );
  IV U2438 ( .A(a[188]), .Z(n1565) );
  IV U2439 ( .A(b[188]), .Z(n813) );
  NOR U2440 ( .A(n1565), .B(n813), .Z(n1567) );
  IV U2441 ( .A(a[187]), .Z(n1562) );
  IV U2442 ( .A(b[187]), .Z(n814) );
  NOR U2443 ( .A(n1562), .B(n814), .Z(n1564) );
  IV U2444 ( .A(a[186]), .Z(n1559) );
  IV U2445 ( .A(b[186]), .Z(n815) );
  NOR U2446 ( .A(n1559), .B(n815), .Z(n1561) );
  IV U2447 ( .A(a[185]), .Z(n1556) );
  IV U2448 ( .A(b[185]), .Z(n816) );
  NOR U2449 ( .A(n1556), .B(n816), .Z(n1558) );
  IV U2450 ( .A(a[184]), .Z(n1553) );
  IV U2451 ( .A(b[184]), .Z(n817) );
  NOR U2452 ( .A(n1553), .B(n817), .Z(n1555) );
  IV U2453 ( .A(a[183]), .Z(n1550) );
  IV U2454 ( .A(b[183]), .Z(n818) );
  NOR U2455 ( .A(n1550), .B(n818), .Z(n1552) );
  IV U2456 ( .A(a[182]), .Z(n1547) );
  IV U2457 ( .A(b[182]), .Z(n819) );
  NOR U2458 ( .A(n1547), .B(n819), .Z(n1549) );
  IV U2459 ( .A(a[181]), .Z(n1544) );
  IV U2460 ( .A(b[181]), .Z(n820) );
  NOR U2461 ( .A(n1544), .B(n820), .Z(n1546) );
  IV U2462 ( .A(a[180]), .Z(n1541) );
  IV U2463 ( .A(b[180]), .Z(n821) );
  NOR U2464 ( .A(n1541), .B(n821), .Z(n1543) );
  IV U2465 ( .A(a[179]), .Z(n1538) );
  IV U2466 ( .A(b[179]), .Z(n822) );
  NOR U2467 ( .A(n1538), .B(n822), .Z(n1540) );
  IV U2468 ( .A(a[178]), .Z(n1535) );
  IV U2469 ( .A(b[178]), .Z(n823) );
  NOR U2470 ( .A(n1535), .B(n823), .Z(n1537) );
  IV U2471 ( .A(a[177]), .Z(n1532) );
  IV U2472 ( .A(b[177]), .Z(n824) );
  NOR U2473 ( .A(n1532), .B(n824), .Z(n1534) );
  IV U2474 ( .A(a[176]), .Z(n1529) );
  IV U2475 ( .A(b[176]), .Z(n825) );
  NOR U2476 ( .A(n1529), .B(n825), .Z(n1531) );
  IV U2477 ( .A(a[175]), .Z(n1526) );
  IV U2478 ( .A(b[175]), .Z(n826) );
  NOR U2479 ( .A(n1526), .B(n826), .Z(n1528) );
  IV U2480 ( .A(a[174]), .Z(n1523) );
  IV U2481 ( .A(b[174]), .Z(n827) );
  NOR U2482 ( .A(n1523), .B(n827), .Z(n1525) );
  IV U2483 ( .A(a[173]), .Z(n1520) );
  IV U2484 ( .A(b[173]), .Z(n828) );
  NOR U2485 ( .A(n1520), .B(n828), .Z(n1522) );
  IV U2486 ( .A(a[172]), .Z(n1517) );
  IV U2487 ( .A(b[172]), .Z(n829) );
  NOR U2488 ( .A(n1517), .B(n829), .Z(n1519) );
  IV U2489 ( .A(a[171]), .Z(n1514) );
  IV U2490 ( .A(b[171]), .Z(n830) );
  NOR U2491 ( .A(n1514), .B(n830), .Z(n1516) );
  IV U2492 ( .A(a[170]), .Z(n1511) );
  IV U2493 ( .A(b[170]), .Z(n831) );
  NOR U2494 ( .A(n1511), .B(n831), .Z(n1513) );
  IV U2495 ( .A(a[169]), .Z(n1508) );
  IV U2496 ( .A(b[169]), .Z(n832) );
  NOR U2497 ( .A(n1508), .B(n832), .Z(n1510) );
  IV U2498 ( .A(a[168]), .Z(n1505) );
  IV U2499 ( .A(b[168]), .Z(n833) );
  NOR U2500 ( .A(n1505), .B(n833), .Z(n1507) );
  IV U2501 ( .A(a[167]), .Z(n1502) );
  IV U2502 ( .A(b[167]), .Z(n834) );
  NOR U2503 ( .A(n1502), .B(n834), .Z(n1504) );
  IV U2504 ( .A(a[166]), .Z(n1499) );
  IV U2505 ( .A(b[166]), .Z(n835) );
  NOR U2506 ( .A(n1499), .B(n835), .Z(n1501) );
  IV U2507 ( .A(a[165]), .Z(n1496) );
  IV U2508 ( .A(b[165]), .Z(n836) );
  NOR U2509 ( .A(n1496), .B(n836), .Z(n1498) );
  IV U2510 ( .A(a[164]), .Z(n1493) );
  IV U2511 ( .A(b[164]), .Z(n837) );
  NOR U2512 ( .A(n1493), .B(n837), .Z(n1495) );
  IV U2513 ( .A(a[163]), .Z(n1490) );
  IV U2514 ( .A(b[163]), .Z(n838) );
  NOR U2515 ( .A(n1490), .B(n838), .Z(n1492) );
  IV U2516 ( .A(a[162]), .Z(n1487) );
  IV U2517 ( .A(b[162]), .Z(n839) );
  NOR U2518 ( .A(n1487), .B(n839), .Z(n1489) );
  IV U2519 ( .A(a[161]), .Z(n1484) );
  IV U2520 ( .A(b[161]), .Z(n840) );
  NOR U2521 ( .A(n1484), .B(n840), .Z(n1486) );
  IV U2522 ( .A(a[160]), .Z(n1481) );
  IV U2523 ( .A(b[160]), .Z(n841) );
  NOR U2524 ( .A(n1481), .B(n841), .Z(n1483) );
  IV U2525 ( .A(a[159]), .Z(n1478) );
  IV U2526 ( .A(b[159]), .Z(n842) );
  NOR U2527 ( .A(n1478), .B(n842), .Z(n1480) );
  IV U2528 ( .A(a[158]), .Z(n1475) );
  IV U2529 ( .A(b[158]), .Z(n843) );
  NOR U2530 ( .A(n1475), .B(n843), .Z(n1477) );
  IV U2531 ( .A(a[157]), .Z(n1472) );
  IV U2532 ( .A(b[157]), .Z(n844) );
  NOR U2533 ( .A(n1472), .B(n844), .Z(n1474) );
  IV U2534 ( .A(a[156]), .Z(n1469) );
  IV U2535 ( .A(b[156]), .Z(n845) );
  NOR U2536 ( .A(n1469), .B(n845), .Z(n1471) );
  IV U2537 ( .A(a[155]), .Z(n1466) );
  IV U2538 ( .A(b[155]), .Z(n846) );
  NOR U2539 ( .A(n1466), .B(n846), .Z(n1468) );
  IV U2540 ( .A(a[154]), .Z(n1463) );
  IV U2541 ( .A(b[154]), .Z(n847) );
  NOR U2542 ( .A(n1463), .B(n847), .Z(n1465) );
  IV U2543 ( .A(a[153]), .Z(n1460) );
  IV U2544 ( .A(b[153]), .Z(n848) );
  NOR U2545 ( .A(n1460), .B(n848), .Z(n1462) );
  IV U2546 ( .A(a[152]), .Z(n1457) );
  IV U2547 ( .A(b[152]), .Z(n849) );
  NOR U2548 ( .A(n1457), .B(n849), .Z(n1459) );
  IV U2549 ( .A(a[151]), .Z(n1454) );
  IV U2550 ( .A(b[151]), .Z(n850) );
  NOR U2551 ( .A(n1454), .B(n850), .Z(n1456) );
  IV U2552 ( .A(a[150]), .Z(n1451) );
  IV U2553 ( .A(b[150]), .Z(n851) );
  NOR U2554 ( .A(n1451), .B(n851), .Z(n1453) );
  IV U2555 ( .A(a[149]), .Z(n1448) );
  IV U2556 ( .A(b[149]), .Z(n852) );
  NOR U2557 ( .A(n1448), .B(n852), .Z(n1450) );
  IV U2558 ( .A(a[148]), .Z(n1445) );
  IV U2559 ( .A(b[148]), .Z(n853) );
  NOR U2560 ( .A(n1445), .B(n853), .Z(n1447) );
  IV U2561 ( .A(a[147]), .Z(n1442) );
  IV U2562 ( .A(b[147]), .Z(n854) );
  NOR U2563 ( .A(n1442), .B(n854), .Z(n1444) );
  IV U2564 ( .A(a[146]), .Z(n1439) );
  IV U2565 ( .A(b[146]), .Z(n855) );
  NOR U2566 ( .A(n1439), .B(n855), .Z(n1441) );
  IV U2567 ( .A(a[145]), .Z(n1436) );
  IV U2568 ( .A(b[145]), .Z(n856) );
  NOR U2569 ( .A(n1436), .B(n856), .Z(n1438) );
  IV U2570 ( .A(a[144]), .Z(n1433) );
  IV U2571 ( .A(b[144]), .Z(n857) );
  NOR U2572 ( .A(n1433), .B(n857), .Z(n1435) );
  IV U2573 ( .A(a[143]), .Z(n1430) );
  IV U2574 ( .A(b[143]), .Z(n858) );
  NOR U2575 ( .A(n1430), .B(n858), .Z(n1432) );
  IV U2576 ( .A(a[142]), .Z(n1427) );
  IV U2577 ( .A(b[142]), .Z(n859) );
  NOR U2578 ( .A(n1427), .B(n859), .Z(n1429) );
  IV U2579 ( .A(a[141]), .Z(n1424) );
  IV U2580 ( .A(b[141]), .Z(n860) );
  NOR U2581 ( .A(n1424), .B(n860), .Z(n1426) );
  IV U2582 ( .A(a[140]), .Z(n1421) );
  IV U2583 ( .A(b[140]), .Z(n861) );
  NOR U2584 ( .A(n1421), .B(n861), .Z(n1423) );
  IV U2585 ( .A(a[139]), .Z(n1418) );
  IV U2586 ( .A(b[139]), .Z(n862) );
  NOR U2587 ( .A(n1418), .B(n862), .Z(n1420) );
  IV U2588 ( .A(a[138]), .Z(n1415) );
  IV U2589 ( .A(b[138]), .Z(n863) );
  NOR U2590 ( .A(n1415), .B(n863), .Z(n1417) );
  IV U2591 ( .A(a[137]), .Z(n1412) );
  IV U2592 ( .A(b[137]), .Z(n864) );
  NOR U2593 ( .A(n1412), .B(n864), .Z(n1414) );
  IV U2594 ( .A(a[136]), .Z(n1409) );
  IV U2595 ( .A(b[136]), .Z(n865) );
  NOR U2596 ( .A(n1409), .B(n865), .Z(n1411) );
  IV U2597 ( .A(a[135]), .Z(n1406) );
  IV U2598 ( .A(b[135]), .Z(n866) );
  NOR U2599 ( .A(n1406), .B(n866), .Z(n1408) );
  IV U2600 ( .A(a[134]), .Z(n1403) );
  IV U2601 ( .A(b[134]), .Z(n867) );
  NOR U2602 ( .A(n1403), .B(n867), .Z(n1405) );
  IV U2603 ( .A(a[133]), .Z(n1400) );
  IV U2604 ( .A(b[133]), .Z(n868) );
  NOR U2605 ( .A(n1400), .B(n868), .Z(n1402) );
  IV U2606 ( .A(a[132]), .Z(n1397) );
  IV U2607 ( .A(b[132]), .Z(n869) );
  NOR U2608 ( .A(n1397), .B(n869), .Z(n1399) );
  IV U2609 ( .A(a[131]), .Z(n1394) );
  IV U2610 ( .A(b[131]), .Z(n870) );
  NOR U2611 ( .A(n1394), .B(n870), .Z(n1396) );
  IV U2612 ( .A(a[130]), .Z(n1391) );
  IV U2613 ( .A(b[130]), .Z(n871) );
  NOR U2614 ( .A(n1391), .B(n871), .Z(n1393) );
  IV U2615 ( .A(a[129]), .Z(n1388) );
  IV U2616 ( .A(b[129]), .Z(n872) );
  NOR U2617 ( .A(n1388), .B(n872), .Z(n1390) );
  IV U2618 ( .A(a[128]), .Z(n1385) );
  IV U2619 ( .A(b[128]), .Z(n873) );
  NOR U2620 ( .A(n1385), .B(n873), .Z(n1387) );
  IV U2621 ( .A(a[127]), .Z(n1382) );
  IV U2622 ( .A(b[127]), .Z(n874) );
  NOR U2623 ( .A(n1382), .B(n874), .Z(n1384) );
  IV U2624 ( .A(a[126]), .Z(n1379) );
  IV U2625 ( .A(b[126]), .Z(n875) );
  NOR U2626 ( .A(n1379), .B(n875), .Z(n1381) );
  IV U2627 ( .A(a[125]), .Z(n1376) );
  IV U2628 ( .A(b[125]), .Z(n876) );
  NOR U2629 ( .A(n1376), .B(n876), .Z(n1378) );
  IV U2630 ( .A(a[124]), .Z(n1373) );
  IV U2631 ( .A(b[124]), .Z(n877) );
  NOR U2632 ( .A(n1373), .B(n877), .Z(n1375) );
  IV U2633 ( .A(a[123]), .Z(n1370) );
  IV U2634 ( .A(b[123]), .Z(n878) );
  NOR U2635 ( .A(n1370), .B(n878), .Z(n1372) );
  IV U2636 ( .A(a[122]), .Z(n1367) );
  IV U2637 ( .A(b[122]), .Z(n879) );
  NOR U2638 ( .A(n1367), .B(n879), .Z(n1369) );
  IV U2639 ( .A(a[121]), .Z(n1364) );
  IV U2640 ( .A(b[121]), .Z(n880) );
  NOR U2641 ( .A(n1364), .B(n880), .Z(n1366) );
  IV U2642 ( .A(a[120]), .Z(n1361) );
  IV U2643 ( .A(b[120]), .Z(n881) );
  NOR U2644 ( .A(n1361), .B(n881), .Z(n1363) );
  IV U2645 ( .A(a[119]), .Z(n1358) );
  IV U2646 ( .A(b[119]), .Z(n882) );
  NOR U2647 ( .A(n1358), .B(n882), .Z(n1360) );
  IV U2648 ( .A(a[118]), .Z(n1355) );
  IV U2649 ( .A(b[118]), .Z(n883) );
  NOR U2650 ( .A(n1355), .B(n883), .Z(n1357) );
  IV U2651 ( .A(a[117]), .Z(n1352) );
  IV U2652 ( .A(b[117]), .Z(n884) );
  NOR U2653 ( .A(n1352), .B(n884), .Z(n1354) );
  IV U2654 ( .A(a[116]), .Z(n1349) );
  IV U2655 ( .A(b[116]), .Z(n885) );
  NOR U2656 ( .A(n1349), .B(n885), .Z(n1351) );
  IV U2657 ( .A(a[115]), .Z(n1346) );
  IV U2658 ( .A(b[115]), .Z(n886) );
  NOR U2659 ( .A(n1346), .B(n886), .Z(n1348) );
  IV U2660 ( .A(a[114]), .Z(n1343) );
  IV U2661 ( .A(b[114]), .Z(n887) );
  NOR U2662 ( .A(n1343), .B(n887), .Z(n1345) );
  IV U2663 ( .A(a[113]), .Z(n1340) );
  IV U2664 ( .A(b[113]), .Z(n888) );
  NOR U2665 ( .A(n1340), .B(n888), .Z(n1342) );
  IV U2666 ( .A(a[112]), .Z(n1337) );
  IV U2667 ( .A(b[112]), .Z(n889) );
  NOR U2668 ( .A(n1337), .B(n889), .Z(n1339) );
  IV U2669 ( .A(a[111]), .Z(n1334) );
  IV U2670 ( .A(b[111]), .Z(n890) );
  NOR U2671 ( .A(n1334), .B(n890), .Z(n1336) );
  IV U2672 ( .A(a[110]), .Z(n1331) );
  IV U2673 ( .A(b[110]), .Z(n891) );
  NOR U2674 ( .A(n1331), .B(n891), .Z(n1333) );
  IV U2675 ( .A(a[109]), .Z(n1328) );
  IV U2676 ( .A(b[109]), .Z(n892) );
  NOR U2677 ( .A(n1328), .B(n892), .Z(n1330) );
  IV U2678 ( .A(a[108]), .Z(n1325) );
  IV U2679 ( .A(b[108]), .Z(n893) );
  NOR U2680 ( .A(n1325), .B(n893), .Z(n1327) );
  IV U2681 ( .A(a[107]), .Z(n1322) );
  IV U2682 ( .A(b[107]), .Z(n894) );
  NOR U2683 ( .A(n1322), .B(n894), .Z(n1324) );
  IV U2684 ( .A(a[106]), .Z(n1319) );
  IV U2685 ( .A(b[106]), .Z(n895) );
  NOR U2686 ( .A(n1319), .B(n895), .Z(n1321) );
  IV U2687 ( .A(a[105]), .Z(n1316) );
  IV U2688 ( .A(b[105]), .Z(n896) );
  NOR U2689 ( .A(n1316), .B(n896), .Z(n1318) );
  IV U2690 ( .A(a[104]), .Z(n1313) );
  IV U2691 ( .A(b[104]), .Z(n897) );
  NOR U2692 ( .A(n1313), .B(n897), .Z(n1315) );
  IV U2693 ( .A(a[103]), .Z(n1310) );
  IV U2694 ( .A(b[103]), .Z(n898) );
  NOR U2695 ( .A(n1310), .B(n898), .Z(n1312) );
  IV U2696 ( .A(a[102]), .Z(n1307) );
  IV U2697 ( .A(b[102]), .Z(n899) );
  NOR U2698 ( .A(n1307), .B(n899), .Z(n1309) );
  IV U2699 ( .A(a[101]), .Z(n1304) );
  IV U2700 ( .A(b[101]), .Z(n900) );
  NOR U2701 ( .A(n1304), .B(n900), .Z(n1306) );
  IV U2702 ( .A(a[100]), .Z(n1301) );
  IV U2703 ( .A(b[100]), .Z(n901) );
  NOR U2704 ( .A(n1301), .B(n901), .Z(n1303) );
  IV U2705 ( .A(b[99]), .Z(n1298) );
  IV U2706 ( .A(a[99]), .Z(n902) );
  NOR U2707 ( .A(n1298), .B(n902), .Z(n1300) );
  IV U2708 ( .A(a[98]), .Z(n1295) );
  IV U2709 ( .A(b[98]), .Z(n903) );
  NOR U2710 ( .A(n1295), .B(n903), .Z(n1297) );
  IV U2711 ( .A(a[97]), .Z(n1292) );
  IV U2712 ( .A(b[97]), .Z(n904) );
  NOR U2713 ( .A(n1292), .B(n904), .Z(n1294) );
  IV U2714 ( .A(a[96]), .Z(n1289) );
  IV U2715 ( .A(b[96]), .Z(n905) );
  NOR U2716 ( .A(n1289), .B(n905), .Z(n1291) );
  IV U2717 ( .A(a[95]), .Z(n1286) );
  IV U2718 ( .A(b[95]), .Z(n906) );
  NOR U2719 ( .A(n1286), .B(n906), .Z(n1288) );
  IV U2720 ( .A(a[94]), .Z(n1283) );
  IV U2721 ( .A(b[94]), .Z(n907) );
  NOR U2722 ( .A(n1283), .B(n907), .Z(n1285) );
  IV U2723 ( .A(a[93]), .Z(n1280) );
  IV U2724 ( .A(b[93]), .Z(n908) );
  NOR U2725 ( .A(n1280), .B(n908), .Z(n1282) );
  IV U2726 ( .A(a[92]), .Z(n1277) );
  IV U2727 ( .A(b[92]), .Z(n909) );
  NOR U2728 ( .A(n1277), .B(n909), .Z(n1279) );
  IV U2729 ( .A(a[91]), .Z(n1274) );
  IV U2730 ( .A(b[91]), .Z(n910) );
  NOR U2731 ( .A(n1274), .B(n910), .Z(n1276) );
  IV U2732 ( .A(a[90]), .Z(n1271) );
  IV U2733 ( .A(b[90]), .Z(n911) );
  NOR U2734 ( .A(n1271), .B(n911), .Z(n1273) );
  IV U2735 ( .A(a[89]), .Z(n1268) );
  IV U2736 ( .A(b[89]), .Z(n912) );
  NOR U2737 ( .A(n1268), .B(n912), .Z(n1270) );
  IV U2738 ( .A(a[88]), .Z(n1265) );
  IV U2739 ( .A(b[88]), .Z(n913) );
  NOR U2740 ( .A(n1265), .B(n913), .Z(n1267) );
  IV U2741 ( .A(a[87]), .Z(n1262) );
  IV U2742 ( .A(b[87]), .Z(n914) );
  NOR U2743 ( .A(n1262), .B(n914), .Z(n1264) );
  IV U2744 ( .A(a[86]), .Z(n1259) );
  IV U2745 ( .A(b[86]), .Z(n915) );
  NOR U2746 ( .A(n1259), .B(n915), .Z(n1261) );
  IV U2747 ( .A(a[85]), .Z(n1256) );
  IV U2748 ( .A(b[85]), .Z(n916) );
  NOR U2749 ( .A(n1256), .B(n916), .Z(n1258) );
  IV U2750 ( .A(a[84]), .Z(n1253) );
  IV U2751 ( .A(b[84]), .Z(n917) );
  NOR U2752 ( .A(n1253), .B(n917), .Z(n1255) );
  IV U2753 ( .A(a[83]), .Z(n1250) );
  IV U2754 ( .A(b[83]), .Z(n918) );
  NOR U2755 ( .A(n1250), .B(n918), .Z(n1252) );
  IV U2756 ( .A(a[82]), .Z(n1247) );
  IV U2757 ( .A(b[82]), .Z(n919) );
  NOR U2758 ( .A(n1247), .B(n919), .Z(n1249) );
  IV U2759 ( .A(a[81]), .Z(n1244) );
  IV U2760 ( .A(b[81]), .Z(n920) );
  NOR U2761 ( .A(n1244), .B(n920), .Z(n1246) );
  IV U2762 ( .A(a[80]), .Z(n1241) );
  IV U2763 ( .A(b[80]), .Z(n921) );
  NOR U2764 ( .A(n1241), .B(n921), .Z(n1243) );
  IV U2765 ( .A(a[79]), .Z(n1238) );
  IV U2766 ( .A(b[79]), .Z(n922) );
  NOR U2767 ( .A(n1238), .B(n922), .Z(n1240) );
  IV U2768 ( .A(a[78]), .Z(n1235) );
  IV U2769 ( .A(b[78]), .Z(n923) );
  NOR U2770 ( .A(n1235), .B(n923), .Z(n1237) );
  IV U2771 ( .A(a[77]), .Z(n1232) );
  IV U2772 ( .A(b[77]), .Z(n924) );
  NOR U2773 ( .A(n1232), .B(n924), .Z(n1234) );
  IV U2774 ( .A(a[76]), .Z(n1229) );
  IV U2775 ( .A(b[76]), .Z(n925) );
  NOR U2776 ( .A(n1229), .B(n925), .Z(n1231) );
  IV U2777 ( .A(a[75]), .Z(n1226) );
  IV U2778 ( .A(b[75]), .Z(n926) );
  NOR U2779 ( .A(n1226), .B(n926), .Z(n1228) );
  IV U2780 ( .A(a[74]), .Z(n1223) );
  IV U2781 ( .A(b[74]), .Z(n927) );
  NOR U2782 ( .A(n1223), .B(n927), .Z(n1225) );
  IV U2783 ( .A(a[73]), .Z(n1220) );
  IV U2784 ( .A(b[73]), .Z(n928) );
  NOR U2785 ( .A(n1220), .B(n928), .Z(n1222) );
  IV U2786 ( .A(a[72]), .Z(n1217) );
  IV U2787 ( .A(b[72]), .Z(n929) );
  NOR U2788 ( .A(n1217), .B(n929), .Z(n1219) );
  IV U2789 ( .A(a[71]), .Z(n1214) );
  IV U2790 ( .A(b[71]), .Z(n930) );
  NOR U2791 ( .A(n1214), .B(n930), .Z(n1216) );
  IV U2792 ( .A(a[70]), .Z(n1211) );
  IV U2793 ( .A(b[70]), .Z(n931) );
  NOR U2794 ( .A(n1211), .B(n931), .Z(n1213) );
  IV U2795 ( .A(a[69]), .Z(n1208) );
  IV U2796 ( .A(b[69]), .Z(n932) );
  NOR U2797 ( .A(n1208), .B(n932), .Z(n1210) );
  IV U2798 ( .A(a[68]), .Z(n1205) );
  IV U2799 ( .A(b[68]), .Z(n933) );
  NOR U2800 ( .A(n1205), .B(n933), .Z(n1207) );
  IV U2801 ( .A(a[67]), .Z(n1202) );
  IV U2802 ( .A(b[67]), .Z(n934) );
  NOR U2803 ( .A(n1202), .B(n934), .Z(n1204) );
  IV U2804 ( .A(a[66]), .Z(n1199) );
  IV U2805 ( .A(b[66]), .Z(n935) );
  NOR U2806 ( .A(n1199), .B(n935), .Z(n1201) );
  IV U2807 ( .A(a[65]), .Z(n1196) );
  IV U2808 ( .A(b[65]), .Z(n936) );
  NOR U2809 ( .A(n1196), .B(n936), .Z(n1198) );
  IV U2810 ( .A(a[64]), .Z(n1193) );
  IV U2811 ( .A(b[64]), .Z(n937) );
  NOR U2812 ( .A(n1193), .B(n937), .Z(n1195) );
  IV U2813 ( .A(a[63]), .Z(n1190) );
  IV U2814 ( .A(b[63]), .Z(n938) );
  NOR U2815 ( .A(n1190), .B(n938), .Z(n1192) );
  IV U2816 ( .A(a[62]), .Z(n1187) );
  IV U2817 ( .A(b[62]), .Z(n939) );
  NOR U2818 ( .A(n1187), .B(n939), .Z(n1189) );
  IV U2819 ( .A(a[61]), .Z(n1184) );
  IV U2820 ( .A(b[61]), .Z(n940) );
  NOR U2821 ( .A(n1184), .B(n940), .Z(n1186) );
  IV U2822 ( .A(a[60]), .Z(n1181) );
  IV U2823 ( .A(b[60]), .Z(n941) );
  NOR U2824 ( .A(n1181), .B(n941), .Z(n1183) );
  IV U2825 ( .A(a[59]), .Z(n1178) );
  IV U2826 ( .A(b[59]), .Z(n942) );
  NOR U2827 ( .A(n1178), .B(n942), .Z(n1180) );
  IV U2828 ( .A(a[58]), .Z(n1175) );
  IV U2829 ( .A(b[58]), .Z(n943) );
  NOR U2830 ( .A(n1175), .B(n943), .Z(n1177) );
  IV U2831 ( .A(a[57]), .Z(n1172) );
  IV U2832 ( .A(b[57]), .Z(n944) );
  NOR U2833 ( .A(n1172), .B(n944), .Z(n1174) );
  IV U2834 ( .A(a[56]), .Z(n1169) );
  IV U2835 ( .A(b[56]), .Z(n945) );
  NOR U2836 ( .A(n1169), .B(n945), .Z(n1171) );
  IV U2837 ( .A(a[55]), .Z(n1166) );
  IV U2838 ( .A(b[55]), .Z(n946) );
  NOR U2839 ( .A(n1166), .B(n946), .Z(n1168) );
  IV U2840 ( .A(a[54]), .Z(n1163) );
  IV U2841 ( .A(b[54]), .Z(n947) );
  NOR U2842 ( .A(n1163), .B(n947), .Z(n1165) );
  IV U2843 ( .A(a[53]), .Z(n1160) );
  IV U2844 ( .A(b[53]), .Z(n948) );
  NOR U2845 ( .A(n1160), .B(n948), .Z(n1162) );
  IV U2846 ( .A(a[52]), .Z(n1157) );
  IV U2847 ( .A(b[52]), .Z(n949) );
  NOR U2848 ( .A(n1157), .B(n949), .Z(n1159) );
  IV U2849 ( .A(a[51]), .Z(n1154) );
  IV U2850 ( .A(b[51]), .Z(n950) );
  NOR U2851 ( .A(n1154), .B(n950), .Z(n1156) );
  IV U2852 ( .A(a[50]), .Z(n1151) );
  IV U2853 ( .A(b[50]), .Z(n951) );
  NOR U2854 ( .A(n1151), .B(n951), .Z(n1153) );
  IV U2855 ( .A(a[49]), .Z(n1148) );
  IV U2856 ( .A(b[49]), .Z(n952) );
  NOR U2857 ( .A(n1148), .B(n952), .Z(n1150) );
  IV U2858 ( .A(a[48]), .Z(n1145) );
  IV U2859 ( .A(b[48]), .Z(n953) );
  NOR U2860 ( .A(n1145), .B(n953), .Z(n1147) );
  IV U2861 ( .A(a[47]), .Z(n1142) );
  IV U2862 ( .A(b[47]), .Z(n954) );
  NOR U2863 ( .A(n1142), .B(n954), .Z(n1144) );
  IV U2864 ( .A(a[46]), .Z(n1139) );
  IV U2865 ( .A(b[46]), .Z(n955) );
  NOR U2866 ( .A(n1139), .B(n955), .Z(n1141) );
  IV U2867 ( .A(a[45]), .Z(n1136) );
  IV U2868 ( .A(b[45]), .Z(n956) );
  NOR U2869 ( .A(n1136), .B(n956), .Z(n1138) );
  IV U2870 ( .A(a[44]), .Z(n1133) );
  IV U2871 ( .A(b[44]), .Z(n957) );
  NOR U2872 ( .A(n1133), .B(n957), .Z(n1135) );
  IV U2873 ( .A(a[43]), .Z(n1130) );
  IV U2874 ( .A(b[43]), .Z(n958) );
  NOR U2875 ( .A(n1130), .B(n958), .Z(n1132) );
  IV U2876 ( .A(a[42]), .Z(n1127) );
  IV U2877 ( .A(b[42]), .Z(n959) );
  NOR U2878 ( .A(n1127), .B(n959), .Z(n1129) );
  IV U2879 ( .A(a[41]), .Z(n1124) );
  IV U2880 ( .A(b[41]), .Z(n960) );
  NOR U2881 ( .A(n1124), .B(n960), .Z(n1126) );
  IV U2882 ( .A(a[40]), .Z(n1121) );
  IV U2883 ( .A(b[40]), .Z(n961) );
  NOR U2884 ( .A(n1121), .B(n961), .Z(n1123) );
  IV U2885 ( .A(a[39]), .Z(n1118) );
  IV U2886 ( .A(b[39]), .Z(n962) );
  NOR U2887 ( .A(n1118), .B(n962), .Z(n1120) );
  IV U2888 ( .A(a[38]), .Z(n1115) );
  IV U2889 ( .A(b[38]), .Z(n963) );
  NOR U2890 ( .A(n1115), .B(n963), .Z(n1117) );
  IV U2891 ( .A(a[37]), .Z(n1112) );
  IV U2892 ( .A(b[37]), .Z(n964) );
  NOR U2893 ( .A(n1112), .B(n964), .Z(n1114) );
  IV U2894 ( .A(a[36]), .Z(n1109) );
  IV U2895 ( .A(b[36]), .Z(n965) );
  NOR U2896 ( .A(n1109), .B(n965), .Z(n1111) );
  IV U2897 ( .A(a[35]), .Z(n1106) );
  IV U2898 ( .A(b[35]), .Z(n966) );
  NOR U2899 ( .A(n1106), .B(n966), .Z(n1108) );
  IV U2900 ( .A(a[34]), .Z(n1103) );
  IV U2901 ( .A(b[34]), .Z(n967) );
  NOR U2902 ( .A(n1103), .B(n967), .Z(n1105) );
  IV U2903 ( .A(a[33]), .Z(n1100) );
  IV U2904 ( .A(b[33]), .Z(n968) );
  NOR U2905 ( .A(n1100), .B(n968), .Z(n1102) );
  IV U2906 ( .A(a[32]), .Z(n1097) );
  IV U2907 ( .A(b[32]), .Z(n969) );
  NOR U2908 ( .A(n1097), .B(n969), .Z(n1099) );
  IV U2909 ( .A(a[31]), .Z(n1094) );
  IV U2910 ( .A(b[31]), .Z(n970) );
  NOR U2911 ( .A(n1094), .B(n970), .Z(n1096) );
  IV U2912 ( .A(a[30]), .Z(n1091) );
  IV U2913 ( .A(b[30]), .Z(n971) );
  NOR U2914 ( .A(n1091), .B(n971), .Z(n1093) );
  IV U2915 ( .A(a[29]), .Z(n1088) );
  IV U2916 ( .A(b[29]), .Z(n972) );
  NOR U2917 ( .A(n1088), .B(n972), .Z(n1090) );
  IV U2918 ( .A(a[28]), .Z(n1085) );
  IV U2919 ( .A(b[28]), .Z(n973) );
  NOR U2920 ( .A(n1085), .B(n973), .Z(n1087) );
  IV U2921 ( .A(a[27]), .Z(n1082) );
  IV U2922 ( .A(b[27]), .Z(n974) );
  NOR U2923 ( .A(n1082), .B(n974), .Z(n1084) );
  IV U2924 ( .A(a[26]), .Z(n1079) );
  IV U2925 ( .A(b[26]), .Z(n975) );
  NOR U2926 ( .A(n1079), .B(n975), .Z(n1081) );
  IV U2927 ( .A(a[25]), .Z(n1076) );
  IV U2928 ( .A(b[25]), .Z(n976) );
  NOR U2929 ( .A(n1076), .B(n976), .Z(n1078) );
  IV U2930 ( .A(a[24]), .Z(n1073) );
  IV U2931 ( .A(b[24]), .Z(n977) );
  NOR U2932 ( .A(n1073), .B(n977), .Z(n1075) );
  IV U2933 ( .A(a[23]), .Z(n1070) );
  IV U2934 ( .A(b[23]), .Z(n978) );
  NOR U2935 ( .A(n1070), .B(n978), .Z(n1072) );
  IV U2936 ( .A(a[22]), .Z(n1067) );
  IV U2937 ( .A(b[22]), .Z(n979) );
  NOR U2938 ( .A(n1067), .B(n979), .Z(n1069) );
  IV U2939 ( .A(a[21]), .Z(n1064) );
  IV U2940 ( .A(b[21]), .Z(n980) );
  NOR U2941 ( .A(n1064), .B(n980), .Z(n1066) );
  IV U2942 ( .A(a[20]), .Z(n1061) );
  IV U2943 ( .A(b[20]), .Z(n981) );
  NOR U2944 ( .A(n1061), .B(n981), .Z(n1063) );
  IV U2945 ( .A(a[19]), .Z(n1058) );
  IV U2946 ( .A(b[19]), .Z(n982) );
  NOR U2947 ( .A(n1058), .B(n982), .Z(n1060) );
  IV U2948 ( .A(a[18]), .Z(n1055) );
  IV U2949 ( .A(b[18]), .Z(n983) );
  NOR U2950 ( .A(n1055), .B(n983), .Z(n1057) );
  IV U2951 ( .A(a[17]), .Z(n1052) );
  IV U2952 ( .A(b[17]), .Z(n984) );
  NOR U2953 ( .A(n1052), .B(n984), .Z(n1054) );
  IV U2954 ( .A(a[16]), .Z(n1049) );
  IV U2955 ( .A(b[16]), .Z(n985) );
  NOR U2956 ( .A(n1049), .B(n985), .Z(n1051) );
  IV U2957 ( .A(a[15]), .Z(n1046) );
  IV U2958 ( .A(b[15]), .Z(n986) );
  NOR U2959 ( .A(n1046), .B(n986), .Z(n1048) );
  IV U2960 ( .A(a[14]), .Z(n1043) );
  IV U2961 ( .A(b[14]), .Z(n987) );
  NOR U2962 ( .A(n1043), .B(n987), .Z(n1045) );
  IV U2963 ( .A(a[13]), .Z(n1040) );
  IV U2964 ( .A(b[13]), .Z(n988) );
  NOR U2965 ( .A(n1040), .B(n988), .Z(n1042) );
  IV U2966 ( .A(a[12]), .Z(n1037) );
  IV U2967 ( .A(b[12]), .Z(n989) );
  NOR U2968 ( .A(n1037), .B(n989), .Z(n1039) );
  IV U2969 ( .A(a[11]), .Z(n1034) );
  IV U2970 ( .A(b[11]), .Z(n990) );
  NOR U2971 ( .A(n1034), .B(n990), .Z(n1036) );
  IV U2972 ( .A(a[10]), .Z(n1031) );
  IV U2973 ( .A(b[10]), .Z(n991) );
  NOR U2974 ( .A(n1031), .B(n991), .Z(n1033) );
  IV U2975 ( .A(b[9]), .Z(n1028) );
  IV U2976 ( .A(a[9]), .Z(n992) );
  NOR U2977 ( .A(n1028), .B(n992), .Z(n1030) );
  IV U2978 ( .A(a[8]), .Z(n1025) );
  IV U2979 ( .A(b[8]), .Z(n993) );
  NOR U2980 ( .A(n1025), .B(n993), .Z(n1027) );
  IV U2981 ( .A(a[7]), .Z(n1022) );
  IV U2982 ( .A(b[7]), .Z(n994) );
  NOR U2983 ( .A(n1022), .B(n994), .Z(n1024) );
  IV U2984 ( .A(a[6]), .Z(n1019) );
  IV U2985 ( .A(b[6]), .Z(n995) );
  NOR U2986 ( .A(n1019), .B(n995), .Z(n1021) );
  IV U2987 ( .A(a[5]), .Z(n1016) );
  IV U2988 ( .A(b[5]), .Z(n996) );
  NOR U2989 ( .A(n1016), .B(n996), .Z(n1018) );
  IV U2990 ( .A(a[4]), .Z(n1013) );
  IV U2991 ( .A(b[4]), .Z(n997) );
  NOR U2992 ( .A(n1013), .B(n997), .Z(n1015) );
  IV U2993 ( .A(a[3]), .Z(n1010) );
  IV U2994 ( .A(b[3]), .Z(n998) );
  NOR U2995 ( .A(n1010), .B(n998), .Z(n1012) );
  IV U2996 ( .A(a[2]), .Z(n1007) );
  IV U2997 ( .A(b[2]), .Z(n999) );
  NOR U2998 ( .A(n1007), .B(n999), .Z(n1009) );
  IV U2999 ( .A(a[1]), .Z(n1001) );
  IV U3000 ( .A(b[1]), .Z(n1000) );
  NOR U3001 ( .A(n1001), .B(n1000), .Z(n1006) );
  XOR U3002 ( .A(n1001), .B(b[1]), .Z(n4360) );
  NOR U3003 ( .A(n1003), .B(n1002), .Z(n1004) );
  IV U3004 ( .A(n1004), .Z(n4359) );
  NOR U3005 ( .A(n4360), .B(n4359), .Z(n1005) );
  NOR U3006 ( .A(n1006), .B(n1005), .Z(n4582) );
  XOR U3007 ( .A(n1007), .B(b[2]), .Z(n4581) );
  NOR U3008 ( .A(n4582), .B(n4581), .Z(n1008) );
  NOR U3009 ( .A(n1009), .B(n1008), .Z(n4804) );
  XOR U3010 ( .A(n1010), .B(b[3]), .Z(n4803) );
  NOR U3011 ( .A(n4804), .B(n4803), .Z(n1011) );
  NOR U3012 ( .A(n1012), .B(n1011), .Z(n5026) );
  XOR U3013 ( .A(n1013), .B(b[4]), .Z(n5025) );
  NOR U3014 ( .A(n5026), .B(n5025), .Z(n1014) );
  NOR U3015 ( .A(n1015), .B(n1014), .Z(n5248) );
  XOR U3016 ( .A(n1016), .B(b[5]), .Z(n5247) );
  NOR U3017 ( .A(n5248), .B(n5247), .Z(n1017) );
  NOR U3018 ( .A(n1018), .B(n1017), .Z(n5470) );
  XOR U3019 ( .A(n1019), .B(b[6]), .Z(n5469) );
  NOR U3020 ( .A(n5470), .B(n5469), .Z(n1020) );
  NOR U3021 ( .A(n1021), .B(n1020), .Z(n5692) );
  XOR U3022 ( .A(n1022), .B(b[7]), .Z(n5691) );
  NOR U3023 ( .A(n5692), .B(n5691), .Z(n1023) );
  NOR U3024 ( .A(n1024), .B(n1023), .Z(n5914) );
  XOR U3025 ( .A(n1025), .B(b[8]), .Z(n5913) );
  NOR U3026 ( .A(n5914), .B(n5913), .Z(n1026) );
  NOR U3027 ( .A(n1027), .B(n1026), .Z(n6136) );
  XOR U3028 ( .A(n1028), .B(a[9]), .Z(n6135) );
  NOR U3029 ( .A(n6136), .B(n6135), .Z(n1029) );
  NOR U3030 ( .A(n1030), .B(n1029), .Z(n4160) );
  XOR U3031 ( .A(n1031), .B(b[10]), .Z(n4159) );
  NOR U3032 ( .A(n4160), .B(n4159), .Z(n1032) );
  NOR U3033 ( .A(n1033), .B(n1032), .Z(n4182) );
  XOR U3034 ( .A(n1034), .B(b[11]), .Z(n4181) );
  NOR U3035 ( .A(n4182), .B(n4181), .Z(n1035) );
  NOR U3036 ( .A(n1036), .B(n1035), .Z(n4204) );
  XOR U3037 ( .A(n1037), .B(b[12]), .Z(n4203) );
  NOR U3038 ( .A(n4204), .B(n4203), .Z(n1038) );
  NOR U3039 ( .A(n1039), .B(n1038), .Z(n4226) );
  XOR U3040 ( .A(n1040), .B(b[13]), .Z(n4225) );
  NOR U3041 ( .A(n4226), .B(n4225), .Z(n1041) );
  NOR U3042 ( .A(n1042), .B(n1041), .Z(n4248) );
  XOR U3043 ( .A(n1043), .B(b[14]), .Z(n4247) );
  NOR U3044 ( .A(n4248), .B(n4247), .Z(n1044) );
  NOR U3045 ( .A(n1045), .B(n1044), .Z(n4270) );
  XOR U3046 ( .A(n1046), .B(b[15]), .Z(n4269) );
  NOR U3047 ( .A(n4270), .B(n4269), .Z(n1047) );
  NOR U3048 ( .A(n1048), .B(n1047), .Z(n4292) );
  XOR U3049 ( .A(n1049), .B(b[16]), .Z(n4291) );
  NOR U3050 ( .A(n4292), .B(n4291), .Z(n1050) );
  NOR U3051 ( .A(n1051), .B(n1050), .Z(n4314) );
  XOR U3052 ( .A(n1052), .B(b[17]), .Z(n4313) );
  NOR U3053 ( .A(n4314), .B(n4313), .Z(n1053) );
  NOR U3054 ( .A(n1054), .B(n1053), .Z(n4336) );
  XOR U3055 ( .A(n1055), .B(b[18]), .Z(n4335) );
  NOR U3056 ( .A(n4336), .B(n4335), .Z(n1056) );
  NOR U3057 ( .A(n1057), .B(n1056), .Z(n4358) );
  XOR U3058 ( .A(n1058), .B(b[19]), .Z(n4357) );
  NOR U3059 ( .A(n4358), .B(n4357), .Z(n1059) );
  NOR U3060 ( .A(n1060), .B(n1059), .Z(n4382) );
  XOR U3061 ( .A(n1061), .B(b[20]), .Z(n4381) );
  NOR U3062 ( .A(n4382), .B(n4381), .Z(n1062) );
  NOR U3063 ( .A(n1063), .B(n1062), .Z(n4404) );
  XOR U3064 ( .A(n1064), .B(b[21]), .Z(n4403) );
  NOR U3065 ( .A(n4404), .B(n4403), .Z(n1065) );
  NOR U3066 ( .A(n1066), .B(n1065), .Z(n4426) );
  XOR U3067 ( .A(n1067), .B(b[22]), .Z(n4425) );
  NOR U3068 ( .A(n4426), .B(n4425), .Z(n1068) );
  NOR U3069 ( .A(n1069), .B(n1068), .Z(n4448) );
  XOR U3070 ( .A(n1070), .B(b[23]), .Z(n4447) );
  NOR U3071 ( .A(n4448), .B(n4447), .Z(n1071) );
  NOR U3072 ( .A(n1072), .B(n1071), .Z(n4470) );
  XOR U3073 ( .A(n1073), .B(b[24]), .Z(n4469) );
  NOR U3074 ( .A(n4470), .B(n4469), .Z(n1074) );
  NOR U3075 ( .A(n1075), .B(n1074), .Z(n4492) );
  XOR U3076 ( .A(n1076), .B(b[25]), .Z(n4491) );
  NOR U3077 ( .A(n4492), .B(n4491), .Z(n1077) );
  NOR U3078 ( .A(n1078), .B(n1077), .Z(n4514) );
  XOR U3079 ( .A(n1079), .B(b[26]), .Z(n4513) );
  NOR U3080 ( .A(n4514), .B(n4513), .Z(n1080) );
  NOR U3081 ( .A(n1081), .B(n1080), .Z(n4536) );
  XOR U3082 ( .A(n1082), .B(b[27]), .Z(n4535) );
  NOR U3083 ( .A(n4536), .B(n4535), .Z(n1083) );
  NOR U3084 ( .A(n1084), .B(n1083), .Z(n4558) );
  XOR U3085 ( .A(n1085), .B(b[28]), .Z(n4557) );
  NOR U3086 ( .A(n4558), .B(n4557), .Z(n1086) );
  NOR U3087 ( .A(n1087), .B(n1086), .Z(n4580) );
  XOR U3088 ( .A(n1088), .B(b[29]), .Z(n4579) );
  NOR U3089 ( .A(n4580), .B(n4579), .Z(n1089) );
  NOR U3090 ( .A(n1090), .B(n1089), .Z(n4604) );
  XOR U3091 ( .A(n1091), .B(b[30]), .Z(n4603) );
  NOR U3092 ( .A(n4604), .B(n4603), .Z(n1092) );
  NOR U3093 ( .A(n1093), .B(n1092), .Z(n4626) );
  XOR U3094 ( .A(n1094), .B(b[31]), .Z(n4625) );
  NOR U3095 ( .A(n4626), .B(n4625), .Z(n1095) );
  NOR U3096 ( .A(n1096), .B(n1095), .Z(n4648) );
  XOR U3097 ( .A(n1097), .B(b[32]), .Z(n4647) );
  NOR U3098 ( .A(n4648), .B(n4647), .Z(n1098) );
  NOR U3099 ( .A(n1099), .B(n1098), .Z(n4670) );
  XOR U3100 ( .A(n1100), .B(b[33]), .Z(n4669) );
  NOR U3101 ( .A(n4670), .B(n4669), .Z(n1101) );
  NOR U3102 ( .A(n1102), .B(n1101), .Z(n4692) );
  XOR U3103 ( .A(n1103), .B(b[34]), .Z(n4691) );
  NOR U3104 ( .A(n4692), .B(n4691), .Z(n1104) );
  NOR U3105 ( .A(n1105), .B(n1104), .Z(n4714) );
  XOR U3106 ( .A(n1106), .B(b[35]), .Z(n4713) );
  NOR U3107 ( .A(n4714), .B(n4713), .Z(n1107) );
  NOR U3108 ( .A(n1108), .B(n1107), .Z(n4736) );
  XOR U3109 ( .A(n1109), .B(b[36]), .Z(n4735) );
  NOR U3110 ( .A(n4736), .B(n4735), .Z(n1110) );
  NOR U3111 ( .A(n1111), .B(n1110), .Z(n4758) );
  XOR U3112 ( .A(n1112), .B(b[37]), .Z(n4757) );
  NOR U3113 ( .A(n4758), .B(n4757), .Z(n1113) );
  NOR U3114 ( .A(n1114), .B(n1113), .Z(n4780) );
  XOR U3115 ( .A(n1115), .B(b[38]), .Z(n4779) );
  NOR U3116 ( .A(n4780), .B(n4779), .Z(n1116) );
  NOR U3117 ( .A(n1117), .B(n1116), .Z(n4802) );
  XOR U3118 ( .A(n1118), .B(b[39]), .Z(n4801) );
  NOR U3119 ( .A(n4802), .B(n4801), .Z(n1119) );
  NOR U3120 ( .A(n1120), .B(n1119), .Z(n4826) );
  XOR U3121 ( .A(n1121), .B(b[40]), .Z(n4825) );
  NOR U3122 ( .A(n4826), .B(n4825), .Z(n1122) );
  NOR U3123 ( .A(n1123), .B(n1122), .Z(n4848) );
  XOR U3124 ( .A(n1124), .B(b[41]), .Z(n4847) );
  NOR U3125 ( .A(n4848), .B(n4847), .Z(n1125) );
  NOR U3126 ( .A(n1126), .B(n1125), .Z(n4870) );
  XOR U3127 ( .A(n1127), .B(b[42]), .Z(n4869) );
  NOR U3128 ( .A(n4870), .B(n4869), .Z(n1128) );
  NOR U3129 ( .A(n1129), .B(n1128), .Z(n4892) );
  XOR U3130 ( .A(n1130), .B(b[43]), .Z(n4891) );
  NOR U3131 ( .A(n4892), .B(n4891), .Z(n1131) );
  NOR U3132 ( .A(n1132), .B(n1131), .Z(n4914) );
  XOR U3133 ( .A(n1133), .B(b[44]), .Z(n4913) );
  NOR U3134 ( .A(n4914), .B(n4913), .Z(n1134) );
  NOR U3135 ( .A(n1135), .B(n1134), .Z(n4936) );
  XOR U3136 ( .A(n1136), .B(b[45]), .Z(n4935) );
  NOR U3137 ( .A(n4936), .B(n4935), .Z(n1137) );
  NOR U3138 ( .A(n1138), .B(n1137), .Z(n4958) );
  XOR U3139 ( .A(n1139), .B(b[46]), .Z(n4957) );
  NOR U3140 ( .A(n4958), .B(n4957), .Z(n1140) );
  NOR U3141 ( .A(n1141), .B(n1140), .Z(n4980) );
  XOR U3142 ( .A(n1142), .B(b[47]), .Z(n4979) );
  NOR U3143 ( .A(n4980), .B(n4979), .Z(n1143) );
  NOR U3144 ( .A(n1144), .B(n1143), .Z(n5002) );
  XOR U3145 ( .A(n1145), .B(b[48]), .Z(n5001) );
  NOR U3146 ( .A(n5002), .B(n5001), .Z(n1146) );
  NOR U3147 ( .A(n1147), .B(n1146), .Z(n5024) );
  XOR U3148 ( .A(n1148), .B(b[49]), .Z(n5023) );
  NOR U3149 ( .A(n5024), .B(n5023), .Z(n1149) );
  NOR U3150 ( .A(n1150), .B(n1149), .Z(n5048) );
  XOR U3151 ( .A(n1151), .B(b[50]), .Z(n5047) );
  NOR U3152 ( .A(n5048), .B(n5047), .Z(n1152) );
  NOR U3153 ( .A(n1153), .B(n1152), .Z(n5070) );
  XOR U3154 ( .A(n1154), .B(b[51]), .Z(n5069) );
  NOR U3155 ( .A(n5070), .B(n5069), .Z(n1155) );
  NOR U3156 ( .A(n1156), .B(n1155), .Z(n5092) );
  XOR U3157 ( .A(n1157), .B(b[52]), .Z(n5091) );
  NOR U3158 ( .A(n5092), .B(n5091), .Z(n1158) );
  NOR U3159 ( .A(n1159), .B(n1158), .Z(n5114) );
  XOR U3160 ( .A(n1160), .B(b[53]), .Z(n5113) );
  NOR U3161 ( .A(n5114), .B(n5113), .Z(n1161) );
  NOR U3162 ( .A(n1162), .B(n1161), .Z(n5136) );
  XOR U3163 ( .A(n1163), .B(b[54]), .Z(n5135) );
  NOR U3164 ( .A(n5136), .B(n5135), .Z(n1164) );
  NOR U3165 ( .A(n1165), .B(n1164), .Z(n5158) );
  XOR U3166 ( .A(n1166), .B(b[55]), .Z(n5157) );
  NOR U3167 ( .A(n5158), .B(n5157), .Z(n1167) );
  NOR U3168 ( .A(n1168), .B(n1167), .Z(n5180) );
  XOR U3169 ( .A(n1169), .B(b[56]), .Z(n5179) );
  NOR U3170 ( .A(n5180), .B(n5179), .Z(n1170) );
  NOR U3171 ( .A(n1171), .B(n1170), .Z(n5202) );
  XOR U3172 ( .A(n1172), .B(b[57]), .Z(n5201) );
  NOR U3173 ( .A(n5202), .B(n5201), .Z(n1173) );
  NOR U3174 ( .A(n1174), .B(n1173), .Z(n5224) );
  XOR U3175 ( .A(n1175), .B(b[58]), .Z(n5223) );
  NOR U3176 ( .A(n5224), .B(n5223), .Z(n1176) );
  NOR U3177 ( .A(n1177), .B(n1176), .Z(n5246) );
  XOR U3178 ( .A(n1178), .B(b[59]), .Z(n5245) );
  NOR U3179 ( .A(n5246), .B(n5245), .Z(n1179) );
  NOR U3180 ( .A(n1180), .B(n1179), .Z(n5270) );
  XOR U3181 ( .A(n1181), .B(b[60]), .Z(n5269) );
  NOR U3182 ( .A(n5270), .B(n5269), .Z(n1182) );
  NOR U3183 ( .A(n1183), .B(n1182), .Z(n5292) );
  XOR U3184 ( .A(n1184), .B(b[61]), .Z(n5291) );
  NOR U3185 ( .A(n5292), .B(n5291), .Z(n1185) );
  NOR U3186 ( .A(n1186), .B(n1185), .Z(n5314) );
  XOR U3187 ( .A(n1187), .B(b[62]), .Z(n5313) );
  NOR U3188 ( .A(n5314), .B(n5313), .Z(n1188) );
  NOR U3189 ( .A(n1189), .B(n1188), .Z(n5336) );
  XOR U3190 ( .A(n1190), .B(b[63]), .Z(n5335) );
  NOR U3191 ( .A(n5336), .B(n5335), .Z(n1191) );
  NOR U3192 ( .A(n1192), .B(n1191), .Z(n5358) );
  XOR U3193 ( .A(n1193), .B(b[64]), .Z(n5357) );
  NOR U3194 ( .A(n5358), .B(n5357), .Z(n1194) );
  NOR U3195 ( .A(n1195), .B(n1194), .Z(n5380) );
  XOR U3196 ( .A(n1196), .B(b[65]), .Z(n5379) );
  NOR U3197 ( .A(n5380), .B(n5379), .Z(n1197) );
  NOR U3198 ( .A(n1198), .B(n1197), .Z(n5402) );
  XOR U3199 ( .A(n1199), .B(b[66]), .Z(n5401) );
  NOR U3200 ( .A(n5402), .B(n5401), .Z(n1200) );
  NOR U3201 ( .A(n1201), .B(n1200), .Z(n5424) );
  XOR U3202 ( .A(n1202), .B(b[67]), .Z(n5423) );
  NOR U3203 ( .A(n5424), .B(n5423), .Z(n1203) );
  NOR U3204 ( .A(n1204), .B(n1203), .Z(n5446) );
  XOR U3205 ( .A(n1205), .B(b[68]), .Z(n5445) );
  NOR U3206 ( .A(n5446), .B(n5445), .Z(n1206) );
  NOR U3207 ( .A(n1207), .B(n1206), .Z(n5468) );
  XOR U3208 ( .A(n1208), .B(b[69]), .Z(n5467) );
  NOR U3209 ( .A(n5468), .B(n5467), .Z(n1209) );
  NOR U3210 ( .A(n1210), .B(n1209), .Z(n5492) );
  XOR U3211 ( .A(n1211), .B(b[70]), .Z(n5491) );
  NOR U3212 ( .A(n5492), .B(n5491), .Z(n1212) );
  NOR U3213 ( .A(n1213), .B(n1212), .Z(n5514) );
  XOR U3214 ( .A(n1214), .B(b[71]), .Z(n5513) );
  NOR U3215 ( .A(n5514), .B(n5513), .Z(n1215) );
  NOR U3216 ( .A(n1216), .B(n1215), .Z(n5536) );
  XOR U3217 ( .A(n1217), .B(b[72]), .Z(n5535) );
  NOR U3218 ( .A(n5536), .B(n5535), .Z(n1218) );
  NOR U3219 ( .A(n1219), .B(n1218), .Z(n5558) );
  XOR U3220 ( .A(n1220), .B(b[73]), .Z(n5557) );
  NOR U3221 ( .A(n5558), .B(n5557), .Z(n1221) );
  NOR U3222 ( .A(n1222), .B(n1221), .Z(n5580) );
  XOR U3223 ( .A(n1223), .B(b[74]), .Z(n5579) );
  NOR U3224 ( .A(n5580), .B(n5579), .Z(n1224) );
  NOR U3225 ( .A(n1225), .B(n1224), .Z(n5602) );
  XOR U3226 ( .A(n1226), .B(b[75]), .Z(n5601) );
  NOR U3227 ( .A(n5602), .B(n5601), .Z(n1227) );
  NOR U3228 ( .A(n1228), .B(n1227), .Z(n5624) );
  XOR U3229 ( .A(n1229), .B(b[76]), .Z(n5623) );
  NOR U3230 ( .A(n5624), .B(n5623), .Z(n1230) );
  NOR U3231 ( .A(n1231), .B(n1230), .Z(n5646) );
  XOR U3232 ( .A(n1232), .B(b[77]), .Z(n5645) );
  NOR U3233 ( .A(n5646), .B(n5645), .Z(n1233) );
  NOR U3234 ( .A(n1234), .B(n1233), .Z(n5668) );
  XOR U3235 ( .A(n1235), .B(b[78]), .Z(n5667) );
  NOR U3236 ( .A(n5668), .B(n5667), .Z(n1236) );
  NOR U3237 ( .A(n1237), .B(n1236), .Z(n5690) );
  XOR U3238 ( .A(n1238), .B(b[79]), .Z(n5689) );
  NOR U3239 ( .A(n5690), .B(n5689), .Z(n1239) );
  NOR U3240 ( .A(n1240), .B(n1239), .Z(n5714) );
  XOR U3241 ( .A(n1241), .B(b[80]), .Z(n5713) );
  NOR U3242 ( .A(n5714), .B(n5713), .Z(n1242) );
  NOR U3243 ( .A(n1243), .B(n1242), .Z(n5736) );
  XOR U3244 ( .A(n1244), .B(b[81]), .Z(n5735) );
  NOR U3245 ( .A(n5736), .B(n5735), .Z(n1245) );
  NOR U3246 ( .A(n1246), .B(n1245), .Z(n5758) );
  XOR U3247 ( .A(n1247), .B(b[82]), .Z(n5757) );
  NOR U3248 ( .A(n5758), .B(n5757), .Z(n1248) );
  NOR U3249 ( .A(n1249), .B(n1248), .Z(n5780) );
  XOR U3250 ( .A(n1250), .B(b[83]), .Z(n5779) );
  NOR U3251 ( .A(n5780), .B(n5779), .Z(n1251) );
  NOR U3252 ( .A(n1252), .B(n1251), .Z(n5802) );
  XOR U3253 ( .A(n1253), .B(b[84]), .Z(n5801) );
  NOR U3254 ( .A(n5802), .B(n5801), .Z(n1254) );
  NOR U3255 ( .A(n1255), .B(n1254), .Z(n5824) );
  XOR U3256 ( .A(n1256), .B(b[85]), .Z(n5823) );
  NOR U3257 ( .A(n5824), .B(n5823), .Z(n1257) );
  NOR U3258 ( .A(n1258), .B(n1257), .Z(n5846) );
  XOR U3259 ( .A(n1259), .B(b[86]), .Z(n5845) );
  NOR U3260 ( .A(n5846), .B(n5845), .Z(n1260) );
  NOR U3261 ( .A(n1261), .B(n1260), .Z(n5868) );
  XOR U3262 ( .A(n1262), .B(b[87]), .Z(n5867) );
  NOR U3263 ( .A(n5868), .B(n5867), .Z(n1263) );
  NOR U3264 ( .A(n1264), .B(n1263), .Z(n5890) );
  XOR U3265 ( .A(n1265), .B(b[88]), .Z(n5889) );
  NOR U3266 ( .A(n5890), .B(n5889), .Z(n1266) );
  NOR U3267 ( .A(n1267), .B(n1266), .Z(n5912) );
  XOR U3268 ( .A(n1268), .B(b[89]), .Z(n5911) );
  NOR U3269 ( .A(n5912), .B(n5911), .Z(n1269) );
  NOR U3270 ( .A(n1270), .B(n1269), .Z(n5936) );
  XOR U3271 ( .A(n1271), .B(b[90]), .Z(n5935) );
  NOR U3272 ( .A(n5936), .B(n5935), .Z(n1272) );
  NOR U3273 ( .A(n1273), .B(n1272), .Z(n5958) );
  XOR U3274 ( .A(n1274), .B(b[91]), .Z(n5957) );
  NOR U3275 ( .A(n5958), .B(n5957), .Z(n1275) );
  NOR U3276 ( .A(n1276), .B(n1275), .Z(n5980) );
  XOR U3277 ( .A(n1277), .B(b[92]), .Z(n5979) );
  NOR U3278 ( .A(n5980), .B(n5979), .Z(n1278) );
  NOR U3279 ( .A(n1279), .B(n1278), .Z(n6002) );
  XOR U3280 ( .A(n1280), .B(b[93]), .Z(n6001) );
  NOR U3281 ( .A(n6002), .B(n6001), .Z(n1281) );
  NOR U3282 ( .A(n1282), .B(n1281), .Z(n6024) );
  XOR U3283 ( .A(n1283), .B(b[94]), .Z(n6023) );
  NOR U3284 ( .A(n6024), .B(n6023), .Z(n1284) );
  NOR U3285 ( .A(n1285), .B(n1284), .Z(n6046) );
  XOR U3286 ( .A(n1286), .B(b[95]), .Z(n6045) );
  NOR U3287 ( .A(n6046), .B(n6045), .Z(n1287) );
  NOR U3288 ( .A(n1288), .B(n1287), .Z(n6068) );
  XOR U3289 ( .A(n1289), .B(b[96]), .Z(n6067) );
  NOR U3290 ( .A(n6068), .B(n6067), .Z(n1290) );
  NOR U3291 ( .A(n1291), .B(n1290), .Z(n6090) );
  XOR U3292 ( .A(n1292), .B(b[97]), .Z(n6089) );
  NOR U3293 ( .A(n6090), .B(n6089), .Z(n1293) );
  NOR U3294 ( .A(n1294), .B(n1293), .Z(n6112) );
  XOR U3295 ( .A(n1295), .B(b[98]), .Z(n6111) );
  NOR U3296 ( .A(n6112), .B(n6111), .Z(n1296) );
  NOR U3297 ( .A(n1297), .B(n1296), .Z(n6134) );
  XOR U3298 ( .A(n1298), .B(a[99]), .Z(n6133) );
  NOR U3299 ( .A(n6134), .B(n6133), .Z(n1299) );
  NOR U3300 ( .A(n1300), .B(n1299), .Z(n4056) );
  XOR U3301 ( .A(n1301), .B(b[100]), .Z(n4055) );
  NOR U3302 ( .A(n4056), .B(n4055), .Z(n1302) );
  NOR U3303 ( .A(n1303), .B(n1302), .Z(n4118) );
  XOR U3304 ( .A(n1304), .B(b[101]), .Z(n4117) );
  NOR U3305 ( .A(n4118), .B(n4117), .Z(n1305) );
  NOR U3306 ( .A(n1306), .B(n1305), .Z(n4144) );
  XOR U3307 ( .A(n1307), .B(b[102]), .Z(n4143) );
  NOR U3308 ( .A(n4144), .B(n4143), .Z(n1308) );
  NOR U3309 ( .A(n1309), .B(n1308), .Z(n4146) );
  XOR U3310 ( .A(n1310), .B(b[103]), .Z(n4145) );
  NOR U3311 ( .A(n4146), .B(n4145), .Z(n1311) );
  NOR U3312 ( .A(n1312), .B(n1311), .Z(n4148) );
  XOR U3313 ( .A(n1313), .B(b[104]), .Z(n4147) );
  NOR U3314 ( .A(n4148), .B(n4147), .Z(n1314) );
  NOR U3315 ( .A(n1315), .B(n1314), .Z(n4150) );
  XOR U3316 ( .A(n1316), .B(b[105]), .Z(n4149) );
  NOR U3317 ( .A(n4150), .B(n4149), .Z(n1317) );
  NOR U3318 ( .A(n1318), .B(n1317), .Z(n4152) );
  XOR U3319 ( .A(n1319), .B(b[106]), .Z(n4151) );
  NOR U3320 ( .A(n4152), .B(n4151), .Z(n1320) );
  NOR U3321 ( .A(n1321), .B(n1320), .Z(n4154) );
  XOR U3322 ( .A(n1322), .B(b[107]), .Z(n4153) );
  NOR U3323 ( .A(n4154), .B(n4153), .Z(n1323) );
  NOR U3324 ( .A(n1324), .B(n1323), .Z(n4156) );
  XOR U3325 ( .A(n1325), .B(b[108]), .Z(n4155) );
  NOR U3326 ( .A(n4156), .B(n4155), .Z(n1326) );
  NOR U3327 ( .A(n1327), .B(n1326), .Z(n4158) );
  XOR U3328 ( .A(n1328), .B(b[109]), .Z(n4157) );
  NOR U3329 ( .A(n4158), .B(n4157), .Z(n1329) );
  NOR U3330 ( .A(n1330), .B(n1329), .Z(n4162) );
  XOR U3331 ( .A(n1331), .B(b[110]), .Z(n4161) );
  NOR U3332 ( .A(n4162), .B(n4161), .Z(n1332) );
  NOR U3333 ( .A(n1333), .B(n1332), .Z(n4164) );
  XOR U3334 ( .A(n1334), .B(b[111]), .Z(n4163) );
  NOR U3335 ( .A(n4164), .B(n4163), .Z(n1335) );
  NOR U3336 ( .A(n1336), .B(n1335), .Z(n4166) );
  XOR U3337 ( .A(n1337), .B(b[112]), .Z(n4165) );
  NOR U3338 ( .A(n4166), .B(n4165), .Z(n1338) );
  NOR U3339 ( .A(n1339), .B(n1338), .Z(n4168) );
  XOR U3340 ( .A(n1340), .B(b[113]), .Z(n4167) );
  NOR U3341 ( .A(n4168), .B(n4167), .Z(n1341) );
  NOR U3342 ( .A(n1342), .B(n1341), .Z(n4170) );
  XOR U3343 ( .A(n1343), .B(b[114]), .Z(n4169) );
  NOR U3344 ( .A(n4170), .B(n4169), .Z(n1344) );
  NOR U3345 ( .A(n1345), .B(n1344), .Z(n4172) );
  XOR U3346 ( .A(n1346), .B(b[115]), .Z(n4171) );
  NOR U3347 ( .A(n4172), .B(n4171), .Z(n1347) );
  NOR U3348 ( .A(n1348), .B(n1347), .Z(n4174) );
  XOR U3349 ( .A(n1349), .B(b[116]), .Z(n4173) );
  NOR U3350 ( .A(n4174), .B(n4173), .Z(n1350) );
  NOR U3351 ( .A(n1351), .B(n1350), .Z(n4176) );
  XOR U3352 ( .A(n1352), .B(b[117]), .Z(n4175) );
  NOR U3353 ( .A(n4176), .B(n4175), .Z(n1353) );
  NOR U3354 ( .A(n1354), .B(n1353), .Z(n4178) );
  XOR U3355 ( .A(n1355), .B(b[118]), .Z(n4177) );
  NOR U3356 ( .A(n4178), .B(n4177), .Z(n1356) );
  NOR U3357 ( .A(n1357), .B(n1356), .Z(n4180) );
  XOR U3358 ( .A(n1358), .B(b[119]), .Z(n4179) );
  NOR U3359 ( .A(n4180), .B(n4179), .Z(n1359) );
  NOR U3360 ( .A(n1360), .B(n1359), .Z(n4184) );
  XOR U3361 ( .A(n1361), .B(b[120]), .Z(n4183) );
  NOR U3362 ( .A(n4184), .B(n4183), .Z(n1362) );
  NOR U3363 ( .A(n1363), .B(n1362), .Z(n4186) );
  XOR U3364 ( .A(n1364), .B(b[121]), .Z(n4185) );
  NOR U3365 ( .A(n4186), .B(n4185), .Z(n1365) );
  NOR U3366 ( .A(n1366), .B(n1365), .Z(n4188) );
  XOR U3367 ( .A(n1367), .B(b[122]), .Z(n4187) );
  NOR U3368 ( .A(n4188), .B(n4187), .Z(n1368) );
  NOR U3369 ( .A(n1369), .B(n1368), .Z(n4190) );
  XOR U3370 ( .A(n1370), .B(b[123]), .Z(n4189) );
  NOR U3371 ( .A(n4190), .B(n4189), .Z(n1371) );
  NOR U3372 ( .A(n1372), .B(n1371), .Z(n4192) );
  XOR U3373 ( .A(n1373), .B(b[124]), .Z(n4191) );
  NOR U3374 ( .A(n4192), .B(n4191), .Z(n1374) );
  NOR U3375 ( .A(n1375), .B(n1374), .Z(n4194) );
  XOR U3376 ( .A(n1376), .B(b[125]), .Z(n4193) );
  NOR U3377 ( .A(n4194), .B(n4193), .Z(n1377) );
  NOR U3378 ( .A(n1378), .B(n1377), .Z(n4196) );
  XOR U3379 ( .A(n1379), .B(b[126]), .Z(n4195) );
  NOR U3380 ( .A(n4196), .B(n4195), .Z(n1380) );
  NOR U3381 ( .A(n1381), .B(n1380), .Z(n4198) );
  XOR U3382 ( .A(n1382), .B(b[127]), .Z(n4197) );
  NOR U3383 ( .A(n4198), .B(n4197), .Z(n1383) );
  NOR U3384 ( .A(n1384), .B(n1383), .Z(n4200) );
  XOR U3385 ( .A(n1385), .B(b[128]), .Z(n4199) );
  NOR U3386 ( .A(n4200), .B(n4199), .Z(n1386) );
  NOR U3387 ( .A(n1387), .B(n1386), .Z(n4202) );
  XOR U3388 ( .A(n1388), .B(b[129]), .Z(n4201) );
  NOR U3389 ( .A(n4202), .B(n4201), .Z(n1389) );
  NOR U3390 ( .A(n1390), .B(n1389), .Z(n4206) );
  XOR U3391 ( .A(n1391), .B(b[130]), .Z(n4205) );
  NOR U3392 ( .A(n4206), .B(n4205), .Z(n1392) );
  NOR U3393 ( .A(n1393), .B(n1392), .Z(n4208) );
  XOR U3394 ( .A(n1394), .B(b[131]), .Z(n4207) );
  NOR U3395 ( .A(n4208), .B(n4207), .Z(n1395) );
  NOR U3396 ( .A(n1396), .B(n1395), .Z(n4210) );
  XOR U3397 ( .A(n1397), .B(b[132]), .Z(n4209) );
  NOR U3398 ( .A(n4210), .B(n4209), .Z(n1398) );
  NOR U3399 ( .A(n1399), .B(n1398), .Z(n4212) );
  XOR U3400 ( .A(n1400), .B(b[133]), .Z(n4211) );
  NOR U3401 ( .A(n4212), .B(n4211), .Z(n1401) );
  NOR U3402 ( .A(n1402), .B(n1401), .Z(n4214) );
  XOR U3403 ( .A(n1403), .B(b[134]), .Z(n4213) );
  NOR U3404 ( .A(n4214), .B(n4213), .Z(n1404) );
  NOR U3405 ( .A(n1405), .B(n1404), .Z(n4216) );
  XOR U3406 ( .A(n1406), .B(b[135]), .Z(n4215) );
  NOR U3407 ( .A(n4216), .B(n4215), .Z(n1407) );
  NOR U3408 ( .A(n1408), .B(n1407), .Z(n4218) );
  XOR U3409 ( .A(n1409), .B(b[136]), .Z(n4217) );
  NOR U3410 ( .A(n4218), .B(n4217), .Z(n1410) );
  NOR U3411 ( .A(n1411), .B(n1410), .Z(n4220) );
  XOR U3412 ( .A(n1412), .B(b[137]), .Z(n4219) );
  NOR U3413 ( .A(n4220), .B(n4219), .Z(n1413) );
  NOR U3414 ( .A(n1414), .B(n1413), .Z(n4222) );
  XOR U3415 ( .A(n1415), .B(b[138]), .Z(n4221) );
  NOR U3416 ( .A(n4222), .B(n4221), .Z(n1416) );
  NOR U3417 ( .A(n1417), .B(n1416), .Z(n4224) );
  XOR U3418 ( .A(n1418), .B(b[139]), .Z(n4223) );
  NOR U3419 ( .A(n4224), .B(n4223), .Z(n1419) );
  NOR U3420 ( .A(n1420), .B(n1419), .Z(n4228) );
  XOR U3421 ( .A(n1421), .B(b[140]), .Z(n4227) );
  NOR U3422 ( .A(n4228), .B(n4227), .Z(n1422) );
  NOR U3423 ( .A(n1423), .B(n1422), .Z(n4230) );
  XOR U3424 ( .A(n1424), .B(b[141]), .Z(n4229) );
  NOR U3425 ( .A(n4230), .B(n4229), .Z(n1425) );
  NOR U3426 ( .A(n1426), .B(n1425), .Z(n4232) );
  XOR U3427 ( .A(n1427), .B(b[142]), .Z(n4231) );
  NOR U3428 ( .A(n4232), .B(n4231), .Z(n1428) );
  NOR U3429 ( .A(n1429), .B(n1428), .Z(n4234) );
  XOR U3430 ( .A(n1430), .B(b[143]), .Z(n4233) );
  NOR U3431 ( .A(n4234), .B(n4233), .Z(n1431) );
  NOR U3432 ( .A(n1432), .B(n1431), .Z(n4236) );
  XOR U3433 ( .A(n1433), .B(b[144]), .Z(n4235) );
  NOR U3434 ( .A(n4236), .B(n4235), .Z(n1434) );
  NOR U3435 ( .A(n1435), .B(n1434), .Z(n4238) );
  XOR U3436 ( .A(n1436), .B(b[145]), .Z(n4237) );
  NOR U3437 ( .A(n4238), .B(n4237), .Z(n1437) );
  NOR U3438 ( .A(n1438), .B(n1437), .Z(n4240) );
  XOR U3439 ( .A(n1439), .B(b[146]), .Z(n4239) );
  NOR U3440 ( .A(n4240), .B(n4239), .Z(n1440) );
  NOR U3441 ( .A(n1441), .B(n1440), .Z(n4242) );
  XOR U3442 ( .A(n1442), .B(b[147]), .Z(n4241) );
  NOR U3443 ( .A(n4242), .B(n4241), .Z(n1443) );
  NOR U3444 ( .A(n1444), .B(n1443), .Z(n4244) );
  XOR U3445 ( .A(n1445), .B(b[148]), .Z(n4243) );
  NOR U3446 ( .A(n4244), .B(n4243), .Z(n1446) );
  NOR U3447 ( .A(n1447), .B(n1446), .Z(n4246) );
  XOR U3448 ( .A(n1448), .B(b[149]), .Z(n4245) );
  NOR U3449 ( .A(n4246), .B(n4245), .Z(n1449) );
  NOR U3450 ( .A(n1450), .B(n1449), .Z(n4250) );
  XOR U3451 ( .A(n1451), .B(b[150]), .Z(n4249) );
  NOR U3452 ( .A(n4250), .B(n4249), .Z(n1452) );
  NOR U3453 ( .A(n1453), .B(n1452), .Z(n4252) );
  XOR U3454 ( .A(n1454), .B(b[151]), .Z(n4251) );
  NOR U3455 ( .A(n4252), .B(n4251), .Z(n1455) );
  NOR U3456 ( .A(n1456), .B(n1455), .Z(n4254) );
  XOR U3457 ( .A(n1457), .B(b[152]), .Z(n4253) );
  NOR U3458 ( .A(n4254), .B(n4253), .Z(n1458) );
  NOR U3459 ( .A(n1459), .B(n1458), .Z(n4256) );
  XOR U3460 ( .A(n1460), .B(b[153]), .Z(n4255) );
  NOR U3461 ( .A(n4256), .B(n4255), .Z(n1461) );
  NOR U3462 ( .A(n1462), .B(n1461), .Z(n4258) );
  XOR U3463 ( .A(n1463), .B(b[154]), .Z(n4257) );
  NOR U3464 ( .A(n4258), .B(n4257), .Z(n1464) );
  NOR U3465 ( .A(n1465), .B(n1464), .Z(n4260) );
  XOR U3466 ( .A(n1466), .B(b[155]), .Z(n4259) );
  NOR U3467 ( .A(n4260), .B(n4259), .Z(n1467) );
  NOR U3468 ( .A(n1468), .B(n1467), .Z(n4262) );
  XOR U3469 ( .A(n1469), .B(b[156]), .Z(n4261) );
  NOR U3470 ( .A(n4262), .B(n4261), .Z(n1470) );
  NOR U3471 ( .A(n1471), .B(n1470), .Z(n4264) );
  XOR U3472 ( .A(n1472), .B(b[157]), .Z(n4263) );
  NOR U3473 ( .A(n4264), .B(n4263), .Z(n1473) );
  NOR U3474 ( .A(n1474), .B(n1473), .Z(n4266) );
  XOR U3475 ( .A(n1475), .B(b[158]), .Z(n4265) );
  NOR U3476 ( .A(n4266), .B(n4265), .Z(n1476) );
  NOR U3477 ( .A(n1477), .B(n1476), .Z(n4268) );
  XOR U3478 ( .A(n1478), .B(b[159]), .Z(n4267) );
  NOR U3479 ( .A(n4268), .B(n4267), .Z(n1479) );
  NOR U3480 ( .A(n1480), .B(n1479), .Z(n4272) );
  XOR U3481 ( .A(n1481), .B(b[160]), .Z(n4271) );
  NOR U3482 ( .A(n4272), .B(n4271), .Z(n1482) );
  NOR U3483 ( .A(n1483), .B(n1482), .Z(n4274) );
  XOR U3484 ( .A(n1484), .B(b[161]), .Z(n4273) );
  NOR U3485 ( .A(n4274), .B(n4273), .Z(n1485) );
  NOR U3486 ( .A(n1486), .B(n1485), .Z(n4276) );
  XOR U3487 ( .A(n1487), .B(b[162]), .Z(n4275) );
  NOR U3488 ( .A(n4276), .B(n4275), .Z(n1488) );
  NOR U3489 ( .A(n1489), .B(n1488), .Z(n4278) );
  XOR U3490 ( .A(n1490), .B(b[163]), .Z(n4277) );
  NOR U3491 ( .A(n4278), .B(n4277), .Z(n1491) );
  NOR U3492 ( .A(n1492), .B(n1491), .Z(n4280) );
  XOR U3493 ( .A(n1493), .B(b[164]), .Z(n4279) );
  NOR U3494 ( .A(n4280), .B(n4279), .Z(n1494) );
  NOR U3495 ( .A(n1495), .B(n1494), .Z(n4282) );
  XOR U3496 ( .A(n1496), .B(b[165]), .Z(n4281) );
  NOR U3497 ( .A(n4282), .B(n4281), .Z(n1497) );
  NOR U3498 ( .A(n1498), .B(n1497), .Z(n4284) );
  XOR U3499 ( .A(n1499), .B(b[166]), .Z(n4283) );
  NOR U3500 ( .A(n4284), .B(n4283), .Z(n1500) );
  NOR U3501 ( .A(n1501), .B(n1500), .Z(n4286) );
  XOR U3502 ( .A(n1502), .B(b[167]), .Z(n4285) );
  NOR U3503 ( .A(n4286), .B(n4285), .Z(n1503) );
  NOR U3504 ( .A(n1504), .B(n1503), .Z(n4288) );
  XOR U3505 ( .A(n1505), .B(b[168]), .Z(n4287) );
  NOR U3506 ( .A(n4288), .B(n4287), .Z(n1506) );
  NOR U3507 ( .A(n1507), .B(n1506), .Z(n4290) );
  XOR U3508 ( .A(n1508), .B(b[169]), .Z(n4289) );
  NOR U3509 ( .A(n4290), .B(n4289), .Z(n1509) );
  NOR U3510 ( .A(n1510), .B(n1509), .Z(n4294) );
  XOR U3511 ( .A(n1511), .B(b[170]), .Z(n4293) );
  NOR U3512 ( .A(n4294), .B(n4293), .Z(n1512) );
  NOR U3513 ( .A(n1513), .B(n1512), .Z(n4296) );
  XOR U3514 ( .A(n1514), .B(b[171]), .Z(n4295) );
  NOR U3515 ( .A(n4296), .B(n4295), .Z(n1515) );
  NOR U3516 ( .A(n1516), .B(n1515), .Z(n4298) );
  XOR U3517 ( .A(n1517), .B(b[172]), .Z(n4297) );
  NOR U3518 ( .A(n4298), .B(n4297), .Z(n1518) );
  NOR U3519 ( .A(n1519), .B(n1518), .Z(n4300) );
  XOR U3520 ( .A(n1520), .B(b[173]), .Z(n4299) );
  NOR U3521 ( .A(n4300), .B(n4299), .Z(n1521) );
  NOR U3522 ( .A(n1522), .B(n1521), .Z(n4302) );
  XOR U3523 ( .A(n1523), .B(b[174]), .Z(n4301) );
  NOR U3524 ( .A(n4302), .B(n4301), .Z(n1524) );
  NOR U3525 ( .A(n1525), .B(n1524), .Z(n4304) );
  XOR U3526 ( .A(n1526), .B(b[175]), .Z(n4303) );
  NOR U3527 ( .A(n4304), .B(n4303), .Z(n1527) );
  NOR U3528 ( .A(n1528), .B(n1527), .Z(n4306) );
  XOR U3529 ( .A(n1529), .B(b[176]), .Z(n4305) );
  NOR U3530 ( .A(n4306), .B(n4305), .Z(n1530) );
  NOR U3531 ( .A(n1531), .B(n1530), .Z(n4308) );
  XOR U3532 ( .A(n1532), .B(b[177]), .Z(n4307) );
  NOR U3533 ( .A(n4308), .B(n4307), .Z(n1533) );
  NOR U3534 ( .A(n1534), .B(n1533), .Z(n4310) );
  XOR U3535 ( .A(n1535), .B(b[178]), .Z(n4309) );
  NOR U3536 ( .A(n4310), .B(n4309), .Z(n1536) );
  NOR U3537 ( .A(n1537), .B(n1536), .Z(n4312) );
  XOR U3538 ( .A(n1538), .B(b[179]), .Z(n4311) );
  NOR U3539 ( .A(n4312), .B(n4311), .Z(n1539) );
  NOR U3540 ( .A(n1540), .B(n1539), .Z(n4316) );
  XOR U3541 ( .A(n1541), .B(b[180]), .Z(n4315) );
  NOR U3542 ( .A(n4316), .B(n4315), .Z(n1542) );
  NOR U3543 ( .A(n1543), .B(n1542), .Z(n4318) );
  XOR U3544 ( .A(n1544), .B(b[181]), .Z(n4317) );
  NOR U3545 ( .A(n4318), .B(n4317), .Z(n1545) );
  NOR U3546 ( .A(n1546), .B(n1545), .Z(n4320) );
  XOR U3547 ( .A(n1547), .B(b[182]), .Z(n4319) );
  NOR U3548 ( .A(n4320), .B(n4319), .Z(n1548) );
  NOR U3549 ( .A(n1549), .B(n1548), .Z(n4322) );
  XOR U3550 ( .A(n1550), .B(b[183]), .Z(n4321) );
  NOR U3551 ( .A(n4322), .B(n4321), .Z(n1551) );
  NOR U3552 ( .A(n1552), .B(n1551), .Z(n4324) );
  XOR U3553 ( .A(n1553), .B(b[184]), .Z(n4323) );
  NOR U3554 ( .A(n4324), .B(n4323), .Z(n1554) );
  NOR U3555 ( .A(n1555), .B(n1554), .Z(n4326) );
  XOR U3556 ( .A(n1556), .B(b[185]), .Z(n4325) );
  NOR U3557 ( .A(n4326), .B(n4325), .Z(n1557) );
  NOR U3558 ( .A(n1558), .B(n1557), .Z(n4328) );
  XOR U3559 ( .A(n1559), .B(b[186]), .Z(n4327) );
  NOR U3560 ( .A(n4328), .B(n4327), .Z(n1560) );
  NOR U3561 ( .A(n1561), .B(n1560), .Z(n4330) );
  XOR U3562 ( .A(n1562), .B(b[187]), .Z(n4329) );
  NOR U3563 ( .A(n4330), .B(n4329), .Z(n1563) );
  NOR U3564 ( .A(n1564), .B(n1563), .Z(n4332) );
  XOR U3565 ( .A(n1565), .B(b[188]), .Z(n4331) );
  NOR U3566 ( .A(n4332), .B(n4331), .Z(n1566) );
  NOR U3567 ( .A(n1567), .B(n1566), .Z(n4334) );
  XOR U3568 ( .A(n1568), .B(b[189]), .Z(n4333) );
  NOR U3569 ( .A(n4334), .B(n4333), .Z(n1569) );
  NOR U3570 ( .A(n1570), .B(n1569), .Z(n4338) );
  XOR U3571 ( .A(n1571), .B(b[190]), .Z(n4337) );
  NOR U3572 ( .A(n4338), .B(n4337), .Z(n1572) );
  NOR U3573 ( .A(n1573), .B(n1572), .Z(n4340) );
  XOR U3574 ( .A(n1574), .B(b[191]), .Z(n4339) );
  NOR U3575 ( .A(n4340), .B(n4339), .Z(n1575) );
  NOR U3576 ( .A(n1576), .B(n1575), .Z(n4342) );
  XOR U3577 ( .A(n1577), .B(b[192]), .Z(n4341) );
  NOR U3578 ( .A(n4342), .B(n4341), .Z(n1578) );
  NOR U3579 ( .A(n1579), .B(n1578), .Z(n4344) );
  XOR U3580 ( .A(n1580), .B(b[193]), .Z(n4343) );
  NOR U3581 ( .A(n4344), .B(n4343), .Z(n1581) );
  NOR U3582 ( .A(n1582), .B(n1581), .Z(n4346) );
  XOR U3583 ( .A(n1583), .B(b[194]), .Z(n4345) );
  NOR U3584 ( .A(n4346), .B(n4345), .Z(n1584) );
  NOR U3585 ( .A(n1585), .B(n1584), .Z(n4348) );
  XOR U3586 ( .A(n1586), .B(b[195]), .Z(n4347) );
  NOR U3587 ( .A(n4348), .B(n4347), .Z(n1587) );
  NOR U3588 ( .A(n1588), .B(n1587), .Z(n4350) );
  XOR U3589 ( .A(n1589), .B(b[196]), .Z(n4349) );
  NOR U3590 ( .A(n4350), .B(n4349), .Z(n1590) );
  NOR U3591 ( .A(n1591), .B(n1590), .Z(n4352) );
  XOR U3592 ( .A(n1592), .B(b[197]), .Z(n4351) );
  NOR U3593 ( .A(n4352), .B(n4351), .Z(n1593) );
  NOR U3594 ( .A(n1594), .B(n1593), .Z(n4354) );
  XOR U3595 ( .A(n1595), .B(b[198]), .Z(n4353) );
  NOR U3596 ( .A(n4354), .B(n4353), .Z(n1596) );
  NOR U3597 ( .A(n1597), .B(n1596), .Z(n4356) );
  XOR U3598 ( .A(n1598), .B(b[199]), .Z(n4355) );
  NOR U3599 ( .A(n4356), .B(n4355), .Z(n1599) );
  NOR U3600 ( .A(n1600), .B(n1599), .Z(n4362) );
  XOR U3601 ( .A(n1601), .B(b[200]), .Z(n4361) );
  NOR U3602 ( .A(n4362), .B(n4361), .Z(n1602) );
  NOR U3603 ( .A(n1603), .B(n1602), .Z(n4364) );
  XOR U3604 ( .A(n1604), .B(b[201]), .Z(n4363) );
  NOR U3605 ( .A(n4364), .B(n4363), .Z(n1605) );
  NOR U3606 ( .A(n1606), .B(n1605), .Z(n4366) );
  XOR U3607 ( .A(n1607), .B(b[202]), .Z(n4365) );
  NOR U3608 ( .A(n4366), .B(n4365), .Z(n1608) );
  NOR U3609 ( .A(n1609), .B(n1608), .Z(n4368) );
  XOR U3610 ( .A(n1610), .B(b[203]), .Z(n4367) );
  NOR U3611 ( .A(n4368), .B(n4367), .Z(n1611) );
  NOR U3612 ( .A(n1612), .B(n1611), .Z(n4370) );
  XOR U3613 ( .A(n1613), .B(b[204]), .Z(n4369) );
  NOR U3614 ( .A(n4370), .B(n4369), .Z(n1614) );
  NOR U3615 ( .A(n1615), .B(n1614), .Z(n4372) );
  XOR U3616 ( .A(n1616), .B(b[205]), .Z(n4371) );
  NOR U3617 ( .A(n4372), .B(n4371), .Z(n1617) );
  NOR U3618 ( .A(n1618), .B(n1617), .Z(n4374) );
  XOR U3619 ( .A(n1619), .B(b[206]), .Z(n4373) );
  NOR U3620 ( .A(n4374), .B(n4373), .Z(n1620) );
  NOR U3621 ( .A(n1621), .B(n1620), .Z(n4376) );
  XOR U3622 ( .A(n1622), .B(b[207]), .Z(n4375) );
  NOR U3623 ( .A(n4376), .B(n4375), .Z(n1623) );
  NOR U3624 ( .A(n1624), .B(n1623), .Z(n4378) );
  XOR U3625 ( .A(n1625), .B(b[208]), .Z(n4377) );
  NOR U3626 ( .A(n4378), .B(n4377), .Z(n1626) );
  NOR U3627 ( .A(n1627), .B(n1626), .Z(n4380) );
  XOR U3628 ( .A(n1628), .B(b[209]), .Z(n4379) );
  NOR U3629 ( .A(n4380), .B(n4379), .Z(n1629) );
  NOR U3630 ( .A(n1630), .B(n1629), .Z(n4384) );
  XOR U3631 ( .A(n1631), .B(b[210]), .Z(n4383) );
  NOR U3632 ( .A(n4384), .B(n4383), .Z(n1632) );
  NOR U3633 ( .A(n1633), .B(n1632), .Z(n4386) );
  XOR U3634 ( .A(n1634), .B(b[211]), .Z(n4385) );
  NOR U3635 ( .A(n4386), .B(n4385), .Z(n1635) );
  NOR U3636 ( .A(n1636), .B(n1635), .Z(n4388) );
  XOR U3637 ( .A(n1637), .B(b[212]), .Z(n4387) );
  NOR U3638 ( .A(n4388), .B(n4387), .Z(n1638) );
  NOR U3639 ( .A(n1639), .B(n1638), .Z(n4390) );
  XOR U3640 ( .A(n1640), .B(b[213]), .Z(n4389) );
  NOR U3641 ( .A(n4390), .B(n4389), .Z(n1641) );
  NOR U3642 ( .A(n1642), .B(n1641), .Z(n4392) );
  XOR U3643 ( .A(n1643), .B(b[214]), .Z(n4391) );
  NOR U3644 ( .A(n4392), .B(n4391), .Z(n1644) );
  NOR U3645 ( .A(n1645), .B(n1644), .Z(n4394) );
  XOR U3646 ( .A(n1646), .B(b[215]), .Z(n4393) );
  NOR U3647 ( .A(n4394), .B(n4393), .Z(n1647) );
  NOR U3648 ( .A(n1648), .B(n1647), .Z(n4396) );
  XOR U3649 ( .A(n1649), .B(b[216]), .Z(n4395) );
  NOR U3650 ( .A(n4396), .B(n4395), .Z(n1650) );
  NOR U3651 ( .A(n1651), .B(n1650), .Z(n4398) );
  XOR U3652 ( .A(n1652), .B(b[217]), .Z(n4397) );
  NOR U3653 ( .A(n4398), .B(n4397), .Z(n1653) );
  NOR U3654 ( .A(n1654), .B(n1653), .Z(n4400) );
  XOR U3655 ( .A(n1655), .B(b[218]), .Z(n4399) );
  NOR U3656 ( .A(n4400), .B(n4399), .Z(n1656) );
  NOR U3657 ( .A(n1657), .B(n1656), .Z(n4402) );
  XOR U3658 ( .A(n1658), .B(b[219]), .Z(n4401) );
  NOR U3659 ( .A(n4402), .B(n4401), .Z(n1659) );
  NOR U3660 ( .A(n1660), .B(n1659), .Z(n4406) );
  XOR U3661 ( .A(n1661), .B(b[220]), .Z(n4405) );
  NOR U3662 ( .A(n4406), .B(n4405), .Z(n1662) );
  NOR U3663 ( .A(n1663), .B(n1662), .Z(n4408) );
  XOR U3664 ( .A(n1664), .B(b[221]), .Z(n4407) );
  NOR U3665 ( .A(n4408), .B(n4407), .Z(n1665) );
  NOR U3666 ( .A(n1666), .B(n1665), .Z(n4410) );
  XOR U3667 ( .A(n1667), .B(b[222]), .Z(n4409) );
  NOR U3668 ( .A(n4410), .B(n4409), .Z(n1668) );
  NOR U3669 ( .A(n1669), .B(n1668), .Z(n4412) );
  XOR U3670 ( .A(n1670), .B(b[223]), .Z(n4411) );
  NOR U3671 ( .A(n4412), .B(n4411), .Z(n1671) );
  NOR U3672 ( .A(n1672), .B(n1671), .Z(n4414) );
  XOR U3673 ( .A(n1673), .B(b[224]), .Z(n4413) );
  NOR U3674 ( .A(n4414), .B(n4413), .Z(n1674) );
  NOR U3675 ( .A(n1675), .B(n1674), .Z(n4416) );
  XOR U3676 ( .A(n1676), .B(b[225]), .Z(n4415) );
  NOR U3677 ( .A(n4416), .B(n4415), .Z(n1677) );
  NOR U3678 ( .A(n1678), .B(n1677), .Z(n4418) );
  XOR U3679 ( .A(n1679), .B(b[226]), .Z(n4417) );
  NOR U3680 ( .A(n4418), .B(n4417), .Z(n1680) );
  NOR U3681 ( .A(n1681), .B(n1680), .Z(n4420) );
  XOR U3682 ( .A(n1682), .B(b[227]), .Z(n4419) );
  NOR U3683 ( .A(n4420), .B(n4419), .Z(n1683) );
  NOR U3684 ( .A(n1684), .B(n1683), .Z(n4422) );
  XOR U3685 ( .A(n1685), .B(b[228]), .Z(n4421) );
  NOR U3686 ( .A(n4422), .B(n4421), .Z(n1686) );
  NOR U3687 ( .A(n1687), .B(n1686), .Z(n4424) );
  XOR U3688 ( .A(n1688), .B(b[229]), .Z(n4423) );
  NOR U3689 ( .A(n4424), .B(n4423), .Z(n1689) );
  NOR U3690 ( .A(n1690), .B(n1689), .Z(n4428) );
  XOR U3691 ( .A(n1691), .B(b[230]), .Z(n4427) );
  NOR U3692 ( .A(n4428), .B(n4427), .Z(n1692) );
  NOR U3693 ( .A(n1693), .B(n1692), .Z(n4430) );
  XOR U3694 ( .A(n1694), .B(b[231]), .Z(n4429) );
  NOR U3695 ( .A(n4430), .B(n4429), .Z(n1695) );
  NOR U3696 ( .A(n1696), .B(n1695), .Z(n4432) );
  XOR U3697 ( .A(n1697), .B(b[232]), .Z(n4431) );
  NOR U3698 ( .A(n4432), .B(n4431), .Z(n1698) );
  NOR U3699 ( .A(n1699), .B(n1698), .Z(n4434) );
  XOR U3700 ( .A(n1700), .B(b[233]), .Z(n4433) );
  NOR U3701 ( .A(n4434), .B(n4433), .Z(n1701) );
  NOR U3702 ( .A(n1702), .B(n1701), .Z(n4436) );
  XOR U3703 ( .A(n1703), .B(b[234]), .Z(n4435) );
  NOR U3704 ( .A(n4436), .B(n4435), .Z(n1704) );
  NOR U3705 ( .A(n1705), .B(n1704), .Z(n4438) );
  XOR U3706 ( .A(n1706), .B(b[235]), .Z(n4437) );
  NOR U3707 ( .A(n4438), .B(n4437), .Z(n1707) );
  NOR U3708 ( .A(n1708), .B(n1707), .Z(n4440) );
  XOR U3709 ( .A(n1709), .B(b[236]), .Z(n4439) );
  NOR U3710 ( .A(n4440), .B(n4439), .Z(n1710) );
  NOR U3711 ( .A(n1711), .B(n1710), .Z(n4442) );
  XOR U3712 ( .A(n1712), .B(b[237]), .Z(n4441) );
  NOR U3713 ( .A(n4442), .B(n4441), .Z(n1713) );
  NOR U3714 ( .A(n1714), .B(n1713), .Z(n4444) );
  XOR U3715 ( .A(n1715), .B(b[238]), .Z(n4443) );
  NOR U3716 ( .A(n4444), .B(n4443), .Z(n1716) );
  NOR U3717 ( .A(n1717), .B(n1716), .Z(n4446) );
  XOR U3718 ( .A(n1718), .B(b[239]), .Z(n4445) );
  NOR U3719 ( .A(n4446), .B(n4445), .Z(n1719) );
  NOR U3720 ( .A(n1720), .B(n1719), .Z(n4450) );
  XOR U3721 ( .A(n1721), .B(b[240]), .Z(n4449) );
  NOR U3722 ( .A(n4450), .B(n4449), .Z(n1722) );
  NOR U3723 ( .A(n1723), .B(n1722), .Z(n4452) );
  XOR U3724 ( .A(n1724), .B(b[241]), .Z(n4451) );
  NOR U3725 ( .A(n4452), .B(n4451), .Z(n1725) );
  NOR U3726 ( .A(n1726), .B(n1725), .Z(n4454) );
  XOR U3727 ( .A(n1727), .B(b[242]), .Z(n4453) );
  NOR U3728 ( .A(n4454), .B(n4453), .Z(n1728) );
  NOR U3729 ( .A(n1729), .B(n1728), .Z(n4456) );
  XOR U3730 ( .A(n1730), .B(b[243]), .Z(n4455) );
  NOR U3731 ( .A(n4456), .B(n4455), .Z(n1731) );
  NOR U3732 ( .A(n1732), .B(n1731), .Z(n4458) );
  XOR U3733 ( .A(n1733), .B(b[244]), .Z(n4457) );
  NOR U3734 ( .A(n4458), .B(n4457), .Z(n1734) );
  NOR U3735 ( .A(n1735), .B(n1734), .Z(n4460) );
  XOR U3736 ( .A(n1736), .B(b[245]), .Z(n4459) );
  NOR U3737 ( .A(n4460), .B(n4459), .Z(n1737) );
  NOR U3738 ( .A(n1738), .B(n1737), .Z(n4462) );
  XOR U3739 ( .A(n1739), .B(b[246]), .Z(n4461) );
  NOR U3740 ( .A(n4462), .B(n4461), .Z(n1740) );
  NOR U3741 ( .A(n1741), .B(n1740), .Z(n4464) );
  XOR U3742 ( .A(n1742), .B(b[247]), .Z(n4463) );
  NOR U3743 ( .A(n4464), .B(n4463), .Z(n1743) );
  NOR U3744 ( .A(n1744), .B(n1743), .Z(n4466) );
  XOR U3745 ( .A(n1745), .B(b[248]), .Z(n4465) );
  NOR U3746 ( .A(n4466), .B(n4465), .Z(n1746) );
  NOR U3747 ( .A(n1747), .B(n1746), .Z(n4468) );
  XOR U3748 ( .A(n1748), .B(b[249]), .Z(n4467) );
  NOR U3749 ( .A(n4468), .B(n4467), .Z(n1749) );
  NOR U3750 ( .A(n1750), .B(n1749), .Z(n4472) );
  XOR U3751 ( .A(n1751), .B(b[250]), .Z(n4471) );
  NOR U3752 ( .A(n4472), .B(n4471), .Z(n1752) );
  NOR U3753 ( .A(n1753), .B(n1752), .Z(n4474) );
  XOR U3754 ( .A(n1754), .B(b[251]), .Z(n4473) );
  NOR U3755 ( .A(n4474), .B(n4473), .Z(n1755) );
  NOR U3756 ( .A(n1756), .B(n1755), .Z(n4476) );
  XOR U3757 ( .A(n1757), .B(b[252]), .Z(n4475) );
  NOR U3758 ( .A(n4476), .B(n4475), .Z(n1758) );
  NOR U3759 ( .A(n1759), .B(n1758), .Z(n4478) );
  XOR U3760 ( .A(n1760), .B(b[253]), .Z(n4477) );
  NOR U3761 ( .A(n4478), .B(n4477), .Z(n1761) );
  NOR U3762 ( .A(n1762), .B(n1761), .Z(n4480) );
  XOR U3763 ( .A(n1763), .B(b[254]), .Z(n4479) );
  NOR U3764 ( .A(n4480), .B(n4479), .Z(n1764) );
  NOR U3765 ( .A(n1765), .B(n1764), .Z(n4482) );
  XOR U3766 ( .A(n1766), .B(b[255]), .Z(n4481) );
  NOR U3767 ( .A(n4482), .B(n4481), .Z(n1767) );
  NOR U3768 ( .A(n1768), .B(n1767), .Z(n4484) );
  XOR U3769 ( .A(n1769), .B(b[256]), .Z(n4483) );
  NOR U3770 ( .A(n4484), .B(n4483), .Z(n1770) );
  NOR U3771 ( .A(n1771), .B(n1770), .Z(n4486) );
  XOR U3772 ( .A(n1772), .B(b[257]), .Z(n4485) );
  NOR U3773 ( .A(n4486), .B(n4485), .Z(n1773) );
  NOR U3774 ( .A(n1774), .B(n1773), .Z(n4488) );
  XOR U3775 ( .A(n1775), .B(b[258]), .Z(n4487) );
  NOR U3776 ( .A(n4488), .B(n4487), .Z(n1776) );
  NOR U3777 ( .A(n1777), .B(n1776), .Z(n4490) );
  XOR U3778 ( .A(n1778), .B(b[259]), .Z(n4489) );
  NOR U3779 ( .A(n4490), .B(n4489), .Z(n1779) );
  NOR U3780 ( .A(n1780), .B(n1779), .Z(n4494) );
  XOR U3781 ( .A(n1781), .B(b[260]), .Z(n4493) );
  NOR U3782 ( .A(n4494), .B(n4493), .Z(n1782) );
  NOR U3783 ( .A(n1783), .B(n1782), .Z(n4496) );
  XOR U3784 ( .A(n1784), .B(b[261]), .Z(n4495) );
  NOR U3785 ( .A(n4496), .B(n4495), .Z(n1785) );
  NOR U3786 ( .A(n1786), .B(n1785), .Z(n4498) );
  XOR U3787 ( .A(n1787), .B(b[262]), .Z(n4497) );
  NOR U3788 ( .A(n4498), .B(n4497), .Z(n1788) );
  NOR U3789 ( .A(n1789), .B(n1788), .Z(n4500) );
  XOR U3790 ( .A(n1790), .B(b[263]), .Z(n4499) );
  NOR U3791 ( .A(n4500), .B(n4499), .Z(n1791) );
  NOR U3792 ( .A(n1792), .B(n1791), .Z(n4502) );
  XOR U3793 ( .A(n1793), .B(b[264]), .Z(n4501) );
  NOR U3794 ( .A(n4502), .B(n4501), .Z(n1794) );
  NOR U3795 ( .A(n1795), .B(n1794), .Z(n4504) );
  XOR U3796 ( .A(n1796), .B(b[265]), .Z(n4503) );
  NOR U3797 ( .A(n4504), .B(n4503), .Z(n1797) );
  NOR U3798 ( .A(n1798), .B(n1797), .Z(n4506) );
  XOR U3799 ( .A(n1799), .B(b[266]), .Z(n4505) );
  NOR U3800 ( .A(n4506), .B(n4505), .Z(n1800) );
  NOR U3801 ( .A(n1801), .B(n1800), .Z(n4508) );
  XOR U3802 ( .A(n1802), .B(b[267]), .Z(n4507) );
  NOR U3803 ( .A(n4508), .B(n4507), .Z(n1803) );
  NOR U3804 ( .A(n1804), .B(n1803), .Z(n4510) );
  XOR U3805 ( .A(n1805), .B(b[268]), .Z(n4509) );
  NOR U3806 ( .A(n4510), .B(n4509), .Z(n1806) );
  NOR U3807 ( .A(n1807), .B(n1806), .Z(n4512) );
  XOR U3808 ( .A(n1808), .B(b[269]), .Z(n4511) );
  NOR U3809 ( .A(n4512), .B(n4511), .Z(n1809) );
  NOR U3810 ( .A(n1810), .B(n1809), .Z(n4516) );
  XOR U3811 ( .A(n1811), .B(b[270]), .Z(n4515) );
  NOR U3812 ( .A(n4516), .B(n4515), .Z(n1812) );
  NOR U3813 ( .A(n1813), .B(n1812), .Z(n4518) );
  XOR U3814 ( .A(n1814), .B(b[271]), .Z(n4517) );
  NOR U3815 ( .A(n4518), .B(n4517), .Z(n1815) );
  NOR U3816 ( .A(n1816), .B(n1815), .Z(n4520) );
  XOR U3817 ( .A(n1817), .B(b[272]), .Z(n4519) );
  NOR U3818 ( .A(n4520), .B(n4519), .Z(n1818) );
  NOR U3819 ( .A(n1819), .B(n1818), .Z(n4522) );
  XOR U3820 ( .A(n1820), .B(b[273]), .Z(n4521) );
  NOR U3821 ( .A(n4522), .B(n4521), .Z(n1821) );
  NOR U3822 ( .A(n1822), .B(n1821), .Z(n4524) );
  XOR U3823 ( .A(n1823), .B(b[274]), .Z(n4523) );
  NOR U3824 ( .A(n4524), .B(n4523), .Z(n1824) );
  NOR U3825 ( .A(n1825), .B(n1824), .Z(n4526) );
  XOR U3826 ( .A(n1826), .B(b[275]), .Z(n4525) );
  NOR U3827 ( .A(n4526), .B(n4525), .Z(n1827) );
  NOR U3828 ( .A(n1828), .B(n1827), .Z(n4528) );
  XOR U3829 ( .A(n1829), .B(b[276]), .Z(n4527) );
  NOR U3830 ( .A(n4528), .B(n4527), .Z(n1830) );
  NOR U3831 ( .A(n1831), .B(n1830), .Z(n4530) );
  XOR U3832 ( .A(n1832), .B(b[277]), .Z(n4529) );
  NOR U3833 ( .A(n4530), .B(n4529), .Z(n1833) );
  NOR U3834 ( .A(n1834), .B(n1833), .Z(n4532) );
  XOR U3835 ( .A(n1835), .B(b[278]), .Z(n4531) );
  NOR U3836 ( .A(n4532), .B(n4531), .Z(n1836) );
  NOR U3837 ( .A(n1837), .B(n1836), .Z(n4534) );
  XOR U3838 ( .A(n1838), .B(b[279]), .Z(n4533) );
  NOR U3839 ( .A(n4534), .B(n4533), .Z(n1839) );
  NOR U3840 ( .A(n1840), .B(n1839), .Z(n4538) );
  XOR U3841 ( .A(n1841), .B(b[280]), .Z(n4537) );
  NOR U3842 ( .A(n4538), .B(n4537), .Z(n1842) );
  NOR U3843 ( .A(n1843), .B(n1842), .Z(n4540) );
  XOR U3844 ( .A(n1844), .B(b[281]), .Z(n4539) );
  NOR U3845 ( .A(n4540), .B(n4539), .Z(n1845) );
  NOR U3846 ( .A(n1846), .B(n1845), .Z(n4542) );
  XOR U3847 ( .A(n1847), .B(b[282]), .Z(n4541) );
  NOR U3848 ( .A(n4542), .B(n4541), .Z(n1848) );
  NOR U3849 ( .A(n1849), .B(n1848), .Z(n4544) );
  XOR U3850 ( .A(n1850), .B(b[283]), .Z(n4543) );
  NOR U3851 ( .A(n4544), .B(n4543), .Z(n1851) );
  NOR U3852 ( .A(n1852), .B(n1851), .Z(n4546) );
  XOR U3853 ( .A(n1853), .B(b[284]), .Z(n4545) );
  NOR U3854 ( .A(n4546), .B(n4545), .Z(n1854) );
  NOR U3855 ( .A(n1855), .B(n1854), .Z(n4548) );
  XOR U3856 ( .A(n1856), .B(b[285]), .Z(n4547) );
  NOR U3857 ( .A(n4548), .B(n4547), .Z(n1857) );
  NOR U3858 ( .A(n1858), .B(n1857), .Z(n4550) );
  XOR U3859 ( .A(n1859), .B(b[286]), .Z(n4549) );
  NOR U3860 ( .A(n4550), .B(n4549), .Z(n1860) );
  NOR U3861 ( .A(n1861), .B(n1860), .Z(n4552) );
  XOR U3862 ( .A(n1862), .B(b[287]), .Z(n4551) );
  NOR U3863 ( .A(n4552), .B(n4551), .Z(n1863) );
  NOR U3864 ( .A(n1864), .B(n1863), .Z(n4554) );
  XOR U3865 ( .A(n1865), .B(b[288]), .Z(n4553) );
  NOR U3866 ( .A(n4554), .B(n4553), .Z(n1866) );
  NOR U3867 ( .A(n1867), .B(n1866), .Z(n4556) );
  XOR U3868 ( .A(n1868), .B(b[289]), .Z(n4555) );
  NOR U3869 ( .A(n4556), .B(n4555), .Z(n1869) );
  NOR U3870 ( .A(n1870), .B(n1869), .Z(n4560) );
  XOR U3871 ( .A(n1871), .B(b[290]), .Z(n4559) );
  NOR U3872 ( .A(n4560), .B(n4559), .Z(n1872) );
  NOR U3873 ( .A(n1873), .B(n1872), .Z(n4562) );
  XOR U3874 ( .A(n1874), .B(b[291]), .Z(n4561) );
  NOR U3875 ( .A(n4562), .B(n4561), .Z(n1875) );
  NOR U3876 ( .A(n1876), .B(n1875), .Z(n4564) );
  XOR U3877 ( .A(n1877), .B(b[292]), .Z(n4563) );
  NOR U3878 ( .A(n4564), .B(n4563), .Z(n1878) );
  NOR U3879 ( .A(n1879), .B(n1878), .Z(n4566) );
  XOR U3880 ( .A(n1880), .B(b[293]), .Z(n4565) );
  NOR U3881 ( .A(n4566), .B(n4565), .Z(n1881) );
  NOR U3882 ( .A(n1882), .B(n1881), .Z(n4568) );
  XOR U3883 ( .A(n1883), .B(b[294]), .Z(n4567) );
  NOR U3884 ( .A(n4568), .B(n4567), .Z(n1884) );
  NOR U3885 ( .A(n1885), .B(n1884), .Z(n4570) );
  XOR U3886 ( .A(n1886), .B(b[295]), .Z(n4569) );
  NOR U3887 ( .A(n4570), .B(n4569), .Z(n1887) );
  NOR U3888 ( .A(n1888), .B(n1887), .Z(n4572) );
  XOR U3889 ( .A(n1889), .B(b[296]), .Z(n4571) );
  NOR U3890 ( .A(n4572), .B(n4571), .Z(n1890) );
  NOR U3891 ( .A(n1891), .B(n1890), .Z(n4574) );
  XOR U3892 ( .A(n1892), .B(b[297]), .Z(n4573) );
  NOR U3893 ( .A(n4574), .B(n4573), .Z(n1893) );
  NOR U3894 ( .A(n1894), .B(n1893), .Z(n4576) );
  XOR U3895 ( .A(n1895), .B(b[298]), .Z(n4575) );
  NOR U3896 ( .A(n4576), .B(n4575), .Z(n1896) );
  NOR U3897 ( .A(n1897), .B(n1896), .Z(n4578) );
  XOR U3898 ( .A(n1898), .B(b[299]), .Z(n4577) );
  NOR U3899 ( .A(n4578), .B(n4577), .Z(n1899) );
  NOR U3900 ( .A(n1900), .B(n1899), .Z(n4584) );
  XOR U3901 ( .A(n1901), .B(b[300]), .Z(n4583) );
  NOR U3902 ( .A(n4584), .B(n4583), .Z(n1902) );
  NOR U3903 ( .A(n1903), .B(n1902), .Z(n4586) );
  XOR U3904 ( .A(n1904), .B(b[301]), .Z(n4585) );
  NOR U3905 ( .A(n4586), .B(n4585), .Z(n1905) );
  NOR U3906 ( .A(n1906), .B(n1905), .Z(n4588) );
  XOR U3907 ( .A(n1907), .B(b[302]), .Z(n4587) );
  NOR U3908 ( .A(n4588), .B(n4587), .Z(n1908) );
  NOR U3909 ( .A(n1909), .B(n1908), .Z(n4590) );
  XOR U3910 ( .A(n1910), .B(b[303]), .Z(n4589) );
  NOR U3911 ( .A(n4590), .B(n4589), .Z(n1911) );
  NOR U3912 ( .A(n1912), .B(n1911), .Z(n4592) );
  XOR U3913 ( .A(n1913), .B(b[304]), .Z(n4591) );
  NOR U3914 ( .A(n4592), .B(n4591), .Z(n1914) );
  NOR U3915 ( .A(n1915), .B(n1914), .Z(n4594) );
  XOR U3916 ( .A(n1916), .B(b[305]), .Z(n4593) );
  NOR U3917 ( .A(n4594), .B(n4593), .Z(n1917) );
  NOR U3918 ( .A(n1918), .B(n1917), .Z(n4596) );
  XOR U3919 ( .A(n1919), .B(b[306]), .Z(n4595) );
  NOR U3920 ( .A(n4596), .B(n4595), .Z(n1920) );
  NOR U3921 ( .A(n1921), .B(n1920), .Z(n4598) );
  XOR U3922 ( .A(n1922), .B(b[307]), .Z(n4597) );
  NOR U3923 ( .A(n4598), .B(n4597), .Z(n1923) );
  NOR U3924 ( .A(n1924), .B(n1923), .Z(n4600) );
  XOR U3925 ( .A(n1925), .B(b[308]), .Z(n4599) );
  NOR U3926 ( .A(n4600), .B(n4599), .Z(n1926) );
  NOR U3927 ( .A(n1927), .B(n1926), .Z(n4602) );
  XOR U3928 ( .A(n1928), .B(b[309]), .Z(n4601) );
  NOR U3929 ( .A(n4602), .B(n4601), .Z(n1929) );
  NOR U3930 ( .A(n1930), .B(n1929), .Z(n4606) );
  XOR U3931 ( .A(n1931), .B(b[310]), .Z(n4605) );
  NOR U3932 ( .A(n4606), .B(n4605), .Z(n1932) );
  NOR U3933 ( .A(n1933), .B(n1932), .Z(n4608) );
  XOR U3934 ( .A(n1934), .B(b[311]), .Z(n4607) );
  NOR U3935 ( .A(n4608), .B(n4607), .Z(n1935) );
  NOR U3936 ( .A(n1936), .B(n1935), .Z(n4610) );
  XOR U3937 ( .A(n1937), .B(b[312]), .Z(n4609) );
  NOR U3938 ( .A(n4610), .B(n4609), .Z(n1938) );
  NOR U3939 ( .A(n1939), .B(n1938), .Z(n4612) );
  XOR U3940 ( .A(n1940), .B(b[313]), .Z(n4611) );
  NOR U3941 ( .A(n4612), .B(n4611), .Z(n1941) );
  NOR U3942 ( .A(n1942), .B(n1941), .Z(n4614) );
  XOR U3943 ( .A(n1943), .B(b[314]), .Z(n4613) );
  NOR U3944 ( .A(n4614), .B(n4613), .Z(n1944) );
  NOR U3945 ( .A(n1945), .B(n1944), .Z(n4616) );
  XOR U3946 ( .A(n1946), .B(b[315]), .Z(n4615) );
  NOR U3947 ( .A(n4616), .B(n4615), .Z(n1947) );
  NOR U3948 ( .A(n1948), .B(n1947), .Z(n4618) );
  XOR U3949 ( .A(n1949), .B(b[316]), .Z(n4617) );
  NOR U3950 ( .A(n4618), .B(n4617), .Z(n1950) );
  NOR U3951 ( .A(n1951), .B(n1950), .Z(n4620) );
  XOR U3952 ( .A(n1952), .B(b[317]), .Z(n4619) );
  NOR U3953 ( .A(n4620), .B(n4619), .Z(n1953) );
  NOR U3954 ( .A(n1954), .B(n1953), .Z(n4622) );
  XOR U3955 ( .A(n1955), .B(b[318]), .Z(n4621) );
  NOR U3956 ( .A(n4622), .B(n4621), .Z(n1956) );
  NOR U3957 ( .A(n1957), .B(n1956), .Z(n4624) );
  XOR U3958 ( .A(n1958), .B(b[319]), .Z(n4623) );
  NOR U3959 ( .A(n4624), .B(n4623), .Z(n1959) );
  NOR U3960 ( .A(n1960), .B(n1959), .Z(n4628) );
  XOR U3961 ( .A(n1961), .B(b[320]), .Z(n4627) );
  NOR U3962 ( .A(n4628), .B(n4627), .Z(n1962) );
  NOR U3963 ( .A(n1963), .B(n1962), .Z(n4630) );
  XOR U3964 ( .A(n1964), .B(b[321]), .Z(n4629) );
  NOR U3965 ( .A(n4630), .B(n4629), .Z(n1965) );
  NOR U3966 ( .A(n1966), .B(n1965), .Z(n4632) );
  XOR U3967 ( .A(n1967), .B(b[322]), .Z(n4631) );
  NOR U3968 ( .A(n4632), .B(n4631), .Z(n1968) );
  NOR U3969 ( .A(n1969), .B(n1968), .Z(n4634) );
  XOR U3970 ( .A(n1970), .B(b[323]), .Z(n4633) );
  NOR U3971 ( .A(n4634), .B(n4633), .Z(n1971) );
  NOR U3972 ( .A(n1972), .B(n1971), .Z(n4636) );
  XOR U3973 ( .A(n1973), .B(b[324]), .Z(n4635) );
  NOR U3974 ( .A(n4636), .B(n4635), .Z(n1974) );
  NOR U3975 ( .A(n1975), .B(n1974), .Z(n4638) );
  XOR U3976 ( .A(n1976), .B(b[325]), .Z(n4637) );
  NOR U3977 ( .A(n4638), .B(n4637), .Z(n1977) );
  NOR U3978 ( .A(n1978), .B(n1977), .Z(n4640) );
  XOR U3979 ( .A(n1979), .B(b[326]), .Z(n4639) );
  NOR U3980 ( .A(n4640), .B(n4639), .Z(n1980) );
  NOR U3981 ( .A(n1981), .B(n1980), .Z(n4642) );
  XOR U3982 ( .A(n1982), .B(b[327]), .Z(n4641) );
  NOR U3983 ( .A(n4642), .B(n4641), .Z(n1983) );
  NOR U3984 ( .A(n1984), .B(n1983), .Z(n4644) );
  XOR U3985 ( .A(n1985), .B(b[328]), .Z(n4643) );
  NOR U3986 ( .A(n4644), .B(n4643), .Z(n1986) );
  NOR U3987 ( .A(n1987), .B(n1986), .Z(n4646) );
  XOR U3988 ( .A(n1988), .B(b[329]), .Z(n4645) );
  NOR U3989 ( .A(n4646), .B(n4645), .Z(n1989) );
  NOR U3990 ( .A(n1990), .B(n1989), .Z(n4650) );
  XOR U3991 ( .A(n1991), .B(b[330]), .Z(n4649) );
  NOR U3992 ( .A(n4650), .B(n4649), .Z(n1992) );
  NOR U3993 ( .A(n1993), .B(n1992), .Z(n4652) );
  XOR U3994 ( .A(n1994), .B(b[331]), .Z(n4651) );
  NOR U3995 ( .A(n4652), .B(n4651), .Z(n1995) );
  NOR U3996 ( .A(n1996), .B(n1995), .Z(n4654) );
  XOR U3997 ( .A(n1997), .B(b[332]), .Z(n4653) );
  NOR U3998 ( .A(n4654), .B(n4653), .Z(n1998) );
  NOR U3999 ( .A(n1999), .B(n1998), .Z(n4656) );
  XOR U4000 ( .A(n2000), .B(b[333]), .Z(n4655) );
  NOR U4001 ( .A(n4656), .B(n4655), .Z(n2001) );
  NOR U4002 ( .A(n2002), .B(n2001), .Z(n4658) );
  XOR U4003 ( .A(n2003), .B(b[334]), .Z(n4657) );
  NOR U4004 ( .A(n4658), .B(n4657), .Z(n2004) );
  NOR U4005 ( .A(n2005), .B(n2004), .Z(n4660) );
  XOR U4006 ( .A(n2006), .B(b[335]), .Z(n4659) );
  NOR U4007 ( .A(n4660), .B(n4659), .Z(n2007) );
  NOR U4008 ( .A(n2008), .B(n2007), .Z(n4662) );
  XOR U4009 ( .A(n2009), .B(b[336]), .Z(n4661) );
  NOR U4010 ( .A(n4662), .B(n4661), .Z(n2010) );
  NOR U4011 ( .A(n2011), .B(n2010), .Z(n4664) );
  XOR U4012 ( .A(n2012), .B(b[337]), .Z(n4663) );
  NOR U4013 ( .A(n4664), .B(n4663), .Z(n2013) );
  NOR U4014 ( .A(n2014), .B(n2013), .Z(n4666) );
  XOR U4015 ( .A(n2015), .B(b[338]), .Z(n4665) );
  NOR U4016 ( .A(n4666), .B(n4665), .Z(n2016) );
  NOR U4017 ( .A(n2017), .B(n2016), .Z(n4668) );
  XOR U4018 ( .A(n2018), .B(b[339]), .Z(n4667) );
  NOR U4019 ( .A(n4668), .B(n4667), .Z(n2019) );
  NOR U4020 ( .A(n2020), .B(n2019), .Z(n4672) );
  XOR U4021 ( .A(n2021), .B(b[340]), .Z(n4671) );
  NOR U4022 ( .A(n4672), .B(n4671), .Z(n2022) );
  NOR U4023 ( .A(n2023), .B(n2022), .Z(n4674) );
  XOR U4024 ( .A(n2024), .B(b[341]), .Z(n4673) );
  NOR U4025 ( .A(n4674), .B(n4673), .Z(n2025) );
  NOR U4026 ( .A(n2026), .B(n2025), .Z(n4676) );
  XOR U4027 ( .A(n2027), .B(b[342]), .Z(n4675) );
  NOR U4028 ( .A(n4676), .B(n4675), .Z(n2028) );
  NOR U4029 ( .A(n2029), .B(n2028), .Z(n4678) );
  XOR U4030 ( .A(n2030), .B(b[343]), .Z(n4677) );
  NOR U4031 ( .A(n4678), .B(n4677), .Z(n2031) );
  NOR U4032 ( .A(n2032), .B(n2031), .Z(n4680) );
  XOR U4033 ( .A(n2033), .B(b[344]), .Z(n4679) );
  NOR U4034 ( .A(n4680), .B(n4679), .Z(n2034) );
  NOR U4035 ( .A(n2035), .B(n2034), .Z(n4682) );
  XOR U4036 ( .A(n2036), .B(b[345]), .Z(n4681) );
  NOR U4037 ( .A(n4682), .B(n4681), .Z(n2037) );
  NOR U4038 ( .A(n2038), .B(n2037), .Z(n4684) );
  XOR U4039 ( .A(n2039), .B(b[346]), .Z(n4683) );
  NOR U4040 ( .A(n4684), .B(n4683), .Z(n2040) );
  NOR U4041 ( .A(n2041), .B(n2040), .Z(n4686) );
  XOR U4042 ( .A(n2042), .B(b[347]), .Z(n4685) );
  NOR U4043 ( .A(n4686), .B(n4685), .Z(n2043) );
  NOR U4044 ( .A(n2044), .B(n2043), .Z(n4688) );
  XOR U4045 ( .A(n2045), .B(b[348]), .Z(n4687) );
  NOR U4046 ( .A(n4688), .B(n4687), .Z(n2046) );
  NOR U4047 ( .A(n2047), .B(n2046), .Z(n4690) );
  XOR U4048 ( .A(n2048), .B(b[349]), .Z(n4689) );
  NOR U4049 ( .A(n4690), .B(n4689), .Z(n2049) );
  NOR U4050 ( .A(n2050), .B(n2049), .Z(n4694) );
  XOR U4051 ( .A(n2051), .B(b[350]), .Z(n4693) );
  NOR U4052 ( .A(n4694), .B(n4693), .Z(n2052) );
  NOR U4053 ( .A(n2053), .B(n2052), .Z(n4696) );
  XOR U4054 ( .A(n2054), .B(b[351]), .Z(n4695) );
  NOR U4055 ( .A(n4696), .B(n4695), .Z(n2055) );
  NOR U4056 ( .A(n2056), .B(n2055), .Z(n4698) );
  XOR U4057 ( .A(n2057), .B(b[352]), .Z(n4697) );
  NOR U4058 ( .A(n4698), .B(n4697), .Z(n2058) );
  NOR U4059 ( .A(n2059), .B(n2058), .Z(n4700) );
  XOR U4060 ( .A(n2060), .B(b[353]), .Z(n4699) );
  NOR U4061 ( .A(n4700), .B(n4699), .Z(n2061) );
  NOR U4062 ( .A(n2062), .B(n2061), .Z(n4702) );
  XOR U4063 ( .A(n2063), .B(b[354]), .Z(n4701) );
  NOR U4064 ( .A(n4702), .B(n4701), .Z(n2064) );
  NOR U4065 ( .A(n2065), .B(n2064), .Z(n4704) );
  XOR U4066 ( .A(n2066), .B(b[355]), .Z(n4703) );
  NOR U4067 ( .A(n4704), .B(n4703), .Z(n2067) );
  NOR U4068 ( .A(n2068), .B(n2067), .Z(n4706) );
  XOR U4069 ( .A(n2069), .B(b[356]), .Z(n4705) );
  NOR U4070 ( .A(n4706), .B(n4705), .Z(n2070) );
  NOR U4071 ( .A(n2071), .B(n2070), .Z(n4708) );
  XOR U4072 ( .A(n2072), .B(b[357]), .Z(n4707) );
  NOR U4073 ( .A(n4708), .B(n4707), .Z(n2073) );
  NOR U4074 ( .A(n2074), .B(n2073), .Z(n4710) );
  XOR U4075 ( .A(n2075), .B(b[358]), .Z(n4709) );
  NOR U4076 ( .A(n4710), .B(n4709), .Z(n2076) );
  NOR U4077 ( .A(n2077), .B(n2076), .Z(n4712) );
  XOR U4078 ( .A(n2078), .B(b[359]), .Z(n4711) );
  NOR U4079 ( .A(n4712), .B(n4711), .Z(n2079) );
  NOR U4080 ( .A(n2080), .B(n2079), .Z(n4716) );
  XOR U4081 ( .A(n2081), .B(b[360]), .Z(n4715) );
  NOR U4082 ( .A(n4716), .B(n4715), .Z(n2082) );
  NOR U4083 ( .A(n2083), .B(n2082), .Z(n4718) );
  XOR U4084 ( .A(n2084), .B(b[361]), .Z(n4717) );
  NOR U4085 ( .A(n4718), .B(n4717), .Z(n2085) );
  NOR U4086 ( .A(n2086), .B(n2085), .Z(n4720) );
  XOR U4087 ( .A(n2087), .B(b[362]), .Z(n4719) );
  NOR U4088 ( .A(n4720), .B(n4719), .Z(n2088) );
  NOR U4089 ( .A(n2089), .B(n2088), .Z(n4722) );
  XOR U4090 ( .A(n2090), .B(b[363]), .Z(n4721) );
  NOR U4091 ( .A(n4722), .B(n4721), .Z(n2091) );
  NOR U4092 ( .A(n2092), .B(n2091), .Z(n4724) );
  XOR U4093 ( .A(n2093), .B(b[364]), .Z(n4723) );
  NOR U4094 ( .A(n4724), .B(n4723), .Z(n2094) );
  NOR U4095 ( .A(n2095), .B(n2094), .Z(n4726) );
  XOR U4096 ( .A(n2096), .B(b[365]), .Z(n4725) );
  NOR U4097 ( .A(n4726), .B(n4725), .Z(n2097) );
  NOR U4098 ( .A(n2098), .B(n2097), .Z(n4728) );
  XOR U4099 ( .A(n2099), .B(b[366]), .Z(n4727) );
  NOR U4100 ( .A(n4728), .B(n4727), .Z(n2100) );
  NOR U4101 ( .A(n2101), .B(n2100), .Z(n4730) );
  XOR U4102 ( .A(n2102), .B(b[367]), .Z(n4729) );
  NOR U4103 ( .A(n4730), .B(n4729), .Z(n2103) );
  NOR U4104 ( .A(n2104), .B(n2103), .Z(n4732) );
  XOR U4105 ( .A(n2105), .B(b[368]), .Z(n4731) );
  NOR U4106 ( .A(n4732), .B(n4731), .Z(n2106) );
  NOR U4107 ( .A(n2107), .B(n2106), .Z(n4734) );
  XOR U4108 ( .A(n2108), .B(b[369]), .Z(n4733) );
  NOR U4109 ( .A(n4734), .B(n4733), .Z(n2109) );
  NOR U4110 ( .A(n2110), .B(n2109), .Z(n4738) );
  XOR U4111 ( .A(n2111), .B(b[370]), .Z(n4737) );
  NOR U4112 ( .A(n4738), .B(n4737), .Z(n2112) );
  NOR U4113 ( .A(n2113), .B(n2112), .Z(n4740) );
  XOR U4114 ( .A(n2114), .B(b[371]), .Z(n4739) );
  NOR U4115 ( .A(n4740), .B(n4739), .Z(n2115) );
  NOR U4116 ( .A(n2116), .B(n2115), .Z(n4742) );
  XOR U4117 ( .A(n2117), .B(b[372]), .Z(n4741) );
  NOR U4118 ( .A(n4742), .B(n4741), .Z(n2118) );
  NOR U4119 ( .A(n2119), .B(n2118), .Z(n4744) );
  XOR U4120 ( .A(n2120), .B(b[373]), .Z(n4743) );
  NOR U4121 ( .A(n4744), .B(n4743), .Z(n2121) );
  NOR U4122 ( .A(n2122), .B(n2121), .Z(n4746) );
  XOR U4123 ( .A(n2123), .B(b[374]), .Z(n4745) );
  NOR U4124 ( .A(n4746), .B(n4745), .Z(n2124) );
  NOR U4125 ( .A(n2125), .B(n2124), .Z(n4748) );
  XOR U4126 ( .A(n2126), .B(b[375]), .Z(n4747) );
  NOR U4127 ( .A(n4748), .B(n4747), .Z(n2127) );
  NOR U4128 ( .A(n2128), .B(n2127), .Z(n4750) );
  XOR U4129 ( .A(n2129), .B(b[376]), .Z(n4749) );
  NOR U4130 ( .A(n4750), .B(n4749), .Z(n2130) );
  NOR U4131 ( .A(n2131), .B(n2130), .Z(n4752) );
  XOR U4132 ( .A(n2132), .B(b[377]), .Z(n4751) );
  NOR U4133 ( .A(n4752), .B(n4751), .Z(n2133) );
  NOR U4134 ( .A(n2134), .B(n2133), .Z(n4754) );
  XOR U4135 ( .A(n2135), .B(b[378]), .Z(n4753) );
  NOR U4136 ( .A(n4754), .B(n4753), .Z(n2136) );
  NOR U4137 ( .A(n2137), .B(n2136), .Z(n4756) );
  XOR U4138 ( .A(n2138), .B(b[379]), .Z(n4755) );
  NOR U4139 ( .A(n4756), .B(n4755), .Z(n2139) );
  NOR U4140 ( .A(n2140), .B(n2139), .Z(n4760) );
  XOR U4141 ( .A(n2141), .B(b[380]), .Z(n4759) );
  NOR U4142 ( .A(n4760), .B(n4759), .Z(n2142) );
  NOR U4143 ( .A(n2143), .B(n2142), .Z(n4762) );
  XOR U4144 ( .A(n2144), .B(b[381]), .Z(n4761) );
  NOR U4145 ( .A(n4762), .B(n4761), .Z(n2145) );
  NOR U4146 ( .A(n2146), .B(n2145), .Z(n4764) );
  XOR U4147 ( .A(n2147), .B(b[382]), .Z(n4763) );
  NOR U4148 ( .A(n4764), .B(n4763), .Z(n2148) );
  NOR U4149 ( .A(n2149), .B(n2148), .Z(n4766) );
  XOR U4150 ( .A(n2150), .B(b[383]), .Z(n4765) );
  NOR U4151 ( .A(n4766), .B(n4765), .Z(n2151) );
  NOR U4152 ( .A(n2152), .B(n2151), .Z(n4768) );
  XOR U4153 ( .A(n2153), .B(b[384]), .Z(n4767) );
  NOR U4154 ( .A(n4768), .B(n4767), .Z(n2154) );
  NOR U4155 ( .A(n2155), .B(n2154), .Z(n4770) );
  XOR U4156 ( .A(n2156), .B(b[385]), .Z(n4769) );
  NOR U4157 ( .A(n4770), .B(n4769), .Z(n2157) );
  NOR U4158 ( .A(n2158), .B(n2157), .Z(n4772) );
  XOR U4159 ( .A(n2159), .B(b[386]), .Z(n4771) );
  NOR U4160 ( .A(n4772), .B(n4771), .Z(n2160) );
  NOR U4161 ( .A(n2161), .B(n2160), .Z(n4774) );
  XOR U4162 ( .A(n2162), .B(b[387]), .Z(n4773) );
  NOR U4163 ( .A(n4774), .B(n4773), .Z(n2163) );
  NOR U4164 ( .A(n2164), .B(n2163), .Z(n4776) );
  XOR U4165 ( .A(n2165), .B(b[388]), .Z(n4775) );
  NOR U4166 ( .A(n4776), .B(n4775), .Z(n2166) );
  NOR U4167 ( .A(n2167), .B(n2166), .Z(n4778) );
  XOR U4168 ( .A(n2168), .B(b[389]), .Z(n4777) );
  NOR U4169 ( .A(n4778), .B(n4777), .Z(n2169) );
  NOR U4170 ( .A(n2170), .B(n2169), .Z(n4782) );
  XOR U4171 ( .A(n2171), .B(b[390]), .Z(n4781) );
  NOR U4172 ( .A(n4782), .B(n4781), .Z(n2172) );
  NOR U4173 ( .A(n2173), .B(n2172), .Z(n4784) );
  XOR U4174 ( .A(n2174), .B(b[391]), .Z(n4783) );
  NOR U4175 ( .A(n4784), .B(n4783), .Z(n2175) );
  NOR U4176 ( .A(n2176), .B(n2175), .Z(n4786) );
  XOR U4177 ( .A(n2177), .B(b[392]), .Z(n4785) );
  NOR U4178 ( .A(n4786), .B(n4785), .Z(n2178) );
  NOR U4179 ( .A(n2179), .B(n2178), .Z(n4788) );
  XOR U4180 ( .A(n2180), .B(b[393]), .Z(n4787) );
  NOR U4181 ( .A(n4788), .B(n4787), .Z(n2181) );
  NOR U4182 ( .A(n2182), .B(n2181), .Z(n4790) );
  XOR U4183 ( .A(n2183), .B(b[394]), .Z(n4789) );
  NOR U4184 ( .A(n4790), .B(n4789), .Z(n2184) );
  NOR U4185 ( .A(n2185), .B(n2184), .Z(n4792) );
  XOR U4186 ( .A(n2186), .B(b[395]), .Z(n4791) );
  NOR U4187 ( .A(n4792), .B(n4791), .Z(n2187) );
  NOR U4188 ( .A(n2188), .B(n2187), .Z(n4794) );
  XOR U4189 ( .A(n2189), .B(b[396]), .Z(n4793) );
  NOR U4190 ( .A(n4794), .B(n4793), .Z(n2190) );
  NOR U4191 ( .A(n2191), .B(n2190), .Z(n4796) );
  XOR U4192 ( .A(n2192), .B(b[397]), .Z(n4795) );
  NOR U4193 ( .A(n4796), .B(n4795), .Z(n2193) );
  NOR U4194 ( .A(n2194), .B(n2193), .Z(n4798) );
  XOR U4195 ( .A(n2195), .B(b[398]), .Z(n4797) );
  NOR U4196 ( .A(n4798), .B(n4797), .Z(n2196) );
  NOR U4197 ( .A(n2197), .B(n2196), .Z(n4800) );
  XOR U4198 ( .A(n2198), .B(b[399]), .Z(n4799) );
  NOR U4199 ( .A(n4800), .B(n4799), .Z(n2199) );
  NOR U4200 ( .A(n2200), .B(n2199), .Z(n4806) );
  XOR U4201 ( .A(n2201), .B(b[400]), .Z(n4805) );
  NOR U4202 ( .A(n4806), .B(n4805), .Z(n2202) );
  NOR U4203 ( .A(n2203), .B(n2202), .Z(n4808) );
  XOR U4204 ( .A(n2204), .B(b[401]), .Z(n4807) );
  NOR U4205 ( .A(n4808), .B(n4807), .Z(n2205) );
  NOR U4206 ( .A(n2206), .B(n2205), .Z(n4810) );
  XOR U4207 ( .A(n2207), .B(b[402]), .Z(n4809) );
  NOR U4208 ( .A(n4810), .B(n4809), .Z(n2208) );
  NOR U4209 ( .A(n2209), .B(n2208), .Z(n4812) );
  XOR U4210 ( .A(n2210), .B(b[403]), .Z(n4811) );
  NOR U4211 ( .A(n4812), .B(n4811), .Z(n2211) );
  NOR U4212 ( .A(n2212), .B(n2211), .Z(n4814) );
  XOR U4213 ( .A(n2213), .B(b[404]), .Z(n4813) );
  NOR U4214 ( .A(n4814), .B(n4813), .Z(n2214) );
  NOR U4215 ( .A(n2215), .B(n2214), .Z(n4816) );
  XOR U4216 ( .A(n2216), .B(b[405]), .Z(n4815) );
  NOR U4217 ( .A(n4816), .B(n4815), .Z(n2217) );
  NOR U4218 ( .A(n2218), .B(n2217), .Z(n4818) );
  XOR U4219 ( .A(n2219), .B(b[406]), .Z(n4817) );
  NOR U4220 ( .A(n4818), .B(n4817), .Z(n2220) );
  NOR U4221 ( .A(n2221), .B(n2220), .Z(n4820) );
  XOR U4222 ( .A(n2222), .B(b[407]), .Z(n4819) );
  NOR U4223 ( .A(n4820), .B(n4819), .Z(n2223) );
  NOR U4224 ( .A(n2224), .B(n2223), .Z(n4822) );
  XOR U4225 ( .A(n2225), .B(b[408]), .Z(n4821) );
  NOR U4226 ( .A(n4822), .B(n4821), .Z(n2226) );
  NOR U4227 ( .A(n2227), .B(n2226), .Z(n4824) );
  XOR U4228 ( .A(n2228), .B(b[409]), .Z(n4823) );
  NOR U4229 ( .A(n4824), .B(n4823), .Z(n2229) );
  NOR U4230 ( .A(n2230), .B(n2229), .Z(n4828) );
  XOR U4231 ( .A(n2231), .B(b[410]), .Z(n4827) );
  NOR U4232 ( .A(n4828), .B(n4827), .Z(n2232) );
  NOR U4233 ( .A(n2233), .B(n2232), .Z(n4830) );
  XOR U4234 ( .A(n2234), .B(b[411]), .Z(n4829) );
  NOR U4235 ( .A(n4830), .B(n4829), .Z(n2235) );
  NOR U4236 ( .A(n2236), .B(n2235), .Z(n4832) );
  XOR U4237 ( .A(n2237), .B(b[412]), .Z(n4831) );
  NOR U4238 ( .A(n4832), .B(n4831), .Z(n2238) );
  NOR U4239 ( .A(n2239), .B(n2238), .Z(n4834) );
  XOR U4240 ( .A(n2240), .B(b[413]), .Z(n4833) );
  NOR U4241 ( .A(n4834), .B(n4833), .Z(n2241) );
  NOR U4242 ( .A(n2242), .B(n2241), .Z(n4836) );
  XOR U4243 ( .A(n2243), .B(b[414]), .Z(n4835) );
  NOR U4244 ( .A(n4836), .B(n4835), .Z(n2244) );
  NOR U4245 ( .A(n2245), .B(n2244), .Z(n4838) );
  XOR U4246 ( .A(n2246), .B(b[415]), .Z(n4837) );
  NOR U4247 ( .A(n4838), .B(n4837), .Z(n2247) );
  NOR U4248 ( .A(n2248), .B(n2247), .Z(n4840) );
  XOR U4249 ( .A(n2249), .B(b[416]), .Z(n4839) );
  NOR U4250 ( .A(n4840), .B(n4839), .Z(n2250) );
  NOR U4251 ( .A(n2251), .B(n2250), .Z(n4842) );
  XOR U4252 ( .A(n2252), .B(b[417]), .Z(n4841) );
  NOR U4253 ( .A(n4842), .B(n4841), .Z(n2253) );
  NOR U4254 ( .A(n2254), .B(n2253), .Z(n4844) );
  XOR U4255 ( .A(n2255), .B(b[418]), .Z(n4843) );
  NOR U4256 ( .A(n4844), .B(n4843), .Z(n2256) );
  NOR U4257 ( .A(n2257), .B(n2256), .Z(n4846) );
  XOR U4258 ( .A(n2258), .B(b[419]), .Z(n4845) );
  NOR U4259 ( .A(n4846), .B(n4845), .Z(n2259) );
  NOR U4260 ( .A(n2260), .B(n2259), .Z(n4850) );
  XOR U4261 ( .A(n2261), .B(b[420]), .Z(n4849) );
  NOR U4262 ( .A(n4850), .B(n4849), .Z(n2262) );
  NOR U4263 ( .A(n2263), .B(n2262), .Z(n4852) );
  XOR U4264 ( .A(n2264), .B(b[421]), .Z(n4851) );
  NOR U4265 ( .A(n4852), .B(n4851), .Z(n2265) );
  NOR U4266 ( .A(n2266), .B(n2265), .Z(n4854) );
  XOR U4267 ( .A(n2267), .B(b[422]), .Z(n4853) );
  NOR U4268 ( .A(n4854), .B(n4853), .Z(n2268) );
  NOR U4269 ( .A(n2269), .B(n2268), .Z(n4856) );
  XOR U4270 ( .A(n2270), .B(b[423]), .Z(n4855) );
  NOR U4271 ( .A(n4856), .B(n4855), .Z(n2271) );
  NOR U4272 ( .A(n2272), .B(n2271), .Z(n4858) );
  XOR U4273 ( .A(n2273), .B(b[424]), .Z(n4857) );
  NOR U4274 ( .A(n4858), .B(n4857), .Z(n2274) );
  NOR U4275 ( .A(n2275), .B(n2274), .Z(n4860) );
  XOR U4276 ( .A(n2276), .B(b[425]), .Z(n4859) );
  NOR U4277 ( .A(n4860), .B(n4859), .Z(n2277) );
  NOR U4278 ( .A(n2278), .B(n2277), .Z(n4862) );
  XOR U4279 ( .A(n2279), .B(b[426]), .Z(n4861) );
  NOR U4280 ( .A(n4862), .B(n4861), .Z(n2280) );
  NOR U4281 ( .A(n2281), .B(n2280), .Z(n4864) );
  XOR U4282 ( .A(n2282), .B(b[427]), .Z(n4863) );
  NOR U4283 ( .A(n4864), .B(n4863), .Z(n2283) );
  NOR U4284 ( .A(n2284), .B(n2283), .Z(n4866) );
  XOR U4285 ( .A(n2285), .B(b[428]), .Z(n4865) );
  NOR U4286 ( .A(n4866), .B(n4865), .Z(n2286) );
  NOR U4287 ( .A(n2287), .B(n2286), .Z(n4868) );
  XOR U4288 ( .A(n2288), .B(b[429]), .Z(n4867) );
  NOR U4289 ( .A(n4868), .B(n4867), .Z(n2289) );
  NOR U4290 ( .A(n2290), .B(n2289), .Z(n4872) );
  XOR U4291 ( .A(n2291), .B(b[430]), .Z(n4871) );
  NOR U4292 ( .A(n4872), .B(n4871), .Z(n2292) );
  NOR U4293 ( .A(n2293), .B(n2292), .Z(n4874) );
  XOR U4294 ( .A(n2294), .B(b[431]), .Z(n4873) );
  NOR U4295 ( .A(n4874), .B(n4873), .Z(n2295) );
  NOR U4296 ( .A(n2296), .B(n2295), .Z(n4876) );
  XOR U4297 ( .A(n2297), .B(b[432]), .Z(n4875) );
  NOR U4298 ( .A(n4876), .B(n4875), .Z(n2298) );
  NOR U4299 ( .A(n2299), .B(n2298), .Z(n4878) );
  XOR U4300 ( .A(n2300), .B(b[433]), .Z(n4877) );
  NOR U4301 ( .A(n4878), .B(n4877), .Z(n2301) );
  NOR U4302 ( .A(n2302), .B(n2301), .Z(n4880) );
  XOR U4303 ( .A(n2303), .B(b[434]), .Z(n4879) );
  NOR U4304 ( .A(n4880), .B(n4879), .Z(n2304) );
  NOR U4305 ( .A(n2305), .B(n2304), .Z(n4882) );
  XOR U4306 ( .A(n2306), .B(b[435]), .Z(n4881) );
  NOR U4307 ( .A(n4882), .B(n4881), .Z(n2307) );
  NOR U4308 ( .A(n2308), .B(n2307), .Z(n4884) );
  XOR U4309 ( .A(n2309), .B(b[436]), .Z(n4883) );
  NOR U4310 ( .A(n4884), .B(n4883), .Z(n2310) );
  NOR U4311 ( .A(n2311), .B(n2310), .Z(n4886) );
  XOR U4312 ( .A(n2312), .B(b[437]), .Z(n4885) );
  NOR U4313 ( .A(n4886), .B(n4885), .Z(n2313) );
  NOR U4314 ( .A(n2314), .B(n2313), .Z(n4888) );
  XOR U4315 ( .A(n2315), .B(b[438]), .Z(n4887) );
  NOR U4316 ( .A(n4888), .B(n4887), .Z(n2316) );
  NOR U4317 ( .A(n2317), .B(n2316), .Z(n4890) );
  XOR U4318 ( .A(n2318), .B(b[439]), .Z(n4889) );
  NOR U4319 ( .A(n4890), .B(n4889), .Z(n2319) );
  NOR U4320 ( .A(n2320), .B(n2319), .Z(n4894) );
  XOR U4321 ( .A(n2321), .B(b[440]), .Z(n4893) );
  NOR U4322 ( .A(n4894), .B(n4893), .Z(n2322) );
  NOR U4323 ( .A(n2323), .B(n2322), .Z(n4896) );
  XOR U4324 ( .A(n2324), .B(b[441]), .Z(n4895) );
  NOR U4325 ( .A(n4896), .B(n4895), .Z(n2325) );
  NOR U4326 ( .A(n2326), .B(n2325), .Z(n4898) );
  XOR U4327 ( .A(n2327), .B(b[442]), .Z(n4897) );
  NOR U4328 ( .A(n4898), .B(n4897), .Z(n2328) );
  NOR U4329 ( .A(n2329), .B(n2328), .Z(n4900) );
  XOR U4330 ( .A(n2330), .B(b[443]), .Z(n4899) );
  NOR U4331 ( .A(n4900), .B(n4899), .Z(n2331) );
  NOR U4332 ( .A(n2332), .B(n2331), .Z(n4902) );
  XOR U4333 ( .A(n2333), .B(b[444]), .Z(n4901) );
  NOR U4334 ( .A(n4902), .B(n4901), .Z(n2334) );
  NOR U4335 ( .A(n2335), .B(n2334), .Z(n4904) );
  XOR U4336 ( .A(n2336), .B(b[445]), .Z(n4903) );
  NOR U4337 ( .A(n4904), .B(n4903), .Z(n2337) );
  NOR U4338 ( .A(n2338), .B(n2337), .Z(n4906) );
  XOR U4339 ( .A(n2339), .B(b[446]), .Z(n4905) );
  NOR U4340 ( .A(n4906), .B(n4905), .Z(n2340) );
  NOR U4341 ( .A(n2341), .B(n2340), .Z(n4908) );
  XOR U4342 ( .A(n2342), .B(b[447]), .Z(n4907) );
  NOR U4343 ( .A(n4908), .B(n4907), .Z(n2343) );
  NOR U4344 ( .A(n2344), .B(n2343), .Z(n4910) );
  XOR U4345 ( .A(n2345), .B(b[448]), .Z(n4909) );
  NOR U4346 ( .A(n4910), .B(n4909), .Z(n2346) );
  NOR U4347 ( .A(n2347), .B(n2346), .Z(n4912) );
  XOR U4348 ( .A(n2348), .B(b[449]), .Z(n4911) );
  NOR U4349 ( .A(n4912), .B(n4911), .Z(n2349) );
  NOR U4350 ( .A(n2350), .B(n2349), .Z(n4916) );
  XOR U4351 ( .A(n2351), .B(b[450]), .Z(n4915) );
  NOR U4352 ( .A(n4916), .B(n4915), .Z(n2352) );
  NOR U4353 ( .A(n2353), .B(n2352), .Z(n4918) );
  XOR U4354 ( .A(n2354), .B(b[451]), .Z(n4917) );
  NOR U4355 ( .A(n4918), .B(n4917), .Z(n2355) );
  NOR U4356 ( .A(n2356), .B(n2355), .Z(n4920) );
  XOR U4357 ( .A(n2357), .B(b[452]), .Z(n4919) );
  NOR U4358 ( .A(n4920), .B(n4919), .Z(n2358) );
  NOR U4359 ( .A(n2359), .B(n2358), .Z(n4922) );
  XOR U4360 ( .A(n2360), .B(b[453]), .Z(n4921) );
  NOR U4361 ( .A(n4922), .B(n4921), .Z(n2361) );
  NOR U4362 ( .A(n2362), .B(n2361), .Z(n4924) );
  XOR U4363 ( .A(n2363), .B(b[454]), .Z(n4923) );
  NOR U4364 ( .A(n4924), .B(n4923), .Z(n2364) );
  NOR U4365 ( .A(n2365), .B(n2364), .Z(n4926) );
  XOR U4366 ( .A(n2366), .B(b[455]), .Z(n4925) );
  NOR U4367 ( .A(n4926), .B(n4925), .Z(n2367) );
  NOR U4368 ( .A(n2368), .B(n2367), .Z(n4928) );
  XOR U4369 ( .A(n2369), .B(b[456]), .Z(n4927) );
  NOR U4370 ( .A(n4928), .B(n4927), .Z(n2370) );
  NOR U4371 ( .A(n2371), .B(n2370), .Z(n4930) );
  XOR U4372 ( .A(n2372), .B(b[457]), .Z(n4929) );
  NOR U4373 ( .A(n4930), .B(n4929), .Z(n2373) );
  NOR U4374 ( .A(n2374), .B(n2373), .Z(n4932) );
  XOR U4375 ( .A(n2375), .B(b[458]), .Z(n4931) );
  NOR U4376 ( .A(n4932), .B(n4931), .Z(n2376) );
  NOR U4377 ( .A(n2377), .B(n2376), .Z(n4934) );
  XOR U4378 ( .A(n2378), .B(b[459]), .Z(n4933) );
  NOR U4379 ( .A(n4934), .B(n4933), .Z(n2379) );
  NOR U4380 ( .A(n2380), .B(n2379), .Z(n4938) );
  XOR U4381 ( .A(n2381), .B(b[460]), .Z(n4937) );
  NOR U4382 ( .A(n4938), .B(n4937), .Z(n2382) );
  NOR U4383 ( .A(n2383), .B(n2382), .Z(n4940) );
  XOR U4384 ( .A(n2384), .B(b[461]), .Z(n4939) );
  NOR U4385 ( .A(n4940), .B(n4939), .Z(n2385) );
  NOR U4386 ( .A(n2386), .B(n2385), .Z(n4942) );
  XOR U4387 ( .A(n2387), .B(b[462]), .Z(n4941) );
  NOR U4388 ( .A(n4942), .B(n4941), .Z(n2388) );
  NOR U4389 ( .A(n2389), .B(n2388), .Z(n4944) );
  XOR U4390 ( .A(n2390), .B(b[463]), .Z(n4943) );
  NOR U4391 ( .A(n4944), .B(n4943), .Z(n2391) );
  NOR U4392 ( .A(n2392), .B(n2391), .Z(n4946) );
  XOR U4393 ( .A(n2393), .B(b[464]), .Z(n4945) );
  NOR U4394 ( .A(n4946), .B(n4945), .Z(n2394) );
  NOR U4395 ( .A(n2395), .B(n2394), .Z(n4948) );
  XOR U4396 ( .A(n2396), .B(b[465]), .Z(n4947) );
  NOR U4397 ( .A(n4948), .B(n4947), .Z(n2397) );
  NOR U4398 ( .A(n2398), .B(n2397), .Z(n4950) );
  XOR U4399 ( .A(n2399), .B(b[466]), .Z(n4949) );
  NOR U4400 ( .A(n4950), .B(n4949), .Z(n2400) );
  NOR U4401 ( .A(n2401), .B(n2400), .Z(n4952) );
  XOR U4402 ( .A(n2402), .B(b[467]), .Z(n4951) );
  NOR U4403 ( .A(n4952), .B(n4951), .Z(n2403) );
  NOR U4404 ( .A(n2404), .B(n2403), .Z(n4954) );
  XOR U4405 ( .A(n2405), .B(b[468]), .Z(n4953) );
  NOR U4406 ( .A(n4954), .B(n4953), .Z(n2406) );
  NOR U4407 ( .A(n2407), .B(n2406), .Z(n4956) );
  XOR U4408 ( .A(n2408), .B(b[469]), .Z(n4955) );
  NOR U4409 ( .A(n4956), .B(n4955), .Z(n2409) );
  NOR U4410 ( .A(n2410), .B(n2409), .Z(n4960) );
  XOR U4411 ( .A(n2411), .B(b[470]), .Z(n4959) );
  NOR U4412 ( .A(n4960), .B(n4959), .Z(n2412) );
  NOR U4413 ( .A(n2413), .B(n2412), .Z(n4962) );
  XOR U4414 ( .A(n2414), .B(b[471]), .Z(n4961) );
  NOR U4415 ( .A(n4962), .B(n4961), .Z(n2415) );
  NOR U4416 ( .A(n2416), .B(n2415), .Z(n4964) );
  XOR U4417 ( .A(n2417), .B(b[472]), .Z(n4963) );
  NOR U4418 ( .A(n4964), .B(n4963), .Z(n2418) );
  NOR U4419 ( .A(n2419), .B(n2418), .Z(n4966) );
  XOR U4420 ( .A(n2420), .B(b[473]), .Z(n4965) );
  NOR U4421 ( .A(n4966), .B(n4965), .Z(n2421) );
  NOR U4422 ( .A(n2422), .B(n2421), .Z(n4968) );
  XOR U4423 ( .A(n2423), .B(b[474]), .Z(n4967) );
  NOR U4424 ( .A(n4968), .B(n4967), .Z(n2424) );
  NOR U4425 ( .A(n2425), .B(n2424), .Z(n4970) );
  XOR U4426 ( .A(n2426), .B(b[475]), .Z(n4969) );
  NOR U4427 ( .A(n4970), .B(n4969), .Z(n2427) );
  NOR U4428 ( .A(n2428), .B(n2427), .Z(n4972) );
  XOR U4429 ( .A(n2429), .B(b[476]), .Z(n4971) );
  NOR U4430 ( .A(n4972), .B(n4971), .Z(n2430) );
  NOR U4431 ( .A(n2431), .B(n2430), .Z(n4974) );
  XOR U4432 ( .A(n2432), .B(b[477]), .Z(n4973) );
  NOR U4433 ( .A(n4974), .B(n4973), .Z(n2433) );
  NOR U4434 ( .A(n2434), .B(n2433), .Z(n4976) );
  XOR U4435 ( .A(n2435), .B(b[478]), .Z(n4975) );
  NOR U4436 ( .A(n4976), .B(n4975), .Z(n2436) );
  NOR U4437 ( .A(n2437), .B(n2436), .Z(n4978) );
  XOR U4438 ( .A(n2438), .B(b[479]), .Z(n4977) );
  NOR U4439 ( .A(n4978), .B(n4977), .Z(n2439) );
  NOR U4440 ( .A(n2440), .B(n2439), .Z(n4982) );
  XOR U4441 ( .A(n2441), .B(b[480]), .Z(n4981) );
  NOR U4442 ( .A(n4982), .B(n4981), .Z(n2442) );
  NOR U4443 ( .A(n2443), .B(n2442), .Z(n4984) );
  XOR U4444 ( .A(n2444), .B(b[481]), .Z(n4983) );
  NOR U4445 ( .A(n4984), .B(n4983), .Z(n2445) );
  NOR U4446 ( .A(n2446), .B(n2445), .Z(n4986) );
  XOR U4447 ( .A(n2447), .B(b[482]), .Z(n4985) );
  NOR U4448 ( .A(n4986), .B(n4985), .Z(n2448) );
  NOR U4449 ( .A(n2449), .B(n2448), .Z(n4988) );
  XOR U4450 ( .A(n2450), .B(b[483]), .Z(n4987) );
  NOR U4451 ( .A(n4988), .B(n4987), .Z(n2451) );
  NOR U4452 ( .A(n2452), .B(n2451), .Z(n4990) );
  XOR U4453 ( .A(n2453), .B(b[484]), .Z(n4989) );
  NOR U4454 ( .A(n4990), .B(n4989), .Z(n2454) );
  NOR U4455 ( .A(n2455), .B(n2454), .Z(n4992) );
  XOR U4456 ( .A(n2456), .B(b[485]), .Z(n4991) );
  NOR U4457 ( .A(n4992), .B(n4991), .Z(n2457) );
  NOR U4458 ( .A(n2458), .B(n2457), .Z(n4994) );
  XOR U4459 ( .A(n2459), .B(b[486]), .Z(n4993) );
  NOR U4460 ( .A(n4994), .B(n4993), .Z(n2460) );
  NOR U4461 ( .A(n2461), .B(n2460), .Z(n4996) );
  XOR U4462 ( .A(n2462), .B(b[487]), .Z(n4995) );
  NOR U4463 ( .A(n4996), .B(n4995), .Z(n2463) );
  NOR U4464 ( .A(n2464), .B(n2463), .Z(n4998) );
  XOR U4465 ( .A(n2465), .B(b[488]), .Z(n4997) );
  NOR U4466 ( .A(n4998), .B(n4997), .Z(n2466) );
  NOR U4467 ( .A(n2467), .B(n2466), .Z(n5000) );
  XOR U4468 ( .A(n2468), .B(b[489]), .Z(n4999) );
  NOR U4469 ( .A(n5000), .B(n4999), .Z(n2469) );
  NOR U4470 ( .A(n2470), .B(n2469), .Z(n5004) );
  XOR U4471 ( .A(n2471), .B(b[490]), .Z(n5003) );
  NOR U4472 ( .A(n5004), .B(n5003), .Z(n2472) );
  NOR U4473 ( .A(n2473), .B(n2472), .Z(n5006) );
  XOR U4474 ( .A(n2474), .B(b[491]), .Z(n5005) );
  NOR U4475 ( .A(n5006), .B(n5005), .Z(n2475) );
  NOR U4476 ( .A(n2476), .B(n2475), .Z(n5008) );
  XOR U4477 ( .A(n2477), .B(b[492]), .Z(n5007) );
  NOR U4478 ( .A(n5008), .B(n5007), .Z(n2478) );
  NOR U4479 ( .A(n2479), .B(n2478), .Z(n5010) );
  XOR U4480 ( .A(n2480), .B(b[493]), .Z(n5009) );
  NOR U4481 ( .A(n5010), .B(n5009), .Z(n2481) );
  NOR U4482 ( .A(n2482), .B(n2481), .Z(n5012) );
  XOR U4483 ( .A(n2483), .B(b[494]), .Z(n5011) );
  NOR U4484 ( .A(n5012), .B(n5011), .Z(n2484) );
  NOR U4485 ( .A(n2485), .B(n2484), .Z(n5014) );
  XOR U4486 ( .A(n2486), .B(b[495]), .Z(n5013) );
  NOR U4487 ( .A(n5014), .B(n5013), .Z(n2487) );
  NOR U4488 ( .A(n2488), .B(n2487), .Z(n5016) );
  XOR U4489 ( .A(n2489), .B(b[496]), .Z(n5015) );
  NOR U4490 ( .A(n5016), .B(n5015), .Z(n2490) );
  NOR U4491 ( .A(n2491), .B(n2490), .Z(n5018) );
  XOR U4492 ( .A(n2492), .B(b[497]), .Z(n5017) );
  NOR U4493 ( .A(n5018), .B(n5017), .Z(n2493) );
  NOR U4494 ( .A(n2494), .B(n2493), .Z(n5020) );
  XOR U4495 ( .A(n2495), .B(b[498]), .Z(n5019) );
  NOR U4496 ( .A(n5020), .B(n5019), .Z(n2496) );
  NOR U4497 ( .A(n2497), .B(n2496), .Z(n5022) );
  XOR U4498 ( .A(n2498), .B(b[499]), .Z(n5021) );
  NOR U4499 ( .A(n5022), .B(n5021), .Z(n2499) );
  NOR U4500 ( .A(n2500), .B(n2499), .Z(n5028) );
  XOR U4501 ( .A(n2501), .B(b[500]), .Z(n5027) );
  NOR U4502 ( .A(n5028), .B(n5027), .Z(n2502) );
  NOR U4503 ( .A(n2503), .B(n2502), .Z(n5030) );
  XOR U4504 ( .A(n2504), .B(b[501]), .Z(n5029) );
  NOR U4505 ( .A(n5030), .B(n5029), .Z(n2505) );
  NOR U4506 ( .A(n2506), .B(n2505), .Z(n5032) );
  XOR U4507 ( .A(n2507), .B(b[502]), .Z(n5031) );
  NOR U4508 ( .A(n5032), .B(n5031), .Z(n2508) );
  NOR U4509 ( .A(n2509), .B(n2508), .Z(n5034) );
  XOR U4510 ( .A(n2510), .B(b[503]), .Z(n5033) );
  NOR U4511 ( .A(n5034), .B(n5033), .Z(n2511) );
  NOR U4512 ( .A(n2512), .B(n2511), .Z(n5036) );
  XOR U4513 ( .A(n2513), .B(b[504]), .Z(n5035) );
  NOR U4514 ( .A(n5036), .B(n5035), .Z(n2514) );
  NOR U4515 ( .A(n2515), .B(n2514), .Z(n5038) );
  XOR U4516 ( .A(n2516), .B(b[505]), .Z(n5037) );
  NOR U4517 ( .A(n5038), .B(n5037), .Z(n2517) );
  NOR U4518 ( .A(n2518), .B(n2517), .Z(n5040) );
  XOR U4519 ( .A(n2519), .B(b[506]), .Z(n5039) );
  NOR U4520 ( .A(n5040), .B(n5039), .Z(n2520) );
  NOR U4521 ( .A(n2521), .B(n2520), .Z(n5042) );
  XOR U4522 ( .A(n2522), .B(b[507]), .Z(n5041) );
  NOR U4523 ( .A(n5042), .B(n5041), .Z(n2523) );
  NOR U4524 ( .A(n2524), .B(n2523), .Z(n5044) );
  XOR U4525 ( .A(n2525), .B(b[508]), .Z(n5043) );
  NOR U4526 ( .A(n5044), .B(n5043), .Z(n2526) );
  NOR U4527 ( .A(n2527), .B(n2526), .Z(n5046) );
  XOR U4528 ( .A(n2528), .B(b[509]), .Z(n5045) );
  NOR U4529 ( .A(n5046), .B(n5045), .Z(n2529) );
  NOR U4530 ( .A(n2530), .B(n2529), .Z(n5050) );
  XOR U4531 ( .A(n2531), .B(b[510]), .Z(n5049) );
  NOR U4532 ( .A(n5050), .B(n5049), .Z(n2532) );
  NOR U4533 ( .A(n2533), .B(n2532), .Z(n5052) );
  XOR U4534 ( .A(n2534), .B(b[511]), .Z(n5051) );
  NOR U4535 ( .A(n5052), .B(n5051), .Z(n2535) );
  NOR U4536 ( .A(n2536), .B(n2535), .Z(n5054) );
  XOR U4537 ( .A(n2537), .B(b[512]), .Z(n5053) );
  NOR U4538 ( .A(n5054), .B(n5053), .Z(n2538) );
  NOR U4539 ( .A(n2539), .B(n2538), .Z(n5056) );
  XOR U4540 ( .A(n2540), .B(b[513]), .Z(n5055) );
  NOR U4541 ( .A(n5056), .B(n5055), .Z(n2541) );
  NOR U4542 ( .A(n2542), .B(n2541), .Z(n5058) );
  XOR U4543 ( .A(n2543), .B(b[514]), .Z(n5057) );
  NOR U4544 ( .A(n5058), .B(n5057), .Z(n2544) );
  NOR U4545 ( .A(n2545), .B(n2544), .Z(n5060) );
  XOR U4546 ( .A(n2546), .B(b[515]), .Z(n5059) );
  NOR U4547 ( .A(n5060), .B(n5059), .Z(n2547) );
  NOR U4548 ( .A(n2548), .B(n2547), .Z(n5062) );
  XOR U4549 ( .A(n2549), .B(b[516]), .Z(n5061) );
  NOR U4550 ( .A(n5062), .B(n5061), .Z(n2550) );
  NOR U4551 ( .A(n2551), .B(n2550), .Z(n5064) );
  XOR U4552 ( .A(n2552), .B(b[517]), .Z(n5063) );
  NOR U4553 ( .A(n5064), .B(n5063), .Z(n2553) );
  NOR U4554 ( .A(n2554), .B(n2553), .Z(n5066) );
  XOR U4555 ( .A(n2555), .B(b[518]), .Z(n5065) );
  NOR U4556 ( .A(n5066), .B(n5065), .Z(n2556) );
  NOR U4557 ( .A(n2557), .B(n2556), .Z(n5068) );
  XOR U4558 ( .A(n2558), .B(b[519]), .Z(n5067) );
  NOR U4559 ( .A(n5068), .B(n5067), .Z(n2559) );
  NOR U4560 ( .A(n2560), .B(n2559), .Z(n5072) );
  XOR U4561 ( .A(n2561), .B(b[520]), .Z(n5071) );
  NOR U4562 ( .A(n5072), .B(n5071), .Z(n2562) );
  NOR U4563 ( .A(n2563), .B(n2562), .Z(n5074) );
  XOR U4564 ( .A(n2564), .B(b[521]), .Z(n5073) );
  NOR U4565 ( .A(n5074), .B(n5073), .Z(n2565) );
  NOR U4566 ( .A(n2566), .B(n2565), .Z(n5076) );
  XOR U4567 ( .A(n2567), .B(b[522]), .Z(n5075) );
  NOR U4568 ( .A(n5076), .B(n5075), .Z(n2568) );
  NOR U4569 ( .A(n2569), .B(n2568), .Z(n5078) );
  XOR U4570 ( .A(n2570), .B(b[523]), .Z(n5077) );
  NOR U4571 ( .A(n5078), .B(n5077), .Z(n2571) );
  NOR U4572 ( .A(n2572), .B(n2571), .Z(n5080) );
  XOR U4573 ( .A(n2573), .B(b[524]), .Z(n5079) );
  NOR U4574 ( .A(n5080), .B(n5079), .Z(n2574) );
  NOR U4575 ( .A(n2575), .B(n2574), .Z(n5082) );
  XOR U4576 ( .A(n2576), .B(b[525]), .Z(n5081) );
  NOR U4577 ( .A(n5082), .B(n5081), .Z(n2577) );
  NOR U4578 ( .A(n2578), .B(n2577), .Z(n5084) );
  XOR U4579 ( .A(n2579), .B(b[526]), .Z(n5083) );
  NOR U4580 ( .A(n5084), .B(n5083), .Z(n2580) );
  NOR U4581 ( .A(n2581), .B(n2580), .Z(n5086) );
  XOR U4582 ( .A(n2582), .B(b[527]), .Z(n5085) );
  NOR U4583 ( .A(n5086), .B(n5085), .Z(n2583) );
  NOR U4584 ( .A(n2584), .B(n2583), .Z(n5088) );
  XOR U4585 ( .A(n2585), .B(b[528]), .Z(n5087) );
  NOR U4586 ( .A(n5088), .B(n5087), .Z(n2586) );
  NOR U4587 ( .A(n2587), .B(n2586), .Z(n5090) );
  XOR U4588 ( .A(n2588), .B(b[529]), .Z(n5089) );
  NOR U4589 ( .A(n5090), .B(n5089), .Z(n2589) );
  NOR U4590 ( .A(n2590), .B(n2589), .Z(n5094) );
  XOR U4591 ( .A(n2591), .B(b[530]), .Z(n5093) );
  NOR U4592 ( .A(n5094), .B(n5093), .Z(n2592) );
  NOR U4593 ( .A(n2593), .B(n2592), .Z(n5096) );
  XOR U4594 ( .A(n2594), .B(b[531]), .Z(n5095) );
  NOR U4595 ( .A(n5096), .B(n5095), .Z(n2595) );
  NOR U4596 ( .A(n2596), .B(n2595), .Z(n5098) );
  XOR U4597 ( .A(n2597), .B(b[532]), .Z(n5097) );
  NOR U4598 ( .A(n5098), .B(n5097), .Z(n2598) );
  NOR U4599 ( .A(n2599), .B(n2598), .Z(n5100) );
  XOR U4600 ( .A(n2600), .B(b[533]), .Z(n5099) );
  NOR U4601 ( .A(n5100), .B(n5099), .Z(n2601) );
  NOR U4602 ( .A(n2602), .B(n2601), .Z(n5102) );
  XOR U4603 ( .A(n2603), .B(b[534]), .Z(n5101) );
  NOR U4604 ( .A(n5102), .B(n5101), .Z(n2604) );
  NOR U4605 ( .A(n2605), .B(n2604), .Z(n5104) );
  XOR U4606 ( .A(n2606), .B(b[535]), .Z(n5103) );
  NOR U4607 ( .A(n5104), .B(n5103), .Z(n2607) );
  NOR U4608 ( .A(n2608), .B(n2607), .Z(n5106) );
  XOR U4609 ( .A(n2609), .B(b[536]), .Z(n5105) );
  NOR U4610 ( .A(n5106), .B(n5105), .Z(n2610) );
  NOR U4611 ( .A(n2611), .B(n2610), .Z(n5108) );
  XOR U4612 ( .A(n2612), .B(b[537]), .Z(n5107) );
  NOR U4613 ( .A(n5108), .B(n5107), .Z(n2613) );
  NOR U4614 ( .A(n2614), .B(n2613), .Z(n5110) );
  XOR U4615 ( .A(n2615), .B(b[538]), .Z(n5109) );
  NOR U4616 ( .A(n5110), .B(n5109), .Z(n2616) );
  NOR U4617 ( .A(n2617), .B(n2616), .Z(n5112) );
  XOR U4618 ( .A(n2618), .B(b[539]), .Z(n5111) );
  NOR U4619 ( .A(n5112), .B(n5111), .Z(n2619) );
  NOR U4620 ( .A(n2620), .B(n2619), .Z(n5116) );
  XOR U4621 ( .A(n2621), .B(b[540]), .Z(n5115) );
  NOR U4622 ( .A(n5116), .B(n5115), .Z(n2622) );
  NOR U4623 ( .A(n2623), .B(n2622), .Z(n5118) );
  XOR U4624 ( .A(n2624), .B(b[541]), .Z(n5117) );
  NOR U4625 ( .A(n5118), .B(n5117), .Z(n2625) );
  NOR U4626 ( .A(n2626), .B(n2625), .Z(n5120) );
  XOR U4627 ( .A(n2627), .B(b[542]), .Z(n5119) );
  NOR U4628 ( .A(n5120), .B(n5119), .Z(n2628) );
  NOR U4629 ( .A(n2629), .B(n2628), .Z(n5122) );
  XOR U4630 ( .A(n2630), .B(b[543]), .Z(n5121) );
  NOR U4631 ( .A(n5122), .B(n5121), .Z(n2631) );
  NOR U4632 ( .A(n2632), .B(n2631), .Z(n5124) );
  XOR U4633 ( .A(n2633), .B(b[544]), .Z(n5123) );
  NOR U4634 ( .A(n5124), .B(n5123), .Z(n2634) );
  NOR U4635 ( .A(n2635), .B(n2634), .Z(n5126) );
  XOR U4636 ( .A(n2636), .B(b[545]), .Z(n5125) );
  NOR U4637 ( .A(n5126), .B(n5125), .Z(n2637) );
  NOR U4638 ( .A(n2638), .B(n2637), .Z(n5128) );
  XOR U4639 ( .A(n2639), .B(b[546]), .Z(n5127) );
  NOR U4640 ( .A(n5128), .B(n5127), .Z(n2640) );
  NOR U4641 ( .A(n2641), .B(n2640), .Z(n5130) );
  XOR U4642 ( .A(n2642), .B(b[547]), .Z(n5129) );
  NOR U4643 ( .A(n5130), .B(n5129), .Z(n2643) );
  NOR U4644 ( .A(n2644), .B(n2643), .Z(n5132) );
  XOR U4645 ( .A(n2645), .B(b[548]), .Z(n5131) );
  NOR U4646 ( .A(n5132), .B(n5131), .Z(n2646) );
  NOR U4647 ( .A(n2647), .B(n2646), .Z(n5134) );
  XOR U4648 ( .A(n2648), .B(b[549]), .Z(n5133) );
  NOR U4649 ( .A(n5134), .B(n5133), .Z(n2649) );
  NOR U4650 ( .A(n2650), .B(n2649), .Z(n5138) );
  XOR U4651 ( .A(n2651), .B(b[550]), .Z(n5137) );
  NOR U4652 ( .A(n5138), .B(n5137), .Z(n2652) );
  NOR U4653 ( .A(n2653), .B(n2652), .Z(n5140) );
  XOR U4654 ( .A(n2654), .B(b[551]), .Z(n5139) );
  NOR U4655 ( .A(n5140), .B(n5139), .Z(n2655) );
  NOR U4656 ( .A(n2656), .B(n2655), .Z(n5142) );
  XOR U4657 ( .A(n2657), .B(b[552]), .Z(n5141) );
  NOR U4658 ( .A(n5142), .B(n5141), .Z(n2658) );
  NOR U4659 ( .A(n2659), .B(n2658), .Z(n5144) );
  XOR U4660 ( .A(n2660), .B(b[553]), .Z(n5143) );
  NOR U4661 ( .A(n5144), .B(n5143), .Z(n2661) );
  NOR U4662 ( .A(n2662), .B(n2661), .Z(n5146) );
  XOR U4663 ( .A(n2663), .B(b[554]), .Z(n5145) );
  NOR U4664 ( .A(n5146), .B(n5145), .Z(n2664) );
  NOR U4665 ( .A(n2665), .B(n2664), .Z(n5148) );
  XOR U4666 ( .A(n2666), .B(b[555]), .Z(n5147) );
  NOR U4667 ( .A(n5148), .B(n5147), .Z(n2667) );
  NOR U4668 ( .A(n2668), .B(n2667), .Z(n5150) );
  XOR U4669 ( .A(n2669), .B(b[556]), .Z(n5149) );
  NOR U4670 ( .A(n5150), .B(n5149), .Z(n2670) );
  NOR U4671 ( .A(n2671), .B(n2670), .Z(n5152) );
  XOR U4672 ( .A(n2672), .B(b[557]), .Z(n5151) );
  NOR U4673 ( .A(n5152), .B(n5151), .Z(n2673) );
  NOR U4674 ( .A(n2674), .B(n2673), .Z(n5154) );
  XOR U4675 ( .A(n2675), .B(b[558]), .Z(n5153) );
  NOR U4676 ( .A(n5154), .B(n5153), .Z(n2676) );
  NOR U4677 ( .A(n2677), .B(n2676), .Z(n5156) );
  XOR U4678 ( .A(n2678), .B(b[559]), .Z(n5155) );
  NOR U4679 ( .A(n5156), .B(n5155), .Z(n2679) );
  NOR U4680 ( .A(n2680), .B(n2679), .Z(n5160) );
  XOR U4681 ( .A(n2681), .B(b[560]), .Z(n5159) );
  NOR U4682 ( .A(n5160), .B(n5159), .Z(n2682) );
  NOR U4683 ( .A(n2683), .B(n2682), .Z(n5162) );
  XOR U4684 ( .A(n2684), .B(b[561]), .Z(n5161) );
  NOR U4685 ( .A(n5162), .B(n5161), .Z(n2685) );
  NOR U4686 ( .A(n2686), .B(n2685), .Z(n5164) );
  XOR U4687 ( .A(n2687), .B(b[562]), .Z(n5163) );
  NOR U4688 ( .A(n5164), .B(n5163), .Z(n2688) );
  NOR U4689 ( .A(n2689), .B(n2688), .Z(n5166) );
  XOR U4690 ( .A(n2690), .B(b[563]), .Z(n5165) );
  NOR U4691 ( .A(n5166), .B(n5165), .Z(n2691) );
  NOR U4692 ( .A(n2692), .B(n2691), .Z(n5168) );
  XOR U4693 ( .A(n2693), .B(b[564]), .Z(n5167) );
  NOR U4694 ( .A(n5168), .B(n5167), .Z(n2694) );
  NOR U4695 ( .A(n2695), .B(n2694), .Z(n5170) );
  XOR U4696 ( .A(n2696), .B(b[565]), .Z(n5169) );
  NOR U4697 ( .A(n5170), .B(n5169), .Z(n2697) );
  NOR U4698 ( .A(n2698), .B(n2697), .Z(n5172) );
  XOR U4699 ( .A(n2699), .B(b[566]), .Z(n5171) );
  NOR U4700 ( .A(n5172), .B(n5171), .Z(n2700) );
  NOR U4701 ( .A(n2701), .B(n2700), .Z(n5174) );
  XOR U4702 ( .A(n2702), .B(b[567]), .Z(n5173) );
  NOR U4703 ( .A(n5174), .B(n5173), .Z(n2703) );
  NOR U4704 ( .A(n2704), .B(n2703), .Z(n5176) );
  XOR U4705 ( .A(n2705), .B(b[568]), .Z(n5175) );
  NOR U4706 ( .A(n5176), .B(n5175), .Z(n2706) );
  NOR U4707 ( .A(n2707), .B(n2706), .Z(n5178) );
  XOR U4708 ( .A(n2708), .B(b[569]), .Z(n5177) );
  NOR U4709 ( .A(n5178), .B(n5177), .Z(n2709) );
  NOR U4710 ( .A(n2710), .B(n2709), .Z(n5182) );
  XOR U4711 ( .A(n2711), .B(b[570]), .Z(n5181) );
  NOR U4712 ( .A(n5182), .B(n5181), .Z(n2712) );
  NOR U4713 ( .A(n2713), .B(n2712), .Z(n5184) );
  XOR U4714 ( .A(n2714), .B(b[571]), .Z(n5183) );
  NOR U4715 ( .A(n5184), .B(n5183), .Z(n2715) );
  NOR U4716 ( .A(n2716), .B(n2715), .Z(n5186) );
  XOR U4717 ( .A(n2717), .B(b[572]), .Z(n5185) );
  NOR U4718 ( .A(n5186), .B(n5185), .Z(n2718) );
  NOR U4719 ( .A(n2719), .B(n2718), .Z(n5188) );
  XOR U4720 ( .A(n2720), .B(b[573]), .Z(n5187) );
  NOR U4721 ( .A(n5188), .B(n5187), .Z(n2721) );
  NOR U4722 ( .A(n2722), .B(n2721), .Z(n5190) );
  XOR U4723 ( .A(n2723), .B(b[574]), .Z(n5189) );
  NOR U4724 ( .A(n5190), .B(n5189), .Z(n2724) );
  NOR U4725 ( .A(n2725), .B(n2724), .Z(n5192) );
  XOR U4726 ( .A(n2726), .B(b[575]), .Z(n5191) );
  NOR U4727 ( .A(n5192), .B(n5191), .Z(n2727) );
  NOR U4728 ( .A(n2728), .B(n2727), .Z(n5194) );
  XOR U4729 ( .A(n2729), .B(b[576]), .Z(n5193) );
  NOR U4730 ( .A(n5194), .B(n5193), .Z(n2730) );
  NOR U4731 ( .A(n2731), .B(n2730), .Z(n5196) );
  XOR U4732 ( .A(n2732), .B(b[577]), .Z(n5195) );
  NOR U4733 ( .A(n5196), .B(n5195), .Z(n2733) );
  NOR U4734 ( .A(n2734), .B(n2733), .Z(n5198) );
  XOR U4735 ( .A(n2735), .B(b[578]), .Z(n5197) );
  NOR U4736 ( .A(n5198), .B(n5197), .Z(n2736) );
  NOR U4737 ( .A(n2737), .B(n2736), .Z(n5200) );
  XOR U4738 ( .A(n2738), .B(b[579]), .Z(n5199) );
  NOR U4739 ( .A(n5200), .B(n5199), .Z(n2739) );
  NOR U4740 ( .A(n2740), .B(n2739), .Z(n5204) );
  XOR U4741 ( .A(n2741), .B(b[580]), .Z(n5203) );
  NOR U4742 ( .A(n5204), .B(n5203), .Z(n2742) );
  NOR U4743 ( .A(n2743), .B(n2742), .Z(n5206) );
  XOR U4744 ( .A(n2744), .B(b[581]), .Z(n5205) );
  NOR U4745 ( .A(n5206), .B(n5205), .Z(n2745) );
  NOR U4746 ( .A(n2746), .B(n2745), .Z(n5208) );
  XOR U4747 ( .A(n2747), .B(b[582]), .Z(n5207) );
  NOR U4748 ( .A(n5208), .B(n5207), .Z(n2748) );
  NOR U4749 ( .A(n2749), .B(n2748), .Z(n5210) );
  XOR U4750 ( .A(n2750), .B(b[583]), .Z(n5209) );
  NOR U4751 ( .A(n5210), .B(n5209), .Z(n2751) );
  NOR U4752 ( .A(n2752), .B(n2751), .Z(n5212) );
  XOR U4753 ( .A(n2753), .B(b[584]), .Z(n5211) );
  NOR U4754 ( .A(n5212), .B(n5211), .Z(n2754) );
  NOR U4755 ( .A(n2755), .B(n2754), .Z(n5214) );
  XOR U4756 ( .A(n2756), .B(b[585]), .Z(n5213) );
  NOR U4757 ( .A(n5214), .B(n5213), .Z(n2757) );
  NOR U4758 ( .A(n2758), .B(n2757), .Z(n5216) );
  XOR U4759 ( .A(n2759), .B(b[586]), .Z(n5215) );
  NOR U4760 ( .A(n5216), .B(n5215), .Z(n2760) );
  NOR U4761 ( .A(n2761), .B(n2760), .Z(n5218) );
  XOR U4762 ( .A(n2762), .B(b[587]), .Z(n5217) );
  NOR U4763 ( .A(n5218), .B(n5217), .Z(n2763) );
  NOR U4764 ( .A(n2764), .B(n2763), .Z(n5220) );
  XOR U4765 ( .A(n2765), .B(b[588]), .Z(n5219) );
  NOR U4766 ( .A(n5220), .B(n5219), .Z(n2766) );
  NOR U4767 ( .A(n2767), .B(n2766), .Z(n5222) );
  XOR U4768 ( .A(n2768), .B(b[589]), .Z(n5221) );
  NOR U4769 ( .A(n5222), .B(n5221), .Z(n2769) );
  NOR U4770 ( .A(n2770), .B(n2769), .Z(n5226) );
  XOR U4771 ( .A(n2771), .B(b[590]), .Z(n5225) );
  NOR U4772 ( .A(n5226), .B(n5225), .Z(n2772) );
  NOR U4773 ( .A(n2773), .B(n2772), .Z(n5228) );
  XOR U4774 ( .A(n2774), .B(b[591]), .Z(n5227) );
  NOR U4775 ( .A(n5228), .B(n5227), .Z(n2775) );
  NOR U4776 ( .A(n2776), .B(n2775), .Z(n5230) );
  XOR U4777 ( .A(n2777), .B(b[592]), .Z(n5229) );
  NOR U4778 ( .A(n5230), .B(n5229), .Z(n2778) );
  NOR U4779 ( .A(n2779), .B(n2778), .Z(n5232) );
  XOR U4780 ( .A(n2780), .B(b[593]), .Z(n5231) );
  NOR U4781 ( .A(n5232), .B(n5231), .Z(n2781) );
  NOR U4782 ( .A(n2782), .B(n2781), .Z(n5234) );
  XOR U4783 ( .A(n2783), .B(b[594]), .Z(n5233) );
  NOR U4784 ( .A(n5234), .B(n5233), .Z(n2784) );
  NOR U4785 ( .A(n2785), .B(n2784), .Z(n5236) );
  XOR U4786 ( .A(n2786), .B(b[595]), .Z(n5235) );
  NOR U4787 ( .A(n5236), .B(n5235), .Z(n2787) );
  NOR U4788 ( .A(n2788), .B(n2787), .Z(n5238) );
  XOR U4789 ( .A(n2789), .B(b[596]), .Z(n5237) );
  NOR U4790 ( .A(n5238), .B(n5237), .Z(n2790) );
  NOR U4791 ( .A(n2791), .B(n2790), .Z(n5240) );
  XOR U4792 ( .A(n2792), .B(b[597]), .Z(n5239) );
  NOR U4793 ( .A(n5240), .B(n5239), .Z(n2793) );
  NOR U4794 ( .A(n2794), .B(n2793), .Z(n5242) );
  XOR U4795 ( .A(n2795), .B(b[598]), .Z(n5241) );
  NOR U4796 ( .A(n5242), .B(n5241), .Z(n2796) );
  NOR U4797 ( .A(n2797), .B(n2796), .Z(n5244) );
  XOR U4798 ( .A(n2798), .B(b[599]), .Z(n5243) );
  NOR U4799 ( .A(n5244), .B(n5243), .Z(n2799) );
  NOR U4800 ( .A(n2800), .B(n2799), .Z(n5250) );
  XOR U4801 ( .A(n2801), .B(b[600]), .Z(n5249) );
  NOR U4802 ( .A(n5250), .B(n5249), .Z(n2802) );
  NOR U4803 ( .A(n2803), .B(n2802), .Z(n5252) );
  XOR U4804 ( .A(n2804), .B(b[601]), .Z(n5251) );
  NOR U4805 ( .A(n5252), .B(n5251), .Z(n2805) );
  NOR U4806 ( .A(n2806), .B(n2805), .Z(n5254) );
  XOR U4807 ( .A(n2807), .B(b[602]), .Z(n5253) );
  NOR U4808 ( .A(n5254), .B(n5253), .Z(n2808) );
  NOR U4809 ( .A(n2809), .B(n2808), .Z(n5256) );
  XOR U4810 ( .A(n2810), .B(b[603]), .Z(n5255) );
  NOR U4811 ( .A(n5256), .B(n5255), .Z(n2811) );
  NOR U4812 ( .A(n2812), .B(n2811), .Z(n5258) );
  XOR U4813 ( .A(n2813), .B(b[604]), .Z(n5257) );
  NOR U4814 ( .A(n5258), .B(n5257), .Z(n2814) );
  NOR U4815 ( .A(n2815), .B(n2814), .Z(n5260) );
  XOR U4816 ( .A(n2816), .B(b[605]), .Z(n5259) );
  NOR U4817 ( .A(n5260), .B(n5259), .Z(n2817) );
  NOR U4818 ( .A(n2818), .B(n2817), .Z(n5262) );
  XOR U4819 ( .A(n2819), .B(b[606]), .Z(n5261) );
  NOR U4820 ( .A(n5262), .B(n5261), .Z(n2820) );
  NOR U4821 ( .A(n2821), .B(n2820), .Z(n5264) );
  XOR U4822 ( .A(n2822), .B(b[607]), .Z(n5263) );
  NOR U4823 ( .A(n5264), .B(n5263), .Z(n2823) );
  NOR U4824 ( .A(n2824), .B(n2823), .Z(n5266) );
  XOR U4825 ( .A(n2825), .B(b[608]), .Z(n5265) );
  NOR U4826 ( .A(n5266), .B(n5265), .Z(n2826) );
  NOR U4827 ( .A(n2827), .B(n2826), .Z(n5268) );
  XOR U4828 ( .A(n2828), .B(b[609]), .Z(n5267) );
  NOR U4829 ( .A(n5268), .B(n5267), .Z(n2829) );
  NOR U4830 ( .A(n2830), .B(n2829), .Z(n5272) );
  XOR U4831 ( .A(n2831), .B(b[610]), .Z(n5271) );
  NOR U4832 ( .A(n5272), .B(n5271), .Z(n2832) );
  NOR U4833 ( .A(n2833), .B(n2832), .Z(n5274) );
  XOR U4834 ( .A(n2834), .B(b[611]), .Z(n5273) );
  NOR U4835 ( .A(n5274), .B(n5273), .Z(n2835) );
  NOR U4836 ( .A(n2836), .B(n2835), .Z(n5276) );
  XOR U4837 ( .A(n2837), .B(b[612]), .Z(n5275) );
  NOR U4838 ( .A(n5276), .B(n5275), .Z(n2838) );
  NOR U4839 ( .A(n2839), .B(n2838), .Z(n5278) );
  XOR U4840 ( .A(n2840), .B(b[613]), .Z(n5277) );
  NOR U4841 ( .A(n5278), .B(n5277), .Z(n2841) );
  NOR U4842 ( .A(n2842), .B(n2841), .Z(n5280) );
  XOR U4843 ( .A(n2843), .B(b[614]), .Z(n5279) );
  NOR U4844 ( .A(n5280), .B(n5279), .Z(n2844) );
  NOR U4845 ( .A(n2845), .B(n2844), .Z(n5282) );
  XOR U4846 ( .A(n2846), .B(b[615]), .Z(n5281) );
  NOR U4847 ( .A(n5282), .B(n5281), .Z(n2847) );
  NOR U4848 ( .A(n2848), .B(n2847), .Z(n5284) );
  XOR U4849 ( .A(n2849), .B(b[616]), .Z(n5283) );
  NOR U4850 ( .A(n5284), .B(n5283), .Z(n2850) );
  NOR U4851 ( .A(n2851), .B(n2850), .Z(n5286) );
  XOR U4852 ( .A(n2852), .B(b[617]), .Z(n5285) );
  NOR U4853 ( .A(n5286), .B(n5285), .Z(n2853) );
  NOR U4854 ( .A(n2854), .B(n2853), .Z(n5288) );
  XOR U4855 ( .A(n2855), .B(b[618]), .Z(n5287) );
  NOR U4856 ( .A(n5288), .B(n5287), .Z(n2856) );
  NOR U4857 ( .A(n2857), .B(n2856), .Z(n5290) );
  XOR U4858 ( .A(n2858), .B(b[619]), .Z(n5289) );
  NOR U4859 ( .A(n5290), .B(n5289), .Z(n2859) );
  NOR U4860 ( .A(n2860), .B(n2859), .Z(n5294) );
  XOR U4861 ( .A(n2861), .B(b[620]), .Z(n5293) );
  NOR U4862 ( .A(n5294), .B(n5293), .Z(n2862) );
  NOR U4863 ( .A(n2863), .B(n2862), .Z(n5296) );
  XOR U4864 ( .A(n2864), .B(b[621]), .Z(n5295) );
  NOR U4865 ( .A(n5296), .B(n5295), .Z(n2865) );
  NOR U4866 ( .A(n2866), .B(n2865), .Z(n5298) );
  XOR U4867 ( .A(n2867), .B(b[622]), .Z(n5297) );
  NOR U4868 ( .A(n5298), .B(n5297), .Z(n2868) );
  NOR U4869 ( .A(n2869), .B(n2868), .Z(n5300) );
  XOR U4870 ( .A(n2870), .B(b[623]), .Z(n5299) );
  NOR U4871 ( .A(n5300), .B(n5299), .Z(n2871) );
  NOR U4872 ( .A(n2872), .B(n2871), .Z(n5302) );
  XOR U4873 ( .A(n2873), .B(b[624]), .Z(n5301) );
  NOR U4874 ( .A(n5302), .B(n5301), .Z(n2874) );
  NOR U4875 ( .A(n2875), .B(n2874), .Z(n5304) );
  XOR U4876 ( .A(n2876), .B(b[625]), .Z(n5303) );
  NOR U4877 ( .A(n5304), .B(n5303), .Z(n2877) );
  NOR U4878 ( .A(n2878), .B(n2877), .Z(n5306) );
  XOR U4879 ( .A(n2879), .B(b[626]), .Z(n5305) );
  NOR U4880 ( .A(n5306), .B(n5305), .Z(n2880) );
  NOR U4881 ( .A(n2881), .B(n2880), .Z(n5308) );
  XOR U4882 ( .A(n2882), .B(b[627]), .Z(n5307) );
  NOR U4883 ( .A(n5308), .B(n5307), .Z(n2883) );
  NOR U4884 ( .A(n2884), .B(n2883), .Z(n5310) );
  XOR U4885 ( .A(n2885), .B(b[628]), .Z(n5309) );
  NOR U4886 ( .A(n5310), .B(n5309), .Z(n2886) );
  NOR U4887 ( .A(n2887), .B(n2886), .Z(n5312) );
  XOR U4888 ( .A(n2888), .B(b[629]), .Z(n5311) );
  NOR U4889 ( .A(n5312), .B(n5311), .Z(n2889) );
  NOR U4890 ( .A(n2890), .B(n2889), .Z(n5316) );
  XOR U4891 ( .A(n2891), .B(b[630]), .Z(n5315) );
  NOR U4892 ( .A(n5316), .B(n5315), .Z(n2892) );
  NOR U4893 ( .A(n2893), .B(n2892), .Z(n5318) );
  XOR U4894 ( .A(n2894), .B(b[631]), .Z(n5317) );
  NOR U4895 ( .A(n5318), .B(n5317), .Z(n2895) );
  NOR U4896 ( .A(n2896), .B(n2895), .Z(n5320) );
  XOR U4897 ( .A(n2897), .B(b[632]), .Z(n5319) );
  NOR U4898 ( .A(n5320), .B(n5319), .Z(n2898) );
  NOR U4899 ( .A(n2899), .B(n2898), .Z(n5322) );
  XOR U4900 ( .A(n2900), .B(b[633]), .Z(n5321) );
  NOR U4901 ( .A(n5322), .B(n5321), .Z(n2901) );
  NOR U4902 ( .A(n2902), .B(n2901), .Z(n5324) );
  XOR U4903 ( .A(n2903), .B(b[634]), .Z(n5323) );
  NOR U4904 ( .A(n5324), .B(n5323), .Z(n2904) );
  NOR U4905 ( .A(n2905), .B(n2904), .Z(n5326) );
  XOR U4906 ( .A(n2906), .B(b[635]), .Z(n5325) );
  NOR U4907 ( .A(n5326), .B(n5325), .Z(n2907) );
  NOR U4908 ( .A(n2908), .B(n2907), .Z(n5328) );
  XOR U4909 ( .A(n2909), .B(b[636]), .Z(n5327) );
  NOR U4910 ( .A(n5328), .B(n5327), .Z(n2910) );
  NOR U4911 ( .A(n2911), .B(n2910), .Z(n5330) );
  XOR U4912 ( .A(n2912), .B(b[637]), .Z(n5329) );
  NOR U4913 ( .A(n5330), .B(n5329), .Z(n2913) );
  NOR U4914 ( .A(n2914), .B(n2913), .Z(n5332) );
  XOR U4915 ( .A(n2915), .B(b[638]), .Z(n5331) );
  NOR U4916 ( .A(n5332), .B(n5331), .Z(n2916) );
  NOR U4917 ( .A(n2917), .B(n2916), .Z(n5334) );
  XOR U4918 ( .A(n2918), .B(b[639]), .Z(n5333) );
  NOR U4919 ( .A(n5334), .B(n5333), .Z(n2919) );
  NOR U4920 ( .A(n2920), .B(n2919), .Z(n5338) );
  XOR U4921 ( .A(n2921), .B(b[640]), .Z(n5337) );
  NOR U4922 ( .A(n5338), .B(n5337), .Z(n2922) );
  NOR U4923 ( .A(n2923), .B(n2922), .Z(n5340) );
  XOR U4924 ( .A(n2924), .B(b[641]), .Z(n5339) );
  NOR U4925 ( .A(n5340), .B(n5339), .Z(n2925) );
  NOR U4926 ( .A(n2926), .B(n2925), .Z(n5342) );
  XOR U4927 ( .A(n2927), .B(b[642]), .Z(n5341) );
  NOR U4928 ( .A(n5342), .B(n5341), .Z(n2928) );
  NOR U4929 ( .A(n2929), .B(n2928), .Z(n5344) );
  XOR U4930 ( .A(n2930), .B(b[643]), .Z(n5343) );
  NOR U4931 ( .A(n5344), .B(n5343), .Z(n2931) );
  NOR U4932 ( .A(n2932), .B(n2931), .Z(n5346) );
  XOR U4933 ( .A(n2933), .B(b[644]), .Z(n5345) );
  NOR U4934 ( .A(n5346), .B(n5345), .Z(n2934) );
  NOR U4935 ( .A(n2935), .B(n2934), .Z(n5348) );
  XOR U4936 ( .A(n2936), .B(b[645]), .Z(n5347) );
  NOR U4937 ( .A(n5348), .B(n5347), .Z(n2937) );
  NOR U4938 ( .A(n2938), .B(n2937), .Z(n5350) );
  XOR U4939 ( .A(n2939), .B(b[646]), .Z(n5349) );
  NOR U4940 ( .A(n5350), .B(n5349), .Z(n2940) );
  NOR U4941 ( .A(n2941), .B(n2940), .Z(n5352) );
  XOR U4942 ( .A(n2942), .B(b[647]), .Z(n5351) );
  NOR U4943 ( .A(n5352), .B(n5351), .Z(n2943) );
  NOR U4944 ( .A(n2944), .B(n2943), .Z(n5354) );
  XOR U4945 ( .A(n2945), .B(b[648]), .Z(n5353) );
  NOR U4946 ( .A(n5354), .B(n5353), .Z(n2946) );
  NOR U4947 ( .A(n2947), .B(n2946), .Z(n5356) );
  XOR U4948 ( .A(n2948), .B(b[649]), .Z(n5355) );
  NOR U4949 ( .A(n5356), .B(n5355), .Z(n2949) );
  NOR U4950 ( .A(n2950), .B(n2949), .Z(n5360) );
  XOR U4951 ( .A(n2951), .B(b[650]), .Z(n5359) );
  NOR U4952 ( .A(n5360), .B(n5359), .Z(n2952) );
  NOR U4953 ( .A(n2953), .B(n2952), .Z(n5362) );
  XOR U4954 ( .A(n2954), .B(b[651]), .Z(n5361) );
  NOR U4955 ( .A(n5362), .B(n5361), .Z(n2955) );
  NOR U4956 ( .A(n2956), .B(n2955), .Z(n5364) );
  XOR U4957 ( .A(n2957), .B(b[652]), .Z(n5363) );
  NOR U4958 ( .A(n5364), .B(n5363), .Z(n2958) );
  NOR U4959 ( .A(n2959), .B(n2958), .Z(n5366) );
  XOR U4960 ( .A(n2960), .B(b[653]), .Z(n5365) );
  NOR U4961 ( .A(n5366), .B(n5365), .Z(n2961) );
  NOR U4962 ( .A(n2962), .B(n2961), .Z(n5368) );
  XOR U4963 ( .A(n2963), .B(b[654]), .Z(n5367) );
  NOR U4964 ( .A(n5368), .B(n5367), .Z(n2964) );
  NOR U4965 ( .A(n2965), .B(n2964), .Z(n5370) );
  XOR U4966 ( .A(n2966), .B(b[655]), .Z(n5369) );
  NOR U4967 ( .A(n5370), .B(n5369), .Z(n2967) );
  NOR U4968 ( .A(n2968), .B(n2967), .Z(n5372) );
  XOR U4969 ( .A(n2969), .B(b[656]), .Z(n5371) );
  NOR U4970 ( .A(n5372), .B(n5371), .Z(n2970) );
  NOR U4971 ( .A(n2971), .B(n2970), .Z(n5374) );
  XOR U4972 ( .A(n2972), .B(b[657]), .Z(n5373) );
  NOR U4973 ( .A(n5374), .B(n5373), .Z(n2973) );
  NOR U4974 ( .A(n2974), .B(n2973), .Z(n5376) );
  XOR U4975 ( .A(n2975), .B(b[658]), .Z(n5375) );
  NOR U4976 ( .A(n5376), .B(n5375), .Z(n2976) );
  NOR U4977 ( .A(n2977), .B(n2976), .Z(n5378) );
  XOR U4978 ( .A(n2978), .B(b[659]), .Z(n5377) );
  NOR U4979 ( .A(n5378), .B(n5377), .Z(n2979) );
  NOR U4980 ( .A(n2980), .B(n2979), .Z(n5382) );
  XOR U4981 ( .A(n2981), .B(b[660]), .Z(n5381) );
  NOR U4982 ( .A(n5382), .B(n5381), .Z(n2982) );
  NOR U4983 ( .A(n2983), .B(n2982), .Z(n5384) );
  XOR U4984 ( .A(n2984), .B(b[661]), .Z(n5383) );
  NOR U4985 ( .A(n5384), .B(n5383), .Z(n2985) );
  NOR U4986 ( .A(n2986), .B(n2985), .Z(n5386) );
  XOR U4987 ( .A(n2987), .B(b[662]), .Z(n5385) );
  NOR U4988 ( .A(n5386), .B(n5385), .Z(n2988) );
  NOR U4989 ( .A(n2989), .B(n2988), .Z(n5388) );
  XOR U4990 ( .A(n2990), .B(b[663]), .Z(n5387) );
  NOR U4991 ( .A(n5388), .B(n5387), .Z(n2991) );
  NOR U4992 ( .A(n2992), .B(n2991), .Z(n5390) );
  XOR U4993 ( .A(n2993), .B(b[664]), .Z(n5389) );
  NOR U4994 ( .A(n5390), .B(n5389), .Z(n2994) );
  NOR U4995 ( .A(n2995), .B(n2994), .Z(n5392) );
  XOR U4996 ( .A(n2996), .B(b[665]), .Z(n5391) );
  NOR U4997 ( .A(n5392), .B(n5391), .Z(n2997) );
  NOR U4998 ( .A(n2998), .B(n2997), .Z(n5394) );
  XOR U4999 ( .A(n2999), .B(b[666]), .Z(n5393) );
  NOR U5000 ( .A(n5394), .B(n5393), .Z(n3000) );
  NOR U5001 ( .A(n3001), .B(n3000), .Z(n5396) );
  XOR U5002 ( .A(n3002), .B(b[667]), .Z(n5395) );
  NOR U5003 ( .A(n5396), .B(n5395), .Z(n3003) );
  NOR U5004 ( .A(n3004), .B(n3003), .Z(n5398) );
  XOR U5005 ( .A(n3005), .B(b[668]), .Z(n5397) );
  NOR U5006 ( .A(n5398), .B(n5397), .Z(n3006) );
  NOR U5007 ( .A(n3007), .B(n3006), .Z(n5400) );
  XOR U5008 ( .A(n3008), .B(b[669]), .Z(n5399) );
  NOR U5009 ( .A(n5400), .B(n5399), .Z(n3009) );
  NOR U5010 ( .A(n3010), .B(n3009), .Z(n5404) );
  XOR U5011 ( .A(n3011), .B(b[670]), .Z(n5403) );
  NOR U5012 ( .A(n5404), .B(n5403), .Z(n3012) );
  NOR U5013 ( .A(n3013), .B(n3012), .Z(n5406) );
  XOR U5014 ( .A(n3014), .B(b[671]), .Z(n5405) );
  NOR U5015 ( .A(n5406), .B(n5405), .Z(n3015) );
  NOR U5016 ( .A(n3016), .B(n3015), .Z(n5408) );
  XOR U5017 ( .A(n3017), .B(b[672]), .Z(n5407) );
  NOR U5018 ( .A(n5408), .B(n5407), .Z(n3018) );
  NOR U5019 ( .A(n3019), .B(n3018), .Z(n5410) );
  XOR U5020 ( .A(n3020), .B(b[673]), .Z(n5409) );
  NOR U5021 ( .A(n5410), .B(n5409), .Z(n3021) );
  NOR U5022 ( .A(n3022), .B(n3021), .Z(n5412) );
  XOR U5023 ( .A(n3023), .B(b[674]), .Z(n5411) );
  NOR U5024 ( .A(n5412), .B(n5411), .Z(n3024) );
  NOR U5025 ( .A(n3025), .B(n3024), .Z(n5414) );
  XOR U5026 ( .A(n3026), .B(b[675]), .Z(n5413) );
  NOR U5027 ( .A(n5414), .B(n5413), .Z(n3027) );
  NOR U5028 ( .A(n3028), .B(n3027), .Z(n5416) );
  XOR U5029 ( .A(n3029), .B(b[676]), .Z(n5415) );
  NOR U5030 ( .A(n5416), .B(n5415), .Z(n3030) );
  NOR U5031 ( .A(n3031), .B(n3030), .Z(n5418) );
  XOR U5032 ( .A(n3032), .B(b[677]), .Z(n5417) );
  NOR U5033 ( .A(n5418), .B(n5417), .Z(n3033) );
  NOR U5034 ( .A(n3034), .B(n3033), .Z(n5420) );
  XOR U5035 ( .A(n3035), .B(b[678]), .Z(n5419) );
  NOR U5036 ( .A(n5420), .B(n5419), .Z(n3036) );
  NOR U5037 ( .A(n3037), .B(n3036), .Z(n5422) );
  XOR U5038 ( .A(n3038), .B(b[679]), .Z(n5421) );
  NOR U5039 ( .A(n5422), .B(n5421), .Z(n3039) );
  NOR U5040 ( .A(n3040), .B(n3039), .Z(n5426) );
  XOR U5041 ( .A(n3041), .B(b[680]), .Z(n5425) );
  NOR U5042 ( .A(n5426), .B(n5425), .Z(n3042) );
  NOR U5043 ( .A(n3043), .B(n3042), .Z(n5428) );
  XOR U5044 ( .A(n3044), .B(b[681]), .Z(n5427) );
  NOR U5045 ( .A(n5428), .B(n5427), .Z(n3045) );
  NOR U5046 ( .A(n3046), .B(n3045), .Z(n5430) );
  XOR U5047 ( .A(n3047), .B(b[682]), .Z(n5429) );
  NOR U5048 ( .A(n5430), .B(n5429), .Z(n3048) );
  NOR U5049 ( .A(n3049), .B(n3048), .Z(n5432) );
  XOR U5050 ( .A(n3050), .B(b[683]), .Z(n5431) );
  NOR U5051 ( .A(n5432), .B(n5431), .Z(n3051) );
  NOR U5052 ( .A(n3052), .B(n3051), .Z(n5434) );
  XOR U5053 ( .A(n3053), .B(b[684]), .Z(n5433) );
  NOR U5054 ( .A(n5434), .B(n5433), .Z(n3054) );
  NOR U5055 ( .A(n3055), .B(n3054), .Z(n5436) );
  XOR U5056 ( .A(n3056), .B(b[685]), .Z(n5435) );
  NOR U5057 ( .A(n5436), .B(n5435), .Z(n3057) );
  NOR U5058 ( .A(n3058), .B(n3057), .Z(n5438) );
  XOR U5059 ( .A(n3059), .B(b[686]), .Z(n5437) );
  NOR U5060 ( .A(n5438), .B(n5437), .Z(n3060) );
  NOR U5061 ( .A(n3061), .B(n3060), .Z(n5440) );
  XOR U5062 ( .A(n3062), .B(b[687]), .Z(n5439) );
  NOR U5063 ( .A(n5440), .B(n5439), .Z(n3063) );
  NOR U5064 ( .A(n3064), .B(n3063), .Z(n5442) );
  XOR U5065 ( .A(n3065), .B(b[688]), .Z(n5441) );
  NOR U5066 ( .A(n5442), .B(n5441), .Z(n3066) );
  NOR U5067 ( .A(n3067), .B(n3066), .Z(n5444) );
  XOR U5068 ( .A(n3068), .B(b[689]), .Z(n5443) );
  NOR U5069 ( .A(n5444), .B(n5443), .Z(n3069) );
  NOR U5070 ( .A(n3070), .B(n3069), .Z(n5448) );
  XOR U5071 ( .A(n3071), .B(b[690]), .Z(n5447) );
  NOR U5072 ( .A(n5448), .B(n5447), .Z(n3072) );
  NOR U5073 ( .A(n3073), .B(n3072), .Z(n5450) );
  XOR U5074 ( .A(n3074), .B(b[691]), .Z(n5449) );
  NOR U5075 ( .A(n5450), .B(n5449), .Z(n3075) );
  NOR U5076 ( .A(n3076), .B(n3075), .Z(n5452) );
  XOR U5077 ( .A(n3077), .B(b[692]), .Z(n5451) );
  NOR U5078 ( .A(n5452), .B(n5451), .Z(n3078) );
  NOR U5079 ( .A(n3079), .B(n3078), .Z(n5454) );
  XOR U5080 ( .A(n3080), .B(b[693]), .Z(n5453) );
  NOR U5081 ( .A(n5454), .B(n5453), .Z(n3081) );
  NOR U5082 ( .A(n3082), .B(n3081), .Z(n5456) );
  XOR U5083 ( .A(n3083), .B(b[694]), .Z(n5455) );
  NOR U5084 ( .A(n5456), .B(n5455), .Z(n3084) );
  NOR U5085 ( .A(n3085), .B(n3084), .Z(n5458) );
  XOR U5086 ( .A(n3086), .B(b[695]), .Z(n5457) );
  NOR U5087 ( .A(n5458), .B(n5457), .Z(n3087) );
  NOR U5088 ( .A(n3088), .B(n3087), .Z(n5460) );
  XOR U5089 ( .A(n3089), .B(b[696]), .Z(n5459) );
  NOR U5090 ( .A(n5460), .B(n5459), .Z(n3090) );
  NOR U5091 ( .A(n3091), .B(n3090), .Z(n5462) );
  XOR U5092 ( .A(n3092), .B(b[697]), .Z(n5461) );
  NOR U5093 ( .A(n5462), .B(n5461), .Z(n3093) );
  NOR U5094 ( .A(n3094), .B(n3093), .Z(n5464) );
  XOR U5095 ( .A(n3095), .B(b[698]), .Z(n5463) );
  NOR U5096 ( .A(n5464), .B(n5463), .Z(n3096) );
  NOR U5097 ( .A(n3097), .B(n3096), .Z(n5466) );
  XOR U5098 ( .A(n3098), .B(b[699]), .Z(n5465) );
  NOR U5099 ( .A(n5466), .B(n5465), .Z(n3099) );
  NOR U5100 ( .A(n3100), .B(n3099), .Z(n5472) );
  XOR U5101 ( .A(n3101), .B(b[700]), .Z(n5471) );
  NOR U5102 ( .A(n5472), .B(n5471), .Z(n3102) );
  NOR U5103 ( .A(n3103), .B(n3102), .Z(n5474) );
  XOR U5104 ( .A(n3104), .B(b[701]), .Z(n5473) );
  NOR U5105 ( .A(n5474), .B(n5473), .Z(n3105) );
  NOR U5106 ( .A(n3106), .B(n3105), .Z(n5476) );
  XOR U5107 ( .A(n3107), .B(b[702]), .Z(n5475) );
  NOR U5108 ( .A(n5476), .B(n5475), .Z(n3108) );
  NOR U5109 ( .A(n3109), .B(n3108), .Z(n5478) );
  XOR U5110 ( .A(n3110), .B(b[703]), .Z(n5477) );
  NOR U5111 ( .A(n5478), .B(n5477), .Z(n3111) );
  NOR U5112 ( .A(n3112), .B(n3111), .Z(n5480) );
  XOR U5113 ( .A(n3113), .B(b[704]), .Z(n5479) );
  NOR U5114 ( .A(n5480), .B(n5479), .Z(n3114) );
  NOR U5115 ( .A(n3115), .B(n3114), .Z(n5482) );
  XOR U5116 ( .A(n3116), .B(b[705]), .Z(n5481) );
  NOR U5117 ( .A(n5482), .B(n5481), .Z(n3117) );
  NOR U5118 ( .A(n3118), .B(n3117), .Z(n5484) );
  XOR U5119 ( .A(n3119), .B(b[706]), .Z(n5483) );
  NOR U5120 ( .A(n5484), .B(n5483), .Z(n3120) );
  NOR U5121 ( .A(n3121), .B(n3120), .Z(n5486) );
  XOR U5122 ( .A(n3122), .B(b[707]), .Z(n5485) );
  NOR U5123 ( .A(n5486), .B(n5485), .Z(n3123) );
  NOR U5124 ( .A(n3124), .B(n3123), .Z(n5488) );
  XOR U5125 ( .A(n3125), .B(b[708]), .Z(n5487) );
  NOR U5126 ( .A(n5488), .B(n5487), .Z(n3126) );
  NOR U5127 ( .A(n3127), .B(n3126), .Z(n5490) );
  XOR U5128 ( .A(n3128), .B(b[709]), .Z(n5489) );
  NOR U5129 ( .A(n5490), .B(n5489), .Z(n3129) );
  NOR U5130 ( .A(n3130), .B(n3129), .Z(n5494) );
  XOR U5131 ( .A(n3131), .B(b[710]), .Z(n5493) );
  NOR U5132 ( .A(n5494), .B(n5493), .Z(n3132) );
  NOR U5133 ( .A(n3133), .B(n3132), .Z(n5496) );
  XOR U5134 ( .A(n3134), .B(b[711]), .Z(n5495) );
  NOR U5135 ( .A(n5496), .B(n5495), .Z(n3135) );
  NOR U5136 ( .A(n3136), .B(n3135), .Z(n5498) );
  XOR U5137 ( .A(n3137), .B(b[712]), .Z(n5497) );
  NOR U5138 ( .A(n5498), .B(n5497), .Z(n3138) );
  NOR U5139 ( .A(n3139), .B(n3138), .Z(n5500) );
  XOR U5140 ( .A(n3140), .B(b[713]), .Z(n5499) );
  NOR U5141 ( .A(n5500), .B(n5499), .Z(n3141) );
  NOR U5142 ( .A(n3142), .B(n3141), .Z(n5502) );
  XOR U5143 ( .A(n3143), .B(b[714]), .Z(n5501) );
  NOR U5144 ( .A(n5502), .B(n5501), .Z(n3144) );
  NOR U5145 ( .A(n3145), .B(n3144), .Z(n5504) );
  XOR U5146 ( .A(n3146), .B(b[715]), .Z(n5503) );
  NOR U5147 ( .A(n5504), .B(n5503), .Z(n3147) );
  NOR U5148 ( .A(n3148), .B(n3147), .Z(n5506) );
  XOR U5149 ( .A(n3149), .B(b[716]), .Z(n5505) );
  NOR U5150 ( .A(n5506), .B(n5505), .Z(n3150) );
  NOR U5151 ( .A(n3151), .B(n3150), .Z(n5508) );
  XOR U5152 ( .A(n3152), .B(b[717]), .Z(n5507) );
  NOR U5153 ( .A(n5508), .B(n5507), .Z(n3153) );
  NOR U5154 ( .A(n3154), .B(n3153), .Z(n5510) );
  XOR U5155 ( .A(n3155), .B(b[718]), .Z(n5509) );
  NOR U5156 ( .A(n5510), .B(n5509), .Z(n3156) );
  NOR U5157 ( .A(n3157), .B(n3156), .Z(n5512) );
  XOR U5158 ( .A(n3158), .B(b[719]), .Z(n5511) );
  NOR U5159 ( .A(n5512), .B(n5511), .Z(n3159) );
  NOR U5160 ( .A(n3160), .B(n3159), .Z(n5516) );
  XOR U5161 ( .A(n3161), .B(b[720]), .Z(n5515) );
  NOR U5162 ( .A(n5516), .B(n5515), .Z(n3162) );
  NOR U5163 ( .A(n3163), .B(n3162), .Z(n5518) );
  XOR U5164 ( .A(n3164), .B(b[721]), .Z(n5517) );
  NOR U5165 ( .A(n5518), .B(n5517), .Z(n3165) );
  NOR U5166 ( .A(n3166), .B(n3165), .Z(n5520) );
  XOR U5167 ( .A(n3167), .B(b[722]), .Z(n5519) );
  NOR U5168 ( .A(n5520), .B(n5519), .Z(n3168) );
  NOR U5169 ( .A(n3169), .B(n3168), .Z(n5522) );
  XOR U5170 ( .A(n3170), .B(b[723]), .Z(n5521) );
  NOR U5171 ( .A(n5522), .B(n5521), .Z(n3171) );
  NOR U5172 ( .A(n3172), .B(n3171), .Z(n5524) );
  XOR U5173 ( .A(n3173), .B(b[724]), .Z(n5523) );
  NOR U5174 ( .A(n5524), .B(n5523), .Z(n3174) );
  NOR U5175 ( .A(n3175), .B(n3174), .Z(n5526) );
  XOR U5176 ( .A(n3176), .B(b[725]), .Z(n5525) );
  NOR U5177 ( .A(n5526), .B(n5525), .Z(n3177) );
  NOR U5178 ( .A(n3178), .B(n3177), .Z(n5528) );
  XOR U5179 ( .A(n3179), .B(b[726]), .Z(n5527) );
  NOR U5180 ( .A(n5528), .B(n5527), .Z(n3180) );
  NOR U5181 ( .A(n3181), .B(n3180), .Z(n5530) );
  XOR U5182 ( .A(n3182), .B(b[727]), .Z(n5529) );
  NOR U5183 ( .A(n5530), .B(n5529), .Z(n3183) );
  NOR U5184 ( .A(n3184), .B(n3183), .Z(n5532) );
  XOR U5185 ( .A(n3185), .B(b[728]), .Z(n5531) );
  NOR U5186 ( .A(n5532), .B(n5531), .Z(n3186) );
  NOR U5187 ( .A(n3187), .B(n3186), .Z(n5534) );
  XOR U5188 ( .A(n3188), .B(b[729]), .Z(n5533) );
  NOR U5189 ( .A(n5534), .B(n5533), .Z(n3189) );
  NOR U5190 ( .A(n3190), .B(n3189), .Z(n5538) );
  XOR U5191 ( .A(n3191), .B(b[730]), .Z(n5537) );
  NOR U5192 ( .A(n5538), .B(n5537), .Z(n3192) );
  NOR U5193 ( .A(n3193), .B(n3192), .Z(n5540) );
  XOR U5194 ( .A(n3194), .B(b[731]), .Z(n5539) );
  NOR U5195 ( .A(n5540), .B(n5539), .Z(n3195) );
  NOR U5196 ( .A(n3196), .B(n3195), .Z(n5542) );
  XOR U5197 ( .A(n3197), .B(b[732]), .Z(n5541) );
  NOR U5198 ( .A(n5542), .B(n5541), .Z(n3198) );
  NOR U5199 ( .A(n3199), .B(n3198), .Z(n5544) );
  XOR U5200 ( .A(n3200), .B(b[733]), .Z(n5543) );
  NOR U5201 ( .A(n5544), .B(n5543), .Z(n3201) );
  NOR U5202 ( .A(n3202), .B(n3201), .Z(n5546) );
  XOR U5203 ( .A(n3203), .B(b[734]), .Z(n5545) );
  NOR U5204 ( .A(n5546), .B(n5545), .Z(n3204) );
  NOR U5205 ( .A(n3205), .B(n3204), .Z(n5548) );
  XOR U5206 ( .A(n3206), .B(b[735]), .Z(n5547) );
  NOR U5207 ( .A(n5548), .B(n5547), .Z(n3207) );
  NOR U5208 ( .A(n3208), .B(n3207), .Z(n5550) );
  XOR U5209 ( .A(n3209), .B(b[736]), .Z(n5549) );
  NOR U5210 ( .A(n5550), .B(n5549), .Z(n3210) );
  NOR U5211 ( .A(n3211), .B(n3210), .Z(n5552) );
  XOR U5212 ( .A(n3212), .B(b[737]), .Z(n5551) );
  NOR U5213 ( .A(n5552), .B(n5551), .Z(n3213) );
  NOR U5214 ( .A(n3214), .B(n3213), .Z(n5554) );
  XOR U5215 ( .A(n3215), .B(b[738]), .Z(n5553) );
  NOR U5216 ( .A(n5554), .B(n5553), .Z(n3216) );
  NOR U5217 ( .A(n3217), .B(n3216), .Z(n5556) );
  XOR U5218 ( .A(n3218), .B(b[739]), .Z(n5555) );
  NOR U5219 ( .A(n5556), .B(n5555), .Z(n3219) );
  NOR U5220 ( .A(n3220), .B(n3219), .Z(n5560) );
  XOR U5221 ( .A(n3221), .B(b[740]), .Z(n5559) );
  NOR U5222 ( .A(n5560), .B(n5559), .Z(n3222) );
  NOR U5223 ( .A(n3223), .B(n3222), .Z(n5562) );
  XOR U5224 ( .A(n3224), .B(b[741]), .Z(n5561) );
  NOR U5225 ( .A(n5562), .B(n5561), .Z(n3225) );
  NOR U5226 ( .A(n3226), .B(n3225), .Z(n5564) );
  XOR U5227 ( .A(n3227), .B(b[742]), .Z(n5563) );
  NOR U5228 ( .A(n5564), .B(n5563), .Z(n3228) );
  NOR U5229 ( .A(n3229), .B(n3228), .Z(n5566) );
  XOR U5230 ( .A(n3230), .B(b[743]), .Z(n5565) );
  NOR U5231 ( .A(n5566), .B(n5565), .Z(n3231) );
  NOR U5232 ( .A(n3232), .B(n3231), .Z(n5568) );
  XOR U5233 ( .A(n3233), .B(b[744]), .Z(n5567) );
  NOR U5234 ( .A(n5568), .B(n5567), .Z(n3234) );
  NOR U5235 ( .A(n3235), .B(n3234), .Z(n5570) );
  XOR U5236 ( .A(n3236), .B(b[745]), .Z(n5569) );
  NOR U5237 ( .A(n5570), .B(n5569), .Z(n3237) );
  NOR U5238 ( .A(n3238), .B(n3237), .Z(n5572) );
  XOR U5239 ( .A(n3239), .B(b[746]), .Z(n5571) );
  NOR U5240 ( .A(n5572), .B(n5571), .Z(n3240) );
  NOR U5241 ( .A(n3241), .B(n3240), .Z(n5574) );
  XOR U5242 ( .A(n3242), .B(b[747]), .Z(n5573) );
  NOR U5243 ( .A(n5574), .B(n5573), .Z(n3243) );
  NOR U5244 ( .A(n3244), .B(n3243), .Z(n5576) );
  XOR U5245 ( .A(n3245), .B(b[748]), .Z(n5575) );
  NOR U5246 ( .A(n5576), .B(n5575), .Z(n3246) );
  NOR U5247 ( .A(n3247), .B(n3246), .Z(n5578) );
  XOR U5248 ( .A(n3248), .B(b[749]), .Z(n5577) );
  NOR U5249 ( .A(n5578), .B(n5577), .Z(n3249) );
  NOR U5250 ( .A(n3250), .B(n3249), .Z(n5582) );
  XOR U5251 ( .A(n3251), .B(b[750]), .Z(n5581) );
  NOR U5252 ( .A(n5582), .B(n5581), .Z(n3252) );
  NOR U5253 ( .A(n3253), .B(n3252), .Z(n5584) );
  XOR U5254 ( .A(n3254), .B(b[751]), .Z(n5583) );
  NOR U5255 ( .A(n5584), .B(n5583), .Z(n3255) );
  NOR U5256 ( .A(n3256), .B(n3255), .Z(n5586) );
  XOR U5257 ( .A(n3257), .B(b[752]), .Z(n5585) );
  NOR U5258 ( .A(n5586), .B(n5585), .Z(n3258) );
  NOR U5259 ( .A(n3259), .B(n3258), .Z(n5588) );
  XOR U5260 ( .A(n3260), .B(b[753]), .Z(n5587) );
  NOR U5261 ( .A(n5588), .B(n5587), .Z(n3261) );
  NOR U5262 ( .A(n3262), .B(n3261), .Z(n5590) );
  XOR U5263 ( .A(n3263), .B(b[754]), .Z(n5589) );
  NOR U5264 ( .A(n5590), .B(n5589), .Z(n3264) );
  NOR U5265 ( .A(n3265), .B(n3264), .Z(n5592) );
  XOR U5266 ( .A(n3266), .B(b[755]), .Z(n5591) );
  NOR U5267 ( .A(n5592), .B(n5591), .Z(n3267) );
  NOR U5268 ( .A(n3268), .B(n3267), .Z(n5594) );
  XOR U5269 ( .A(n3269), .B(b[756]), .Z(n5593) );
  NOR U5270 ( .A(n5594), .B(n5593), .Z(n3270) );
  NOR U5271 ( .A(n3271), .B(n3270), .Z(n5596) );
  XOR U5272 ( .A(n3272), .B(b[757]), .Z(n5595) );
  NOR U5273 ( .A(n5596), .B(n5595), .Z(n3273) );
  NOR U5274 ( .A(n3274), .B(n3273), .Z(n5598) );
  XOR U5275 ( .A(n3275), .B(b[758]), .Z(n5597) );
  NOR U5276 ( .A(n5598), .B(n5597), .Z(n3276) );
  NOR U5277 ( .A(n3277), .B(n3276), .Z(n5600) );
  XOR U5278 ( .A(n3278), .B(b[759]), .Z(n5599) );
  NOR U5279 ( .A(n5600), .B(n5599), .Z(n3279) );
  NOR U5280 ( .A(n3280), .B(n3279), .Z(n5604) );
  XOR U5281 ( .A(n3281), .B(b[760]), .Z(n5603) );
  NOR U5282 ( .A(n5604), .B(n5603), .Z(n3282) );
  NOR U5283 ( .A(n3283), .B(n3282), .Z(n5606) );
  XOR U5284 ( .A(n3284), .B(b[761]), .Z(n5605) );
  NOR U5285 ( .A(n5606), .B(n5605), .Z(n3285) );
  NOR U5286 ( .A(n3286), .B(n3285), .Z(n5608) );
  XOR U5287 ( .A(n3287), .B(b[762]), .Z(n5607) );
  NOR U5288 ( .A(n5608), .B(n5607), .Z(n3288) );
  NOR U5289 ( .A(n3289), .B(n3288), .Z(n5610) );
  XOR U5290 ( .A(n3290), .B(b[763]), .Z(n5609) );
  NOR U5291 ( .A(n5610), .B(n5609), .Z(n3291) );
  NOR U5292 ( .A(n3292), .B(n3291), .Z(n5612) );
  XOR U5293 ( .A(n3293), .B(b[764]), .Z(n5611) );
  NOR U5294 ( .A(n5612), .B(n5611), .Z(n3294) );
  NOR U5295 ( .A(n3295), .B(n3294), .Z(n5614) );
  XOR U5296 ( .A(n3296), .B(b[765]), .Z(n5613) );
  NOR U5297 ( .A(n5614), .B(n5613), .Z(n3297) );
  NOR U5298 ( .A(n3298), .B(n3297), .Z(n5616) );
  XOR U5299 ( .A(n3299), .B(b[766]), .Z(n5615) );
  NOR U5300 ( .A(n5616), .B(n5615), .Z(n3300) );
  NOR U5301 ( .A(n3301), .B(n3300), .Z(n5618) );
  XOR U5302 ( .A(n3302), .B(b[767]), .Z(n5617) );
  NOR U5303 ( .A(n5618), .B(n5617), .Z(n3303) );
  NOR U5304 ( .A(n3304), .B(n3303), .Z(n5620) );
  XOR U5305 ( .A(n3305), .B(b[768]), .Z(n5619) );
  NOR U5306 ( .A(n5620), .B(n5619), .Z(n3306) );
  NOR U5307 ( .A(n3307), .B(n3306), .Z(n5622) );
  XOR U5308 ( .A(n3308), .B(b[769]), .Z(n5621) );
  NOR U5309 ( .A(n5622), .B(n5621), .Z(n3309) );
  NOR U5310 ( .A(n3310), .B(n3309), .Z(n5626) );
  XOR U5311 ( .A(n3311), .B(b[770]), .Z(n5625) );
  NOR U5312 ( .A(n5626), .B(n5625), .Z(n3312) );
  NOR U5313 ( .A(n3313), .B(n3312), .Z(n5628) );
  XOR U5314 ( .A(n3314), .B(b[771]), .Z(n5627) );
  NOR U5315 ( .A(n5628), .B(n5627), .Z(n3315) );
  NOR U5316 ( .A(n3316), .B(n3315), .Z(n5630) );
  XOR U5317 ( .A(n3317), .B(b[772]), .Z(n5629) );
  NOR U5318 ( .A(n5630), .B(n5629), .Z(n3318) );
  NOR U5319 ( .A(n3319), .B(n3318), .Z(n5632) );
  XOR U5320 ( .A(n3320), .B(b[773]), .Z(n5631) );
  NOR U5321 ( .A(n5632), .B(n5631), .Z(n3321) );
  NOR U5322 ( .A(n3322), .B(n3321), .Z(n5634) );
  XOR U5323 ( .A(n3323), .B(b[774]), .Z(n5633) );
  NOR U5324 ( .A(n5634), .B(n5633), .Z(n3324) );
  NOR U5325 ( .A(n3325), .B(n3324), .Z(n5636) );
  XOR U5326 ( .A(n3326), .B(b[775]), .Z(n5635) );
  NOR U5327 ( .A(n5636), .B(n5635), .Z(n3327) );
  NOR U5328 ( .A(n3328), .B(n3327), .Z(n5638) );
  XOR U5329 ( .A(n3329), .B(b[776]), .Z(n5637) );
  NOR U5330 ( .A(n5638), .B(n5637), .Z(n3330) );
  NOR U5331 ( .A(n3331), .B(n3330), .Z(n5640) );
  XOR U5332 ( .A(n3332), .B(b[777]), .Z(n5639) );
  NOR U5333 ( .A(n5640), .B(n5639), .Z(n3333) );
  NOR U5334 ( .A(n3334), .B(n3333), .Z(n5642) );
  XOR U5335 ( .A(n3335), .B(b[778]), .Z(n5641) );
  NOR U5336 ( .A(n5642), .B(n5641), .Z(n3336) );
  NOR U5337 ( .A(n3337), .B(n3336), .Z(n5644) );
  XOR U5338 ( .A(n3338), .B(b[779]), .Z(n5643) );
  NOR U5339 ( .A(n5644), .B(n5643), .Z(n3339) );
  NOR U5340 ( .A(n3340), .B(n3339), .Z(n5648) );
  XOR U5341 ( .A(n3341), .B(b[780]), .Z(n5647) );
  NOR U5342 ( .A(n5648), .B(n5647), .Z(n3342) );
  NOR U5343 ( .A(n3343), .B(n3342), .Z(n5650) );
  XOR U5344 ( .A(n3344), .B(b[781]), .Z(n5649) );
  NOR U5345 ( .A(n5650), .B(n5649), .Z(n3345) );
  NOR U5346 ( .A(n3346), .B(n3345), .Z(n5652) );
  XOR U5347 ( .A(n3347), .B(b[782]), .Z(n5651) );
  NOR U5348 ( .A(n5652), .B(n5651), .Z(n3348) );
  NOR U5349 ( .A(n3349), .B(n3348), .Z(n5654) );
  XOR U5350 ( .A(n3350), .B(b[783]), .Z(n5653) );
  NOR U5351 ( .A(n5654), .B(n5653), .Z(n3351) );
  NOR U5352 ( .A(n3352), .B(n3351), .Z(n5656) );
  XOR U5353 ( .A(n3353), .B(b[784]), .Z(n5655) );
  NOR U5354 ( .A(n5656), .B(n5655), .Z(n3354) );
  NOR U5355 ( .A(n3355), .B(n3354), .Z(n5658) );
  XOR U5356 ( .A(n3356), .B(b[785]), .Z(n5657) );
  NOR U5357 ( .A(n5658), .B(n5657), .Z(n3357) );
  NOR U5358 ( .A(n3358), .B(n3357), .Z(n5660) );
  XOR U5359 ( .A(n3359), .B(b[786]), .Z(n5659) );
  NOR U5360 ( .A(n5660), .B(n5659), .Z(n3360) );
  NOR U5361 ( .A(n3361), .B(n3360), .Z(n5662) );
  XOR U5362 ( .A(n3362), .B(b[787]), .Z(n5661) );
  NOR U5363 ( .A(n5662), .B(n5661), .Z(n3363) );
  NOR U5364 ( .A(n3364), .B(n3363), .Z(n5664) );
  XOR U5365 ( .A(n3365), .B(b[788]), .Z(n5663) );
  NOR U5366 ( .A(n5664), .B(n5663), .Z(n3366) );
  NOR U5367 ( .A(n3367), .B(n3366), .Z(n5666) );
  XOR U5368 ( .A(n3368), .B(b[789]), .Z(n5665) );
  NOR U5369 ( .A(n5666), .B(n5665), .Z(n3369) );
  NOR U5370 ( .A(n3370), .B(n3369), .Z(n5670) );
  XOR U5371 ( .A(n3371), .B(b[790]), .Z(n5669) );
  NOR U5372 ( .A(n5670), .B(n5669), .Z(n3372) );
  NOR U5373 ( .A(n3373), .B(n3372), .Z(n5672) );
  XOR U5374 ( .A(n3374), .B(b[791]), .Z(n5671) );
  NOR U5375 ( .A(n5672), .B(n5671), .Z(n3375) );
  NOR U5376 ( .A(n3376), .B(n3375), .Z(n5674) );
  XOR U5377 ( .A(n3377), .B(b[792]), .Z(n5673) );
  NOR U5378 ( .A(n5674), .B(n5673), .Z(n3378) );
  NOR U5379 ( .A(n3379), .B(n3378), .Z(n5676) );
  XOR U5380 ( .A(n3380), .B(b[793]), .Z(n5675) );
  NOR U5381 ( .A(n5676), .B(n5675), .Z(n3381) );
  NOR U5382 ( .A(n3382), .B(n3381), .Z(n5678) );
  XOR U5383 ( .A(n3383), .B(b[794]), .Z(n5677) );
  NOR U5384 ( .A(n5678), .B(n5677), .Z(n3384) );
  NOR U5385 ( .A(n3385), .B(n3384), .Z(n5680) );
  XOR U5386 ( .A(n3386), .B(b[795]), .Z(n5679) );
  NOR U5387 ( .A(n5680), .B(n5679), .Z(n3387) );
  NOR U5388 ( .A(n3388), .B(n3387), .Z(n5682) );
  XOR U5389 ( .A(n3389), .B(b[796]), .Z(n5681) );
  NOR U5390 ( .A(n5682), .B(n5681), .Z(n3390) );
  NOR U5391 ( .A(n3391), .B(n3390), .Z(n5684) );
  XOR U5392 ( .A(n3392), .B(b[797]), .Z(n5683) );
  NOR U5393 ( .A(n5684), .B(n5683), .Z(n3393) );
  NOR U5394 ( .A(n3394), .B(n3393), .Z(n5686) );
  XOR U5395 ( .A(n3395), .B(b[798]), .Z(n5685) );
  NOR U5396 ( .A(n5686), .B(n5685), .Z(n3396) );
  NOR U5397 ( .A(n3397), .B(n3396), .Z(n5688) );
  XOR U5398 ( .A(n3398), .B(b[799]), .Z(n5687) );
  NOR U5399 ( .A(n5688), .B(n5687), .Z(n3399) );
  NOR U5400 ( .A(n3400), .B(n3399), .Z(n5694) );
  XOR U5401 ( .A(n3401), .B(b[800]), .Z(n5693) );
  NOR U5402 ( .A(n5694), .B(n5693), .Z(n3402) );
  NOR U5403 ( .A(n3403), .B(n3402), .Z(n5696) );
  XOR U5404 ( .A(n3404), .B(b[801]), .Z(n5695) );
  NOR U5405 ( .A(n5696), .B(n5695), .Z(n3405) );
  NOR U5406 ( .A(n3406), .B(n3405), .Z(n5698) );
  XOR U5407 ( .A(n3407), .B(b[802]), .Z(n5697) );
  NOR U5408 ( .A(n5698), .B(n5697), .Z(n3408) );
  NOR U5409 ( .A(n3409), .B(n3408), .Z(n5700) );
  XOR U5410 ( .A(n3410), .B(b[803]), .Z(n5699) );
  NOR U5411 ( .A(n5700), .B(n5699), .Z(n3411) );
  NOR U5412 ( .A(n3412), .B(n3411), .Z(n5702) );
  XOR U5413 ( .A(n3413), .B(b[804]), .Z(n5701) );
  NOR U5414 ( .A(n5702), .B(n5701), .Z(n3414) );
  NOR U5415 ( .A(n3415), .B(n3414), .Z(n5704) );
  XOR U5416 ( .A(n3416), .B(b[805]), .Z(n5703) );
  NOR U5417 ( .A(n5704), .B(n5703), .Z(n3417) );
  NOR U5418 ( .A(n3418), .B(n3417), .Z(n5706) );
  XOR U5419 ( .A(n3419), .B(b[806]), .Z(n5705) );
  NOR U5420 ( .A(n5706), .B(n5705), .Z(n3420) );
  NOR U5421 ( .A(n3421), .B(n3420), .Z(n5708) );
  XOR U5422 ( .A(n3422), .B(b[807]), .Z(n5707) );
  NOR U5423 ( .A(n5708), .B(n5707), .Z(n3423) );
  NOR U5424 ( .A(n3424), .B(n3423), .Z(n5710) );
  XOR U5425 ( .A(n3425), .B(b[808]), .Z(n5709) );
  NOR U5426 ( .A(n5710), .B(n5709), .Z(n3426) );
  NOR U5427 ( .A(n3427), .B(n3426), .Z(n5712) );
  XOR U5428 ( .A(n3428), .B(b[809]), .Z(n5711) );
  NOR U5429 ( .A(n5712), .B(n5711), .Z(n3429) );
  NOR U5430 ( .A(n3430), .B(n3429), .Z(n5716) );
  XOR U5431 ( .A(n3431), .B(b[810]), .Z(n5715) );
  NOR U5432 ( .A(n5716), .B(n5715), .Z(n3432) );
  NOR U5433 ( .A(n3433), .B(n3432), .Z(n5718) );
  XOR U5434 ( .A(n3434), .B(b[811]), .Z(n5717) );
  NOR U5435 ( .A(n5718), .B(n5717), .Z(n3435) );
  NOR U5436 ( .A(n3436), .B(n3435), .Z(n5720) );
  XOR U5437 ( .A(n3437), .B(b[812]), .Z(n5719) );
  NOR U5438 ( .A(n5720), .B(n5719), .Z(n3438) );
  NOR U5439 ( .A(n3439), .B(n3438), .Z(n5722) );
  XOR U5440 ( .A(n3440), .B(b[813]), .Z(n5721) );
  NOR U5441 ( .A(n5722), .B(n5721), .Z(n3441) );
  NOR U5442 ( .A(n3442), .B(n3441), .Z(n5724) );
  XOR U5443 ( .A(n3443), .B(b[814]), .Z(n5723) );
  NOR U5444 ( .A(n5724), .B(n5723), .Z(n3444) );
  NOR U5445 ( .A(n3445), .B(n3444), .Z(n5726) );
  XOR U5446 ( .A(n3446), .B(b[815]), .Z(n5725) );
  NOR U5447 ( .A(n5726), .B(n5725), .Z(n3447) );
  NOR U5448 ( .A(n3448), .B(n3447), .Z(n5728) );
  XOR U5449 ( .A(n3449), .B(b[816]), .Z(n5727) );
  NOR U5450 ( .A(n5728), .B(n5727), .Z(n3450) );
  NOR U5451 ( .A(n3451), .B(n3450), .Z(n5730) );
  XOR U5452 ( .A(n3452), .B(b[817]), .Z(n5729) );
  NOR U5453 ( .A(n5730), .B(n5729), .Z(n3453) );
  NOR U5454 ( .A(n3454), .B(n3453), .Z(n5732) );
  XOR U5455 ( .A(n3455), .B(b[818]), .Z(n5731) );
  NOR U5456 ( .A(n5732), .B(n5731), .Z(n3456) );
  NOR U5457 ( .A(n3457), .B(n3456), .Z(n5734) );
  XOR U5458 ( .A(n3458), .B(b[819]), .Z(n5733) );
  NOR U5459 ( .A(n5734), .B(n5733), .Z(n3459) );
  NOR U5460 ( .A(n3460), .B(n3459), .Z(n5738) );
  XOR U5461 ( .A(n3461), .B(b[820]), .Z(n5737) );
  NOR U5462 ( .A(n5738), .B(n5737), .Z(n3462) );
  NOR U5463 ( .A(n3463), .B(n3462), .Z(n5740) );
  XOR U5464 ( .A(n3464), .B(b[821]), .Z(n5739) );
  NOR U5465 ( .A(n5740), .B(n5739), .Z(n3465) );
  NOR U5466 ( .A(n3466), .B(n3465), .Z(n5742) );
  XOR U5467 ( .A(n3467), .B(b[822]), .Z(n5741) );
  NOR U5468 ( .A(n5742), .B(n5741), .Z(n3468) );
  NOR U5469 ( .A(n3469), .B(n3468), .Z(n5744) );
  XOR U5470 ( .A(n3470), .B(b[823]), .Z(n5743) );
  NOR U5471 ( .A(n5744), .B(n5743), .Z(n3471) );
  NOR U5472 ( .A(n3472), .B(n3471), .Z(n5746) );
  XOR U5473 ( .A(n3473), .B(b[824]), .Z(n5745) );
  NOR U5474 ( .A(n5746), .B(n5745), .Z(n3474) );
  NOR U5475 ( .A(n3475), .B(n3474), .Z(n5748) );
  XOR U5476 ( .A(n3476), .B(b[825]), .Z(n5747) );
  NOR U5477 ( .A(n5748), .B(n5747), .Z(n3477) );
  NOR U5478 ( .A(n3478), .B(n3477), .Z(n5750) );
  XOR U5479 ( .A(n3479), .B(b[826]), .Z(n5749) );
  NOR U5480 ( .A(n5750), .B(n5749), .Z(n3480) );
  NOR U5481 ( .A(n3481), .B(n3480), .Z(n5752) );
  XOR U5482 ( .A(n3482), .B(b[827]), .Z(n5751) );
  NOR U5483 ( .A(n5752), .B(n5751), .Z(n3483) );
  NOR U5484 ( .A(n3484), .B(n3483), .Z(n5754) );
  XOR U5485 ( .A(n3485), .B(b[828]), .Z(n5753) );
  NOR U5486 ( .A(n5754), .B(n5753), .Z(n3486) );
  NOR U5487 ( .A(n3487), .B(n3486), .Z(n5756) );
  XOR U5488 ( .A(n3488), .B(b[829]), .Z(n5755) );
  NOR U5489 ( .A(n5756), .B(n5755), .Z(n3489) );
  NOR U5490 ( .A(n3490), .B(n3489), .Z(n5760) );
  XOR U5491 ( .A(n3491), .B(b[830]), .Z(n5759) );
  NOR U5492 ( .A(n5760), .B(n5759), .Z(n3492) );
  NOR U5493 ( .A(n3493), .B(n3492), .Z(n5762) );
  XOR U5494 ( .A(n3494), .B(b[831]), .Z(n5761) );
  NOR U5495 ( .A(n5762), .B(n5761), .Z(n3495) );
  NOR U5496 ( .A(n3496), .B(n3495), .Z(n5764) );
  XOR U5497 ( .A(n3497), .B(b[832]), .Z(n5763) );
  NOR U5498 ( .A(n5764), .B(n5763), .Z(n3498) );
  NOR U5499 ( .A(n3499), .B(n3498), .Z(n5766) );
  XOR U5500 ( .A(n3500), .B(b[833]), .Z(n5765) );
  NOR U5501 ( .A(n5766), .B(n5765), .Z(n3501) );
  NOR U5502 ( .A(n3502), .B(n3501), .Z(n5768) );
  XOR U5503 ( .A(n3503), .B(b[834]), .Z(n5767) );
  NOR U5504 ( .A(n5768), .B(n5767), .Z(n3504) );
  NOR U5505 ( .A(n3505), .B(n3504), .Z(n5770) );
  XOR U5506 ( .A(n3506), .B(b[835]), .Z(n5769) );
  NOR U5507 ( .A(n5770), .B(n5769), .Z(n3507) );
  NOR U5508 ( .A(n3508), .B(n3507), .Z(n5772) );
  XOR U5509 ( .A(n3509), .B(b[836]), .Z(n5771) );
  NOR U5510 ( .A(n5772), .B(n5771), .Z(n3510) );
  NOR U5511 ( .A(n3511), .B(n3510), .Z(n5774) );
  XOR U5512 ( .A(n3512), .B(b[837]), .Z(n5773) );
  NOR U5513 ( .A(n5774), .B(n5773), .Z(n3513) );
  NOR U5514 ( .A(n3514), .B(n3513), .Z(n5776) );
  XOR U5515 ( .A(n3515), .B(b[838]), .Z(n5775) );
  NOR U5516 ( .A(n5776), .B(n5775), .Z(n3516) );
  NOR U5517 ( .A(n3517), .B(n3516), .Z(n5778) );
  XOR U5518 ( .A(n3518), .B(b[839]), .Z(n5777) );
  NOR U5519 ( .A(n5778), .B(n5777), .Z(n3519) );
  NOR U5520 ( .A(n3520), .B(n3519), .Z(n5782) );
  XOR U5521 ( .A(n3521), .B(b[840]), .Z(n5781) );
  NOR U5522 ( .A(n5782), .B(n5781), .Z(n3522) );
  NOR U5523 ( .A(n3523), .B(n3522), .Z(n5784) );
  XOR U5524 ( .A(n3524), .B(b[841]), .Z(n5783) );
  NOR U5525 ( .A(n5784), .B(n5783), .Z(n3525) );
  NOR U5526 ( .A(n3526), .B(n3525), .Z(n5786) );
  XOR U5527 ( .A(n3527), .B(b[842]), .Z(n5785) );
  NOR U5528 ( .A(n5786), .B(n5785), .Z(n3528) );
  NOR U5529 ( .A(n3529), .B(n3528), .Z(n5788) );
  XOR U5530 ( .A(n3530), .B(b[843]), .Z(n5787) );
  NOR U5531 ( .A(n5788), .B(n5787), .Z(n3531) );
  NOR U5532 ( .A(n3532), .B(n3531), .Z(n5790) );
  XOR U5533 ( .A(n3533), .B(b[844]), .Z(n5789) );
  NOR U5534 ( .A(n5790), .B(n5789), .Z(n3534) );
  NOR U5535 ( .A(n3535), .B(n3534), .Z(n5792) );
  XOR U5536 ( .A(n3536), .B(b[845]), .Z(n5791) );
  NOR U5537 ( .A(n5792), .B(n5791), .Z(n3537) );
  NOR U5538 ( .A(n3538), .B(n3537), .Z(n5794) );
  XOR U5539 ( .A(n3539), .B(b[846]), .Z(n5793) );
  NOR U5540 ( .A(n5794), .B(n5793), .Z(n3540) );
  NOR U5541 ( .A(n3541), .B(n3540), .Z(n5796) );
  XOR U5542 ( .A(n3542), .B(b[847]), .Z(n5795) );
  NOR U5543 ( .A(n5796), .B(n5795), .Z(n3543) );
  NOR U5544 ( .A(n3544), .B(n3543), .Z(n5798) );
  XOR U5545 ( .A(n3545), .B(b[848]), .Z(n5797) );
  NOR U5546 ( .A(n5798), .B(n5797), .Z(n3546) );
  NOR U5547 ( .A(n3547), .B(n3546), .Z(n5800) );
  XOR U5548 ( .A(n3548), .B(b[849]), .Z(n5799) );
  NOR U5549 ( .A(n5800), .B(n5799), .Z(n3549) );
  NOR U5550 ( .A(n3550), .B(n3549), .Z(n5804) );
  XOR U5551 ( .A(n3551), .B(b[850]), .Z(n5803) );
  NOR U5552 ( .A(n5804), .B(n5803), .Z(n3552) );
  NOR U5553 ( .A(n3553), .B(n3552), .Z(n5806) );
  XOR U5554 ( .A(n3554), .B(b[851]), .Z(n5805) );
  NOR U5555 ( .A(n5806), .B(n5805), .Z(n3555) );
  NOR U5556 ( .A(n3556), .B(n3555), .Z(n5808) );
  XOR U5557 ( .A(n3557), .B(b[852]), .Z(n5807) );
  NOR U5558 ( .A(n5808), .B(n5807), .Z(n3558) );
  NOR U5559 ( .A(n3559), .B(n3558), .Z(n5810) );
  XOR U5560 ( .A(n3560), .B(b[853]), .Z(n5809) );
  NOR U5561 ( .A(n5810), .B(n5809), .Z(n3561) );
  NOR U5562 ( .A(n3562), .B(n3561), .Z(n5812) );
  XOR U5563 ( .A(n3563), .B(b[854]), .Z(n5811) );
  NOR U5564 ( .A(n5812), .B(n5811), .Z(n3564) );
  NOR U5565 ( .A(n3565), .B(n3564), .Z(n5814) );
  XOR U5566 ( .A(n3566), .B(b[855]), .Z(n5813) );
  NOR U5567 ( .A(n5814), .B(n5813), .Z(n3567) );
  NOR U5568 ( .A(n3568), .B(n3567), .Z(n5816) );
  XOR U5569 ( .A(n3569), .B(b[856]), .Z(n5815) );
  NOR U5570 ( .A(n5816), .B(n5815), .Z(n3570) );
  NOR U5571 ( .A(n3571), .B(n3570), .Z(n5818) );
  XOR U5572 ( .A(n3572), .B(b[857]), .Z(n5817) );
  NOR U5573 ( .A(n5818), .B(n5817), .Z(n3573) );
  NOR U5574 ( .A(n3574), .B(n3573), .Z(n5820) );
  XOR U5575 ( .A(n3575), .B(b[858]), .Z(n5819) );
  NOR U5576 ( .A(n5820), .B(n5819), .Z(n3576) );
  NOR U5577 ( .A(n3577), .B(n3576), .Z(n5822) );
  XOR U5578 ( .A(n3578), .B(b[859]), .Z(n5821) );
  NOR U5579 ( .A(n5822), .B(n5821), .Z(n3579) );
  NOR U5580 ( .A(n3580), .B(n3579), .Z(n5826) );
  XOR U5581 ( .A(n3581), .B(b[860]), .Z(n5825) );
  NOR U5582 ( .A(n5826), .B(n5825), .Z(n3582) );
  NOR U5583 ( .A(n3583), .B(n3582), .Z(n5828) );
  XOR U5584 ( .A(n3584), .B(b[861]), .Z(n5827) );
  NOR U5585 ( .A(n5828), .B(n5827), .Z(n3585) );
  NOR U5586 ( .A(n3586), .B(n3585), .Z(n5830) );
  XOR U5587 ( .A(n3587), .B(b[862]), .Z(n5829) );
  NOR U5588 ( .A(n5830), .B(n5829), .Z(n3588) );
  NOR U5589 ( .A(n3589), .B(n3588), .Z(n5832) );
  XOR U5590 ( .A(n3590), .B(b[863]), .Z(n5831) );
  NOR U5591 ( .A(n5832), .B(n5831), .Z(n3591) );
  NOR U5592 ( .A(n3592), .B(n3591), .Z(n5834) );
  XOR U5593 ( .A(n3593), .B(b[864]), .Z(n5833) );
  NOR U5594 ( .A(n5834), .B(n5833), .Z(n3594) );
  NOR U5595 ( .A(n3595), .B(n3594), .Z(n5836) );
  XOR U5596 ( .A(n3596), .B(b[865]), .Z(n5835) );
  NOR U5597 ( .A(n5836), .B(n5835), .Z(n3597) );
  NOR U5598 ( .A(n3598), .B(n3597), .Z(n5838) );
  XOR U5599 ( .A(n3599), .B(b[866]), .Z(n5837) );
  NOR U5600 ( .A(n5838), .B(n5837), .Z(n3600) );
  NOR U5601 ( .A(n3601), .B(n3600), .Z(n5840) );
  XOR U5602 ( .A(n3602), .B(b[867]), .Z(n5839) );
  NOR U5603 ( .A(n5840), .B(n5839), .Z(n3603) );
  NOR U5604 ( .A(n3604), .B(n3603), .Z(n5842) );
  XOR U5605 ( .A(n3605), .B(b[868]), .Z(n5841) );
  NOR U5606 ( .A(n5842), .B(n5841), .Z(n3606) );
  NOR U5607 ( .A(n3607), .B(n3606), .Z(n5844) );
  XOR U5608 ( .A(n3608), .B(b[869]), .Z(n5843) );
  NOR U5609 ( .A(n5844), .B(n5843), .Z(n3609) );
  NOR U5610 ( .A(n3610), .B(n3609), .Z(n5848) );
  XOR U5611 ( .A(n3611), .B(b[870]), .Z(n5847) );
  NOR U5612 ( .A(n5848), .B(n5847), .Z(n3612) );
  NOR U5613 ( .A(n3613), .B(n3612), .Z(n5850) );
  XOR U5614 ( .A(n3614), .B(b[871]), .Z(n5849) );
  NOR U5615 ( .A(n5850), .B(n5849), .Z(n3615) );
  NOR U5616 ( .A(n3616), .B(n3615), .Z(n5852) );
  XOR U5617 ( .A(n3617), .B(b[872]), .Z(n5851) );
  NOR U5618 ( .A(n5852), .B(n5851), .Z(n3618) );
  NOR U5619 ( .A(n3619), .B(n3618), .Z(n5854) );
  XOR U5620 ( .A(n3620), .B(b[873]), .Z(n5853) );
  NOR U5621 ( .A(n5854), .B(n5853), .Z(n3621) );
  NOR U5622 ( .A(n3622), .B(n3621), .Z(n5856) );
  XOR U5623 ( .A(n3623), .B(b[874]), .Z(n5855) );
  NOR U5624 ( .A(n5856), .B(n5855), .Z(n3624) );
  NOR U5625 ( .A(n3625), .B(n3624), .Z(n5858) );
  XOR U5626 ( .A(n3626), .B(b[875]), .Z(n5857) );
  NOR U5627 ( .A(n5858), .B(n5857), .Z(n3627) );
  NOR U5628 ( .A(n3628), .B(n3627), .Z(n5860) );
  XOR U5629 ( .A(n3629), .B(b[876]), .Z(n5859) );
  NOR U5630 ( .A(n5860), .B(n5859), .Z(n3630) );
  NOR U5631 ( .A(n3631), .B(n3630), .Z(n5862) );
  XOR U5632 ( .A(n3632), .B(b[877]), .Z(n5861) );
  NOR U5633 ( .A(n5862), .B(n5861), .Z(n3633) );
  NOR U5634 ( .A(n3634), .B(n3633), .Z(n5864) );
  XOR U5635 ( .A(n3635), .B(b[878]), .Z(n5863) );
  NOR U5636 ( .A(n5864), .B(n5863), .Z(n3636) );
  NOR U5637 ( .A(n3637), .B(n3636), .Z(n5866) );
  XOR U5638 ( .A(n3638), .B(b[879]), .Z(n5865) );
  NOR U5639 ( .A(n5866), .B(n5865), .Z(n3639) );
  NOR U5640 ( .A(n3640), .B(n3639), .Z(n5870) );
  XOR U5641 ( .A(n3641), .B(b[880]), .Z(n5869) );
  NOR U5642 ( .A(n5870), .B(n5869), .Z(n3642) );
  NOR U5643 ( .A(n3643), .B(n3642), .Z(n5872) );
  XOR U5644 ( .A(n3644), .B(b[881]), .Z(n5871) );
  NOR U5645 ( .A(n5872), .B(n5871), .Z(n3645) );
  NOR U5646 ( .A(n3646), .B(n3645), .Z(n5874) );
  XOR U5647 ( .A(n3647), .B(b[882]), .Z(n5873) );
  NOR U5648 ( .A(n5874), .B(n5873), .Z(n3648) );
  NOR U5649 ( .A(n3649), .B(n3648), .Z(n5876) );
  XOR U5650 ( .A(n3650), .B(b[883]), .Z(n5875) );
  NOR U5651 ( .A(n5876), .B(n5875), .Z(n3651) );
  NOR U5652 ( .A(n3652), .B(n3651), .Z(n5878) );
  XOR U5653 ( .A(n3653), .B(b[884]), .Z(n5877) );
  NOR U5654 ( .A(n5878), .B(n5877), .Z(n3654) );
  NOR U5655 ( .A(n3655), .B(n3654), .Z(n5880) );
  XOR U5656 ( .A(n3656), .B(b[885]), .Z(n5879) );
  NOR U5657 ( .A(n5880), .B(n5879), .Z(n3657) );
  NOR U5658 ( .A(n3658), .B(n3657), .Z(n5882) );
  XOR U5659 ( .A(n3659), .B(b[886]), .Z(n5881) );
  NOR U5660 ( .A(n5882), .B(n5881), .Z(n3660) );
  NOR U5661 ( .A(n3661), .B(n3660), .Z(n5884) );
  XOR U5662 ( .A(n3662), .B(b[887]), .Z(n5883) );
  NOR U5663 ( .A(n5884), .B(n5883), .Z(n3663) );
  NOR U5664 ( .A(n3664), .B(n3663), .Z(n5886) );
  XOR U5665 ( .A(n3665), .B(b[888]), .Z(n5885) );
  NOR U5666 ( .A(n5886), .B(n5885), .Z(n3666) );
  NOR U5667 ( .A(n3667), .B(n3666), .Z(n5888) );
  XOR U5668 ( .A(n3668), .B(b[889]), .Z(n5887) );
  NOR U5669 ( .A(n5888), .B(n5887), .Z(n3669) );
  NOR U5670 ( .A(n3670), .B(n3669), .Z(n5892) );
  XOR U5671 ( .A(n3671), .B(b[890]), .Z(n5891) );
  NOR U5672 ( .A(n5892), .B(n5891), .Z(n3672) );
  NOR U5673 ( .A(n3673), .B(n3672), .Z(n5894) );
  XOR U5674 ( .A(n3674), .B(b[891]), .Z(n5893) );
  NOR U5675 ( .A(n5894), .B(n5893), .Z(n3675) );
  NOR U5676 ( .A(n3676), .B(n3675), .Z(n5896) );
  XOR U5677 ( .A(n3677), .B(b[892]), .Z(n5895) );
  NOR U5678 ( .A(n5896), .B(n5895), .Z(n3678) );
  NOR U5679 ( .A(n3679), .B(n3678), .Z(n5898) );
  XOR U5680 ( .A(n3680), .B(b[893]), .Z(n5897) );
  NOR U5681 ( .A(n5898), .B(n5897), .Z(n3681) );
  NOR U5682 ( .A(n3682), .B(n3681), .Z(n5900) );
  XOR U5683 ( .A(n3683), .B(b[894]), .Z(n5899) );
  NOR U5684 ( .A(n5900), .B(n5899), .Z(n3684) );
  NOR U5685 ( .A(n3685), .B(n3684), .Z(n5902) );
  XOR U5686 ( .A(n3686), .B(b[895]), .Z(n5901) );
  NOR U5687 ( .A(n5902), .B(n5901), .Z(n3687) );
  NOR U5688 ( .A(n3688), .B(n3687), .Z(n5904) );
  XOR U5689 ( .A(n3689), .B(b[896]), .Z(n5903) );
  NOR U5690 ( .A(n5904), .B(n5903), .Z(n3690) );
  NOR U5691 ( .A(n3691), .B(n3690), .Z(n5906) );
  XOR U5692 ( .A(n3692), .B(b[897]), .Z(n5905) );
  NOR U5693 ( .A(n5906), .B(n5905), .Z(n3693) );
  NOR U5694 ( .A(n3694), .B(n3693), .Z(n5908) );
  XOR U5695 ( .A(n3695), .B(b[898]), .Z(n5907) );
  NOR U5696 ( .A(n5908), .B(n5907), .Z(n3696) );
  NOR U5697 ( .A(n3697), .B(n3696), .Z(n5910) );
  XOR U5698 ( .A(n3698), .B(b[899]), .Z(n5909) );
  NOR U5699 ( .A(n5910), .B(n5909), .Z(n3699) );
  NOR U5700 ( .A(n3700), .B(n3699), .Z(n5916) );
  XOR U5701 ( .A(n3701), .B(b[900]), .Z(n5915) );
  NOR U5702 ( .A(n5916), .B(n5915), .Z(n3702) );
  NOR U5703 ( .A(n3703), .B(n3702), .Z(n5918) );
  XOR U5704 ( .A(n3704), .B(b[901]), .Z(n5917) );
  NOR U5705 ( .A(n5918), .B(n5917), .Z(n3705) );
  NOR U5706 ( .A(n3706), .B(n3705), .Z(n5920) );
  XOR U5707 ( .A(n3707), .B(b[902]), .Z(n5919) );
  NOR U5708 ( .A(n5920), .B(n5919), .Z(n3708) );
  NOR U5709 ( .A(n3709), .B(n3708), .Z(n5922) );
  XOR U5710 ( .A(n3710), .B(b[903]), .Z(n5921) );
  NOR U5711 ( .A(n5922), .B(n5921), .Z(n3711) );
  NOR U5712 ( .A(n3712), .B(n3711), .Z(n5924) );
  XOR U5713 ( .A(n3713), .B(b[904]), .Z(n5923) );
  NOR U5714 ( .A(n5924), .B(n5923), .Z(n3714) );
  NOR U5715 ( .A(n3715), .B(n3714), .Z(n5926) );
  XOR U5716 ( .A(n3716), .B(b[905]), .Z(n5925) );
  NOR U5717 ( .A(n5926), .B(n5925), .Z(n3717) );
  NOR U5718 ( .A(n3718), .B(n3717), .Z(n5928) );
  XOR U5719 ( .A(n3719), .B(b[906]), .Z(n5927) );
  NOR U5720 ( .A(n5928), .B(n5927), .Z(n3720) );
  NOR U5721 ( .A(n3721), .B(n3720), .Z(n5930) );
  XOR U5722 ( .A(n3722), .B(b[907]), .Z(n5929) );
  NOR U5723 ( .A(n5930), .B(n5929), .Z(n3723) );
  NOR U5724 ( .A(n3724), .B(n3723), .Z(n5932) );
  XOR U5725 ( .A(n3725), .B(b[908]), .Z(n5931) );
  NOR U5726 ( .A(n5932), .B(n5931), .Z(n3726) );
  NOR U5727 ( .A(n3727), .B(n3726), .Z(n5934) );
  XOR U5728 ( .A(n3728), .B(b[909]), .Z(n5933) );
  NOR U5729 ( .A(n5934), .B(n5933), .Z(n3729) );
  NOR U5730 ( .A(n3730), .B(n3729), .Z(n5938) );
  XOR U5731 ( .A(n3731), .B(b[910]), .Z(n5937) );
  NOR U5732 ( .A(n5938), .B(n5937), .Z(n3732) );
  NOR U5733 ( .A(n3733), .B(n3732), .Z(n5940) );
  XOR U5734 ( .A(n3734), .B(b[911]), .Z(n5939) );
  NOR U5735 ( .A(n5940), .B(n5939), .Z(n3735) );
  NOR U5736 ( .A(n3736), .B(n3735), .Z(n5942) );
  XOR U5737 ( .A(n3737), .B(b[912]), .Z(n5941) );
  NOR U5738 ( .A(n5942), .B(n5941), .Z(n3738) );
  NOR U5739 ( .A(n3739), .B(n3738), .Z(n5944) );
  XOR U5740 ( .A(n3740), .B(b[913]), .Z(n5943) );
  NOR U5741 ( .A(n5944), .B(n5943), .Z(n3741) );
  NOR U5742 ( .A(n3742), .B(n3741), .Z(n5946) );
  XOR U5743 ( .A(n3743), .B(b[914]), .Z(n5945) );
  NOR U5744 ( .A(n5946), .B(n5945), .Z(n3744) );
  NOR U5745 ( .A(n3745), .B(n3744), .Z(n5948) );
  XOR U5746 ( .A(n3746), .B(b[915]), .Z(n5947) );
  NOR U5747 ( .A(n5948), .B(n5947), .Z(n3747) );
  NOR U5748 ( .A(n3748), .B(n3747), .Z(n5950) );
  XOR U5749 ( .A(n3749), .B(b[916]), .Z(n5949) );
  NOR U5750 ( .A(n5950), .B(n5949), .Z(n3750) );
  NOR U5751 ( .A(n3751), .B(n3750), .Z(n5952) );
  XOR U5752 ( .A(n3752), .B(b[917]), .Z(n5951) );
  NOR U5753 ( .A(n5952), .B(n5951), .Z(n3753) );
  NOR U5754 ( .A(n3754), .B(n3753), .Z(n5954) );
  XOR U5755 ( .A(n3755), .B(b[918]), .Z(n5953) );
  NOR U5756 ( .A(n5954), .B(n5953), .Z(n3756) );
  NOR U5757 ( .A(n3757), .B(n3756), .Z(n5956) );
  XOR U5758 ( .A(n3758), .B(b[919]), .Z(n5955) );
  NOR U5759 ( .A(n5956), .B(n5955), .Z(n3759) );
  NOR U5760 ( .A(n3760), .B(n3759), .Z(n5960) );
  XOR U5761 ( .A(n3761), .B(b[920]), .Z(n5959) );
  NOR U5762 ( .A(n5960), .B(n5959), .Z(n3762) );
  NOR U5763 ( .A(n3763), .B(n3762), .Z(n5962) );
  XOR U5764 ( .A(n3764), .B(b[921]), .Z(n5961) );
  NOR U5765 ( .A(n5962), .B(n5961), .Z(n3765) );
  NOR U5766 ( .A(n3766), .B(n3765), .Z(n5964) );
  XOR U5767 ( .A(n3767), .B(b[922]), .Z(n5963) );
  NOR U5768 ( .A(n5964), .B(n5963), .Z(n3768) );
  NOR U5769 ( .A(n3769), .B(n3768), .Z(n5966) );
  XOR U5770 ( .A(n3770), .B(b[923]), .Z(n5965) );
  NOR U5771 ( .A(n5966), .B(n5965), .Z(n3771) );
  NOR U5772 ( .A(n3772), .B(n3771), .Z(n5968) );
  XOR U5773 ( .A(n3773), .B(b[924]), .Z(n5967) );
  NOR U5774 ( .A(n5968), .B(n5967), .Z(n3774) );
  NOR U5775 ( .A(n3775), .B(n3774), .Z(n5970) );
  XOR U5776 ( .A(n3776), .B(b[925]), .Z(n5969) );
  NOR U5777 ( .A(n5970), .B(n5969), .Z(n3777) );
  NOR U5778 ( .A(n3778), .B(n3777), .Z(n5972) );
  XOR U5779 ( .A(n3779), .B(b[926]), .Z(n5971) );
  NOR U5780 ( .A(n5972), .B(n5971), .Z(n3780) );
  NOR U5781 ( .A(n3781), .B(n3780), .Z(n5974) );
  XOR U5782 ( .A(n3782), .B(b[927]), .Z(n5973) );
  NOR U5783 ( .A(n5974), .B(n5973), .Z(n3783) );
  NOR U5784 ( .A(n3784), .B(n3783), .Z(n5976) );
  XOR U5785 ( .A(n3785), .B(b[928]), .Z(n5975) );
  NOR U5786 ( .A(n5976), .B(n5975), .Z(n3786) );
  NOR U5787 ( .A(n3787), .B(n3786), .Z(n5978) );
  XOR U5788 ( .A(n3788), .B(b[929]), .Z(n5977) );
  NOR U5789 ( .A(n5978), .B(n5977), .Z(n3789) );
  NOR U5790 ( .A(n3790), .B(n3789), .Z(n5982) );
  XOR U5791 ( .A(n3791), .B(b[930]), .Z(n5981) );
  NOR U5792 ( .A(n5982), .B(n5981), .Z(n3792) );
  NOR U5793 ( .A(n3793), .B(n3792), .Z(n5984) );
  XOR U5794 ( .A(n3794), .B(b[931]), .Z(n5983) );
  NOR U5795 ( .A(n5984), .B(n5983), .Z(n3795) );
  NOR U5796 ( .A(n3796), .B(n3795), .Z(n5986) );
  XOR U5797 ( .A(n3797), .B(b[932]), .Z(n5985) );
  NOR U5798 ( .A(n5986), .B(n5985), .Z(n3798) );
  NOR U5799 ( .A(n3799), .B(n3798), .Z(n5988) );
  XOR U5800 ( .A(n3800), .B(b[933]), .Z(n5987) );
  NOR U5801 ( .A(n5988), .B(n5987), .Z(n3801) );
  NOR U5802 ( .A(n3802), .B(n3801), .Z(n5990) );
  XOR U5803 ( .A(n3803), .B(b[934]), .Z(n5989) );
  NOR U5804 ( .A(n5990), .B(n5989), .Z(n3804) );
  NOR U5805 ( .A(n3805), .B(n3804), .Z(n5992) );
  XOR U5806 ( .A(n3806), .B(b[935]), .Z(n5991) );
  NOR U5807 ( .A(n5992), .B(n5991), .Z(n3807) );
  NOR U5808 ( .A(n3808), .B(n3807), .Z(n5994) );
  XOR U5809 ( .A(n3809), .B(b[936]), .Z(n5993) );
  NOR U5810 ( .A(n5994), .B(n5993), .Z(n3810) );
  NOR U5811 ( .A(n3811), .B(n3810), .Z(n5996) );
  XOR U5812 ( .A(n3812), .B(b[937]), .Z(n5995) );
  NOR U5813 ( .A(n5996), .B(n5995), .Z(n3813) );
  NOR U5814 ( .A(n3814), .B(n3813), .Z(n5998) );
  XOR U5815 ( .A(n3815), .B(b[938]), .Z(n5997) );
  NOR U5816 ( .A(n5998), .B(n5997), .Z(n3816) );
  NOR U5817 ( .A(n3817), .B(n3816), .Z(n6000) );
  XOR U5818 ( .A(n3818), .B(b[939]), .Z(n5999) );
  NOR U5819 ( .A(n6000), .B(n5999), .Z(n3819) );
  NOR U5820 ( .A(n3820), .B(n3819), .Z(n6004) );
  XOR U5821 ( .A(n3821), .B(b[940]), .Z(n6003) );
  NOR U5822 ( .A(n6004), .B(n6003), .Z(n3822) );
  NOR U5823 ( .A(n3823), .B(n3822), .Z(n6006) );
  XOR U5824 ( .A(n3824), .B(b[941]), .Z(n6005) );
  NOR U5825 ( .A(n6006), .B(n6005), .Z(n3825) );
  NOR U5826 ( .A(n3826), .B(n3825), .Z(n6008) );
  XOR U5827 ( .A(n3827), .B(b[942]), .Z(n6007) );
  NOR U5828 ( .A(n6008), .B(n6007), .Z(n3828) );
  NOR U5829 ( .A(n3829), .B(n3828), .Z(n6010) );
  XOR U5830 ( .A(n3830), .B(b[943]), .Z(n6009) );
  NOR U5831 ( .A(n6010), .B(n6009), .Z(n3831) );
  NOR U5832 ( .A(n3832), .B(n3831), .Z(n6012) );
  XOR U5833 ( .A(n3833), .B(b[944]), .Z(n6011) );
  NOR U5834 ( .A(n6012), .B(n6011), .Z(n3834) );
  NOR U5835 ( .A(n3835), .B(n3834), .Z(n6014) );
  XOR U5836 ( .A(n3836), .B(b[945]), .Z(n6013) );
  NOR U5837 ( .A(n6014), .B(n6013), .Z(n3837) );
  NOR U5838 ( .A(n3838), .B(n3837), .Z(n6016) );
  XOR U5839 ( .A(n3839), .B(b[946]), .Z(n6015) );
  NOR U5840 ( .A(n6016), .B(n6015), .Z(n3840) );
  NOR U5841 ( .A(n3841), .B(n3840), .Z(n6018) );
  XOR U5842 ( .A(n3842), .B(b[947]), .Z(n6017) );
  NOR U5843 ( .A(n6018), .B(n6017), .Z(n3843) );
  NOR U5844 ( .A(n3844), .B(n3843), .Z(n6020) );
  XOR U5845 ( .A(n3845), .B(b[948]), .Z(n6019) );
  NOR U5846 ( .A(n6020), .B(n6019), .Z(n3846) );
  NOR U5847 ( .A(n3847), .B(n3846), .Z(n6022) );
  XOR U5848 ( .A(n3848), .B(b[949]), .Z(n6021) );
  NOR U5849 ( .A(n6022), .B(n6021), .Z(n3849) );
  NOR U5850 ( .A(n3850), .B(n3849), .Z(n6026) );
  XOR U5851 ( .A(n3851), .B(b[950]), .Z(n6025) );
  NOR U5852 ( .A(n6026), .B(n6025), .Z(n3852) );
  NOR U5853 ( .A(n3853), .B(n3852), .Z(n6028) );
  XOR U5854 ( .A(n3854), .B(b[951]), .Z(n6027) );
  NOR U5855 ( .A(n6028), .B(n6027), .Z(n3855) );
  NOR U5856 ( .A(n3856), .B(n3855), .Z(n6030) );
  XOR U5857 ( .A(n3857), .B(b[952]), .Z(n6029) );
  NOR U5858 ( .A(n6030), .B(n6029), .Z(n3858) );
  NOR U5859 ( .A(n3859), .B(n3858), .Z(n6032) );
  XOR U5860 ( .A(n3860), .B(b[953]), .Z(n6031) );
  NOR U5861 ( .A(n6032), .B(n6031), .Z(n3861) );
  NOR U5862 ( .A(n3862), .B(n3861), .Z(n6034) );
  XOR U5863 ( .A(n3863), .B(b[954]), .Z(n6033) );
  NOR U5864 ( .A(n6034), .B(n6033), .Z(n3864) );
  NOR U5865 ( .A(n3865), .B(n3864), .Z(n6036) );
  XOR U5866 ( .A(n3866), .B(b[955]), .Z(n6035) );
  NOR U5867 ( .A(n6036), .B(n6035), .Z(n3867) );
  NOR U5868 ( .A(n3868), .B(n3867), .Z(n6038) );
  XOR U5869 ( .A(n3869), .B(b[956]), .Z(n6037) );
  NOR U5870 ( .A(n6038), .B(n6037), .Z(n3870) );
  NOR U5871 ( .A(n3871), .B(n3870), .Z(n6040) );
  XOR U5872 ( .A(n3872), .B(b[957]), .Z(n6039) );
  NOR U5873 ( .A(n6040), .B(n6039), .Z(n3873) );
  NOR U5874 ( .A(n3874), .B(n3873), .Z(n6042) );
  XOR U5875 ( .A(n3875), .B(b[958]), .Z(n6041) );
  NOR U5876 ( .A(n6042), .B(n6041), .Z(n3876) );
  NOR U5877 ( .A(n3877), .B(n3876), .Z(n6044) );
  XOR U5878 ( .A(n3878), .B(b[959]), .Z(n6043) );
  NOR U5879 ( .A(n6044), .B(n6043), .Z(n3879) );
  NOR U5880 ( .A(n3880), .B(n3879), .Z(n6048) );
  XOR U5881 ( .A(n3881), .B(b[960]), .Z(n6047) );
  NOR U5882 ( .A(n6048), .B(n6047), .Z(n3882) );
  NOR U5883 ( .A(n3883), .B(n3882), .Z(n6050) );
  XOR U5884 ( .A(n3884), .B(b[961]), .Z(n6049) );
  NOR U5885 ( .A(n6050), .B(n6049), .Z(n3885) );
  NOR U5886 ( .A(n3886), .B(n3885), .Z(n6052) );
  XOR U5887 ( .A(n3887), .B(b[962]), .Z(n6051) );
  NOR U5888 ( .A(n6052), .B(n6051), .Z(n3888) );
  NOR U5889 ( .A(n3889), .B(n3888), .Z(n6054) );
  XOR U5890 ( .A(n3890), .B(b[963]), .Z(n6053) );
  NOR U5891 ( .A(n6054), .B(n6053), .Z(n3891) );
  NOR U5892 ( .A(n3892), .B(n3891), .Z(n6056) );
  XOR U5893 ( .A(n3893), .B(b[964]), .Z(n6055) );
  NOR U5894 ( .A(n6056), .B(n6055), .Z(n3894) );
  NOR U5895 ( .A(n3895), .B(n3894), .Z(n6058) );
  XOR U5896 ( .A(n3896), .B(b[965]), .Z(n6057) );
  NOR U5897 ( .A(n6058), .B(n6057), .Z(n3897) );
  NOR U5898 ( .A(n3898), .B(n3897), .Z(n6060) );
  XOR U5899 ( .A(n3899), .B(b[966]), .Z(n6059) );
  NOR U5900 ( .A(n6060), .B(n6059), .Z(n3900) );
  NOR U5901 ( .A(n3901), .B(n3900), .Z(n6062) );
  XOR U5902 ( .A(n3902), .B(b[967]), .Z(n6061) );
  NOR U5903 ( .A(n6062), .B(n6061), .Z(n3903) );
  NOR U5904 ( .A(n3904), .B(n3903), .Z(n6064) );
  XOR U5905 ( .A(n3905), .B(b[968]), .Z(n6063) );
  NOR U5906 ( .A(n6064), .B(n6063), .Z(n3906) );
  NOR U5907 ( .A(n3907), .B(n3906), .Z(n6066) );
  XOR U5908 ( .A(n3908), .B(b[969]), .Z(n6065) );
  NOR U5909 ( .A(n6066), .B(n6065), .Z(n3909) );
  NOR U5910 ( .A(n3910), .B(n3909), .Z(n6070) );
  XOR U5911 ( .A(n3911), .B(b[970]), .Z(n6069) );
  NOR U5912 ( .A(n6070), .B(n6069), .Z(n3912) );
  NOR U5913 ( .A(n3913), .B(n3912), .Z(n6072) );
  XOR U5914 ( .A(n3914), .B(b[971]), .Z(n6071) );
  NOR U5915 ( .A(n6072), .B(n6071), .Z(n3915) );
  NOR U5916 ( .A(n3916), .B(n3915), .Z(n6074) );
  XOR U5917 ( .A(n3917), .B(b[972]), .Z(n6073) );
  NOR U5918 ( .A(n6074), .B(n6073), .Z(n3918) );
  NOR U5919 ( .A(n3919), .B(n3918), .Z(n6076) );
  XOR U5920 ( .A(n3920), .B(b[973]), .Z(n6075) );
  NOR U5921 ( .A(n6076), .B(n6075), .Z(n3921) );
  NOR U5922 ( .A(n3922), .B(n3921), .Z(n6078) );
  XOR U5923 ( .A(n3923), .B(b[974]), .Z(n6077) );
  NOR U5924 ( .A(n6078), .B(n6077), .Z(n3924) );
  NOR U5925 ( .A(n3925), .B(n3924), .Z(n6080) );
  XOR U5926 ( .A(n3926), .B(b[975]), .Z(n6079) );
  NOR U5927 ( .A(n6080), .B(n6079), .Z(n3927) );
  NOR U5928 ( .A(n3928), .B(n3927), .Z(n6082) );
  XOR U5929 ( .A(n3929), .B(b[976]), .Z(n6081) );
  NOR U5930 ( .A(n6082), .B(n6081), .Z(n3930) );
  NOR U5931 ( .A(n3931), .B(n3930), .Z(n6084) );
  XOR U5932 ( .A(n3932), .B(b[977]), .Z(n6083) );
  NOR U5933 ( .A(n6084), .B(n6083), .Z(n3933) );
  NOR U5934 ( .A(n3934), .B(n3933), .Z(n6086) );
  XOR U5935 ( .A(n3935), .B(b[978]), .Z(n6085) );
  NOR U5936 ( .A(n6086), .B(n6085), .Z(n3936) );
  NOR U5937 ( .A(n3937), .B(n3936), .Z(n6088) );
  XOR U5938 ( .A(n3938), .B(b[979]), .Z(n6087) );
  NOR U5939 ( .A(n6088), .B(n6087), .Z(n3939) );
  NOR U5940 ( .A(n3940), .B(n3939), .Z(n6092) );
  XOR U5941 ( .A(n3941), .B(b[980]), .Z(n6091) );
  NOR U5942 ( .A(n6092), .B(n6091), .Z(n3942) );
  NOR U5943 ( .A(n3943), .B(n3942), .Z(n6094) );
  XOR U5944 ( .A(n3944), .B(b[981]), .Z(n6093) );
  NOR U5945 ( .A(n6094), .B(n6093), .Z(n3945) );
  NOR U5946 ( .A(n3946), .B(n3945), .Z(n6096) );
  XOR U5947 ( .A(n3947), .B(b[982]), .Z(n6095) );
  NOR U5948 ( .A(n6096), .B(n6095), .Z(n3948) );
  NOR U5949 ( .A(n3949), .B(n3948), .Z(n6098) );
  XOR U5950 ( .A(n3950), .B(b[983]), .Z(n6097) );
  NOR U5951 ( .A(n6098), .B(n6097), .Z(n3951) );
  NOR U5952 ( .A(n3952), .B(n3951), .Z(n6100) );
  XOR U5953 ( .A(n3953), .B(b[984]), .Z(n6099) );
  NOR U5954 ( .A(n6100), .B(n6099), .Z(n3954) );
  NOR U5955 ( .A(n3955), .B(n3954), .Z(n6102) );
  XOR U5956 ( .A(n3956), .B(b[985]), .Z(n6101) );
  NOR U5957 ( .A(n6102), .B(n6101), .Z(n3957) );
  NOR U5958 ( .A(n3958), .B(n3957), .Z(n6104) );
  XOR U5959 ( .A(n3959), .B(b[986]), .Z(n6103) );
  NOR U5960 ( .A(n6104), .B(n6103), .Z(n3960) );
  NOR U5961 ( .A(n3961), .B(n3960), .Z(n6106) );
  XOR U5962 ( .A(n3962), .B(b[987]), .Z(n6105) );
  NOR U5963 ( .A(n6106), .B(n6105), .Z(n3963) );
  NOR U5964 ( .A(n3964), .B(n3963), .Z(n6108) );
  XOR U5965 ( .A(n3965), .B(b[988]), .Z(n6107) );
  NOR U5966 ( .A(n6108), .B(n6107), .Z(n3966) );
  NOR U5967 ( .A(n3967), .B(n3966), .Z(n6110) );
  XOR U5968 ( .A(n3968), .B(b[989]), .Z(n6109) );
  NOR U5969 ( .A(n6110), .B(n6109), .Z(n3969) );
  NOR U5970 ( .A(n3970), .B(n3969), .Z(n6114) );
  XOR U5971 ( .A(n3971), .B(b[990]), .Z(n6113) );
  NOR U5972 ( .A(n6114), .B(n6113), .Z(n3972) );
  NOR U5973 ( .A(n3973), .B(n3972), .Z(n6116) );
  XOR U5974 ( .A(n3974), .B(b[991]), .Z(n6115) );
  NOR U5975 ( .A(n6116), .B(n6115), .Z(n3975) );
  NOR U5976 ( .A(n3976), .B(n3975), .Z(n6118) );
  XOR U5977 ( .A(n3977), .B(b[992]), .Z(n6117) );
  NOR U5978 ( .A(n6118), .B(n6117), .Z(n3978) );
  NOR U5979 ( .A(n3979), .B(n3978), .Z(n6120) );
  XOR U5980 ( .A(n3980), .B(b[993]), .Z(n6119) );
  NOR U5981 ( .A(n6120), .B(n6119), .Z(n3981) );
  NOR U5982 ( .A(n3982), .B(n3981), .Z(n6122) );
  XOR U5983 ( .A(n3983), .B(b[994]), .Z(n6121) );
  NOR U5984 ( .A(n6122), .B(n6121), .Z(n3984) );
  NOR U5985 ( .A(n3985), .B(n3984), .Z(n6124) );
  XOR U5986 ( .A(n3986), .B(b[995]), .Z(n6123) );
  NOR U5987 ( .A(n6124), .B(n6123), .Z(n3987) );
  NOR U5988 ( .A(n3988), .B(n3987), .Z(n6126) );
  XOR U5989 ( .A(n3989), .B(b[996]), .Z(n6125) );
  NOR U5990 ( .A(n6126), .B(n6125), .Z(n3990) );
  NOR U5991 ( .A(n3991), .B(n3990), .Z(n6128) );
  XOR U5992 ( .A(n3992), .B(b[997]), .Z(n6127) );
  NOR U5993 ( .A(n6128), .B(n6127), .Z(n3993) );
  NOR U5994 ( .A(n3994), .B(n3993), .Z(n6130) );
  XOR U5995 ( .A(n3995), .B(b[998]), .Z(n6129) );
  NOR U5996 ( .A(n6130), .B(n6129), .Z(n3996) );
  NOR U5997 ( .A(n3997), .B(n3996), .Z(n6132) );
  XOR U5998 ( .A(n3998), .B(a[999]), .Z(n6131) );
  NOR U5999 ( .A(n6132), .B(n6131), .Z(n3999) );
  NOR U6000 ( .A(n4000), .B(n3999), .Z(n4004) );
  IV U6001 ( .A(a[1000]), .Z(n4002) );
  XOR U6002 ( .A(n4002), .B(b[1000]), .Z(n4003) );
  XOR U6003 ( .A(n4004), .B(n4003), .Z(c[1000]) );
  IV U6004 ( .A(b[1000]), .Z(n4001) );
  NOR U6005 ( .A(n4002), .B(n4001), .Z(n4006) );
  NOR U6006 ( .A(n4004), .B(n4003), .Z(n4005) );
  NOR U6007 ( .A(n4006), .B(n4005), .Z(n4010) );
  IV U6008 ( .A(a[1001]), .Z(n4008) );
  XOR U6009 ( .A(n4008), .B(b[1001]), .Z(n4009) );
  XOR U6010 ( .A(n4010), .B(n4009), .Z(c[1001]) );
  IV U6011 ( .A(b[1001]), .Z(n4007) );
  NOR U6012 ( .A(n4008), .B(n4007), .Z(n4012) );
  NOR U6013 ( .A(n4010), .B(n4009), .Z(n4011) );
  NOR U6014 ( .A(n4012), .B(n4011), .Z(n4016) );
  IV U6015 ( .A(a[1002]), .Z(n4014) );
  XOR U6016 ( .A(n4014), .B(b[1002]), .Z(n4015) );
  XOR U6017 ( .A(n4016), .B(n4015), .Z(c[1002]) );
  IV U6018 ( .A(b[1002]), .Z(n4013) );
  NOR U6019 ( .A(n4014), .B(n4013), .Z(n4018) );
  NOR U6020 ( .A(n4016), .B(n4015), .Z(n4017) );
  NOR U6021 ( .A(n4018), .B(n4017), .Z(n4022) );
  IV U6022 ( .A(a[1003]), .Z(n4020) );
  XOR U6023 ( .A(n4020), .B(b[1003]), .Z(n4021) );
  XOR U6024 ( .A(n4022), .B(n4021), .Z(c[1003]) );
  IV U6025 ( .A(b[1003]), .Z(n4019) );
  NOR U6026 ( .A(n4020), .B(n4019), .Z(n4024) );
  NOR U6027 ( .A(n4022), .B(n4021), .Z(n4023) );
  NOR U6028 ( .A(n4024), .B(n4023), .Z(n4028) );
  IV U6029 ( .A(a[1004]), .Z(n4026) );
  XOR U6030 ( .A(n4026), .B(b[1004]), .Z(n4027) );
  XOR U6031 ( .A(n4028), .B(n4027), .Z(c[1004]) );
  IV U6032 ( .A(b[1004]), .Z(n4025) );
  NOR U6033 ( .A(n4026), .B(n4025), .Z(n4030) );
  NOR U6034 ( .A(n4028), .B(n4027), .Z(n4029) );
  NOR U6035 ( .A(n4030), .B(n4029), .Z(n4034) );
  IV U6036 ( .A(a[1005]), .Z(n4032) );
  XOR U6037 ( .A(n4032), .B(b[1005]), .Z(n4033) );
  XOR U6038 ( .A(n4034), .B(n4033), .Z(c[1005]) );
  IV U6039 ( .A(b[1005]), .Z(n4031) );
  NOR U6040 ( .A(n4032), .B(n4031), .Z(n4036) );
  NOR U6041 ( .A(n4034), .B(n4033), .Z(n4035) );
  NOR U6042 ( .A(n4036), .B(n4035), .Z(n4040) );
  IV U6043 ( .A(a[1006]), .Z(n4038) );
  XOR U6044 ( .A(n4038), .B(b[1006]), .Z(n4039) );
  XOR U6045 ( .A(n4040), .B(n4039), .Z(c[1006]) );
  IV U6046 ( .A(b[1006]), .Z(n4037) );
  NOR U6047 ( .A(n4038), .B(n4037), .Z(n4042) );
  NOR U6048 ( .A(n4040), .B(n4039), .Z(n4041) );
  NOR U6049 ( .A(n4042), .B(n4041), .Z(n4046) );
  IV U6050 ( .A(a[1007]), .Z(n4044) );
  XOR U6051 ( .A(n4044), .B(b[1007]), .Z(n4045) );
  XOR U6052 ( .A(n4046), .B(n4045), .Z(c[1007]) );
  IV U6053 ( .A(b[1007]), .Z(n4043) );
  NOR U6054 ( .A(n4044), .B(n4043), .Z(n4048) );
  NOR U6055 ( .A(n4046), .B(n4045), .Z(n4047) );
  NOR U6056 ( .A(n4048), .B(n4047), .Z(n4052) );
  IV U6057 ( .A(a[1008]), .Z(n4050) );
  XOR U6058 ( .A(n4050), .B(b[1008]), .Z(n4051) );
  XOR U6059 ( .A(n4052), .B(n4051), .Z(c[1008]) );
  IV U6060 ( .A(b[1008]), .Z(n4049) );
  NOR U6061 ( .A(n4050), .B(n4049), .Z(n4054) );
  NOR U6062 ( .A(n4052), .B(n4051), .Z(n4053) );
  NOR U6063 ( .A(n4054), .B(n4053), .Z(n4060) );
  IV U6064 ( .A(a[1009]), .Z(n4058) );
  XOR U6065 ( .A(n4058), .B(b[1009]), .Z(n4059) );
  XOR U6066 ( .A(n4060), .B(n4059), .Z(c[1009]) );
  XOR U6067 ( .A(n4056), .B(n4055), .Z(c[100]) );
  IV U6068 ( .A(b[1009]), .Z(n4057) );
  NOR U6069 ( .A(n4058), .B(n4057), .Z(n4062) );
  NOR U6070 ( .A(n4060), .B(n4059), .Z(n4061) );
  NOR U6071 ( .A(n4062), .B(n4061), .Z(n4066) );
  IV U6072 ( .A(a[1010]), .Z(n4064) );
  XOR U6073 ( .A(n4064), .B(b[1010]), .Z(n4065) );
  XOR U6074 ( .A(n4066), .B(n4065), .Z(c[1010]) );
  IV U6075 ( .A(b[1010]), .Z(n4063) );
  NOR U6076 ( .A(n4064), .B(n4063), .Z(n4068) );
  NOR U6077 ( .A(n4066), .B(n4065), .Z(n4067) );
  NOR U6078 ( .A(n4068), .B(n4067), .Z(n4072) );
  IV U6079 ( .A(a[1011]), .Z(n4070) );
  XOR U6080 ( .A(n4070), .B(b[1011]), .Z(n4071) );
  XOR U6081 ( .A(n4072), .B(n4071), .Z(c[1011]) );
  IV U6082 ( .A(b[1011]), .Z(n4069) );
  NOR U6083 ( .A(n4070), .B(n4069), .Z(n4074) );
  NOR U6084 ( .A(n4072), .B(n4071), .Z(n4073) );
  NOR U6085 ( .A(n4074), .B(n4073), .Z(n4078) );
  IV U6086 ( .A(a[1012]), .Z(n4076) );
  XOR U6087 ( .A(n4076), .B(b[1012]), .Z(n4077) );
  XOR U6088 ( .A(n4078), .B(n4077), .Z(c[1012]) );
  IV U6089 ( .A(b[1012]), .Z(n4075) );
  NOR U6090 ( .A(n4076), .B(n4075), .Z(n4080) );
  NOR U6091 ( .A(n4078), .B(n4077), .Z(n4079) );
  NOR U6092 ( .A(n4080), .B(n4079), .Z(n4084) );
  IV U6093 ( .A(a[1013]), .Z(n4082) );
  XOR U6094 ( .A(n4082), .B(b[1013]), .Z(n4083) );
  XOR U6095 ( .A(n4084), .B(n4083), .Z(c[1013]) );
  IV U6096 ( .A(b[1013]), .Z(n4081) );
  NOR U6097 ( .A(n4082), .B(n4081), .Z(n4086) );
  NOR U6098 ( .A(n4084), .B(n4083), .Z(n4085) );
  NOR U6099 ( .A(n4086), .B(n4085), .Z(n4090) );
  IV U6100 ( .A(a[1014]), .Z(n4088) );
  XOR U6101 ( .A(n4088), .B(b[1014]), .Z(n4089) );
  XOR U6102 ( .A(n4090), .B(n4089), .Z(c[1014]) );
  IV U6103 ( .A(b[1014]), .Z(n4087) );
  NOR U6104 ( .A(n4088), .B(n4087), .Z(n4092) );
  NOR U6105 ( .A(n4090), .B(n4089), .Z(n4091) );
  NOR U6106 ( .A(n4092), .B(n4091), .Z(n4096) );
  IV U6107 ( .A(a[1015]), .Z(n4094) );
  XOR U6108 ( .A(n4094), .B(b[1015]), .Z(n4095) );
  XOR U6109 ( .A(n4096), .B(n4095), .Z(c[1015]) );
  IV U6110 ( .A(b[1015]), .Z(n4093) );
  NOR U6111 ( .A(n4094), .B(n4093), .Z(n4098) );
  NOR U6112 ( .A(n4096), .B(n4095), .Z(n4097) );
  NOR U6113 ( .A(n4098), .B(n4097), .Z(n4102) );
  IV U6114 ( .A(a[1016]), .Z(n4100) );
  XOR U6115 ( .A(n4100), .B(b[1016]), .Z(n4101) );
  XOR U6116 ( .A(n4102), .B(n4101), .Z(c[1016]) );
  IV U6117 ( .A(b[1016]), .Z(n4099) );
  NOR U6118 ( .A(n4100), .B(n4099), .Z(n4104) );
  NOR U6119 ( .A(n4102), .B(n4101), .Z(n4103) );
  NOR U6120 ( .A(n4104), .B(n4103), .Z(n4108) );
  IV U6121 ( .A(a[1017]), .Z(n4106) );
  XOR U6122 ( .A(n4106), .B(b[1017]), .Z(n4107) );
  XOR U6123 ( .A(n4108), .B(n4107), .Z(c[1017]) );
  IV U6124 ( .A(b[1017]), .Z(n4105) );
  NOR U6125 ( .A(n4106), .B(n4105), .Z(n4110) );
  NOR U6126 ( .A(n4108), .B(n4107), .Z(n4109) );
  NOR U6127 ( .A(n4110), .B(n4109), .Z(n4114) );
  IV U6128 ( .A(a[1018]), .Z(n4112) );
  XOR U6129 ( .A(n4112), .B(b[1018]), .Z(n4113) );
  XOR U6130 ( .A(n4114), .B(n4113), .Z(c[1018]) );
  IV U6131 ( .A(b[1018]), .Z(n4111) );
  NOR U6132 ( .A(n4112), .B(n4111), .Z(n4116) );
  NOR U6133 ( .A(n4114), .B(n4113), .Z(n4115) );
  NOR U6134 ( .A(n4116), .B(n4115), .Z(n4122) );
  IV U6135 ( .A(a[1019]), .Z(n4120) );
  XOR U6136 ( .A(n4120), .B(b[1019]), .Z(n4121) );
  XOR U6137 ( .A(n4122), .B(n4121), .Z(c[1019]) );
  XOR U6138 ( .A(n4118), .B(n4117), .Z(c[101]) );
  IV U6139 ( .A(b[1019]), .Z(n4119) );
  NOR U6140 ( .A(n4120), .B(n4119), .Z(n4124) );
  NOR U6141 ( .A(n4122), .B(n4121), .Z(n4123) );
  NOR U6142 ( .A(n4124), .B(n4123), .Z(n4128) );
  IV U6143 ( .A(a[1020]), .Z(n4126) );
  XOR U6144 ( .A(n4126), .B(b[1020]), .Z(n4127) );
  XOR U6145 ( .A(n4128), .B(n4127), .Z(c[1020]) );
  IV U6146 ( .A(b[1020]), .Z(n4125) );
  NOR U6147 ( .A(n4126), .B(n4125), .Z(n4130) );
  NOR U6148 ( .A(n4128), .B(n4127), .Z(n4129) );
  NOR U6149 ( .A(n4130), .B(n4129), .Z(n4134) );
  IV U6150 ( .A(a[1021]), .Z(n4132) );
  XOR U6151 ( .A(n4132), .B(b[1021]), .Z(n4133) );
  XOR U6152 ( .A(n4134), .B(n4133), .Z(c[1021]) );
  IV U6153 ( .A(b[1021]), .Z(n4131) );
  NOR U6154 ( .A(n4132), .B(n4131), .Z(n4136) );
  NOR U6155 ( .A(n4134), .B(n4133), .Z(n4135) );
  NOR U6156 ( .A(n4136), .B(n4135), .Z(n4140) );
  IV U6157 ( .A(a[1022]), .Z(n4138) );
  XOR U6158 ( .A(n4138), .B(b[1022]), .Z(n4139) );
  XOR U6159 ( .A(n4140), .B(n4139), .Z(c[1022]) );
  IV U6160 ( .A(b[1022]), .Z(n4137) );
  NOR U6161 ( .A(n4138), .B(n4137), .Z(n4142) );
  NOR U6162 ( .A(n4140), .B(n4139), .Z(n4141) );
  NOR U6163 ( .A(n4142), .B(n4141), .Z(n6140) );
  XOR U6164 ( .A(n6140), .B(a[1023]), .Z(n6138) );
  IV U6165 ( .A(b[1023]), .Z(n6137) );
  XOR U6166 ( .A(n6138), .B(n6137), .Z(c[1023]) );
  XOR U6167 ( .A(n4144), .B(n4143), .Z(c[102]) );
  XOR U6168 ( .A(n4146), .B(n4145), .Z(c[103]) );
  XOR U6169 ( .A(n4148), .B(n4147), .Z(c[104]) );
  XOR U6170 ( .A(n4150), .B(n4149), .Z(c[105]) );
  XOR U6171 ( .A(n4152), .B(n4151), .Z(c[106]) );
  XOR U6172 ( .A(n4154), .B(n4153), .Z(c[107]) );
  XOR U6173 ( .A(n4156), .B(n4155), .Z(c[108]) );
  XOR U6174 ( .A(n4158), .B(n4157), .Z(c[109]) );
  XOR U6175 ( .A(n4160), .B(n4159), .Z(c[10]) );
  XOR U6176 ( .A(n4162), .B(n4161), .Z(c[110]) );
  XOR U6177 ( .A(n4164), .B(n4163), .Z(c[111]) );
  XOR U6178 ( .A(n4166), .B(n4165), .Z(c[112]) );
  XOR U6179 ( .A(n4168), .B(n4167), .Z(c[113]) );
  XOR U6180 ( .A(n4170), .B(n4169), .Z(c[114]) );
  XOR U6181 ( .A(n4172), .B(n4171), .Z(c[115]) );
  XOR U6182 ( .A(n4174), .B(n4173), .Z(c[116]) );
  XOR U6183 ( .A(n4176), .B(n4175), .Z(c[117]) );
  XOR U6184 ( .A(n4178), .B(n4177), .Z(c[118]) );
  XOR U6185 ( .A(n4180), .B(n4179), .Z(c[119]) );
  XOR U6186 ( .A(n4182), .B(n4181), .Z(c[11]) );
  XOR U6187 ( .A(n4184), .B(n4183), .Z(c[120]) );
  XOR U6188 ( .A(n4186), .B(n4185), .Z(c[121]) );
  XOR U6189 ( .A(n4188), .B(n4187), .Z(c[122]) );
  XOR U6190 ( .A(n4190), .B(n4189), .Z(c[123]) );
  XOR U6191 ( .A(n4192), .B(n4191), .Z(c[124]) );
  XOR U6192 ( .A(n4194), .B(n4193), .Z(c[125]) );
  XOR U6193 ( .A(n4196), .B(n4195), .Z(c[126]) );
  XOR U6194 ( .A(n4198), .B(n4197), .Z(c[127]) );
  XOR U6195 ( .A(n4200), .B(n4199), .Z(c[128]) );
  XOR U6196 ( .A(n4202), .B(n4201), .Z(c[129]) );
  XOR U6197 ( .A(n4204), .B(n4203), .Z(c[12]) );
  XOR U6198 ( .A(n4206), .B(n4205), .Z(c[130]) );
  XOR U6199 ( .A(n4208), .B(n4207), .Z(c[131]) );
  XOR U6200 ( .A(n4210), .B(n4209), .Z(c[132]) );
  XOR U6201 ( .A(n4212), .B(n4211), .Z(c[133]) );
  XOR U6202 ( .A(n4214), .B(n4213), .Z(c[134]) );
  XOR U6203 ( .A(n4216), .B(n4215), .Z(c[135]) );
  XOR U6204 ( .A(n4218), .B(n4217), .Z(c[136]) );
  XOR U6205 ( .A(n4220), .B(n4219), .Z(c[137]) );
  XOR U6206 ( .A(n4222), .B(n4221), .Z(c[138]) );
  XOR U6207 ( .A(n4224), .B(n4223), .Z(c[139]) );
  XOR U6208 ( .A(n4226), .B(n4225), .Z(c[13]) );
  XOR U6209 ( .A(n4228), .B(n4227), .Z(c[140]) );
  XOR U6210 ( .A(n4230), .B(n4229), .Z(c[141]) );
  XOR U6211 ( .A(n4232), .B(n4231), .Z(c[142]) );
  XOR U6212 ( .A(n4234), .B(n4233), .Z(c[143]) );
  XOR U6213 ( .A(n4236), .B(n4235), .Z(c[144]) );
  XOR U6214 ( .A(n4238), .B(n4237), .Z(c[145]) );
  XOR U6215 ( .A(n4240), .B(n4239), .Z(c[146]) );
  XOR U6216 ( .A(n4242), .B(n4241), .Z(c[147]) );
  XOR U6217 ( .A(n4244), .B(n4243), .Z(c[148]) );
  XOR U6218 ( .A(n4246), .B(n4245), .Z(c[149]) );
  XOR U6219 ( .A(n4248), .B(n4247), .Z(c[14]) );
  XOR U6220 ( .A(n4250), .B(n4249), .Z(c[150]) );
  XOR U6221 ( .A(n4252), .B(n4251), .Z(c[151]) );
  XOR U6222 ( .A(n4254), .B(n4253), .Z(c[152]) );
  XOR U6223 ( .A(n4256), .B(n4255), .Z(c[153]) );
  XOR U6224 ( .A(n4258), .B(n4257), .Z(c[154]) );
  XOR U6225 ( .A(n4260), .B(n4259), .Z(c[155]) );
  XOR U6226 ( .A(n4262), .B(n4261), .Z(c[156]) );
  XOR U6227 ( .A(n4264), .B(n4263), .Z(c[157]) );
  XOR U6228 ( .A(n4266), .B(n4265), .Z(c[158]) );
  XOR U6229 ( .A(n4268), .B(n4267), .Z(c[159]) );
  XOR U6230 ( .A(n4270), .B(n4269), .Z(c[15]) );
  XOR U6231 ( .A(n4272), .B(n4271), .Z(c[160]) );
  XOR U6232 ( .A(n4274), .B(n4273), .Z(c[161]) );
  XOR U6233 ( .A(n4276), .B(n4275), .Z(c[162]) );
  XOR U6234 ( .A(n4278), .B(n4277), .Z(c[163]) );
  XOR U6235 ( .A(n4280), .B(n4279), .Z(c[164]) );
  XOR U6236 ( .A(n4282), .B(n4281), .Z(c[165]) );
  XOR U6237 ( .A(n4284), .B(n4283), .Z(c[166]) );
  XOR U6238 ( .A(n4286), .B(n4285), .Z(c[167]) );
  XOR U6239 ( .A(n4288), .B(n4287), .Z(c[168]) );
  XOR U6240 ( .A(n4290), .B(n4289), .Z(c[169]) );
  XOR U6241 ( .A(n4292), .B(n4291), .Z(c[16]) );
  XOR U6242 ( .A(n4294), .B(n4293), .Z(c[170]) );
  XOR U6243 ( .A(n4296), .B(n4295), .Z(c[171]) );
  XOR U6244 ( .A(n4298), .B(n4297), .Z(c[172]) );
  XOR U6245 ( .A(n4300), .B(n4299), .Z(c[173]) );
  XOR U6246 ( .A(n4302), .B(n4301), .Z(c[174]) );
  XOR U6247 ( .A(n4304), .B(n4303), .Z(c[175]) );
  XOR U6248 ( .A(n4306), .B(n4305), .Z(c[176]) );
  XOR U6249 ( .A(n4308), .B(n4307), .Z(c[177]) );
  XOR U6250 ( .A(n4310), .B(n4309), .Z(c[178]) );
  XOR U6251 ( .A(n4312), .B(n4311), .Z(c[179]) );
  XOR U6252 ( .A(n4314), .B(n4313), .Z(c[17]) );
  XOR U6253 ( .A(n4316), .B(n4315), .Z(c[180]) );
  XOR U6254 ( .A(n4318), .B(n4317), .Z(c[181]) );
  XOR U6255 ( .A(n4320), .B(n4319), .Z(c[182]) );
  XOR U6256 ( .A(n4322), .B(n4321), .Z(c[183]) );
  XOR U6257 ( .A(n4324), .B(n4323), .Z(c[184]) );
  XOR U6258 ( .A(n4326), .B(n4325), .Z(c[185]) );
  XOR U6259 ( .A(n4328), .B(n4327), .Z(c[186]) );
  XOR U6260 ( .A(n4330), .B(n4329), .Z(c[187]) );
  XOR U6261 ( .A(n4332), .B(n4331), .Z(c[188]) );
  XOR U6262 ( .A(n4334), .B(n4333), .Z(c[189]) );
  XOR U6263 ( .A(n4336), .B(n4335), .Z(c[18]) );
  XOR U6264 ( .A(n4338), .B(n4337), .Z(c[190]) );
  XOR U6265 ( .A(n4340), .B(n4339), .Z(c[191]) );
  XOR U6266 ( .A(n4342), .B(n4341), .Z(c[192]) );
  XOR U6267 ( .A(n4344), .B(n4343), .Z(c[193]) );
  XOR U6268 ( .A(n4346), .B(n4345), .Z(c[194]) );
  XOR U6269 ( .A(n4348), .B(n4347), .Z(c[195]) );
  XOR U6270 ( .A(n4350), .B(n4349), .Z(c[196]) );
  XOR U6271 ( .A(n4352), .B(n4351), .Z(c[197]) );
  XOR U6272 ( .A(n4354), .B(n4353), .Z(c[198]) );
  XOR U6273 ( .A(n4356), .B(n4355), .Z(c[199]) );
  XOR U6274 ( .A(n4358), .B(n4357), .Z(c[19]) );
  XOR U6275 ( .A(n4360), .B(n4359), .Z(c[1]) );
  XOR U6276 ( .A(n4362), .B(n4361), .Z(c[200]) );
  XOR U6277 ( .A(n4364), .B(n4363), .Z(c[201]) );
  XOR U6278 ( .A(n4366), .B(n4365), .Z(c[202]) );
  XOR U6279 ( .A(n4368), .B(n4367), .Z(c[203]) );
  XOR U6280 ( .A(n4370), .B(n4369), .Z(c[204]) );
  XOR U6281 ( .A(n4372), .B(n4371), .Z(c[205]) );
  XOR U6282 ( .A(n4374), .B(n4373), .Z(c[206]) );
  XOR U6283 ( .A(n4376), .B(n4375), .Z(c[207]) );
  XOR U6284 ( .A(n4378), .B(n4377), .Z(c[208]) );
  XOR U6285 ( .A(n4380), .B(n4379), .Z(c[209]) );
  XOR U6286 ( .A(n4382), .B(n4381), .Z(c[20]) );
  XOR U6287 ( .A(n4384), .B(n4383), .Z(c[210]) );
  XOR U6288 ( .A(n4386), .B(n4385), .Z(c[211]) );
  XOR U6289 ( .A(n4388), .B(n4387), .Z(c[212]) );
  XOR U6290 ( .A(n4390), .B(n4389), .Z(c[213]) );
  XOR U6291 ( .A(n4392), .B(n4391), .Z(c[214]) );
  XOR U6292 ( .A(n4394), .B(n4393), .Z(c[215]) );
  XOR U6293 ( .A(n4396), .B(n4395), .Z(c[216]) );
  XOR U6294 ( .A(n4398), .B(n4397), .Z(c[217]) );
  XOR U6295 ( .A(n4400), .B(n4399), .Z(c[218]) );
  XOR U6296 ( .A(n4402), .B(n4401), .Z(c[219]) );
  XOR U6297 ( .A(n4404), .B(n4403), .Z(c[21]) );
  XOR U6298 ( .A(n4406), .B(n4405), .Z(c[220]) );
  XOR U6299 ( .A(n4408), .B(n4407), .Z(c[221]) );
  XOR U6300 ( .A(n4410), .B(n4409), .Z(c[222]) );
  XOR U6301 ( .A(n4412), .B(n4411), .Z(c[223]) );
  XOR U6302 ( .A(n4414), .B(n4413), .Z(c[224]) );
  XOR U6303 ( .A(n4416), .B(n4415), .Z(c[225]) );
  XOR U6304 ( .A(n4418), .B(n4417), .Z(c[226]) );
  XOR U6305 ( .A(n4420), .B(n4419), .Z(c[227]) );
  XOR U6306 ( .A(n4422), .B(n4421), .Z(c[228]) );
  XOR U6307 ( .A(n4424), .B(n4423), .Z(c[229]) );
  XOR U6308 ( .A(n4426), .B(n4425), .Z(c[22]) );
  XOR U6309 ( .A(n4428), .B(n4427), .Z(c[230]) );
  XOR U6310 ( .A(n4430), .B(n4429), .Z(c[231]) );
  XOR U6311 ( .A(n4432), .B(n4431), .Z(c[232]) );
  XOR U6312 ( .A(n4434), .B(n4433), .Z(c[233]) );
  XOR U6313 ( .A(n4436), .B(n4435), .Z(c[234]) );
  XOR U6314 ( .A(n4438), .B(n4437), .Z(c[235]) );
  XOR U6315 ( .A(n4440), .B(n4439), .Z(c[236]) );
  XOR U6316 ( .A(n4442), .B(n4441), .Z(c[237]) );
  XOR U6317 ( .A(n4444), .B(n4443), .Z(c[238]) );
  XOR U6318 ( .A(n4446), .B(n4445), .Z(c[239]) );
  XOR U6319 ( .A(n4448), .B(n4447), .Z(c[23]) );
  XOR U6320 ( .A(n4450), .B(n4449), .Z(c[240]) );
  XOR U6321 ( .A(n4452), .B(n4451), .Z(c[241]) );
  XOR U6322 ( .A(n4454), .B(n4453), .Z(c[242]) );
  XOR U6323 ( .A(n4456), .B(n4455), .Z(c[243]) );
  XOR U6324 ( .A(n4458), .B(n4457), .Z(c[244]) );
  XOR U6325 ( .A(n4460), .B(n4459), .Z(c[245]) );
  XOR U6326 ( .A(n4462), .B(n4461), .Z(c[246]) );
  XOR U6327 ( .A(n4464), .B(n4463), .Z(c[247]) );
  XOR U6328 ( .A(n4466), .B(n4465), .Z(c[248]) );
  XOR U6329 ( .A(n4468), .B(n4467), .Z(c[249]) );
  XOR U6330 ( .A(n4470), .B(n4469), .Z(c[24]) );
  XOR U6331 ( .A(n4472), .B(n4471), .Z(c[250]) );
  XOR U6332 ( .A(n4474), .B(n4473), .Z(c[251]) );
  XOR U6333 ( .A(n4476), .B(n4475), .Z(c[252]) );
  XOR U6334 ( .A(n4478), .B(n4477), .Z(c[253]) );
  XOR U6335 ( .A(n4480), .B(n4479), .Z(c[254]) );
  XOR U6336 ( .A(n4482), .B(n4481), .Z(c[255]) );
  XOR U6337 ( .A(n4484), .B(n4483), .Z(c[256]) );
  XOR U6338 ( .A(n4486), .B(n4485), .Z(c[257]) );
  XOR U6339 ( .A(n4488), .B(n4487), .Z(c[258]) );
  XOR U6340 ( .A(n4490), .B(n4489), .Z(c[259]) );
  XOR U6341 ( .A(n4492), .B(n4491), .Z(c[25]) );
  XOR U6342 ( .A(n4494), .B(n4493), .Z(c[260]) );
  XOR U6343 ( .A(n4496), .B(n4495), .Z(c[261]) );
  XOR U6344 ( .A(n4498), .B(n4497), .Z(c[262]) );
  XOR U6345 ( .A(n4500), .B(n4499), .Z(c[263]) );
  XOR U6346 ( .A(n4502), .B(n4501), .Z(c[264]) );
  XOR U6347 ( .A(n4504), .B(n4503), .Z(c[265]) );
  XOR U6348 ( .A(n4506), .B(n4505), .Z(c[266]) );
  XOR U6349 ( .A(n4508), .B(n4507), .Z(c[267]) );
  XOR U6350 ( .A(n4510), .B(n4509), .Z(c[268]) );
  XOR U6351 ( .A(n4512), .B(n4511), .Z(c[269]) );
  XOR U6352 ( .A(n4514), .B(n4513), .Z(c[26]) );
  XOR U6353 ( .A(n4516), .B(n4515), .Z(c[270]) );
  XOR U6354 ( .A(n4518), .B(n4517), .Z(c[271]) );
  XOR U6355 ( .A(n4520), .B(n4519), .Z(c[272]) );
  XOR U6356 ( .A(n4522), .B(n4521), .Z(c[273]) );
  XOR U6357 ( .A(n4524), .B(n4523), .Z(c[274]) );
  XOR U6358 ( .A(n4526), .B(n4525), .Z(c[275]) );
  XOR U6359 ( .A(n4528), .B(n4527), .Z(c[276]) );
  XOR U6360 ( .A(n4530), .B(n4529), .Z(c[277]) );
  XOR U6361 ( .A(n4532), .B(n4531), .Z(c[278]) );
  XOR U6362 ( .A(n4534), .B(n4533), .Z(c[279]) );
  XOR U6363 ( .A(n4536), .B(n4535), .Z(c[27]) );
  XOR U6364 ( .A(n4538), .B(n4537), .Z(c[280]) );
  XOR U6365 ( .A(n4540), .B(n4539), .Z(c[281]) );
  XOR U6366 ( .A(n4542), .B(n4541), .Z(c[282]) );
  XOR U6367 ( .A(n4544), .B(n4543), .Z(c[283]) );
  XOR U6368 ( .A(n4546), .B(n4545), .Z(c[284]) );
  XOR U6369 ( .A(n4548), .B(n4547), .Z(c[285]) );
  XOR U6370 ( .A(n4550), .B(n4549), .Z(c[286]) );
  XOR U6371 ( .A(n4552), .B(n4551), .Z(c[287]) );
  XOR U6372 ( .A(n4554), .B(n4553), .Z(c[288]) );
  XOR U6373 ( .A(n4556), .B(n4555), .Z(c[289]) );
  XOR U6374 ( .A(n4558), .B(n4557), .Z(c[28]) );
  XOR U6375 ( .A(n4560), .B(n4559), .Z(c[290]) );
  XOR U6376 ( .A(n4562), .B(n4561), .Z(c[291]) );
  XOR U6377 ( .A(n4564), .B(n4563), .Z(c[292]) );
  XOR U6378 ( .A(n4566), .B(n4565), .Z(c[293]) );
  XOR U6379 ( .A(n4568), .B(n4567), .Z(c[294]) );
  XOR U6380 ( .A(n4570), .B(n4569), .Z(c[295]) );
  XOR U6381 ( .A(n4572), .B(n4571), .Z(c[296]) );
  XOR U6382 ( .A(n4574), .B(n4573), .Z(c[297]) );
  XOR U6383 ( .A(n4576), .B(n4575), .Z(c[298]) );
  XOR U6384 ( .A(n4578), .B(n4577), .Z(c[299]) );
  XOR U6385 ( .A(n4580), .B(n4579), .Z(c[29]) );
  XOR U6386 ( .A(n4582), .B(n4581), .Z(c[2]) );
  XOR U6387 ( .A(n4584), .B(n4583), .Z(c[300]) );
  XOR U6388 ( .A(n4586), .B(n4585), .Z(c[301]) );
  XOR U6389 ( .A(n4588), .B(n4587), .Z(c[302]) );
  XOR U6390 ( .A(n4590), .B(n4589), .Z(c[303]) );
  XOR U6391 ( .A(n4592), .B(n4591), .Z(c[304]) );
  XOR U6392 ( .A(n4594), .B(n4593), .Z(c[305]) );
  XOR U6393 ( .A(n4596), .B(n4595), .Z(c[306]) );
  XOR U6394 ( .A(n4598), .B(n4597), .Z(c[307]) );
  XOR U6395 ( .A(n4600), .B(n4599), .Z(c[308]) );
  XOR U6396 ( .A(n4602), .B(n4601), .Z(c[309]) );
  XOR U6397 ( .A(n4604), .B(n4603), .Z(c[30]) );
  XOR U6398 ( .A(n4606), .B(n4605), .Z(c[310]) );
  XOR U6399 ( .A(n4608), .B(n4607), .Z(c[311]) );
  XOR U6400 ( .A(n4610), .B(n4609), .Z(c[312]) );
  XOR U6401 ( .A(n4612), .B(n4611), .Z(c[313]) );
  XOR U6402 ( .A(n4614), .B(n4613), .Z(c[314]) );
  XOR U6403 ( .A(n4616), .B(n4615), .Z(c[315]) );
  XOR U6404 ( .A(n4618), .B(n4617), .Z(c[316]) );
  XOR U6405 ( .A(n4620), .B(n4619), .Z(c[317]) );
  XOR U6406 ( .A(n4622), .B(n4621), .Z(c[318]) );
  XOR U6407 ( .A(n4624), .B(n4623), .Z(c[319]) );
  XOR U6408 ( .A(n4626), .B(n4625), .Z(c[31]) );
  XOR U6409 ( .A(n4628), .B(n4627), .Z(c[320]) );
  XOR U6410 ( .A(n4630), .B(n4629), .Z(c[321]) );
  XOR U6411 ( .A(n4632), .B(n4631), .Z(c[322]) );
  XOR U6412 ( .A(n4634), .B(n4633), .Z(c[323]) );
  XOR U6413 ( .A(n4636), .B(n4635), .Z(c[324]) );
  XOR U6414 ( .A(n4638), .B(n4637), .Z(c[325]) );
  XOR U6415 ( .A(n4640), .B(n4639), .Z(c[326]) );
  XOR U6416 ( .A(n4642), .B(n4641), .Z(c[327]) );
  XOR U6417 ( .A(n4644), .B(n4643), .Z(c[328]) );
  XOR U6418 ( .A(n4646), .B(n4645), .Z(c[329]) );
  XOR U6419 ( .A(n4648), .B(n4647), .Z(c[32]) );
  XOR U6420 ( .A(n4650), .B(n4649), .Z(c[330]) );
  XOR U6421 ( .A(n4652), .B(n4651), .Z(c[331]) );
  XOR U6422 ( .A(n4654), .B(n4653), .Z(c[332]) );
  XOR U6423 ( .A(n4656), .B(n4655), .Z(c[333]) );
  XOR U6424 ( .A(n4658), .B(n4657), .Z(c[334]) );
  XOR U6425 ( .A(n4660), .B(n4659), .Z(c[335]) );
  XOR U6426 ( .A(n4662), .B(n4661), .Z(c[336]) );
  XOR U6427 ( .A(n4664), .B(n4663), .Z(c[337]) );
  XOR U6428 ( .A(n4666), .B(n4665), .Z(c[338]) );
  XOR U6429 ( .A(n4668), .B(n4667), .Z(c[339]) );
  XOR U6430 ( .A(n4670), .B(n4669), .Z(c[33]) );
  XOR U6431 ( .A(n4672), .B(n4671), .Z(c[340]) );
  XOR U6432 ( .A(n4674), .B(n4673), .Z(c[341]) );
  XOR U6433 ( .A(n4676), .B(n4675), .Z(c[342]) );
  XOR U6434 ( .A(n4678), .B(n4677), .Z(c[343]) );
  XOR U6435 ( .A(n4680), .B(n4679), .Z(c[344]) );
  XOR U6436 ( .A(n4682), .B(n4681), .Z(c[345]) );
  XOR U6437 ( .A(n4684), .B(n4683), .Z(c[346]) );
  XOR U6438 ( .A(n4686), .B(n4685), .Z(c[347]) );
  XOR U6439 ( .A(n4688), .B(n4687), .Z(c[348]) );
  XOR U6440 ( .A(n4690), .B(n4689), .Z(c[349]) );
  XOR U6441 ( .A(n4692), .B(n4691), .Z(c[34]) );
  XOR U6442 ( .A(n4694), .B(n4693), .Z(c[350]) );
  XOR U6443 ( .A(n4696), .B(n4695), .Z(c[351]) );
  XOR U6444 ( .A(n4698), .B(n4697), .Z(c[352]) );
  XOR U6445 ( .A(n4700), .B(n4699), .Z(c[353]) );
  XOR U6446 ( .A(n4702), .B(n4701), .Z(c[354]) );
  XOR U6447 ( .A(n4704), .B(n4703), .Z(c[355]) );
  XOR U6448 ( .A(n4706), .B(n4705), .Z(c[356]) );
  XOR U6449 ( .A(n4708), .B(n4707), .Z(c[357]) );
  XOR U6450 ( .A(n4710), .B(n4709), .Z(c[358]) );
  XOR U6451 ( .A(n4712), .B(n4711), .Z(c[359]) );
  XOR U6452 ( .A(n4714), .B(n4713), .Z(c[35]) );
  XOR U6453 ( .A(n4716), .B(n4715), .Z(c[360]) );
  XOR U6454 ( .A(n4718), .B(n4717), .Z(c[361]) );
  XOR U6455 ( .A(n4720), .B(n4719), .Z(c[362]) );
  XOR U6456 ( .A(n4722), .B(n4721), .Z(c[363]) );
  XOR U6457 ( .A(n4724), .B(n4723), .Z(c[364]) );
  XOR U6458 ( .A(n4726), .B(n4725), .Z(c[365]) );
  XOR U6459 ( .A(n4728), .B(n4727), .Z(c[366]) );
  XOR U6460 ( .A(n4730), .B(n4729), .Z(c[367]) );
  XOR U6461 ( .A(n4732), .B(n4731), .Z(c[368]) );
  XOR U6462 ( .A(n4734), .B(n4733), .Z(c[369]) );
  XOR U6463 ( .A(n4736), .B(n4735), .Z(c[36]) );
  XOR U6464 ( .A(n4738), .B(n4737), .Z(c[370]) );
  XOR U6465 ( .A(n4740), .B(n4739), .Z(c[371]) );
  XOR U6466 ( .A(n4742), .B(n4741), .Z(c[372]) );
  XOR U6467 ( .A(n4744), .B(n4743), .Z(c[373]) );
  XOR U6468 ( .A(n4746), .B(n4745), .Z(c[374]) );
  XOR U6469 ( .A(n4748), .B(n4747), .Z(c[375]) );
  XOR U6470 ( .A(n4750), .B(n4749), .Z(c[376]) );
  XOR U6471 ( .A(n4752), .B(n4751), .Z(c[377]) );
  XOR U6472 ( .A(n4754), .B(n4753), .Z(c[378]) );
  XOR U6473 ( .A(n4756), .B(n4755), .Z(c[379]) );
  XOR U6474 ( .A(n4758), .B(n4757), .Z(c[37]) );
  XOR U6475 ( .A(n4760), .B(n4759), .Z(c[380]) );
  XOR U6476 ( .A(n4762), .B(n4761), .Z(c[381]) );
  XOR U6477 ( .A(n4764), .B(n4763), .Z(c[382]) );
  XOR U6478 ( .A(n4766), .B(n4765), .Z(c[383]) );
  XOR U6479 ( .A(n4768), .B(n4767), .Z(c[384]) );
  XOR U6480 ( .A(n4770), .B(n4769), .Z(c[385]) );
  XOR U6481 ( .A(n4772), .B(n4771), .Z(c[386]) );
  XOR U6482 ( .A(n4774), .B(n4773), .Z(c[387]) );
  XOR U6483 ( .A(n4776), .B(n4775), .Z(c[388]) );
  XOR U6484 ( .A(n4778), .B(n4777), .Z(c[389]) );
  XOR U6485 ( .A(n4780), .B(n4779), .Z(c[38]) );
  XOR U6486 ( .A(n4782), .B(n4781), .Z(c[390]) );
  XOR U6487 ( .A(n4784), .B(n4783), .Z(c[391]) );
  XOR U6488 ( .A(n4786), .B(n4785), .Z(c[392]) );
  XOR U6489 ( .A(n4788), .B(n4787), .Z(c[393]) );
  XOR U6490 ( .A(n4790), .B(n4789), .Z(c[394]) );
  XOR U6491 ( .A(n4792), .B(n4791), .Z(c[395]) );
  XOR U6492 ( .A(n4794), .B(n4793), .Z(c[396]) );
  XOR U6493 ( .A(n4796), .B(n4795), .Z(c[397]) );
  XOR U6494 ( .A(n4798), .B(n4797), .Z(c[398]) );
  XOR U6495 ( .A(n4800), .B(n4799), .Z(c[399]) );
  XOR U6496 ( .A(n4802), .B(n4801), .Z(c[39]) );
  XOR U6497 ( .A(n4804), .B(n4803), .Z(c[3]) );
  XOR U6498 ( .A(n4806), .B(n4805), .Z(c[400]) );
  XOR U6499 ( .A(n4808), .B(n4807), .Z(c[401]) );
  XOR U6500 ( .A(n4810), .B(n4809), .Z(c[402]) );
  XOR U6501 ( .A(n4812), .B(n4811), .Z(c[403]) );
  XOR U6502 ( .A(n4814), .B(n4813), .Z(c[404]) );
  XOR U6503 ( .A(n4816), .B(n4815), .Z(c[405]) );
  XOR U6504 ( .A(n4818), .B(n4817), .Z(c[406]) );
  XOR U6505 ( .A(n4820), .B(n4819), .Z(c[407]) );
  XOR U6506 ( .A(n4822), .B(n4821), .Z(c[408]) );
  XOR U6507 ( .A(n4824), .B(n4823), .Z(c[409]) );
  XOR U6508 ( .A(n4826), .B(n4825), .Z(c[40]) );
  XOR U6509 ( .A(n4828), .B(n4827), .Z(c[410]) );
  XOR U6510 ( .A(n4830), .B(n4829), .Z(c[411]) );
  XOR U6511 ( .A(n4832), .B(n4831), .Z(c[412]) );
  XOR U6512 ( .A(n4834), .B(n4833), .Z(c[413]) );
  XOR U6513 ( .A(n4836), .B(n4835), .Z(c[414]) );
  XOR U6514 ( .A(n4838), .B(n4837), .Z(c[415]) );
  XOR U6515 ( .A(n4840), .B(n4839), .Z(c[416]) );
  XOR U6516 ( .A(n4842), .B(n4841), .Z(c[417]) );
  XOR U6517 ( .A(n4844), .B(n4843), .Z(c[418]) );
  XOR U6518 ( .A(n4846), .B(n4845), .Z(c[419]) );
  XOR U6519 ( .A(n4848), .B(n4847), .Z(c[41]) );
  XOR U6520 ( .A(n4850), .B(n4849), .Z(c[420]) );
  XOR U6521 ( .A(n4852), .B(n4851), .Z(c[421]) );
  XOR U6522 ( .A(n4854), .B(n4853), .Z(c[422]) );
  XOR U6523 ( .A(n4856), .B(n4855), .Z(c[423]) );
  XOR U6524 ( .A(n4858), .B(n4857), .Z(c[424]) );
  XOR U6525 ( .A(n4860), .B(n4859), .Z(c[425]) );
  XOR U6526 ( .A(n4862), .B(n4861), .Z(c[426]) );
  XOR U6527 ( .A(n4864), .B(n4863), .Z(c[427]) );
  XOR U6528 ( .A(n4866), .B(n4865), .Z(c[428]) );
  XOR U6529 ( .A(n4868), .B(n4867), .Z(c[429]) );
  XOR U6530 ( .A(n4870), .B(n4869), .Z(c[42]) );
  XOR U6531 ( .A(n4872), .B(n4871), .Z(c[430]) );
  XOR U6532 ( .A(n4874), .B(n4873), .Z(c[431]) );
  XOR U6533 ( .A(n4876), .B(n4875), .Z(c[432]) );
  XOR U6534 ( .A(n4878), .B(n4877), .Z(c[433]) );
  XOR U6535 ( .A(n4880), .B(n4879), .Z(c[434]) );
  XOR U6536 ( .A(n4882), .B(n4881), .Z(c[435]) );
  XOR U6537 ( .A(n4884), .B(n4883), .Z(c[436]) );
  XOR U6538 ( .A(n4886), .B(n4885), .Z(c[437]) );
  XOR U6539 ( .A(n4888), .B(n4887), .Z(c[438]) );
  XOR U6540 ( .A(n4890), .B(n4889), .Z(c[439]) );
  XOR U6541 ( .A(n4892), .B(n4891), .Z(c[43]) );
  XOR U6542 ( .A(n4894), .B(n4893), .Z(c[440]) );
  XOR U6543 ( .A(n4896), .B(n4895), .Z(c[441]) );
  XOR U6544 ( .A(n4898), .B(n4897), .Z(c[442]) );
  XOR U6545 ( .A(n4900), .B(n4899), .Z(c[443]) );
  XOR U6546 ( .A(n4902), .B(n4901), .Z(c[444]) );
  XOR U6547 ( .A(n4904), .B(n4903), .Z(c[445]) );
  XOR U6548 ( .A(n4906), .B(n4905), .Z(c[446]) );
  XOR U6549 ( .A(n4908), .B(n4907), .Z(c[447]) );
  XOR U6550 ( .A(n4910), .B(n4909), .Z(c[448]) );
  XOR U6551 ( .A(n4912), .B(n4911), .Z(c[449]) );
  XOR U6552 ( .A(n4914), .B(n4913), .Z(c[44]) );
  XOR U6553 ( .A(n4916), .B(n4915), .Z(c[450]) );
  XOR U6554 ( .A(n4918), .B(n4917), .Z(c[451]) );
  XOR U6555 ( .A(n4920), .B(n4919), .Z(c[452]) );
  XOR U6556 ( .A(n4922), .B(n4921), .Z(c[453]) );
  XOR U6557 ( .A(n4924), .B(n4923), .Z(c[454]) );
  XOR U6558 ( .A(n4926), .B(n4925), .Z(c[455]) );
  XOR U6559 ( .A(n4928), .B(n4927), .Z(c[456]) );
  XOR U6560 ( .A(n4930), .B(n4929), .Z(c[457]) );
  XOR U6561 ( .A(n4932), .B(n4931), .Z(c[458]) );
  XOR U6562 ( .A(n4934), .B(n4933), .Z(c[459]) );
  XOR U6563 ( .A(n4936), .B(n4935), .Z(c[45]) );
  XOR U6564 ( .A(n4938), .B(n4937), .Z(c[460]) );
  XOR U6565 ( .A(n4940), .B(n4939), .Z(c[461]) );
  XOR U6566 ( .A(n4942), .B(n4941), .Z(c[462]) );
  XOR U6567 ( .A(n4944), .B(n4943), .Z(c[463]) );
  XOR U6568 ( .A(n4946), .B(n4945), .Z(c[464]) );
  XOR U6569 ( .A(n4948), .B(n4947), .Z(c[465]) );
  XOR U6570 ( .A(n4950), .B(n4949), .Z(c[466]) );
  XOR U6571 ( .A(n4952), .B(n4951), .Z(c[467]) );
  XOR U6572 ( .A(n4954), .B(n4953), .Z(c[468]) );
  XOR U6573 ( .A(n4956), .B(n4955), .Z(c[469]) );
  XOR U6574 ( .A(n4958), .B(n4957), .Z(c[46]) );
  XOR U6575 ( .A(n4960), .B(n4959), .Z(c[470]) );
  XOR U6576 ( .A(n4962), .B(n4961), .Z(c[471]) );
  XOR U6577 ( .A(n4964), .B(n4963), .Z(c[472]) );
  XOR U6578 ( .A(n4966), .B(n4965), .Z(c[473]) );
  XOR U6579 ( .A(n4968), .B(n4967), .Z(c[474]) );
  XOR U6580 ( .A(n4970), .B(n4969), .Z(c[475]) );
  XOR U6581 ( .A(n4972), .B(n4971), .Z(c[476]) );
  XOR U6582 ( .A(n4974), .B(n4973), .Z(c[477]) );
  XOR U6583 ( .A(n4976), .B(n4975), .Z(c[478]) );
  XOR U6584 ( .A(n4978), .B(n4977), .Z(c[479]) );
  XOR U6585 ( .A(n4980), .B(n4979), .Z(c[47]) );
  XOR U6586 ( .A(n4982), .B(n4981), .Z(c[480]) );
  XOR U6587 ( .A(n4984), .B(n4983), .Z(c[481]) );
  XOR U6588 ( .A(n4986), .B(n4985), .Z(c[482]) );
  XOR U6589 ( .A(n4988), .B(n4987), .Z(c[483]) );
  XOR U6590 ( .A(n4990), .B(n4989), .Z(c[484]) );
  XOR U6591 ( .A(n4992), .B(n4991), .Z(c[485]) );
  XOR U6592 ( .A(n4994), .B(n4993), .Z(c[486]) );
  XOR U6593 ( .A(n4996), .B(n4995), .Z(c[487]) );
  XOR U6594 ( .A(n4998), .B(n4997), .Z(c[488]) );
  XOR U6595 ( .A(n5000), .B(n4999), .Z(c[489]) );
  XOR U6596 ( .A(n5002), .B(n5001), .Z(c[48]) );
  XOR U6597 ( .A(n5004), .B(n5003), .Z(c[490]) );
  XOR U6598 ( .A(n5006), .B(n5005), .Z(c[491]) );
  XOR U6599 ( .A(n5008), .B(n5007), .Z(c[492]) );
  XOR U6600 ( .A(n5010), .B(n5009), .Z(c[493]) );
  XOR U6601 ( .A(n5012), .B(n5011), .Z(c[494]) );
  XOR U6602 ( .A(n5014), .B(n5013), .Z(c[495]) );
  XOR U6603 ( .A(n5016), .B(n5015), .Z(c[496]) );
  XOR U6604 ( .A(n5018), .B(n5017), .Z(c[497]) );
  XOR U6605 ( .A(n5020), .B(n5019), .Z(c[498]) );
  XOR U6606 ( .A(n5022), .B(n5021), .Z(c[499]) );
  XOR U6607 ( .A(n5024), .B(n5023), .Z(c[49]) );
  XOR U6608 ( .A(n5026), .B(n5025), .Z(c[4]) );
  XOR U6609 ( .A(n5028), .B(n5027), .Z(c[500]) );
  XOR U6610 ( .A(n5030), .B(n5029), .Z(c[501]) );
  XOR U6611 ( .A(n5032), .B(n5031), .Z(c[502]) );
  XOR U6612 ( .A(n5034), .B(n5033), .Z(c[503]) );
  XOR U6613 ( .A(n5036), .B(n5035), .Z(c[504]) );
  XOR U6614 ( .A(n5038), .B(n5037), .Z(c[505]) );
  XOR U6615 ( .A(n5040), .B(n5039), .Z(c[506]) );
  XOR U6616 ( .A(n5042), .B(n5041), .Z(c[507]) );
  XOR U6617 ( .A(n5044), .B(n5043), .Z(c[508]) );
  XOR U6618 ( .A(n5046), .B(n5045), .Z(c[509]) );
  XOR U6619 ( .A(n5048), .B(n5047), .Z(c[50]) );
  XOR U6620 ( .A(n5050), .B(n5049), .Z(c[510]) );
  XOR U6621 ( .A(n5052), .B(n5051), .Z(c[511]) );
  XOR U6622 ( .A(n5054), .B(n5053), .Z(c[512]) );
  XOR U6623 ( .A(n5056), .B(n5055), .Z(c[513]) );
  XOR U6624 ( .A(n5058), .B(n5057), .Z(c[514]) );
  XOR U6625 ( .A(n5060), .B(n5059), .Z(c[515]) );
  XOR U6626 ( .A(n5062), .B(n5061), .Z(c[516]) );
  XOR U6627 ( .A(n5064), .B(n5063), .Z(c[517]) );
  XOR U6628 ( .A(n5066), .B(n5065), .Z(c[518]) );
  XOR U6629 ( .A(n5068), .B(n5067), .Z(c[519]) );
  XOR U6630 ( .A(n5070), .B(n5069), .Z(c[51]) );
  XOR U6631 ( .A(n5072), .B(n5071), .Z(c[520]) );
  XOR U6632 ( .A(n5074), .B(n5073), .Z(c[521]) );
  XOR U6633 ( .A(n5076), .B(n5075), .Z(c[522]) );
  XOR U6634 ( .A(n5078), .B(n5077), .Z(c[523]) );
  XOR U6635 ( .A(n5080), .B(n5079), .Z(c[524]) );
  XOR U6636 ( .A(n5082), .B(n5081), .Z(c[525]) );
  XOR U6637 ( .A(n5084), .B(n5083), .Z(c[526]) );
  XOR U6638 ( .A(n5086), .B(n5085), .Z(c[527]) );
  XOR U6639 ( .A(n5088), .B(n5087), .Z(c[528]) );
  XOR U6640 ( .A(n5090), .B(n5089), .Z(c[529]) );
  XOR U6641 ( .A(n5092), .B(n5091), .Z(c[52]) );
  XOR U6642 ( .A(n5094), .B(n5093), .Z(c[530]) );
  XOR U6643 ( .A(n5096), .B(n5095), .Z(c[531]) );
  XOR U6644 ( .A(n5098), .B(n5097), .Z(c[532]) );
  XOR U6645 ( .A(n5100), .B(n5099), .Z(c[533]) );
  XOR U6646 ( .A(n5102), .B(n5101), .Z(c[534]) );
  XOR U6647 ( .A(n5104), .B(n5103), .Z(c[535]) );
  XOR U6648 ( .A(n5106), .B(n5105), .Z(c[536]) );
  XOR U6649 ( .A(n5108), .B(n5107), .Z(c[537]) );
  XOR U6650 ( .A(n5110), .B(n5109), .Z(c[538]) );
  XOR U6651 ( .A(n5112), .B(n5111), .Z(c[539]) );
  XOR U6652 ( .A(n5114), .B(n5113), .Z(c[53]) );
  XOR U6653 ( .A(n5116), .B(n5115), .Z(c[540]) );
  XOR U6654 ( .A(n5118), .B(n5117), .Z(c[541]) );
  XOR U6655 ( .A(n5120), .B(n5119), .Z(c[542]) );
  XOR U6656 ( .A(n5122), .B(n5121), .Z(c[543]) );
  XOR U6657 ( .A(n5124), .B(n5123), .Z(c[544]) );
  XOR U6658 ( .A(n5126), .B(n5125), .Z(c[545]) );
  XOR U6659 ( .A(n5128), .B(n5127), .Z(c[546]) );
  XOR U6660 ( .A(n5130), .B(n5129), .Z(c[547]) );
  XOR U6661 ( .A(n5132), .B(n5131), .Z(c[548]) );
  XOR U6662 ( .A(n5134), .B(n5133), .Z(c[549]) );
  XOR U6663 ( .A(n5136), .B(n5135), .Z(c[54]) );
  XOR U6664 ( .A(n5138), .B(n5137), .Z(c[550]) );
  XOR U6665 ( .A(n5140), .B(n5139), .Z(c[551]) );
  XOR U6666 ( .A(n5142), .B(n5141), .Z(c[552]) );
  XOR U6667 ( .A(n5144), .B(n5143), .Z(c[553]) );
  XOR U6668 ( .A(n5146), .B(n5145), .Z(c[554]) );
  XOR U6669 ( .A(n5148), .B(n5147), .Z(c[555]) );
  XOR U6670 ( .A(n5150), .B(n5149), .Z(c[556]) );
  XOR U6671 ( .A(n5152), .B(n5151), .Z(c[557]) );
  XOR U6672 ( .A(n5154), .B(n5153), .Z(c[558]) );
  XOR U6673 ( .A(n5156), .B(n5155), .Z(c[559]) );
  XOR U6674 ( .A(n5158), .B(n5157), .Z(c[55]) );
  XOR U6675 ( .A(n5160), .B(n5159), .Z(c[560]) );
  XOR U6676 ( .A(n5162), .B(n5161), .Z(c[561]) );
  XOR U6677 ( .A(n5164), .B(n5163), .Z(c[562]) );
  XOR U6678 ( .A(n5166), .B(n5165), .Z(c[563]) );
  XOR U6679 ( .A(n5168), .B(n5167), .Z(c[564]) );
  XOR U6680 ( .A(n5170), .B(n5169), .Z(c[565]) );
  XOR U6681 ( .A(n5172), .B(n5171), .Z(c[566]) );
  XOR U6682 ( .A(n5174), .B(n5173), .Z(c[567]) );
  XOR U6683 ( .A(n5176), .B(n5175), .Z(c[568]) );
  XOR U6684 ( .A(n5178), .B(n5177), .Z(c[569]) );
  XOR U6685 ( .A(n5180), .B(n5179), .Z(c[56]) );
  XOR U6686 ( .A(n5182), .B(n5181), .Z(c[570]) );
  XOR U6687 ( .A(n5184), .B(n5183), .Z(c[571]) );
  XOR U6688 ( .A(n5186), .B(n5185), .Z(c[572]) );
  XOR U6689 ( .A(n5188), .B(n5187), .Z(c[573]) );
  XOR U6690 ( .A(n5190), .B(n5189), .Z(c[574]) );
  XOR U6691 ( .A(n5192), .B(n5191), .Z(c[575]) );
  XOR U6692 ( .A(n5194), .B(n5193), .Z(c[576]) );
  XOR U6693 ( .A(n5196), .B(n5195), .Z(c[577]) );
  XOR U6694 ( .A(n5198), .B(n5197), .Z(c[578]) );
  XOR U6695 ( .A(n5200), .B(n5199), .Z(c[579]) );
  XOR U6696 ( .A(n5202), .B(n5201), .Z(c[57]) );
  XOR U6697 ( .A(n5204), .B(n5203), .Z(c[580]) );
  XOR U6698 ( .A(n5206), .B(n5205), .Z(c[581]) );
  XOR U6699 ( .A(n5208), .B(n5207), .Z(c[582]) );
  XOR U6700 ( .A(n5210), .B(n5209), .Z(c[583]) );
  XOR U6701 ( .A(n5212), .B(n5211), .Z(c[584]) );
  XOR U6702 ( .A(n5214), .B(n5213), .Z(c[585]) );
  XOR U6703 ( .A(n5216), .B(n5215), .Z(c[586]) );
  XOR U6704 ( .A(n5218), .B(n5217), .Z(c[587]) );
  XOR U6705 ( .A(n5220), .B(n5219), .Z(c[588]) );
  XOR U6706 ( .A(n5222), .B(n5221), .Z(c[589]) );
  XOR U6707 ( .A(n5224), .B(n5223), .Z(c[58]) );
  XOR U6708 ( .A(n5226), .B(n5225), .Z(c[590]) );
  XOR U6709 ( .A(n5228), .B(n5227), .Z(c[591]) );
  XOR U6710 ( .A(n5230), .B(n5229), .Z(c[592]) );
  XOR U6711 ( .A(n5232), .B(n5231), .Z(c[593]) );
  XOR U6712 ( .A(n5234), .B(n5233), .Z(c[594]) );
  XOR U6713 ( .A(n5236), .B(n5235), .Z(c[595]) );
  XOR U6714 ( .A(n5238), .B(n5237), .Z(c[596]) );
  XOR U6715 ( .A(n5240), .B(n5239), .Z(c[597]) );
  XOR U6716 ( .A(n5242), .B(n5241), .Z(c[598]) );
  XOR U6717 ( .A(n5244), .B(n5243), .Z(c[599]) );
  XOR U6718 ( .A(n5246), .B(n5245), .Z(c[59]) );
  XOR U6719 ( .A(n5248), .B(n5247), .Z(c[5]) );
  XOR U6720 ( .A(n5250), .B(n5249), .Z(c[600]) );
  XOR U6721 ( .A(n5252), .B(n5251), .Z(c[601]) );
  XOR U6722 ( .A(n5254), .B(n5253), .Z(c[602]) );
  XOR U6723 ( .A(n5256), .B(n5255), .Z(c[603]) );
  XOR U6724 ( .A(n5258), .B(n5257), .Z(c[604]) );
  XOR U6725 ( .A(n5260), .B(n5259), .Z(c[605]) );
  XOR U6726 ( .A(n5262), .B(n5261), .Z(c[606]) );
  XOR U6727 ( .A(n5264), .B(n5263), .Z(c[607]) );
  XOR U6728 ( .A(n5266), .B(n5265), .Z(c[608]) );
  XOR U6729 ( .A(n5268), .B(n5267), .Z(c[609]) );
  XOR U6730 ( .A(n5270), .B(n5269), .Z(c[60]) );
  XOR U6731 ( .A(n5272), .B(n5271), .Z(c[610]) );
  XOR U6732 ( .A(n5274), .B(n5273), .Z(c[611]) );
  XOR U6733 ( .A(n5276), .B(n5275), .Z(c[612]) );
  XOR U6734 ( .A(n5278), .B(n5277), .Z(c[613]) );
  XOR U6735 ( .A(n5280), .B(n5279), .Z(c[614]) );
  XOR U6736 ( .A(n5282), .B(n5281), .Z(c[615]) );
  XOR U6737 ( .A(n5284), .B(n5283), .Z(c[616]) );
  XOR U6738 ( .A(n5286), .B(n5285), .Z(c[617]) );
  XOR U6739 ( .A(n5288), .B(n5287), .Z(c[618]) );
  XOR U6740 ( .A(n5290), .B(n5289), .Z(c[619]) );
  XOR U6741 ( .A(n5292), .B(n5291), .Z(c[61]) );
  XOR U6742 ( .A(n5294), .B(n5293), .Z(c[620]) );
  XOR U6743 ( .A(n5296), .B(n5295), .Z(c[621]) );
  XOR U6744 ( .A(n5298), .B(n5297), .Z(c[622]) );
  XOR U6745 ( .A(n5300), .B(n5299), .Z(c[623]) );
  XOR U6746 ( .A(n5302), .B(n5301), .Z(c[624]) );
  XOR U6747 ( .A(n5304), .B(n5303), .Z(c[625]) );
  XOR U6748 ( .A(n5306), .B(n5305), .Z(c[626]) );
  XOR U6749 ( .A(n5308), .B(n5307), .Z(c[627]) );
  XOR U6750 ( .A(n5310), .B(n5309), .Z(c[628]) );
  XOR U6751 ( .A(n5312), .B(n5311), .Z(c[629]) );
  XOR U6752 ( .A(n5314), .B(n5313), .Z(c[62]) );
  XOR U6753 ( .A(n5316), .B(n5315), .Z(c[630]) );
  XOR U6754 ( .A(n5318), .B(n5317), .Z(c[631]) );
  XOR U6755 ( .A(n5320), .B(n5319), .Z(c[632]) );
  XOR U6756 ( .A(n5322), .B(n5321), .Z(c[633]) );
  XOR U6757 ( .A(n5324), .B(n5323), .Z(c[634]) );
  XOR U6758 ( .A(n5326), .B(n5325), .Z(c[635]) );
  XOR U6759 ( .A(n5328), .B(n5327), .Z(c[636]) );
  XOR U6760 ( .A(n5330), .B(n5329), .Z(c[637]) );
  XOR U6761 ( .A(n5332), .B(n5331), .Z(c[638]) );
  XOR U6762 ( .A(n5334), .B(n5333), .Z(c[639]) );
  XOR U6763 ( .A(n5336), .B(n5335), .Z(c[63]) );
  XOR U6764 ( .A(n5338), .B(n5337), .Z(c[640]) );
  XOR U6765 ( .A(n5340), .B(n5339), .Z(c[641]) );
  XOR U6766 ( .A(n5342), .B(n5341), .Z(c[642]) );
  XOR U6767 ( .A(n5344), .B(n5343), .Z(c[643]) );
  XOR U6768 ( .A(n5346), .B(n5345), .Z(c[644]) );
  XOR U6769 ( .A(n5348), .B(n5347), .Z(c[645]) );
  XOR U6770 ( .A(n5350), .B(n5349), .Z(c[646]) );
  XOR U6771 ( .A(n5352), .B(n5351), .Z(c[647]) );
  XOR U6772 ( .A(n5354), .B(n5353), .Z(c[648]) );
  XOR U6773 ( .A(n5356), .B(n5355), .Z(c[649]) );
  XOR U6774 ( .A(n5358), .B(n5357), .Z(c[64]) );
  XOR U6775 ( .A(n5360), .B(n5359), .Z(c[650]) );
  XOR U6776 ( .A(n5362), .B(n5361), .Z(c[651]) );
  XOR U6777 ( .A(n5364), .B(n5363), .Z(c[652]) );
  XOR U6778 ( .A(n5366), .B(n5365), .Z(c[653]) );
  XOR U6779 ( .A(n5368), .B(n5367), .Z(c[654]) );
  XOR U6780 ( .A(n5370), .B(n5369), .Z(c[655]) );
  XOR U6781 ( .A(n5372), .B(n5371), .Z(c[656]) );
  XOR U6782 ( .A(n5374), .B(n5373), .Z(c[657]) );
  XOR U6783 ( .A(n5376), .B(n5375), .Z(c[658]) );
  XOR U6784 ( .A(n5378), .B(n5377), .Z(c[659]) );
  XOR U6785 ( .A(n5380), .B(n5379), .Z(c[65]) );
  XOR U6786 ( .A(n5382), .B(n5381), .Z(c[660]) );
  XOR U6787 ( .A(n5384), .B(n5383), .Z(c[661]) );
  XOR U6788 ( .A(n5386), .B(n5385), .Z(c[662]) );
  XOR U6789 ( .A(n5388), .B(n5387), .Z(c[663]) );
  XOR U6790 ( .A(n5390), .B(n5389), .Z(c[664]) );
  XOR U6791 ( .A(n5392), .B(n5391), .Z(c[665]) );
  XOR U6792 ( .A(n5394), .B(n5393), .Z(c[666]) );
  XOR U6793 ( .A(n5396), .B(n5395), .Z(c[667]) );
  XOR U6794 ( .A(n5398), .B(n5397), .Z(c[668]) );
  XOR U6795 ( .A(n5400), .B(n5399), .Z(c[669]) );
  XOR U6796 ( .A(n5402), .B(n5401), .Z(c[66]) );
  XOR U6797 ( .A(n5404), .B(n5403), .Z(c[670]) );
  XOR U6798 ( .A(n5406), .B(n5405), .Z(c[671]) );
  XOR U6799 ( .A(n5408), .B(n5407), .Z(c[672]) );
  XOR U6800 ( .A(n5410), .B(n5409), .Z(c[673]) );
  XOR U6801 ( .A(n5412), .B(n5411), .Z(c[674]) );
  XOR U6802 ( .A(n5414), .B(n5413), .Z(c[675]) );
  XOR U6803 ( .A(n5416), .B(n5415), .Z(c[676]) );
  XOR U6804 ( .A(n5418), .B(n5417), .Z(c[677]) );
  XOR U6805 ( .A(n5420), .B(n5419), .Z(c[678]) );
  XOR U6806 ( .A(n5422), .B(n5421), .Z(c[679]) );
  XOR U6807 ( .A(n5424), .B(n5423), .Z(c[67]) );
  XOR U6808 ( .A(n5426), .B(n5425), .Z(c[680]) );
  XOR U6809 ( .A(n5428), .B(n5427), .Z(c[681]) );
  XOR U6810 ( .A(n5430), .B(n5429), .Z(c[682]) );
  XOR U6811 ( .A(n5432), .B(n5431), .Z(c[683]) );
  XOR U6812 ( .A(n5434), .B(n5433), .Z(c[684]) );
  XOR U6813 ( .A(n5436), .B(n5435), .Z(c[685]) );
  XOR U6814 ( .A(n5438), .B(n5437), .Z(c[686]) );
  XOR U6815 ( .A(n5440), .B(n5439), .Z(c[687]) );
  XOR U6816 ( .A(n5442), .B(n5441), .Z(c[688]) );
  XOR U6817 ( .A(n5444), .B(n5443), .Z(c[689]) );
  XOR U6818 ( .A(n5446), .B(n5445), .Z(c[68]) );
  XOR U6819 ( .A(n5448), .B(n5447), .Z(c[690]) );
  XOR U6820 ( .A(n5450), .B(n5449), .Z(c[691]) );
  XOR U6821 ( .A(n5452), .B(n5451), .Z(c[692]) );
  XOR U6822 ( .A(n5454), .B(n5453), .Z(c[693]) );
  XOR U6823 ( .A(n5456), .B(n5455), .Z(c[694]) );
  XOR U6824 ( .A(n5458), .B(n5457), .Z(c[695]) );
  XOR U6825 ( .A(n5460), .B(n5459), .Z(c[696]) );
  XOR U6826 ( .A(n5462), .B(n5461), .Z(c[697]) );
  XOR U6827 ( .A(n5464), .B(n5463), .Z(c[698]) );
  XOR U6828 ( .A(n5466), .B(n5465), .Z(c[699]) );
  XOR U6829 ( .A(n5468), .B(n5467), .Z(c[69]) );
  XOR U6830 ( .A(n5470), .B(n5469), .Z(c[6]) );
  XOR U6831 ( .A(n5472), .B(n5471), .Z(c[700]) );
  XOR U6832 ( .A(n5474), .B(n5473), .Z(c[701]) );
  XOR U6833 ( .A(n5476), .B(n5475), .Z(c[702]) );
  XOR U6834 ( .A(n5478), .B(n5477), .Z(c[703]) );
  XOR U6835 ( .A(n5480), .B(n5479), .Z(c[704]) );
  XOR U6836 ( .A(n5482), .B(n5481), .Z(c[705]) );
  XOR U6837 ( .A(n5484), .B(n5483), .Z(c[706]) );
  XOR U6838 ( .A(n5486), .B(n5485), .Z(c[707]) );
  XOR U6839 ( .A(n5488), .B(n5487), .Z(c[708]) );
  XOR U6840 ( .A(n5490), .B(n5489), .Z(c[709]) );
  XOR U6841 ( .A(n5492), .B(n5491), .Z(c[70]) );
  XOR U6842 ( .A(n5494), .B(n5493), .Z(c[710]) );
  XOR U6843 ( .A(n5496), .B(n5495), .Z(c[711]) );
  XOR U6844 ( .A(n5498), .B(n5497), .Z(c[712]) );
  XOR U6845 ( .A(n5500), .B(n5499), .Z(c[713]) );
  XOR U6846 ( .A(n5502), .B(n5501), .Z(c[714]) );
  XOR U6847 ( .A(n5504), .B(n5503), .Z(c[715]) );
  XOR U6848 ( .A(n5506), .B(n5505), .Z(c[716]) );
  XOR U6849 ( .A(n5508), .B(n5507), .Z(c[717]) );
  XOR U6850 ( .A(n5510), .B(n5509), .Z(c[718]) );
  XOR U6851 ( .A(n5512), .B(n5511), .Z(c[719]) );
  XOR U6852 ( .A(n5514), .B(n5513), .Z(c[71]) );
  XOR U6853 ( .A(n5516), .B(n5515), .Z(c[720]) );
  XOR U6854 ( .A(n5518), .B(n5517), .Z(c[721]) );
  XOR U6855 ( .A(n5520), .B(n5519), .Z(c[722]) );
  XOR U6856 ( .A(n5522), .B(n5521), .Z(c[723]) );
  XOR U6857 ( .A(n5524), .B(n5523), .Z(c[724]) );
  XOR U6858 ( .A(n5526), .B(n5525), .Z(c[725]) );
  XOR U6859 ( .A(n5528), .B(n5527), .Z(c[726]) );
  XOR U6860 ( .A(n5530), .B(n5529), .Z(c[727]) );
  XOR U6861 ( .A(n5532), .B(n5531), .Z(c[728]) );
  XOR U6862 ( .A(n5534), .B(n5533), .Z(c[729]) );
  XOR U6863 ( .A(n5536), .B(n5535), .Z(c[72]) );
  XOR U6864 ( .A(n5538), .B(n5537), .Z(c[730]) );
  XOR U6865 ( .A(n5540), .B(n5539), .Z(c[731]) );
  XOR U6866 ( .A(n5542), .B(n5541), .Z(c[732]) );
  XOR U6867 ( .A(n5544), .B(n5543), .Z(c[733]) );
  XOR U6868 ( .A(n5546), .B(n5545), .Z(c[734]) );
  XOR U6869 ( .A(n5548), .B(n5547), .Z(c[735]) );
  XOR U6870 ( .A(n5550), .B(n5549), .Z(c[736]) );
  XOR U6871 ( .A(n5552), .B(n5551), .Z(c[737]) );
  XOR U6872 ( .A(n5554), .B(n5553), .Z(c[738]) );
  XOR U6873 ( .A(n5556), .B(n5555), .Z(c[739]) );
  XOR U6874 ( .A(n5558), .B(n5557), .Z(c[73]) );
  XOR U6875 ( .A(n5560), .B(n5559), .Z(c[740]) );
  XOR U6876 ( .A(n5562), .B(n5561), .Z(c[741]) );
  XOR U6877 ( .A(n5564), .B(n5563), .Z(c[742]) );
  XOR U6878 ( .A(n5566), .B(n5565), .Z(c[743]) );
  XOR U6879 ( .A(n5568), .B(n5567), .Z(c[744]) );
  XOR U6880 ( .A(n5570), .B(n5569), .Z(c[745]) );
  XOR U6881 ( .A(n5572), .B(n5571), .Z(c[746]) );
  XOR U6882 ( .A(n5574), .B(n5573), .Z(c[747]) );
  XOR U6883 ( .A(n5576), .B(n5575), .Z(c[748]) );
  XOR U6884 ( .A(n5578), .B(n5577), .Z(c[749]) );
  XOR U6885 ( .A(n5580), .B(n5579), .Z(c[74]) );
  XOR U6886 ( .A(n5582), .B(n5581), .Z(c[750]) );
  XOR U6887 ( .A(n5584), .B(n5583), .Z(c[751]) );
  XOR U6888 ( .A(n5586), .B(n5585), .Z(c[752]) );
  XOR U6889 ( .A(n5588), .B(n5587), .Z(c[753]) );
  XOR U6890 ( .A(n5590), .B(n5589), .Z(c[754]) );
  XOR U6891 ( .A(n5592), .B(n5591), .Z(c[755]) );
  XOR U6892 ( .A(n5594), .B(n5593), .Z(c[756]) );
  XOR U6893 ( .A(n5596), .B(n5595), .Z(c[757]) );
  XOR U6894 ( .A(n5598), .B(n5597), .Z(c[758]) );
  XOR U6895 ( .A(n5600), .B(n5599), .Z(c[759]) );
  XOR U6896 ( .A(n5602), .B(n5601), .Z(c[75]) );
  XOR U6897 ( .A(n5604), .B(n5603), .Z(c[760]) );
  XOR U6898 ( .A(n5606), .B(n5605), .Z(c[761]) );
  XOR U6899 ( .A(n5608), .B(n5607), .Z(c[762]) );
  XOR U6900 ( .A(n5610), .B(n5609), .Z(c[763]) );
  XOR U6901 ( .A(n5612), .B(n5611), .Z(c[764]) );
  XOR U6902 ( .A(n5614), .B(n5613), .Z(c[765]) );
  XOR U6903 ( .A(n5616), .B(n5615), .Z(c[766]) );
  XOR U6904 ( .A(n5618), .B(n5617), .Z(c[767]) );
  XOR U6905 ( .A(n5620), .B(n5619), .Z(c[768]) );
  XOR U6906 ( .A(n5622), .B(n5621), .Z(c[769]) );
  XOR U6907 ( .A(n5624), .B(n5623), .Z(c[76]) );
  XOR U6908 ( .A(n5626), .B(n5625), .Z(c[770]) );
  XOR U6909 ( .A(n5628), .B(n5627), .Z(c[771]) );
  XOR U6910 ( .A(n5630), .B(n5629), .Z(c[772]) );
  XOR U6911 ( .A(n5632), .B(n5631), .Z(c[773]) );
  XOR U6912 ( .A(n5634), .B(n5633), .Z(c[774]) );
  XOR U6913 ( .A(n5636), .B(n5635), .Z(c[775]) );
  XOR U6914 ( .A(n5638), .B(n5637), .Z(c[776]) );
  XOR U6915 ( .A(n5640), .B(n5639), .Z(c[777]) );
  XOR U6916 ( .A(n5642), .B(n5641), .Z(c[778]) );
  XOR U6917 ( .A(n5644), .B(n5643), .Z(c[779]) );
  XOR U6918 ( .A(n5646), .B(n5645), .Z(c[77]) );
  XOR U6919 ( .A(n5648), .B(n5647), .Z(c[780]) );
  XOR U6920 ( .A(n5650), .B(n5649), .Z(c[781]) );
  XOR U6921 ( .A(n5652), .B(n5651), .Z(c[782]) );
  XOR U6922 ( .A(n5654), .B(n5653), .Z(c[783]) );
  XOR U6923 ( .A(n5656), .B(n5655), .Z(c[784]) );
  XOR U6924 ( .A(n5658), .B(n5657), .Z(c[785]) );
  XOR U6925 ( .A(n5660), .B(n5659), .Z(c[786]) );
  XOR U6926 ( .A(n5662), .B(n5661), .Z(c[787]) );
  XOR U6927 ( .A(n5664), .B(n5663), .Z(c[788]) );
  XOR U6928 ( .A(n5666), .B(n5665), .Z(c[789]) );
  XOR U6929 ( .A(n5668), .B(n5667), .Z(c[78]) );
  XOR U6930 ( .A(n5670), .B(n5669), .Z(c[790]) );
  XOR U6931 ( .A(n5672), .B(n5671), .Z(c[791]) );
  XOR U6932 ( .A(n5674), .B(n5673), .Z(c[792]) );
  XOR U6933 ( .A(n5676), .B(n5675), .Z(c[793]) );
  XOR U6934 ( .A(n5678), .B(n5677), .Z(c[794]) );
  XOR U6935 ( .A(n5680), .B(n5679), .Z(c[795]) );
  XOR U6936 ( .A(n5682), .B(n5681), .Z(c[796]) );
  XOR U6937 ( .A(n5684), .B(n5683), .Z(c[797]) );
  XOR U6938 ( .A(n5686), .B(n5685), .Z(c[798]) );
  XOR U6939 ( .A(n5688), .B(n5687), .Z(c[799]) );
  XOR U6940 ( .A(n5690), .B(n5689), .Z(c[79]) );
  XOR U6941 ( .A(n5692), .B(n5691), .Z(c[7]) );
  XOR U6942 ( .A(n5694), .B(n5693), .Z(c[800]) );
  XOR U6943 ( .A(n5696), .B(n5695), .Z(c[801]) );
  XOR U6944 ( .A(n5698), .B(n5697), .Z(c[802]) );
  XOR U6945 ( .A(n5700), .B(n5699), .Z(c[803]) );
  XOR U6946 ( .A(n5702), .B(n5701), .Z(c[804]) );
  XOR U6947 ( .A(n5704), .B(n5703), .Z(c[805]) );
  XOR U6948 ( .A(n5706), .B(n5705), .Z(c[806]) );
  XOR U6949 ( .A(n5708), .B(n5707), .Z(c[807]) );
  XOR U6950 ( .A(n5710), .B(n5709), .Z(c[808]) );
  XOR U6951 ( .A(n5712), .B(n5711), .Z(c[809]) );
  XOR U6952 ( .A(n5714), .B(n5713), .Z(c[80]) );
  XOR U6953 ( .A(n5716), .B(n5715), .Z(c[810]) );
  XOR U6954 ( .A(n5718), .B(n5717), .Z(c[811]) );
  XOR U6955 ( .A(n5720), .B(n5719), .Z(c[812]) );
  XOR U6956 ( .A(n5722), .B(n5721), .Z(c[813]) );
  XOR U6957 ( .A(n5724), .B(n5723), .Z(c[814]) );
  XOR U6958 ( .A(n5726), .B(n5725), .Z(c[815]) );
  XOR U6959 ( .A(n5728), .B(n5727), .Z(c[816]) );
  XOR U6960 ( .A(n5730), .B(n5729), .Z(c[817]) );
  XOR U6961 ( .A(n5732), .B(n5731), .Z(c[818]) );
  XOR U6962 ( .A(n5734), .B(n5733), .Z(c[819]) );
  XOR U6963 ( .A(n5736), .B(n5735), .Z(c[81]) );
  XOR U6964 ( .A(n5738), .B(n5737), .Z(c[820]) );
  XOR U6965 ( .A(n5740), .B(n5739), .Z(c[821]) );
  XOR U6966 ( .A(n5742), .B(n5741), .Z(c[822]) );
  XOR U6967 ( .A(n5744), .B(n5743), .Z(c[823]) );
  XOR U6968 ( .A(n5746), .B(n5745), .Z(c[824]) );
  XOR U6969 ( .A(n5748), .B(n5747), .Z(c[825]) );
  XOR U6970 ( .A(n5750), .B(n5749), .Z(c[826]) );
  XOR U6971 ( .A(n5752), .B(n5751), .Z(c[827]) );
  XOR U6972 ( .A(n5754), .B(n5753), .Z(c[828]) );
  XOR U6973 ( .A(n5756), .B(n5755), .Z(c[829]) );
  XOR U6974 ( .A(n5758), .B(n5757), .Z(c[82]) );
  XOR U6975 ( .A(n5760), .B(n5759), .Z(c[830]) );
  XOR U6976 ( .A(n5762), .B(n5761), .Z(c[831]) );
  XOR U6977 ( .A(n5764), .B(n5763), .Z(c[832]) );
  XOR U6978 ( .A(n5766), .B(n5765), .Z(c[833]) );
  XOR U6979 ( .A(n5768), .B(n5767), .Z(c[834]) );
  XOR U6980 ( .A(n5770), .B(n5769), .Z(c[835]) );
  XOR U6981 ( .A(n5772), .B(n5771), .Z(c[836]) );
  XOR U6982 ( .A(n5774), .B(n5773), .Z(c[837]) );
  XOR U6983 ( .A(n5776), .B(n5775), .Z(c[838]) );
  XOR U6984 ( .A(n5778), .B(n5777), .Z(c[839]) );
  XOR U6985 ( .A(n5780), .B(n5779), .Z(c[83]) );
  XOR U6986 ( .A(n5782), .B(n5781), .Z(c[840]) );
  XOR U6987 ( .A(n5784), .B(n5783), .Z(c[841]) );
  XOR U6988 ( .A(n5786), .B(n5785), .Z(c[842]) );
  XOR U6989 ( .A(n5788), .B(n5787), .Z(c[843]) );
  XOR U6990 ( .A(n5790), .B(n5789), .Z(c[844]) );
  XOR U6991 ( .A(n5792), .B(n5791), .Z(c[845]) );
  XOR U6992 ( .A(n5794), .B(n5793), .Z(c[846]) );
  XOR U6993 ( .A(n5796), .B(n5795), .Z(c[847]) );
  XOR U6994 ( .A(n5798), .B(n5797), .Z(c[848]) );
  XOR U6995 ( .A(n5800), .B(n5799), .Z(c[849]) );
  XOR U6996 ( .A(n5802), .B(n5801), .Z(c[84]) );
  XOR U6997 ( .A(n5804), .B(n5803), .Z(c[850]) );
  XOR U6998 ( .A(n5806), .B(n5805), .Z(c[851]) );
  XOR U6999 ( .A(n5808), .B(n5807), .Z(c[852]) );
  XOR U7000 ( .A(n5810), .B(n5809), .Z(c[853]) );
  XOR U7001 ( .A(n5812), .B(n5811), .Z(c[854]) );
  XOR U7002 ( .A(n5814), .B(n5813), .Z(c[855]) );
  XOR U7003 ( .A(n5816), .B(n5815), .Z(c[856]) );
  XOR U7004 ( .A(n5818), .B(n5817), .Z(c[857]) );
  XOR U7005 ( .A(n5820), .B(n5819), .Z(c[858]) );
  XOR U7006 ( .A(n5822), .B(n5821), .Z(c[859]) );
  XOR U7007 ( .A(n5824), .B(n5823), .Z(c[85]) );
  XOR U7008 ( .A(n5826), .B(n5825), .Z(c[860]) );
  XOR U7009 ( .A(n5828), .B(n5827), .Z(c[861]) );
  XOR U7010 ( .A(n5830), .B(n5829), .Z(c[862]) );
  XOR U7011 ( .A(n5832), .B(n5831), .Z(c[863]) );
  XOR U7012 ( .A(n5834), .B(n5833), .Z(c[864]) );
  XOR U7013 ( .A(n5836), .B(n5835), .Z(c[865]) );
  XOR U7014 ( .A(n5838), .B(n5837), .Z(c[866]) );
  XOR U7015 ( .A(n5840), .B(n5839), .Z(c[867]) );
  XOR U7016 ( .A(n5842), .B(n5841), .Z(c[868]) );
  XOR U7017 ( .A(n5844), .B(n5843), .Z(c[869]) );
  XOR U7018 ( .A(n5846), .B(n5845), .Z(c[86]) );
  XOR U7019 ( .A(n5848), .B(n5847), .Z(c[870]) );
  XOR U7020 ( .A(n5850), .B(n5849), .Z(c[871]) );
  XOR U7021 ( .A(n5852), .B(n5851), .Z(c[872]) );
  XOR U7022 ( .A(n5854), .B(n5853), .Z(c[873]) );
  XOR U7023 ( .A(n5856), .B(n5855), .Z(c[874]) );
  XOR U7024 ( .A(n5858), .B(n5857), .Z(c[875]) );
  XOR U7025 ( .A(n5860), .B(n5859), .Z(c[876]) );
  XOR U7026 ( .A(n5862), .B(n5861), .Z(c[877]) );
  XOR U7027 ( .A(n5864), .B(n5863), .Z(c[878]) );
  XOR U7028 ( .A(n5866), .B(n5865), .Z(c[879]) );
  XOR U7029 ( .A(n5868), .B(n5867), .Z(c[87]) );
  XOR U7030 ( .A(n5870), .B(n5869), .Z(c[880]) );
  XOR U7031 ( .A(n5872), .B(n5871), .Z(c[881]) );
  XOR U7032 ( .A(n5874), .B(n5873), .Z(c[882]) );
  XOR U7033 ( .A(n5876), .B(n5875), .Z(c[883]) );
  XOR U7034 ( .A(n5878), .B(n5877), .Z(c[884]) );
  XOR U7035 ( .A(n5880), .B(n5879), .Z(c[885]) );
  XOR U7036 ( .A(n5882), .B(n5881), .Z(c[886]) );
  XOR U7037 ( .A(n5884), .B(n5883), .Z(c[887]) );
  XOR U7038 ( .A(n5886), .B(n5885), .Z(c[888]) );
  XOR U7039 ( .A(n5888), .B(n5887), .Z(c[889]) );
  XOR U7040 ( .A(n5890), .B(n5889), .Z(c[88]) );
  XOR U7041 ( .A(n5892), .B(n5891), .Z(c[890]) );
  XOR U7042 ( .A(n5894), .B(n5893), .Z(c[891]) );
  XOR U7043 ( .A(n5896), .B(n5895), .Z(c[892]) );
  XOR U7044 ( .A(n5898), .B(n5897), .Z(c[893]) );
  XOR U7045 ( .A(n5900), .B(n5899), .Z(c[894]) );
  XOR U7046 ( .A(n5902), .B(n5901), .Z(c[895]) );
  XOR U7047 ( .A(n5904), .B(n5903), .Z(c[896]) );
  XOR U7048 ( .A(n5906), .B(n5905), .Z(c[897]) );
  XOR U7049 ( .A(n5908), .B(n5907), .Z(c[898]) );
  XOR U7050 ( .A(n5910), .B(n5909), .Z(c[899]) );
  XOR U7051 ( .A(n5912), .B(n5911), .Z(c[89]) );
  XOR U7052 ( .A(n5914), .B(n5913), .Z(c[8]) );
  XOR U7053 ( .A(n5916), .B(n5915), .Z(c[900]) );
  XOR U7054 ( .A(n5918), .B(n5917), .Z(c[901]) );
  XOR U7055 ( .A(n5920), .B(n5919), .Z(c[902]) );
  XOR U7056 ( .A(n5922), .B(n5921), .Z(c[903]) );
  XOR U7057 ( .A(n5924), .B(n5923), .Z(c[904]) );
  XOR U7058 ( .A(n5926), .B(n5925), .Z(c[905]) );
  XOR U7059 ( .A(n5928), .B(n5927), .Z(c[906]) );
  XOR U7060 ( .A(n5930), .B(n5929), .Z(c[907]) );
  XOR U7061 ( .A(n5932), .B(n5931), .Z(c[908]) );
  XOR U7062 ( .A(n5934), .B(n5933), .Z(c[909]) );
  XOR U7063 ( .A(n5936), .B(n5935), .Z(c[90]) );
  XOR U7064 ( .A(n5938), .B(n5937), .Z(c[910]) );
  XOR U7065 ( .A(n5940), .B(n5939), .Z(c[911]) );
  XOR U7066 ( .A(n5942), .B(n5941), .Z(c[912]) );
  XOR U7067 ( .A(n5944), .B(n5943), .Z(c[913]) );
  XOR U7068 ( .A(n5946), .B(n5945), .Z(c[914]) );
  XOR U7069 ( .A(n5948), .B(n5947), .Z(c[915]) );
  XOR U7070 ( .A(n5950), .B(n5949), .Z(c[916]) );
  XOR U7071 ( .A(n5952), .B(n5951), .Z(c[917]) );
  XOR U7072 ( .A(n5954), .B(n5953), .Z(c[918]) );
  XOR U7073 ( .A(n5956), .B(n5955), .Z(c[919]) );
  XOR U7074 ( .A(n5958), .B(n5957), .Z(c[91]) );
  XOR U7075 ( .A(n5960), .B(n5959), .Z(c[920]) );
  XOR U7076 ( .A(n5962), .B(n5961), .Z(c[921]) );
  XOR U7077 ( .A(n5964), .B(n5963), .Z(c[922]) );
  XOR U7078 ( .A(n5966), .B(n5965), .Z(c[923]) );
  XOR U7079 ( .A(n5968), .B(n5967), .Z(c[924]) );
  XOR U7080 ( .A(n5970), .B(n5969), .Z(c[925]) );
  XOR U7081 ( .A(n5972), .B(n5971), .Z(c[926]) );
  XOR U7082 ( .A(n5974), .B(n5973), .Z(c[927]) );
  XOR U7083 ( .A(n5976), .B(n5975), .Z(c[928]) );
  XOR U7084 ( .A(n5978), .B(n5977), .Z(c[929]) );
  XOR U7085 ( .A(n5980), .B(n5979), .Z(c[92]) );
  XOR U7086 ( .A(n5982), .B(n5981), .Z(c[930]) );
  XOR U7087 ( .A(n5984), .B(n5983), .Z(c[931]) );
  XOR U7088 ( .A(n5986), .B(n5985), .Z(c[932]) );
  XOR U7089 ( .A(n5988), .B(n5987), .Z(c[933]) );
  XOR U7090 ( .A(n5990), .B(n5989), .Z(c[934]) );
  XOR U7091 ( .A(n5992), .B(n5991), .Z(c[935]) );
  XOR U7092 ( .A(n5994), .B(n5993), .Z(c[936]) );
  XOR U7093 ( .A(n5996), .B(n5995), .Z(c[937]) );
  XOR U7094 ( .A(n5998), .B(n5997), .Z(c[938]) );
  XOR U7095 ( .A(n6000), .B(n5999), .Z(c[939]) );
  XOR U7096 ( .A(n6002), .B(n6001), .Z(c[93]) );
  XOR U7097 ( .A(n6004), .B(n6003), .Z(c[940]) );
  XOR U7098 ( .A(n6006), .B(n6005), .Z(c[941]) );
  XOR U7099 ( .A(n6008), .B(n6007), .Z(c[942]) );
  XOR U7100 ( .A(n6010), .B(n6009), .Z(c[943]) );
  XOR U7101 ( .A(n6012), .B(n6011), .Z(c[944]) );
  XOR U7102 ( .A(n6014), .B(n6013), .Z(c[945]) );
  XOR U7103 ( .A(n6016), .B(n6015), .Z(c[946]) );
  XOR U7104 ( .A(n6018), .B(n6017), .Z(c[947]) );
  XOR U7105 ( .A(n6020), .B(n6019), .Z(c[948]) );
  XOR U7106 ( .A(n6022), .B(n6021), .Z(c[949]) );
  XOR U7107 ( .A(n6024), .B(n6023), .Z(c[94]) );
  XOR U7108 ( .A(n6026), .B(n6025), .Z(c[950]) );
  XOR U7109 ( .A(n6028), .B(n6027), .Z(c[951]) );
  XOR U7110 ( .A(n6030), .B(n6029), .Z(c[952]) );
  XOR U7111 ( .A(n6032), .B(n6031), .Z(c[953]) );
  XOR U7112 ( .A(n6034), .B(n6033), .Z(c[954]) );
  XOR U7113 ( .A(n6036), .B(n6035), .Z(c[955]) );
  XOR U7114 ( .A(n6038), .B(n6037), .Z(c[956]) );
  XOR U7115 ( .A(n6040), .B(n6039), .Z(c[957]) );
  XOR U7116 ( .A(n6042), .B(n6041), .Z(c[958]) );
  XOR U7117 ( .A(n6044), .B(n6043), .Z(c[959]) );
  XOR U7118 ( .A(n6046), .B(n6045), .Z(c[95]) );
  XOR U7119 ( .A(n6048), .B(n6047), .Z(c[960]) );
  XOR U7120 ( .A(n6050), .B(n6049), .Z(c[961]) );
  XOR U7121 ( .A(n6052), .B(n6051), .Z(c[962]) );
  XOR U7122 ( .A(n6054), .B(n6053), .Z(c[963]) );
  XOR U7123 ( .A(n6056), .B(n6055), .Z(c[964]) );
  XOR U7124 ( .A(n6058), .B(n6057), .Z(c[965]) );
  XOR U7125 ( .A(n6060), .B(n6059), .Z(c[966]) );
  XOR U7126 ( .A(n6062), .B(n6061), .Z(c[967]) );
  XOR U7127 ( .A(n6064), .B(n6063), .Z(c[968]) );
  XOR U7128 ( .A(n6066), .B(n6065), .Z(c[969]) );
  XOR U7129 ( .A(n6068), .B(n6067), .Z(c[96]) );
  XOR U7130 ( .A(n6070), .B(n6069), .Z(c[970]) );
  XOR U7131 ( .A(n6072), .B(n6071), .Z(c[971]) );
  XOR U7132 ( .A(n6074), .B(n6073), .Z(c[972]) );
  XOR U7133 ( .A(n6076), .B(n6075), .Z(c[973]) );
  XOR U7134 ( .A(n6078), .B(n6077), .Z(c[974]) );
  XOR U7135 ( .A(n6080), .B(n6079), .Z(c[975]) );
  XOR U7136 ( .A(n6082), .B(n6081), .Z(c[976]) );
  XOR U7137 ( .A(n6084), .B(n6083), .Z(c[977]) );
  XOR U7138 ( .A(n6086), .B(n6085), .Z(c[978]) );
  XOR U7139 ( .A(n6088), .B(n6087), .Z(c[979]) );
  XOR U7140 ( .A(n6090), .B(n6089), .Z(c[97]) );
  XOR U7141 ( .A(n6092), .B(n6091), .Z(c[980]) );
  XOR U7142 ( .A(n6094), .B(n6093), .Z(c[981]) );
  XOR U7143 ( .A(n6096), .B(n6095), .Z(c[982]) );
  XOR U7144 ( .A(n6098), .B(n6097), .Z(c[983]) );
  XOR U7145 ( .A(n6100), .B(n6099), .Z(c[984]) );
  XOR U7146 ( .A(n6102), .B(n6101), .Z(c[985]) );
  XOR U7147 ( .A(n6104), .B(n6103), .Z(c[986]) );
  XOR U7148 ( .A(n6106), .B(n6105), .Z(c[987]) );
  XOR U7149 ( .A(n6108), .B(n6107), .Z(c[988]) );
  XOR U7150 ( .A(n6110), .B(n6109), .Z(c[989]) );
  XOR U7151 ( .A(n6112), .B(n6111), .Z(c[98]) );
  XOR U7152 ( .A(n6114), .B(n6113), .Z(c[990]) );
  XOR U7153 ( .A(n6116), .B(n6115), .Z(c[991]) );
  XOR U7154 ( .A(n6118), .B(n6117), .Z(c[992]) );
  XOR U7155 ( .A(n6120), .B(n6119), .Z(c[993]) );
  XOR U7156 ( .A(n6122), .B(n6121), .Z(c[994]) );
  XOR U7157 ( .A(n6124), .B(n6123), .Z(c[995]) );
  XOR U7158 ( .A(n6126), .B(n6125), .Z(c[996]) );
  XOR U7159 ( .A(n6128), .B(n6127), .Z(c[997]) );
  XOR U7160 ( .A(n6130), .B(n6129), .Z(c[998]) );
  XOR U7161 ( .A(n6132), .B(n6131), .Z(c[999]) );
  XOR U7162 ( .A(n6134), .B(n6133), .Z(c[99]) );
  XOR U7163 ( .A(n6136), .B(n6135), .Z(c[9]) );
  NOR U7164 ( .A(n6138), .B(n6137), .Z(n6142) );
  IV U7165 ( .A(a[1023]), .Z(n6139) );
  NOR U7166 ( .A(n6140), .B(n6139), .Z(n6141) );
  NOR U7167 ( .A(n6142), .B(n6141), .Z(n6143) );
  IV U7168 ( .A(n6143), .Z(c[1024]) );
endmodule

