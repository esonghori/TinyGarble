
module compare_N16384_CC4 ( clk, rst, x, y, g, e );
  input [4095:0] x;
  input [4095:0] y;
  input clk, rst;
  output g, e;
  wire   ebreg, n4, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626,
         n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
         n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
         n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,
         n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
         n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666,
         n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674,
         n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
         n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
         n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706,
         n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
         n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,
         n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
         n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,
         n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746,
         n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
         n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,
         n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770,
         n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778,
         n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786,
         n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794,
         n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802,
         n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810,
         n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818,
         n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826,
         n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834,
         n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842,
         n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850,
         n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858,
         n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866,
         n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874,
         n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882,
         n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890,
         n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898,
         n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906,
         n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914,
         n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922,
         n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930,
         n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938,
         n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946,
         n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954,
         n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962,
         n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970,
         n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978,
         n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986,
         n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994,
         n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002,
         n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010,
         n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
         n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,
         n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034,
         n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,
         n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050,
         n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058,
         n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066,
         n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
         n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082,
         n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,
         n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,
         n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106,
         n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114,
         n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122,
         n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130,
         n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
         n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146,
         n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154,
         n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,
         n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170,
         n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178,
         n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186,
         n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194,
         n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202,
         n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
         n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218,
         n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226,
         n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
         n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242,
         n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250,
         n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258,
         n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266,
         n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274,
         n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282,
         n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290,
         n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298,
         n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
         n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314,
         n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322,
         n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330,
         n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
         n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346,
         n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354,
         n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,
         n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370,
         n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
         n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386,
         n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394,
         n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402,
         n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
         n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,
         n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,
         n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,
         n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442,
         n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
         n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458,
         n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466,
         n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,
         n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
         n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490,
         n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
         n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
         n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
         n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
         n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538,
         n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546,
         n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
         n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562,
         n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,
         n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
         n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,
         n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
         n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602,
         n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610,
         n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618,
         n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626,
         n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634,
         n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642,
         n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650,
         n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658,
         n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
         n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674,
         n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682,
         n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690,
         n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
         n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706,
         n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714,
         n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722,
         n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730,
         n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,
         n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746,
         n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754,
         n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762,
         n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770,
         n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778,
         n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786,
         n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794,
         n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802,
         n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,
         n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818,
         n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826,
         n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834,
         n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842,
         n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850,
         n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858,
         n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866,
         n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874,
         n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,
         n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890,
         n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898,
         n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906,
         n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914,
         n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922,
         n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930,
         n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938,
         n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946,
         n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,
         n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962,
         n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970,
         n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978,
         n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986,
         n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994,
         n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002,
         n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010,
         n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018,
         n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
         n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034,
         n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042,
         n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050,
         n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058,
         n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
         n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074,
         n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082,
         n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090,
         n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
         n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106,
         n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114,
         n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122,
         n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130,
         n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,
         n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,
         n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
         n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
         n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
         n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178,
         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,
         n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194,
         n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,
         n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,
         n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218,
         n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
         n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234,
         n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
         n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250,
         n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258,
         n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266,
         n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
         n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282,
         n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290,
         n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
         n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306,
         n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314,
         n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322,
         n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330,
         n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338,
         n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346,
         n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
         n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362,
         n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,
         n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378,
         n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386,
         n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394,
         n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402,
         n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410,
         n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418,
         n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426,
         n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434,
         n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,
         n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450,
         n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458,
         n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466,
         n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474,
         n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482,
         n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490,
         n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498,
         n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506,
         n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514,
         n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522,
         n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530,
         n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538,
         n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546,
         n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554,
         n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562,
         n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570,
         n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578,
         n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586,
         n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594,
         n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602,
         n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610,
         n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618,
         n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626,
         n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634,
         n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642,
         n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650,
         n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658,
         n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666,
         n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674,
         n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682,
         n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690,
         n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698,
         n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706,
         n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714,
         n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722,
         n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730,
         n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738,
         n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746,
         n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754,
         n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762,
         n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770,
         n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778,
         n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786,
         n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794,
         n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802,
         n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810,
         n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818,
         n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826,
         n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834,
         n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842,
         n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850,
         n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858,
         n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866,
         n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874,
         n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882,
         n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890,
         n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898,
         n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906,
         n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914,
         n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922,
         n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930,
         n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938,
         n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946,
         n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954,
         n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962,
         n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970,
         n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978,
         n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986,
         n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994,
         n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002,
         n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010,
         n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018,
         n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026,
         n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034,
         n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042,
         n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050,
         n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058,
         n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066,
         n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074,
         n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082,
         n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090,
         n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098,
         n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106,
         n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114,
         n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122,
         n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130,
         n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138,
         n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146,
         n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154,
         n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162,
         n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170,
         n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178,
         n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186,
         n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194,
         n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202,
         n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210,
         n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218,
         n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226,
         n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234,
         n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242,
         n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250,
         n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258,
         n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266,
         n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274,
         n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282,
         n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290,
         n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298,
         n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306,
         n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314,
         n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322,
         n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330,
         n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338,
         n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346,
         n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354,
         n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362,
         n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370,
         n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378,
         n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386,
         n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394,
         n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402,
         n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410,
         n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418,
         n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426,
         n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434,
         n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442,
         n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450,
         n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458,
         n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466,
         n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474,
         n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482,
         n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490,
         n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498,
         n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506,
         n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514,
         n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522,
         n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530,
         n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538,
         n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546,
         n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554,
         n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562,
         n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570,
         n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578,
         n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586,
         n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594,
         n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602,
         n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610,
         n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618,
         n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626,
         n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634,
         n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642,
         n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650,
         n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658,
         n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666,
         n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674,
         n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682,
         n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690,
         n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698,
         n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706,
         n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714,
         n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722,
         n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730,
         n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738,
         n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746,
         n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754,
         n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762,
         n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770,
         n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778,
         n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786,
         n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794,
         n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802,
         n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810,
         n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818,
         n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826,
         n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834,
         n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842,
         n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850,
         n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858,
         n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866,
         n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874,
         n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882,
         n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890,
         n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898,
         n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906,
         n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914,
         n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922,
         n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930,
         n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938,
         n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946,
         n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954,
         n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962,
         n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970,
         n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978,
         n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986,
         n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994,
         n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002,
         n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010,
         n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018,
         n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026,
         n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034,
         n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042,
         n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050,
         n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058,
         n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066,
         n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074,
         n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082,
         n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090,
         n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098,
         n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106,
         n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114,
         n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122,
         n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130,
         n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138,
         n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146,
         n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154,
         n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162,
         n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170,
         n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178,
         n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186,
         n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194,
         n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202,
         n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210,
         n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218,
         n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226,
         n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234,
         n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242,
         n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250,
         n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258,
         n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266,
         n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274,
         n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282,
         n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290,
         n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298,
         n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306,
         n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314,
         n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322,
         n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330,
         n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338,
         n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346,
         n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354,
         n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362,
         n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370,
         n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378,
         n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386,
         n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394,
         n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402,
         n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410,
         n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418,
         n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426,
         n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434,
         n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442,
         n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450,
         n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458,
         n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466,
         n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474,
         n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482,
         n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490,
         n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498,
         n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506,
         n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514,
         n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522,
         n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530,
         n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538,
         n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546,
         n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554,
         n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562,
         n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570,
         n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578,
         n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586,
         n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594,
         n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602,
         n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610,
         n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618,
         n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626,
         n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634,
         n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642,
         n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650,
         n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658,
         n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666,
         n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674,
         n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682,
         n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690,
         n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698,
         n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706,
         n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714,
         n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
         n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730,
         n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738,
         n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746,
         n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754,
         n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762,
         n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770,
         n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778,
         n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786,
         n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794,
         n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802,
         n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810,
         n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818,
         n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826,
         n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834,
         n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842,
         n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850,
         n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858,
         n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866,
         n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874,
         n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882,
         n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890,
         n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898,
         n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906,
         n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914,
         n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922,
         n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930,
         n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
         n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946,
         n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954,
         n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962,
         n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970,
         n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978,
         n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986,
         n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994,
         n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002,
         n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010,
         n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018,
         n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026,
         n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034,
         n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042,
         n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050,
         n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058,
         n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066,
         n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074,
         n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082,
         n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090,
         n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098,
         n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106,
         n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114,
         n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122,
         n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130,
         n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138,
         n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146,
         n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154,
         n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162,
         n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170,
         n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178,
         n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186,
         n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194,
         n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202,
         n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210,
         n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218,
         n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226,
         n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234,
         n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242,
         n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250,
         n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258,
         n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266,
         n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274,
         n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282,
         n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290,
         n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298,
         n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306,
         n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314,
         n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322,
         n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330,
         n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338,
         n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346,
         n21347, n21348, n21349, n21350, n21351, n21352, n21353, n21354,
         n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362,
         n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370,
         n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378,
         n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386,
         n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394,
         n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402,
         n21403, n21404, n21405, n21406, n21407, n21408, n21409, n21410,
         n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418,
         n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426,
         n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434,
         n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442,
         n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450,
         n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458,
         n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466,
         n21467, n21468, n21469, n21470, n21471, n21472, n21473, n21474,
         n21475, n21476, n21477, n21478, n21479, n21480, n21481, n21482,
         n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490,
         n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498,
         n21499, n21500, n21501, n21502, n21503, n21504, n21505, n21506,
         n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514,
         n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522,
         n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530,
         n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538,
         n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546,
         n21547, n21548, n21549, n21550, n21551, n21552, n21553, n21554,
         n21555, n21556, n21557, n21558, n21559, n21560, n21561, n21562,
         n21563, n21564, n21565, n21566, n21567, n21568, n21569, n21570,
         n21571, n21572, n21573, n21574, n21575, n21576, n21577, n21578,
         n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586,
         n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594,
         n21595, n21596, n21597, n21598, n21599, n21600, n21601, n21602,
         n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610,
         n21611, n21612, n21613, n21614, n21615, n21616, n21617, n21618,
         n21619, n21620, n21621, n21622, n21623, n21624, n21625, n21626,
         n21627, n21628, n21629, n21630, n21631, n21632, n21633, n21634,
         n21635, n21636, n21637, n21638, n21639, n21640, n21641, n21642,
         n21643, n21644, n21645, n21646, n21647, n21648, n21649, n21650,
         n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658,
         n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666,
         n21667, n21668, n21669, n21670, n21671, n21672, n21673, n21674,
         n21675, n21676, n21677, n21678, n21679, n21680, n21681, n21682,
         n21683, n21684, n21685, n21686, n21687, n21688, n21689, n21690,
         n21691, n21692, n21693, n21694, n21695, n21696, n21697, n21698,
         n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706,
         n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21714,
         n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722,
         n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730,
         n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738,
         n21739, n21740, n21741, n21742, n21743, n21744, n21745, n21746,
         n21747, n21748, n21749, n21750, n21751, n21752, n21753, n21754,
         n21755, n21756, n21757, n21758, n21759, n21760, n21761, n21762,
         n21763, n21764, n21765, n21766, n21767, n21768, n21769, n21770,
         n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778,
         n21779, n21780, n21781, n21782, n21783, n21784, n21785, n21786,
         n21787, n21788, n21789, n21790, n21791, n21792, n21793, n21794,
         n21795, n21796, n21797, n21798, n21799, n21800, n21801, n21802,
         n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810,
         n21811, n21812, n21813, n21814, n21815, n21816, n21817, n21818,
         n21819, n21820, n21821, n21822, n21823, n21824, n21825, n21826,
         n21827, n21828, n21829, n21830, n21831, n21832, n21833, n21834,
         n21835, n21836, n21837, n21838, n21839, n21840, n21841, n21842,
         n21843, n21844, n21845, n21846, n21847, n21848, n21849, n21850,
         n21851, n21852, n21853, n21854, n21855, n21856, n21857, n21858,
         n21859, n21860, n21861, n21862, n21863, n21864, n21865, n21866,
         n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21874,
         n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882,
         n21883, n21884, n21885, n21886, n21887, n21888, n21889, n21890,
         n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21898,
         n21899, n21900, n21901, n21902, n21903, n21904, n21905, n21906,
         n21907, n21908, n21909, n21910, n21911, n21912, n21913, n21914,
         n21915, n21916, n21917, n21918, n21919, n21920, n21921, n21922,
         n21923, n21924, n21925, n21926, n21927, n21928, n21929, n21930,
         n21931, n21932, n21933, n21934, n21935, n21936, n21937, n21938,
         n21939, n21940, n21941, n21942, n21943, n21944, n21945, n21946,
         n21947, n21948, n21949, n21950, n21951, n21952, n21953, n21954,
         n21955, n21956, n21957, n21958, n21959, n21960, n21961, n21962,
         n21963, n21964, n21965, n21966, n21967, n21968, n21969, n21970,
         n21971, n21972, n21973, n21974, n21975, n21976, n21977, n21978,
         n21979, n21980, n21981, n21982, n21983, n21984, n21985, n21986,
         n21987, n21988, n21989, n21990, n21991, n21992, n21993, n21994,
         n21995, n21996, n21997, n21998, n21999, n22000, n22001, n22002,
         n22003, n22004, n22005, n22006, n22007, n22008, n22009, n22010,
         n22011, n22012, n22013, n22014, n22015, n22016, n22017, n22018,
         n22019, n22020, n22021, n22022, n22023, n22024, n22025, n22026,
         n22027, n22028, n22029, n22030, n22031, n22032, n22033, n22034,
         n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042,
         n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050,
         n22051, n22052, n22053, n22054, n22055, n22056, n22057, n22058,
         n22059, n22060, n22061, n22062, n22063, n22064, n22065, n22066,
         n22067, n22068, n22069, n22070, n22071, n22072, n22073, n22074,
         n22075, n22076, n22077, n22078, n22079, n22080, n22081, n22082,
         n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090,
         n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098,
         n22099, n22100, n22101, n22102, n22103, n22104, n22105, n22106,
         n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114,
         n22115, n22116, n22117, n22118, n22119, n22120, n22121, n22122,
         n22123, n22124, n22125, n22126, n22127, n22128, n22129, n22130,
         n22131, n22132, n22133, n22134, n22135, n22136, n22137, n22138,
         n22139, n22140, n22141, n22142, n22143, n22144, n22145, n22146,
         n22147, n22148, n22149, n22150, n22151, n22152, n22153, n22154,
         n22155, n22156, n22157, n22158, n22159, n22160, n22161, n22162,
         n22163, n22164, n22165, n22166, n22167, n22168, n22169, n22170,
         n22171, n22172, n22173, n22174, n22175, n22176, n22177, n22178,
         n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22186,
         n22187, n22188, n22189, n22190, n22191, n22192, n22193, n22194,
         n22195, n22196, n22197, n22198, n22199, n22200, n22201, n22202,
         n22203, n22204, n22205, n22206, n22207, n22208, n22209, n22210,
         n22211, n22212, n22213, n22214, n22215, n22216, n22217, n22218,
         n22219, n22220, n22221, n22222, n22223, n22224, n22225, n22226,
         n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22234,
         n22235, n22236, n22237, n22238, n22239, n22240, n22241, n22242,
         n22243, n22244, n22245, n22246, n22247, n22248, n22249, n22250,
         n22251, n22252, n22253, n22254, n22255, n22256, n22257, n22258,
         n22259, n22260, n22261, n22262, n22263, n22264, n22265, n22266,
         n22267, n22268, n22269, n22270, n22271, n22272, n22273, n22274,
         n22275, n22276, n22277, n22278, n22279, n22280, n22281, n22282,
         n22283, n22284, n22285, n22286, n22287, n22288, n22289, n22290,
         n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298,
         n22299, n22300, n22301, n22302, n22303, n22304, n22305, n22306,
         n22307, n22308, n22309, n22310, n22311, n22312, n22313, n22314,
         n22315, n22316, n22317, n22318, n22319, n22320, n22321, n22322,
         n22323, n22324, n22325, n22326, n22327, n22328, n22329, n22330,
         n22331, n22332, n22333, n22334, n22335, n22336, n22337, n22338,
         n22339, n22340, n22341, n22342, n22343, n22344, n22345, n22346,
         n22347, n22348, n22349, n22350, n22351, n22352, n22353, n22354,
         n22355, n22356, n22357, n22358, n22359, n22360, n22361, n22362,
         n22363, n22364, n22365, n22366, n22367, n22368, n22369, n22370,
         n22371, n22372, n22373, n22374, n22375, n22376, n22377, n22378,
         n22379, n22380, n22381, n22382, n22383, n22384, n22385, n22386,
         n22387, n22388, n22389, n22390, n22391, n22392, n22393, n22394,
         n22395, n22396, n22397, n22398, n22399, n22400, n22401, n22402,
         n22403, n22404, n22405, n22406, n22407, n22408, n22409, n22410,
         n22411, n22412, n22413, n22414, n22415, n22416, n22417, n22418,
         n22419, n22420, n22421, n22422, n22423, n22424, n22425, n22426,
         n22427, n22428, n22429, n22430, n22431, n22432, n22433, n22434,
         n22435, n22436, n22437, n22438, n22439, n22440, n22441, n22442,
         n22443, n22444, n22445, n22446, n22447, n22448, n22449, n22450,
         n22451, n22452, n22453, n22454, n22455, n22456, n22457, n22458,
         n22459, n22460, n22461, n22462, n22463, n22464, n22465, n22466,
         n22467, n22468, n22469, n22470, n22471, n22472, n22473, n22474,
         n22475, n22476, n22477, n22478, n22479, n22480, n22481, n22482,
         n22483, n22484, n22485, n22486, n22487, n22488, n22489, n22490,
         n22491, n22492, n22493, n22494, n22495, n22496, n22497, n22498,
         n22499, n22500, n22501, n22502, n22503, n22504, n22505, n22506,
         n22507, n22508, n22509, n22510, n22511, n22512, n22513, n22514,
         n22515, n22516, n22517, n22518, n22519, n22520, n22521, n22522,
         n22523, n22524, n22525, n22526, n22527, n22528, n22529, n22530,
         n22531, n22532, n22533, n22534, n22535, n22536, n22537, n22538,
         n22539, n22540, n22541, n22542, n22543, n22544, n22545, n22546,
         n22547, n22548, n22549, n22550, n22551, n22552, n22553, n22554,
         n22555, n22556, n22557, n22558, n22559, n22560, n22561, n22562,
         n22563, n22564, n22565, n22566, n22567, n22568, n22569, n22570,
         n22571, n22572, n22573, n22574, n22575, n22576, n22577, n22578,
         n22579, n22580, n22581, n22582, n22583, n22584, n22585, n22586,
         n22587, n22588, n22589, n22590, n22591, n22592, n22593, n22594,
         n22595, n22596, n22597, n22598, n22599, n22600, n22601, n22602,
         n22603, n22604, n22605, n22606, n22607, n22608, n22609, n22610,
         n22611, n22612, n22613, n22614, n22615, n22616, n22617, n22618,
         n22619, n22620, n22621, n22622, n22623, n22624, n22625, n22626,
         n22627, n22628, n22629, n22630, n22631, n22632, n22633, n22634,
         n22635, n22636, n22637, n22638, n22639, n22640, n22641, n22642,
         n22643, n22644, n22645, n22646, n22647, n22648, n22649, n22650,
         n22651, n22652, n22653, n22654, n22655, n22656, n22657, n22658,
         n22659, n22660, n22661, n22662, n22663, n22664, n22665, n22666,
         n22667, n22668, n22669, n22670, n22671, n22672, n22673, n22674,
         n22675, n22676, n22677, n22678, n22679, n22680, n22681, n22682,
         n22683, n22684, n22685, n22686, n22687, n22688, n22689, n22690,
         n22691, n22692, n22693, n22694, n22695, n22696, n22697, n22698,
         n22699, n22700, n22701, n22702, n22703, n22704, n22705, n22706,
         n22707, n22708, n22709, n22710, n22711, n22712, n22713, n22714,
         n22715, n22716, n22717, n22718, n22719, n22720, n22721, n22722,
         n22723, n22724, n22725, n22726, n22727, n22728, n22729, n22730,
         n22731, n22732, n22733, n22734, n22735, n22736, n22737, n22738,
         n22739, n22740, n22741, n22742, n22743, n22744, n22745, n22746,
         n22747, n22748, n22749, n22750, n22751, n22752, n22753, n22754,
         n22755, n22756, n22757, n22758, n22759, n22760, n22761, n22762,
         n22763, n22764, n22765, n22766, n22767, n22768, n22769, n22770,
         n22771, n22772, n22773, n22774, n22775, n22776, n22777, n22778,
         n22779, n22780, n22781, n22782, n22783, n22784, n22785, n22786,
         n22787, n22788, n22789, n22790, n22791, n22792, n22793, n22794,
         n22795, n22796, n22797, n22798, n22799, n22800, n22801, n22802,
         n22803, n22804, n22805, n22806, n22807, n22808, n22809, n22810,
         n22811, n22812, n22813, n22814, n22815, n22816, n22817, n22818,
         n22819, n22820, n22821, n22822, n22823, n22824, n22825, n22826,
         n22827, n22828, n22829, n22830, n22831, n22832, n22833, n22834,
         n22835, n22836, n22837, n22838, n22839, n22840, n22841, n22842,
         n22843, n22844, n22845, n22846, n22847, n22848, n22849, n22850,
         n22851, n22852, n22853, n22854, n22855, n22856, n22857, n22858,
         n22859, n22860, n22861, n22862, n22863, n22864, n22865, n22866,
         n22867, n22868, n22869, n22870, n22871, n22872, n22873, n22874,
         n22875, n22876, n22877, n22878, n22879, n22880, n22881, n22882,
         n22883, n22884, n22885, n22886, n22887, n22888, n22889, n22890,
         n22891, n22892, n22893, n22894, n22895, n22896, n22897, n22898,
         n22899, n22900, n22901, n22902, n22903, n22904, n22905, n22906,
         n22907, n22908, n22909, n22910, n22911, n22912, n22913, n22914,
         n22915, n22916, n22917, n22918, n22919, n22920, n22921, n22922,
         n22923, n22924, n22925, n22926, n22927, n22928, n22929, n22930,
         n22931, n22932, n22933, n22934, n22935, n22936, n22937, n22938,
         n22939, n22940, n22941, n22942, n22943, n22944, n22945, n22946,
         n22947, n22948, n22949, n22950, n22951, n22952, n22953, n22954,
         n22955, n22956, n22957, n22958, n22959, n22960, n22961, n22962,
         n22963, n22964, n22965, n22966, n22967, n22968, n22969, n22970,
         n22971, n22972, n22973, n22974, n22975, n22976, n22977, n22978,
         n22979, n22980, n22981, n22982, n22983, n22984, n22985, n22986,
         n22987, n22988, n22989, n22990, n22991, n22992, n22993, n22994,
         n22995, n22996, n22997, n22998, n22999, n23000, n23001, n23002,
         n23003, n23004, n23005, n23006, n23007, n23008, n23009, n23010,
         n23011, n23012, n23013, n23014, n23015, n23016, n23017, n23018,
         n23019, n23020, n23021, n23022, n23023, n23024, n23025, n23026,
         n23027, n23028, n23029, n23030, n23031, n23032, n23033, n23034,
         n23035, n23036, n23037, n23038, n23039, n23040, n23041, n23042,
         n23043, n23044, n23045, n23046, n23047, n23048, n23049, n23050,
         n23051, n23052, n23053, n23054, n23055, n23056, n23057, n23058,
         n23059, n23060, n23061, n23062, n23063, n23064, n23065, n23066,
         n23067, n23068, n23069, n23070, n23071, n23072, n23073, n23074,
         n23075, n23076, n23077, n23078, n23079, n23080, n23081, n23082,
         n23083, n23084, n23085, n23086, n23087, n23088, n23089, n23090,
         n23091, n23092, n23093, n23094, n23095, n23096, n23097, n23098,
         n23099, n23100, n23101, n23102, n23103, n23104, n23105, n23106,
         n23107, n23108, n23109, n23110, n23111, n23112, n23113, n23114,
         n23115, n23116, n23117, n23118, n23119, n23120, n23121, n23122,
         n23123, n23124, n23125, n23126, n23127, n23128, n23129, n23130,
         n23131, n23132, n23133, n23134, n23135, n23136, n23137, n23138,
         n23139, n23140, n23141, n23142, n23143, n23144, n23145, n23146,
         n23147, n23148, n23149, n23150, n23151, n23152, n23153, n23154,
         n23155, n23156, n23157, n23158, n23159, n23160, n23161, n23162,
         n23163, n23164, n23165, n23166, n23167, n23168, n23169, n23170,
         n23171, n23172, n23173, n23174, n23175, n23176, n23177, n23178,
         n23179, n23180, n23181, n23182, n23183, n23184, n23185, n23186,
         n23187, n23188, n23189, n23190, n23191, n23192, n23193, n23194,
         n23195, n23196, n23197, n23198, n23199, n23200, n23201, n23202,
         n23203, n23204, n23205, n23206, n23207, n23208, n23209, n23210,
         n23211, n23212, n23213, n23214, n23215, n23216, n23217, n23218,
         n23219, n23220, n23221, n23222, n23223, n23224, n23225, n23226,
         n23227, n23228, n23229, n23230, n23231, n23232, n23233, n23234,
         n23235, n23236, n23237, n23238, n23239, n23240, n23241, n23242,
         n23243, n23244, n23245, n23246, n23247, n23248, n23249, n23250,
         n23251, n23252, n23253, n23254, n23255, n23256, n23257, n23258,
         n23259, n23260, n23261, n23262, n23263, n23264, n23265, n23266,
         n23267, n23268, n23269, n23270, n23271, n23272, n23273, n23274,
         n23275, n23276, n23277, n23278, n23279, n23280, n23281, n23282,
         n23283, n23284, n23285, n23286, n23287, n23288, n23289, n23290,
         n23291, n23292, n23293, n23294, n23295, n23296, n23297, n23298,
         n23299, n23300, n23301, n23302, n23303, n23304, n23305, n23306,
         n23307, n23308, n23309, n23310, n23311, n23312, n23313, n23314,
         n23315, n23316, n23317, n23318, n23319, n23320, n23321, n23322,
         n23323, n23324, n23325, n23326, n23327, n23328, n23329, n23330,
         n23331, n23332, n23333, n23334, n23335, n23336, n23337, n23338,
         n23339, n23340, n23341, n23342, n23343, n23344, n23345, n23346,
         n23347, n23348, n23349, n23350, n23351, n23352, n23353, n23354,
         n23355, n23356, n23357, n23358, n23359, n23360, n23361, n23362,
         n23363, n23364, n23365, n23366, n23367, n23368, n23369, n23370,
         n23371, n23372, n23373, n23374, n23375, n23376, n23377, n23378,
         n23379, n23380, n23381, n23382, n23383, n23384, n23385, n23386,
         n23387, n23388, n23389, n23390, n23391, n23392, n23393, n23394,
         n23395, n23396, n23397, n23398, n23399, n23400, n23401, n23402,
         n23403, n23404, n23405, n23406, n23407, n23408, n23409, n23410,
         n23411, n23412, n23413, n23414, n23415, n23416, n23417, n23418,
         n23419, n23420, n23421, n23422, n23423, n23424, n23425, n23426,
         n23427, n23428, n23429, n23430, n23431, n23432, n23433, n23434,
         n23435, n23436, n23437, n23438, n23439, n23440, n23441, n23442,
         n23443, n23444, n23445, n23446, n23447, n23448, n23449, n23450,
         n23451, n23452, n23453, n23454, n23455, n23456, n23457, n23458,
         n23459, n23460, n23461, n23462, n23463, n23464, n23465, n23466,
         n23467, n23468, n23469, n23470, n23471, n23472, n23473, n23474,
         n23475, n23476, n23477, n23478, n23479, n23480, n23481, n23482,
         n23483, n23484, n23485, n23486, n23487, n23488, n23489, n23490,
         n23491, n23492, n23493, n23494, n23495, n23496, n23497, n23498,
         n23499, n23500, n23501, n23502, n23503, n23504, n23505, n23506,
         n23507, n23508, n23509, n23510, n23511, n23512, n23513, n23514,
         n23515, n23516, n23517, n23518, n23519, n23520, n23521, n23522,
         n23523, n23524, n23525, n23526, n23527, n23528, n23529, n23530,
         n23531, n23532, n23533, n23534, n23535, n23536, n23537, n23538,
         n23539, n23540, n23541, n23542, n23543, n23544, n23545, n23546,
         n23547, n23548, n23549, n23550, n23551, n23552, n23553, n23554,
         n23555, n23556, n23557, n23558, n23559, n23560, n23561, n23562,
         n23563, n23564, n23565, n23566, n23567, n23568, n23569, n23570,
         n23571, n23572, n23573, n23574, n23575, n23576, n23577, n23578,
         n23579, n23580, n23581, n23582, n23583, n23584, n23585, n23586,
         n23587, n23588, n23589, n23590, n23591, n23592, n23593, n23594,
         n23595, n23596, n23597, n23598, n23599, n23600, n23601, n23602,
         n23603, n23604, n23605, n23606, n23607, n23608, n23609, n23610,
         n23611, n23612, n23613, n23614, n23615, n23616, n23617, n23618,
         n23619, n23620, n23621, n23622, n23623, n23624, n23625, n23626,
         n23627, n23628, n23629, n23630, n23631, n23632, n23633, n23634,
         n23635, n23636, n23637, n23638, n23639, n23640, n23641, n23642,
         n23643, n23644, n23645, n23646, n23647, n23648, n23649, n23650,
         n23651, n23652, n23653, n23654, n23655, n23656, n23657, n23658,
         n23659, n23660, n23661, n23662, n23663, n23664, n23665, n23666,
         n23667, n23668, n23669, n23670, n23671, n23672, n23673, n23674,
         n23675, n23676, n23677, n23678, n23679, n23680, n23681, n23682,
         n23683, n23684, n23685, n23686, n23687, n23688, n23689, n23690,
         n23691, n23692, n23693, n23694, n23695, n23696, n23697, n23698,
         n23699, n23700, n23701, n23702, n23703, n23704, n23705, n23706,
         n23707, n23708, n23709, n23710, n23711, n23712, n23713, n23714,
         n23715, n23716, n23717, n23718, n23719, n23720, n23721, n23722,
         n23723, n23724, n23725, n23726, n23727, n23728, n23729, n23730,
         n23731, n23732, n23733, n23734, n23735, n23736, n23737, n23738,
         n23739, n23740, n23741, n23742, n23743, n23744, n23745, n23746,
         n23747, n23748, n23749, n23750, n23751, n23752, n23753, n23754,
         n23755, n23756, n23757, n23758, n23759, n23760, n23761, n23762,
         n23763, n23764, n23765, n23766, n23767, n23768, n23769, n23770,
         n23771, n23772, n23773, n23774, n23775, n23776, n23777, n23778,
         n23779, n23780, n23781, n23782, n23783, n23784, n23785, n23786,
         n23787, n23788, n23789, n23790, n23791, n23792, n23793, n23794,
         n23795, n23796, n23797, n23798, n23799, n23800, n23801, n23802,
         n23803, n23804, n23805, n23806, n23807, n23808, n23809, n23810,
         n23811, n23812, n23813, n23814, n23815, n23816, n23817, n23818,
         n23819, n23820, n23821, n23822, n23823, n23824, n23825, n23826,
         n23827, n23828, n23829, n23830, n23831, n23832, n23833, n23834,
         n23835, n23836, n23837, n23838, n23839, n23840, n23841, n23842,
         n23843, n23844, n23845, n23846, n23847, n23848, n23849, n23850,
         n23851, n23852, n23853, n23854, n23855, n23856, n23857, n23858,
         n23859, n23860, n23861, n23862, n23863, n23864, n23865, n23866,
         n23867, n23868, n23869, n23870, n23871, n23872, n23873, n23874,
         n23875, n23876, n23877, n23878, n23879, n23880, n23881, n23882,
         n23883, n23884, n23885, n23886, n23887, n23888, n23889, n23890,
         n23891, n23892, n23893, n23894, n23895, n23896, n23897, n23898,
         n23899, n23900, n23901, n23902, n23903, n23904, n23905, n23906,
         n23907, n23908, n23909, n23910, n23911, n23912, n23913, n23914,
         n23915, n23916, n23917, n23918, n23919, n23920, n23921, n23922,
         n23923, n23924, n23925, n23926, n23927, n23928, n23929, n23930,
         n23931, n23932, n23933, n23934, n23935, n23936, n23937, n23938,
         n23939, n23940, n23941, n23942, n23943, n23944, n23945, n23946,
         n23947, n23948, n23949, n23950, n23951, n23952, n23953, n23954,
         n23955, n23956, n23957, n23958, n23959, n23960, n23961, n23962,
         n23963, n23964, n23965, n23966, n23967, n23968, n23969, n23970,
         n23971, n23972, n23973, n23974, n23975, n23976, n23977, n23978,
         n23979, n23980, n23981, n23982, n23983, n23984, n23985, n23986,
         n23987, n23988, n23989, n23990, n23991, n23992, n23993, n23994,
         n23995, n23996, n23997, n23998, n23999, n24000, n24001, n24002,
         n24003, n24004, n24005, n24006, n24007, n24008, n24009, n24010,
         n24011, n24012, n24013, n24014, n24015, n24016, n24017, n24018,
         n24019, n24020, n24021, n24022, n24023, n24024, n24025, n24026,
         n24027, n24028, n24029, n24030, n24031, n24032, n24033, n24034,
         n24035, n24036, n24037, n24038, n24039, n24040, n24041, n24042,
         n24043, n24044, n24045, n24046, n24047, n24048, n24049, n24050,
         n24051, n24052, n24053, n24054, n24055, n24056, n24057, n24058,
         n24059, n24060, n24061, n24062, n24063, n24064, n24065, n24066,
         n24067, n24068, n24069, n24070, n24071, n24072, n24073, n24074,
         n24075, n24076, n24077, n24078, n24079, n24080, n24081, n24082,
         n24083, n24084, n24085, n24086, n24087, n24088, n24089, n24090,
         n24091, n24092, n24093, n24094, n24095, n24096, n24097, n24098,
         n24099, n24100, n24101, n24102, n24103, n24104, n24105, n24106,
         n24107, n24108, n24109, n24110, n24111, n24112, n24113, n24114,
         n24115, n24116, n24117, n24118, n24119, n24120, n24121, n24122,
         n24123, n24124, n24125, n24126, n24127, n24128, n24129, n24130,
         n24131, n24132, n24133, n24134, n24135, n24136, n24137, n24138,
         n24139, n24140, n24141, n24142, n24143, n24144, n24145, n24146,
         n24147, n24148, n24149, n24150, n24151, n24152, n24153, n24154,
         n24155, n24156, n24157, n24158, n24159, n24160, n24161, n24162,
         n24163, n24164, n24165, n24166, n24167, n24168, n24169, n24170,
         n24171, n24172, n24173, n24174, n24175, n24176, n24177, n24178,
         n24179, n24180, n24181, n24182, n24183, n24184, n24185, n24186,
         n24187, n24188, n24189, n24190, n24191, n24192, n24193, n24194,
         n24195, n24196, n24197, n24198, n24199, n24200, n24201, n24202,
         n24203, n24204, n24205, n24206, n24207, n24208, n24209, n24210,
         n24211, n24212, n24213, n24214, n24215, n24216, n24217, n24218,
         n24219, n24220, n24221, n24222, n24223, n24224, n24225, n24226,
         n24227, n24228, n24229, n24230, n24231, n24232, n24233, n24234,
         n24235, n24236, n24237, n24238, n24239, n24240, n24241, n24242,
         n24243, n24244, n24245, n24246, n24247, n24248, n24249, n24250,
         n24251, n24252, n24253, n24254, n24255, n24256, n24257, n24258,
         n24259, n24260, n24261, n24262, n24263, n24264, n24265, n24266,
         n24267, n24268, n24269, n24270, n24271, n24272, n24273, n24274,
         n24275, n24276, n24277, n24278, n24279, n24280, n24281, n24282,
         n24283, n24284, n24285, n24286, n24287, n24288, n24289, n24290,
         n24291, n24292, n24293, n24294, n24295, n24296, n24297, n24298,
         n24299, n24300, n24301, n24302, n24303, n24304, n24305, n24306,
         n24307, n24308, n24309, n24310, n24311, n24312, n24313, n24314,
         n24315, n24316, n24317, n24318, n24319, n24320, n24321, n24322,
         n24323, n24324, n24325, n24326, n24327, n24328, n24329, n24330,
         n24331, n24332, n24333, n24334, n24335, n24336, n24337, n24338,
         n24339, n24340, n24341, n24342, n24343, n24344, n24345, n24346,
         n24347, n24348, n24349, n24350, n24351, n24352, n24353, n24354,
         n24355, n24356, n24357, n24358, n24359, n24360, n24361, n24362,
         n24363, n24364, n24365, n24366, n24367, n24368, n24369, n24370,
         n24371, n24372, n24373, n24374, n24375, n24376, n24377, n24378,
         n24379, n24380, n24381, n24382, n24383, n24384, n24385, n24386,
         n24387, n24388, n24389, n24390, n24391, n24392, n24393, n24394,
         n24395, n24396, n24397, n24398, n24399, n24400, n24401, n24402,
         n24403, n24404, n24405, n24406, n24407, n24408, n24409, n24410,
         n24411, n24412, n24413, n24414, n24415, n24416, n24417, n24418,
         n24419, n24420, n24421, n24422, n24423, n24424, n24425, n24426,
         n24427, n24428, n24429, n24430, n24431, n24432, n24433, n24434,
         n24435, n24436, n24437, n24438, n24439, n24440, n24441, n24442,
         n24443, n24444, n24445, n24446, n24447, n24448, n24449, n24450,
         n24451, n24452, n24453, n24454, n24455, n24456, n24457, n24458,
         n24459, n24460, n24461, n24462, n24463, n24464, n24465, n24466,
         n24467, n24468, n24469, n24470, n24471, n24472, n24473, n24474,
         n24475, n24476, n24477, n24478, n24479, n24480, n24481, n24482,
         n24483, n24484, n24485, n24486, n24487, n24488, n24489, n24490,
         n24491, n24492, n24493, n24494, n24495, n24496, n24497, n24498,
         n24499, n24500, n24501, n24502, n24503, n24504, n24505, n24506,
         n24507, n24508, n24509, n24510, n24511, n24512, n24513, n24514,
         n24515, n24516, n24517, n24518, n24519, n24520, n24521, n24522,
         n24523, n24524, n24525, n24526, n24527, n24528, n24529, n24530,
         n24531, n24532, n24533, n24534, n24535, n24536, n24537, n24538,
         n24539, n24540, n24541, n24542, n24543, n24544, n24545, n24546,
         n24547, n24548, n24549, n24550, n24551, n24552, n24553, n24554,
         n24555, n24556, n24557, n24558, n24559, n24560, n24561, n24562,
         n24563, n24564, n24565, n24566, n24567, n24568, n24569, n24570,
         n24571, n24572, n24573, n24574, n24575, n24576, n24577, n24578,
         n24579, n24580, n24581, n24582, n24583, n24584, n24585, n24586,
         n24587, n24588, n24589, n24590, n24591, n24592, n24593, n24594,
         n24595, n24596, n24597, n24598, n24599, n24600, n24601, n24602,
         n24603, n24604, n24605, n24606, n24607, n24608, n24609, n24610,
         n24611, n24612, n24613, n24614, n24615, n24616, n24617, n24618,
         n24619, n24620, n24621, n24622, n24623, n24624, n24625, n24626,
         n24627, n24628, n24629, n24630, n24631, n24632, n24633, n24634,
         n24635, n24636, n24637, n24638, n24639, n24640, n24641, n24642,
         n24643, n24644, n24645, n24646, n24647, n24648, n24649, n24650,
         n24651, n24652, n24653, n24654, n24655, n24656, n24657, n24658,
         n24659, n24660, n24661, n24662, n24663, n24664, n24665, n24666,
         n24667, n24668, n24669, n24670, n24671, n24672, n24673, n24674,
         n24675, n24676, n24677, n24678, n24679, n24680, n24681, n24682,
         n24683, n24684, n24685, n24686, n24687, n24688, n24689, n24690,
         n24691, n24692, n24693, n24694, n24695, n24696, n24697, n24698,
         n24699, n24700, n24701, n24702, n24703, n24704, n24705, n24706,
         n24707, n24708, n24709, n24710, n24711, n24712, n24713, n24714,
         n24715, n24716, n24717, n24718, n24719, n24720, n24721, n24722,
         n24723, n24724, n24725, n24726, n24727, n24728, n24729, n24730,
         n24731, n24732, n24733, n24734, n24735, n24736, n24737, n24738,
         n24739, n24740, n24741, n24742, n24743, n24744, n24745, n24746,
         n24747, n24748, n24749, n24750, n24751, n24752, n24753, n24754,
         n24755, n24756, n24757, n24758, n24759, n24760, n24761, n24762,
         n24763, n24764, n24765, n24766, n24767, n24768, n24769, n24770,
         n24771, n24772, n24773, n24774, n24775, n24776, n24777, n24778,
         n24779, n24780, n24781, n24782, n24783, n24784, n24785, n24786,
         n24787, n24788, n24789, n24790, n24791, n24792, n24793, n24794,
         n24795, n24796, n24797, n24798, n24799, n24800, n24801, n24802,
         n24803, n24804, n24805, n24806, n24807, n24808, n24809, n24810,
         n24811, n24812, n24813, n24814, n24815, n24816, n24817, n24818,
         n24819, n24820, n24821, n24822, n24823, n24824, n24825, n24826,
         n24827, n24828, n24829, n24830, n24831, n24832, n24833, n24834,
         n24835, n24836, n24837, n24838, n24839, n24840, n24841, n24842,
         n24843, n24844, n24845, n24846, n24847, n24848, n24849, n24850,
         n24851, n24852, n24853, n24854, n24855, n24856, n24857, n24858,
         n24859, n24860, n24861, n24862, n24863, n24864, n24865, n24866,
         n24867, n24868, n24869, n24870, n24871, n24872, n24873, n24874,
         n24875, n24876, n24877, n24878, n24879, n24880, n24881, n24882,
         n24883, n24884, n24885, n24886, n24887, n24888, n24889, n24890,
         n24891, n24892, n24893, n24894, n24895, n24896, n24897, n24898,
         n24899, n24900, n24901, n24902, n24903, n24904, n24905, n24906,
         n24907, n24908, n24909, n24910, n24911, n24912, n24913, n24914,
         n24915, n24916, n24917, n24918, n24919, n24920, n24921, n24922,
         n24923, n24924, n24925, n24926, n24927, n24928, n24929, n24930,
         n24931, n24932, n24933, n24934, n24935, n24936, n24937, n24938,
         n24939, n24940, n24941, n24942, n24943, n24944, n24945, n24946,
         n24947, n24948, n24949, n24950, n24951, n24952, n24953, n24954,
         n24955, n24956, n24957, n24958, n24959, n24960, n24961, n24962,
         n24963, n24964, n24965, n24966, n24967, n24968, n24969, n24970,
         n24971, n24972, n24973, n24974, n24975, n24976, n24977, n24978,
         n24979, n24980, n24981, n24982, n24983, n24984, n24985, n24986,
         n24987, n24988, n24989, n24990, n24991, n24992, n24993, n24994,
         n24995, n24996, n24997, n24998, n24999, n25000, n25001, n25002,
         n25003, n25004, n25005, n25006, n25007, n25008, n25009, n25010,
         n25011, n25012, n25013, n25014, n25015, n25016, n25017, n25018,
         n25019, n25020, n25021, n25022, n25023, n25024, n25025, n25026,
         n25027, n25028, n25029, n25030, n25031, n25032, n25033, n25034,
         n25035, n25036, n25037, n25038, n25039, n25040, n25041, n25042,
         n25043, n25044, n25045, n25046, n25047, n25048, n25049, n25050,
         n25051, n25052, n25053, n25054, n25055, n25056, n25057, n25058,
         n25059, n25060, n25061, n25062, n25063, n25064, n25065, n25066,
         n25067, n25068, n25069, n25070, n25071, n25072, n25073, n25074,
         n25075, n25076, n25077, n25078, n25079, n25080, n25081, n25082,
         n25083, n25084, n25085, n25086, n25087, n25088, n25089, n25090,
         n25091, n25092, n25093, n25094, n25095, n25096, n25097, n25098,
         n25099, n25100, n25101, n25102, n25103, n25104, n25105, n25106,
         n25107, n25108, n25109, n25110, n25111, n25112, n25113, n25114,
         n25115, n25116, n25117, n25118, n25119, n25120, n25121, n25122,
         n25123, n25124, n25125, n25126, n25127, n25128, n25129, n25130,
         n25131, n25132, n25133, n25134, n25135, n25136, n25137, n25138,
         n25139, n25140, n25141, n25142, n25143, n25144, n25145, n25146,
         n25147, n25148, n25149, n25150, n25151, n25152, n25153, n25154,
         n25155, n25156, n25157, n25158, n25159, n25160, n25161, n25162,
         n25163, n25164, n25165, n25166, n25167, n25168, n25169, n25170,
         n25171, n25172, n25173, n25174, n25175, n25176, n25177, n25178,
         n25179, n25180, n25181, n25182, n25183, n25184, n25185, n25186,
         n25187, n25188, n25189, n25190, n25191, n25192, n25193, n25194,
         n25195, n25196, n25197, n25198, n25199, n25200, n25201, n25202,
         n25203, n25204, n25205, n25206, n25207, n25208, n25209, n25210,
         n25211, n25212, n25213, n25214, n25215, n25216, n25217, n25218,
         n25219, n25220, n25221, n25222, n25223, n25224, n25225, n25226,
         n25227, n25228, n25229, n25230, n25231, n25232, n25233, n25234,
         n25235, n25236, n25237, n25238, n25239, n25240, n25241, n25242,
         n25243, n25244, n25245, n25246, n25247, n25248, n25249, n25250,
         n25251, n25252, n25253, n25254, n25255, n25256, n25257, n25258,
         n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266,
         n25267, n25268, n25269, n25270, n25271, n25272, n25273, n25274,
         n25275, n25276, n25277, n25278, n25279, n25280, n25281, n25282,
         n25283, n25284, n25285, n25286, n25287, n25288, n25289, n25290,
         n25291, n25292, n25293, n25294, n25295, n25296, n25297, n25298,
         n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25306,
         n25307, n25308, n25309, n25310, n25311, n25312, n25313, n25314,
         n25315, n25316, n25317, n25318, n25319, n25320, n25321, n25322,
         n25323, n25324, n25325, n25326, n25327, n25328, n25329, n25330,
         n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338,
         n25339, n25340, n25341, n25342, n25343, n25344, n25345, n25346,
         n25347, n25348, n25349, n25350, n25351, n25352, n25353, n25354,
         n25355, n25356, n25357, n25358, n25359, n25360, n25361, n25362,
         n25363, n25364, n25365, n25366, n25367, n25368, n25369, n25370,
         n25371, n25372, n25373, n25374, n25375, n25376, n25377, n25378,
         n25379, n25380, n25381, n25382, n25383, n25384, n25385, n25386,
         n25387, n25388, n25389, n25390, n25391, n25392, n25393, n25394,
         n25395, n25396, n25397, n25398, n25399, n25400, n25401, n25402,
         n25403, n25404, n25405, n25406, n25407, n25408, n25409, n25410,
         n25411, n25412, n25413, n25414, n25415, n25416, n25417, n25418,
         n25419, n25420, n25421, n25422, n25423, n25424, n25425, n25426,
         n25427, n25428, n25429, n25430, n25431, n25432, n25433, n25434,
         n25435, n25436, n25437, n25438, n25439, n25440, n25441, n25442,
         n25443, n25444, n25445, n25446, n25447, n25448, n25449, n25450,
         n25451, n25452, n25453, n25454, n25455, n25456, n25457, n25458,
         n25459, n25460, n25461, n25462, n25463, n25464, n25465, n25466,
         n25467, n25468, n25469, n25470, n25471, n25472, n25473, n25474,
         n25475, n25476, n25477, n25478, n25479, n25480, n25481, n25482,
         n25483, n25484, n25485, n25486, n25487, n25488, n25489, n25490,
         n25491, n25492, n25493, n25494, n25495, n25496, n25497, n25498,
         n25499, n25500, n25501, n25502, n25503, n25504, n25505, n25506,
         n25507, n25508, n25509, n25510, n25511, n25512, n25513, n25514,
         n25515, n25516, n25517, n25518, n25519, n25520, n25521, n25522,
         n25523, n25524, n25525, n25526, n25527, n25528, n25529, n25530,
         n25531, n25532, n25533, n25534, n25535, n25536, n25537, n25538,
         n25539, n25540, n25541, n25542, n25543, n25544, n25545, n25546,
         n25547, n25548, n25549, n25550, n25551, n25552, n25553, n25554,
         n25555, n25556, n25557, n25558, n25559, n25560, n25561, n25562,
         n25563, n25564, n25565, n25566, n25567, n25568, n25569, n25570,
         n25571, n25572, n25573, n25574, n25575, n25576, n25577, n25578,
         n25579, n25580, n25581, n25582, n25583, n25584, n25585, n25586,
         n25587, n25588, n25589, n25590, n25591, n25592, n25593, n25594,
         n25595, n25596, n25597, n25598, n25599, n25600, n25601, n25602,
         n25603, n25604, n25605, n25606, n25607, n25608, n25609, n25610,
         n25611, n25612, n25613, n25614, n25615, n25616, n25617, n25618,
         n25619, n25620, n25621, n25622, n25623, n25624, n25625, n25626,
         n25627, n25628, n25629, n25630, n25631, n25632, n25633, n25634,
         n25635, n25636, n25637, n25638, n25639, n25640, n25641, n25642,
         n25643, n25644, n25645, n25646, n25647, n25648, n25649, n25650,
         n25651, n25652, n25653, n25654, n25655, n25656, n25657, n25658,
         n25659, n25660, n25661, n25662, n25663, n25664, n25665, n25666,
         n25667, n25668, n25669, n25670, n25671, n25672, n25673, n25674,
         n25675, n25676, n25677, n25678, n25679, n25680, n25681, n25682,
         n25683, n25684, n25685, n25686, n25687, n25688, n25689, n25690,
         n25691, n25692, n25693, n25694, n25695, n25696, n25697, n25698,
         n25699, n25700, n25701, n25702, n25703, n25704, n25705, n25706,
         n25707, n25708, n25709, n25710, n25711, n25712, n25713, n25714,
         n25715, n25716, n25717, n25718, n25719, n25720, n25721, n25722,
         n25723, n25724, n25725, n25726, n25727, n25728, n25729, n25730,
         n25731, n25732, n25733, n25734, n25735, n25736, n25737, n25738,
         n25739, n25740, n25741, n25742, n25743, n25744, n25745, n25746,
         n25747, n25748, n25749, n25750, n25751, n25752, n25753, n25754,
         n25755, n25756, n25757, n25758, n25759, n25760, n25761, n25762,
         n25763, n25764, n25765, n25766, n25767, n25768, n25769, n25770,
         n25771, n25772, n25773, n25774, n25775, n25776, n25777, n25778,
         n25779, n25780, n25781, n25782, n25783, n25784, n25785, n25786,
         n25787, n25788, n25789, n25790, n25791, n25792, n25793, n25794,
         n25795, n25796, n25797, n25798, n25799, n25800, n25801, n25802,
         n25803, n25804, n25805, n25806, n25807, n25808, n25809, n25810,
         n25811, n25812, n25813, n25814, n25815, n25816, n25817, n25818,
         n25819, n25820, n25821, n25822, n25823, n25824, n25825, n25826,
         n25827, n25828, n25829, n25830, n25831, n25832, n25833, n25834,
         n25835, n25836, n25837, n25838, n25839, n25840, n25841, n25842,
         n25843, n25844, n25845, n25846, n25847, n25848, n25849, n25850,
         n25851, n25852, n25853, n25854, n25855, n25856, n25857, n25858,
         n25859, n25860, n25861, n25862, n25863, n25864, n25865, n25866,
         n25867, n25868, n25869, n25870, n25871, n25872, n25873, n25874,
         n25875, n25876, n25877, n25878, n25879, n25880, n25881, n25882,
         n25883, n25884, n25885, n25886, n25887, n25888, n25889, n25890,
         n25891, n25892, n25893, n25894, n25895, n25896, n25897, n25898,
         n25899, n25900, n25901, n25902, n25903, n25904, n25905, n25906,
         n25907, n25908, n25909, n25910, n25911, n25912, n25913, n25914,
         n25915, n25916, n25917, n25918, n25919, n25920, n25921, n25922,
         n25923, n25924, n25925, n25926, n25927, n25928, n25929, n25930,
         n25931, n25932, n25933, n25934, n25935, n25936, n25937, n25938,
         n25939, n25940, n25941, n25942, n25943, n25944, n25945, n25946,
         n25947, n25948, n25949, n25950, n25951, n25952, n25953, n25954,
         n25955, n25956, n25957, n25958, n25959, n25960, n25961, n25962,
         n25963, n25964, n25965, n25966, n25967, n25968, n25969, n25970,
         n25971, n25972, n25973, n25974, n25975, n25976, n25977, n25978,
         n25979, n25980, n25981, n25982, n25983, n25984, n25985, n25986,
         n25987, n25988, n25989, n25990, n25991, n25992, n25993, n25994,
         n25995, n25996, n25997, n25998, n25999, n26000, n26001, n26002,
         n26003, n26004, n26005, n26006, n26007, n26008, n26009, n26010,
         n26011, n26012, n26013, n26014, n26015, n26016, n26017, n26018,
         n26019, n26020, n26021, n26022, n26023, n26024, n26025, n26026,
         n26027, n26028, n26029, n26030, n26031, n26032, n26033, n26034,
         n26035, n26036, n26037, n26038, n26039, n26040, n26041, n26042,
         n26043, n26044, n26045, n26046, n26047, n26048, n26049, n26050,
         n26051, n26052, n26053, n26054, n26055, n26056, n26057, n26058,
         n26059, n26060, n26061, n26062, n26063, n26064, n26065, n26066,
         n26067, n26068, n26069, n26070, n26071, n26072, n26073, n26074,
         n26075, n26076, n26077, n26078, n26079, n26080, n26081, n26082,
         n26083, n26084, n26085, n26086, n26087, n26088, n26089, n26090,
         n26091, n26092, n26093, n26094, n26095, n26096, n26097, n26098,
         n26099, n26100, n26101, n26102, n26103, n26104, n26105, n26106,
         n26107, n26108, n26109, n26110, n26111, n26112, n26113, n26114,
         n26115, n26116, n26117, n26118, n26119, n26120, n26121, n26122,
         n26123, n26124, n26125, n26126, n26127, n26128, n26129, n26130,
         n26131, n26132, n26133, n26134, n26135, n26136, n26137, n26138,
         n26139, n26140, n26141, n26142, n26143, n26144, n26145, n26146,
         n26147, n26148, n26149, n26150, n26151, n26152, n26153, n26154,
         n26155, n26156, n26157, n26158, n26159, n26160, n26161, n26162,
         n26163, n26164, n26165, n26166, n26167, n26168, n26169, n26170,
         n26171, n26172, n26173, n26174, n26175, n26176, n26177, n26178,
         n26179, n26180, n26181, n26182, n26183, n26184, n26185, n26186,
         n26187, n26188, n26189, n26190, n26191, n26192, n26193, n26194,
         n26195, n26196, n26197, n26198, n26199, n26200, n26201, n26202,
         n26203, n26204, n26205, n26206, n26207, n26208, n26209, n26210,
         n26211, n26212, n26213, n26214, n26215, n26216, n26217, n26218,
         n26219, n26220, n26221, n26222, n26223, n26224, n26225, n26226,
         n26227, n26228, n26229, n26230, n26231, n26232, n26233, n26234,
         n26235, n26236, n26237, n26238, n26239, n26240, n26241, n26242,
         n26243, n26244, n26245, n26246, n26247, n26248, n26249, n26250,
         n26251, n26252, n26253, n26254, n26255, n26256, n26257, n26258,
         n26259, n26260, n26261, n26262, n26263, n26264, n26265, n26266,
         n26267, n26268, n26269, n26270, n26271, n26272, n26273, n26274,
         n26275, n26276, n26277, n26278, n26279, n26280, n26281, n26282,
         n26283, n26284, n26285, n26286, n26287, n26288, n26289, n26290,
         n26291, n26292, n26293, n26294, n26295, n26296, n26297, n26298,
         n26299, n26300, n26301, n26302, n26303, n26304, n26305, n26306,
         n26307, n26308, n26309, n26310, n26311, n26312, n26313, n26314,
         n26315, n26316, n26317, n26318, n26319, n26320, n26321, n26322,
         n26323, n26324, n26325, n26326, n26327, n26328, n26329, n26330,
         n26331, n26332, n26333, n26334, n26335, n26336, n26337, n26338,
         n26339, n26340, n26341, n26342, n26343, n26344, n26345, n26346,
         n26347, n26348, n26349, n26350, n26351, n26352, n26353, n26354,
         n26355, n26356, n26357, n26358, n26359, n26360, n26361, n26362,
         n26363, n26364, n26365, n26366, n26367, n26368, n26369, n26370,
         n26371, n26372, n26373, n26374, n26375, n26376, n26377, n26378,
         n26379, n26380, n26381, n26382, n26383, n26384, n26385, n26386,
         n26387, n26388, n26389, n26390, n26391, n26392, n26393, n26394,
         n26395, n26396, n26397, n26398, n26399, n26400, n26401, n26402,
         n26403, n26404, n26405, n26406, n26407, n26408, n26409, n26410,
         n26411, n26412, n26413, n26414, n26415, n26416, n26417, n26418,
         n26419, n26420, n26421, n26422, n26423, n26424, n26425, n26426,
         n26427, n26428, n26429, n26430, n26431, n26432, n26433, n26434,
         n26435, n26436, n26437, n26438, n26439, n26440, n26441, n26442,
         n26443, n26444, n26445, n26446, n26447, n26448, n26449, n26450,
         n26451, n26452, n26453, n26454, n26455, n26456, n26457, n26458,
         n26459, n26460, n26461, n26462, n26463, n26464, n26465, n26466,
         n26467, n26468, n26469, n26470, n26471, n26472, n26473, n26474,
         n26475, n26476, n26477, n26478, n26479, n26480, n26481, n26482,
         n26483, n26484, n26485, n26486, n26487, n26488, n26489, n26490,
         n26491, n26492, n26493, n26494, n26495, n26496, n26497, n26498,
         n26499, n26500, n26501, n26502, n26503, n26504, n26505, n26506,
         n26507, n26508, n26509, n26510, n26511, n26512, n26513, n26514,
         n26515, n26516, n26517, n26518, n26519, n26520, n26521, n26522,
         n26523, n26524, n26525, n26526, n26527, n26528, n26529, n26530,
         n26531, n26532, n26533, n26534, n26535, n26536, n26537, n26538,
         n26539, n26540, n26541, n26542, n26543, n26544, n26545, n26546,
         n26547, n26548, n26549, n26550, n26551, n26552, n26553, n26554,
         n26555, n26556, n26557, n26558, n26559, n26560, n26561, n26562,
         n26563, n26564, n26565, n26566, n26567, n26568, n26569, n26570,
         n26571, n26572, n26573, n26574, n26575, n26576, n26577, n26578,
         n26579, n26580, n26581, n26582, n26583, n26584, n26585, n26586,
         n26587, n26588, n26589, n26590, n26591, n26592, n26593, n26594,
         n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602,
         n26603, n26604, n26605, n26606, n26607, n26608, n26609, n26610,
         n26611, n26612, n26613, n26614, n26615, n26616, n26617, n26618,
         n26619, n26620, n26621, n26622, n26623, n26624, n26625, n26626,
         n26627, n26628, n26629, n26630, n26631, n26632, n26633, n26634,
         n26635, n26636, n26637, n26638, n26639, n26640, n26641, n26642,
         n26643, n26644, n26645, n26646, n26647, n26648, n26649, n26650,
         n26651, n26652, n26653, n26654, n26655, n26656, n26657, n26658,
         n26659, n26660, n26661, n26662, n26663, n26664, n26665, n26666,
         n26667, n26668, n26669, n26670, n26671, n26672, n26673, n26674,
         n26675, n26676, n26677, n26678, n26679, n26680, n26681, n26682,
         n26683, n26684, n26685, n26686, n26687, n26688, n26689, n26690,
         n26691, n26692, n26693, n26694, n26695, n26696, n26697, n26698,
         n26699, n26700, n26701, n26702, n26703, n26704, n26705, n26706,
         n26707, n26708, n26709, n26710, n26711, n26712, n26713, n26714,
         n26715, n26716, n26717, n26718, n26719, n26720, n26721, n26722,
         n26723, n26724, n26725, n26726, n26727, n26728, n26729, n26730,
         n26731, n26732, n26733, n26734, n26735, n26736, n26737, n26738,
         n26739, n26740, n26741, n26742, n26743, n26744, n26745, n26746,
         n26747, n26748, n26749, n26750, n26751, n26752, n26753, n26754,
         n26755, n26756, n26757, n26758, n26759, n26760, n26761, n26762,
         n26763, n26764, n26765, n26766, n26767, n26768, n26769, n26770,
         n26771, n26772, n26773, n26774, n26775, n26776, n26777, n26778,
         n26779, n26780, n26781, n26782, n26783, n26784, n26785, n26786,
         n26787, n26788, n26789, n26790, n26791, n26792, n26793, n26794,
         n26795, n26796, n26797, n26798, n26799, n26800, n26801, n26802,
         n26803, n26804, n26805, n26806, n26807, n26808, n26809, n26810,
         n26811, n26812, n26813, n26814, n26815, n26816, n26817, n26818,
         n26819, n26820, n26821, n26822, n26823, n26824, n26825, n26826,
         n26827, n26828, n26829, n26830, n26831, n26832, n26833, n26834,
         n26835, n26836, n26837, n26838, n26839, n26840, n26841, n26842,
         n26843, n26844, n26845, n26846, n26847, n26848, n26849, n26850,
         n26851, n26852, n26853, n26854, n26855, n26856, n26857, n26858,
         n26859, n26860, n26861, n26862, n26863, n26864, n26865, n26866,
         n26867, n26868, n26869, n26870, n26871, n26872, n26873, n26874,
         n26875, n26876, n26877, n26878, n26879, n26880, n26881, n26882,
         n26883, n26884, n26885, n26886, n26887, n26888, n26889, n26890,
         n26891, n26892, n26893, n26894, n26895, n26896, n26897, n26898,
         n26899, n26900, n26901, n26902, n26903, n26904, n26905, n26906,
         n26907, n26908, n26909, n26910, n26911, n26912, n26913, n26914,
         n26915, n26916, n26917, n26918, n26919, n26920, n26921, n26922,
         n26923, n26924, n26925, n26926, n26927, n26928, n26929, n26930,
         n26931, n26932, n26933, n26934, n26935, n26936, n26937, n26938,
         n26939, n26940, n26941, n26942, n26943, n26944, n26945, n26946,
         n26947, n26948, n26949, n26950, n26951, n26952, n26953, n26954,
         n26955, n26956, n26957, n26958, n26959, n26960, n26961, n26962,
         n26963, n26964, n26965, n26966, n26967, n26968, n26969, n26970,
         n26971, n26972, n26973, n26974, n26975, n26976, n26977, n26978,
         n26979, n26980, n26981, n26982, n26983, n26984, n26985, n26986,
         n26987, n26988, n26989, n26990, n26991, n26992, n26993, n26994,
         n26995, n26996, n26997, n26998, n26999, n27000, n27001, n27002,
         n27003, n27004, n27005, n27006, n27007, n27008, n27009, n27010,
         n27011, n27012, n27013, n27014, n27015, n27016, n27017, n27018,
         n27019, n27020, n27021, n27022, n27023, n27024, n27025, n27026,
         n27027, n27028, n27029, n27030, n27031, n27032, n27033, n27034,
         n27035, n27036, n27037, n27038, n27039, n27040, n27041, n27042,
         n27043, n27044, n27045, n27046, n27047, n27048, n27049, n27050,
         n27051, n27052, n27053, n27054, n27055, n27056, n27057, n27058,
         n27059, n27060, n27061, n27062, n27063, n27064, n27065, n27066,
         n27067, n27068, n27069, n27070, n27071, n27072, n27073, n27074,
         n27075, n27076, n27077, n27078, n27079, n27080, n27081, n27082,
         n27083, n27084, n27085, n27086, n27087, n27088, n27089, n27090,
         n27091, n27092, n27093, n27094, n27095, n27096, n27097, n27098,
         n27099, n27100, n27101, n27102, n27103, n27104, n27105, n27106,
         n27107, n27108, n27109, n27110, n27111, n27112, n27113, n27114,
         n27115, n27116, n27117, n27118, n27119, n27120, n27121, n27122,
         n27123, n27124, n27125, n27126, n27127, n27128, n27129, n27130,
         n27131, n27132, n27133, n27134, n27135, n27136, n27137, n27138,
         n27139, n27140, n27141, n27142, n27143, n27144, n27145, n27146,
         n27147, n27148, n27149, n27150, n27151, n27152, n27153, n27154,
         n27155, n27156, n27157, n27158, n27159, n27160, n27161, n27162,
         n27163, n27164, n27165, n27166, n27167, n27168, n27169, n27170,
         n27171, n27172, n27173, n27174, n27175, n27176, n27177, n27178,
         n27179, n27180, n27181, n27182, n27183, n27184, n27185, n27186,
         n27187, n27188, n27189, n27190, n27191, n27192, n27193, n27194,
         n27195, n27196, n27197, n27198, n27199, n27200, n27201, n27202,
         n27203, n27204, n27205, n27206, n27207, n27208, n27209, n27210,
         n27211, n27212, n27213, n27214, n27215, n27216, n27217, n27218,
         n27219, n27220, n27221, n27222, n27223, n27224, n27225, n27226,
         n27227, n27228, n27229, n27230, n27231, n27232, n27233, n27234,
         n27235, n27236, n27237, n27238, n27239, n27240, n27241, n27242,
         n27243, n27244, n27245, n27246, n27247, n27248, n27249, n27250,
         n27251, n27252, n27253, n27254, n27255, n27256, n27257, n27258,
         n27259, n27260, n27261, n27262, n27263, n27264, n27265, n27266,
         n27267, n27268, n27269, n27270, n27271, n27272, n27273, n27274,
         n27275, n27276, n27277, n27278, n27279, n27280, n27281, n27282,
         n27283, n27284, n27285, n27286, n27287, n27288, n27289, n27290,
         n27291, n27292, n27293, n27294, n27295, n27296, n27297, n27298,
         n27299, n27300, n27301, n27302, n27303, n27304, n27305, n27306,
         n27307, n27308, n27309, n27310, n27311, n27312, n27313, n27314,
         n27315, n27316, n27317, n27318, n27319, n27320, n27321, n27322,
         n27323, n27324, n27325, n27326, n27327, n27328, n27329, n27330,
         n27331, n27332, n27333, n27334, n27335, n27336, n27337, n27338,
         n27339, n27340, n27341, n27342, n27343, n27344, n27345, n27346,
         n27347, n27348, n27349, n27350, n27351, n27352, n27353, n27354,
         n27355, n27356, n27357, n27358, n27359, n27360, n27361, n27362,
         n27363, n27364, n27365, n27366, n27367, n27368, n27369, n27370,
         n27371, n27372, n27373, n27374, n27375, n27376, n27377, n27378,
         n27379, n27380, n27381, n27382, n27383, n27384, n27385, n27386,
         n27387, n27388, n27389, n27390, n27391, n27392, n27393, n27394,
         n27395, n27396, n27397, n27398, n27399, n27400, n27401, n27402,
         n27403, n27404, n27405, n27406, n27407, n27408, n27409, n27410,
         n27411, n27412, n27413, n27414, n27415, n27416, n27417, n27418,
         n27419, n27420, n27421, n27422, n27423, n27424, n27425, n27426,
         n27427, n27428, n27429, n27430, n27431, n27432, n27433, n27434,
         n27435, n27436, n27437, n27438, n27439, n27440, n27441, n27442,
         n27443, n27444, n27445, n27446, n27447, n27448, n27449, n27450,
         n27451, n27452, n27453, n27454, n27455, n27456, n27457, n27458,
         n27459, n27460, n27461, n27462, n27463, n27464, n27465, n27466,
         n27467, n27468, n27469, n27470, n27471, n27472, n27473, n27474,
         n27475, n27476, n27477, n27478, n27479, n27480, n27481, n27482,
         n27483, n27484, n27485, n27486, n27487, n27488, n27489, n27490,
         n27491, n27492, n27493, n27494, n27495, n27496, n27497, n27498,
         n27499, n27500, n27501, n27502, n27503, n27504, n27505, n27506,
         n27507, n27508, n27509, n27510, n27511, n27512, n27513, n27514,
         n27515, n27516, n27517, n27518, n27519, n27520, n27521, n27522,
         n27523, n27524, n27525, n27526, n27527, n27528, n27529, n27530,
         n27531, n27532, n27533, n27534, n27535, n27536, n27537, n27538,
         n27539, n27540, n27541, n27542, n27543, n27544, n27545, n27546,
         n27547, n27548, n27549, n27550, n27551, n27552, n27553, n27554,
         n27555, n27556, n27557, n27558, n27559, n27560, n27561, n27562,
         n27563, n27564, n27565, n27566, n27567, n27568, n27569, n27570,
         n27571, n27572, n27573, n27574, n27575, n27576, n27577, n27578,
         n27579, n27580, n27581, n27582, n27583, n27584, n27585, n27586,
         n27587, n27588, n27589, n27590, n27591, n27592, n27593, n27594,
         n27595, n27596, n27597, n27598, n27599, n27600, n27601, n27602,
         n27603, n27604, n27605, n27606, n27607, n27608, n27609, n27610,
         n27611, n27612, n27613, n27614, n27615, n27616, n27617, n27618,
         n27619, n27620, n27621, n27622, n27623, n27624, n27625, n27626,
         n27627, n27628, n27629, n27630, n27631, n27632, n27633, n27634,
         n27635, n27636, n27637, n27638, n27639, n27640, n27641, n27642,
         n27643, n27644, n27645, n27646, n27647, n27648, n27649, n27650,
         n27651, n27652, n27653, n27654, n27655, n27656, n27657, n27658,
         n27659, n27660, n27661, n27662, n27663, n27664, n27665, n27666,
         n27667, n27668, n27669, n27670, n27671, n27672, n27673, n27674,
         n27675, n27676, n27677, n27678, n27679, n27680, n27681, n27682,
         n27683, n27684, n27685, n27686, n27687, n27688, n27689, n27690,
         n27691, n27692, n27693, n27694, n27695, n27696, n27697, n27698,
         n27699, n27700, n27701, n27702, n27703, n27704, n27705, n27706,
         n27707, n27708, n27709, n27710, n27711, n27712, n27713, n27714,
         n27715, n27716, n27717, n27718, n27719, n27720, n27721, n27722,
         n27723, n27724, n27725, n27726, n27727, n27728, n27729, n27730,
         n27731, n27732, n27733, n27734, n27735, n27736, n27737, n27738,
         n27739, n27740, n27741, n27742, n27743, n27744, n27745, n27746,
         n27747, n27748, n27749, n27750, n27751, n27752, n27753, n27754,
         n27755, n27756, n27757, n27758, n27759, n27760, n27761, n27762,
         n27763, n27764, n27765, n27766, n27767, n27768, n27769, n27770,
         n27771, n27772, n27773, n27774, n27775, n27776, n27777, n27778,
         n27779, n27780, n27781, n27782, n27783, n27784, n27785, n27786,
         n27787, n27788, n27789, n27790, n27791, n27792, n27793, n27794,
         n27795, n27796, n27797, n27798, n27799, n27800, n27801, n27802,
         n27803, n27804, n27805, n27806, n27807, n27808, n27809, n27810,
         n27811, n27812, n27813, n27814, n27815, n27816, n27817, n27818,
         n27819, n27820, n27821, n27822, n27823, n27824, n27825, n27826,
         n27827, n27828, n27829, n27830, n27831, n27832, n27833, n27834,
         n27835, n27836, n27837, n27838, n27839, n27840, n27841, n27842,
         n27843, n27844, n27845, n27846, n27847, n27848, n27849, n27850,
         n27851, n27852, n27853, n27854, n27855, n27856, n27857, n27858,
         n27859, n27860, n27861, n27862, n27863, n27864, n27865, n27866,
         n27867, n27868, n27869, n27870, n27871, n27872, n27873, n27874,
         n27875, n27876, n27877, n27878, n27879, n27880, n27881, n27882,
         n27883, n27884, n27885, n27886, n27887, n27888, n27889, n27890,
         n27891, n27892, n27893, n27894, n27895, n27896, n27897, n27898,
         n27899, n27900, n27901, n27902, n27903, n27904, n27905, n27906,
         n27907, n27908, n27909, n27910, n27911, n27912, n27913, n27914,
         n27915, n27916, n27917, n27918, n27919, n27920, n27921, n27922,
         n27923, n27924, n27925, n27926, n27927, n27928, n27929, n27930,
         n27931, n27932, n27933, n27934, n27935, n27936, n27937, n27938,
         n27939, n27940, n27941, n27942, n27943, n27944, n27945, n27946,
         n27947, n27948, n27949, n27950, n27951, n27952, n27953, n27954,
         n27955, n27956, n27957, n27958, n27959, n27960, n27961, n27962,
         n27963, n27964, n27965, n27966, n27967, n27968, n27969, n27970,
         n27971, n27972, n27973, n27974, n27975, n27976, n27977, n27978,
         n27979, n27980, n27981, n27982, n27983, n27984, n27985, n27986,
         n27987, n27988, n27989, n27990, n27991, n27992, n27993, n27994,
         n27995, n27996, n27997, n27998, n27999, n28000, n28001, n28002,
         n28003, n28004, n28005, n28006, n28007, n28008, n28009, n28010,
         n28011, n28012, n28013, n28014, n28015, n28016, n28017, n28018,
         n28019, n28020, n28021, n28022, n28023, n28024, n28025, n28026,
         n28027, n28028, n28029, n28030, n28031, n28032, n28033, n28034,
         n28035, n28036, n28037, n28038, n28039, n28040, n28041, n28042,
         n28043, n28044, n28045, n28046, n28047, n28048, n28049, n28050,
         n28051, n28052, n28053, n28054, n28055, n28056, n28057, n28058,
         n28059, n28060, n28061, n28062, n28063, n28064, n28065, n28066,
         n28067, n28068, n28069, n28070, n28071, n28072, n28073, n28074,
         n28075, n28076, n28077, n28078, n28079, n28080, n28081, n28082,
         n28083, n28084, n28085, n28086, n28087, n28088, n28089, n28090,
         n28091, n28092, n28093, n28094, n28095, n28096, n28097, n28098,
         n28099, n28100, n28101, n28102, n28103, n28104, n28105, n28106,
         n28107, n28108, n28109, n28110, n28111, n28112, n28113, n28114,
         n28115, n28116, n28117, n28118, n28119, n28120, n28121, n28122,
         n28123, n28124, n28125, n28126, n28127, n28128, n28129, n28130,
         n28131, n28132, n28133, n28134, n28135, n28136, n28137, n28138,
         n28139, n28140, n28141, n28142, n28143, n28144, n28145, n28146,
         n28147, n28148, n28149, n28150, n28151, n28152, n28153, n28154,
         n28155, n28156, n28157, n28158, n28159, n28160, n28161, n28162,
         n28163, n28164, n28165, n28166, n28167, n28168, n28169, n28170,
         n28171, n28172, n28173, n28174, n28175, n28176, n28177, n28178,
         n28179, n28180, n28181, n28182, n28183, n28184, n28185, n28186,
         n28187, n28188, n28189, n28190, n28191, n28192, n28193, n28194,
         n28195, n28196, n28197, n28198, n28199, n28200, n28201, n28202,
         n28203, n28204, n28205, n28206, n28207, n28208, n28209, n28210,
         n28211, n28212, n28213, n28214, n28215, n28216, n28217, n28218,
         n28219, n28220, n28221, n28222, n28223, n28224, n28225, n28226,
         n28227, n28228, n28229, n28230, n28231, n28232, n28233, n28234,
         n28235, n28236, n28237, n28238, n28239, n28240, n28241, n28242,
         n28243, n28244, n28245, n28246, n28247, n28248, n28249, n28250,
         n28251, n28252, n28253, n28254, n28255, n28256, n28257, n28258,
         n28259, n28260, n28261, n28262, n28263, n28264, n28265, n28266,
         n28267, n28268, n28269, n28270, n28271, n28272, n28273, n28274,
         n28275, n28276, n28277, n28278, n28279, n28280, n28281, n28282,
         n28283, n28284, n28285, n28286, n28287, n28288, n28289, n28290,
         n28291, n28292, n28293, n28294, n28295, n28296, n28297, n28298,
         n28299, n28300, n28301, n28302, n28303, n28304, n28305, n28306,
         n28307, n28308, n28309, n28310, n28311, n28312, n28313, n28314,
         n28315, n28316, n28317, n28318, n28319, n28320, n28321, n28322,
         n28323, n28324, n28325, n28326, n28327, n28328, n28329, n28330,
         n28331, n28332, n28333, n28334, n28335, n28336, n28337, n28338,
         n28339, n28340, n28341, n28342, n28343, n28344, n28345, n28346,
         n28347, n28348, n28349, n28350, n28351, n28352, n28353, n28354,
         n28355, n28356, n28357, n28358, n28359, n28360, n28361, n28362,
         n28363, n28364, n28365, n28366, n28367, n28368, n28369, n28370,
         n28371, n28372, n28373, n28374, n28375, n28376, n28377, n28378,
         n28379, n28380, n28381, n28382, n28383, n28384, n28385, n28386,
         n28387, n28388, n28389, n28390, n28391, n28392, n28393, n28394,
         n28395, n28396, n28397, n28398, n28399, n28400, n28401, n28402,
         n28403, n28404, n28405, n28406, n28407, n28408, n28409, n28410,
         n28411, n28412, n28413, n28414, n28415, n28416, n28417, n28418,
         n28419, n28420, n28421, n28422, n28423, n28424, n28425, n28426,
         n28427, n28428, n28429, n28430, n28431, n28432, n28433, n28434,
         n28435, n28436, n28437, n28438, n28439, n28440, n28441, n28442,
         n28443, n28444, n28445, n28446, n28447, n28448, n28449, n28450,
         n28451, n28452, n28453, n28454, n28455, n28456, n28457, n28458,
         n28459, n28460, n28461, n28462, n28463, n28464, n28465, n28466,
         n28467, n28468, n28469, n28470, n28471, n28472, n28473, n28474,
         n28475, n28476, n28477, n28478, n28479, n28480, n28481, n28482,
         n28483, n28484, n28485, n28486, n28487, n28488, n28489, n28490,
         n28491, n28492, n28493, n28494, n28495, n28496, n28497, n28498,
         n28499, n28500, n28501, n28502, n28503, n28504, n28505, n28506,
         n28507, n28508, n28509, n28510, n28511, n28512, n28513, n28514,
         n28515, n28516, n28517, n28518, n28519, n28520, n28521, n28522,
         n28523, n28524, n28525, n28526, n28527, n28528, n28529, n28530,
         n28531, n28532, n28533, n28534, n28535, n28536, n28537, n28538,
         n28539, n28540, n28541, n28542, n28543, n28544, n28545, n28546,
         n28547, n28548, n28549, n28550, n28551, n28552, n28553, n28554,
         n28555, n28556, n28557, n28558, n28559, n28560, n28561, n28562,
         n28563, n28564, n28565, n28566, n28567, n28568, n28569, n28570,
         n28571, n28572, n28573, n28574, n28575, n28576, n28577, n28578,
         n28579, n28580, n28581, n28582, n28583, n28584, n28585, n28586,
         n28587, n28588, n28589, n28590, n28591, n28592, n28593, n28594,
         n28595, n28596, n28597, n28598, n28599, n28600, n28601, n28602,
         n28603, n28604, n28605, n28606, n28607, n28608, n28609, n28610,
         n28611, n28612, n28613, n28614, n28615, n28616, n28617, n28618,
         n28619, n28620, n28621, n28622, n28623, n28624, n28625, n28626,
         n28627, n28628, n28629, n28630, n28631, n28632, n28633, n28634,
         n28635, n28636, n28637, n28638, n28639, n28640, n28641, n28642,
         n28643, n28644, n28645, n28646, n28647, n28648, n28649, n28650,
         n28651, n28652, n28653, n28654, n28655, n28656, n28657, n28658,
         n28659, n28660, n28661, n28662, n28663, n28664, n28665, n28666,
         n28667, n28668, n28669, n28670, n28671, n28672, n28673, n28674,
         n28675, n28676, n28677, n28678, n28679, n28680, n28681, n28682,
         n28683, n28684, n28685, n28686, n28687, n28688, n28689, n28690,
         n28691, n28692, n28693, n28694, n28695, n28696, n28697, n28698,
         n28699, n28700, n28701, n28702, n28703, n28704, n28705, n28706,
         n28707, n28708, n28709, n28710, n28711, n28712, n28713, n28714,
         n28715, n28716, n28717, n28718, n28719, n28720, n28721, n28722,
         n28723, n28724, n28725, n28726, n28727, n28728, n28729, n28730,
         n28731, n28732, n28733, n28734, n28735, n28736, n28737, n28738,
         n28739, n28740, n28741, n28742, n28743, n28744, n28745, n28746,
         n28747, n28748, n28749, n28750, n28751, n28752, n28753, n28754,
         n28755, n28756, n28757, n28758, n28759, n28760, n28761, n28762,
         n28763, n28764, n28765, n28766, n28767, n28768, n28769, n28770,
         n28771, n28772, n28773, n28774, n28775, n28776, n28777, n28778,
         n28779, n28780, n28781, n28782, n28783, n28784, n28785, n28786,
         n28787, n28788, n28789, n28790, n28791, n28792, n28793, n28794,
         n28795, n28796, n28797, n28798, n28799, n28800, n28801, n28802,
         n28803, n28804, n28805, n28806, n28807, n28808, n28809, n28810,
         n28811, n28812, n28813, n28814, n28815, n28816, n28817, n28818,
         n28819, n28820, n28821, n28822, n28823, n28824, n28825, n28826,
         n28827, n28828, n28829, n28830, n28831, n28832, n28833, n28834,
         n28835, n28836, n28837, n28838, n28839, n28840, n28841, n28842,
         n28843, n28844, n28845, n28846, n28847, n28848, n28849, n28850,
         n28851, n28852, n28853, n28854, n28855, n28856, n28857, n28858,
         n28859, n28860, n28861, n28862, n28863, n28864, n28865, n28866,
         n28867, n28868, n28869, n28870, n28871, n28872, n28873, n28874,
         n28875, n28876, n28877, n28878, n28879, n28880, n28881, n28882,
         n28883, n28884, n28885, n28886, n28887, n28888, n28889, n28890,
         n28891, n28892, n28893, n28894, n28895, n28896, n28897, n28898,
         n28899, n28900, n28901, n28902, n28903, n28904, n28905, n28906,
         n28907, n28908, n28909, n28910, n28911, n28912, n28913, n28914,
         n28915, n28916, n28917, n28918, n28919, n28920, n28921, n28922,
         n28923, n28924, n28925, n28926, n28927, n28928, n28929, n28930,
         n28931, n28932, n28933, n28934, n28935, n28936, n28937, n28938,
         n28939, n28940, n28941, n28942, n28943, n28944, n28945, n28946,
         n28947, n28948, n28949, n28950, n28951, n28952, n28953, n28954,
         n28955, n28956, n28957, n28958, n28959, n28960, n28961, n28962,
         n28963, n28964, n28965, n28966, n28967, n28968, n28969, n28970,
         n28971, n28972, n28973, n28974, n28975, n28976, n28977, n28978,
         n28979, n28980, n28981, n28982, n28983, n28984, n28985, n28986,
         n28987, n28988, n28989, n28990, n28991, n28992, n28993, n28994,
         n28995, n28996, n28997, n28998, n28999, n29000, n29001, n29002,
         n29003, n29004, n29005, n29006, n29007, n29008, n29009, n29010,
         n29011, n29012, n29013, n29014, n29015, n29016, n29017, n29018,
         n29019, n29020, n29021, n29022, n29023, n29024, n29025, n29026,
         n29027, n29028, n29029, n29030, n29031, n29032, n29033, n29034,
         n29035, n29036, n29037, n29038, n29039, n29040, n29041, n29042,
         n29043, n29044, n29045, n29046, n29047, n29048, n29049, n29050,
         n29051, n29052, n29053, n29054, n29055, n29056, n29057, n29058,
         n29059, n29060, n29061, n29062, n29063, n29064, n29065, n29066,
         n29067, n29068, n29069, n29070, n29071, n29072, n29073, n29074,
         n29075, n29076, n29077, n29078, n29079, n29080, n29081, n29082,
         n29083, n29084, n29085, n29086, n29087, n29088, n29089, n29090,
         n29091, n29092, n29093, n29094, n29095, n29096, n29097, n29098,
         n29099, n29100, n29101, n29102, n29103, n29104, n29105, n29106,
         n29107, n29108, n29109, n29110, n29111, n29112, n29113, n29114,
         n29115, n29116, n29117, n29118, n29119, n29120, n29121, n29122,
         n29123, n29124, n29125, n29126, n29127, n29128, n29129, n29130,
         n29131, n29132, n29133, n29134, n29135, n29136, n29137, n29138,
         n29139, n29140, n29141, n29142, n29143, n29144, n29145, n29146,
         n29147, n29148, n29149, n29150, n29151, n29152, n29153, n29154,
         n29155, n29156, n29157, n29158, n29159, n29160, n29161, n29162,
         n29163, n29164, n29165, n29166, n29167, n29168, n29169, n29170,
         n29171, n29172, n29173, n29174, n29175, n29176, n29177, n29178,
         n29179, n29180, n29181, n29182, n29183, n29184, n29185, n29186,
         n29187, n29188, n29189, n29190, n29191, n29192, n29193, n29194,
         n29195, n29196, n29197, n29198, n29199, n29200, n29201, n29202,
         n29203, n29204, n29205, n29206, n29207, n29208, n29209, n29210,
         n29211, n29212, n29213, n29214, n29215, n29216, n29217, n29218,
         n29219, n29220, n29221, n29222, n29223, n29224, n29225, n29226,
         n29227, n29228, n29229, n29230, n29231, n29232, n29233, n29234,
         n29235, n29236, n29237, n29238, n29239, n29240, n29241, n29242,
         n29243, n29244, n29245, n29246, n29247, n29248, n29249, n29250,
         n29251, n29252, n29253, n29254, n29255, n29256, n29257, n29258,
         n29259, n29260, n29261, n29262, n29263, n29264, n29265, n29266,
         n29267, n29268, n29269, n29270, n29271, n29272, n29273, n29274,
         n29275, n29276, n29277, n29278, n29279, n29280, n29281, n29282,
         n29283, n29284, n29285, n29286, n29287, n29288, n29289, n29290,
         n29291, n29292, n29293, n29294, n29295, n29296, n29297, n29298,
         n29299, n29300, n29301, n29302, n29303, n29304, n29305, n29306,
         n29307, n29308, n29309, n29310, n29311, n29312, n29313, n29314,
         n29315, n29316, n29317, n29318, n29319, n29320, n29321, n29322,
         n29323, n29324, n29325, n29326, n29327, n29328, n29329, n29330,
         n29331, n29332, n29333, n29334, n29335, n29336, n29337, n29338,
         n29339, n29340, n29341, n29342, n29343, n29344, n29345, n29346,
         n29347, n29348, n29349, n29350, n29351, n29352, n29353, n29354,
         n29355, n29356, n29357, n29358, n29359, n29360, n29361, n29362,
         n29363, n29364, n29365, n29366, n29367, n29368, n29369, n29370,
         n29371, n29372, n29373, n29374, n29375, n29376, n29377, n29378,
         n29379, n29380, n29381, n29382, n29383, n29384, n29385, n29386,
         n29387, n29388, n29389, n29390, n29391, n29392, n29393, n29394,
         n29395, n29396, n29397, n29398, n29399, n29400, n29401, n29402,
         n29403, n29404, n29405, n29406, n29407, n29408, n29409, n29410,
         n29411, n29412, n29413, n29414, n29415, n29416, n29417, n29418,
         n29419, n29420, n29421, n29422, n29423, n29424, n29425, n29426,
         n29427, n29428, n29429, n29430, n29431, n29432, n29433, n29434,
         n29435, n29436, n29437, n29438, n29439, n29440, n29441, n29442,
         n29443, n29444, n29445, n29446, n29447, n29448, n29449, n29450,
         n29451, n29452, n29453, n29454, n29455, n29456, n29457, n29458,
         n29459, n29460, n29461, n29462, n29463, n29464, n29465, n29466,
         n29467, n29468, n29469, n29470, n29471, n29472, n29473, n29474,
         n29475, n29476, n29477, n29478, n29479, n29480, n29481, n29482,
         n29483, n29484, n29485, n29486, n29487, n29488, n29489, n29490,
         n29491, n29492, n29493, n29494, n29495, n29496, n29497, n29498,
         n29499, n29500, n29501, n29502, n29503, n29504, n29505, n29506,
         n29507, n29508, n29509, n29510, n29511, n29512, n29513, n29514,
         n29515, n29516, n29517, n29518, n29519, n29520, n29521, n29522,
         n29523, n29524, n29525, n29526, n29527, n29528, n29529, n29530,
         n29531;

  DFF ebreg_reg ( .D(n5), .CLK(clk), .RST(rst), .Q(ebreg) );
  DFF greg_reg ( .D(n4), .CLK(clk), .RST(rst), .Q(g) );
  ANDN U10 ( .B(n15287), .A(n15286), .Z(n24763) );
  ANDN U11 ( .B(n15229), .A(n15228), .Z(n24827) );
  ANDN U12 ( .B(n15185), .A(n15184), .Z(n24871) );
  ANDN U13 ( .B(n15143), .A(n15142), .Z(n24911) );
  ANDN U14 ( .B(n15103), .A(n15102), .Z(n24951) );
  ANDN U15 ( .B(n15063), .A(n15062), .Z(n24991) );
  ANDN U16 ( .B(n15025), .A(n15024), .Z(n25031) );
  ANDN U17 ( .B(n14946), .A(n14945), .Z(n25123) );
  ANDN U18 ( .B(n14906), .A(n14905), .Z(n25163) );
  ANDN U19 ( .B(n14873), .A(n14872), .Z(n25199) );
  NANDN U20 ( .A(n14648), .B(n14649), .Z(n25449) );
  NANDN U21 ( .A(n14595), .B(n14596), .Z(n25501) );
  ANDN U22 ( .B(n14199), .A(n14198), .Z(n25871) );
  ANDN U23 ( .B(n14165), .A(n14164), .Z(n25891) );
  ANDN U24 ( .B(n14140), .A(n14139), .Z(n25902) );
  ANDN U25 ( .B(n14110), .A(n14109), .Z(n25919) );
  ANDN U26 ( .B(n14044), .A(n14043), .Z(n25973) );
  ANDN U27 ( .B(n13915), .A(n13914), .Z(n26155) );
  NANDN U28 ( .A(n13892), .B(n13893), .Z(n26176) );
  ANDN U29 ( .B(n13421), .A(n13420), .Z(n26913) );
  ANDN U30 ( .B(n12881), .A(n12880), .Z(n8) );
  NANDN U31 ( .A(n12883), .B(n12882), .Z(n9) );
  AND U32 ( .A(n8), .B(n9), .Z(n27557) );
  ANDN U33 ( .B(n12771), .A(n12770), .Z(n27700) );
  NOR U34 ( .A(n12592), .B(n12593), .Z(n27962) );
  NANDN U35 ( .A(n15473), .B(n15474), .Z(n24557) );
  NANDN U36 ( .A(n15326), .B(n15327), .Z(n24721) );
  ANDN U37 ( .B(n15263), .A(n15262), .Z(n24787) );
  ANDN U38 ( .B(n15225), .A(n15224), .Z(n24831) );
  ANDN U39 ( .B(n15166), .A(n15165), .Z(n24887) );
  ANDN U40 ( .B(n15135), .A(n15134), .Z(n24919) );
  ANDN U41 ( .B(n15096), .A(n15095), .Z(n24959) );
  ANDN U42 ( .B(n15056), .A(n15055), .Z(n24999) );
  ANDN U43 ( .B(n15017), .A(n15016), .Z(n25039) );
  ANDN U44 ( .B(n14991), .A(n14990), .Z(n25079) );
  XNOR U45 ( .A(y[296]), .B(x[296]), .Z(n10) );
  NAND U46 ( .A(n14944), .B(n10), .Z(n25125) );
  ANDN U47 ( .B(n14902), .A(n14901), .Z(n25167) );
  ANDN U48 ( .B(n14869), .A(n14868), .Z(n25203) );
  NANDN U49 ( .A(n14810), .B(n14811), .Z(n25257) );
  NANDN U50 ( .A(n14640), .B(n14641), .Z(n25457) );
  NANDN U51 ( .A(n14591), .B(n14592), .Z(n25505) );
  NANDN U52 ( .A(n14521), .B(n14522), .Z(n25560) );
  NANDN U53 ( .A(n14307), .B(n14308), .Z(n25774) );
  XNOR U54 ( .A(y[684]), .B(x[684]), .Z(n11) );
  NAND U55 ( .A(n14232), .B(n11), .Z(n25852) );
  ANDN U56 ( .B(n16238), .A(n16237), .Z(n25872) );
  ANDN U57 ( .B(n14163), .A(n14162), .Z(n25892) );
  ANDN U58 ( .B(n14136), .A(n14135), .Z(n25904) );
  ANDN U59 ( .B(n14108), .A(n14107), .Z(n25920) );
  XNOR U60 ( .A(y[812]), .B(x[812]), .Z(n12) );
  NAND U61 ( .A(n14042), .B(n12), .Z(n25975) );
  ANDN U62 ( .B(n13911), .A(n13910), .Z(n26157) );
  NANDN U63 ( .A(n13888), .B(n13889), .Z(n26178) );
  ANDN U64 ( .B(n16772), .A(n16771), .Z(n26208) );
  ANDN U65 ( .B(n13854), .A(n13853), .Z(n26221) );
  ANDN U66 ( .B(n13756), .A(n13755), .Z(n24452) );
  NANDN U67 ( .A(n13501), .B(n13502), .Z(n26773) );
  ANDN U68 ( .B(n13480), .A(n13479), .Z(n26811) );
  ANDN U69 ( .B(n13419), .A(n13418), .Z(n26914) );
  ANDN U70 ( .B(n18391), .A(n18390), .Z(n27097) );
  ANDN U71 ( .B(n13194), .A(n13193), .Z(n27182) );
  NAND U72 ( .A(n12881), .B(n12878), .Z(n13) );
  ANDN U73 ( .B(n13), .A(n12879), .Z(n27558) );
  ANDN U74 ( .B(n12849), .A(n19217), .Z(n27587) );
  ANDN U75 ( .B(n12767), .A(n12766), .Z(n27704) );
  NANDN U76 ( .A(n24222), .B(n12591), .Z(n27964) );
  ANDN U77 ( .B(n12539), .A(n12538), .Z(n28044) );
  ANDN U78 ( .B(n24173), .A(n12444), .Z(n28158) );
  NANDN U79 ( .A(n15469), .B(n15470), .Z(n24561) );
  NANDN U80 ( .A(n15429), .B(n15430), .Z(n24601) );
  ANDN U81 ( .B(n15305), .A(n15304), .Z(n24747) );
  XNOR U82 ( .A(y[128]), .B(x[128]), .Z(n14) );
  NAND U83 ( .A(n15261), .B(n14), .Z(n24789) );
  ANDN U84 ( .B(n15218), .A(n15217), .Z(n24839) );
  ANDN U85 ( .B(n15162), .A(n15161), .Z(n24891) );
  ANDN U86 ( .B(n15131), .A(n15130), .Z(n24923) );
  ANDN U87 ( .B(n15092), .A(n15091), .Z(n24963) );
  ANDN U88 ( .B(n15052), .A(n15051), .Z(n25003) );
  XNOR U89 ( .A(y[254]), .B(x[254]), .Z(n15) );
  NAND U90 ( .A(n15015), .B(n15), .Z(n25041) );
  ANDN U91 ( .B(n14987), .A(n14986), .Z(n25083) );
  ANDN U92 ( .B(n14943), .A(n14942), .Z(n25127) );
  NANDN U93 ( .A(n14899), .B(n14900), .Z(n25169) );
  NANDN U94 ( .A(x[337]), .B(y[337]), .Z(n16) );
  ANDN U95 ( .B(n16), .A(n14865), .Z(n25207) );
  NANDN U96 ( .A(n14806), .B(n14807), .Z(n25261) );
  NANDN U97 ( .A(n14636), .B(n14637), .Z(n25461) );
  NANDN U98 ( .A(n14587), .B(n14588), .Z(n25509) );
  NANDN U99 ( .A(n14517), .B(n14518), .Z(n25564) );
  NANDN U100 ( .A(n14485), .B(n14486), .Z(n25596) );
  NANDN U101 ( .A(n14387), .B(n14388), .Z(n25694) );
  NANDN U102 ( .A(n14347), .B(n14348), .Z(n25734) );
  NANDN U103 ( .A(n14299), .B(n14300), .Z(n25782) );
  XNOR U104 ( .A(x[686]), .B(y[686]), .Z(n17) );
  ANDN U105 ( .B(n17), .A(n16195), .Z(n25854) );
  NANDN U106 ( .A(x[712]), .B(y[712]), .Z(n18) );
  ANDN U107 ( .B(n18), .A(n14191), .Z(n25877) );
  NOR U108 ( .A(n16276), .B(n16277), .Z(n25893) );
  ANDN U109 ( .B(n14134), .A(n14133), .Z(n25905) );
  ANDN U110 ( .B(n14106), .A(n14105), .Z(n25921) );
  ANDN U111 ( .B(n14041), .A(n14040), .Z(n25977) );
  NANDN U112 ( .A(n13992), .B(n13993), .Z(n26068) );
  NANDN U113 ( .A(n13908), .B(n13909), .Z(n26158) );
  NANDN U114 ( .A(n13884), .B(n13885), .Z(n26180) );
  NANDN U115 ( .A(n13867), .B(n13868), .Z(n26209) );
  ANDN U116 ( .B(n13851), .A(n13850), .Z(n19) );
  AND U117 ( .A(n13852), .B(n19), .Z(n26222) );
  NANDN U118 ( .A(n13753), .B(n13754), .Z(n26337) );
  NOR U119 ( .A(n13499), .B(n13498), .Z(n20) );
  NANDN U120 ( .A(n13496), .B(n13497), .Z(n21) );
  NAND U121 ( .A(n20), .B(n21), .Z(n26778) );
  ANDN U122 ( .B(n17884), .A(n17883), .Z(n26812) );
  ANDN U123 ( .B(n13417), .A(n13416), .Z(n26915) );
  ANDN U124 ( .B(n13343), .A(n13342), .Z(n26995) );
  NOR U125 ( .A(n18290), .B(n18291), .Z(n27039) );
  ANDN U126 ( .B(n13291), .A(n13290), .Z(n27061) );
  ANDN U127 ( .B(n13260), .A(n13259), .Z(n27098) );
  ANDN U128 ( .B(n13222), .A(n13221), .Z(n27141) );
  NANDN U129 ( .A(n13191), .B(n13192), .Z(n27183) );
  NOR U130 ( .A(n18586), .B(n18587), .Z(n27237) );
  ANDN U131 ( .B(n13124), .A(n13123), .Z(n27255) );
  ANDN U132 ( .B(n12877), .A(n12876), .Z(n27559) );
  ANDN U133 ( .B(n12848), .A(n12847), .Z(n27589) );
  ANDN U134 ( .B(n12761), .A(n12760), .Z(n27710) );
  ANDN U135 ( .B(n12590), .A(n12589), .Z(n24224) );
  ANDN U136 ( .B(n12522), .A(n12521), .Z(n28058) );
  ANDN U137 ( .B(n20269), .A(n20268), .Z(n22) );
  NANDN U138 ( .A(n20271), .B(n20270), .Z(n23) );
  AND U139 ( .A(n22), .B(n23), .Z(n28170) );
  NANDN U140 ( .A(n15465), .B(n15466), .Z(n24565) );
  NANDN U141 ( .A(n15425), .B(n15426), .Z(n24605) );
  NANDN U142 ( .A(n15393), .B(n15394), .Z(n24637) );
  NANDN U143 ( .A(n15338), .B(n15339), .Z(n24709) );
  ANDN U144 ( .B(n15301), .A(n15300), .Z(n24751) );
  ANDN U145 ( .B(n15260), .A(n15259), .Z(n24791) );
  ANDN U146 ( .B(n15214), .A(n15213), .Z(n24843) );
  XNOR U147 ( .A(y[180]), .B(x[180]), .Z(n24) );
  NAND U148 ( .A(n15160), .B(n24), .Z(n24893) );
  ANDN U149 ( .B(n15127), .A(n15126), .Z(n24927) );
  ANDN U150 ( .B(n15088), .A(n15087), .Z(n24967) );
  ANDN U151 ( .B(n15048), .A(n15047), .Z(n25007) );
  ANDN U152 ( .B(n15014), .A(n15013), .Z(n25043) );
  ANDN U153 ( .B(n14983), .A(n14982), .Z(n25087) );
  ANDN U154 ( .B(n14935), .A(n14934), .Z(n25135) );
  NANDN U155 ( .A(x[318]), .B(y[318]), .Z(n25) );
  ANDN U156 ( .B(n25), .A(n14898), .Z(n25171) );
  NANDN U157 ( .A(y[337]), .B(x[337]), .Z(n26) );
  ANDN U158 ( .B(n26), .A(n14864), .Z(n25209) );
  NANDN U159 ( .A(n14802), .B(n14803), .Z(n25265) );
  NANDN U160 ( .A(n14758), .B(n14759), .Z(n25329) );
  NANDN U161 ( .A(n14688), .B(n14689), .Z(n25409) );
  NANDN U162 ( .A(n14632), .B(n14633), .Z(n25465) );
  NANDN U163 ( .A(n14567), .B(n14568), .Z(n25529) );
  NANDN U164 ( .A(n14513), .B(n14514), .Z(n25568) );
  NANDN U165 ( .A(n14481), .B(n14482), .Z(n25600) );
  NANDN U166 ( .A(n14383), .B(n14384), .Z(n25698) );
  NANDN U167 ( .A(n14339), .B(n14340), .Z(n25742) );
  NANDN U168 ( .A(n14295), .B(n14296), .Z(n25786) );
  NANDN U169 ( .A(n14267), .B(n14268), .Z(n25818) );
  ANDN U170 ( .B(n14227), .A(n14226), .Z(n25855) );
  ANDN U171 ( .B(n16248), .A(n16247), .Z(n25878) );
  NOR U172 ( .A(n14158), .B(n14159), .Z(n25894) );
  NANDN U173 ( .A(x[748]), .B(y[748]), .Z(n27) );
  ANDN U174 ( .B(n27), .A(n14132), .Z(n25906) );
  ANDN U175 ( .B(n14102), .A(n14101), .Z(n25922) );
  ANDN U176 ( .B(n14086), .A(n14085), .Z(n25938) );
  NANDN U177 ( .A(n14038), .B(n14039), .Z(n25979) );
  NANDN U178 ( .A(n13988), .B(n13989), .Z(n26070) );
  ANDN U179 ( .B(n13960), .A(n13959), .Z(n26106) );
  ANDN U180 ( .B(n13907), .A(n13906), .Z(n26159) );
  NOR U181 ( .A(n13882), .B(n13883), .Z(n26181) );
  ANDN U182 ( .B(n13866), .A(n13865), .Z(n26210) );
  NAND U183 ( .A(n13848), .B(n13849), .Z(n28) );
  NANDN U184 ( .A(n13847), .B(n28), .Z(n29) );
  NAND U185 ( .A(n13852), .B(n29), .Z(n30) );
  NANDN U186 ( .A(n13846), .B(n30), .Z(n26223) );
  ANDN U187 ( .B(n13839), .A(n13838), .Z(n26243) );
  NANDN U188 ( .A(n13810), .B(n13811), .Z(n26280) );
  ANDN U189 ( .B(n13792), .A(n13791), .Z(n31) );
  NANDN U190 ( .A(n13794), .B(n13793), .Z(n32) );
  AND U191 ( .A(n31), .B(n32), .Z(n26293) );
  NANDN U192 ( .A(n13749), .B(n13750), .Z(n26339) );
  ANDN U193 ( .B(n13725), .A(n13724), .Z(n26371) );
  ANDN U194 ( .B(n13646), .A(x[1286]), .Z(n33) );
  NAND U195 ( .A(y[1286]), .B(n33), .Z(n34) );
  ANDN U196 ( .B(n34), .A(n13645), .Z(n35) );
  NAND U197 ( .A(n13644), .B(n35), .Z(n26510) );
  NANDN U198 ( .A(n13625), .B(n13626), .Z(n26523) );
  ANDN U199 ( .B(n13585), .A(n13584), .Z(n26590) );
  NAND U200 ( .A(n13544), .B(n13545), .Z(n36) );
  ANDN U201 ( .B(n36), .A(n13546), .Z(n26692) );
  OR U202 ( .A(n13498), .B(n13494), .Z(n37) );
  AND U203 ( .A(n13495), .B(n37), .Z(n26779) );
  ANDN U204 ( .B(n13478), .A(n13477), .Z(n26813) );
  ANDN U205 ( .B(n13453), .A(n13452), .Z(n26843) );
  ANDN U206 ( .B(n13442), .A(n13441), .Z(n26874) );
  NOR U207 ( .A(n13412), .B(n13413), .Z(n26921) );
  ANDN U208 ( .B(n13341), .A(n13340), .Z(n26996) );
  NOR U209 ( .A(n18247), .B(n18248), .Z(n27011) );
  NANDN U210 ( .A(n13309), .B(n13310), .Z(n27046) );
  NANDN U211 ( .A(n13288), .B(n13289), .Z(n27062) );
  ANDN U212 ( .B(n13268), .A(n13267), .Z(n27086) );
  ANDN U213 ( .B(n13253), .A(n13252), .Z(n27107) );
  ANDN U214 ( .B(n13243), .A(n13242), .Z(n27114) );
  ANDN U215 ( .B(n13220), .A(n13219), .Z(n27145) );
  ANDN U216 ( .B(n13202), .A(n13201), .Z(n27170) );
  NOR U217 ( .A(n18511), .B(n18512), .Z(n27193) );
  ANDN U218 ( .B(n13170), .A(n13169), .Z(n27209) );
  ANDN U219 ( .B(n13136), .A(n13135), .Z(n27245) );
  ANDN U220 ( .B(n13120), .A(n13119), .Z(n27257) );
  NANDN U221 ( .A(n13084), .B(n13085), .Z(n27311) );
  NAND U222 ( .A(n13064), .B(n13063), .Z(n38) );
  ANDN U223 ( .B(n38), .A(n13065), .Z(n27333) );
  ANDN U224 ( .B(n13008), .A(n13007), .Z(n27405) );
  ANDN U225 ( .B(n12982), .A(n12981), .Z(n27436) );
  ANDN U226 ( .B(n12954), .A(n12953), .Z(n27473) );
  ANDN U227 ( .B(n12875), .A(n12874), .Z(n27560) );
  NANDN U228 ( .A(n12845), .B(n12846), .Z(n27590) );
  ANDN U229 ( .B(n12813), .A(n12812), .Z(n27633) );
  NANDN U230 ( .A(n12758), .B(n12759), .Z(n27712) );
  NANDN U231 ( .A(n12704), .B(n12703), .Z(n39) );
  NAND U232 ( .A(n12705), .B(n39), .Z(n40) );
  NAND U233 ( .A(n12702), .B(n40), .Z(n27812) );
  NANDN U234 ( .A(n19861), .B(n19862), .Z(n27965) );
  NAND U235 ( .A(n12533), .B(n12534), .Z(n41) );
  ANDN U236 ( .B(n41), .A(n12535), .Z(n28046) );
  ANDN U237 ( .B(n12519), .A(n12518), .Z(n28064) );
  ANDN U238 ( .B(n12471), .A(n12470), .Z(n28118) );
  ANDN U239 ( .B(n12451), .A(n12450), .Z(n24179) );
  NAND U240 ( .A(n12433), .B(n20269), .Z(n42) );
  AND U241 ( .A(n12434), .B(n42), .Z(n28171) );
  NANDN U242 ( .A(n12356), .B(n12357), .Z(n28306) );
  NANDN U243 ( .A(n12314), .B(n12315), .Z(n28353) );
  AND U244 ( .A(n20811), .B(n12229), .Z(n43) );
  NANDN U245 ( .A(n12227), .B(n12228), .Z(n44) );
  NAND U246 ( .A(n43), .B(n44), .Z(n28461) );
  NANDN U247 ( .A(n15441), .B(n15442), .Z(n24589) );
  NANDN U248 ( .A(n15401), .B(n15402), .Z(n24629) );
  NANDN U249 ( .A(n15369), .B(n15370), .Z(n24669) );
  NANDN U250 ( .A(n15322), .B(n15323), .Z(n24725) );
  ANDN U251 ( .B(n15283), .A(n15282), .Z(n24767) );
  ANDN U252 ( .B(n15252), .A(n15251), .Z(n24799) );
  ANDN U253 ( .B(n15206), .A(n15205), .Z(n24851) );
  ANDN U254 ( .B(n15159), .A(n15158), .Z(n24895) );
  XNOR U255 ( .A(y[198]), .B(x[198]), .Z(n45) );
  NAND U256 ( .A(n15125), .B(n45), .Z(n24929) );
  ANDN U257 ( .B(n15084), .A(n15083), .Z(n24971) );
  ANDN U258 ( .B(n15044), .A(n15043), .Z(n25011) );
  ANDN U259 ( .B(n15010), .A(n15009), .Z(n25047) );
  XNOR U260 ( .A(y[278]), .B(x[278]), .Z(n46) );
  NAND U261 ( .A(n14981), .B(n46), .Z(n25089) );
  XNOR U262 ( .A(y[302]), .B(x[302]), .Z(n47) );
  NAND U263 ( .A(n14933), .B(n47), .Z(n25137) );
  XNOR U264 ( .A(y[320]), .B(x[320]), .Z(n48) );
  NAND U265 ( .A(n14897), .B(n48), .Z(n25173) );
  NANDN U266 ( .A(n14862), .B(n14863), .Z(n25217) );
  NANDN U267 ( .A(n14838), .B(n14839), .Z(n25240) );
  NANDN U268 ( .A(n14794), .B(n14795), .Z(n25273) );
  NANDN U269 ( .A(n14746), .B(n14747), .Z(n25341) );
  NANDN U270 ( .A(n14676), .B(n14677), .Z(n25421) );
  NANDN U271 ( .A(n14628), .B(n14629), .Z(n25469) );
  NANDN U272 ( .A(n14583), .B(n14584), .Z(n25513) );
  NANDN U273 ( .A(n14557), .B(n14558), .Z(n25537) );
  NANDN U274 ( .A(n14509), .B(n14510), .Z(n25572) );
  NANDN U275 ( .A(n14469), .B(n14470), .Z(n25612) );
  NANDN U276 ( .A(n14417), .B(n14418), .Z(n25658) );
  NANDN U277 ( .A(n14379), .B(n14380), .Z(n25702) );
  NANDN U278 ( .A(n14335), .B(n14336), .Z(n25746) );
  NANDN U279 ( .A(n14291), .B(n14292), .Z(n25790) );
  NANDN U280 ( .A(n14263), .B(n14264), .Z(n25822) );
  NOR U281 ( .A(n14224), .B(n14225), .Z(n25860) );
  ANDN U282 ( .B(n14190), .A(n14189), .Z(n25879) );
  ANDN U283 ( .B(n14153), .A(n14152), .Z(n25896) );
  NOR U284 ( .A(n16302), .B(n16303), .Z(n25907) );
  NOR U285 ( .A(n16329), .B(n16330), .Z(n25923) );
  NANDN U286 ( .A(n14078), .B(n14079), .Z(n25947) );
  ANDN U287 ( .B(n14037), .A(n14036), .Z(n25981) );
  ANDN U288 ( .B(n13987), .A(n13986), .Z(n26071) );
  ANDN U289 ( .B(n13978), .A(n13977), .Z(n26087) );
  ANDN U290 ( .B(n13956), .A(n13955), .Z(n26111) );
  ANDN U291 ( .B(n13937), .A(n13936), .Z(n26124) );
  NANDN U292 ( .A(n13900), .B(n13901), .Z(n26162) );
  NOR U293 ( .A(n16695), .B(n16696), .Z(n26182) );
  NOR U294 ( .A(n13876), .B(n13877), .Z(n26191) );
  ANDN U295 ( .B(n13862), .A(n13861), .Z(n26212) );
  ANDN U296 ( .B(n13845), .A(n13844), .Z(n26224) );
  NOR U297 ( .A(n13834), .B(n13835), .Z(n26245) );
  ANDN U298 ( .B(n13821), .A(n13820), .Z(n26263) );
  ANDN U299 ( .B(n13809), .A(n13808), .Z(n26281) );
  ANDN U300 ( .B(n13787), .A(n13786), .Z(n26295) );
  ANDN U301 ( .B(n17030), .A(n17029), .Z(n26340) );
  ANDN U302 ( .B(n13741), .A(n13740), .Z(n26349) );
  NANDN U303 ( .A(n13722), .B(n13723), .Z(n26372) );
  NANDN U304 ( .A(n13705), .B(n13704), .Z(n49) );
  ANDN U305 ( .B(n49), .A(n13706), .Z(n26391) );
  NANDN U306 ( .A(n13645), .B(n13642), .Z(n50) );
  ANDN U307 ( .B(n50), .A(n13643), .Z(n26511) );
  ANDN U308 ( .B(n13624), .A(n13623), .Z(n26524) );
  ANDN U309 ( .B(n13581), .A(n13580), .Z(n26597) );
  NANDN U310 ( .A(n13540), .B(n13539), .Z(n51) );
  ANDN U311 ( .B(n51), .A(n13541), .Z(n26699) );
  ANDN U312 ( .B(n13532), .A(n13531), .Z(n26718) );
  NANDN U313 ( .A(n13521), .B(n13520), .Z(n52) );
  ANDN U314 ( .B(n52), .A(n13522), .Z(n26732) );
  NANDN U315 ( .A(n13509), .B(n13510), .Z(n26753) );
  NANDN U316 ( .A(n17822), .B(n17823), .Z(n26783) );
  ANDN U317 ( .B(n13474), .A(n13473), .Z(n26815) );
  ANDN U318 ( .B(n13451), .A(n13450), .Z(n26847) );
  NANDN U319 ( .A(n17959), .B(n17958), .Z(n53) );
  AND U320 ( .A(n17960), .B(n53), .Z(n26856) );
  ANDN U321 ( .B(n13440), .A(n13439), .Z(n26878) );
  ANDN U322 ( .B(n13409), .A(n13408), .Z(n26923) );
  NANDN U323 ( .A(n13400), .B(n13401), .Z(n26935) );
  ANDN U324 ( .B(n13366), .A(n13365), .Z(n26972) );
  ANDN U325 ( .B(n13339), .A(n13338), .Z(n26997) );
  NOR U326 ( .A(n13325), .B(n13326), .Z(n27013) );
  ANDN U327 ( .B(n13319), .A(n13318), .Z(n27033) );
  NANDN U328 ( .A(n13305), .B(n13306), .Z(n27048) );
  NANDN U329 ( .A(n13281), .B(n13282), .Z(n27071) );
  ANDN U330 ( .B(n18367), .A(n18366), .Z(n27087) );
  ANDN U331 ( .B(n13251), .A(n13250), .Z(n27108) );
  ANDN U332 ( .B(n13234), .A(n13233), .Z(n27122) );
  NANDN U333 ( .A(n13217), .B(n13218), .Z(n27147) );
  ANDN U334 ( .B(n13200), .A(n13199), .Z(n27179) );
  ANDN U335 ( .B(n13181), .A(n13180), .Z(n27195) );
  ANDN U336 ( .B(n13164), .A(n13163), .Z(n27211) );
  ANDN U337 ( .B(n18581), .A(n18580), .Z(n27231) );
  ANDN U338 ( .B(n13134), .A(n13133), .Z(n27246) );
  NANDN U339 ( .A(n13117), .B(n13118), .Z(n27258) );
  ANDN U340 ( .B(n13075), .A(n13074), .Z(n27320) );
  NANDN U341 ( .A(n18757), .B(n18756), .Z(n54) );
  ANDN U342 ( .B(n54), .A(n18758), .Z(n27337) );
  ANDN U343 ( .B(n13015), .A(n13014), .Z(n27396) );
  ANDN U344 ( .B(n13005), .A(n13004), .Z(n27409) );
  NOR U345 ( .A(n12975), .B(n12976), .Z(n27441) );
  ANDN U346 ( .B(n12952), .A(n12951), .Z(n27477) );
  AND U347 ( .A(n12939), .B(n12940), .Z(n55) );
  NAND U348 ( .A(n12942), .B(n12941), .Z(n56) );
  AND U349 ( .A(n55), .B(n56), .Z(n27492) );
  NANDN U350 ( .A(y[2218]), .B(x[2218]), .Z(n57) );
  ANDN U351 ( .B(n57), .A(n12873), .Z(n27564) );
  ANDN U352 ( .B(n12859), .A(n12858), .Z(n58) );
  NANDN U353 ( .A(n12861), .B(n12860), .Z(n59) );
  AND U354 ( .A(n58), .B(n59), .Z(n27577) );
  ANDN U355 ( .B(n19237), .A(n19236), .Z(n60) );
  NAND U356 ( .A(n19238), .B(n19239), .Z(n61) );
  AND U357 ( .A(n60), .B(n61), .Z(n24269) );
  ANDN U358 ( .B(n19289), .A(n19288), .Z(n27624) );
  NOR U359 ( .A(n19300), .B(n19301), .Z(n27634) );
  ANDN U360 ( .B(n12757), .A(n12756), .Z(n27714) );
  ANDN U361 ( .B(n19457), .A(n19456), .Z(n27740) );
  ANDN U362 ( .B(n12736), .A(n12735), .Z(n27754) );
  ANDN U363 ( .B(n12698), .A(n12697), .Z(n27815) );
  NANDN U364 ( .A(n12666), .B(n27862), .Z(n27860) );
  NANDN U365 ( .A(n12608), .B(n12609), .Z(n27943) );
  ANDN U366 ( .B(n12585), .A(n12584), .Z(n27972) );
  NANDN U367 ( .A(n12530), .B(n12529), .Z(n62) );
  ANDN U368 ( .B(n62), .A(n12531), .Z(n28050) );
  ANDN U369 ( .B(n12515), .A(n12514), .Z(n28069) );
  NANDN U370 ( .A(x[2708]), .B(y[2708]), .Z(n63) );
  ANDN U371 ( .B(n63), .A(n20167), .Z(n28119) );
  ANDN U372 ( .B(n24176), .A(n12448), .Z(n28150) );
  ANDN U373 ( .B(n12442), .A(n12441), .Z(n28160) );
  ANDN U374 ( .B(n12425), .A(n12424), .Z(n28181) );
  ANDN U375 ( .B(n12411), .A(n12410), .Z(n28204) );
  NANDN U376 ( .A(x[2796]), .B(y[2796]), .Z(n64) );
  ANDN U377 ( .B(n64), .A(n20360), .Z(n28214) );
  NOR U378 ( .A(n20402), .B(n20403), .Z(n28232) );
  NANDN U379 ( .A(x[2858]), .B(y[2858]), .Z(n65) );
  ANDN U380 ( .B(n65), .A(n12355), .Z(n28307) );
  NANDN U381 ( .A(n12310), .B(n12311), .Z(n28357) );
  NAND U382 ( .A(n20810), .B(n20811), .Z(n28462) );
  ANDN U383 ( .B(n12216), .A(n12215), .Z(n28475) );
  NANDN U384 ( .A(n15461), .B(n15462), .Z(n24569) );
  NANDN U385 ( .A(n15417), .B(n15418), .Z(n24613) );
  NANDN U386 ( .A(n15385), .B(n15386), .Z(n24645) );
  NANDN U387 ( .A(n15362), .B(n15363), .Z(n24681) );
  NANDN U388 ( .A(n15318), .B(n15319), .Z(n24729) );
  ANDN U389 ( .B(n15279), .A(n15278), .Z(n24771) );
  ANDN U390 ( .B(n15244), .A(n15243), .Z(n24807) );
  ANDN U391 ( .B(n15202), .A(n15201), .Z(n24855) );
  XNOR U392 ( .A(y[182]), .B(x[182]), .Z(n66) );
  NAND U393 ( .A(n15157), .B(n66), .Z(n24897) );
  ANDN U394 ( .B(n15124), .A(n15123), .Z(n24931) );
  ANDN U395 ( .B(n15080), .A(n15079), .Z(n24975) );
  XNOR U396 ( .A(y[242]), .B(x[242]), .Z(n67) );
  NAND U397 ( .A(n15038), .B(n67), .Z(n25017) );
  ANDN U398 ( .B(n15006), .A(n15005), .Z(n25051) );
  ANDN U399 ( .B(n14980), .A(n14979), .Z(n25091) );
  ANDN U400 ( .B(n14932), .A(n14931), .Z(n25139) );
  ANDN U401 ( .B(n14896), .A(n14895), .Z(n25175) );
  NANDN U402 ( .A(n14858), .B(n14859), .Z(n25221) );
  NANDN U403 ( .A(n14834), .B(n14835), .Z(n25242) );
  NANDN U404 ( .A(n14790), .B(n14791), .Z(n25277) );
  NANDN U405 ( .A(n14742), .B(n14743), .Z(n25345) );
  NANDN U406 ( .A(n14672), .B(n14673), .Z(n25425) );
  NANDN U407 ( .A(n14624), .B(n14625), .Z(n25473) );
  NANDN U408 ( .A(n14579), .B(n14580), .Z(n25517) );
  NANDN U409 ( .A(n14553), .B(n14554), .Z(n25539) );
  NANDN U410 ( .A(n14505), .B(n14506), .Z(n25576) );
  NANDN U411 ( .A(n14465), .B(n14466), .Z(n25616) );
  NANDN U412 ( .A(n14409), .B(n14410), .Z(n25666) );
  NANDN U413 ( .A(n14375), .B(n14376), .Z(n25706) );
  NANDN U414 ( .A(n14331), .B(n14332), .Z(n25750) );
  NANDN U415 ( .A(n14287), .B(n14288), .Z(n25794) );
  NANDN U416 ( .A(n14259), .B(n14260), .Z(n25826) );
  ANDN U417 ( .B(n14221), .A(n14220), .Z(n25862) );
  ANDN U418 ( .B(n14188), .A(n14187), .Z(n25880) );
  ANDN U419 ( .B(n14177), .A(n14176), .Z(n25885) );
  ANDN U420 ( .B(n14120), .A(n14119), .Z(n25914) );
  ANDN U421 ( .B(n14094), .A(n14093), .Z(n25928) );
  NANDN U422 ( .A(n14074), .B(n14075), .Z(n25949) );
  NANDN U423 ( .A(n14030), .B(n14031), .Z(n25987) );
  NANDN U424 ( .A(x[870]), .B(y[870]), .Z(n68) );
  NANDN U425 ( .A(n13985), .B(n68), .Z(n26072) );
  ANDN U426 ( .B(n16531), .A(n16530), .Z(n26088) );
  ANDN U427 ( .B(n13954), .A(n13953), .Z(n26112) );
  NAND U428 ( .A(n13931), .B(n13930), .Z(n69) );
  NAND U429 ( .A(n13932), .B(n69), .Z(n70) );
  AND U430 ( .A(n13933), .B(n70), .Z(n26133) );
  NAND U431 ( .A(n26151), .B(n26150), .Z(n71) );
  NANDN U432 ( .A(n26152), .B(n71), .Z(n72) );
  AND U433 ( .A(n26153), .B(n72), .Z(n73) );
  OR U434 ( .A(n26154), .B(n73), .Z(n74) );
  NAND U435 ( .A(n26155), .B(n74), .Z(n75) );
  NANDN U436 ( .A(n26156), .B(n75), .Z(n76) );
  NAND U437 ( .A(n26157), .B(n76), .Z(n77) );
  NANDN U438 ( .A(n26158), .B(n77), .Z(n78) );
  AND U439 ( .A(n26159), .B(n78), .Z(n79) );
  OR U440 ( .A(n26160), .B(n79), .Z(n80) );
  NAND U441 ( .A(n26161), .B(n80), .Z(n81) );
  NANDN U442 ( .A(n26162), .B(n81), .Z(n82) );
  NAND U443 ( .A(n26163), .B(n82), .Z(n83) );
  NANDN U444 ( .A(n26164), .B(n83), .Z(n84) );
  AND U445 ( .A(n26165), .B(n84), .Z(n85) );
  OR U446 ( .A(n26166), .B(n85), .Z(n86) );
  NAND U447 ( .A(n26167), .B(n86), .Z(n87) );
  NANDN U448 ( .A(n26168), .B(n87), .Z(n88) );
  NANDN U449 ( .A(n26169), .B(n88), .Z(n26170) );
  ANDN U450 ( .B(n13873), .A(n13872), .Z(n26193) );
  ANDN U451 ( .B(n26219), .A(n26218), .Z(n89) );
  NANDN U452 ( .A(n26217), .B(n26216), .Z(n90) );
  NAND U453 ( .A(n89), .B(n90), .Z(n91) );
  NANDN U454 ( .A(n24478), .B(n91), .Z(n92) );
  NAND U455 ( .A(n24477), .B(n92), .Z(n93) );
  AND U456 ( .A(n26220), .B(n93), .Z(n94) );
  OR U457 ( .A(n24476), .B(n94), .Z(n95) );
  NAND U458 ( .A(n26221), .B(n95), .Z(n96) );
  NANDN U459 ( .A(n24475), .B(n96), .Z(n97) );
  NAND U460 ( .A(n26222), .B(n97), .Z(n98) );
  NANDN U461 ( .A(n26223), .B(n98), .Z(n99) );
  AND U462 ( .A(n26224), .B(n99), .Z(n100) );
  OR U463 ( .A(n26225), .B(n100), .Z(n101) );
  NAND U464 ( .A(n26226), .B(n101), .Z(n102) );
  NAND U465 ( .A(n26227), .B(n102), .Z(n103) );
  AND U466 ( .A(n26228), .B(n103), .Z(n26231) );
  ANDN U467 ( .B(n13828), .A(n13827), .Z(n26254) );
  NAND U468 ( .A(n26276), .B(n26275), .Z(n104) );
  NAND U469 ( .A(n26277), .B(n104), .Z(n105) );
  ANDN U470 ( .B(n105), .A(n24466), .Z(n106) );
  OR U471 ( .A(n26278), .B(n106), .Z(n107) );
  NAND U472 ( .A(n26279), .B(n107), .Z(n108) );
  NANDN U473 ( .A(n26280), .B(n108), .Z(n109) );
  NAND U474 ( .A(n26281), .B(n109), .Z(n110) );
  NANDN U475 ( .A(n26282), .B(n110), .Z(n111) );
  AND U476 ( .A(n26283), .B(n111), .Z(n112) );
  OR U477 ( .A(n24465), .B(n112), .Z(n113) );
  NANDN U478 ( .A(n26284), .B(n113), .Z(n114) );
  NAND U479 ( .A(n26285), .B(n114), .Z(n115) );
  AND U480 ( .A(n24463), .B(n24464), .Z(n116) );
  NAND U481 ( .A(n115), .B(n116), .Z(n117) );
  NANDN U482 ( .A(n26286), .B(n117), .Z(n118) );
  NAND U483 ( .A(n26287), .B(n118), .Z(n119) );
  NANDN U484 ( .A(n26288), .B(n119), .Z(n120) );
  AND U485 ( .A(n26289), .B(n120), .Z(n26290) );
  NOR U486 ( .A(n16996), .B(n16997), .Z(n26328) );
  NAND U487 ( .A(n13745), .B(n13744), .Z(n121) );
  AND U488 ( .A(n13746), .B(n121), .Z(n24449) );
  ANDN U489 ( .B(n13721), .A(n13720), .Z(n26373) );
  NAND U490 ( .A(n13709), .B(n13710), .Z(n122) );
  ANDN U491 ( .B(n122), .A(n13711), .Z(n26385) );
  NOR U492 ( .A(n13700), .B(n13701), .Z(n24440) );
  NANDN U493 ( .A(n13679), .B(n13680), .Z(n26459) );
  NANDN U494 ( .A(n17262), .B(n17263), .Z(n26474) );
  ANDN U495 ( .B(n13656), .A(n13655), .Z(n26492) );
  ANDN U496 ( .B(n13638), .A(n13637), .Z(n26513) );
  NANDN U497 ( .A(n13616), .B(n13617), .Z(n26534) );
  ANDN U498 ( .B(n17552), .A(n13574), .Z(n123) );
  NANDN U499 ( .A(n13576), .B(n13575), .Z(n124) );
  AND U500 ( .A(n123), .B(n124), .Z(n26603) );
  NANDN U501 ( .A(n13537), .B(n13536), .Z(n125) );
  AND U502 ( .A(n13538), .B(n125), .Z(n26705) );
  NANDN U503 ( .A(n26730), .B(n26729), .Z(n126) );
  NAND U504 ( .A(n26731), .B(n126), .Z(n127) );
  AND U505 ( .A(n26732), .B(n127), .Z(n128) );
  NANDN U506 ( .A(n128), .B(n26733), .Z(n129) );
  NANDN U507 ( .A(n26734), .B(n129), .Z(n130) );
  NANDN U508 ( .A(n26735), .B(n130), .Z(n131) );
  NANDN U509 ( .A(n26736), .B(n131), .Z(n132) );
  NAND U510 ( .A(n26737), .B(n132), .Z(n133) );
  AND U511 ( .A(n26738), .B(n133), .Z(n134) );
  NANDN U512 ( .A(n134), .B(n26739), .Z(n135) );
  NANDN U513 ( .A(n26740), .B(n135), .Z(n136) );
  NAND U514 ( .A(n26741), .B(n136), .Z(n137) );
  NANDN U515 ( .A(n24400), .B(n137), .Z(n138) );
  NANDN U516 ( .A(n26742), .B(n138), .Z(n139) );
  AND U517 ( .A(n26743), .B(n139), .Z(n140) );
  NANDN U518 ( .A(n140), .B(n26744), .Z(n141) );
  NAND U519 ( .A(n26745), .B(n141), .Z(n142) );
  NANDN U520 ( .A(n26746), .B(n142), .Z(n143) );
  NAND U521 ( .A(n26747), .B(n143), .Z(n26748) );
  NANDN U522 ( .A(n13492), .B(n13493), .Z(n26781) );
  NAND U523 ( .A(n26822), .B(n24386), .Z(n144) );
  NAND U524 ( .A(n26823), .B(n144), .Z(n145) );
  AND U525 ( .A(n24385), .B(n145), .Z(n146) );
  NANDN U526 ( .A(n146), .B(n26824), .Z(n147) );
  NAND U527 ( .A(n26825), .B(n147), .Z(n148) );
  NAND U528 ( .A(n26826), .B(n148), .Z(n149) );
  NAND U529 ( .A(n24384), .B(n149), .Z(n150) );
  NAND U530 ( .A(n26827), .B(n150), .Z(n151) );
  ANDN U531 ( .B(n151), .A(n26828), .Z(n152) );
  NANDN U532 ( .A(n152), .B(n26829), .Z(n153) );
  NANDN U533 ( .A(n26830), .B(n153), .Z(n154) );
  NANDN U534 ( .A(n26831), .B(n154), .Z(n155) );
  NAND U535 ( .A(n26832), .B(n155), .Z(n156) );
  AND U536 ( .A(n26834), .B(n156), .Z(n157) );
  NANDN U537 ( .A(n26833), .B(n157), .Z(n158) );
  AND U538 ( .A(n26835), .B(n158), .Z(n26836) );
  NANDN U539 ( .A(n17965), .B(n17966), .Z(n159) );
  ANDN U540 ( .B(n159), .A(n17967), .Z(n26860) );
  ANDN U541 ( .B(n13438), .A(n13437), .Z(n26879) );
  ANDN U542 ( .B(n13405), .A(n13404), .Z(n26925) );
  ANDN U543 ( .B(n13399), .A(n13398), .Z(n26936) );
  ANDN U544 ( .B(n13383), .A(n13382), .Z(n26950) );
  NANDN U545 ( .A(n13363), .B(n13364), .Z(n26973) );
  ANDN U546 ( .B(n13351), .A(n13350), .Z(n26984) );
  ANDN U547 ( .B(n13330), .A(n13329), .Z(n27006) );
  ANDN U548 ( .B(n13322), .A(n13321), .Z(n27018) );
  ANDN U549 ( .B(n18283), .A(n18282), .Z(n27034) );
  NANDN U550 ( .A(n13301), .B(n13302), .Z(n27050) );
  NANDN U551 ( .A(n13277), .B(n13278), .Z(n27073) );
  NANDN U552 ( .A(n13263), .B(n13264), .Z(n27088) );
  ANDN U553 ( .B(n13249), .A(n13248), .Z(n27110) );
  NANDN U554 ( .A(n13231), .B(n13232), .Z(n27123) );
  ANDN U555 ( .B(n13216), .A(n13215), .Z(n27149) );
  NANDN U556 ( .A(n13197), .B(n13198), .Z(n27180) );
  NANDN U557 ( .A(n13178), .B(n13179), .Z(n27196) );
  NANDN U558 ( .A(n13161), .B(n13162), .Z(n27212) );
  ANDN U559 ( .B(n13146), .A(n13145), .Z(n27232) );
  ANDN U560 ( .B(n13132), .A(n13131), .Z(n27247) );
  ANDN U561 ( .B(n13116), .A(n13115), .Z(n27259) );
  NAND U562 ( .A(n18675), .B(n18676), .Z(n160) );
  ANDN U563 ( .B(n160), .A(n18677), .Z(n27288) );
  ANDN U564 ( .B(n13093), .A(n13092), .Z(n27300) );
  NANDN U565 ( .A(n13072), .B(n13073), .Z(n27321) );
  ANDN U566 ( .B(n13061), .A(n13060), .Z(n27341) );
  NANDN U567 ( .A(n13047), .B(n13048), .Z(n27351) );
  ANDN U568 ( .B(n13027), .A(n13026), .Z(n27376) );
  ANDN U569 ( .B(n27403), .A(n13010), .Z(n27399) );
  NANDN U570 ( .A(n12999), .B(n12998), .Z(n161) );
  ANDN U571 ( .B(n161), .A(n13000), .Z(n27417) );
  ANDN U572 ( .B(n12987), .A(n12986), .Z(n27431) );
  NOR U573 ( .A(n18944), .B(n18945), .Z(n27443) );
  ANDN U574 ( .B(n12958), .A(n12957), .Z(n27470) );
  NOR U575 ( .A(n12934), .B(n12935), .Z(n27494) );
  ANDN U576 ( .B(n12923), .A(n12922), .Z(n27514) );
  AND U577 ( .A(n27554), .B(n27553), .Z(n162) );
  NAND U578 ( .A(n27556), .B(n27555), .Z(n163) );
  AND U579 ( .A(n162), .B(n163), .Z(n164) );
  NANDN U580 ( .A(n164), .B(n27557), .Z(n165) );
  NAND U581 ( .A(n27558), .B(n165), .Z(n166) );
  NAND U582 ( .A(n27559), .B(n166), .Z(n167) );
  NAND U583 ( .A(n27560), .B(n167), .Z(n168) );
  NANDN U584 ( .A(n27561), .B(n168), .Z(n169) );
  AND U585 ( .A(n27562), .B(n169), .Z(n170) );
  NANDN U586 ( .A(n170), .B(n27563), .Z(n171) );
  NAND U587 ( .A(n27564), .B(n171), .Z(n172) );
  NAND U588 ( .A(n24274), .B(n172), .Z(n173) );
  NAND U589 ( .A(n27565), .B(n173), .Z(n174) );
  NAND U590 ( .A(n27566), .B(n174), .Z(n175) );
  AND U591 ( .A(n27567), .B(n175), .Z(n176) );
  NANDN U592 ( .A(n176), .B(n27568), .Z(n177) );
  ANDN U593 ( .B(n177), .A(n27569), .Z(n27572) );
  NAND U594 ( .A(n12839), .B(n19237), .Z(n178) );
  AND U595 ( .A(n12840), .B(n178), .Z(n27597) );
  ANDN U596 ( .B(n12816), .A(n12815), .Z(n27625) );
  ANDN U597 ( .B(n12801), .A(n12800), .Z(n27646) );
  NANDN U598 ( .A(n12754), .B(n12755), .Z(n27716) );
  XNOR U599 ( .A(x[2362]), .B(y[2362]), .Z(n179) );
  NAND U600 ( .A(n27735), .B(n179), .Z(n180) );
  ANDN U601 ( .B(n180), .A(n24255), .Z(n181) );
  NANDN U602 ( .A(y[2362]), .B(x[2362]), .Z(n182) );
  AND U603 ( .A(n181), .B(n182), .Z(n183) );
  OR U604 ( .A(n183), .B(n27736), .Z(n184) );
  NAND U605 ( .A(n27737), .B(n184), .Z(n185) );
  NANDN U606 ( .A(n27738), .B(n185), .Z(n186) );
  NAND U607 ( .A(n27739), .B(n186), .Z(n187) );
  NAND U608 ( .A(n27740), .B(n187), .Z(n188) );
  AND U609 ( .A(n27741), .B(n188), .Z(n189) );
  NANDN U610 ( .A(n189), .B(n27742), .Z(n190) );
  NAND U611 ( .A(n24254), .B(n190), .Z(n191) );
  NANDN U612 ( .A(n24253), .B(n191), .Z(n192) );
  NAND U613 ( .A(n27743), .B(n192), .Z(n27744) );
  NAND U614 ( .A(n12693), .B(n12692), .Z(n193) );
  AND U615 ( .A(n12694), .B(n193), .Z(n24243) );
  ANDN U616 ( .B(n12684), .A(n12683), .Z(n27833) );
  NANDN U617 ( .A(n12662), .B(n12663), .Z(n27865) );
  ANDN U618 ( .B(n12638), .A(n12637), .Z(n27912) );
  NANDN U619 ( .A(n12598), .B(n12599), .Z(n27959) );
  ANDN U620 ( .B(n12581), .A(n12580), .Z(n27974) );
  ANDN U621 ( .B(n12541), .A(n24203), .Z(n28036) );
  NAND U622 ( .A(n28038), .B(n28039), .Z(n28040) );
  NANDN U623 ( .A(n12527), .B(n12528), .Z(n28055) );
  ANDN U624 ( .B(n12498), .A(n12497), .Z(n28094) );
  NANDN U625 ( .A(n12478), .B(n12479), .Z(n28111) );
  NANDN U626 ( .A(n20171), .B(n20172), .Z(n28120) );
  NANDN U627 ( .A(x[2742]), .B(y[2742]), .Z(n194) );
  ANDN U628 ( .B(n194), .A(n12445), .Z(n28157) );
  ANDN U629 ( .B(n12439), .A(n12438), .Z(n28167) );
  ANDN U630 ( .B(n24163), .A(n20354), .Z(n28209) );
  ANDN U631 ( .B(n12402), .A(n12401), .Z(n24159) );
  ANDN U632 ( .B(n12393), .A(n12392), .Z(n28233) );
  ANDN U633 ( .B(n20436), .A(n20435), .Z(n28252) );
  ANDN U634 ( .B(n12376), .A(n12375), .Z(n28265) );
  ANDN U635 ( .B(n12352), .A(n12351), .Z(n28309) );
  ANDN U636 ( .B(n12333), .A(n12332), .Z(n28331) );
  ANDN U637 ( .B(n12308), .A(n12307), .Z(n28365) );
  NANDN U638 ( .A(n12254), .B(n12255), .Z(n28433) );
  ANDN U639 ( .B(n12222), .A(n12221), .Z(n28470) );
  ANDN U640 ( .B(n20834), .A(n20833), .Z(n28477) );
  ANDN U641 ( .B(n12174), .A(n12173), .Z(n24097) );
  ANDN U642 ( .B(n12165), .A(n12164), .Z(n28545) );
  NANDN U643 ( .A(n15457), .B(n15458), .Z(n24573) );
  NANDN U644 ( .A(n15413), .B(n15414), .Z(n24617) );
  NANDN U645 ( .A(n15381), .B(n15382), .Z(n24649) );
  NANDN U646 ( .A(n15358), .B(n15359), .Z(n24685) );
  NANDN U647 ( .A(y[100]), .B(x[100]), .Z(n195) );
  NANDN U648 ( .A(n15315), .B(n195), .Z(n24733) );
  ANDN U649 ( .B(n15275), .A(n15274), .Z(n24775) );
  ANDN U650 ( .B(n15240), .A(n15239), .Z(n24811) );
  ANDN U651 ( .B(n15198), .A(n15197), .Z(n24859) );
  ANDN U652 ( .B(n15156), .A(n15155), .Z(n24899) );
  ANDN U653 ( .B(n15120), .A(n15119), .Z(n24935) );
  ANDN U654 ( .B(n15076), .A(n15075), .Z(n24979) );
  ANDN U655 ( .B(n15037), .A(n15036), .Z(n25019) );
  XNOR U656 ( .A(x[260]), .B(y[260]), .Z(n196) );
  NAND U657 ( .A(n15004), .B(n196), .Z(n25053) );
  ANDN U658 ( .B(n14958), .A(n14957), .Z(n25111) );
  ANDN U659 ( .B(n14919), .A(n14918), .Z(n25151) );
  ANDN U660 ( .B(n14885), .A(n14884), .Z(n25187) );
  NANDN U661 ( .A(n14850), .B(n14851), .Z(n25229) );
  NANDN U662 ( .A(n14818), .B(n14819), .Z(n25250) );
  NANDN U663 ( .A(n14778), .B(n14779), .Z(n25289) );
  NANDN U664 ( .A(n14734), .B(n14735), .Z(n25353) );
  NANDN U665 ( .A(n14708), .B(n14709), .Z(n25389) );
  NANDN U666 ( .A(n14664), .B(n14665), .Z(n25433) );
  NANDN U667 ( .A(n14620), .B(n14621), .Z(n25477) );
  NANDN U668 ( .A(n14575), .B(n14576), .Z(n25521) );
  NANDN U669 ( .A(n14549), .B(n14550), .Z(n25541) );
  NANDN U670 ( .A(n14501), .B(n14502), .Z(n25580) );
  NANDN U671 ( .A(n14457), .B(n14458), .Z(n25624) );
  NANDN U672 ( .A(n14403), .B(n14404), .Z(n25678) );
  NANDN U673 ( .A(n14363), .B(n14364), .Z(n25718) );
  NANDN U674 ( .A(n14327), .B(n14328), .Z(n25754) );
  NANDN U675 ( .A(n14283), .B(n14284), .Z(n25798) );
  NANDN U676 ( .A(n14251), .B(n14252), .Z(n25834) );
  ANDN U677 ( .B(n14234), .A(n14233), .Z(n25851) );
  NAND U678 ( .A(n25874), .B(n25873), .Z(n197) );
  NAND U679 ( .A(n25875), .B(n197), .Z(n198) );
  NAND U680 ( .A(n25876), .B(n198), .Z(n199) );
  NAND U681 ( .A(n25877), .B(n199), .Z(n200) );
  NAND U682 ( .A(n24529), .B(n200), .Z(n201) );
  AND U683 ( .A(n25878), .B(n201), .Z(n202) );
  NANDN U684 ( .A(n202), .B(n25879), .Z(n203) );
  NAND U685 ( .A(n25880), .B(n203), .Z(n204) );
  NAND U686 ( .A(n25881), .B(n204), .Z(n205) );
  NAND U687 ( .A(n25882), .B(n205), .Z(n206) );
  NAND U688 ( .A(n24528), .B(n206), .Z(n207) );
  AND U689 ( .A(n25883), .B(n207), .Z(n208) );
  NANDN U690 ( .A(n208), .B(n24527), .Z(n209) );
  ANDN U691 ( .B(n209), .A(n25884), .Z(n25886) );
  OR U692 ( .A(n25910), .B(n25911), .Z(n210) );
  NAND U693 ( .A(n25912), .B(n210), .Z(n211) );
  NAND U694 ( .A(n25913), .B(n211), .Z(n212) );
  NANDN U695 ( .A(n24518), .B(n212), .Z(n213) );
  NAND U696 ( .A(n25914), .B(n213), .Z(n214) );
  ANDN U697 ( .B(n214), .A(n25915), .Z(n215) );
  NANDN U698 ( .A(n215), .B(n25916), .Z(n216) );
  NAND U699 ( .A(n25917), .B(n216), .Z(n217) );
  NAND U700 ( .A(n24517), .B(n217), .Z(n218) );
  NAND U701 ( .A(n25918), .B(n218), .Z(n219) );
  NAND U702 ( .A(n25919), .B(n219), .Z(n220) );
  AND U703 ( .A(n25920), .B(n220), .Z(n221) );
  NANDN U704 ( .A(n221), .B(n25921), .Z(n222) );
  NANDN U705 ( .A(n24516), .B(n222), .Z(n223) );
  NAND U706 ( .A(n25922), .B(n223), .Z(n224) );
  NAND U707 ( .A(n25923), .B(n224), .Z(n25924) );
  ANDN U708 ( .B(n14073), .A(n14072), .Z(n25950) );
  ANDN U709 ( .B(n14029), .A(n14028), .Z(n25989) );
  ANDN U710 ( .B(n14011), .A(n14010), .Z(n26041) );
  NANDN U711 ( .A(n14002), .B(n14003), .Z(n26052) );
  NOR U712 ( .A(n16499), .B(n16500), .Z(n26077) );
  ANDN U713 ( .B(n13976), .A(n13975), .Z(n26089) );
  NANDN U714 ( .A(n26109), .B(n26108), .Z(n225) );
  NAND U715 ( .A(n26110), .B(n225), .Z(n226) );
  AND U716 ( .A(n26111), .B(n226), .Z(n227) );
  NANDN U717 ( .A(n227), .B(n26112), .Z(n228) );
  NANDN U718 ( .A(n26113), .B(n228), .Z(n229) );
  NAND U719 ( .A(n26114), .B(n229), .Z(n230) );
  NANDN U720 ( .A(n26115), .B(n230), .Z(n231) );
  NAND U721 ( .A(n26116), .B(n231), .Z(n232) );
  ANDN U722 ( .B(n232), .A(n26117), .Z(n233) );
  NANDN U723 ( .A(n233), .B(n26118), .Z(n234) );
  NANDN U724 ( .A(n24495), .B(n234), .Z(n235) );
  NAND U725 ( .A(n24494), .B(n235), .Z(n236) );
  NANDN U726 ( .A(n24493), .B(n236), .Z(n237) );
  NAND U727 ( .A(n24492), .B(n237), .Z(n238) );
  ANDN U728 ( .B(n238), .A(n26119), .Z(n26121) );
  NANDN U729 ( .A(n13928), .B(n13929), .Z(n26139) );
  NAND U730 ( .A(n26171), .B(n26170), .Z(n239) );
  NANDN U731 ( .A(n26172), .B(n239), .Z(n240) );
  AND U732 ( .A(n26173), .B(n240), .Z(n241) );
  OR U733 ( .A(n26174), .B(n241), .Z(n242) );
  NAND U734 ( .A(n26175), .B(n242), .Z(n243) );
  NANDN U735 ( .A(n26176), .B(n243), .Z(n244) );
  NAND U736 ( .A(n26177), .B(n244), .Z(n245) );
  NANDN U737 ( .A(n26178), .B(n245), .Z(n246) );
  AND U738 ( .A(n26179), .B(n246), .Z(n247) );
  OR U739 ( .A(n26180), .B(n247), .Z(n248) );
  NAND U740 ( .A(n26181), .B(n248), .Z(n249) );
  NAND U741 ( .A(n24485), .B(n249), .Z(n250) );
  NAND U742 ( .A(n26182), .B(n250), .Z(n251) );
  NAND U743 ( .A(n26183), .B(n251), .Z(n252) );
  AND U744 ( .A(n26184), .B(n252), .Z(n253) );
  NANDN U745 ( .A(n253), .B(n26185), .Z(n254) );
  NAND U746 ( .A(n26186), .B(n254), .Z(n255) );
  NAND U747 ( .A(n24484), .B(n255), .Z(n26189) );
  NANDN U748 ( .A(n13859), .B(n13860), .Z(n26213) );
  NANDN U749 ( .A(n26231), .B(n26230), .Z(n256) );
  NAND U750 ( .A(n26232), .B(n256), .Z(n257) );
  NANDN U751 ( .A(n26233), .B(n257), .Z(n258) );
  NAND U752 ( .A(n26234), .B(n258), .Z(n259) );
  NAND U753 ( .A(n26235), .B(n259), .Z(n260) );
  AND U754 ( .A(n26236), .B(n260), .Z(n261) );
  OR U755 ( .A(n26237), .B(n261), .Z(n262) );
  NAND U756 ( .A(n26238), .B(n262), .Z(n263) );
  NANDN U757 ( .A(n26239), .B(n263), .Z(n264) );
  NAND U758 ( .A(n26240), .B(n264), .Z(n265) );
  NANDN U759 ( .A(n24474), .B(n265), .Z(n266) );
  AND U760 ( .A(n24473), .B(n266), .Z(n267) );
  NANDN U761 ( .A(n267), .B(n26241), .Z(n268) );
  ANDN U762 ( .B(n268), .A(n26242), .Z(n269) );
  NANDN U763 ( .A(n269), .B(n26243), .Z(n270) );
  NAND U764 ( .A(n26244), .B(n270), .Z(n271) );
  NAND U765 ( .A(n26245), .B(n271), .Z(n26246) );
  NAND U766 ( .A(n13816), .B(n13817), .Z(n272) );
  ANDN U767 ( .B(n272), .A(n13818), .Z(n26271) );
  NAND U768 ( .A(n26290), .B(n24462), .Z(n273) );
  NAND U769 ( .A(n26291), .B(n273), .Z(n274) );
  NAND U770 ( .A(n24461), .B(n274), .Z(n275) );
  NAND U771 ( .A(n26292), .B(n275), .Z(n276) );
  NAND U772 ( .A(n26293), .B(n276), .Z(n277) );
  AND U773 ( .A(n26294), .B(n277), .Z(n278) );
  NANDN U774 ( .A(n278), .B(n26295), .Z(n279) );
  NANDN U775 ( .A(n26296), .B(n279), .Z(n280) );
  NAND U776 ( .A(n26297), .B(n280), .Z(n281) );
  NANDN U777 ( .A(n26298), .B(n281), .Z(n282) );
  NAND U778 ( .A(n26299), .B(n282), .Z(n283) );
  AND U779 ( .A(n26300), .B(n283), .Z(n284) );
  NANDN U780 ( .A(n284), .B(n24460), .Z(n285) );
  NANDN U781 ( .A(n26301), .B(n285), .Z(n286) );
  NAND U782 ( .A(n26302), .B(n286), .Z(n26305) );
  NANDN U783 ( .A(n13768), .B(n13763), .Z(n287) );
  ANDN U784 ( .B(n287), .A(n13764), .Z(n26321) );
  NANDN U785 ( .A(n24449), .B(n26342), .Z(n288) );
  NAND U786 ( .A(n24448), .B(n288), .Z(n289) );
  ANDN U787 ( .B(n289), .A(n26343), .Z(n290) );
  NAND U788 ( .A(n290), .B(n26344), .Z(n291) );
  NAND U789 ( .A(n26345), .B(n291), .Z(n292) );
  ANDN U790 ( .B(n292), .A(n26346), .Z(n293) );
  OR U791 ( .A(n26347), .B(n293), .Z(n294) );
  NANDN U792 ( .A(n26348), .B(n294), .Z(n295) );
  NAND U793 ( .A(n26349), .B(n295), .Z(n296) );
  NANDN U794 ( .A(n24447), .B(n296), .Z(n297) );
  NAND U795 ( .A(n26350), .B(n297), .Z(n298) );
  ANDN U796 ( .B(n298), .A(n26351), .Z(n299) );
  OR U797 ( .A(n26352), .B(n299), .Z(n300) );
  NAND U798 ( .A(n26353), .B(n300), .Z(n301) );
  NAND U799 ( .A(n26354), .B(n301), .Z(n26357) );
  NOR U800 ( .A(n13714), .B(n13715), .Z(n26375) );
  NANDN U801 ( .A(n13696), .B(n13697), .Z(n26402) );
  NOR U802 ( .A(n13675), .B(n13676), .Z(n26462) );
  NAND U803 ( .A(n26503), .B(n26504), .Z(n302) );
  NANDN U804 ( .A(n26505), .B(n302), .Z(n303) );
  NAND U805 ( .A(n26506), .B(n303), .Z(n304) );
  NANDN U806 ( .A(n24425), .B(n304), .Z(n305) );
  NAND U807 ( .A(n26507), .B(n305), .Z(n306) );
  ANDN U808 ( .B(n306), .A(n24424), .Z(n307) );
  OR U809 ( .A(n26508), .B(n307), .Z(n308) );
  NANDN U810 ( .A(n26509), .B(n308), .Z(n309) );
  NANDN U811 ( .A(n26510), .B(n309), .Z(n310) );
  NAND U812 ( .A(n26511), .B(n310), .Z(n311) );
  NANDN U813 ( .A(n26512), .B(n311), .Z(n312) );
  AND U814 ( .A(n26513), .B(n312), .Z(n313) );
  NANDN U815 ( .A(n313), .B(n26514), .Z(n314) );
  NAND U816 ( .A(n24423), .B(n314), .Z(n315) );
  NAND U817 ( .A(n26515), .B(n315), .Z(n316) );
  NAND U818 ( .A(n26516), .B(n316), .Z(n26519) );
  NANDN U819 ( .A(n13611), .B(n13612), .Z(n317) );
  NAND U820 ( .A(n13610), .B(n317), .Z(n318) );
  ANDN U821 ( .B(n318), .A(n13613), .Z(n26539) );
  NANDN U822 ( .A(x[1331]), .B(y[1331]), .Z(n319) );
  ANDN U823 ( .B(n319), .A(n13606), .Z(n26551) );
  NOR U824 ( .A(n17521), .B(n17522), .Z(n26588) );
  ANDN U825 ( .B(n13567), .A(n13566), .Z(n26635) );
  NANDN U826 ( .A(n13564), .B(n13565), .Z(n26647) );
  NANDN U827 ( .A(n26679), .B(n26680), .Z(n320) );
  NANDN U828 ( .A(n26681), .B(n320), .Z(n321) );
  NAND U829 ( .A(n26682), .B(n321), .Z(n322) );
  NAND U830 ( .A(n24404), .B(n322), .Z(n323) );
  NANDN U831 ( .A(n26683), .B(n323), .Z(n324) );
  AND U832 ( .A(n26684), .B(n324), .Z(n325) );
  OR U833 ( .A(n26685), .B(n325), .Z(n326) );
  NAND U834 ( .A(n26686), .B(n326), .Z(n327) );
  NANDN U835 ( .A(n26687), .B(n327), .Z(n328) );
  NAND U836 ( .A(n26688), .B(n328), .Z(n329) );
  NANDN U837 ( .A(n26689), .B(n329), .Z(n330) );
  AND U838 ( .A(n26690), .B(n330), .Z(n331) );
  NANDN U839 ( .A(n331), .B(n26691), .Z(n332) );
  NAND U840 ( .A(n26692), .B(n332), .Z(n333) );
  NANDN U841 ( .A(n26693), .B(n333), .Z(n334) );
  NAND U842 ( .A(n26694), .B(n334), .Z(n26695) );
  ANDN U843 ( .B(n13530), .A(n13529), .Z(n26719) );
  NANDN U844 ( .A(n17739), .B(n17740), .Z(n26734) );
  NAND U845 ( .A(n26765), .B(n26766), .Z(n335) );
  NANDN U846 ( .A(n26767), .B(n335), .Z(n336) );
  NAND U847 ( .A(n26768), .B(n336), .Z(n337) );
  ANDN U848 ( .B(n337), .A(n24397), .Z(n338) );
  NANDN U849 ( .A(n26770), .B(n26769), .Z(n339) );
  AND U850 ( .A(n338), .B(n339), .Z(n340) );
  NANDN U851 ( .A(n340), .B(n24396), .Z(n341) );
  NANDN U852 ( .A(n26771), .B(n341), .Z(n342) );
  NAND U853 ( .A(n26772), .B(n342), .Z(n343) );
  NANDN U854 ( .A(n26773), .B(n343), .Z(n344) );
  NAND U855 ( .A(n26774), .B(n344), .Z(n345) );
  ANDN U856 ( .B(n345), .A(n26775), .Z(n346) );
  OR U857 ( .A(n24395), .B(n346), .Z(n347) );
  ANDN U858 ( .B(n347), .A(n26776), .Z(n348) );
  NANDN U859 ( .A(n348), .B(n26777), .Z(n349) );
  NANDN U860 ( .A(n26778), .B(n349), .Z(n350) );
  NAND U861 ( .A(n26779), .B(n350), .Z(n26780) );
  NANDN U862 ( .A(n13485), .B(n13486), .Z(n26799) );
  NOR U863 ( .A(n13470), .B(n13471), .Z(n26821) );
  NAND U864 ( .A(n26853), .B(n26854), .Z(n351) );
  NANDN U865 ( .A(n26855), .B(n351), .Z(n352) );
  NAND U866 ( .A(n26856), .B(n352), .Z(n353) );
  NAND U867 ( .A(n26857), .B(n353), .Z(n354) );
  NANDN U868 ( .A(n26858), .B(n354), .Z(n355) );
  AND U869 ( .A(n26859), .B(n355), .Z(n356) );
  NANDN U870 ( .A(n356), .B(n26860), .Z(n357) );
  NAND U871 ( .A(n26861), .B(n357), .Z(n358) );
  NAND U872 ( .A(n26862), .B(n358), .Z(n359) );
  NAND U873 ( .A(n26863), .B(n359), .Z(n360) );
  NANDN U874 ( .A(n24381), .B(n360), .Z(n361) );
  AND U875 ( .A(n26864), .B(n361), .Z(n362) );
  OR U876 ( .A(n362), .B(n26865), .Z(n363) );
  NANDN U877 ( .A(n26866), .B(n363), .Z(n364) );
  AND U878 ( .A(n26867), .B(n364), .Z(n365) );
  OR U879 ( .A(n26868), .B(n365), .Z(n366) );
  AND U880 ( .A(n26869), .B(n366), .Z(n26871) );
  NANDN U881 ( .A(n13427), .B(n13428), .Z(n26897) );
  ANDN U882 ( .B(n18070), .A(n18069), .Z(n26904) );
  ANDN U883 ( .B(n13423), .A(n13422), .Z(n26911) );
  NANDN U884 ( .A(x[1672]), .B(y[1672]), .Z(n367) );
  ANDN U885 ( .B(n367), .A(n13395), .Z(n26938) );
  ANDN U886 ( .B(n13376), .A(n13375), .Z(n26957) );
  NANDN U887 ( .A(n13359), .B(n13360), .Z(n26975) );
  ANDN U888 ( .B(n13347), .A(n13346), .Z(n26986) );
  ANDN U889 ( .B(n18238), .A(n18237), .Z(n27008) );
  ANDN U890 ( .B(n13315), .A(n13314), .Z(n27035) );
  ANDN U891 ( .B(n13295), .A(n13294), .Z(n27058) );
  NANDN U892 ( .A(n13273), .B(n13274), .Z(n27075) );
  ANDN U893 ( .B(n13262), .A(n13261), .Z(n27089) );
  ANDN U894 ( .B(n13258), .A(n13257), .Z(n27100) );
  ANDN U895 ( .B(n13228), .A(n13227), .Z(n27124) );
  ANDN U896 ( .B(n13214), .A(n13213), .Z(n27150) );
  OR U897 ( .A(n27187), .B(n27188), .Z(n368) );
  NANDN U898 ( .A(n27189), .B(n368), .Z(n369) );
  AND U899 ( .A(n27190), .B(n369), .Z(n370) );
  NANDN U900 ( .A(n370), .B(n27191), .Z(n371) );
  NAND U901 ( .A(n27192), .B(n371), .Z(n372) );
  NAND U902 ( .A(n27193), .B(n372), .Z(n373) );
  NAND U903 ( .A(n27194), .B(n373), .Z(n374) );
  NAND U904 ( .A(n27195), .B(n374), .Z(n375) );
  ANDN U905 ( .B(n375), .A(n27196), .Z(n376) );
  NANDN U906 ( .A(n376), .B(n27197), .Z(n377) );
  NAND U907 ( .A(n27198), .B(n377), .Z(n378) );
  NAND U908 ( .A(n27199), .B(n378), .Z(n379) );
  NAND U909 ( .A(n27200), .B(n379), .Z(n380) );
  NAND U910 ( .A(n27201), .B(n380), .Z(n381) );
  AND U911 ( .A(n27202), .B(n381), .Z(n382) );
  OR U912 ( .A(n27203), .B(n382), .Z(n383) );
  AND U913 ( .A(n27204), .B(n383), .Z(n27206) );
  ANDN U914 ( .B(n13144), .A(n13143), .Z(n27233) );
  ANDN U915 ( .B(n13112), .A(n13111), .Z(n27261) );
  OR U916 ( .A(n13108), .B(n13109), .Z(n384) );
  NAND U917 ( .A(n13110), .B(n384), .Z(n385) );
  NAND U918 ( .A(n13107), .B(n385), .Z(n27269) );
  NAND U919 ( .A(n13097), .B(n13098), .Z(n386) );
  ANDN U920 ( .B(n386), .A(n13099), .Z(n27290) );
  ANDN U921 ( .B(n13089), .A(n13088), .Z(n27302) );
  NANDN U922 ( .A(n13070), .B(n24318), .Z(n27323) );
  NANDN U923 ( .A(n27325), .B(n27324), .Z(n387) );
  ANDN U924 ( .B(n387), .A(n27326), .Z(n27327) );
  ANDN U925 ( .B(n13057), .A(n13056), .Z(n27344) );
  ANDN U926 ( .B(n13031), .A(n13030), .Z(n27370) );
  NAND U927 ( .A(n27387), .B(n27388), .Z(n388) );
  NANDN U928 ( .A(n27389), .B(n388), .Z(n389) );
  NANDN U929 ( .A(n27390), .B(n389), .Z(n390) );
  NAND U930 ( .A(n27391), .B(n390), .Z(n391) );
  NANDN U931 ( .A(n27392), .B(n391), .Z(n392) );
  AND U932 ( .A(n27393), .B(n392), .Z(n393) );
  OR U933 ( .A(n24310), .B(n393), .Z(n394) );
  NAND U934 ( .A(n24308), .B(n24309), .Z(n395) );
  AND U935 ( .A(n394), .B(n395), .Z(n396) );
  NAND U936 ( .A(n396), .B(n27394), .Z(n397) );
  NANDN U937 ( .A(n27395), .B(n397), .Z(n398) );
  AND U938 ( .A(n27396), .B(n398), .Z(n399) );
  OR U939 ( .A(n24307), .B(n399), .Z(n400) );
  NAND U940 ( .A(n27397), .B(n400), .Z(n401) );
  NAND U941 ( .A(n27398), .B(n401), .Z(n402) );
  NAND U942 ( .A(n27399), .B(n402), .Z(n27400) );
  NAND U943 ( .A(n12992), .B(n12991), .Z(n403) );
  AND U944 ( .A(n12993), .B(n403), .Z(n27425) );
  NANDN U945 ( .A(n27438), .B(n27437), .Z(n404) );
  NANDN U946 ( .A(n27439), .B(n404), .Z(n405) );
  NAND U947 ( .A(n27440), .B(n405), .Z(n406) );
  NAND U948 ( .A(n27441), .B(n406), .Z(n407) );
  NAND U949 ( .A(n27442), .B(n407), .Z(n408) );
  AND U950 ( .A(n27443), .B(n408), .Z(n409) );
  NANDN U951 ( .A(n409), .B(n24294), .Z(n410) );
  NAND U952 ( .A(n27444), .B(n410), .Z(n411) );
  NAND U953 ( .A(n27445), .B(n411), .Z(n412) );
  NANDN U954 ( .A(n27446), .B(n412), .Z(n413) );
  NAND U955 ( .A(n27447), .B(n413), .Z(n414) );
  AND U956 ( .A(n27448), .B(n414), .Z(n415) );
  ANDN U957 ( .B(n27449), .A(n415), .Z(n416) );
  OR U958 ( .A(n24293), .B(n24292), .Z(n417) );
  NAND U959 ( .A(n416), .B(n417), .Z(n418) );
  NAND U960 ( .A(n27450), .B(n418), .Z(n419) );
  NANDN U961 ( .A(n27451), .B(n419), .Z(n27452) );
  NANDN U962 ( .A(x[2140]), .B(n27490), .Z(n420) );
  AND U963 ( .A(n27489), .B(n420), .Z(n421) );
  XNOR U964 ( .A(x[2140]), .B(n27490), .Z(n422) );
  NAND U965 ( .A(y[2140]), .B(n422), .Z(n423) );
  NAND U966 ( .A(n421), .B(n423), .Z(n424) );
  NAND U967 ( .A(n27491), .B(n424), .Z(n425) );
  NAND U968 ( .A(n27492), .B(n425), .Z(n426) );
  AND U969 ( .A(n27493), .B(n426), .Z(n427) );
  NANDN U970 ( .A(n427), .B(n27494), .Z(n428) );
  NAND U971 ( .A(n27495), .B(n428), .Z(n429) );
  NAND U972 ( .A(n27496), .B(n429), .Z(n430) );
  NAND U973 ( .A(n24289), .B(n430), .Z(n431) );
  NAND U974 ( .A(n27497), .B(n431), .Z(n432) );
  AND U975 ( .A(n27498), .B(n432), .Z(n433) );
  NANDN U976 ( .A(n433), .B(n27499), .Z(n434) );
  NAND U977 ( .A(n27500), .B(n434), .Z(n435) );
  NAND U978 ( .A(n27501), .B(n435), .Z(n436) );
  ANDN U979 ( .B(n436), .A(n27502), .Z(n27503) );
  ANDN U980 ( .B(n12914), .A(n12913), .Z(n27525) );
  ANDN U981 ( .B(n19119), .A(n19118), .Z(n24279) );
  NOR U982 ( .A(n19153), .B(n19152), .Z(n437) );
  NANDN U983 ( .A(n19150), .B(n19151), .Z(n438) );
  NAND U984 ( .A(n437), .B(n438), .Z(n27547) );
  ANDN U985 ( .B(n19181), .A(n19180), .Z(n27565) );
  NAND U986 ( .A(n27585), .B(n27584), .Z(n439) );
  NAND U987 ( .A(n27586), .B(n439), .Z(n440) );
  NAND U988 ( .A(n27587), .B(n440), .Z(n441) );
  NAND U989 ( .A(n27588), .B(n441), .Z(n442) );
  NAND U990 ( .A(n27589), .B(n442), .Z(n443) );
  ANDN U991 ( .B(n443), .A(n27590), .Z(n444) );
  NANDN U992 ( .A(n444), .B(n27591), .Z(n445) );
  NANDN U993 ( .A(n27592), .B(n445), .Z(n446) );
  NAND U994 ( .A(n24270), .B(n446), .Z(n447) );
  NANDN U995 ( .A(n27593), .B(n447), .Z(n448) );
  NAND U996 ( .A(n27594), .B(n448), .Z(n449) );
  ANDN U997 ( .B(n449), .A(n27595), .Z(n450) );
  NANDN U998 ( .A(n450), .B(n27596), .Z(n451) );
  NAND U999 ( .A(n24269), .B(n451), .Z(n452) );
  NAND U1000 ( .A(n27597), .B(n452), .Z(n453) );
  NANDN U1001 ( .A(n27598), .B(n453), .Z(n27599) );
  NANDN U1002 ( .A(n19267), .B(n19266), .Z(n454) );
  ANDN U1003 ( .B(n454), .A(n19268), .Z(n27617) );
  AND U1004 ( .A(n19317), .B(n19318), .Z(n455) );
  NAND U1005 ( .A(n19320), .B(n19319), .Z(n456) );
  AND U1006 ( .A(n455), .B(n456), .Z(n27642) );
  NOR U1007 ( .A(n19343), .B(n19344), .Z(n27653) );
  NAND U1008 ( .A(n12790), .B(n12791), .Z(n457) );
  ANDN U1009 ( .B(n457), .A(n12792), .Z(n27662) );
  ANDN U1010 ( .B(n12779), .A(n12778), .Z(n27682) );
  ANDN U1011 ( .B(n12751), .A(n12750), .Z(n27721) );
  ANDN U1012 ( .B(n12745), .A(n12744), .Z(n27741) );
  NAND U1013 ( .A(n27764), .B(n27765), .Z(n458) );
  NANDN U1014 ( .A(n27766), .B(n458), .Z(n459) );
  AND U1015 ( .A(n24252), .B(n459), .Z(n460) );
  OR U1016 ( .A(n24251), .B(n460), .Z(n461) );
  NAND U1017 ( .A(n24250), .B(n461), .Z(n462) );
  NAND U1018 ( .A(n27767), .B(n462), .Z(n463) );
  NANDN U1019 ( .A(n27768), .B(n463), .Z(n464) );
  NAND U1020 ( .A(n27769), .B(n464), .Z(n465) );
  ANDN U1021 ( .B(n465), .A(n27770), .Z(n466) );
  NANDN U1022 ( .A(n466), .B(n27771), .Z(n467) );
  AND U1023 ( .A(n27772), .B(n467), .Z(n468) );
  NANDN U1024 ( .A(n468), .B(n24249), .Z(n469) );
  NANDN U1025 ( .A(n27773), .B(n469), .Z(n470) );
  NAND U1026 ( .A(n27774), .B(n470), .Z(n27777) );
  NANDN U1027 ( .A(n12710), .B(n12711), .Z(n27805) );
  NANDN U1028 ( .A(n19597), .B(n19598), .Z(n471) );
  NAND U1029 ( .A(n19599), .B(n471), .Z(n27820) );
  NANDN U1030 ( .A(n12680), .B(n12681), .Z(n27837) );
  NAND U1031 ( .A(n12668), .B(n12667), .Z(n472) );
  AND U1032 ( .A(n12669), .B(n472), .Z(n27852) );
  ANDN U1033 ( .B(n12658), .A(n12657), .Z(n27872) );
  NANDN U1034 ( .A(n12648), .B(n12649), .Z(n27891) );
  NANDN U1035 ( .A(n24234), .B(n27911), .Z(n473) );
  NAND U1036 ( .A(n27912), .B(n473), .Z(n474) );
  NAND U1037 ( .A(n24233), .B(n474), .Z(n475) );
  NAND U1038 ( .A(n24232), .B(n24231), .Z(n476) );
  NAND U1039 ( .A(n27913), .B(n475), .Z(n477) );
  NAND U1040 ( .A(n476), .B(n477), .Z(n478) );
  OR U1041 ( .A(n478), .B(n27914), .Z(n479) );
  NAND U1042 ( .A(n24230), .B(n479), .Z(n480) );
  NAND U1043 ( .A(n27915), .B(n480), .Z(n481) );
  NANDN U1044 ( .A(n27916), .B(n481), .Z(n482) );
  NAND U1045 ( .A(n27917), .B(n482), .Z(n483) );
  ANDN U1046 ( .B(n483), .A(n27918), .Z(n484) );
  NANDN U1047 ( .A(n484), .B(n27919), .Z(n485) );
  NAND U1048 ( .A(n27920), .B(n485), .Z(n486) );
  NAND U1049 ( .A(n24229), .B(n486), .Z(n27921) );
  ANDN U1050 ( .B(n12597), .A(n12596), .Z(n27960) );
  ANDN U1051 ( .B(n19873), .A(n12579), .Z(n487) );
  NANDN U1052 ( .A(n12577), .B(n12578), .Z(n488) );
  NAND U1053 ( .A(n487), .B(n488), .Z(n24220) );
  NAND U1054 ( .A(n28022), .B(n28023), .Z(n489) );
  AND U1055 ( .A(n28028), .B(n489), .Z(n490) );
  NAND U1056 ( .A(n490), .B(n28027), .Z(n491) );
  NAND U1057 ( .A(n28029), .B(n491), .Z(n492) );
  NANDN U1058 ( .A(n28030), .B(n492), .Z(n493) );
  AND U1059 ( .A(n28031), .B(n493), .Z(n494) );
  OR U1060 ( .A(n28032), .B(n494), .Z(n495) );
  NAND U1061 ( .A(n24206), .B(n495), .Z(n496) );
  NAND U1062 ( .A(n28033), .B(n496), .Z(n497) );
  NAND U1063 ( .A(n28034), .B(n497), .Z(n498) );
  NANDN U1064 ( .A(n28035), .B(n498), .Z(n499) );
  AND U1065 ( .A(n28036), .B(n499), .Z(n500) );
  ANDN U1066 ( .B(n24205), .A(n500), .Z(n501) );
  OR U1067 ( .A(n24203), .B(n24204), .Z(n502) );
  NAND U1068 ( .A(n501), .B(n502), .Z(n503) );
  NAND U1069 ( .A(n28037), .B(n503), .Z(n28041) );
  OR U1070 ( .A(n28072), .B(n28073), .Z(n504) );
  NANDN U1071 ( .A(n28074), .B(n504), .Z(n505) );
  AND U1072 ( .A(n28075), .B(n505), .Z(n506) );
  OR U1073 ( .A(n28076), .B(n506), .Z(n507) );
  NAND U1074 ( .A(n28077), .B(n507), .Z(n508) );
  NAND U1075 ( .A(n28078), .B(n508), .Z(n509) );
  NOR U1076 ( .A(n28080), .B(n28079), .Z(n510) );
  NAND U1077 ( .A(n509), .B(n510), .Z(n511) );
  NAND U1078 ( .A(n28081), .B(n511), .Z(n512) );
  NANDN U1079 ( .A(n28082), .B(n512), .Z(n513) );
  NANDN U1080 ( .A(n24199), .B(n513), .Z(n514) );
  AND U1081 ( .A(n28083), .B(n514), .Z(n515) );
  OR U1082 ( .A(n28084), .B(n515), .Z(n516) );
  AND U1083 ( .A(n28085), .B(n516), .Z(n517) );
  OR U1084 ( .A(n28086), .B(n517), .Z(n518) );
  NAND U1085 ( .A(n28087), .B(n518), .Z(n519) );
  NAND U1086 ( .A(n28088), .B(n519), .Z(n28089) );
  NANDN U1087 ( .A(n12473), .B(n12474), .Z(n28114) );
  NANDN U1088 ( .A(n12461), .B(n12462), .Z(n28122) );
  NANDN U1089 ( .A(n28152), .B(n28153), .Z(n520) );
  NAND U1090 ( .A(n28154), .B(n520), .Z(n521) );
  AND U1091 ( .A(n28155), .B(n521), .Z(n522) );
  NANDN U1092 ( .A(n28156), .B(n522), .Z(n523) );
  NAND U1093 ( .A(n28157), .B(n523), .Z(n524) );
  ANDN U1094 ( .B(n524), .A(n24175), .Z(n525) );
  NANDN U1095 ( .A(n525), .B(n24174), .Z(n526) );
  NAND U1096 ( .A(n28158), .B(n526), .Z(n527) );
  NAND U1097 ( .A(n28159), .B(n527), .Z(n528) );
  NANDN U1098 ( .A(n24172), .B(n24173), .Z(n529) );
  NANDN U1099 ( .A(n528), .B(n529), .Z(n530) );
  AND U1100 ( .A(n28160), .B(n530), .Z(n531) );
  OR U1101 ( .A(n28161), .B(n531), .Z(n532) );
  AND U1102 ( .A(n28162), .B(n532), .Z(n533) );
  OR U1103 ( .A(n28163), .B(n533), .Z(n534) );
  NAND U1104 ( .A(n28164), .B(n534), .Z(n535) );
  NAND U1105 ( .A(n28165), .B(n535), .Z(n28166) );
  NANDN U1106 ( .A(n24168), .B(n28201), .Z(n536) );
  NAND U1107 ( .A(n28202), .B(n536), .Z(n537) );
  NAND U1108 ( .A(n28203), .B(n537), .Z(n538) );
  NANDN U1109 ( .A(n24167), .B(n538), .Z(n539) );
  NAND U1110 ( .A(n28204), .B(n539), .Z(n540) );
  AND U1111 ( .A(n28205), .B(n540), .Z(n541) );
  NANDN U1112 ( .A(n541), .B(n28206), .Z(n542) );
  NANDN U1113 ( .A(n24166), .B(n542), .Z(n543) );
  NAND U1114 ( .A(n24165), .B(n543), .Z(n544) );
  NANDN U1115 ( .A(n28207), .B(n544), .Z(n545) );
  NAND U1116 ( .A(n28208), .B(n545), .Z(n546) );
  AND U1117 ( .A(n24164), .B(n546), .Z(n547) );
  NANDN U1118 ( .A(n547), .B(n28209), .Z(n548) );
  AND U1119 ( .A(n28210), .B(n548), .Z(n28211) );
  XNOR U1120 ( .A(x[2818]), .B(y[2818]), .Z(n549) );
  ANDN U1121 ( .B(n549), .A(n12389), .Z(n28239) );
  ANDN U1122 ( .B(n12380), .A(n12379), .Z(n28253) );
  ANDN U1123 ( .B(n12373), .A(n12372), .Z(n28277) );
  ANDN U1124 ( .B(n12350), .A(n12349), .Z(n28310) );
  ANDN U1125 ( .B(n12331), .A(n12330), .Z(n28337) );
  NANDN U1126 ( .A(x[2906]), .B(y[2906]), .Z(n550) );
  ANDN U1127 ( .B(n550), .A(n20607), .Z(n28366) );
  ANDN U1128 ( .B(n12298), .A(n12297), .Z(n28378) );
  ANDN U1129 ( .B(n12271), .A(n12270), .Z(n24130) );
  NANDN U1130 ( .A(n20732), .B(n20733), .Z(n28427) );
  ANDN U1131 ( .B(n12243), .A(n24121), .Z(n28443) );
  NOR U1132 ( .A(n20824), .B(n20825), .Z(n28472) );
  NANDN U1133 ( .A(x[3016]), .B(y[3016]), .Z(n551) );
  ANDN U1134 ( .B(n551), .A(n12212), .Z(n28482) );
  NAND U1135 ( .A(n28529), .B(n28528), .Z(n552) );
  NAND U1136 ( .A(n24099), .B(n552), .Z(n553) );
  NAND U1137 ( .A(n28530), .B(n553), .Z(n554) );
  NAND U1138 ( .A(n24098), .B(n554), .Z(n555) );
  NANDN U1139 ( .A(n28531), .B(n555), .Z(n556) );
  AND U1140 ( .A(n28532), .B(n556), .Z(n557) );
  NANDN U1141 ( .A(n24097), .B(n24096), .Z(n558) );
  NANDN U1142 ( .A(n557), .B(n28533), .Z(n559) );
  NAND U1143 ( .A(n558), .B(n559), .Z(n560) );
  NANDN U1144 ( .A(n560), .B(n28534), .Z(n561) );
  NANDN U1145 ( .A(n28535), .B(n561), .Z(n562) );
  NAND U1146 ( .A(n28536), .B(n562), .Z(n563) );
  NANDN U1147 ( .A(n28537), .B(n563), .Z(n564) );
  NAND U1148 ( .A(n28538), .B(n564), .Z(n565) );
  ANDN U1149 ( .B(n565), .A(n28539), .Z(n566) );
  NANDN U1150 ( .A(n566), .B(n28540), .Z(n567) );
  NANDN U1151 ( .A(n28541), .B(n567), .Z(n568) );
  NAND U1152 ( .A(n28542), .B(n568), .Z(n28543) );
  AND U1153 ( .A(n29050), .B(n29051), .Z(n29052) );
  ANDN U1154 ( .B(n29212), .A(n29213), .Z(n29214) );
  NAND U1155 ( .A(n29252), .B(n29251), .Z(n569) );
  NANDN U1156 ( .A(n29253), .B(n569), .Z(n570) );
  AND U1157 ( .A(n29254), .B(n570), .Z(n571) );
  OR U1158 ( .A(n29255), .B(n571), .Z(n572) );
  NAND U1159 ( .A(n29256), .B(n572), .Z(n573) );
  NANDN U1160 ( .A(n29257), .B(n573), .Z(n574) );
  ANDN U1161 ( .B(n23920), .A(n23919), .Z(n575) );
  NAND U1162 ( .A(n574), .B(n575), .Z(n576) );
  NAND U1163 ( .A(n29258), .B(n576), .Z(n577) );
  ANDN U1164 ( .B(n29259), .A(n29260), .Z(n578) );
  NAND U1165 ( .A(n577), .B(n578), .Z(n579) );
  NANDN U1166 ( .A(n29261), .B(n579), .Z(n580) );
  AND U1167 ( .A(n23918), .B(n29262), .Z(n581) );
  NAND U1168 ( .A(n580), .B(n581), .Z(n582) );
  NANDN U1169 ( .A(n23917), .B(n582), .Z(n583) );
  NAND U1170 ( .A(n23916), .B(n583), .Z(n29265) );
  AND U1171 ( .A(n29317), .B(n29318), .Z(n29319) );
  NANDN U1172 ( .A(n29483), .B(n29484), .Z(n584) );
  NAND U1173 ( .A(n29485), .B(n584), .Z(n585) );
  ANDN U1174 ( .B(n585), .A(n29486), .Z(n586) );
  NANDN U1175 ( .A(n29487), .B(n586), .Z(n587) );
  NANDN U1176 ( .A(n29488), .B(n587), .Z(n588) );
  AND U1177 ( .A(n29489), .B(n588), .Z(n589) );
  AND U1178 ( .A(n23861), .B(n23862), .Z(n590) );
  NANDN U1179 ( .A(n589), .B(n29490), .Z(n591) );
  AND U1180 ( .A(n590), .B(n591), .Z(n592) );
  AND U1181 ( .A(n29493), .B(n29492), .Z(n593) );
  NANDN U1182 ( .A(n592), .B(n29491), .Z(n594) );
  AND U1183 ( .A(n593), .B(n594), .Z(n595) );
  AND U1184 ( .A(n29496), .B(n29495), .Z(n596) );
  NANDN U1185 ( .A(n595), .B(n29494), .Z(n597) );
  AND U1186 ( .A(n596), .B(n597), .Z(n29499) );
  NANDN U1187 ( .A(n15453), .B(n15454), .Z(n24577) );
  NANDN U1188 ( .A(n15409), .B(n15410), .Z(n24621) );
  NANDN U1189 ( .A(n15377), .B(n15378), .Z(n24653) );
  NANDN U1190 ( .A(n15350), .B(n15351), .Z(n24697) );
  NANDN U1191 ( .A(x[100]), .B(y[100]), .Z(n598) );
  ANDN U1192 ( .B(n598), .A(n15314), .Z(n24735) );
  ANDN U1193 ( .B(n15271), .A(n15270), .Z(n24779) );
  ANDN U1194 ( .B(n15232), .A(n15231), .Z(n24823) );
  ANDN U1195 ( .B(n15194), .A(n15193), .Z(n24863) );
  ANDN U1196 ( .B(n15152), .A(n15151), .Z(n24903) );
  ANDN U1197 ( .B(n15116), .A(n15115), .Z(n24939) );
  ANDN U1198 ( .B(n15072), .A(n15071), .Z(n24983) );
  ANDN U1199 ( .B(n15033), .A(n15032), .Z(n25023) );
  ANDN U1200 ( .B(n15003), .A(n15002), .Z(n25055) );
  ANDN U1201 ( .B(n14976), .A(n14975), .Z(n25095) );
  ANDN U1202 ( .B(n14928), .A(n14927), .Z(n25143) );
  NANDN U1203 ( .A(n14889), .B(n14890), .Z(n25181) );
  NANDN U1204 ( .A(n14854), .B(n14855), .Z(n25225) );
  NANDN U1205 ( .A(n14822), .B(n14823), .Z(n25248) );
  NANDN U1206 ( .A(n14786), .B(n14787), .Z(n25281) );
  NANDN U1207 ( .A(n14770), .B(n14771), .Z(n25297) );
  NANDN U1208 ( .A(n14730), .B(n14731), .Z(n25361) );
  NANDN U1209 ( .A(n14700), .B(n14701), .Z(n25397) );
  NANDN U1210 ( .A(n14660), .B(n14661), .Z(n25437) );
  NANDN U1211 ( .A(n14616), .B(n14617), .Z(n25481) );
  NANDN U1212 ( .A(n14571), .B(n14572), .Z(n25525) );
  NANDN U1213 ( .A(n14541), .B(n14542), .Z(n25545) );
  NANDN U1214 ( .A(n14493), .B(n14494), .Z(n25588) );
  NANDN U1215 ( .A(n14453), .B(n14454), .Z(n25628) );
  NANDN U1216 ( .A(n14443), .B(n14444), .Z(n25636) );
  NANDN U1217 ( .A(n14399), .B(n14400), .Z(n25682) );
  NANDN U1218 ( .A(n14359), .B(n14360), .Z(n25722) );
  NANDN U1219 ( .A(n14323), .B(n14324), .Z(n25758) );
  NANDN U1220 ( .A(n14279), .B(n14280), .Z(n25802) );
  NANDN U1221 ( .A(n14239), .B(n14240), .Z(n25846) );
  ANDN U1222 ( .B(n16219), .A(n16218), .Z(n25864) );
  ANDN U1223 ( .B(n14197), .A(n14196), .Z(n25874) );
  NANDN U1224 ( .A(n24522), .B(n25897), .Z(n599) );
  NAND U1225 ( .A(n25898), .B(n599), .Z(n600) );
  ANDN U1226 ( .B(n600), .A(n25899), .Z(n601) );
  NANDN U1227 ( .A(n601), .B(n25900), .Z(n602) );
  NAND U1228 ( .A(n25901), .B(n602), .Z(n603) );
  NAND U1229 ( .A(n25902), .B(n603), .Z(n604) );
  NAND U1230 ( .A(n25903), .B(n604), .Z(n605) );
  NAND U1231 ( .A(n24521), .B(n605), .Z(n606) );
  AND U1232 ( .A(n25904), .B(n606), .Z(n607) );
  NANDN U1233 ( .A(n607), .B(n25905), .Z(n608) );
  NAND U1234 ( .A(n25906), .B(n608), .Z(n609) );
  NAND U1235 ( .A(n24520), .B(n609), .Z(n610) );
  NAND U1236 ( .A(n25907), .B(n610), .Z(n611) );
  NAND U1237 ( .A(n24519), .B(n611), .Z(n612) );
  AND U1238 ( .A(n25908), .B(n612), .Z(n25911) );
  NOR U1239 ( .A(n14097), .B(n14098), .Z(n25926) );
  XNOR U1240 ( .A(x[782]), .B(y[782]), .Z(n613) );
  ANDN U1241 ( .B(n613), .A(n14090), .Z(n25933) );
  NANDN U1242 ( .A(n14026), .B(n14027), .Z(n25990) );
  NANDN U1243 ( .A(n14016), .B(n14017), .Z(n26027) );
  NANDN U1244 ( .A(n26049), .B(n26048), .Z(n614) );
  NANDN U1245 ( .A(n26050), .B(n614), .Z(n615) );
  NAND U1246 ( .A(n26051), .B(n615), .Z(n616) );
  NANDN U1247 ( .A(n26052), .B(n616), .Z(n617) );
  NAND U1248 ( .A(n26053), .B(n617), .Z(n618) );
  ANDN U1249 ( .B(n618), .A(n26054), .Z(n619) );
  ANDN U1250 ( .B(n26055), .A(n619), .Z(n620) );
  NAND U1251 ( .A(n26056), .B(n620), .Z(n621) );
  ANDN U1252 ( .B(n621), .A(n26057), .Z(n622) );
  NANDN U1253 ( .A(n622), .B(n26058), .Z(n623) );
  NAND U1254 ( .A(n26059), .B(n623), .Z(n624) );
  NANDN U1255 ( .A(n24507), .B(n624), .Z(n625) );
  NAND U1256 ( .A(n26060), .B(n625), .Z(n626) );
  NANDN U1257 ( .A(n24506), .B(n626), .Z(n627) );
  AND U1258 ( .A(n26061), .B(n627), .Z(n628) );
  NANDN U1259 ( .A(n628), .B(n26062), .Z(n629) );
  NANDN U1260 ( .A(n26063), .B(n629), .Z(n630) );
  NAND U1261 ( .A(n26064), .B(n630), .Z(n26065) );
  OR U1262 ( .A(n26094), .B(n26095), .Z(n631) );
  NAND U1263 ( .A(n26096), .B(n631), .Z(n632) );
  NAND U1264 ( .A(n24499), .B(n632), .Z(n633) );
  NAND U1265 ( .A(n26097), .B(n633), .Z(n634) );
  NANDN U1266 ( .A(n26098), .B(n634), .Z(n635) );
  AND U1267 ( .A(n26099), .B(n635), .Z(n636) );
  NANDN U1268 ( .A(n636), .B(n26100), .Z(n637) );
  NANDN U1269 ( .A(n24498), .B(n637), .Z(n638) );
  NAND U1270 ( .A(n24497), .B(n638), .Z(n639) );
  NAND U1271 ( .A(n26101), .B(n639), .Z(n640) );
  NANDN U1272 ( .A(n26102), .B(n640), .Z(n641) );
  AND U1273 ( .A(n26103), .B(n641), .Z(n642) );
  ANDN U1274 ( .B(n26106), .A(n642), .Z(n643) );
  NANDN U1275 ( .A(n26105), .B(n26104), .Z(n644) );
  NAND U1276 ( .A(n643), .B(n644), .Z(n645) );
  NAND U1277 ( .A(n26107), .B(n645), .Z(n26108) );
  ANDN U1278 ( .B(n13941), .A(n13940), .Z(n26122) );
  ANDN U1279 ( .B(n13925), .A(n13924), .Z(n26140) );
  ANDN U1280 ( .B(n13899), .A(n13898), .Z(n26163) );
  NAND U1281 ( .A(n26188), .B(n26189), .Z(n646) );
  NAND U1282 ( .A(n26190), .B(n646), .Z(n647) );
  AND U1283 ( .A(n26191), .B(n647), .Z(n648) );
  NANDN U1284 ( .A(n648), .B(n26192), .Z(n649) );
  NAND U1285 ( .A(n26193), .B(n649), .Z(n650) );
  NAND U1286 ( .A(n24483), .B(n650), .Z(n651) );
  NANDN U1287 ( .A(n26194), .B(n651), .Z(n652) );
  NANDN U1288 ( .A(n26195), .B(n652), .Z(n653) );
  AND U1289 ( .A(n26196), .B(n653), .Z(n654) );
  OR U1290 ( .A(n654), .B(n26197), .Z(n655) );
  NANDN U1291 ( .A(n24482), .B(n655), .Z(n656) );
  AND U1292 ( .A(n26198), .B(n656), .Z(n657) );
  NANDN U1293 ( .A(n657), .B(n26199), .Z(n658) );
  NAND U1294 ( .A(n26200), .B(n658), .Z(n659) );
  NAND U1295 ( .A(n26201), .B(n659), .Z(n660) );
  NAND U1296 ( .A(n26202), .B(n660), .Z(n26203) );
  NANDN U1297 ( .A(n13842), .B(n13843), .Z(n26225) );
  NANDN U1298 ( .A(n26247), .B(n26246), .Z(n661) );
  NAND U1299 ( .A(n26248), .B(n661), .Z(n662) );
  ANDN U1300 ( .B(n662), .A(n26249), .Z(n663) );
  OR U1301 ( .A(n26250), .B(n663), .Z(n664) );
  NAND U1302 ( .A(n26251), .B(n664), .Z(n665) );
  NAND U1303 ( .A(n26252), .B(n665), .Z(n666) );
  NAND U1304 ( .A(n26253), .B(n666), .Z(n667) );
  NAND U1305 ( .A(n26254), .B(n667), .Z(n668) );
  AND U1306 ( .A(n24471), .B(n668), .Z(n669) );
  OR U1307 ( .A(n26255), .B(n669), .Z(n670) );
  ANDN U1308 ( .B(n670), .A(n26256), .Z(n671) );
  OR U1309 ( .A(n26257), .B(n671), .Z(n672) );
  NAND U1310 ( .A(n26258), .B(n672), .Z(n673) );
  NANDN U1311 ( .A(n24470), .B(n673), .Z(n26259) );
  NAND U1312 ( .A(n13802), .B(n13801), .Z(n674) );
  AND U1313 ( .A(n13803), .B(n674), .Z(n26284) );
  NAND U1314 ( .A(n26305), .B(n26304), .Z(n675) );
  NAND U1315 ( .A(n26306), .B(n675), .Z(n676) );
  NAND U1316 ( .A(n26307), .B(n676), .Z(n677) );
  NAND U1317 ( .A(n24459), .B(n677), .Z(n678) );
  NAND U1318 ( .A(n26308), .B(n678), .Z(n679) );
  AND U1319 ( .A(n26309), .B(n679), .Z(n680) );
  OR U1320 ( .A(n26310), .B(n680), .Z(n681) );
  NAND U1321 ( .A(n26311), .B(n681), .Z(n682) );
  NAND U1322 ( .A(n26312), .B(n682), .Z(n683) );
  NANDN U1323 ( .A(n26313), .B(n683), .Z(n684) );
  NAND U1324 ( .A(n26314), .B(n684), .Z(n685) );
  AND U1325 ( .A(n26315), .B(n685), .Z(n686) );
  NAND U1326 ( .A(n26316), .B(n26317), .Z(n687) );
  AND U1327 ( .A(n26318), .B(n687), .Z(n688) );
  NANDN U1328 ( .A(n686), .B(n688), .Z(n689) );
  NANDN U1329 ( .A(n26319), .B(n689), .Z(n26320) );
  ANDN U1330 ( .B(n13748), .A(n13747), .Z(n26341) );
  OR U1331 ( .A(n26356), .B(n26357), .Z(n690) );
  NAND U1332 ( .A(n26358), .B(n690), .Z(n691) );
  ANDN U1333 ( .B(n691), .A(n26359), .Z(n692) );
  NANDN U1334 ( .A(n692), .B(n26360), .Z(n693) );
  NAND U1335 ( .A(n26361), .B(n693), .Z(n694) );
  NANDN U1336 ( .A(n26362), .B(n694), .Z(n695) );
  NAND U1337 ( .A(n26363), .B(n695), .Z(n696) );
  NAND U1338 ( .A(n26364), .B(n696), .Z(n697) );
  ANDN U1339 ( .B(n697), .A(n26365), .Z(n698) );
  OR U1340 ( .A(n26366), .B(n698), .Z(n699) );
  NAND U1341 ( .A(n26367), .B(n699), .Z(n700) );
  NANDN U1342 ( .A(n26368), .B(n700), .Z(n701) );
  NAND U1343 ( .A(n26369), .B(n701), .Z(n702) );
  NANDN U1344 ( .A(n26370), .B(n702), .Z(n703) );
  AND U1345 ( .A(n26371), .B(n703), .Z(n704) );
  OR U1346 ( .A(n26372), .B(n704), .Z(n705) );
  NAND U1347 ( .A(n26373), .B(n705), .Z(n706) );
  NANDN U1348 ( .A(n26374), .B(n706), .Z(n707) );
  NAND U1349 ( .A(n24446), .B(n707), .Z(n26376) );
  ANDN U1350 ( .B(n13695), .A(n13694), .Z(n26403) );
  ANDN U1351 ( .B(n13690), .A(n13689), .Z(n26434) );
  NAND U1352 ( .A(n26461), .B(n26462), .Z(n708) );
  NANDN U1353 ( .A(n26463), .B(n708), .Z(n709) );
  ANDN U1354 ( .B(n709), .A(n24436), .Z(n710) );
  OR U1355 ( .A(n710), .B(n26464), .Z(n711) );
  NANDN U1356 ( .A(n26465), .B(n711), .Z(n712) );
  AND U1357 ( .A(n26466), .B(n712), .Z(n713) );
  NANDN U1358 ( .A(n713), .B(n26467), .Z(n714) );
  NANDN U1359 ( .A(n26468), .B(n714), .Z(n715) );
  NAND U1360 ( .A(n26469), .B(n715), .Z(n716) );
  NANDN U1361 ( .A(n26470), .B(n716), .Z(n717) );
  NANDN U1362 ( .A(n26471), .B(n717), .Z(n718) );
  ANDN U1363 ( .B(n718), .A(n26472), .Z(n719) );
  NANDN U1364 ( .A(n719), .B(n26473), .Z(n720) );
  ANDN U1365 ( .B(n720), .A(n26474), .Z(n721) );
  NANDN U1366 ( .A(n721), .B(n26475), .Z(n722) );
  NAND U1367 ( .A(n26476), .B(n722), .Z(n723) );
  NAND U1368 ( .A(n26477), .B(n723), .Z(n26478) );
  ANDN U1369 ( .B(n13651), .A(n13650), .Z(n26499) );
  NOR U1370 ( .A(n17363), .B(n17364), .Z(n26515) );
  OR U1371 ( .A(n26531), .B(n26532), .Z(n724) );
  NAND U1372 ( .A(n26533), .B(n724), .Z(n725) );
  NANDN U1373 ( .A(n26534), .B(n725), .Z(n726) );
  NAND U1374 ( .A(n26535), .B(n726), .Z(n727) );
  NANDN U1375 ( .A(n24419), .B(n727), .Z(n728) );
  AND U1376 ( .A(n24418), .B(n728), .Z(n729) );
  OR U1377 ( .A(n24417), .B(n729), .Z(n730) );
  NAND U1378 ( .A(n26536), .B(n730), .Z(n731) );
  NANDN U1379 ( .A(n26537), .B(n731), .Z(n732) );
  NAND U1380 ( .A(n26538), .B(n732), .Z(n733) );
  NAND U1381 ( .A(n26539), .B(n733), .Z(n734) );
  ANDN U1382 ( .B(n734), .A(n26540), .Z(n735) );
  NANDN U1383 ( .A(n735), .B(n26541), .Z(n736) );
  NANDN U1384 ( .A(n26542), .B(n736), .Z(n737) );
  NAND U1385 ( .A(n26543), .B(n737), .Z(n738) );
  NANDN U1386 ( .A(n26544), .B(n738), .Z(n26546) );
  NAND U1387 ( .A(n26575), .B(n26574), .Z(n739) );
  NAND U1388 ( .A(n24410), .B(n24411), .Z(n740) );
  NAND U1389 ( .A(n739), .B(n740), .Z(n741) );
  OR U1390 ( .A(n741), .B(n26576), .Z(n742) );
  NAND U1391 ( .A(n26578), .B(n26577), .Z(n743) );
  AND U1392 ( .A(n742), .B(n743), .Z(n744) );
  NAND U1393 ( .A(n26579), .B(n744), .Z(n745) );
  NANDN U1394 ( .A(n26580), .B(n745), .Z(n746) );
  NAND U1395 ( .A(n26581), .B(n746), .Z(n747) );
  NANDN U1396 ( .A(n26582), .B(n747), .Z(n748) );
  NAND U1397 ( .A(n26583), .B(n748), .Z(n749) );
  ANDN U1398 ( .B(n749), .A(n26584), .Z(n750) );
  NANDN U1399 ( .A(n750), .B(n24409), .Z(n751) );
  NANDN U1400 ( .A(n26585), .B(n751), .Z(n752) );
  NAND U1401 ( .A(n26586), .B(n752), .Z(n26587) );
  ANDN U1402 ( .B(n17552), .A(n17551), .Z(n26605) );
  NANDN U1403 ( .A(n13560), .B(n13561), .Z(n26649) );
  NANDN U1404 ( .A(n13547), .B(n13548), .Z(n26670) );
  NANDN U1405 ( .A(n26696), .B(n26695), .Z(n753) );
  NAND U1406 ( .A(n26697), .B(n753), .Z(n754) );
  ANDN U1407 ( .B(n754), .A(n26698), .Z(n755) );
  NANDN U1408 ( .A(n755), .B(n26699), .Z(n756) );
  NAND U1409 ( .A(n26700), .B(n756), .Z(n757) );
  NANDN U1410 ( .A(n26701), .B(n757), .Z(n758) );
  NAND U1411 ( .A(n26702), .B(n758), .Z(n759) );
  NAND U1412 ( .A(n26703), .B(n759), .Z(n760) );
  ANDN U1413 ( .B(n760), .A(n26704), .Z(n761) );
  NANDN U1414 ( .A(n761), .B(n26705), .Z(n762) );
  NANDN U1415 ( .A(n26706), .B(n762), .Z(n763) );
  NAND U1416 ( .A(n26707), .B(n763), .Z(n764) );
  NANDN U1417 ( .A(n26708), .B(n764), .Z(n765) );
  NAND U1418 ( .A(n26709), .B(n765), .Z(n766) );
  ANDN U1419 ( .B(n766), .A(n26710), .Z(n767) );
  NANDN U1420 ( .A(n767), .B(n26711), .Z(n768) );
  NANDN U1421 ( .A(n26712), .B(n768), .Z(n769) );
  NAND U1422 ( .A(n26713), .B(n769), .Z(n770) );
  NANDN U1423 ( .A(n26714), .B(n770), .Z(n26715) );
  NANDN U1424 ( .A(n13518), .B(n13519), .Z(n26740) );
  NANDN U1425 ( .A(n13511), .B(n13512), .Z(n771) );
  NAND U1426 ( .A(n13513), .B(n771), .Z(n772) );
  ANDN U1427 ( .B(n772), .A(n13514), .Z(n26750) );
  NANDN U1428 ( .A(n26781), .B(n26780), .Z(n773) );
  NAND U1429 ( .A(n26782), .B(n773), .Z(n774) );
  ANDN U1430 ( .B(n774), .A(n26783), .Z(n775) );
  NANDN U1431 ( .A(n775), .B(n26784), .Z(n776) );
  NANDN U1432 ( .A(n26785), .B(n776), .Z(n777) );
  NANDN U1433 ( .A(n26786), .B(n777), .Z(n778) );
  NAND U1434 ( .A(n26787), .B(n778), .Z(n779) );
  NANDN U1435 ( .A(n24394), .B(n779), .Z(n780) );
  ANDN U1436 ( .B(n780), .A(n26788), .Z(n781) );
  NANDN U1437 ( .A(n781), .B(n26789), .Z(n782) );
  NAND U1438 ( .A(n24393), .B(n782), .Z(n783) );
  NANDN U1439 ( .A(n26790), .B(n783), .Z(n784) );
  NAND U1440 ( .A(n26791), .B(n784), .Z(n785) );
  NANDN U1441 ( .A(n26792), .B(n785), .Z(n786) );
  AND U1442 ( .A(n26793), .B(n786), .Z(n787) );
  OR U1443 ( .A(n26794), .B(n787), .Z(n788) );
  AND U1444 ( .A(n26795), .B(n788), .Z(n26796) );
  ANDN U1445 ( .B(n17893), .A(n17892), .Z(n26816) );
  NAND U1446 ( .A(n13463), .B(n13464), .Z(n789) );
  ANDN U1447 ( .B(n789), .A(n13465), .Z(n26826) );
  NAND U1448 ( .A(n13457), .B(n13458), .Z(n790) );
  NANDN U1449 ( .A(n13456), .B(n790), .Z(n26838) );
  OR U1450 ( .A(n26870), .B(n26871), .Z(n791) );
  NAND U1451 ( .A(n26872), .B(n791), .Z(n792) );
  NANDN U1452 ( .A(n26873), .B(n792), .Z(n793) );
  NAND U1453 ( .A(n26874), .B(n793), .Z(n794) );
  NAND U1454 ( .A(n26875), .B(n794), .Z(n795) );
  ANDN U1455 ( .B(n795), .A(n26876), .Z(n796) );
  NANDN U1456 ( .A(n796), .B(n24380), .Z(n797) );
  NANDN U1457 ( .A(n24379), .B(n797), .Z(n798) );
  NAND U1458 ( .A(n24378), .B(n798), .Z(n799) );
  NANDN U1459 ( .A(n26877), .B(n799), .Z(n800) );
  NAND U1460 ( .A(n26878), .B(n800), .Z(n801) );
  ANDN U1461 ( .B(n801), .A(n24377), .Z(n802) );
  NANDN U1462 ( .A(n802), .B(n26879), .Z(n803) );
  NAND U1463 ( .A(n26880), .B(n803), .Z(n804) );
  NAND U1464 ( .A(n24376), .B(n804), .Z(n26883) );
  NANDN U1465 ( .A(n26912), .B(n26911), .Z(n805) );
  NANDN U1466 ( .A(n24369), .B(n805), .Z(n806) );
  NAND U1467 ( .A(n26913), .B(n806), .Z(n807) );
  NAND U1468 ( .A(n26914), .B(n807), .Z(n808) );
  NAND U1469 ( .A(n26915), .B(n808), .Z(n809) );
  AND U1470 ( .A(n26916), .B(n809), .Z(n810) );
  NANDN U1471 ( .A(n810), .B(n26917), .Z(n811) );
  NANDN U1472 ( .A(n26918), .B(n811), .Z(n812) );
  NANDN U1473 ( .A(n26919), .B(n812), .Z(n813) );
  NANDN U1474 ( .A(n26920), .B(n813), .Z(n814) );
  NAND U1475 ( .A(n24368), .B(n814), .Z(n815) );
  AND U1476 ( .A(n26921), .B(n815), .Z(n816) );
  OR U1477 ( .A(n26922), .B(n816), .Z(n817) );
  NAND U1478 ( .A(n26923), .B(n817), .Z(n818) );
  NANDN U1479 ( .A(n26924), .B(n818), .Z(n819) );
  NAND U1480 ( .A(n26925), .B(n819), .Z(n820) );
  NANDN U1481 ( .A(n26926), .B(n820), .Z(n821) );
  AND U1482 ( .A(n26927), .B(n821), .Z(n26928) );
  AND U1483 ( .A(n26960), .B(n26961), .Z(n822) );
  OR U1484 ( .A(n26958), .B(n26959), .Z(n823) );
  NAND U1485 ( .A(n822), .B(n823), .Z(n824) );
  ANDN U1486 ( .B(n24364), .A(n26962), .Z(n825) );
  NAND U1487 ( .A(n824), .B(n825), .Z(n826) );
  NAND U1488 ( .A(n26963), .B(n826), .Z(n827) );
  ANDN U1489 ( .B(n26965), .A(n26966), .Z(n828) );
  NANDN U1490 ( .A(n827), .B(n26964), .Z(n829) );
  AND U1491 ( .A(n828), .B(n829), .Z(n830) );
  NANDN U1492 ( .A(n830), .B(n26967), .Z(n831) );
  NAND U1493 ( .A(n26968), .B(n831), .Z(n832) );
  NAND U1494 ( .A(n26969), .B(n832), .Z(n833) );
  NANDN U1495 ( .A(n26970), .B(n833), .Z(n834) );
  NANDN U1496 ( .A(n26971), .B(n834), .Z(n835) );
  AND U1497 ( .A(n26972), .B(n835), .Z(n836) );
  OR U1498 ( .A(n26973), .B(n836), .Z(n837) );
  NAND U1499 ( .A(n26974), .B(n837), .Z(n838) );
  NANDN U1500 ( .A(n26975), .B(n838), .Z(n26976) );
  NAND U1501 ( .A(n27007), .B(n27008), .Z(n839) );
  AND U1502 ( .A(n27010), .B(n839), .Z(n840) );
  NANDN U1503 ( .A(n27009), .B(n840), .Z(n841) );
  NAND U1504 ( .A(n24358), .B(n841), .Z(n842) );
  NAND U1505 ( .A(n27011), .B(n842), .Z(n843) );
  AND U1506 ( .A(n27012), .B(n843), .Z(n844) );
  NANDN U1507 ( .A(n844), .B(n27013), .Z(n845) );
  NAND U1508 ( .A(n24357), .B(n845), .Z(n846) );
  NANDN U1509 ( .A(n24356), .B(n846), .Z(n847) );
  NANDN U1510 ( .A(n27014), .B(n847), .Z(n848) );
  NAND U1511 ( .A(n27015), .B(n848), .Z(n849) );
  AND U1512 ( .A(n27016), .B(n849), .Z(n850) );
  NANDN U1513 ( .A(n850), .B(n27017), .Z(n851) );
  NAND U1514 ( .A(n27018), .B(n851), .Z(n852) );
  NANDN U1515 ( .A(n27019), .B(n852), .Z(n27020) );
  OR U1516 ( .A(n27055), .B(n27056), .Z(n853) );
  NANDN U1517 ( .A(n24352), .B(n853), .Z(n854) );
  AND U1518 ( .A(n24351), .B(n854), .Z(n855) );
  NANDN U1519 ( .A(n855), .B(n27057), .Z(n856) );
  NAND U1520 ( .A(n24350), .B(n856), .Z(n857) );
  NAND U1521 ( .A(n27058), .B(n857), .Z(n858) );
  NAND U1522 ( .A(n27059), .B(n858), .Z(n859) );
  NANDN U1523 ( .A(n24349), .B(n859), .Z(n860) );
  AND U1524 ( .A(n24348), .B(n860), .Z(n861) );
  OR U1525 ( .A(n27060), .B(n861), .Z(n862) );
  AND U1526 ( .A(n27061), .B(n862), .Z(n863) );
  OR U1527 ( .A(n27062), .B(n863), .Z(n864) );
  NAND U1528 ( .A(n27063), .B(n864), .Z(n865) );
  NAND U1529 ( .A(n27064), .B(n865), .Z(n27065) );
  NAND U1530 ( .A(n27099), .B(n27100), .Z(n866) );
  NAND U1531 ( .A(n24344), .B(n866), .Z(n867) );
  AND U1532 ( .A(n27101), .B(n867), .Z(n868) );
  OR U1533 ( .A(n24343), .B(n868), .Z(n869) );
  NAND U1534 ( .A(n24342), .B(n869), .Z(n870) );
  NANDN U1535 ( .A(n27102), .B(n870), .Z(n871) );
  NAND U1536 ( .A(n27103), .B(n871), .Z(n872) );
  NAND U1537 ( .A(n27104), .B(n872), .Z(n873) );
  AND U1538 ( .A(n27105), .B(n873), .Z(n874) );
  OR U1539 ( .A(n27106), .B(n874), .Z(n875) );
  AND U1540 ( .A(n27107), .B(n875), .Z(n876) );
  NANDN U1541 ( .A(n876), .B(n27108), .Z(n877) );
  NANDN U1542 ( .A(n27109), .B(n877), .Z(n878) );
  NAND U1543 ( .A(n27110), .B(n878), .Z(n27111) );
  NANDN U1544 ( .A(n13209), .B(n13210), .Z(n27164) );
  NANDN U1545 ( .A(n13187), .B(n13188), .Z(n27185) );
  NANDN U1546 ( .A(n27206), .B(n27205), .Z(n879) );
  NAND U1547 ( .A(n27208), .B(n879), .Z(n880) );
  NAND U1548 ( .A(n27209), .B(n880), .Z(n881) );
  NANDN U1549 ( .A(n24338), .B(n881), .Z(n882) );
  NAND U1550 ( .A(n24337), .B(n882), .Z(n883) );
  ANDN U1551 ( .B(n883), .A(n27210), .Z(n884) );
  NANDN U1552 ( .A(n884), .B(n27211), .Z(n885) );
  NANDN U1553 ( .A(n27212), .B(n885), .Z(n886) );
  NAND U1554 ( .A(n27213), .B(n886), .Z(n887) );
  NANDN U1555 ( .A(n27214), .B(n887), .Z(n888) );
  NAND U1556 ( .A(n27215), .B(n888), .Z(n889) );
  ANDN U1557 ( .B(n889), .A(n27216), .Z(n890) );
  OR U1558 ( .A(n27217), .B(n890), .Z(n891) );
  AND U1559 ( .A(n27218), .B(n891), .Z(n892) );
  ANDN U1560 ( .B(n24336), .A(n24335), .Z(n893) );
  OR U1561 ( .A(n892), .B(n27219), .Z(n894) );
  AND U1562 ( .A(n893), .B(n894), .Z(n27221) );
  NAND U1563 ( .A(n27249), .B(n24329), .Z(n895) );
  NANDN U1564 ( .A(n27250), .B(n895), .Z(n896) );
  NAND U1565 ( .A(n27251), .B(n896), .Z(n897) );
  NANDN U1566 ( .A(n24328), .B(n897), .Z(n898) );
  NAND U1567 ( .A(n27252), .B(n898), .Z(n899) );
  AND U1568 ( .A(n27253), .B(n899), .Z(n900) );
  OR U1569 ( .A(n27254), .B(n900), .Z(n901) );
  NAND U1570 ( .A(n27255), .B(n901), .Z(n902) );
  NANDN U1571 ( .A(n27256), .B(n902), .Z(n903) );
  NAND U1572 ( .A(n27257), .B(n903), .Z(n904) );
  NANDN U1573 ( .A(n27258), .B(n904), .Z(n905) );
  AND U1574 ( .A(n27259), .B(n905), .Z(n906) );
  OR U1575 ( .A(n27260), .B(n906), .Z(n907) );
  NAND U1576 ( .A(n27261), .B(n907), .Z(n908) );
  NANDN U1577 ( .A(n27262), .B(n908), .Z(n909) );
  AND U1578 ( .A(n27263), .B(n909), .Z(n27265) );
  NAND U1579 ( .A(n27292), .B(n27293), .Z(n910) );
  NAND U1580 ( .A(n24321), .B(n910), .Z(n911) );
  NANDN U1581 ( .A(n27294), .B(n911), .Z(n912) );
  NAND U1582 ( .A(n27295), .B(n912), .Z(n913) );
  NANDN U1583 ( .A(n24320), .B(n913), .Z(n914) );
  AND U1584 ( .A(n27296), .B(n914), .Z(n915) );
  NANDN U1585 ( .A(n915), .B(n27297), .Z(n916) );
  NAND U1586 ( .A(n27298), .B(n916), .Z(n917) );
  NANDN U1587 ( .A(n27299), .B(n917), .Z(n918) );
  NAND U1588 ( .A(n27300), .B(n918), .Z(n919) );
  NANDN U1589 ( .A(n27301), .B(n919), .Z(n920) );
  AND U1590 ( .A(n27302), .B(n920), .Z(n921) );
  OR U1591 ( .A(n27303), .B(n921), .Z(n922) );
  NAND U1592 ( .A(n27304), .B(n922), .Z(n923) );
  NAND U1593 ( .A(n27305), .B(n923), .Z(n924) );
  NANDN U1594 ( .A(n27306), .B(n924), .Z(n27308) );
  NAND U1595 ( .A(n27344), .B(n27343), .Z(n925) );
  ANDN U1596 ( .B(n925), .A(n27345), .Z(n926) );
  NANDN U1597 ( .A(n926), .B(n27346), .Z(n927) );
  NANDN U1598 ( .A(n27347), .B(n927), .Z(n928) );
  NAND U1599 ( .A(n27348), .B(n928), .Z(n929) );
  NAND U1600 ( .A(n27350), .B(n27349), .Z(n930) );
  NANDN U1601 ( .A(n929), .B(n930), .Z(n931) );
  ANDN U1602 ( .B(n931), .A(n27351), .Z(n932) );
  NANDN U1603 ( .A(n932), .B(n27352), .Z(n933) );
  NANDN U1604 ( .A(n27353), .B(n933), .Z(n934) );
  NANDN U1605 ( .A(n27354), .B(n934), .Z(n935) );
  NAND U1606 ( .A(n27355), .B(n935), .Z(n936) );
  NANDN U1607 ( .A(n24314), .B(n936), .Z(n937) );
  AND U1608 ( .A(n27356), .B(n937), .Z(n938) );
  OR U1609 ( .A(n938), .B(n27357), .Z(n939) );
  ANDN U1610 ( .B(n939), .A(n27358), .Z(n27360) );
  ANDN U1611 ( .B(n13024), .A(n13023), .Z(n27383) );
  ANDN U1612 ( .B(n27400), .A(n27404), .Z(n940) );
  NAND U1613 ( .A(n27401), .B(n940), .Z(n941) );
  AND U1614 ( .A(n27405), .B(n941), .Z(n942) );
  OR U1615 ( .A(n942), .B(n27406), .Z(n943) );
  NAND U1616 ( .A(n27407), .B(n943), .Z(n944) );
  NANDN U1617 ( .A(n27408), .B(n944), .Z(n945) );
  NAND U1618 ( .A(n24306), .B(n24305), .Z(n946) );
  NANDN U1619 ( .A(n945), .B(n946), .Z(n947) );
  AND U1620 ( .A(n27409), .B(n947), .Z(n948) );
  OR U1621 ( .A(n948), .B(n27410), .Z(n949) );
  NAND U1622 ( .A(n24304), .B(n949), .Z(n950) );
  NANDN U1623 ( .A(n27411), .B(n950), .Z(n951) );
  NANDN U1624 ( .A(n27412), .B(n951), .Z(n952) );
  NAND U1625 ( .A(n27413), .B(n952), .Z(n953) );
  ANDN U1626 ( .B(n953), .A(n27414), .Z(n954) );
  NANDN U1627 ( .A(n954), .B(n27415), .Z(n955) );
  NANDN U1628 ( .A(n27416), .B(n955), .Z(n956) );
  NAND U1629 ( .A(n27417), .B(n956), .Z(n27418) );
  ANDN U1630 ( .B(n12985), .A(n12984), .Z(n27432) );
  ANDN U1631 ( .B(n12970), .A(n12969), .Z(n24292) );
  NAND U1632 ( .A(n27470), .B(n27469), .Z(n957) );
  NAND U1633 ( .A(n27472), .B(n957), .Z(n958) );
  AND U1634 ( .A(n27473), .B(n958), .Z(n959) );
  OR U1635 ( .A(n27474), .B(n959), .Z(n960) );
  NAND U1636 ( .A(n27475), .B(n960), .Z(n961) );
  NAND U1637 ( .A(n27476), .B(n961), .Z(n962) );
  NAND U1638 ( .A(n27477), .B(n962), .Z(n963) );
  NANDN U1639 ( .A(n27478), .B(n963), .Z(n964) );
  AND U1640 ( .A(n27479), .B(n964), .Z(n965) );
  NANDN U1641 ( .A(n965), .B(n27480), .Z(n966) );
  NANDN U1642 ( .A(n27481), .B(n966), .Z(n967) );
  NAND U1643 ( .A(n27482), .B(n967), .Z(n968) );
  NAND U1644 ( .A(n27483), .B(n968), .Z(n969) );
  AND U1645 ( .A(n27484), .B(n969), .Z(n970) );
  NAND U1646 ( .A(n970), .B(n27485), .Z(n971) );
  AND U1647 ( .A(n27487), .B(n27486), .Z(n972) );
  NAND U1648 ( .A(n971), .B(n972), .Z(n973) );
  NAND U1649 ( .A(n27488), .B(n973), .Z(n27490) );
  NANDN U1650 ( .A(n24286), .B(n27519), .Z(n974) );
  NAND U1651 ( .A(n24285), .B(n974), .Z(n975) );
  ANDN U1652 ( .B(n975), .A(n27520), .Z(n976) );
  NANDN U1653 ( .A(n976), .B(n27521), .Z(n977) );
  NANDN U1654 ( .A(n24284), .B(n977), .Z(n978) );
  NAND U1655 ( .A(n27522), .B(n978), .Z(n979) );
  NAND U1656 ( .A(n27523), .B(n979), .Z(n980) );
  NAND U1657 ( .A(n27524), .B(n980), .Z(n981) );
  AND U1658 ( .A(n27525), .B(n981), .Z(n982) );
  OR U1659 ( .A(n27526), .B(n982), .Z(n983) );
  NAND U1660 ( .A(n27527), .B(n983), .Z(n984) );
  NANDN U1661 ( .A(n24283), .B(n984), .Z(n985) );
  NAND U1662 ( .A(n24282), .B(n985), .Z(n27529) );
  ANDN U1663 ( .B(n12887), .A(n12886), .Z(n27549) );
  OR U1664 ( .A(n27571), .B(n27572), .Z(n986) );
  NAND U1665 ( .A(n27573), .B(n986), .Z(n987) );
  NAND U1666 ( .A(n24273), .B(n987), .Z(n988) );
  NANDN U1667 ( .A(n27574), .B(n988), .Z(n989) );
  NAND U1668 ( .A(n27575), .B(n989), .Z(n990) );
  ANDN U1669 ( .B(n990), .A(n24272), .Z(n991) );
  NANDN U1670 ( .A(n991), .B(n24271), .Z(n992) );
  NAND U1671 ( .A(n27576), .B(n992), .Z(n993) );
  NAND U1672 ( .A(n27577), .B(n993), .Z(n994) );
  NAND U1673 ( .A(n27578), .B(n994), .Z(n995) );
  NAND U1674 ( .A(n27579), .B(n995), .Z(n996) );
  ANDN U1675 ( .B(n996), .A(n27580), .Z(n997) );
  NANDN U1676 ( .A(n997), .B(n27581), .Z(n998) );
  NANDN U1677 ( .A(n27582), .B(n998), .Z(n999) );
  NAND U1678 ( .A(n27583), .B(n999), .Z(n27585) );
  NANDN U1679 ( .A(n12833), .B(n12834), .Z(n27601) );
  OR U1680 ( .A(n27628), .B(n27629), .Z(n1000) );
  NAND U1681 ( .A(n27630), .B(n1000), .Z(n1001) );
  NAND U1682 ( .A(n27631), .B(n1001), .Z(n1002) );
  NANDN U1683 ( .A(n27632), .B(n1002), .Z(n1003) );
  NAND U1684 ( .A(n27633), .B(n1003), .Z(n1004) );
  AND U1685 ( .A(n27634), .B(n1004), .Z(n1005) );
  OR U1686 ( .A(n27635), .B(n1005), .Z(n1006) );
  NAND U1687 ( .A(n27636), .B(n1006), .Z(n1007) );
  NAND U1688 ( .A(n27637), .B(n1007), .Z(n1008) );
  NANDN U1689 ( .A(n27638), .B(n1008), .Z(n1009) );
  NAND U1690 ( .A(n27639), .B(n1009), .Z(n1010) );
  AND U1691 ( .A(n27640), .B(n1010), .Z(n1011) );
  NANDN U1692 ( .A(n1011), .B(n27641), .Z(n1012) );
  NAND U1693 ( .A(n27642), .B(n1012), .Z(n1013) );
  NANDN U1694 ( .A(n27643), .B(n1013), .Z(n1014) );
  NAND U1695 ( .A(n27644), .B(n1014), .Z(n1015) );
  NANDN U1696 ( .A(n27645), .B(n1015), .Z(n1016) );
  AND U1697 ( .A(n27646), .B(n1016), .Z(n27649) );
  NANDN U1698 ( .A(n19374), .B(n19375), .Z(n1017) );
  NAND U1699 ( .A(n19376), .B(n1017), .Z(n24257) );
  ANDN U1700 ( .B(n27675), .A(n12780), .Z(n27674) );
  ANDN U1701 ( .B(n12749), .A(n12748), .Z(n27727) );
  NANDN U1702 ( .A(n27745), .B(n27744), .Z(n1018) );
  NAND U1703 ( .A(n27746), .B(n1018), .Z(n1019) );
  ANDN U1704 ( .B(n1019), .A(n27747), .Z(n1020) );
  NANDN U1705 ( .A(n1020), .B(n27748), .Z(n1021) );
  NAND U1706 ( .A(n27749), .B(n1021), .Z(n1022) );
  NAND U1707 ( .A(n27750), .B(n1022), .Z(n1023) );
  NANDN U1708 ( .A(n27751), .B(n1023), .Z(n1024) );
  NAND U1709 ( .A(n27752), .B(n1024), .Z(n1025) );
  ANDN U1710 ( .B(n1025), .A(n27753), .Z(n1026) );
  NANDN U1711 ( .A(n1026), .B(n27754), .Z(n1027) );
  NANDN U1712 ( .A(n27755), .B(n1027), .Z(n1028) );
  NANDN U1713 ( .A(n27756), .B(n1028), .Z(n1029) );
  NAND U1714 ( .A(n27757), .B(n1029), .Z(n1030) );
  NAND U1715 ( .A(n27758), .B(n1030), .Z(n1031) );
  AND U1716 ( .A(n27759), .B(n1031), .Z(n1032) );
  NANDN U1717 ( .A(n1032), .B(n27760), .Z(n1033) );
  NAND U1718 ( .A(n27761), .B(n1033), .Z(n1034) );
  NAND U1719 ( .A(n27762), .B(n1034), .Z(n1035) );
  NANDN U1720 ( .A(n27763), .B(n1035), .Z(n27764) );
  NAND U1721 ( .A(n24247), .B(n24248), .Z(n1036) );
  NAND U1722 ( .A(n27796), .B(n27797), .Z(n1037) );
  NAND U1723 ( .A(n1036), .B(n1037), .Z(n1038) );
  OR U1724 ( .A(n1038), .B(n27798), .Z(n1039) );
  NAND U1725 ( .A(n27799), .B(n1039), .Z(n1040) );
  NANDN U1726 ( .A(n27800), .B(n1040), .Z(n1041) );
  AND U1727 ( .A(n27801), .B(n24246), .Z(n1042) );
  NAND U1728 ( .A(n1041), .B(n1042), .Z(n1043) );
  NANDN U1729 ( .A(n24245), .B(n1043), .Z(n1044) );
  NANDN U1730 ( .A(n27802), .B(n1044), .Z(n1045) );
  NANDN U1731 ( .A(n27803), .B(n1045), .Z(n1046) );
  AND U1732 ( .A(n27804), .B(n1046), .Z(n1047) );
  OR U1733 ( .A(n27805), .B(n1047), .Z(n1048) );
  NAND U1734 ( .A(n27806), .B(n1048), .Z(n1049) );
  NANDN U1735 ( .A(n27807), .B(n1049), .Z(n27808) );
  NAND U1736 ( .A(n27838), .B(n27839), .Z(n1050) );
  NANDN U1737 ( .A(n27840), .B(n1050), .Z(n1051) );
  ANDN U1738 ( .B(n1051), .A(n24238), .Z(n1052) );
  NANDN U1739 ( .A(n1052), .B(n27841), .Z(n1053) );
  NAND U1740 ( .A(n27842), .B(n1053), .Z(n1054) );
  NANDN U1741 ( .A(n27843), .B(n1054), .Z(n1055) );
  NAND U1742 ( .A(n27844), .B(n1055), .Z(n1056) );
  NANDN U1743 ( .A(n27845), .B(n1056), .Z(n1057) );
  AND U1744 ( .A(n27846), .B(n1057), .Z(n1058) );
  OR U1745 ( .A(n27847), .B(n1058), .Z(n1059) );
  AND U1746 ( .A(n27848), .B(n1059), .Z(n1060) );
  ANDN U1747 ( .B(n27851), .A(n1060), .Z(n1061) );
  OR U1748 ( .A(n27850), .B(n27849), .Z(n1062) );
  NAND U1749 ( .A(n1061), .B(n1062), .Z(n1063) );
  NAND U1750 ( .A(n27852), .B(n1063), .Z(n1064) );
  NANDN U1751 ( .A(n27853), .B(n1064), .Z(n1065) );
  AND U1752 ( .A(n27854), .B(n1065), .Z(n1066) );
  OR U1753 ( .A(n27855), .B(n1066), .Z(n1067) );
  AND U1754 ( .A(n27856), .B(n1067), .Z(n27857) );
  NANDN U1755 ( .A(n27896), .B(n27897), .Z(n1068) );
  NAND U1756 ( .A(n27898), .B(n1068), .Z(n1069) );
  NANDN U1757 ( .A(n27899), .B(n1069), .Z(n1070) );
  NAND U1758 ( .A(n27900), .B(n1070), .Z(n1071) );
  NANDN U1759 ( .A(n27901), .B(n1071), .Z(n1072) );
  ANDN U1760 ( .B(n1072), .A(n27902), .Z(n1073) );
  NANDN U1761 ( .A(n1073), .B(n27903), .Z(n1074) );
  NANDN U1762 ( .A(n27904), .B(n1074), .Z(n1075) );
  NANDN U1763 ( .A(n27905), .B(n1075), .Z(n1076) );
  NAND U1764 ( .A(n27906), .B(n1076), .Z(n1077) );
  NAND U1765 ( .A(n27907), .B(n1077), .Z(n1078) );
  ANDN U1766 ( .B(n1078), .A(n27908), .Z(n1079) );
  NANDN U1767 ( .A(n1079), .B(n27909), .Z(n1080) );
  NAND U1768 ( .A(n27910), .B(n1080), .Z(n1081) );
  NANDN U1769 ( .A(n24236), .B(n1081), .Z(n1082) );
  NAND U1770 ( .A(n24235), .B(n1082), .Z(n27911) );
  NANDN U1771 ( .A(n27935), .B(n27934), .Z(n1083) );
  NAND U1772 ( .A(n27936), .B(n1083), .Z(n1084) );
  NANDN U1773 ( .A(n27937), .B(n1084), .Z(n1085) );
  NAND U1774 ( .A(n27938), .B(n1085), .Z(n1086) );
  NANDN U1775 ( .A(n27939), .B(n1086), .Z(n1087) );
  AND U1776 ( .A(n27940), .B(n1087), .Z(n1088) );
  NAND U1777 ( .A(n27941), .B(n27942), .Z(n1089) );
  NAND U1778 ( .A(n1088), .B(n1089), .Z(n1090) );
  NANDN U1779 ( .A(n27943), .B(n1090), .Z(n1091) );
  NAND U1780 ( .A(n27944), .B(n1091), .Z(n1092) );
  NAND U1781 ( .A(n27945), .B(n1092), .Z(n1093) );
  AND U1782 ( .A(n27946), .B(n1093), .Z(n1094) );
  OR U1783 ( .A(n27947), .B(n1094), .Z(n1095) );
  AND U1784 ( .A(n27948), .B(n1095), .Z(n1096) );
  OR U1785 ( .A(n27949), .B(n1096), .Z(n1097) );
  NAND U1786 ( .A(n27950), .B(n1097), .Z(n1098) );
  NANDN U1787 ( .A(n27951), .B(n1098), .Z(n27952) );
  NAND U1788 ( .A(n27980), .B(n24218), .Z(n1099) );
  NANDN U1789 ( .A(n27981), .B(n1099), .Z(n1100) );
  AND U1790 ( .A(n27982), .B(n1100), .Z(n1101) );
  OR U1791 ( .A(n27983), .B(n1101), .Z(n1102) );
  NAND U1792 ( .A(n27984), .B(n1102), .Z(n1103) );
  NAND U1793 ( .A(n24217), .B(n1103), .Z(n1104) );
  NAND U1794 ( .A(n27985), .B(n1104), .Z(n1105) );
  NAND U1795 ( .A(n27986), .B(n1105), .Z(n1106) );
  AND U1796 ( .A(n27987), .B(n1106), .Z(n1107) );
  NANDN U1797 ( .A(n1107), .B(n27988), .Z(n1108) );
  ANDN U1798 ( .B(n1108), .A(n27989), .Z(n1109) );
  NANDN U1799 ( .A(n1109), .B(n27990), .Z(n1110) );
  NAND U1800 ( .A(n27991), .B(n1110), .Z(n1111) );
  NANDN U1801 ( .A(n27992), .B(n1111), .Z(n27993) );
  ANDN U1802 ( .B(n12551), .A(n12550), .Z(n28008) );
  NANDN U1803 ( .A(n28041), .B(n28040), .Z(n1112) );
  NAND U1804 ( .A(n24202), .B(n1112), .Z(n1113) );
  ANDN U1805 ( .B(n1113), .A(n28042), .Z(n1114) );
  NANDN U1806 ( .A(n1114), .B(n28043), .Z(n1115) );
  NANDN U1807 ( .A(n24201), .B(n1115), .Z(n1116) );
  NAND U1808 ( .A(n28044), .B(n1116), .Z(n1117) );
  NANDN U1809 ( .A(n28045), .B(n1117), .Z(n1118) );
  NAND U1810 ( .A(n28046), .B(n1118), .Z(n1119) );
  ANDN U1811 ( .B(n1119), .A(n28047), .Z(n1120) );
  NANDN U1812 ( .A(n1120), .B(n28048), .Z(n1121) );
  NAND U1813 ( .A(n28049), .B(n1121), .Z(n1122) );
  NAND U1814 ( .A(n28050), .B(n1122), .Z(n1123) );
  NANDN U1815 ( .A(n28051), .B(n1123), .Z(n1124) );
  NAND U1816 ( .A(n28052), .B(n1124), .Z(n1125) );
  ANDN U1817 ( .B(n1125), .A(n28053), .Z(n28054) );
  ANDN U1818 ( .B(n12508), .A(n12507), .Z(n28079) );
  NAND U1819 ( .A(n28105), .B(n28104), .Z(n1126) );
  NAND U1820 ( .A(n28106), .B(n1126), .Z(n1127) );
  ANDN U1821 ( .B(n1127), .A(n28107), .Z(n1128) );
  NANDN U1822 ( .A(n1128), .B(n28108), .Z(n1129) );
  NANDN U1823 ( .A(n24196), .B(n1129), .Z(n1130) );
  NANDN U1824 ( .A(n28109), .B(n1130), .Z(n1131) );
  NAND U1825 ( .A(n28110), .B(n1131), .Z(n1132) );
  NANDN U1826 ( .A(n28111), .B(n1132), .Z(n1133) );
  AND U1827 ( .A(n28112), .B(n1133), .Z(n1134) );
  NAND U1828 ( .A(n24194), .B(n24193), .Z(n1135) );
  AND U1829 ( .A(n24195), .B(n1135), .Z(n1136) );
  OR U1830 ( .A(n28113), .B(n1134), .Z(n1137) );
  NAND U1831 ( .A(n1136), .B(n1137), .Z(n1138) );
  NANDN U1832 ( .A(n28114), .B(n1138), .Z(n1139) );
  ANDN U1833 ( .B(n1139), .A(n28115), .Z(n28117) );
  NAND U1834 ( .A(n28142), .B(n28141), .Z(n1140) );
  NANDN U1835 ( .A(n28143), .B(n1140), .Z(n1141) );
  NANDN U1836 ( .A(n28144), .B(n1141), .Z(n1142) );
  NAND U1837 ( .A(n28145), .B(n1142), .Z(n1143) );
  NANDN U1838 ( .A(n24181), .B(n1143), .Z(n1144) );
  AND U1839 ( .A(n24180), .B(n1144), .Z(n1145) );
  NAND U1840 ( .A(n1145), .B(n28146), .Z(n1146) );
  NAND U1841 ( .A(n28147), .B(n1146), .Z(n1147) );
  AND U1842 ( .A(n28148), .B(n1147), .Z(n1148) );
  OR U1843 ( .A(n28149), .B(n1148), .Z(n1149) );
  AND U1844 ( .A(n28150), .B(n1149), .Z(n1150) );
  NANDN U1845 ( .A(n24179), .B(n24178), .Z(n1151) );
  NAND U1846 ( .A(n1150), .B(n1151), .Z(n1152) );
  NAND U1847 ( .A(n28151), .B(n1152), .Z(n28152) );
  NANDN U1848 ( .A(x[2752]), .B(y[2752]), .Z(n1153) );
  NANDN U1849 ( .A(n12437), .B(n1153), .Z(n28168) );
  NAND U1850 ( .A(n12421), .B(n12420), .Z(n1154) );
  ANDN U1851 ( .B(n1154), .A(n12422), .Z(n28191) );
  ANDN U1852 ( .B(n12405), .A(n12404), .Z(n28213) );
  NANDN U1853 ( .A(n28241), .B(n28242), .Z(n1155) );
  NANDN U1854 ( .A(n28243), .B(n1155), .Z(n1156) );
  NAND U1855 ( .A(n28244), .B(n1156), .Z(n1157) );
  NANDN U1856 ( .A(n28245), .B(n1157), .Z(n1158) );
  NAND U1857 ( .A(n28246), .B(n1158), .Z(n1159) );
  AND U1858 ( .A(n28247), .B(n1159), .Z(n1160) );
  ANDN U1859 ( .B(n28250), .A(n1160), .Z(n1161) );
  NANDN U1860 ( .A(n28248), .B(n28249), .Z(n1162) );
  NAND U1861 ( .A(n1161), .B(n1162), .Z(n1163) );
  NAND U1862 ( .A(n28251), .B(n1163), .Z(n1164) );
  NAND U1863 ( .A(n28252), .B(n1164), .Z(n1165) );
  ANDN U1864 ( .B(n1165), .A(n24152), .Z(n1166) );
  NANDN U1865 ( .A(n1166), .B(n28253), .Z(n1167) );
  NANDN U1866 ( .A(n28254), .B(n1167), .Z(n1168) );
  NANDN U1867 ( .A(n28255), .B(n1168), .Z(n28256) );
  NANDN U1868 ( .A(n28312), .B(n28313), .Z(n1169) );
  NANDN U1869 ( .A(n28314), .B(n1169), .Z(n1170) );
  AND U1870 ( .A(n28315), .B(n1170), .Z(n1171) );
  OR U1871 ( .A(n1171), .B(n28316), .Z(n1172) );
  NAND U1872 ( .A(n28317), .B(n1172), .Z(n1173) );
  AND U1873 ( .A(n28318), .B(n1173), .Z(n1174) );
  OR U1874 ( .A(n1174), .B(n28319), .Z(n1175) );
  NAND U1875 ( .A(n28320), .B(n1175), .Z(n1176) );
  ANDN U1876 ( .B(n1176), .A(n28321), .Z(n1177) );
  NANDN U1877 ( .A(n1177), .B(n28322), .Z(n1178) );
  NANDN U1878 ( .A(n28323), .B(n1178), .Z(n1179) );
  NAND U1879 ( .A(n28324), .B(n1179), .Z(n1180) );
  NANDN U1880 ( .A(n28325), .B(n1180), .Z(n1181) );
  NAND U1881 ( .A(n24149), .B(n1181), .Z(n1182) );
  ANDN U1882 ( .B(n1182), .A(n28326), .Z(n1183) );
  OR U1883 ( .A(n1183), .B(n28327), .Z(n1184) );
  NAND U1884 ( .A(n28328), .B(n1184), .Z(n1185) );
  NANDN U1885 ( .A(n28329), .B(n1185), .Z(n28330) );
  OR U1886 ( .A(n28359), .B(n28360), .Z(n1186) );
  NAND U1887 ( .A(n28362), .B(n1186), .Z(n1187) );
  NANDN U1888 ( .A(n28363), .B(n1187), .Z(n1188) );
  NANDN U1889 ( .A(n28364), .B(n1188), .Z(n1189) );
  NAND U1890 ( .A(n28365), .B(n1189), .Z(n1190) );
  AND U1891 ( .A(n28366), .B(n1190), .Z(n1191) );
  NANDN U1892 ( .A(n1191), .B(n28367), .Z(n1192) );
  ANDN U1893 ( .B(n1192), .A(n28368), .Z(n1193) );
  ANDN U1894 ( .B(n28371), .A(n28370), .Z(n1194) );
  NANDN U1895 ( .A(n1193), .B(n28369), .Z(n1195) );
  AND U1896 ( .A(n1194), .B(n1195), .Z(n1196) );
  ANDN U1897 ( .B(n24142), .A(n1196), .Z(n1197) );
  NANDN U1898 ( .A(n28372), .B(n28373), .Z(n1198) );
  NAND U1899 ( .A(n1197), .B(n1198), .Z(n1199) );
  NANDN U1900 ( .A(n24141), .B(n1199), .Z(n28374) );
  NAND U1901 ( .A(n28401), .B(n24132), .Z(n1200) );
  NANDN U1902 ( .A(n28402), .B(n1200), .Z(n1201) );
  NAND U1903 ( .A(n28403), .B(n1201), .Z(n1202) );
  NANDN U1904 ( .A(n28404), .B(n1202), .Z(n1203) );
  NAND U1905 ( .A(n28405), .B(n1203), .Z(n1204) );
  AND U1906 ( .A(n28406), .B(n1204), .Z(n1205) );
  OR U1907 ( .A(n28407), .B(n1205), .Z(n1206) );
  AND U1908 ( .A(n28408), .B(n1206), .Z(n1207) );
  NOR U1909 ( .A(n1207), .B(n24131), .Z(n1208) );
  OR U1910 ( .A(n24129), .B(n24130), .Z(n1209) );
  AND U1911 ( .A(n1208), .B(n1209), .Z(n1210) );
  NANDN U1912 ( .A(n1210), .B(n28409), .Z(n1211) );
  NANDN U1913 ( .A(n28410), .B(n1211), .Z(n1212) );
  NAND U1914 ( .A(n28411), .B(n1212), .Z(n1213) );
  NANDN U1915 ( .A(n24128), .B(n1213), .Z(n28412) );
  AND U1916 ( .A(n28443), .B(n28442), .Z(n1214) );
  OR U1917 ( .A(n24121), .B(n24122), .Z(n1215) );
  NANDN U1918 ( .A(n28444), .B(n1214), .Z(n1216) );
  NAND U1919 ( .A(n1215), .B(n1216), .Z(n1217) );
  AND U1920 ( .A(n28446), .B(n28447), .Z(n1218) );
  NANDN U1921 ( .A(n1217), .B(n28445), .Z(n1219) );
  AND U1922 ( .A(n1218), .B(n1219), .Z(n1220) );
  NANDN U1923 ( .A(n1220), .B(n28448), .Z(n1221) );
  NANDN U1924 ( .A(n28449), .B(n1221), .Z(n1222) );
  NAND U1925 ( .A(n28450), .B(n1222), .Z(n1223) );
  NANDN U1926 ( .A(n24120), .B(n1223), .Z(n1224) );
  NAND U1927 ( .A(n24119), .B(n1224), .Z(n1225) );
  ANDN U1928 ( .B(n1225), .A(n28451), .Z(n1226) );
  NANDN U1929 ( .A(n1226), .B(n28452), .Z(n1227) );
  NAND U1930 ( .A(n28453), .B(n1227), .Z(n1228) );
  NAND U1931 ( .A(n28454), .B(n1228), .Z(n1229) );
  NANDN U1932 ( .A(n28455), .B(n1229), .Z(n28456) );
  NANDN U1933 ( .A(n24110), .B(n28486), .Z(n1230) );
  NAND U1934 ( .A(n28487), .B(n1230), .Z(n1231) );
  AND U1935 ( .A(n28488), .B(n1231), .Z(n1232) );
  OR U1936 ( .A(n28489), .B(n1232), .Z(n1233) );
  AND U1937 ( .A(n28490), .B(n1233), .Z(n1234) );
  OR U1938 ( .A(n28491), .B(n28492), .Z(n1235) );
  NAND U1939 ( .A(n1234), .B(n1235), .Z(n1236) );
  NANDN U1940 ( .A(n28493), .B(n1236), .Z(n1237) );
  NAND U1941 ( .A(n28494), .B(n1237), .Z(n1238) );
  NANDN U1942 ( .A(n28495), .B(n1238), .Z(n1239) );
  AND U1943 ( .A(n24109), .B(n1239), .Z(n1240) );
  OR U1944 ( .A(n28496), .B(n1240), .Z(n1241) );
  AND U1945 ( .A(n28497), .B(n1241), .Z(n1242) );
  NANDN U1946 ( .A(n1242), .B(n28498), .Z(n1243) );
  NANDN U1947 ( .A(n28499), .B(n1243), .Z(n1244) );
  NAND U1948 ( .A(n28500), .B(n1244), .Z(n28501) );
  NOR U1949 ( .A(n12177), .B(n12178), .Z(n28526) );
  NAND U1950 ( .A(n28543), .B(n24095), .Z(n1245) );
  NANDN U1951 ( .A(n28544), .B(n1245), .Z(n1246) );
  NAND U1952 ( .A(n28545), .B(n1246), .Z(n1247) );
  NAND U1953 ( .A(n28546), .B(n1247), .Z(n1248) );
  NAND U1954 ( .A(n28547), .B(n1248), .Z(n1249) );
  ANDN U1955 ( .B(n1249), .A(n28548), .Z(n1250) );
  NANDN U1956 ( .A(n1250), .B(n28549), .Z(n1251) );
  NANDN U1957 ( .A(n28550), .B(n1251), .Z(n1252) );
  NAND U1958 ( .A(n28551), .B(n1252), .Z(n1253) );
  NAND U1959 ( .A(n28552), .B(n1253), .Z(n1254) );
  NAND U1960 ( .A(n28553), .B(n1254), .Z(n1255) );
  ANDN U1961 ( .B(n1255), .A(n28554), .Z(n1256) );
  OR U1962 ( .A(n1256), .B(n28555), .Z(n1257) );
  NAND U1963 ( .A(n28556), .B(n1257), .Z(n1258) );
  NANDN U1964 ( .A(n28557), .B(n1258), .Z(n1259) );
  AND U1965 ( .A(n28558), .B(n1259), .Z(n28560) );
  NANDN U1966 ( .A(n24090), .B(n28587), .Z(n1260) );
  NAND U1967 ( .A(n24089), .B(n1260), .Z(n1261) );
  NAND U1968 ( .A(n28588), .B(n1261), .Z(n1262) );
  NANDN U1969 ( .A(n28589), .B(n1262), .Z(n1263) );
  NAND U1970 ( .A(n28590), .B(n1263), .Z(n1264) );
  ANDN U1971 ( .B(n1264), .A(n24088), .Z(n1265) );
  NANDN U1972 ( .A(n1265), .B(n28591), .Z(n1266) );
  NANDN U1973 ( .A(n28592), .B(n1266), .Z(n1267) );
  NAND U1974 ( .A(n28593), .B(n1267), .Z(n1268) );
  NAND U1975 ( .A(n28594), .B(n1268), .Z(n1269) );
  NAND U1976 ( .A(n28595), .B(n1269), .Z(n1270) );
  ANDN U1977 ( .B(n1270), .A(n28596), .Z(n1271) );
  NANDN U1978 ( .A(n1271), .B(n28597), .Z(n1272) );
  ANDN U1979 ( .B(n1272), .A(n28598), .Z(n28600) );
  NAND U1980 ( .A(n28629), .B(n28630), .Z(n1273) );
  NAND U1981 ( .A(n28631), .B(n1273), .Z(n1274) );
  NANDN U1982 ( .A(n24082), .B(n1274), .Z(n1275) );
  NAND U1983 ( .A(n24081), .B(n1275), .Z(n1276) );
  NANDN U1984 ( .A(n28632), .B(n1276), .Z(n1277) );
  AND U1985 ( .A(n28633), .B(n1277), .Z(n1278) );
  OR U1986 ( .A(n1278), .B(n28634), .Z(n1279) );
  NAND U1987 ( .A(n28635), .B(n1279), .Z(n1280) );
  ANDN U1988 ( .B(n1280), .A(n28636), .Z(n1281) );
  NANDN U1989 ( .A(n1281), .B(n24080), .Z(n1282) );
  ANDN U1990 ( .B(n1282), .A(n28637), .Z(n1283) );
  NANDN U1991 ( .A(n1283), .B(n28638), .Z(n1284) );
  NAND U1992 ( .A(n28639), .B(n1284), .Z(n1285) );
  NANDN U1993 ( .A(n28640), .B(n1285), .Z(n28641) );
  NANDN U1994 ( .A(n28668), .B(n28667), .Z(n1286) );
  NANDN U1995 ( .A(n28669), .B(n1286), .Z(n1287) );
  AND U1996 ( .A(n28670), .B(n1287), .Z(n1288) );
  OR U1997 ( .A(n24071), .B(n1288), .Z(n1289) );
  NAND U1998 ( .A(n24070), .B(n1289), .Z(n1290) );
  NANDN U1999 ( .A(n28671), .B(n1290), .Z(n1291) );
  NAND U2000 ( .A(n28672), .B(n1291), .Z(n1292) );
  NAND U2001 ( .A(n28673), .B(n1292), .Z(n1293) );
  ANDN U2002 ( .B(n1293), .A(n24069), .Z(n1294) );
  NANDN U2003 ( .A(n1294), .B(n24068), .Z(n1295) );
  NANDN U2004 ( .A(n28674), .B(n1295), .Z(n1296) );
  NAND U2005 ( .A(n28675), .B(n1296), .Z(n1297) );
  NANDN U2006 ( .A(n28676), .B(n1297), .Z(n28677) );
  NANDN U2007 ( .A(n24059), .B(n28697), .Z(n1298) );
  NAND U2008 ( .A(n24058), .B(n1298), .Z(n1299) );
  NANDN U2009 ( .A(n28698), .B(n1299), .Z(n1300) );
  NAND U2010 ( .A(n28699), .B(n1300), .Z(n1301) );
  NANDN U2011 ( .A(n28700), .B(n1301), .Z(n1302) );
  AND U2012 ( .A(n28701), .B(n1302), .Z(n1303) );
  AND U2013 ( .A(n28704), .B(n28703), .Z(n1304) );
  OR U2014 ( .A(n1303), .B(n28702), .Z(n1305) );
  AND U2015 ( .A(n1304), .B(n1305), .Z(n1306) );
  OR U2016 ( .A(n28705), .B(n1306), .Z(n1307) );
  AND U2017 ( .A(n28706), .B(n1307), .Z(n1308) );
  OR U2018 ( .A(n24057), .B(n1308), .Z(n1309) );
  NAND U2019 ( .A(n24056), .B(n1309), .Z(n1310) );
  NANDN U2020 ( .A(n28707), .B(n1310), .Z(n28708) );
  OR U2021 ( .A(n28734), .B(n28735), .Z(n1311) );
  NANDN U2022 ( .A(n28736), .B(n1311), .Z(n1312) );
  AND U2023 ( .A(n28737), .B(n1312), .Z(n1313) );
  OR U2024 ( .A(n1313), .B(n28738), .Z(n1314) );
  NAND U2025 ( .A(n28739), .B(n1314), .Z(n1315) );
  NANDN U2026 ( .A(n28740), .B(n1315), .Z(n1316) );
  NAND U2027 ( .A(n24048), .B(n1316), .Z(n1317) );
  NANDN U2028 ( .A(n28741), .B(n1317), .Z(n1318) );
  AND U2029 ( .A(n28742), .B(n1318), .Z(n1319) );
  OR U2030 ( .A(n24047), .B(n1319), .Z(n1320) );
  AND U2031 ( .A(n24046), .B(n1320), .Z(n1321) );
  AND U2032 ( .A(n24043), .B(n24044), .Z(n1322) );
  OR U2033 ( .A(n24045), .B(n1321), .Z(n1323) );
  AND U2034 ( .A(n1322), .B(n1323), .Z(n28743) );
  NAND U2035 ( .A(n28772), .B(n28771), .Z(n1324) );
  NAND U2036 ( .A(n28773), .B(n1324), .Z(n1325) );
  ANDN U2037 ( .B(n1325), .A(n24036), .Z(n1326) );
  NANDN U2038 ( .A(n1326), .B(n28774), .Z(n1327) );
  NAND U2039 ( .A(n24035), .B(n1327), .Z(n1328) );
  NANDN U2040 ( .A(n28775), .B(n1328), .Z(n1329) );
  NAND U2041 ( .A(n28776), .B(n1329), .Z(n1330) );
  NANDN U2042 ( .A(n24034), .B(n1330), .Z(n1331) );
  AND U2043 ( .A(n24033), .B(n1331), .Z(n1332) );
  OR U2044 ( .A(n1332), .B(n28777), .Z(n1333) );
  NAND U2045 ( .A(n28778), .B(n1333), .Z(n1334) );
  NANDN U2046 ( .A(n28779), .B(n1334), .Z(n1335) );
  NAND U2047 ( .A(n28780), .B(n1335), .Z(n28781) );
  NAND U2048 ( .A(n28802), .B(n28803), .Z(n1336) );
  NANDN U2049 ( .A(n28804), .B(n1336), .Z(n1337) );
  AND U2050 ( .A(n28805), .B(n1337), .Z(n1338) );
  OR U2051 ( .A(n1338), .B(n28806), .Z(n1339) );
  NAND U2052 ( .A(n28807), .B(n1339), .Z(n1340) );
  ANDN U2053 ( .B(n1340), .A(n28808), .Z(n1341) );
  NANDN U2054 ( .A(n1341), .B(n24022), .Z(n1342) );
  NAND U2055 ( .A(n28809), .B(n1342), .Z(n1343) );
  NANDN U2056 ( .A(n28810), .B(n1343), .Z(n1344) );
  NAND U2057 ( .A(n28811), .B(n1344), .Z(n1345) );
  NANDN U2058 ( .A(n28812), .B(n1345), .Z(n1346) );
  AND U2059 ( .A(n24021), .B(n1346), .Z(n1347) );
  OR U2060 ( .A(n28813), .B(n1347), .Z(n1348) );
  NAND U2061 ( .A(n28814), .B(n1348), .Z(n1349) );
  NAND U2062 ( .A(n28815), .B(n1349), .Z(n1350) );
  NANDN U2063 ( .A(n28816), .B(n1350), .Z(n28817) );
  NAND U2064 ( .A(n28837), .B(n24008), .Z(n1351) );
  NANDN U2065 ( .A(n28838), .B(n1351), .Z(n1352) );
  NAND U2066 ( .A(n28839), .B(n1352), .Z(n1353) );
  NAND U2067 ( .A(n28840), .B(n1353), .Z(n1354) );
  NANDN U2068 ( .A(n28841), .B(n1354), .Z(n1355) );
  AND U2069 ( .A(n24007), .B(n1355), .Z(n1356) );
  OR U2070 ( .A(n28842), .B(n1356), .Z(n1357) );
  NAND U2071 ( .A(n28843), .B(n1357), .Z(n1358) );
  NANDN U2072 ( .A(n24006), .B(n1358), .Z(n1359) );
  NAND U2073 ( .A(n24005), .B(n1359), .Z(n1360) );
  NANDN U2074 ( .A(n28844), .B(n1360), .Z(n1361) );
  AND U2075 ( .A(n28845), .B(n1361), .Z(n28846) );
  AND U2076 ( .A(n23996), .B(n23997), .Z(n1362) );
  OR U2077 ( .A(n28869), .B(n28870), .Z(n1363) );
  AND U2078 ( .A(n1362), .B(n1363), .Z(n1364) );
  OR U2079 ( .A(n28871), .B(n1364), .Z(n1365) );
  NAND U2080 ( .A(n28872), .B(n1365), .Z(n1366) );
  NANDN U2081 ( .A(n23995), .B(n1366), .Z(n1367) );
  NAND U2082 ( .A(n28873), .B(n1367), .Z(n1368) );
  NANDN U2083 ( .A(n23994), .B(n1368), .Z(n1369) );
  AND U2084 ( .A(n28874), .B(n1369), .Z(n1370) );
  NANDN U2085 ( .A(n1370), .B(n28875), .Z(n1371) );
  NANDN U2086 ( .A(n28876), .B(n1371), .Z(n1372) );
  NAND U2087 ( .A(n28877), .B(n1372), .Z(n1373) );
  NAND U2088 ( .A(n28878), .B(n1373), .Z(n1374) );
  NAND U2089 ( .A(n28879), .B(n1374), .Z(n1375) );
  ANDN U2090 ( .B(n1375), .A(n28880), .Z(n1376) );
  NANDN U2091 ( .A(n1376), .B(n28881), .Z(n1377) );
  NANDN U2092 ( .A(n28882), .B(n1377), .Z(n1378) );
  NAND U2093 ( .A(n28883), .B(n1378), .Z(n28884) );
  NAND U2094 ( .A(n28907), .B(n28908), .Z(n1379) );
  NANDN U2095 ( .A(n28909), .B(n1379), .Z(n1380) );
  AND U2096 ( .A(n28910), .B(n1380), .Z(n1381) );
  OR U2097 ( .A(n1381), .B(n28911), .Z(n1382) );
  NAND U2098 ( .A(n23988), .B(n1382), .Z(n1383) );
  NANDN U2099 ( .A(n28912), .B(n1383), .Z(n1384) );
  NAND U2100 ( .A(n28913), .B(n1384), .Z(n1385) );
  NANDN U2101 ( .A(n23987), .B(n1385), .Z(n1386) );
  AND U2102 ( .A(n23986), .B(n1386), .Z(n1387) );
  NANDN U2103 ( .A(n1387), .B(n28914), .Z(n1388) );
  ANDN U2104 ( .B(n1388), .A(n28915), .Z(n1389) );
  NANDN U2105 ( .A(n1389), .B(n28916), .Z(n1390) );
  NANDN U2106 ( .A(n28917), .B(n1390), .Z(n1391) );
  NAND U2107 ( .A(n28918), .B(n1391), .Z(n28919) );
  AND U2108 ( .A(n28941), .B(n23975), .Z(n1392) );
  NAND U2109 ( .A(n23976), .B(n1392), .Z(n1393) );
  AND U2110 ( .A(n28942), .B(n1393), .Z(n1394) );
  ANDN U2111 ( .B(n28943), .A(n1394), .Z(n1395) );
  NAND U2112 ( .A(n28944), .B(n1395), .Z(n1396) );
  ANDN U2113 ( .B(n1396), .A(n28945), .Z(n1397) );
  NANDN U2114 ( .A(n1397), .B(n28946), .Z(n1398) );
  ANDN U2115 ( .B(n1398), .A(n28947), .Z(n1399) );
  NOR U2116 ( .A(n23973), .B(n1399), .Z(n1400) );
  NAND U2117 ( .A(n23974), .B(n1400), .Z(n1401) );
  NANDN U2118 ( .A(n28948), .B(n1401), .Z(n1402) );
  NAND U2119 ( .A(n28949), .B(n1402), .Z(n1403) );
  NANDN U2120 ( .A(n28950), .B(n1403), .Z(n1404) );
  AND U2121 ( .A(n28951), .B(n1404), .Z(n1405) );
  OR U2122 ( .A(n28952), .B(n1405), .Z(n1406) );
  NAND U2123 ( .A(n28953), .B(n1406), .Z(n1407) );
  NANDN U2124 ( .A(n28954), .B(n1407), .Z(n1408) );
  NAND U2125 ( .A(n28955), .B(n1408), .Z(n28956) );
  NAND U2126 ( .A(n28988), .B(n28989), .Z(n1409) );
  NANDN U2127 ( .A(n28990), .B(n1409), .Z(n1410) );
  NAND U2128 ( .A(n28991), .B(n1410), .Z(n1411) );
  NAND U2129 ( .A(n28992), .B(n1411), .Z(n1412) );
  NANDN U2130 ( .A(n28993), .B(n1412), .Z(n1413) );
  AND U2131 ( .A(n28994), .B(n1413), .Z(n1414) );
  OR U2132 ( .A(n1414), .B(n28995), .Z(n1415) );
  NAND U2133 ( .A(n28996), .B(n1415), .Z(n1416) );
  NANDN U2134 ( .A(n28997), .B(n1416), .Z(n1417) );
  NAND U2135 ( .A(n28998), .B(n1417), .Z(n1418) );
  NANDN U2136 ( .A(n28999), .B(n1418), .Z(n1419) );
  AND U2137 ( .A(n29000), .B(n1419), .Z(n1420) );
  OR U2138 ( .A(n1420), .B(n29001), .Z(n1421) );
  AND U2139 ( .A(n29002), .B(n1421), .Z(n1422) );
  OR U2140 ( .A(n29003), .B(n1422), .Z(n1423) );
  NAND U2141 ( .A(n29004), .B(n1423), .Z(n1424) );
  NAND U2142 ( .A(n29005), .B(n1424), .Z(n29006) );
  NAND U2143 ( .A(n29034), .B(n29033), .Z(n1425) );
  NANDN U2144 ( .A(n29035), .B(n1425), .Z(n1426) );
  NAND U2145 ( .A(n29036), .B(n1426), .Z(n1427) );
  OR U2146 ( .A(n1427), .B(n23961), .Z(n1428) );
  NANDN U2147 ( .A(n29037), .B(n1428), .Z(n1429) );
  NANDN U2148 ( .A(n29038), .B(n1429), .Z(n1430) );
  OR U2149 ( .A(n1430), .B(n29039), .Z(n1431) );
  NANDN U2150 ( .A(n29040), .B(n1431), .Z(n1432) );
  NAND U2151 ( .A(n29041), .B(n1432), .Z(n1433) );
  NANDN U2152 ( .A(n29042), .B(n1433), .Z(n1434) );
  NAND U2153 ( .A(n29043), .B(n1434), .Z(n1435) );
  ANDN U2154 ( .B(n1435), .A(n29044), .Z(n1436) );
  ANDN U2155 ( .B(n29046), .A(n1436), .Z(n1437) );
  NAND U2156 ( .A(n29045), .B(n1437), .Z(n1438) );
  ANDN U2157 ( .B(n1438), .A(n29047), .Z(n1439) );
  NANDN U2158 ( .A(n1439), .B(n29048), .Z(n1440) );
  ANDN U2159 ( .B(n1440), .A(n29049), .Z(n29053) );
  NAND U2160 ( .A(n29079), .B(n29078), .Z(n1441) );
  NAND U2161 ( .A(n23952), .B(n1441), .Z(n1442) );
  ANDN U2162 ( .B(n1442), .A(n29080), .Z(n1443) );
  NANDN U2163 ( .A(n1443), .B(n29081), .Z(n1444) );
  AND U2164 ( .A(n29082), .B(n1444), .Z(n1445) );
  AND U2165 ( .A(n29085), .B(n29084), .Z(n1446) );
  OR U2166 ( .A(n29083), .B(n1445), .Z(n1447) );
  AND U2167 ( .A(n1446), .B(n1447), .Z(n1448) );
  ANDN U2168 ( .B(n29086), .A(n29087), .Z(n1449) );
  OR U2169 ( .A(n23951), .B(n1448), .Z(n1450) );
  AND U2170 ( .A(n1449), .B(n1450), .Z(n1451) );
  AND U2171 ( .A(n23949), .B(n23950), .Z(n1452) );
  NANDN U2172 ( .A(n1451), .B(n29088), .Z(n1453) );
  AND U2173 ( .A(n1452), .B(n1453), .Z(n29089) );
  NAND U2174 ( .A(n29118), .B(n29119), .Z(n1454) );
  NANDN U2175 ( .A(n29120), .B(n1454), .Z(n1455) );
  AND U2176 ( .A(n29121), .B(n1455), .Z(n1456) );
  OR U2177 ( .A(n1456), .B(n29122), .Z(n1457) );
  NAND U2178 ( .A(n29123), .B(n1457), .Z(n1458) );
  NAND U2179 ( .A(n23943), .B(n1458), .Z(n1459) );
  AND U2180 ( .A(n29124), .B(n29125), .Z(n1460) );
  NAND U2181 ( .A(n1459), .B(n1460), .Z(n1461) );
  NAND U2182 ( .A(n29126), .B(n1461), .Z(n1462) );
  NAND U2183 ( .A(n29127), .B(n1462), .Z(n1463) );
  NANDN U2184 ( .A(n29128), .B(n1463), .Z(n1464) );
  AND U2185 ( .A(n29129), .B(n1464), .Z(n1465) );
  OR U2186 ( .A(n1465), .B(n29130), .Z(n1466) );
  NAND U2187 ( .A(n29131), .B(n1466), .Z(n1467) );
  NANDN U2188 ( .A(n29132), .B(n1467), .Z(n1468) );
  NAND U2189 ( .A(n23942), .B(n1468), .Z(n29135) );
  NAND U2190 ( .A(n23938), .B(n29166), .Z(n1469) );
  NAND U2191 ( .A(n29167), .B(n1469), .Z(n1470) );
  ANDN U2192 ( .B(n1470), .A(n29168), .Z(n1471) );
  NAND U2193 ( .A(n1471), .B(n29169), .Z(n1472) );
  NANDN U2194 ( .A(n29170), .B(n1472), .Z(n1473) );
  AND U2195 ( .A(n29171), .B(n1473), .Z(n1474) );
  AND U2196 ( .A(n23936), .B(n23937), .Z(n1475) );
  NANDN U2197 ( .A(n1474), .B(n29172), .Z(n1476) );
  AND U2198 ( .A(n1475), .B(n1476), .Z(n1477) );
  NANDN U2199 ( .A(n1477), .B(n29173), .Z(n1478) );
  NANDN U2200 ( .A(n23935), .B(n1478), .Z(n1479) );
  NAND U2201 ( .A(n23934), .B(n1479), .Z(n1480) );
  ANDN U2202 ( .B(n1480), .A(n29174), .Z(n29177) );
  NANDN U2203 ( .A(n23926), .B(n29196), .Z(n1481) );
  NAND U2204 ( .A(n23925), .B(n1481), .Z(n1482) );
  AND U2205 ( .A(n29197), .B(n1482), .Z(n1483) );
  ANDN U2206 ( .B(n29198), .A(n1483), .Z(n1484) );
  NAND U2207 ( .A(n29199), .B(n1484), .Z(n1485) );
  ANDN U2208 ( .B(n1485), .A(n29200), .Z(n1486) );
  NANDN U2209 ( .A(n1486), .B(n29201), .Z(n1487) );
  NANDN U2210 ( .A(n29202), .B(n1487), .Z(n1488) );
  NAND U2211 ( .A(n29203), .B(n1488), .Z(n1489) );
  NANDN U2212 ( .A(n29204), .B(n1489), .Z(n1490) );
  NAND U2213 ( .A(n29205), .B(n1490), .Z(n1491) );
  ANDN U2214 ( .B(n1491), .A(n29206), .Z(n1492) );
  ANDN U2215 ( .B(n29208), .A(n1492), .Z(n1493) );
  NAND U2216 ( .A(n29207), .B(n1493), .Z(n1494) );
  ANDN U2217 ( .B(n1494), .A(n29209), .Z(n1495) );
  NANDN U2218 ( .A(n1495), .B(n29210), .Z(n1496) );
  ANDN U2219 ( .B(n1496), .A(n29211), .Z(n29215) );
  NAND U2220 ( .A(n29264), .B(n29265), .Z(n1497) );
  NAND U2221 ( .A(n29268), .B(n1497), .Z(n1498) );
  NANDN U2222 ( .A(n29269), .B(n1498), .Z(n1499) );
  NAND U2223 ( .A(n29270), .B(n1499), .Z(n1500) );
  NANDN U2224 ( .A(n23915), .B(n1500), .Z(n1501) );
  AND U2225 ( .A(n23914), .B(n1501), .Z(n1502) );
  OR U2226 ( .A(n23913), .B(n1502), .Z(n1503) );
  NAND U2227 ( .A(n29271), .B(n1503), .Z(n1504) );
  NANDN U2228 ( .A(n29272), .B(n1504), .Z(n1505) );
  AND U2229 ( .A(n29274), .B(n29273), .Z(n1506) );
  NAND U2230 ( .A(n1505), .B(n1506), .Z(n1507) );
  NANDN U2231 ( .A(n29275), .B(n1507), .Z(n1508) );
  AND U2232 ( .A(n23912), .B(n23911), .Z(n1509) );
  NAND U2233 ( .A(n1508), .B(n1509), .Z(n1510) );
  NANDN U2234 ( .A(n29276), .B(n1510), .Z(n29277) );
  NAND U2235 ( .A(n29307), .B(n29308), .Z(n1511) );
  NANDN U2236 ( .A(n29309), .B(n1511), .Z(n1512) );
  NAND U2237 ( .A(n29310), .B(n1512), .Z(n1513) );
  NAND U2238 ( .A(n29311), .B(n1513), .Z(n1514) );
  AND U2239 ( .A(n23904), .B(n1514), .Z(n1515) );
  NAND U2240 ( .A(n1515), .B(n23903), .Z(n1516) );
  NAND U2241 ( .A(n29312), .B(n1516), .Z(n1517) );
  NANDN U2242 ( .A(n23902), .B(n1517), .Z(n1518) );
  AND U2243 ( .A(n23901), .B(n1518), .Z(n1519) );
  OR U2244 ( .A(n29313), .B(n1519), .Z(n1520) );
  NAND U2245 ( .A(n29314), .B(n1520), .Z(n1521) );
  NAND U2246 ( .A(n29315), .B(n1521), .Z(n1522) );
  ANDN U2247 ( .B(n1522), .A(n29316), .Z(n29320) );
  NAND U2248 ( .A(n29353), .B(n29352), .Z(n1523) );
  NANDN U2249 ( .A(n29354), .B(n1523), .Z(n1524) );
  NAND U2250 ( .A(n29355), .B(n1524), .Z(n1525) );
  NANDN U2251 ( .A(n1525), .B(n29356), .Z(n1526) );
  NANDN U2252 ( .A(n29357), .B(n1526), .Z(n1527) );
  NAND U2253 ( .A(n29358), .B(n1527), .Z(n1528) );
  NANDN U2254 ( .A(n29359), .B(n1528), .Z(n1529) );
  NAND U2255 ( .A(n29360), .B(n1529), .Z(n1530) );
  ANDN U2256 ( .B(n1530), .A(n29361), .Z(n1531) );
  NANDN U2257 ( .A(n1531), .B(n29362), .Z(n1532) );
  ANDN U2258 ( .B(n1532), .A(n23896), .Z(n1533) );
  NANDN U2259 ( .A(n1533), .B(n23895), .Z(n1534) );
  NANDN U2260 ( .A(n29363), .B(n1534), .Z(n1535) );
  NAND U2261 ( .A(n29364), .B(n1535), .Z(n29365) );
  NAND U2262 ( .A(n29392), .B(n23888), .Z(n1536) );
  NAND U2263 ( .A(n29393), .B(n1536), .Z(n1537) );
  NANDN U2264 ( .A(n29394), .B(n1537), .Z(n1538) );
  NAND U2265 ( .A(n29395), .B(n1538), .Z(n1539) );
  NANDN U2266 ( .A(n29396), .B(n1539), .Z(n1540) );
  AND U2267 ( .A(n29397), .B(n1540), .Z(n1541) );
  OR U2268 ( .A(n1541), .B(n29398), .Z(n1542) );
  NAND U2269 ( .A(n29399), .B(n1542), .Z(n1543) );
  NAND U2270 ( .A(n29400), .B(n1543), .Z(n1544) );
  NANDN U2271 ( .A(n1544), .B(n29401), .Z(n1545) );
  AND U2272 ( .A(n29402), .B(n1545), .Z(n1546) );
  OR U2273 ( .A(n29403), .B(n1546), .Z(n1547) );
  NAND U2274 ( .A(n29404), .B(n1547), .Z(n1548) );
  NANDN U2275 ( .A(n23887), .B(n1548), .Z(n29405) );
  NAND U2276 ( .A(n29432), .B(n29433), .Z(n1549) );
  NAND U2277 ( .A(n29434), .B(n1549), .Z(n1550) );
  NANDN U2278 ( .A(n29435), .B(n1550), .Z(n1551) );
  NAND U2279 ( .A(n29436), .B(n1551), .Z(n1552) );
  NAND U2280 ( .A(n29437), .B(n1552), .Z(n1553) );
  ANDN U2281 ( .B(n1553), .A(n29438), .Z(n1554) );
  NANDN U2282 ( .A(n1554), .B(n29439), .Z(n1555) );
  NANDN U2283 ( .A(n29440), .B(n1555), .Z(n1556) );
  NAND U2284 ( .A(n29441), .B(n1556), .Z(n1557) );
  NANDN U2285 ( .A(n23878), .B(n1557), .Z(n1558) );
  NAND U2286 ( .A(n23877), .B(n1558), .Z(n1559) );
  AND U2287 ( .A(n29442), .B(n1559), .Z(n1560) );
  NAND U2288 ( .A(n23876), .B(n1560), .Z(n29443) );
  NAND U2289 ( .A(n29467), .B(n29468), .Z(n1561) );
  NAND U2290 ( .A(n29469), .B(n1561), .Z(n1562) );
  NANDN U2291 ( .A(n23871), .B(n1562), .Z(n1563) );
  NAND U2292 ( .A(n23870), .B(n1563), .Z(n1564) );
  NAND U2293 ( .A(n29470), .B(n1564), .Z(n1565) );
  ANDN U2294 ( .B(n1565), .A(n29471), .Z(n1566) );
  NANDN U2295 ( .A(n1566), .B(n23869), .Z(n1567) );
  ANDN U2296 ( .B(n1567), .A(n29472), .Z(n1568) );
  NANDN U2297 ( .A(n1568), .B(n29473), .Z(n1569) );
  NANDN U2298 ( .A(n23868), .B(n1569), .Z(n1570) );
  NAND U2299 ( .A(n23867), .B(n1570), .Z(n29476) );
  OR U2300 ( .A(n29498), .B(n29499), .Z(n1571) );
  ANDN U2301 ( .B(n1571), .A(n29500), .Z(n1572) );
  NANDN U2302 ( .A(n1572), .B(n29501), .Z(n1573) );
  NANDN U2303 ( .A(n23860), .B(n1573), .Z(n1574) );
  NAND U2304 ( .A(n23859), .B(n1574), .Z(n1575) );
  AND U2305 ( .A(n29503), .B(n29502), .Z(n1576) );
  NAND U2306 ( .A(n1575), .B(n1576), .Z(n1577) );
  NAND U2307 ( .A(n29504), .B(n1577), .Z(n1578) );
  ANDN U2308 ( .B(n23858), .A(n23857), .Z(n1579) );
  NAND U2309 ( .A(n1578), .B(n1579), .Z(n1580) );
  NANDN U2310 ( .A(n29505), .B(n1580), .Z(n1581) );
  NOR U2311 ( .A(n29507), .B(n29506), .Z(n1582) );
  NAND U2312 ( .A(n1581), .B(n1582), .Z(n1583) );
  NANDN U2313 ( .A(n29508), .B(n1583), .Z(n29509) );
  NANDN U2314 ( .A(n15489), .B(n15490), .Z(n24541) );
  NANDN U2315 ( .A(n15449), .B(n15450), .Z(n24581) );
  NANDN U2316 ( .A(n15405), .B(n15406), .Z(n24625) );
  NANDN U2317 ( .A(n15373), .B(n15374), .Z(n24665) );
  NANDN U2318 ( .A(n15342), .B(n15343), .Z(n24705) );
  ANDN U2319 ( .B(n15313), .A(n15312), .Z(n24739) );
  ANDN U2320 ( .B(n15267), .A(n15266), .Z(n24783) );
  XNOR U2321 ( .A(y[146]), .B(x[146]), .Z(n1584) );
  NAND U2322 ( .A(n15230), .B(n1584), .Z(n24825) );
  XNOR U2323 ( .A(y[150]), .B(x[150]), .Z(n1585) );
  NAND U2324 ( .A(n15223), .B(n1585), .Z(n24833) );
  NANDN U2325 ( .A(n15182), .B(n15183), .Z(n24873) );
  ANDN U2326 ( .B(n15112), .A(n15111), .Z(n24943) );
  XNOR U2327 ( .A(x[210]), .B(y[210]), .Z(n1586) );
  NAND U2328 ( .A(n15101), .B(n1586), .Z(n24953) );
  XNOR U2329 ( .A(x[230]), .B(y[230]), .Z(n1587) );
  NAND U2330 ( .A(n15061), .B(n1587), .Z(n24993) );
  NANDN U2331 ( .A(x[262]), .B(y[262]), .Z(n1588) );
  ANDN U2332 ( .B(n1588), .A(n14999), .Z(n25059) );
  ANDN U2333 ( .B(n14972), .A(n14971), .Z(n25099) );
  XNOR U2334 ( .A(y[306]), .B(x[306]), .Z(n1589) );
  NAND U2335 ( .A(n14926), .B(n1589), .Z(n25145) );
  NANDN U2336 ( .A(x[324]), .B(y[324]), .Z(n1590) );
  ANDN U2337 ( .B(n1590), .A(n14888), .Z(n25183) );
  ANDN U2338 ( .B(n14877), .A(n14876), .Z(n25195) );
  NANDN U2339 ( .A(n14846), .B(n14847), .Z(n25233) );
  NANDN U2340 ( .A(n14782), .B(n14783), .Z(n25285) );
  NANDN U2341 ( .A(n14762), .B(n14763), .Z(n25325) );
  NANDN U2342 ( .A(n14726), .B(n14727), .Z(n25365) );
  NANDN U2343 ( .A(n14696), .B(n14697), .Z(n25401) );
  NANDN U2344 ( .A(n14656), .B(n14657), .Z(n25441) );
  NANDN U2345 ( .A(n14612), .B(n14613), .Z(n25485) );
  NANDN U2346 ( .A(n14604), .B(n14605), .Z(n25493) );
  NANDN U2347 ( .A(n14533), .B(n14534), .Z(n25549) );
  NANDN U2348 ( .A(n14529), .B(n14530), .Z(n25552) );
  NANDN U2349 ( .A(n14489), .B(n14490), .Z(n25592) );
  NANDN U2350 ( .A(n14439), .B(n14440), .Z(n25638) );
  NANDN U2351 ( .A(n14395), .B(n14396), .Z(n25686) );
  NANDN U2352 ( .A(n14355), .B(n14356), .Z(n25726) );
  NANDN U2353 ( .A(n14315), .B(n14316), .Z(n25766) );
  NANDN U2354 ( .A(n14271), .B(n14272), .Z(n25810) );
  NAND U2355 ( .A(n25863), .B(n24534), .Z(n1591) );
  NAND U2356 ( .A(n25864), .B(n1591), .Z(n1592) );
  AND U2357 ( .A(n24533), .B(n1592), .Z(n1593) );
  NANDN U2358 ( .A(n1593), .B(n25865), .Z(n1594) );
  NAND U2359 ( .A(n25866), .B(n1594), .Z(n1595) );
  NAND U2360 ( .A(n25867), .B(n1595), .Z(n1596) );
  NAND U2361 ( .A(n24532), .B(n1596), .Z(n1597) );
  NAND U2362 ( .A(n25868), .B(n1597), .Z(n1598) );
  AND U2363 ( .A(n24531), .B(n1598), .Z(n1599) );
  NANDN U2364 ( .A(n1599), .B(n25869), .Z(n1600) );
  AND U2365 ( .A(n25870), .B(n1600), .Z(n1601) );
  OR U2366 ( .A(n24530), .B(n1601), .Z(n1602) );
  NAND U2367 ( .A(n25871), .B(n1602), .Z(n1603) );
  NAND U2368 ( .A(n25872), .B(n1603), .Z(n25873) );
  ANDN U2369 ( .B(n14175), .A(n14174), .Z(n25887) );
  NOR U2370 ( .A(n14128), .B(n14129), .Z(n25908) );
  NANDN U2371 ( .A(n25925), .B(n25924), .Z(n1604) );
  NAND U2372 ( .A(n25926), .B(n1604), .Z(n1605) );
  AND U2373 ( .A(n25927), .B(n1605), .Z(n1606) );
  NANDN U2374 ( .A(n1606), .B(n25928), .Z(n1607) );
  NAND U2375 ( .A(n25929), .B(n1607), .Z(n1608) );
  NANDN U2376 ( .A(n24514), .B(n1608), .Z(n1609) );
  NAND U2377 ( .A(n24513), .B(n1609), .Z(n1610) );
  NANDN U2378 ( .A(n25930), .B(n1610), .Z(n1611) );
  AND U2379 ( .A(n25931), .B(n1611), .Z(n1612) );
  OR U2380 ( .A(n24512), .B(n1612), .Z(n1613) );
  NAND U2381 ( .A(n24511), .B(n1613), .Z(n1614) );
  NANDN U2382 ( .A(n24510), .B(n1614), .Z(n25932) );
  ANDN U2383 ( .B(n14069), .A(n14068), .Z(n25953) );
  NANDN U2384 ( .A(n14022), .B(n14023), .Z(n25995) );
  NANDN U2385 ( .A(n14008), .B(n14007), .Z(n1615) );
  ANDN U2386 ( .B(n1615), .A(n14009), .Z(n26045) );
  NANDN U2387 ( .A(n26066), .B(n26065), .Z(n1616) );
  NAND U2388 ( .A(n26067), .B(n1616), .Z(n1617) );
  NANDN U2389 ( .A(n26068), .B(n1617), .Z(n1618) );
  NAND U2390 ( .A(n26069), .B(n1618), .Z(n1619) );
  NANDN U2391 ( .A(n26070), .B(n1619), .Z(n1620) );
  AND U2392 ( .A(n26071), .B(n1620), .Z(n1621) );
  OR U2393 ( .A(n1621), .B(n26072), .Z(n1622) );
  NAND U2394 ( .A(n26073), .B(n1622), .Z(n1623) );
  NAND U2395 ( .A(n26074), .B(n1623), .Z(n1624) );
  NAND U2396 ( .A(n24505), .B(n1624), .Z(n1625) );
  NAND U2397 ( .A(n26075), .B(n1625), .Z(n1626) );
  AND U2398 ( .A(n26076), .B(n1626), .Z(n1627) );
  NANDN U2399 ( .A(n1627), .B(n26077), .Z(n1628) );
  NAND U2400 ( .A(n24504), .B(n1628), .Z(n1629) );
  NAND U2401 ( .A(n26078), .B(n1629), .Z(n1630) );
  NAND U2402 ( .A(n24503), .B(n1630), .Z(n26081) );
  NOR U2403 ( .A(n13957), .B(n13958), .Z(n26107) );
  OR U2404 ( .A(n26120), .B(n26121), .Z(n1631) );
  NAND U2405 ( .A(n26122), .B(n1631), .Z(n1632) );
  ANDN U2406 ( .B(n1632), .A(n26123), .Z(n1633) );
  NANDN U2407 ( .A(n1633), .B(n26124), .Z(n1634) );
  NANDN U2408 ( .A(n26125), .B(n1634), .Z(n1635) );
  NAND U2409 ( .A(n26126), .B(n1635), .Z(n1636) );
  NANDN U2410 ( .A(n1636), .B(n26127), .Z(n1637) );
  NAND U2411 ( .A(n24491), .B(n1637), .Z(n1638) );
  NAND U2412 ( .A(n26128), .B(n1638), .Z(n1639) );
  NAND U2413 ( .A(n26129), .B(n1639), .Z(n1640) );
  NANDN U2414 ( .A(n26130), .B(n1640), .Z(n1641) );
  AND U2415 ( .A(n26131), .B(n1641), .Z(n1642) );
  NANDN U2416 ( .A(n1642), .B(n26132), .Z(n1643) );
  NAND U2417 ( .A(n26133), .B(n1643), .Z(n1644) );
  NAND U2418 ( .A(n24490), .B(n1644), .Z(n1645) );
  NANDN U2419 ( .A(n24489), .B(n1645), .Z(n26134) );
  ANDN U2420 ( .B(n13895), .A(n13894), .Z(n26165) );
  NAND U2421 ( .A(n26203), .B(n26204), .Z(n1646) );
  NANDN U2422 ( .A(n26205), .B(n1646), .Z(n1647) );
  NAND U2423 ( .A(n24481), .B(n1647), .Z(n1648) );
  NANDN U2424 ( .A(n26206), .B(n1648), .Z(n1649) );
  NAND U2425 ( .A(n26207), .B(n1649), .Z(n1650) );
  ANDN U2426 ( .B(n1650), .A(n24480), .Z(n1651) );
  NANDN U2427 ( .A(n1651), .B(n24479), .Z(n1652) );
  NAND U2428 ( .A(n26208), .B(n1652), .Z(n1653) );
  NANDN U2429 ( .A(n26209), .B(n1653), .Z(n1654) );
  NAND U2430 ( .A(n26210), .B(n1654), .Z(n1655) );
  NANDN U2431 ( .A(n26211), .B(n1655), .Z(n1656) );
  AND U2432 ( .A(n26212), .B(n1656), .Z(n1657) );
  OR U2433 ( .A(n26213), .B(n1657), .Z(n1658) );
  NAND U2434 ( .A(n26214), .B(n1658), .Z(n1659) );
  NANDN U2435 ( .A(n26215), .B(n1659), .Z(n26216) );
  NOR U2436 ( .A(n13830), .B(n13831), .Z(n26248) );
  NAND U2437 ( .A(n13814), .B(n13813), .Z(n1660) );
  ANDN U2438 ( .B(n1660), .A(n13815), .Z(n26273) );
  NANDN U2439 ( .A(n13798), .B(n13799), .Z(n24464) );
  ANDN U2440 ( .B(n13765), .A(n13768), .Z(n1661) );
  NANDN U2441 ( .A(n13766), .B(n13767), .Z(n1662) );
  NAND U2442 ( .A(n1661), .B(n1662), .Z(n26319) );
  NAND U2443 ( .A(n26332), .B(n26331), .Z(n1663) );
  NAND U2444 ( .A(n24454), .B(n1663), .Z(n1664) );
  ANDN U2445 ( .B(n1664), .A(n26333), .Z(n1665) );
  NANDN U2446 ( .A(n1665), .B(n26334), .Z(n1666) );
  NAND U2447 ( .A(n26335), .B(n1666), .Z(n1667) );
  NAND U2448 ( .A(n24453), .B(n1667), .Z(n1668) );
  NAND U2449 ( .A(n26336), .B(n1668), .Z(n1669) );
  AND U2450 ( .A(n24452), .B(n1669), .Z(n1670) );
  NANDN U2451 ( .A(n24451), .B(n1670), .Z(n1671) );
  NANDN U2452 ( .A(n26337), .B(n1671), .Z(n1672) );
  NAND U2453 ( .A(n26338), .B(n1672), .Z(n1673) );
  ANDN U2454 ( .B(n1673), .A(n26339), .Z(n1674) );
  NANDN U2455 ( .A(n1674), .B(n24450), .Z(n1675) );
  NAND U2456 ( .A(n26340), .B(n1675), .Z(n1676) );
  NAND U2457 ( .A(n26341), .B(n1676), .Z(n26342) );
  NOR U2458 ( .A(n13734), .B(n13735), .Z(n26358) );
  NANDN U2459 ( .A(n13881), .B(n4669), .Z(n1677) );
  AND U2460 ( .A(n16703), .B(n1677), .Z(n26185) );
  NANDN U2461 ( .A(n26393), .B(n26392), .Z(n1678) );
  NAND U2462 ( .A(n26395), .B(n1678), .Z(n1679) );
  NANDN U2463 ( .A(n26396), .B(n1679), .Z(n1680) );
  NANDN U2464 ( .A(n24443), .B(n1680), .Z(n1681) );
  NAND U2465 ( .A(n24442), .B(n1681), .Z(n1682) );
  AND U2466 ( .A(n26397), .B(n1682), .Z(n1683) );
  NANDN U2467 ( .A(n24440), .B(n24439), .Z(n1684) );
  AND U2468 ( .A(n24441), .B(n1684), .Z(n1685) );
  NANDN U2469 ( .A(n1683), .B(n26398), .Z(n1686) );
  NAND U2470 ( .A(n1685), .B(n1686), .Z(n1687) );
  NAND U2471 ( .A(n26399), .B(n1687), .Z(n1688) );
  NANDN U2472 ( .A(n24438), .B(n1688), .Z(n1689) );
  NANDN U2473 ( .A(n26400), .B(n1689), .Z(n1690) );
  AND U2474 ( .A(n26401), .B(n1690), .Z(n1691) );
  OR U2475 ( .A(n1691), .B(n26402), .Z(n1692) );
  NAND U2476 ( .A(n26403), .B(n1692), .Z(n1693) );
  NAND U2477 ( .A(n26404), .B(n1693), .Z(n26405) );
  NANDN U2478 ( .A(n13685), .B(n13686), .Z(n26446) );
  NANDN U2479 ( .A(n16817), .B(n4638), .Z(n1694) );
  AND U2480 ( .A(n16822), .B(n1694), .Z(n26234) );
  NAND U2481 ( .A(n26478), .B(n26479), .Z(n1695) );
  NAND U2482 ( .A(n24434), .B(n1695), .Z(n1696) );
  NANDN U2483 ( .A(n24433), .B(n1696), .Z(n1697) );
  NAND U2484 ( .A(n24432), .B(n1697), .Z(n1698) );
  NAND U2485 ( .A(n26480), .B(n1698), .Z(n1699) );
  ANDN U2486 ( .B(n1699), .A(n26481), .Z(n1700) );
  OR U2487 ( .A(n1700), .B(n26482), .Z(n1701) );
  NANDN U2488 ( .A(n26483), .B(n1701), .Z(n1702) );
  AND U2489 ( .A(n26484), .B(n1702), .Z(n1703) );
  NAND U2490 ( .A(n24429), .B(n24430), .Z(n1704) );
  ANDN U2491 ( .B(n1704), .A(n24431), .Z(n1705) );
  NANDN U2492 ( .A(n1703), .B(n26485), .Z(n1706) );
  NAND U2493 ( .A(n1705), .B(n1706), .Z(n1707) );
  NAND U2494 ( .A(n26486), .B(n1707), .Z(n1708) );
  NANDN U2495 ( .A(n24428), .B(n1708), .Z(n26487) );
  NANDN U2496 ( .A(x[1100]), .B(y[1100]), .Z(n1709) );
  ANDN U2497 ( .B(n1709), .A(n4598), .Z(n26299) );
  AND U2498 ( .A(n26519), .B(n26518), .Z(n1710) );
  NAND U2499 ( .A(n26520), .B(n1710), .Z(n1711) );
  AND U2500 ( .A(n24422), .B(n1711), .Z(n1712) );
  NANDN U2501 ( .A(n1712), .B(n26521), .Z(n1713) );
  NAND U2502 ( .A(n26522), .B(n1713), .Z(n1714) );
  NANDN U2503 ( .A(n26523), .B(n1714), .Z(n1715) );
  NAND U2504 ( .A(n26524), .B(n1715), .Z(n1716) );
  NANDN U2505 ( .A(n26525), .B(n1716), .Z(n1717) );
  AND U2506 ( .A(n26526), .B(n1717), .Z(n1718) );
  NANDN U2507 ( .A(n1718), .B(n26527), .Z(n1719) );
  NANDN U2508 ( .A(n24421), .B(n1719), .Z(n1720) );
  NAND U2509 ( .A(n24420), .B(n1720), .Z(n1721) );
  NAND U2510 ( .A(n26528), .B(n1721), .Z(n1722) );
  NANDN U2511 ( .A(n26529), .B(n1722), .Z(n1723) );
  ANDN U2512 ( .B(n1723), .A(n26530), .Z(n26532) );
  NANDN U2513 ( .A(n26557), .B(n26556), .Z(n1724) );
  NAND U2514 ( .A(n26558), .B(n1724), .Z(n1725) );
  NAND U2515 ( .A(n26559), .B(n1725), .Z(n1726) );
  NAND U2516 ( .A(n26560), .B(n1726), .Z(n1727) );
  NANDN U2517 ( .A(n26561), .B(n1727), .Z(n1728) );
  AND U2518 ( .A(n26562), .B(n1728), .Z(n1729) );
  OR U2519 ( .A(n1729), .B(n26563), .Z(n1730) );
  NAND U2520 ( .A(n26564), .B(n1730), .Z(n1731) );
  NANDN U2521 ( .A(n24413), .B(n1731), .Z(n1732) );
  NAND U2522 ( .A(n26565), .B(n1732), .Z(n1733) );
  NANDN U2523 ( .A(n26566), .B(n1733), .Z(n1734) );
  AND U2524 ( .A(n26567), .B(n1734), .Z(n1735) );
  OR U2525 ( .A(n1735), .B(n26568), .Z(n1736) );
  NAND U2526 ( .A(n26569), .B(n1736), .Z(n1737) );
  ANDN U2527 ( .B(n1737), .A(n24412), .Z(n1738) );
  NANDN U2528 ( .A(n1738), .B(n26570), .Z(n1739) );
  NAND U2529 ( .A(n26571), .B(n1739), .Z(n1740) );
  NANDN U2530 ( .A(n26572), .B(n1740), .Z(n26575) );
  ANDN U2531 ( .B(n13587), .A(n13586), .Z(n26589) );
  NANDN U2532 ( .A(n26645), .B(n26644), .Z(n1741) );
  NAND U2533 ( .A(n26646), .B(n1741), .Z(n1742) );
  NANDN U2534 ( .A(n26647), .B(n1742), .Z(n1743) );
  NAND U2535 ( .A(n26648), .B(n1743), .Z(n1744) );
  NANDN U2536 ( .A(n26649), .B(n1744), .Z(n1745) );
  AND U2537 ( .A(n26650), .B(n1745), .Z(n1746) );
  OR U2538 ( .A(n26651), .B(n1746), .Z(n1747) );
  NAND U2539 ( .A(n26652), .B(n1747), .Z(n1748) );
  NANDN U2540 ( .A(n26653), .B(n1748), .Z(n1749) );
  NAND U2541 ( .A(n26654), .B(n1749), .Z(n1750) );
  NAND U2542 ( .A(n26655), .B(n1750), .Z(n1751) );
  AND U2543 ( .A(n26656), .B(n1751), .Z(n1752) );
  OR U2544 ( .A(n1752), .B(n26657), .Z(n1753) );
  NANDN U2545 ( .A(n26658), .B(n1753), .Z(n1754) );
  AND U2546 ( .A(n26659), .B(n1754), .Z(n1755) );
  OR U2547 ( .A(n1755), .B(n26660), .Z(n1756) );
  NAND U2548 ( .A(n26661), .B(n1756), .Z(n1757) );
  NANDN U2549 ( .A(n26662), .B(n1757), .Z(n1758) );
  NANDN U2550 ( .A(n24407), .B(n1758), .Z(n26663) );
  ANDN U2551 ( .B(n13543), .A(n13542), .Z(n26697) );
  NANDN U2552 ( .A(n13533), .B(n13534), .Z(n26717) );
  NANDN U2553 ( .A(n26749), .B(n26748), .Z(n1759) );
  NAND U2554 ( .A(n26750), .B(n1759), .Z(n1760) );
  ANDN U2555 ( .B(n1760), .A(n26751), .Z(n1761) );
  NANDN U2556 ( .A(n1761), .B(n26752), .Z(n1762) );
  NANDN U2557 ( .A(n26753), .B(n1762), .Z(n1763) );
  NAND U2558 ( .A(n26754), .B(n1763), .Z(n1764) );
  NANDN U2559 ( .A(n26755), .B(n1764), .Z(n1765) );
  NAND U2560 ( .A(n26756), .B(n1765), .Z(n1766) );
  ANDN U2561 ( .B(n1766), .A(n26757), .Z(n1767) );
  NANDN U2562 ( .A(n1767), .B(n26758), .Z(n1768) );
  NANDN U2563 ( .A(n26759), .B(n1768), .Z(n1769) );
  NAND U2564 ( .A(n24399), .B(n1769), .Z(n1770) );
  NANDN U2565 ( .A(n26760), .B(n1770), .Z(n1771) );
  NAND U2566 ( .A(n26761), .B(n1771), .Z(n1772) );
  ANDN U2567 ( .B(n1772), .A(n24398), .Z(n1773) );
  NANDN U2568 ( .A(n1773), .B(n26762), .Z(n1774) );
  NAND U2569 ( .A(n26763), .B(n1774), .Z(n1775) );
  NANDN U2570 ( .A(n26764), .B(n1775), .Z(n26765) );
  OR U2571 ( .A(n26797), .B(n26796), .Z(n1776) );
  NAND U2572 ( .A(n26798), .B(n1776), .Z(n1777) );
  NANDN U2573 ( .A(n26799), .B(n1777), .Z(n1778) );
  NAND U2574 ( .A(n26800), .B(n1778), .Z(n1779) );
  NAND U2575 ( .A(n26801), .B(n1779), .Z(n1780) );
  ANDN U2576 ( .B(n1780), .A(n26802), .Z(n1781) );
  NOR U2577 ( .A(n26804), .B(n26803), .Z(n1782) );
  NANDN U2578 ( .A(n1781), .B(n1782), .Z(n1783) );
  AND U2579 ( .A(n24392), .B(n1783), .Z(n1784) );
  NANDN U2580 ( .A(n1784), .B(n26805), .Z(n1785) );
  AND U2581 ( .A(n26806), .B(n1785), .Z(n1786) );
  OR U2582 ( .A(n26807), .B(n1786), .Z(n1787) );
  NAND U2583 ( .A(n26808), .B(n1787), .Z(n1788) );
  NANDN U2584 ( .A(n24391), .B(n1788), .Z(n26809) );
  NAND U2585 ( .A(n26836), .B(n26837), .Z(n1789) );
  NANDN U2586 ( .A(n26838), .B(n1789), .Z(n1790) );
  NAND U2587 ( .A(n26839), .B(n1790), .Z(n1791) );
  NANDN U2588 ( .A(n26840), .B(n1791), .Z(n1792) );
  NAND U2589 ( .A(n26841), .B(n1792), .Z(n1793) );
  AND U2590 ( .A(n26842), .B(n1793), .Z(n1794) );
  OR U2591 ( .A(n24383), .B(n1794), .Z(n1795) );
  NAND U2592 ( .A(n26843), .B(n1795), .Z(n1796) );
  NAND U2593 ( .A(n26844), .B(n1796), .Z(n1797) );
  OR U2594 ( .A(n1797), .B(n26845), .Z(n1798) );
  NAND U2595 ( .A(n26846), .B(n1798), .Z(n1799) );
  NAND U2596 ( .A(n24382), .B(n1799), .Z(n1800) );
  NAND U2597 ( .A(n26847), .B(n1800), .Z(n1801) );
  NANDN U2598 ( .A(n26848), .B(n1801), .Z(n1802) );
  AND U2599 ( .A(n26849), .B(n1802), .Z(n1803) );
  OR U2600 ( .A(n26850), .B(n1803), .Z(n1804) );
  NAND U2601 ( .A(n26851), .B(n1804), .Z(n1805) );
  NANDN U2602 ( .A(n26852), .B(n1805), .Z(n26853) );
  NAND U2603 ( .A(n26883), .B(n26882), .Z(n1806) );
  NANDN U2604 ( .A(n26885), .B(n1806), .Z(n1807) );
  NANDN U2605 ( .A(n24375), .B(n1807), .Z(n1808) );
  NAND U2606 ( .A(n24374), .B(n1808), .Z(n1809) );
  NAND U2607 ( .A(n26886), .B(n1809), .Z(n1810) );
  AND U2608 ( .A(n26887), .B(n1810), .Z(n1811) );
  NOR U2609 ( .A(n26889), .B(n1811), .Z(n1812) );
  NAND U2610 ( .A(n26888), .B(n1812), .Z(n1813) );
  AND U2611 ( .A(n26890), .B(n1813), .Z(n1814) );
  OR U2612 ( .A(n26891), .B(n1814), .Z(n1815) );
  NAND U2613 ( .A(n26892), .B(n1815), .Z(n1816) );
  NANDN U2614 ( .A(n26893), .B(n1816), .Z(n1817) );
  NAND U2615 ( .A(n26894), .B(n1817), .Z(n1818) );
  NANDN U2616 ( .A(n26895), .B(n1818), .Z(n1819) );
  AND U2617 ( .A(n26896), .B(n1819), .Z(n1820) );
  OR U2618 ( .A(n26897), .B(n1820), .Z(n1821) );
  NAND U2619 ( .A(n26898), .B(n1821), .Z(n1822) );
  NANDN U2620 ( .A(n26899), .B(n1822), .Z(n26900) );
  OR U2621 ( .A(n26929), .B(n26928), .Z(n1823) );
  NANDN U2622 ( .A(n26930), .B(n1823), .Z(n1824) );
  NANDN U2623 ( .A(n26931), .B(n1824), .Z(n1825) );
  NAND U2624 ( .A(n26932), .B(n1825), .Z(n1826) );
  NANDN U2625 ( .A(n26933), .B(n1826), .Z(n1827) );
  AND U2626 ( .A(n26934), .B(n1827), .Z(n1828) );
  OR U2627 ( .A(n26935), .B(n1828), .Z(n1829) );
  NAND U2628 ( .A(n26936), .B(n1829), .Z(n1830) );
  NANDN U2629 ( .A(n26937), .B(n1830), .Z(n1831) );
  NAND U2630 ( .A(n26938), .B(n1831), .Z(n1832) );
  NAND U2631 ( .A(n24367), .B(n1832), .Z(n1833) );
  ANDN U2632 ( .B(n1833), .A(n26939), .Z(n1834) );
  NANDN U2633 ( .A(n1834), .B(n26940), .Z(n1835) );
  NANDN U2634 ( .A(n26941), .B(n1835), .Z(n1836) );
  NAND U2635 ( .A(n26942), .B(n1836), .Z(n1837) );
  NAND U2636 ( .A(n26943), .B(n1837), .Z(n26944) );
  NAND U2637 ( .A(n26976), .B(n26977), .Z(n1838) );
  NANDN U2638 ( .A(n24363), .B(n1838), .Z(n1839) );
  NAND U2639 ( .A(n24362), .B(n1839), .Z(n1840) );
  NANDN U2640 ( .A(n24361), .B(n1840), .Z(n1841) );
  NAND U2641 ( .A(n24360), .B(n1841), .Z(n1842) );
  AND U2642 ( .A(n26978), .B(n1842), .Z(n1843) );
  OR U2643 ( .A(n26979), .B(n1843), .Z(n1844) );
  NAND U2644 ( .A(n26980), .B(n1844), .Z(n1845) );
  NANDN U2645 ( .A(n26981), .B(n1845), .Z(n1846) );
  NAND U2646 ( .A(n26982), .B(n1846), .Z(n1847) );
  NANDN U2647 ( .A(n26983), .B(n1847), .Z(n1848) );
  AND U2648 ( .A(n26984), .B(n1848), .Z(n1849) );
  OR U2649 ( .A(n26985), .B(n1849), .Z(n1850) );
  NAND U2650 ( .A(n26986), .B(n1850), .Z(n1851) );
  NANDN U2651 ( .A(n26987), .B(n1851), .Z(n1852) );
  NAND U2652 ( .A(n26988), .B(n1852), .Z(n26989) );
  NANDN U2653 ( .A(n27021), .B(n27020), .Z(n1853) );
  NANDN U2654 ( .A(n27022), .B(n1853), .Z(n1854) );
  AND U2655 ( .A(n27023), .B(n1854), .Z(n1855) );
  OR U2656 ( .A(n27024), .B(n1855), .Z(n1856) );
  NAND U2657 ( .A(n27025), .B(n1856), .Z(n1857) );
  NAND U2658 ( .A(n27026), .B(n1857), .Z(n1858) );
  AND U2659 ( .A(n27028), .B(n27027), .Z(n1859) );
  NAND U2660 ( .A(n1858), .B(n1859), .Z(n1860) );
  NANDN U2661 ( .A(n27029), .B(n1860), .Z(n1861) );
  NAND U2662 ( .A(n27030), .B(n1861), .Z(n1862) );
  NANDN U2663 ( .A(n27031), .B(n1862), .Z(n1863) );
  ANDN U2664 ( .B(n1863), .A(n27032), .Z(n1864) );
  NANDN U2665 ( .A(n1864), .B(n27033), .Z(n1865) );
  NAND U2666 ( .A(n27034), .B(n1865), .Z(n1866) );
  NAND U2667 ( .A(n24354), .B(n1866), .Z(n27036) );
  NAND U2668 ( .A(n27065), .B(n27066), .Z(n1867) );
  NANDN U2669 ( .A(n27067), .B(n1867), .Z(n1868) );
  AND U2670 ( .A(n27068), .B(n1868), .Z(n1869) );
  NANDN U2671 ( .A(n1869), .B(n27069), .Z(n1870) );
  NAND U2672 ( .A(n27070), .B(n1870), .Z(n1871) );
  NANDN U2673 ( .A(n27071), .B(n1871), .Z(n1872) );
  NAND U2674 ( .A(n27072), .B(n1872), .Z(n1873) );
  NANDN U2675 ( .A(n27073), .B(n1873), .Z(n1874) );
  AND U2676 ( .A(n27074), .B(n1874), .Z(n1875) );
  OR U2677 ( .A(n27075), .B(n1875), .Z(n1876) );
  NAND U2678 ( .A(n24347), .B(n1876), .Z(n1877) );
  NAND U2679 ( .A(n27076), .B(n1877), .Z(n1878) );
  OR U2680 ( .A(n1878), .B(n27077), .Z(n1879) );
  NAND U2681 ( .A(n27078), .B(n1879), .Z(n1880) );
  NAND U2682 ( .A(n24346), .B(n1880), .Z(n1881) );
  NAND U2683 ( .A(n27079), .B(n1881), .Z(n1882) );
  NANDN U2684 ( .A(n27080), .B(n1882), .Z(n1883) );
  AND U2685 ( .A(n27081), .B(n1883), .Z(n27082) );
  NAND U2686 ( .A(n27112), .B(n27111), .Z(n1884) );
  NANDN U2687 ( .A(n27113), .B(n1884), .Z(n1885) );
  NAND U2688 ( .A(n27114), .B(n1885), .Z(n1886) );
  NAND U2689 ( .A(n27115), .B(n1886), .Z(n1887) );
  NANDN U2690 ( .A(n27116), .B(n1887), .Z(n1888) );
  AND U2691 ( .A(n27117), .B(n1888), .Z(n1889) );
  OR U2692 ( .A(n1889), .B(n27118), .Z(n1890) );
  NANDN U2693 ( .A(n27119), .B(n1890), .Z(n1891) );
  AND U2694 ( .A(n27120), .B(n1891), .Z(n1892) );
  OR U2695 ( .A(n1892), .B(n27121), .Z(n1893) );
  NAND U2696 ( .A(n27122), .B(n1893), .Z(n1894) );
  ANDN U2697 ( .B(n1894), .A(n27123), .Z(n1895) );
  NANDN U2698 ( .A(n1895), .B(n24340), .Z(n1896) );
  AND U2699 ( .A(n27124), .B(n1896), .Z(n1897) );
  NANDN U2700 ( .A(n1897), .B(n27125), .Z(n1898) );
  NAND U2701 ( .A(n27126), .B(n1898), .Z(n1899) );
  NANDN U2702 ( .A(n27127), .B(n1899), .Z(n27128) );
  NANDN U2703 ( .A(n13205), .B(n13206), .Z(n27169) );
  AND U2704 ( .A(n24333), .B(n24334), .Z(n1900) );
  NANDN U2705 ( .A(n27221), .B(n27220), .Z(n1901) );
  AND U2706 ( .A(n1900), .B(n1901), .Z(n1902) );
  OR U2707 ( .A(n1902), .B(n27222), .Z(n1903) );
  NAND U2708 ( .A(n27223), .B(n1903), .Z(n1904) );
  NANDN U2709 ( .A(n27224), .B(n1904), .Z(n1905) );
  NANDN U2710 ( .A(n24332), .B(n1905), .Z(n1906) );
  NAND U2711 ( .A(n27225), .B(n1906), .Z(n1907) );
  ANDN U2712 ( .B(n1907), .A(n27226), .Z(n1908) );
  OR U2713 ( .A(n1908), .B(n27227), .Z(n1909) );
  NANDN U2714 ( .A(n27228), .B(n1909), .Z(n1910) );
  ANDN U2715 ( .B(n1910), .A(n27229), .Z(n1911) );
  NANDN U2716 ( .A(n1911), .B(n27230), .Z(n1912) );
  NAND U2717 ( .A(n27231), .B(n1912), .Z(n1913) );
  NAND U2718 ( .A(n27232), .B(n1913), .Z(n27234) );
  NANDN U2719 ( .A(n27265), .B(n27264), .Z(n1914) );
  NAND U2720 ( .A(n27266), .B(n1914), .Z(n1915) );
  ANDN U2721 ( .B(n1915), .A(n27267), .Z(n1916) );
  NANDN U2722 ( .A(n1916), .B(n27268), .Z(n1917) );
  NANDN U2723 ( .A(n27269), .B(n1917), .Z(n1918) );
  NAND U2724 ( .A(n27270), .B(n1918), .Z(n1919) );
  NANDN U2725 ( .A(n27271), .B(n1919), .Z(n1920) );
  NAND U2726 ( .A(n27272), .B(n1920), .Z(n1921) );
  ANDN U2727 ( .B(n1921), .A(n27273), .Z(n1922) );
  NANDN U2728 ( .A(n1922), .B(n24327), .Z(n1923) );
  ANDN U2729 ( .B(n1923), .A(n27274), .Z(n1924) );
  NANDN U2730 ( .A(n1924), .B(n27275), .Z(n1925) );
  NANDN U2731 ( .A(n27276), .B(n1925), .Z(n1926) );
  NAND U2732 ( .A(n27277), .B(n1926), .Z(n27278) );
  NANDN U2733 ( .A(n27307), .B(n27308), .Z(n1927) );
  NANDN U2734 ( .A(n27309), .B(n1927), .Z(n1928) );
  AND U2735 ( .A(n27310), .B(n1928), .Z(n1929) );
  OR U2736 ( .A(n27311), .B(n1929), .Z(n1930) );
  NAND U2737 ( .A(n27312), .B(n1930), .Z(n1931) );
  NAND U2738 ( .A(n27313), .B(n1931), .Z(n1932) );
  NAND U2739 ( .A(n27314), .B(n1932), .Z(n1933) );
  NAND U2740 ( .A(n27315), .B(n1933), .Z(n1934) );
  ANDN U2741 ( .B(n1934), .A(n27316), .Z(n1935) );
  OR U2742 ( .A(n27317), .B(n1935), .Z(n1936) );
  NAND U2743 ( .A(n27318), .B(n1936), .Z(n1937) );
  NANDN U2744 ( .A(n27319), .B(n1937), .Z(n1938) );
  NAND U2745 ( .A(n27320), .B(n1938), .Z(n1939) );
  NANDN U2746 ( .A(n27321), .B(n1939), .Z(n1940) );
  AND U2747 ( .A(n27322), .B(n1940), .Z(n1941) );
  NAND U2748 ( .A(n24317), .B(n24318), .Z(n1942) );
  AND U2749 ( .A(n24319), .B(n1942), .Z(n1943) );
  OR U2750 ( .A(n27323), .B(n1941), .Z(n1944) );
  AND U2751 ( .A(n1943), .B(n1944), .Z(n27328) );
  NANDN U2752 ( .A(n27360), .B(n27359), .Z(n1945) );
  NAND U2753 ( .A(n27361), .B(n1945), .Z(n1946) );
  NANDN U2754 ( .A(n27362), .B(n1946), .Z(n1947) );
  NAND U2755 ( .A(n27363), .B(n1947), .Z(n1948) );
  NANDN U2756 ( .A(n27364), .B(n1948), .Z(n1949) );
  ANDN U2757 ( .B(n1949), .A(n27365), .Z(n1950) );
  NANDN U2758 ( .A(n1950), .B(n27366), .Z(n1951) );
  NANDN U2759 ( .A(n24313), .B(n1951), .Z(n1952) );
  NAND U2760 ( .A(n27367), .B(n1952), .Z(n1953) );
  NAND U2761 ( .A(n27368), .B(n1953), .Z(n1954) );
  NAND U2762 ( .A(n27369), .B(n1954), .Z(n1955) );
  AND U2763 ( .A(n27370), .B(n1955), .Z(n1956) );
  OR U2764 ( .A(n27371), .B(n1956), .Z(n1957) );
  NAND U2765 ( .A(n27372), .B(n1957), .Z(n1958) );
  NANDN U2766 ( .A(n24312), .B(n1958), .Z(n27373) );
  ANDN U2767 ( .B(n13013), .A(n13012), .Z(n27397) );
  ANDN U2768 ( .B(n27403), .A(n27402), .Z(n27404) );
  NAND U2769 ( .A(n27427), .B(n27428), .Z(n1959) );
  NAND U2770 ( .A(n27429), .B(n1959), .Z(n1960) );
  AND U2771 ( .A(n27430), .B(n1960), .Z(n1961) );
  NANDN U2772 ( .A(n1961), .B(n27431), .Z(n1962) );
  NAND U2773 ( .A(n27432), .B(n1962), .Z(n1963) );
  NAND U2774 ( .A(n27433), .B(n1963), .Z(n1964) );
  NANDN U2775 ( .A(n24299), .B(n1964), .Z(n1965) );
  NAND U2776 ( .A(n24298), .B(n1965), .Z(n1966) );
  ANDN U2777 ( .B(n1966), .A(n27434), .Z(n1967) );
  NANDN U2778 ( .A(n1967), .B(n27435), .Z(n1968) );
  NANDN U2779 ( .A(n24297), .B(n1968), .Z(n1969) );
  NAND U2780 ( .A(n24296), .B(n1969), .Z(n1970) );
  NAND U2781 ( .A(n27436), .B(n1970), .Z(n27437) );
  NANDN U2782 ( .A(n18519), .B(n4282), .Z(n1971) );
  AND U2783 ( .A(n13175), .B(n1971), .Z(n27200) );
  NOR U2784 ( .A(n19029), .B(n19030), .Z(n27496) );
  ANDN U2785 ( .B(n12929), .A(n12928), .Z(n24287) );
  NAND U2786 ( .A(n27528), .B(n27529), .Z(n1972) );
  NANDN U2787 ( .A(n27531), .B(n1972), .Z(n1973) );
  NAND U2788 ( .A(n27532), .B(n1973), .Z(n1974) );
  NAND U2789 ( .A(n27533), .B(n1974), .Z(n1975) );
  NAND U2790 ( .A(n27534), .B(n1975), .Z(n1976) );
  AND U2791 ( .A(n24281), .B(n1976), .Z(n1977) );
  NANDN U2792 ( .A(n1977), .B(n27535), .Z(n1978) );
  AND U2793 ( .A(n27536), .B(n1978), .Z(n1979) );
  NOR U2794 ( .A(n24280), .B(n1979), .Z(n1980) );
  NANDN U2795 ( .A(n24279), .B(n24278), .Z(n1981) );
  NAND U2796 ( .A(n1980), .B(n1981), .Z(n1982) );
  NANDN U2797 ( .A(n27537), .B(n1982), .Z(n1983) );
  NAND U2798 ( .A(n27538), .B(n1983), .Z(n1984) );
  ANDN U2799 ( .B(n1984), .A(n27539), .Z(n1985) );
  NANDN U2800 ( .A(n1985), .B(n24277), .Z(n1986) );
  ANDN U2801 ( .B(n1986), .A(n27540), .Z(n27541) );
  ANDN U2802 ( .B(n12854), .A(n12853), .Z(n27579) );
  NANDN U2803 ( .A(n12837), .B(n12838), .Z(n27598) );
  NAND U2804 ( .A(n27616), .B(n27617), .Z(n1987) );
  NAND U2805 ( .A(n24267), .B(n1987), .Z(n1988) );
  ANDN U2806 ( .B(n1988), .A(n27618), .Z(n1989) );
  NANDN U2807 ( .A(n1989), .B(n27619), .Z(n1990) );
  NANDN U2808 ( .A(n24266), .B(n1990), .Z(n1991) );
  NANDN U2809 ( .A(n27620), .B(n1991), .Z(n1992) );
  NANDN U2810 ( .A(n27621), .B(n1992), .Z(n1993) );
  NANDN U2811 ( .A(n24265), .B(n24264), .Z(n1994) );
  NAND U2812 ( .A(n1993), .B(n1994), .Z(n1995) );
  NANDN U2813 ( .A(n27623), .B(n27622), .Z(n1996) );
  AND U2814 ( .A(n27624), .B(n1996), .Z(n1997) );
  NANDN U2815 ( .A(n1995), .B(n24263), .Z(n1998) );
  NAND U2816 ( .A(n1997), .B(n1998), .Z(n1999) );
  NAND U2817 ( .A(n27625), .B(n1999), .Z(n2000) );
  AND U2818 ( .A(n27626), .B(n2000), .Z(n27629) );
  NAND U2819 ( .A(n27658), .B(n27659), .Z(n2001) );
  NANDN U2820 ( .A(n27660), .B(n2001), .Z(n2002) );
  NAND U2821 ( .A(n27661), .B(n2002), .Z(n2003) );
  NAND U2822 ( .A(n27662), .B(n2003), .Z(n2004) );
  NAND U2823 ( .A(n27663), .B(n2004), .Z(n2005) );
  ANDN U2824 ( .B(n2005), .A(n27664), .Z(n2006) );
  NANDN U2825 ( .A(n2006), .B(n27665), .Z(n2007) );
  NANDN U2826 ( .A(n27666), .B(n2007), .Z(n2008) );
  NAND U2827 ( .A(n27667), .B(n2008), .Z(n2009) );
  NAND U2828 ( .A(n27668), .B(n2009), .Z(n2010) );
  NANDN U2829 ( .A(n24257), .B(n2010), .Z(n2011) );
  AND U2830 ( .A(n24256), .B(n2011), .Z(n2012) );
  OR U2831 ( .A(n27669), .B(n2012), .Z(n2013) );
  NAND U2832 ( .A(n27670), .B(n2013), .Z(n2014) );
  NAND U2833 ( .A(n27671), .B(n2014), .Z(n2015) );
  NANDN U2834 ( .A(n27672), .B(n2015), .Z(n27673) );
  ANDN U2835 ( .B(n12753), .A(n12752), .Z(n27718) );
  ANDN U2836 ( .B(n12743), .A(n12742), .Z(n27742) );
  NANDN U2837 ( .A(n12963), .B(n4250), .Z(n2016) );
  AND U2838 ( .A(n18971), .B(n2016), .Z(n27459) );
  OR U2839 ( .A(n12717), .B(n12718), .Z(n2017) );
  ANDN U2840 ( .B(n2017), .A(n12719), .Z(n27784) );
  NAND U2841 ( .A(n18995), .B(n8634), .Z(n2018) );
  ANDN U2842 ( .B(n2018), .A(n18998), .Z(n27476) );
  NAND U2843 ( .A(n27809), .B(n27808), .Z(n2019) );
  NANDN U2844 ( .A(n27810), .B(n2019), .Z(n2020) );
  NAND U2845 ( .A(n27811), .B(n2020), .Z(n2021) );
  NANDN U2846 ( .A(n27812), .B(n2021), .Z(n2022) );
  NAND U2847 ( .A(n27813), .B(n2022), .Z(n2023) );
  ANDN U2848 ( .B(n2023), .A(n27814), .Z(n2024) );
  NANDN U2849 ( .A(n2024), .B(n27815), .Z(n2025) );
  ANDN U2850 ( .B(n2025), .A(n27816), .Z(n2026) );
  ANDN U2851 ( .B(n24243), .A(n2026), .Z(n2027) );
  NAND U2852 ( .A(n24244), .B(n2027), .Z(n2028) );
  AND U2853 ( .A(n27817), .B(n2028), .Z(n2029) );
  ANDN U2854 ( .B(n24241), .A(n27818), .Z(n2030) );
  OR U2855 ( .A(n24242), .B(n2029), .Z(n2031) );
  AND U2856 ( .A(n2030), .B(n2031), .Z(n2032) );
  NANDN U2857 ( .A(n2032), .B(n27819), .Z(n2033) );
  NANDN U2858 ( .A(n27820), .B(n2033), .Z(n2034) );
  NAND U2859 ( .A(n27821), .B(n2034), .Z(n2035) );
  NANDN U2860 ( .A(n27822), .B(n2035), .Z(n27823) );
  OR U2861 ( .A(n27858), .B(n27857), .Z(n2036) );
  NAND U2862 ( .A(n27859), .B(n2036), .Z(n2037) );
  NANDN U2863 ( .A(n27860), .B(n2037), .Z(n2038) );
  AND U2864 ( .A(n2038), .B(n27864), .Z(n2039) );
  NAND U2865 ( .A(n27863), .B(n27862), .Z(n2040) );
  AND U2866 ( .A(n2039), .B(n2040), .Z(n2041) );
  OR U2867 ( .A(n2041), .B(n27865), .Z(n2042) );
  NAND U2868 ( .A(n27866), .B(n2042), .Z(n2043) );
  NANDN U2869 ( .A(n27867), .B(n2043), .Z(n2044) );
  NAND U2870 ( .A(n27868), .B(n2044), .Z(n2045) );
  NAND U2871 ( .A(n27869), .B(n2045), .Z(n2046) );
  AND U2872 ( .A(n27870), .B(n2046), .Z(n2047) );
  NANDN U2873 ( .A(n2047), .B(n27871), .Z(n2048) );
  NAND U2874 ( .A(n27872), .B(n2048), .Z(n2049) );
  NANDN U2875 ( .A(n27873), .B(n2049), .Z(n2050) );
  NAND U2876 ( .A(n27874), .B(n2050), .Z(n2051) );
  NAND U2877 ( .A(n27875), .B(n2051), .Z(n2052) );
  AND U2878 ( .A(n27876), .B(n2052), .Z(n2053) );
  NAND U2879 ( .A(n27877), .B(n2053), .Z(n27878) );
  NANDN U2880 ( .A(n12872), .B(n4226), .Z(n2054) );
  AND U2881 ( .A(n19187), .B(n2054), .Z(n27568) );
  NANDN U2882 ( .A(n12642), .B(n12641), .Z(n2055) );
  ANDN U2883 ( .B(n2055), .A(n12643), .Z(n27907) );
  NANDN U2884 ( .A(n27922), .B(n27921), .Z(n2056) );
  NAND U2885 ( .A(n27923), .B(n2056), .Z(n2057) );
  ANDN U2886 ( .B(n2057), .A(n27924), .Z(n2058) );
  NANDN U2887 ( .A(n2058), .B(n27925), .Z(n2059) );
  NANDN U2888 ( .A(n27926), .B(n2059), .Z(n2060) );
  NAND U2889 ( .A(n27927), .B(n2060), .Z(n2061) );
  NANDN U2890 ( .A(n2061), .B(n24228), .Z(n2062) );
  NAND U2891 ( .A(n24227), .B(n2062), .Z(n2063) );
  NAND U2892 ( .A(n27928), .B(n2063), .Z(n2064) );
  NANDN U2893 ( .A(n27929), .B(n2064), .Z(n2065) );
  NAND U2894 ( .A(n27930), .B(n2065), .Z(n2066) );
  ANDN U2895 ( .B(n2066), .A(n27931), .Z(n2067) );
  OR U2896 ( .A(n27932), .B(n2067), .Z(n2068) );
  NAND U2897 ( .A(n27933), .B(n2068), .Z(n2069) );
  NANDN U2898 ( .A(n24226), .B(n2069), .Z(n27934) );
  ANDN U2899 ( .B(n12562), .A(n12561), .Z(n24214) );
  NANDN U2900 ( .A(n27969), .B(n27968), .Z(n2070) );
  NAND U2901 ( .A(n27970), .B(n2070), .Z(n2071) );
  ANDN U2902 ( .B(n2071), .A(n27971), .Z(n2072) );
  NANDN U2903 ( .A(n2072), .B(n27972), .Z(n2073) );
  ANDN U2904 ( .B(n2073), .A(n27973), .Z(n2074) );
  NANDN U2905 ( .A(n2074), .B(n27974), .Z(n2075) );
  NANDN U2906 ( .A(n24220), .B(n2075), .Z(n2076) );
  NANDN U2907 ( .A(n27975), .B(n2076), .Z(n2077) );
  NAND U2908 ( .A(n2077), .B(x[2582]), .Z(n2078) );
  AND U2909 ( .A(n27976), .B(n2078), .Z(n2079) );
  XOR U2910 ( .A(n2077), .B(x[2582]), .Z(n2080) );
  NANDN U2911 ( .A(y[2582]), .B(n2080), .Z(n2081) );
  AND U2912 ( .A(n2079), .B(n2081), .Z(n2082) );
  OR U2913 ( .A(n27977), .B(n2082), .Z(n2083) );
  NAND U2914 ( .A(n27978), .B(n2083), .Z(n2084) );
  NANDN U2915 ( .A(n27979), .B(n2084), .Z(n2085) );
  NANDN U2916 ( .A(n24219), .B(n2085), .Z(n27980) );
  AND U2917 ( .A(n28004), .B(n28003), .Z(n2086) );
  NANDN U2918 ( .A(n28007), .B(n28006), .Z(n2087) );
  NAND U2919 ( .A(n2086), .B(n2087), .Z(n2088) );
  NAND U2920 ( .A(n28008), .B(n2088), .Z(n2089) );
  NANDN U2921 ( .A(n28009), .B(n2089), .Z(n2090) );
  ANDN U2922 ( .B(n2090), .A(n28010), .Z(n2091) );
  NANDN U2923 ( .A(n2091), .B(n28011), .Z(n2092) );
  NANDN U2924 ( .A(n28012), .B(n2092), .Z(n2093) );
  NAND U2925 ( .A(n28013), .B(n2093), .Z(n2094) );
  NANDN U2926 ( .A(n28014), .B(n2094), .Z(n2095) );
  NAND U2927 ( .A(n28015), .B(n2095), .Z(n2096) );
  AND U2928 ( .A(n28016), .B(n2096), .Z(n2097) );
  OR U2929 ( .A(n28017), .B(n2097), .Z(n2098) );
  AND U2930 ( .A(n28018), .B(n2098), .Z(n2099) );
  OR U2931 ( .A(n2099), .B(n28019), .Z(n2100) );
  NAND U2932 ( .A(n28020), .B(n2100), .Z(n2101) );
  NAND U2933 ( .A(n28021), .B(n2101), .Z(n28022) );
  NANDN U2934 ( .A(n19484), .B(n9012), .Z(n2102) );
  AND U2935 ( .A(n12734), .B(n2102), .Z(n27758) );
  OR U2936 ( .A(n28054), .B(n28055), .Z(n2103) );
  NAND U2937 ( .A(n28056), .B(n2103), .Z(n2104) );
  NANDN U2938 ( .A(n28057), .B(n2104), .Z(n2105) );
  NAND U2939 ( .A(n28058), .B(n2105), .Z(n2106) );
  NAND U2940 ( .A(n28059), .B(n2106), .Z(n2107) );
  AND U2941 ( .A(n28060), .B(n2107), .Z(n2108) );
  NANDN U2942 ( .A(n2108), .B(n28061), .Z(n2109) );
  NAND U2943 ( .A(n28062), .B(n2109), .Z(n2110) );
  NANDN U2944 ( .A(n28063), .B(n2110), .Z(n2111) );
  NAND U2945 ( .A(n28064), .B(n2111), .Z(n2112) );
  NAND U2946 ( .A(n24200), .B(n2112), .Z(n2113) );
  AND U2947 ( .A(n28065), .B(n2113), .Z(n2114) );
  OR U2948 ( .A(n28066), .B(n2114), .Z(n2115) );
  NAND U2949 ( .A(n28067), .B(n2115), .Z(n2116) );
  NANDN U2950 ( .A(n28068), .B(n2116), .Z(n2117) );
  NAND U2951 ( .A(n28069), .B(n2117), .Z(n2118) );
  NANDN U2952 ( .A(n28070), .B(n2118), .Z(n2119) );
  AND U2953 ( .A(n28071), .B(n2119), .Z(n28073) );
  ANDN U2954 ( .B(n12502), .A(n12501), .Z(n28091) );
  NANDN U2955 ( .A(n24190), .B(n24189), .Z(n2120) );
  AND U2956 ( .A(n24192), .B(n2120), .Z(n2121) );
  NANDN U2957 ( .A(n28117), .B(n28116), .Z(n2122) );
  NAND U2958 ( .A(n2121), .B(n2122), .Z(n2123) );
  NAND U2959 ( .A(n28118), .B(n2123), .Z(n2124) );
  NAND U2960 ( .A(n28119), .B(n2124), .Z(n2125) );
  NAND U2961 ( .A(n24187), .B(n2125), .Z(n2126) );
  ANDN U2962 ( .B(n2126), .A(n24186), .Z(n2127) );
  ANDN U2963 ( .B(n28120), .A(n2127), .Z(n2128) );
  NAND U2964 ( .A(n28121), .B(n2128), .Z(n2129) );
  ANDN U2965 ( .B(n2129), .A(n28122), .Z(n2130) );
  NANDN U2966 ( .A(n2130), .B(n28123), .Z(n2131) );
  ANDN U2967 ( .B(n2131), .A(n28124), .Z(n2132) );
  OR U2968 ( .A(n28125), .B(n2132), .Z(n2133) );
  NANDN U2969 ( .A(n28126), .B(n2133), .Z(n2134) );
  NAND U2970 ( .A(n24185), .B(n2134), .Z(n28129) );
  ANDN U2971 ( .B(n12455), .A(n12454), .Z(n28142) );
  ANDN U2972 ( .B(n12447), .A(n12446), .Z(n28154) );
  NAND U2973 ( .A(n28196), .B(n28197), .Z(n2135) );
  ANDN U2974 ( .B(n2135), .A(n28198), .Z(n2136) );
  NAND U2975 ( .A(n28184), .B(n28183), .Z(n2137) );
  NANDN U2976 ( .A(n28186), .B(n2137), .Z(n2138) );
  NAND U2977 ( .A(n28187), .B(n2138), .Z(n2139) );
  NANDN U2978 ( .A(n28188), .B(n2139), .Z(n2140) );
  NANDN U2979 ( .A(n28189), .B(n2140), .Z(n2141) );
  AND U2980 ( .A(n28190), .B(n2141), .Z(n2142) );
  NANDN U2981 ( .A(n2142), .B(n28191), .Z(n2143) );
  NAND U2982 ( .A(n24169), .B(n2143), .Z(n2144) );
  NAND U2983 ( .A(n28192), .B(n2144), .Z(n2145) );
  NAND U2984 ( .A(n28193), .B(n2145), .Z(n2146) );
  NANDN U2985 ( .A(n28194), .B(n2146), .Z(n2147) );
  AND U2986 ( .A(n28195), .B(n2147), .Z(n2148) );
  NANDN U2987 ( .A(n2148), .B(n2136), .Z(n2149) );
  NAND U2988 ( .A(n28199), .B(n2149), .Z(n2150) );
  NANDN U2989 ( .A(n28200), .B(n2150), .Z(n28201) );
  NAND U2990 ( .A(n28226), .B(n28225), .Z(n2151) );
  NANDN U2991 ( .A(n28228), .B(n2151), .Z(n2152) );
  AND U2992 ( .A(n28229), .B(n2152), .Z(n2153) );
  ANDN U2993 ( .B(n24156), .A(n2153), .Z(n2154) );
  OR U2994 ( .A(n24155), .B(n24154), .Z(n2155) );
  NAND U2995 ( .A(n2154), .B(n2155), .Z(n2156) );
  AND U2996 ( .A(n2156), .B(n28232), .Z(n2157) );
  NAND U2997 ( .A(n28231), .B(n28230), .Z(n2158) );
  AND U2998 ( .A(n2157), .B(n2158), .Z(n2159) );
  NANDN U2999 ( .A(n2159), .B(n28233), .Z(n2160) );
  NAND U3000 ( .A(n28234), .B(n2160), .Z(n2161) );
  NAND U3001 ( .A(n28235), .B(n2161), .Z(n2162) );
  NAND U3002 ( .A(n28236), .B(n2162), .Z(n2163) );
  NAND U3003 ( .A(n28237), .B(n2163), .Z(n2164) );
  ANDN U3004 ( .B(n2164), .A(n28238), .Z(n2165) );
  NANDN U3005 ( .A(n2165), .B(n28239), .Z(n2166) );
  NANDN U3006 ( .A(n24153), .B(n2166), .Z(n2167) );
  NAND U3007 ( .A(n28240), .B(n2167), .Z(n28242) );
  NAND U3008 ( .A(n28296), .B(n28297), .Z(n2168) );
  NAND U3009 ( .A(n28298), .B(n2168), .Z(n2169) );
  NAND U3010 ( .A(n28299), .B(n2169), .Z(n2170) );
  NANDN U3011 ( .A(n28300), .B(n2170), .Z(n2171) );
  NAND U3012 ( .A(n28301), .B(n2171), .Z(n2172) );
  ANDN U3013 ( .B(n2172), .A(n28302), .Z(n2173) );
  NANDN U3014 ( .A(n2173), .B(n24151), .Z(n2174) );
  NANDN U3015 ( .A(n28303), .B(n2174), .Z(n2175) );
  NANDN U3016 ( .A(n28304), .B(n2175), .Z(n2176) );
  NAND U3017 ( .A(n28305), .B(n2176), .Z(n2177) );
  NANDN U3018 ( .A(n28306), .B(n2177), .Z(n2178) );
  AND U3019 ( .A(n28307), .B(n2178), .Z(n2179) );
  OR U3020 ( .A(n28308), .B(n2179), .Z(n2180) );
  AND U3021 ( .A(n28309), .B(n2180), .Z(n2181) );
  NANDN U3022 ( .A(n2181), .B(n28310), .Z(n2182) );
  NAND U3023 ( .A(n28311), .B(n2182), .Z(n2183) );
  NAND U3024 ( .A(n24150), .B(n2183), .Z(n28313) );
  OR U3025 ( .A(n28347), .B(n28348), .Z(n2184) );
  NANDN U3026 ( .A(n28349), .B(n2184), .Z(n2185) );
  AND U3027 ( .A(n28350), .B(n2185), .Z(n2186) );
  OR U3028 ( .A(n24146), .B(n2186), .Z(n2187) );
  NAND U3029 ( .A(n24145), .B(n2187), .Z(n2188) );
  NANDN U3030 ( .A(n28351), .B(n2188), .Z(n2189) );
  NAND U3031 ( .A(n28352), .B(n2189), .Z(n2190) );
  NANDN U3032 ( .A(n28353), .B(n2190), .Z(n2191) );
  AND U3033 ( .A(n28354), .B(n2191), .Z(n2192) );
  NANDN U3034 ( .A(n2192), .B(n28355), .Z(n2193) );
  NANDN U3035 ( .A(n24144), .B(n2193), .Z(n2194) );
  NAND U3036 ( .A(n24143), .B(n2194), .Z(n2195) );
  NAND U3037 ( .A(n28356), .B(n2195), .Z(n2196) );
  NANDN U3038 ( .A(n28357), .B(n2196), .Z(n2197) );
  AND U3039 ( .A(n28358), .B(n2197), .Z(n28360) );
  NAND U3040 ( .A(n28389), .B(n28390), .Z(n2198) );
  NANDN U3041 ( .A(n28391), .B(n2198), .Z(n2199) );
  NANDN U3042 ( .A(n28392), .B(n2199), .Z(n2200) );
  NAND U3043 ( .A(n28393), .B(n2200), .Z(n2201) );
  NAND U3044 ( .A(n28394), .B(n2201), .Z(n2202) );
  AND U3045 ( .A(n28395), .B(n2202), .Z(n2203) );
  NAND U3046 ( .A(n2203), .B(n28396), .Z(n2204) );
  NAND U3047 ( .A(n28397), .B(n2204), .Z(n2205) );
  AND U3048 ( .A(n28398), .B(n2205), .Z(n2206) );
  NANDN U3049 ( .A(n24135), .B(n24134), .Z(n2207) );
  ANDN U3050 ( .B(n2207), .A(n24136), .Z(n2208) );
  NANDN U3051 ( .A(n2206), .B(n28399), .Z(n2209) );
  NAND U3052 ( .A(n2208), .B(n2209), .Z(n2210) );
  NAND U3053 ( .A(n28400), .B(n2210), .Z(n2211) );
  NANDN U3054 ( .A(n24133), .B(n2211), .Z(n28401) );
  NANDN U3055 ( .A(n28425), .B(n28424), .Z(n2212) );
  NAND U3056 ( .A(n28426), .B(n2212), .Z(n2213) );
  NANDN U3057 ( .A(n28427), .B(n2213), .Z(n2214) );
  NAND U3058 ( .A(n28428), .B(n2214), .Z(n2215) );
  NANDN U3059 ( .A(n28429), .B(n2215), .Z(n2216) );
  AND U3060 ( .A(n28430), .B(n2216), .Z(n2217) );
  NAND U3061 ( .A(n28432), .B(n28431), .Z(n2218) );
  NAND U3062 ( .A(n2217), .B(n2218), .Z(n2219) );
  NANDN U3063 ( .A(n28433), .B(n2219), .Z(n2220) );
  NAND U3064 ( .A(n28434), .B(n2220), .Z(n2221) );
  NANDN U3065 ( .A(n28435), .B(n2221), .Z(n2222) );
  AND U3066 ( .A(n28436), .B(n2222), .Z(n2223) );
  OR U3067 ( .A(n28437), .B(n2223), .Z(n2224) );
  ANDN U3068 ( .B(n2224), .A(n28438), .Z(n2225) );
  NANDN U3069 ( .A(n2225), .B(n28439), .Z(n2226) );
  NAND U3070 ( .A(n28440), .B(n2226), .Z(n2227) );
  NAND U3071 ( .A(n28441), .B(n2227), .Z(n28442) );
  NOR U3072 ( .A(n12231), .B(n12232), .Z(n24116) );
  NAND U3073 ( .A(n24113), .B(n28473), .Z(n2228) );
  NANDN U3074 ( .A(n28474), .B(n2228), .Z(n2229) );
  NAND U3075 ( .A(n28475), .B(n2229), .Z(n2230) );
  NAND U3076 ( .A(n28476), .B(n2230), .Z(n2231) );
  NAND U3077 ( .A(n28477), .B(n2231), .Z(n2232) );
  AND U3078 ( .A(n24112), .B(n2232), .Z(n2233) );
  NANDN U3079 ( .A(n2233), .B(n28478), .Z(n2234) );
  NAND U3080 ( .A(n24111), .B(n2234), .Z(n2235) );
  NAND U3081 ( .A(n28479), .B(n2235), .Z(n2236) );
  NAND U3082 ( .A(n28480), .B(n2236), .Z(n2237) );
  NAND U3083 ( .A(n28481), .B(n2237), .Z(n2238) );
  AND U3084 ( .A(n28482), .B(n2238), .Z(n2239) );
  NANDN U3085 ( .A(n2239), .B(n28483), .Z(n2240) );
  NAND U3086 ( .A(n28484), .B(n2240), .Z(n2241) );
  NAND U3087 ( .A(n28485), .B(n2241), .Z(n28486) );
  AND U3088 ( .A(n28512), .B(n28513), .Z(n2242) );
  NAND U3089 ( .A(n28516), .B(n2242), .Z(n2243) );
  NAND U3090 ( .A(n28517), .B(n2243), .Z(n2244) );
  NANDN U3091 ( .A(n24103), .B(n2244), .Z(n2245) );
  NAND U3092 ( .A(n24102), .B(n2245), .Z(n2246) );
  ANDN U3093 ( .B(n2246), .A(n28518), .Z(n2247) );
  NANDN U3094 ( .A(n2247), .B(n28519), .Z(n2248) );
  NANDN U3095 ( .A(n28520), .B(n2248), .Z(n2249) );
  NAND U3096 ( .A(n28521), .B(n2249), .Z(n2250) );
  NAND U3097 ( .A(n24101), .B(n2250), .Z(n2251) );
  NAND U3098 ( .A(n28522), .B(n2251), .Z(n2252) );
  ANDN U3099 ( .B(n2252), .A(n28523), .Z(n2253) );
  NOR U3100 ( .A(n28524), .B(n2253), .Z(n2254) );
  NANDN U3101 ( .A(n28526), .B(n28525), .Z(n2255) );
  NAND U3102 ( .A(n2254), .B(n2255), .Z(n2256) );
  NAND U3103 ( .A(n28527), .B(n2256), .Z(n28528) );
  NANDN U3104 ( .A(n28560), .B(n28559), .Z(n2257) );
  NAND U3105 ( .A(n28561), .B(n2257), .Z(n2258) );
  AND U3106 ( .A(n28562), .B(n2258), .Z(n2259) );
  OR U3107 ( .A(n28563), .B(n2259), .Z(n2260) );
  NAND U3108 ( .A(n28564), .B(n2260), .Z(n2261) );
  NANDN U3109 ( .A(n28565), .B(n2261), .Z(n2262) );
  NAND U3110 ( .A(n28566), .B(n2262), .Z(n2263) );
  NAND U3111 ( .A(n28567), .B(n2263), .Z(n2264) );
  AND U3112 ( .A(n28568), .B(n2264), .Z(n2265) );
  OR U3113 ( .A(n2265), .B(n28569), .Z(n2266) );
  NAND U3114 ( .A(n28570), .B(n2266), .Z(n2267) );
  ANDN U3115 ( .B(n2267), .A(n28571), .Z(n2268) );
  NANDN U3116 ( .A(n2268), .B(n28572), .Z(n2269) );
  NANDN U3117 ( .A(n28573), .B(n2269), .Z(n2270) );
  NAND U3118 ( .A(n28574), .B(n2270), .Z(n2271) );
  NANDN U3119 ( .A(n24094), .B(n2271), .Z(n28575) );
  NANDN U3120 ( .A(n28600), .B(n28599), .Z(n2272) );
  NANDN U3121 ( .A(n24087), .B(n2272), .Z(n2273) );
  NAND U3122 ( .A(n28601), .B(n2273), .Z(n2274) );
  NANDN U3123 ( .A(n28602), .B(n2274), .Z(n2275) );
  NAND U3124 ( .A(n28603), .B(n2275), .Z(n2276) );
  ANDN U3125 ( .B(n2276), .A(n28604), .Z(n2277) );
  NANDN U3126 ( .A(n2277), .B(n28605), .Z(n2278) );
  NANDN U3127 ( .A(n28606), .B(n2278), .Z(n2279) );
  NAND U3128 ( .A(n28607), .B(n2279), .Z(n2280) );
  NAND U3129 ( .A(n28608), .B(n2280), .Z(n2281) );
  NANDN U3130 ( .A(n28609), .B(n2281), .Z(n2282) );
  AND U3131 ( .A(n28610), .B(n2282), .Z(n2283) );
  OR U3132 ( .A(n24086), .B(n2283), .Z(n2284) );
  NAND U3133 ( .A(n28611), .B(n2284), .Z(n2285) );
  NANDN U3134 ( .A(n28612), .B(n2285), .Z(n2286) );
  NANDN U3135 ( .A(n28613), .B(n2286), .Z(n28614) );
  NANDN U3136 ( .A(n28642), .B(n28641), .Z(n2287) );
  NANDN U3137 ( .A(n28643), .B(n2287), .Z(n2288) );
  AND U3138 ( .A(n28644), .B(n2288), .Z(n2289) );
  OR U3139 ( .A(n24078), .B(n2289), .Z(n2290) );
  NAND U3140 ( .A(n24077), .B(n2290), .Z(n2291) );
  NANDN U3141 ( .A(n28645), .B(n2291), .Z(n2292) );
  NAND U3142 ( .A(n28646), .B(n2292), .Z(n2293) );
  NANDN U3143 ( .A(n28647), .B(n2293), .Z(n2294) );
  AND U3144 ( .A(n28648), .B(n2294), .Z(n2295) );
  OR U3145 ( .A(n2295), .B(n28649), .Z(n2296) );
  NAND U3146 ( .A(n24076), .B(n2296), .Z(n2297) );
  AND U3147 ( .A(n28650), .B(n2297), .Z(n2298) );
  OR U3148 ( .A(n2298), .B(n28651), .Z(n2299) );
  NAND U3149 ( .A(n28652), .B(n2299), .Z(n2300) );
  NANDN U3150 ( .A(n28653), .B(n2300), .Z(n28654) );
  NAND U3151 ( .A(n28677), .B(n28678), .Z(n2301) );
  NANDN U3152 ( .A(n28679), .B(n2301), .Z(n2302) );
  NAND U3153 ( .A(n24067), .B(n2302), .Z(n2303) );
  NANDN U3154 ( .A(n28680), .B(n2303), .Z(n2304) );
  NAND U3155 ( .A(n28681), .B(n2304), .Z(n2305) );
  ANDN U3156 ( .B(n2305), .A(n24066), .Z(n2306) );
  NANDN U3157 ( .A(n2306), .B(n24065), .Z(n2307) );
  AND U3158 ( .A(n24064), .B(n2307), .Z(n2308) );
  OR U3159 ( .A(n28682), .B(n2308), .Z(n2309) );
  NAND U3160 ( .A(n28683), .B(n2309), .Z(n2310) );
  NANDN U3161 ( .A(n24063), .B(n2310), .Z(n28684) );
  NAND U3162 ( .A(n28708), .B(n28709), .Z(n2311) );
  NANDN U3163 ( .A(n28710), .B(n2311), .Z(n2312) );
  AND U3164 ( .A(n28711), .B(n2312), .Z(n2313) );
  OR U3165 ( .A(n2313), .B(n28712), .Z(n2314) );
  NAND U3166 ( .A(n24055), .B(n2314), .Z(n2315) );
  NANDN U3167 ( .A(n28713), .B(n2315), .Z(n2316) );
  NAND U3168 ( .A(n28714), .B(n2316), .Z(n2317) );
  NAND U3169 ( .A(n28715), .B(n2317), .Z(n2318) );
  ANDN U3170 ( .B(n2318), .A(n28716), .Z(n2319) );
  NANDN U3171 ( .A(n2319), .B(n24054), .Z(n2320) );
  NANDN U3172 ( .A(n28717), .B(n2320), .Z(n2321) );
  NAND U3173 ( .A(n28718), .B(n2321), .Z(n2322) );
  NANDN U3174 ( .A(n24053), .B(n2322), .Z(n28719) );
  OR U3175 ( .A(n28743), .B(n28744), .Z(n2323) );
  NAND U3176 ( .A(n28745), .B(n2323), .Z(n2324) );
  ANDN U3177 ( .B(n2324), .A(n28746), .Z(n2325) );
  NANDN U3178 ( .A(n2325), .B(n24042), .Z(n2326) );
  NAND U3179 ( .A(n28747), .B(n2326), .Z(n2327) );
  NANDN U3180 ( .A(n28748), .B(n2327), .Z(n2328) );
  NAND U3181 ( .A(n28749), .B(n2328), .Z(n2329) );
  NANDN U3182 ( .A(n28750), .B(n2329), .Z(n2330) );
  AND U3183 ( .A(n24041), .B(n2330), .Z(n2331) );
  OR U3184 ( .A(n28751), .B(n2331), .Z(n2332) );
  NAND U3185 ( .A(n28752), .B(n2332), .Z(n2333) );
  NAND U3186 ( .A(n28753), .B(n2333), .Z(n2334) );
  ANDN U3187 ( .B(n28756), .A(n28755), .Z(n2335) );
  NANDN U3188 ( .A(n28754), .B(n2334), .Z(n2336) );
  NAND U3189 ( .A(n2335), .B(n2336), .Z(n28759) );
  NANDN U3190 ( .A(n28782), .B(n28781), .Z(n2337) );
  NAND U3191 ( .A(n24032), .B(n2337), .Z(n2338) );
  ANDN U3192 ( .B(n2338), .A(n28783), .Z(n2339) );
  NANDN U3193 ( .A(n2339), .B(n28784), .Z(n2340) );
  NANDN U3194 ( .A(n24031), .B(n2340), .Z(n2341) );
  NAND U3195 ( .A(n24030), .B(n2341), .Z(n2342) );
  NAND U3196 ( .A(n28785), .B(n2342), .Z(n2343) );
  NAND U3197 ( .A(n24029), .B(n2343), .Z(n2344) );
  ANDN U3198 ( .B(n2344), .A(n28786), .Z(n2345) );
  OR U3199 ( .A(n28787), .B(n2345), .Z(n2346) );
  NAND U3200 ( .A(n28788), .B(n2346), .Z(n2347) );
  NANDN U3201 ( .A(n28789), .B(n2347), .Z(n2348) );
  NAND U3202 ( .A(n24028), .B(n2348), .Z(n28792) );
  NANDN U3203 ( .A(n28818), .B(n28817), .Z(n2349) );
  NAND U3204 ( .A(n28820), .B(n2349), .Z(n2350) );
  NAND U3205 ( .A(n28821), .B(n2350), .Z(n2351) );
  NANDN U3206 ( .A(n24019), .B(n2351), .Z(n2352) );
  NAND U3207 ( .A(n24018), .B(n2352), .Z(n2353) );
  ANDN U3208 ( .B(n2353), .A(n28822), .Z(n2354) );
  NANDN U3209 ( .A(n2354), .B(n28823), .Z(n2355) );
  ANDN U3210 ( .B(n2355), .A(n28824), .Z(n2356) );
  NANDN U3211 ( .A(n2356), .B(n28825), .Z(n2357) );
  NANDN U3212 ( .A(n24017), .B(n2357), .Z(n2358) );
  NAND U3213 ( .A(n24016), .B(n2358), .Z(n28826) );
  OR U3214 ( .A(n28846), .B(n28847), .Z(n2359) );
  NAND U3215 ( .A(n28848), .B(n2359), .Z(n2360) );
  NANDN U3216 ( .A(n28849), .B(n2360), .Z(n2361) );
  NAND U3217 ( .A(n24004), .B(n2361), .Z(n2362) );
  NAND U3218 ( .A(n28850), .B(n2362), .Z(n2363) );
  ANDN U3219 ( .B(n2363), .A(n28851), .Z(n2364) );
  NANDN U3220 ( .A(n2364), .B(n28852), .Z(n2365) );
  ANDN U3221 ( .B(n2365), .A(n28853), .Z(n2366) );
  NANDN U3222 ( .A(n2366), .B(n24003), .Z(n2367) );
  NANDN U3223 ( .A(n28854), .B(n2367), .Z(n2368) );
  NAND U3224 ( .A(n28855), .B(n2368), .Z(n2369) );
  ANDN U3225 ( .B(n24001), .A(n28856), .Z(n2370) );
  NANDN U3226 ( .A(n24002), .B(n2369), .Z(n2371) );
  NAND U3227 ( .A(n2370), .B(n2371), .Z(n28857) );
  NANDN U3228 ( .A(n28885), .B(n28884), .Z(n2372) );
  NAND U3229 ( .A(n28886), .B(n2372), .Z(n2373) );
  AND U3230 ( .A(n28887), .B(n2373), .Z(n2374) );
  AND U3231 ( .A(n23992), .B(n28888), .Z(n2375) );
  OR U3232 ( .A(n23993), .B(n2374), .Z(n2376) );
  AND U3233 ( .A(n2375), .B(n2376), .Z(n2377) );
  OR U3234 ( .A(n28889), .B(n2377), .Z(n2378) );
  AND U3235 ( .A(n28890), .B(n2378), .Z(n2379) );
  OR U3236 ( .A(n28891), .B(n2379), .Z(n2380) );
  NAND U3237 ( .A(n28892), .B(n2380), .Z(n2381) );
  NANDN U3238 ( .A(n23991), .B(n2381), .Z(n28893) );
  NANDN U3239 ( .A(n28920), .B(n28919), .Z(n2382) );
  NAND U3240 ( .A(n28921), .B(n2382), .Z(n2383) );
  NANDN U3241 ( .A(n28922), .B(n2383), .Z(n2384) );
  NAND U3242 ( .A(n23985), .B(n2384), .Z(n2385) );
  NANDN U3243 ( .A(n28923), .B(n2385), .Z(n2386) );
  AND U3244 ( .A(n28924), .B(n2386), .Z(n2387) );
  OR U3245 ( .A(n23984), .B(n2387), .Z(n2388) );
  NAND U3246 ( .A(n23983), .B(n2388), .Z(n2389) );
  NAND U3247 ( .A(n28925), .B(n2389), .Z(n2390) );
  AND U3248 ( .A(n23982), .B(n23981), .Z(n2391) );
  NANDN U3249 ( .A(n28926), .B(n2390), .Z(n2392) );
  NAND U3250 ( .A(n2391), .B(n2392), .Z(n2393) );
  NANDN U3251 ( .A(n28927), .B(n2393), .Z(n2394) );
  NAND U3252 ( .A(n28928), .B(n2394), .Z(n28929) );
  NANDN U3253 ( .A(n28957), .B(n28956), .Z(n2395) );
  NAND U3254 ( .A(n28958), .B(n2395), .Z(n2396) );
  ANDN U3255 ( .B(n2396), .A(n28959), .Z(n2397) );
  NANDN U3256 ( .A(n2397), .B(n23972), .Z(n2398) );
  NAND U3257 ( .A(n28960), .B(n2398), .Z(n2399) );
  NANDN U3258 ( .A(n28961), .B(n2399), .Z(n2400) );
  NAND U3259 ( .A(n28962), .B(n2400), .Z(n2401) );
  NANDN U3260 ( .A(n28963), .B(n2401), .Z(n2402) );
  AND U3261 ( .A(n28964), .B(n2402), .Z(n2403) );
  OR U3262 ( .A(n28965), .B(n2403), .Z(n2404) );
  NAND U3263 ( .A(n28966), .B(n2404), .Z(n2405) );
  NANDN U3264 ( .A(n28967), .B(n2405), .Z(n2406) );
  NAND U3265 ( .A(n28968), .B(n2406), .Z(n2407) );
  NANDN U3266 ( .A(n28969), .B(n2407), .Z(n2408) );
  AND U3267 ( .A(n28970), .B(n2408), .Z(n2409) );
  NANDN U3268 ( .A(n2409), .B(n28971), .Z(n2410) );
  NAND U3269 ( .A(n28972), .B(n2410), .Z(n2411) );
  NANDN U3270 ( .A(n28973), .B(n2411), .Z(n28974) );
  NAND U3271 ( .A(n29007), .B(n29006), .Z(n2412) );
  NAND U3272 ( .A(n23968), .B(n2412), .Z(n2413) );
  ANDN U3273 ( .B(n2413), .A(n29008), .Z(n2414) );
  NANDN U3274 ( .A(n2414), .B(n29009), .Z(n2415) );
  ANDN U3275 ( .B(n2415), .A(n23967), .Z(n2416) );
  NANDN U3276 ( .A(n2416), .B(n23966), .Z(n2417) );
  NAND U3277 ( .A(n29010), .B(n2417), .Z(n2418) );
  NANDN U3278 ( .A(n29011), .B(n2418), .Z(n2419) );
  ANDN U3279 ( .B(n23965), .A(n23964), .Z(n2420) );
  NAND U3280 ( .A(n2419), .B(n2420), .Z(n2421) );
  NANDN U3281 ( .A(n29012), .B(n2421), .Z(n2422) );
  NAND U3282 ( .A(n29013), .B(n2422), .Z(n2423) );
  NANDN U3283 ( .A(n29014), .B(n2423), .Z(n2424) );
  ANDN U3284 ( .B(n2424), .A(n29015), .Z(n29017) );
  NANDN U3285 ( .A(n29053), .B(n29052), .Z(n2425) );
  NANDN U3286 ( .A(n29054), .B(n2425), .Z(n2426) );
  AND U3287 ( .A(n29055), .B(n2426), .Z(n2427) );
  NAND U3288 ( .A(n2427), .B(n29056), .Z(n2428) );
  NANDN U3289 ( .A(n29057), .B(n2428), .Z(n2429) );
  AND U3290 ( .A(n29058), .B(n2429), .Z(n2430) );
  OR U3291 ( .A(n2430), .B(n29059), .Z(n2431) );
  NAND U3292 ( .A(n29060), .B(n2431), .Z(n2432) );
  NANDN U3293 ( .A(n29061), .B(n2432), .Z(n2433) );
  NAND U3294 ( .A(n29062), .B(n2433), .Z(n2434) );
  NAND U3295 ( .A(n29063), .B(n2434), .Z(n2435) );
  ANDN U3296 ( .B(n2435), .A(n29064), .Z(n2436) );
  NANDN U3297 ( .A(n2436), .B(n29065), .Z(n2437) );
  NANDN U3298 ( .A(n23960), .B(n2437), .Z(n2438) );
  NAND U3299 ( .A(n23959), .B(n2438), .Z(n29068) );
  OR U3300 ( .A(n29089), .B(n29090), .Z(n2439) );
  NAND U3301 ( .A(n29091), .B(n2439), .Z(n2440) );
  ANDN U3302 ( .B(n2440), .A(n29092), .Z(n2441) );
  NOR U3303 ( .A(n29093), .B(n29094), .Z(n2442) );
  NANDN U3304 ( .A(n2441), .B(n2442), .Z(n2443) );
  ANDN U3305 ( .B(n2443), .A(n29095), .Z(n2444) );
  NANDN U3306 ( .A(n2444), .B(n29096), .Z(n2445) );
  ANDN U3307 ( .B(n2445), .A(n29097), .Z(n2446) );
  NANDN U3308 ( .A(n2446), .B(n29098), .Z(n2447) );
  NANDN U3309 ( .A(n29099), .B(n2447), .Z(n2448) );
  NAND U3310 ( .A(n29100), .B(n2448), .Z(n2449) );
  AND U3311 ( .A(n23947), .B(n23948), .Z(n2450) );
  NANDN U3312 ( .A(n29101), .B(n2449), .Z(n2451) );
  NAND U3313 ( .A(n2450), .B(n2451), .Z(n2452) );
  AND U3314 ( .A(n29103), .B(n29104), .Z(n2453) );
  NANDN U3315 ( .A(n29102), .B(n2452), .Z(n2454) );
  NAND U3316 ( .A(n2453), .B(n2454), .Z(n29107) );
  NAND U3317 ( .A(n29134), .B(n29135), .Z(n2455) );
  NAND U3318 ( .A(n29136), .B(n2455), .Z(n2456) );
  NANDN U3319 ( .A(n23941), .B(n2456), .Z(n2457) );
  NAND U3320 ( .A(n23940), .B(n2457), .Z(n2458) );
  NANDN U3321 ( .A(n29137), .B(n2458), .Z(n2459) );
  AND U3322 ( .A(n29138), .B(n2459), .Z(n2460) );
  AND U3323 ( .A(n29141), .B(n29140), .Z(n2461) );
  OR U3324 ( .A(n29139), .B(n2460), .Z(n2462) );
  AND U3325 ( .A(n2461), .B(n2462), .Z(n2463) );
  OR U3326 ( .A(n29142), .B(n2463), .Z(n2464) );
  NAND U3327 ( .A(n29143), .B(n2464), .Z(n2465) );
  NANDN U3328 ( .A(n29144), .B(n2465), .Z(n2466) );
  NAND U3329 ( .A(n29145), .B(n2466), .Z(n2467) );
  NANDN U3330 ( .A(n29146), .B(n2467), .Z(n2468) );
  AND U3331 ( .A(n29147), .B(n2468), .Z(n29149) );
  OR U3332 ( .A(n29176), .B(n29177), .Z(n2469) );
  NANDN U3333 ( .A(n29178), .B(n2469), .Z(n2470) );
  NAND U3334 ( .A(n29179), .B(n2470), .Z(n2471) );
  NANDN U3335 ( .A(n23933), .B(n2471), .Z(n2472) );
  NAND U3336 ( .A(n23932), .B(n2472), .Z(n2473) );
  ANDN U3337 ( .B(n2473), .A(n29180), .Z(n2474) );
  NANDN U3338 ( .A(n2474), .B(n29181), .Z(n2475) );
  AND U3339 ( .A(n23931), .B(n2475), .Z(n2476) );
  OR U3340 ( .A(n29182), .B(n2476), .Z(n2477) );
  NAND U3341 ( .A(n29183), .B(n2477), .Z(n2478) );
  NANDN U3342 ( .A(n23930), .B(n2478), .Z(n29184) );
  NANDN U3343 ( .A(n29215), .B(n29214), .Z(n2479) );
  NANDN U3344 ( .A(n29216), .B(n2479), .Z(n2480) );
  ANDN U3345 ( .B(n2480), .A(n29217), .Z(n2481) );
  NANDN U3346 ( .A(n23924), .B(n2481), .Z(n2482) );
  NANDN U3347 ( .A(n29218), .B(n2482), .Z(n2483) );
  AND U3348 ( .A(n29219), .B(n2483), .Z(n2484) );
  OR U3349 ( .A(n29220), .B(n2484), .Z(n2485) );
  NAND U3350 ( .A(n29221), .B(n2485), .Z(n2486) );
  NANDN U3351 ( .A(n29222), .B(n2486), .Z(n2487) );
  NAND U3352 ( .A(n29223), .B(n2487), .Z(n2488) );
  NANDN U3353 ( .A(n29224), .B(n2488), .Z(n2489) );
  AND U3354 ( .A(n29225), .B(n2489), .Z(n2490) );
  OR U3355 ( .A(n29226), .B(n2490), .Z(n2491) );
  NAND U3356 ( .A(n29227), .B(n2491), .Z(n2492) );
  NANDN U3357 ( .A(n29228), .B(n2492), .Z(n2493) );
  AND U3358 ( .A(n29230), .B(n29229), .Z(n2494) );
  NAND U3359 ( .A(n2493), .B(n2494), .Z(n2495) );
  NAND U3360 ( .A(n29231), .B(n2495), .Z(n29232) );
  AND U3361 ( .A(n29266), .B(n29267), .Z(n29268) );
  NAND U3362 ( .A(n29294), .B(n29293), .Z(n2496) );
  NANDN U3363 ( .A(n29295), .B(n2496), .Z(n2497) );
  AND U3364 ( .A(n29296), .B(n2497), .Z(n2498) );
  OR U3365 ( .A(n2498), .B(n23906), .Z(n2499) );
  NAND U3366 ( .A(n29297), .B(n2499), .Z(n2500) );
  AND U3367 ( .A(n29298), .B(n2500), .Z(n2501) );
  OR U3368 ( .A(n2501), .B(n29299), .Z(n2502) );
  NAND U3369 ( .A(n29300), .B(n2502), .Z(n2503) );
  ANDN U3370 ( .B(n2503), .A(n29301), .Z(n2504) );
  NANDN U3371 ( .A(n2504), .B(n29302), .Z(n2505) );
  NANDN U3372 ( .A(n29303), .B(n2505), .Z(n2506) );
  NAND U3373 ( .A(n29304), .B(n2506), .Z(n2507) );
  NAND U3374 ( .A(n23905), .B(n2507), .Z(n2508) );
  NAND U3375 ( .A(n29305), .B(n2508), .Z(n2509) );
  ANDN U3376 ( .B(n2509), .A(n29306), .Z(n29307) );
  NANDN U3377 ( .A(n29333), .B(n29332), .Z(n2510) );
  NAND U3378 ( .A(n29334), .B(n2510), .Z(n2511) );
  NANDN U3379 ( .A(n29335), .B(n2511), .Z(n2512) );
  NAND U3380 ( .A(n29336), .B(n2512), .Z(n2513) );
  NANDN U3381 ( .A(n29337), .B(n2513), .Z(n2514) );
  AND U3382 ( .A(n29338), .B(n2514), .Z(n2515) );
  ANDN U3383 ( .B(n29340), .A(n29341), .Z(n2516) );
  OR U3384 ( .A(n29339), .B(n2515), .Z(n2517) );
  AND U3385 ( .A(n2516), .B(n2517), .Z(n2518) );
  OR U3386 ( .A(n29342), .B(n2518), .Z(n2519) );
  NAND U3387 ( .A(n29343), .B(n2519), .Z(n2520) );
  NANDN U3388 ( .A(n29344), .B(n2520), .Z(n2521) );
  NAND U3389 ( .A(n29345), .B(n2521), .Z(n2522) );
  NANDN U3390 ( .A(n29346), .B(n2522), .Z(n2523) );
  AND U3391 ( .A(n29347), .B(n2523), .Z(n2524) );
  OR U3392 ( .A(n29348), .B(n2524), .Z(n2525) );
  NAND U3393 ( .A(n29349), .B(n2525), .Z(n2526) );
  NANDN U3394 ( .A(n29350), .B(n2526), .Z(n2527) );
  AND U3395 ( .A(n29351), .B(n2527), .Z(n29353) );
  NAND U3396 ( .A(n29375), .B(n29376), .Z(n2528) );
  NAND U3397 ( .A(n29377), .B(n2528), .Z(n2529) );
  AND U3398 ( .A(n29378), .B(n2529), .Z(n2530) );
  NANDN U3399 ( .A(n2530), .B(n29379), .Z(n2531) );
  ANDN U3400 ( .B(n2531), .A(n29380), .Z(n2532) );
  ANDN U3401 ( .B(n23890), .A(n2532), .Z(n2533) );
  NAND U3402 ( .A(n23889), .B(n2533), .Z(n2534) );
  ANDN U3403 ( .B(n2534), .A(n29381), .Z(n2535) );
  NANDN U3404 ( .A(n2535), .B(n29382), .Z(n2536) );
  NANDN U3405 ( .A(n29383), .B(n2536), .Z(n2537) );
  NAND U3406 ( .A(n29384), .B(n2537), .Z(n2538) );
  NANDN U3407 ( .A(n29385), .B(n2538), .Z(n2539) );
  NAND U3408 ( .A(n29386), .B(n2539), .Z(n2540) );
  ANDN U3409 ( .B(n2540), .A(n29387), .Z(n2541) );
  NANDN U3410 ( .A(n2541), .B(n29388), .Z(n2542) );
  NANDN U3411 ( .A(n29389), .B(n2542), .Z(n2543) );
  NAND U3412 ( .A(n29390), .B(n2543), .Z(n2544) );
  NANDN U3413 ( .A(n29391), .B(n2544), .Z(n29392) );
  NAND U3414 ( .A(n29420), .B(n29419), .Z(n2545) );
  AND U3415 ( .A(n29423), .B(n2545), .Z(n2546) );
  NANDN U3416 ( .A(n29422), .B(n2546), .Z(n2547) );
  NAND U3417 ( .A(n23882), .B(n2547), .Z(n2548) );
  AND U3418 ( .A(n29424), .B(n2548), .Z(n2549) );
  NANDN U3419 ( .A(n29425), .B(n2549), .Z(n2550) );
  ANDN U3420 ( .B(n23880), .A(n23881), .Z(n2551) );
  NANDN U3421 ( .A(n29426), .B(n2550), .Z(n2552) );
  NAND U3422 ( .A(n2551), .B(n2552), .Z(n2553) );
  NOR U3423 ( .A(n29429), .B(n29428), .Z(n2554) );
  NANDN U3424 ( .A(n29427), .B(n2553), .Z(n2555) );
  NAND U3425 ( .A(n2554), .B(n2555), .Z(n2556) );
  NANDN U3426 ( .A(n29430), .B(n2556), .Z(n2557) );
  NAND U3427 ( .A(n29431), .B(n2557), .Z(n29432) );
  NANDN U3428 ( .A(n23875), .B(n29458), .Z(n2558) );
  NAND U3429 ( .A(n23874), .B(n2558), .Z(n2559) );
  ANDN U3430 ( .B(n2559), .A(n29459), .Z(n2560) );
  ANDN U3431 ( .B(n29461), .A(n2560), .Z(n2561) );
  NAND U3432 ( .A(n29460), .B(n2561), .Z(n2562) );
  ANDN U3433 ( .B(n2562), .A(n29462), .Z(n2563) );
  NANDN U3434 ( .A(n2563), .B(n29463), .Z(n2564) );
  ANDN U3435 ( .B(n2564), .A(n23873), .Z(n2565) );
  NANDN U3436 ( .A(n2565), .B(n23872), .Z(n2566) );
  NANDN U3437 ( .A(n29464), .B(n2566), .Z(n2567) );
  NAND U3438 ( .A(n29465), .B(n2567), .Z(n29468) );
  NANDN U3439 ( .A(n29471), .B(n11210), .Z(n2568) );
  NAND U3440 ( .A(n23869), .B(n2568), .Z(n2569) );
  NANDN U3441 ( .A(n29472), .B(n2569), .Z(n2570) );
  NAND U3442 ( .A(n29473), .B(n2570), .Z(n2571) );
  NANDN U3443 ( .A(n23868), .B(n2571), .Z(n2572) );
  AND U3444 ( .A(n23867), .B(n2572), .Z(n2573) );
  OR U3445 ( .A(n29474), .B(n2573), .Z(n2574) );
  NAND U3446 ( .A(n29477), .B(n2574), .Z(n2575) );
  NANDN U3447 ( .A(n29478), .B(n2575), .Z(n2576) );
  NAND U3448 ( .A(n29479), .B(n2576), .Z(n2577) );
  NANDN U3449 ( .A(n23866), .B(n2577), .Z(n2578) );
  AND U3450 ( .A(n23865), .B(n2578), .Z(n2579) );
  OR U3451 ( .A(n29480), .B(n2579), .Z(n2580) );
  AND U3452 ( .A(n29481), .B(n2580), .Z(n2581) );
  OR U3453 ( .A(n23864), .B(n2581), .Z(n2582) );
  NAND U3454 ( .A(n23863), .B(n2582), .Z(n2583) );
  NANDN U3455 ( .A(n11276), .B(n2583), .Z(n2584) );
  XNOR U3456 ( .A(y[4052]), .B(x[4052]), .Z(n2585) );
  NANDN U3457 ( .A(n2584), .B(n2585), .Z(n11212) );
  NAND U3458 ( .A(n29510), .B(n29509), .Z(n2586) );
  AND U3459 ( .A(n29512), .B(n2586), .Z(n2587) );
  NOR U3460 ( .A(n2587), .B(n23856), .Z(n2588) );
  NAND U3461 ( .A(n23855), .B(n2588), .Z(n2589) );
  ANDN U3462 ( .B(n2589), .A(n29513), .Z(n2590) );
  NOR U3463 ( .A(n29514), .B(n2590), .Z(n2591) );
  NAND U3464 ( .A(n29515), .B(n2591), .Z(n2592) );
  ANDN U3465 ( .B(n2592), .A(n29516), .Z(n2593) );
  NANDN U3466 ( .A(n2593), .B(n29517), .Z(n2594) );
  ANDN U3467 ( .B(n2594), .A(n23854), .Z(n2595) );
  NANDN U3468 ( .A(n2595), .B(n23853), .Z(n2596) );
  NANDN U3469 ( .A(n29518), .B(n2596), .Z(n2597) );
  NAND U3470 ( .A(n29519), .B(n2597), .Z(n29520) );
  NANDN U3471 ( .A(n15485), .B(n15486), .Z(n24545) );
  NANDN U3472 ( .A(n15477), .B(n15478), .Z(n24553) );
  NANDN U3473 ( .A(n15437), .B(n15438), .Z(n24593) );
  NANDN U3474 ( .A(n15397), .B(n15398), .Z(n24633) );
  NANDN U3475 ( .A(y[69]), .B(x[69]), .Z(n2598) );
  ANDN U3476 ( .B(n2598), .A(n15366), .Z(n24672) );
  NANDN U3477 ( .A(n15334), .B(n15335), .Z(n24713) );
  ANDN U3478 ( .B(n15297), .A(n15296), .Z(n24755) );
  ANDN U3479 ( .B(n15256), .A(n15255), .Z(n24795) );
  ANDN U3480 ( .B(n15222), .A(n15221), .Z(n24835) );
  NANDN U3481 ( .A(x[170]), .B(y[170]), .Z(n2599) );
  ANDN U3482 ( .B(n2599), .A(n15181), .Z(n24875) );
  ANDN U3483 ( .B(n15139), .A(n15138), .Z(n24915) );
  ANDN U3484 ( .B(n15100), .A(n15099), .Z(n24955) );
  ANDN U3485 ( .B(n15060), .A(n15059), .Z(n24995) );
  ANDN U3486 ( .B(n15021), .A(n15020), .Z(n25035) );
  ANDN U3487 ( .B(n14968), .A(n14967), .Z(n25103) );
  ANDN U3488 ( .B(n14954), .A(n14953), .Z(n25115) );
  ANDN U3489 ( .B(n14881), .A(n14880), .Z(n25191) );
  NANDN U3490 ( .A(n25233), .B(n25232), .Z(n2600) );
  AND U3491 ( .A(n25234), .B(n2600), .Z(n2601) );
  ANDN U3492 ( .B(n25235), .A(n2601), .Z(n2602) );
  NAND U3493 ( .A(n25236), .B(n2602), .Z(n2603) );
  AND U3494 ( .A(n25237), .B(n2603), .Z(n2604) );
  OR U3495 ( .A(n2604), .B(n25238), .Z(n2605) );
  NAND U3496 ( .A(n25239), .B(n2605), .Z(n2606) );
  NANDN U3497 ( .A(n25240), .B(n2606), .Z(n2607) );
  NAND U3498 ( .A(n25241), .B(n2607), .Z(n2608) );
  NANDN U3499 ( .A(n25242), .B(n2608), .Z(n2609) );
  AND U3500 ( .A(n25243), .B(n2609), .Z(n2610) );
  OR U3501 ( .A(n2610), .B(n25244), .Z(n2611) );
  NAND U3502 ( .A(n25245), .B(n2611), .Z(n2612) );
  ANDN U3503 ( .B(n2612), .A(n25246), .Z(n2613) );
  NANDN U3504 ( .A(n2613), .B(n25247), .Z(n2614) );
  ANDN U3505 ( .B(n2614), .A(n25248), .Z(n2615) );
  NANDN U3506 ( .A(n2615), .B(n25249), .Z(n2616) );
  NANDN U3507 ( .A(n25250), .B(n2616), .Z(n2617) );
  NAND U3508 ( .A(n25251), .B(n2617), .Z(n25252) );
  NANDN U3509 ( .A(n14774), .B(n14775), .Z(n25293) );
  NANDN U3510 ( .A(n14754), .B(n14755), .Z(n25333) );
  NANDN U3511 ( .A(n14692), .B(n14693), .Z(n25405) );
  NANDN U3512 ( .A(n14684), .B(n14685), .Z(n25413) );
  NANDN U3513 ( .A(n14644), .B(n14645), .Z(n25453) );
  ANDN U3514 ( .B(n25533), .A(n25532), .Z(n2618) );
  NAND U3515 ( .A(n24539), .B(n2618), .Z(n2619) );
  AND U3516 ( .A(n25534), .B(n2619), .Z(n2620) );
  OR U3517 ( .A(n2620), .B(n25535), .Z(n2621) );
  NAND U3518 ( .A(n25536), .B(n2621), .Z(n2622) );
  NANDN U3519 ( .A(n25537), .B(n2622), .Z(n2623) );
  NAND U3520 ( .A(n25538), .B(n2623), .Z(n2624) );
  NANDN U3521 ( .A(n25539), .B(n2624), .Z(n2625) );
  AND U3522 ( .A(n25540), .B(n2625), .Z(n2626) );
  OR U3523 ( .A(n2626), .B(n25541), .Z(n2627) );
  NAND U3524 ( .A(n25542), .B(n2627), .Z(n2628) );
  NANDN U3525 ( .A(n25543), .B(n2628), .Z(n2629) );
  NAND U3526 ( .A(n25544), .B(n2629), .Z(n2630) );
  NANDN U3527 ( .A(n25545), .B(n2630), .Z(n2631) );
  AND U3528 ( .A(n25546), .B(n2631), .Z(n2632) );
  OR U3529 ( .A(n2632), .B(n25547), .Z(n2633) );
  NAND U3530 ( .A(n25548), .B(n2633), .Z(n2634) );
  NANDN U3531 ( .A(n25549), .B(n2634), .Z(n2635) );
  NAND U3532 ( .A(n25550), .B(n2635), .Z(n25551) );
  OR U3533 ( .A(n25632), .B(n25631), .Z(n2636) );
  NAND U3534 ( .A(n25633), .B(n2636), .Z(n2637) );
  NAND U3535 ( .A(n24538), .B(n2637), .Z(n2638) );
  OR U3536 ( .A(n2638), .B(n25634), .Z(n2639) );
  NAND U3537 ( .A(n25635), .B(n2639), .Z(n2640) );
  NANDN U3538 ( .A(n25636), .B(n2640), .Z(n2641) );
  NAND U3539 ( .A(n25637), .B(n2641), .Z(n2642) );
  NANDN U3540 ( .A(n25638), .B(n2642), .Z(n2643) );
  AND U3541 ( .A(n25639), .B(n2643), .Z(n2644) );
  OR U3542 ( .A(n25640), .B(n2644), .Z(n2645) );
  NAND U3543 ( .A(n25641), .B(n2645), .Z(n2646) );
  NANDN U3544 ( .A(n25642), .B(n2646), .Z(n2647) );
  NAND U3545 ( .A(n25643), .B(n2647), .Z(n2648) );
  NANDN U3546 ( .A(n25644), .B(n2648), .Z(n2649) );
  AND U3547 ( .A(n25645), .B(n2649), .Z(n2650) );
  NOR U3548 ( .A(n25647), .B(n2650), .Z(n2651) );
  NAND U3549 ( .A(n25646), .B(n2651), .Z(n2652) );
  AND U3550 ( .A(n25648), .B(n2652), .Z(n25649) );
  NANDN U3551 ( .A(n14391), .B(n14392), .Z(n25690) );
  NANDN U3552 ( .A(n14351), .B(n14352), .Z(n25730) );
  NANDN U3553 ( .A(n14311), .B(n14312), .Z(n25770) );
  NANDN U3554 ( .A(n25850), .B(n25849), .Z(n2653) );
  NAND U3555 ( .A(n25851), .B(n2653), .Z(n2654) );
  NANDN U3556 ( .A(n25852), .B(n2654), .Z(n2655) );
  NAND U3557 ( .A(n25853), .B(n2655), .Z(n2656) );
  NAND U3558 ( .A(n25854), .B(n2656), .Z(n2657) );
  ANDN U3559 ( .B(n2657), .A(n24537), .Z(n2658) );
  NANDN U3560 ( .A(n2658), .B(n25855), .Z(n2659) );
  NANDN U3561 ( .A(n25856), .B(n2659), .Z(n2660) );
  NAND U3562 ( .A(n25857), .B(n2660), .Z(n2661) );
  NAND U3563 ( .A(n25858), .B(n2661), .Z(n2662) );
  NAND U3564 ( .A(n24536), .B(n2662), .Z(n2663) );
  AND U3565 ( .A(n25859), .B(n2663), .Z(n2664) );
  NANDN U3566 ( .A(n2664), .B(n24535), .Z(n2665) );
  NAND U3567 ( .A(n25860), .B(n2665), .Z(n2666) );
  NAND U3568 ( .A(n25861), .B(n2666), .Z(n2667) );
  NAND U3569 ( .A(n25862), .B(n2667), .Z(n25863) );
  NANDN U3570 ( .A(n25886), .B(n25885), .Z(n2668) );
  NAND U3571 ( .A(n25887), .B(n2668), .Z(n2669) );
  NAND U3572 ( .A(n25888), .B(n2669), .Z(n2670) );
  NAND U3573 ( .A(n25889), .B(n2670), .Z(n2671) );
  NAND U3574 ( .A(n24526), .B(n2671), .Z(n2672) );
  AND U3575 ( .A(n25890), .B(n2672), .Z(n2673) );
  NANDN U3576 ( .A(n2673), .B(n25891), .Z(n2674) );
  NAND U3577 ( .A(n25892), .B(n2674), .Z(n2675) );
  NAND U3578 ( .A(n24525), .B(n2675), .Z(n2676) );
  NAND U3579 ( .A(n25893), .B(n2676), .Z(n2677) );
  NAND U3580 ( .A(n24524), .B(n2677), .Z(n2678) );
  AND U3581 ( .A(n25894), .B(n2678), .Z(n2679) );
  NANDN U3582 ( .A(n2679), .B(n25895), .Z(n2680) );
  NANDN U3583 ( .A(n24523), .B(n2680), .Z(n2681) );
  NAND U3584 ( .A(n25896), .B(n2681), .Z(n25897) );
  ANDN U3585 ( .B(n14125), .A(n14124), .Z(n25912) );
  NAND U3586 ( .A(n25933), .B(n25932), .Z(n2682) );
  NAND U3587 ( .A(n25934), .B(n2682), .Z(n2683) );
  AND U3588 ( .A(n25935), .B(n2683), .Z(n2684) );
  NANDN U3589 ( .A(n2684), .B(n25936), .Z(n2685) );
  NANDN U3590 ( .A(n25937), .B(n2685), .Z(n2686) );
  NAND U3591 ( .A(n25938), .B(n2686), .Z(n2687) );
  NANDN U3592 ( .A(n25939), .B(n2687), .Z(n2688) );
  NAND U3593 ( .A(n25940), .B(n2688), .Z(n2689) );
  ANDN U3594 ( .B(n2689), .A(n25941), .Z(n2690) );
  NANDN U3595 ( .A(n2690), .B(n25942), .Z(n2691) );
  NANDN U3596 ( .A(n25943), .B(n2691), .Z(n2692) );
  NAND U3597 ( .A(n25944), .B(n2692), .Z(n2693) );
  NANDN U3598 ( .A(n25945), .B(n2693), .Z(n2694) );
  NAND U3599 ( .A(n25946), .B(n2694), .Z(n2695) );
  ANDN U3600 ( .B(n2695), .A(n25947), .Z(n2696) );
  NANDN U3601 ( .A(n2696), .B(n25948), .Z(n2697) );
  NANDN U3602 ( .A(n25949), .B(n2697), .Z(n2698) );
  NAND U3603 ( .A(n25950), .B(n2698), .Z(n2699) );
  NANDN U3604 ( .A(n25951), .B(n2699), .Z(n25952) );
  NAND U3605 ( .A(n26032), .B(n26033), .Z(n2700) );
  NANDN U3606 ( .A(n26034), .B(n2700), .Z(n2701) );
  NAND U3607 ( .A(n26035), .B(n2701), .Z(n2702) );
  NANDN U3608 ( .A(n26036), .B(n2702), .Z(n2703) );
  NAND U3609 ( .A(n26037), .B(n2703), .Z(n2704) );
  AND U3610 ( .A(n26038), .B(n2704), .Z(n2705) );
  NANDN U3611 ( .A(n2705), .B(n26039), .Z(n2706) );
  NAND U3612 ( .A(n26040), .B(n2706), .Z(n2707) );
  NAND U3613 ( .A(n26041), .B(n2707), .Z(n2708) );
  NANDN U3614 ( .A(n26042), .B(n2708), .Z(n2709) );
  NAND U3615 ( .A(n26043), .B(n2709), .Z(n2710) );
  ANDN U3616 ( .B(n2710), .A(n24509), .Z(n2711) );
  NANDN U3617 ( .A(n2711), .B(n24508), .Z(n2712) );
  AND U3618 ( .A(n26044), .B(n2712), .Z(n2713) );
  NANDN U3619 ( .A(n2713), .B(n26045), .Z(n2714) );
  NANDN U3620 ( .A(n26046), .B(n2714), .Z(n2715) );
  NANDN U3621 ( .A(n26047), .B(n2715), .Z(n26048) );
  NAND U3622 ( .A(n26081), .B(n26080), .Z(n2716) );
  NAND U3623 ( .A(n26082), .B(n2716), .Z(n2717) );
  ANDN U3624 ( .B(n2717), .A(n24502), .Z(n2718) );
  OR U3625 ( .A(n26083), .B(n2718), .Z(n2719) );
  NAND U3626 ( .A(n26084), .B(n2719), .Z(n2720) );
  NAND U3627 ( .A(n26085), .B(n2720), .Z(n2721) );
  NANDN U3628 ( .A(n26086), .B(n2721), .Z(n2722) );
  NAND U3629 ( .A(n26087), .B(n2722), .Z(n2723) );
  AND U3630 ( .A(n26088), .B(n2723), .Z(n2724) );
  NANDN U3631 ( .A(n2724), .B(n26089), .Z(n2725) );
  NANDN U3632 ( .A(n24501), .B(n2725), .Z(n2726) );
  NAND U3633 ( .A(n26090), .B(n2726), .Z(n2727) );
  NAND U3634 ( .A(n26091), .B(n2727), .Z(n2728) );
  NAND U3635 ( .A(n24500), .B(n2728), .Z(n2729) );
  AND U3636 ( .A(n26092), .B(n2729), .Z(n26095) );
  NOR U3637 ( .A(n16564), .B(n16565), .Z(n26110) );
  NAND U3638 ( .A(n26134), .B(n24488), .Z(n2730) );
  NANDN U3639 ( .A(n26135), .B(n2730), .Z(n2731) );
  AND U3640 ( .A(n26136), .B(n2731), .Z(n2732) );
  OR U3641 ( .A(n26137), .B(n2732), .Z(n2733) );
  NAND U3642 ( .A(n26138), .B(n2733), .Z(n2734) );
  NANDN U3643 ( .A(n26139), .B(n2734), .Z(n2735) );
  NANDN U3644 ( .A(n24487), .B(n2735), .Z(n2736) );
  NAND U3645 ( .A(n26140), .B(n2736), .Z(n2737) );
  AND U3646 ( .A(n26141), .B(n2737), .Z(n2738) );
  OR U3647 ( .A(n26142), .B(n2738), .Z(n2739) );
  AND U3648 ( .A(n26143), .B(n2739), .Z(n2740) );
  ANDN U3649 ( .B(n26146), .A(n26145), .Z(n2741) );
  NANDN U3650 ( .A(n2740), .B(n26144), .Z(n2742) );
  AND U3651 ( .A(n2741), .B(n2742), .Z(n2743) );
  OR U3652 ( .A(n2743), .B(n26147), .Z(n2744) );
  NAND U3653 ( .A(n26148), .B(n2744), .Z(n2745) );
  NANDN U3654 ( .A(n26149), .B(n2745), .Z(n26150) );
  NAND U3655 ( .A(n13869), .B(n13870), .Z(n2746) );
  ANDN U3656 ( .B(n2746), .A(n13871), .Z(n26201) );
  NAND U3657 ( .A(n26260), .B(n26259), .Z(n2747) );
  NAND U3658 ( .A(n26261), .B(n2747), .Z(n2748) );
  NANDN U3659 ( .A(n26262), .B(n2748), .Z(n2749) );
  NAND U3660 ( .A(n26263), .B(n2749), .Z(n2750) );
  NANDN U3661 ( .A(n26264), .B(n2750), .Z(n2751) );
  AND U3662 ( .A(n26265), .B(n2751), .Z(n2752) );
  NANDN U3663 ( .A(n2752), .B(n26266), .Z(n2753) );
  NANDN U3664 ( .A(n26267), .B(n2753), .Z(n2754) );
  NAND U3665 ( .A(n26268), .B(n2754), .Z(n2755) );
  NAND U3666 ( .A(n26269), .B(n2755), .Z(n2756) );
  NAND U3667 ( .A(n26270), .B(n2756), .Z(n2757) );
  AND U3668 ( .A(n26271), .B(n2757), .Z(n2758) );
  NANDN U3669 ( .A(n2758), .B(n24469), .Z(n2759) );
  ANDN U3670 ( .B(n2759), .A(n24468), .Z(n2760) );
  NANDN U3671 ( .A(n2760), .B(n26272), .Z(n2761) );
  NAND U3672 ( .A(n26273), .B(n2761), .Z(n2762) );
  NAND U3673 ( .A(n26274), .B(n2762), .Z(n26275) );
  NAND U3674 ( .A(n26321), .B(n26320), .Z(n2763) );
  NANDN U3675 ( .A(n26322), .B(n2763), .Z(n2764) );
  AND U3676 ( .A(n26323), .B(n2764), .Z(n2765) );
  OR U3677 ( .A(n26324), .B(n2765), .Z(n2766) );
  NANDN U3678 ( .A(n26325), .B(n2766), .Z(n2767) );
  NANDN U3679 ( .A(n26326), .B(n2767), .Z(n2768) );
  NAND U3680 ( .A(n26327), .B(n2768), .Z(n2769) );
  NANDN U3681 ( .A(n24458), .B(n2769), .Z(n2770) );
  AND U3682 ( .A(n24457), .B(n2770), .Z(n2771) );
  NANDN U3683 ( .A(n2771), .B(n26328), .Z(n2772) );
  NAND U3684 ( .A(n24456), .B(n2772), .Z(n2773) );
  NANDN U3685 ( .A(n26329), .B(n2773), .Z(n2774) );
  NAND U3686 ( .A(n26330), .B(n2774), .Z(n26331) );
  NAND U3687 ( .A(n16707), .B(n16711), .Z(n2775) );
  AND U3688 ( .A(n4663), .B(n2775), .Z(n2776) );
  NAND U3689 ( .A(n2776), .B(n16715), .Z(n2777) );
  AND U3690 ( .A(n16710), .B(n2777), .Z(n24484) );
  NAND U3691 ( .A(n26376), .B(n26375), .Z(n2778) );
  NAND U3692 ( .A(n26377), .B(n2778), .Z(n2779) );
  NAND U3693 ( .A(n26378), .B(n2779), .Z(n2780) );
  NAND U3694 ( .A(n26379), .B(n2780), .Z(n2781) );
  NANDN U3695 ( .A(n24445), .B(n2781), .Z(n2782) );
  AND U3696 ( .A(n26380), .B(n2782), .Z(n2783) );
  OR U3697 ( .A(n2783), .B(n26381), .Z(n2784) );
  NAND U3698 ( .A(n26382), .B(n2784), .Z(n2785) );
  NAND U3699 ( .A(n26383), .B(n2785), .Z(n2786) );
  NAND U3700 ( .A(n26384), .B(n2786), .Z(n2787) );
  NAND U3701 ( .A(n26385), .B(n2787), .Z(n2788) );
  ANDN U3702 ( .B(n2788), .A(n26386), .Z(n2789) );
  NANDN U3703 ( .A(n2789), .B(n26387), .Z(n2790) );
  ANDN U3704 ( .B(n2790), .A(n26388), .Z(n2791) );
  OR U3705 ( .A(n2791), .B(n26389), .Z(n2792) );
  NAND U3706 ( .A(n26390), .B(n2792), .Z(n2793) );
  NAND U3707 ( .A(n26391), .B(n2793), .Z(n26392) );
  NANDN U3708 ( .A(n16749), .B(n16751), .Z(n2794) );
  AND U3709 ( .A(n16756), .B(n2794), .Z(n26204) );
  AND U3710 ( .A(n16810), .B(n16805), .Z(n2795) );
  NANDN U3711 ( .A(n16800), .B(n4645), .Z(n2796) );
  AND U3712 ( .A(n2795), .B(n2796), .Z(n26228) );
  NANDN U3713 ( .A(n26446), .B(n26445), .Z(n2797) );
  NAND U3714 ( .A(n26447), .B(n2797), .Z(n2798) );
  NANDN U3715 ( .A(n26448), .B(n2798), .Z(n2799) );
  NANDN U3716 ( .A(n26449), .B(n2799), .Z(n2800) );
  NAND U3717 ( .A(n26450), .B(n2800), .Z(n2801) );
  ANDN U3718 ( .B(n2801), .A(n24437), .Z(n2802) );
  NANDN U3719 ( .A(n2802), .B(n26451), .Z(n2803) );
  ANDN U3720 ( .B(n2803), .A(n26452), .Z(n2804) );
  ANDN U3721 ( .B(n26453), .A(n2804), .Z(n2805) );
  NAND U3722 ( .A(n26454), .B(n2805), .Z(n2806) );
  ANDN U3723 ( .B(n2806), .A(n26455), .Z(n2807) );
  NANDN U3724 ( .A(n2807), .B(n26456), .Z(n2808) );
  ANDN U3725 ( .B(n2808), .A(n26457), .Z(n2809) );
  NANDN U3726 ( .A(n2809), .B(n26458), .Z(n2810) );
  NANDN U3727 ( .A(n26459), .B(n2810), .Z(n2811) );
  NAND U3728 ( .A(n26460), .B(n2811), .Z(n26461) );
  NANDN U3729 ( .A(n16823), .B(n6850), .Z(n2812) );
  AND U3730 ( .A(n16828), .B(n2812), .Z(n26236) );
  NAND U3731 ( .A(n26487), .B(n26488), .Z(n2813) );
  NANDN U3732 ( .A(n24427), .B(n2813), .Z(n2814) );
  NANDN U3733 ( .A(n26489), .B(n2814), .Z(n2815) );
  NAND U3734 ( .A(n26490), .B(n2815), .Z(n2816) );
  NANDN U3735 ( .A(n26491), .B(n2816), .Z(n2817) );
  AND U3736 ( .A(n26492), .B(n2817), .Z(n2818) );
  OR U3737 ( .A(n26493), .B(n2818), .Z(n2819) );
  NAND U3738 ( .A(n26494), .B(n2819), .Z(n2820) );
  NAND U3739 ( .A(n24426), .B(n2820), .Z(n2821) );
  NAND U3740 ( .A(n26495), .B(n2821), .Z(n2822) );
  NAND U3741 ( .A(n26496), .B(n2822), .Z(n2823) );
  AND U3742 ( .A(n26497), .B(n2823), .Z(n2824) );
  OR U3743 ( .A(n26498), .B(n2824), .Z(n2825) );
  AND U3744 ( .A(n26499), .B(n2825), .Z(n2826) );
  OR U3745 ( .A(n26500), .B(n2826), .Z(n2827) );
  NAND U3746 ( .A(n26501), .B(n2827), .Z(n2828) );
  NANDN U3747 ( .A(n26502), .B(n2828), .Z(n26503) );
  AND U3748 ( .A(n6943), .B(n24462), .Z(n2829) );
  NAND U3749 ( .A(n26289), .B(n2829), .Z(n2830) );
  ANDN U3750 ( .B(n2830), .A(n13795), .Z(n2831) );
  ANDN U3751 ( .B(n13794), .A(n2831), .Z(n2832) );
  NAND U3752 ( .A(n24461), .B(n2832), .Z(n2833) );
  AND U3753 ( .A(n26292), .B(n2833), .Z(n2834) );
  OR U3754 ( .A(n2834), .B(n13791), .Z(n2835) );
  ANDN U3755 ( .B(n2835), .A(n13788), .Z(n2836) );
  NOR U3756 ( .A(n13786), .B(n2836), .Z(n2837) );
  NAND U3757 ( .A(n13792), .B(n2837), .Z(n2838) );
  AND U3758 ( .A(n16944), .B(n2838), .Z(n2839) );
  AND U3759 ( .A(n26297), .B(n13787), .Z(n2840) );
  NAND U3760 ( .A(n13790), .B(n2839), .Z(n2841) );
  AND U3761 ( .A(n2840), .B(n2841), .Z(n2842) );
  OR U3762 ( .A(n2842), .B(n26298), .Z(n2843) );
  AND U3763 ( .A(n26299), .B(n2843), .Z(n2844) );
  NANDN U3764 ( .A(n2844), .B(n26300), .Z(n2845) );
  NAND U3765 ( .A(n24460), .B(n2845), .Z(n2846) );
  NANDN U3766 ( .A(n26301), .B(n2846), .Z(n6954) );
  NANDN U3767 ( .A(n26545), .B(n26546), .Z(n2847) );
  NAND U3768 ( .A(n26547), .B(n2847), .Z(n2848) );
  ANDN U3769 ( .B(n2848), .A(n24416), .Z(n2849) );
  NANDN U3770 ( .A(n2849), .B(n24415), .Z(n2850) );
  NAND U3771 ( .A(n26548), .B(n2850), .Z(n2851) );
  NANDN U3772 ( .A(n24414), .B(n2851), .Z(n2852) );
  NAND U3773 ( .A(n26549), .B(n2852), .Z(n2853) );
  NAND U3774 ( .A(n26550), .B(n2853), .Z(n2854) );
  AND U3775 ( .A(n26551), .B(n2854), .Z(n2855) );
  NANDN U3776 ( .A(n2855), .B(n26552), .Z(n2856) );
  NANDN U3777 ( .A(n26553), .B(n2856), .Z(n2857) );
  NAND U3778 ( .A(n26554), .B(n2857), .Z(n2858) );
  NAND U3779 ( .A(n26555), .B(n2858), .Z(n26556) );
  NANDN U3780 ( .A(n13736), .B(n4572), .Z(n2859) );
  AND U3781 ( .A(n17063), .B(n2859), .Z(n26354) );
  NAND U3782 ( .A(n26587), .B(n26588), .Z(n2860) );
  NAND U3783 ( .A(n26589), .B(n2860), .Z(n2861) );
  NAND U3784 ( .A(n26590), .B(n2861), .Z(n2862) );
  NAND U3785 ( .A(n26591), .B(n2862), .Z(n2863) );
  NANDN U3786 ( .A(n26592), .B(n2863), .Z(n2864) );
  ANDN U3787 ( .B(n2864), .A(n26593), .Z(n2865) );
  OR U3788 ( .A(n24408), .B(n2865), .Z(n2866) );
  NAND U3789 ( .A(n26594), .B(n2866), .Z(n2867) );
  NAND U3790 ( .A(n26595), .B(n2867), .Z(n2868) );
  NANDN U3791 ( .A(n26596), .B(n2868), .Z(n2869) );
  NAND U3792 ( .A(n26597), .B(n2869), .Z(n2870) );
  AND U3793 ( .A(n26598), .B(n2870), .Z(n2871) );
  NANDN U3794 ( .A(n26601), .B(n26600), .Z(n2872) );
  ANDN U3795 ( .B(n2872), .A(n26602), .Z(n2873) );
  NANDN U3796 ( .A(n2871), .B(n26599), .Z(n2874) );
  NAND U3797 ( .A(n2873), .B(n2874), .Z(n2875) );
  NAND U3798 ( .A(n26603), .B(n2875), .Z(n26604) );
  NANDN U3799 ( .A(n26664), .B(n26663), .Z(n2876) );
  NAND U3800 ( .A(n26665), .B(n2876), .Z(n2877) );
  NANDN U3801 ( .A(n26666), .B(n2877), .Z(n2878) );
  NAND U3802 ( .A(n26667), .B(n2878), .Z(n2879) );
  NAND U3803 ( .A(n26668), .B(n2879), .Z(n2880) );
  ANDN U3804 ( .B(n2880), .A(n24406), .Z(n2881) );
  NANDN U3805 ( .A(n2881), .B(n24405), .Z(n2882) );
  NAND U3806 ( .A(n26669), .B(n2882), .Z(n2883) );
  NANDN U3807 ( .A(n26670), .B(n2883), .Z(n2884) );
  NAND U3808 ( .A(n26671), .B(n2884), .Z(n2885) );
  NANDN U3809 ( .A(n26672), .B(n2885), .Z(n2886) );
  AND U3810 ( .A(n26673), .B(n2886), .Z(n2887) );
  OR U3811 ( .A(n2887), .B(n26674), .Z(n2888) );
  AND U3812 ( .A(n26675), .B(n2888), .Z(n2889) );
  OR U3813 ( .A(n26676), .B(n2889), .Z(n2890) );
  NAND U3814 ( .A(n26677), .B(n2890), .Z(n2891) );
  NANDN U3815 ( .A(n26678), .B(n2891), .Z(n26680) );
  NAND U3816 ( .A(n26715), .B(n26716), .Z(n2892) );
  NANDN U3817 ( .A(n26717), .B(n2892), .Z(n2893) );
  NAND U3818 ( .A(n26718), .B(n2893), .Z(n2894) );
  NAND U3819 ( .A(n26719), .B(n2894), .Z(n2895) );
  NAND U3820 ( .A(n24403), .B(n2895), .Z(n2896) );
  AND U3821 ( .A(n26720), .B(n2896), .Z(n2897) );
  NANDN U3822 ( .A(n2897), .B(n26721), .Z(n2898) );
  NAND U3823 ( .A(n24402), .B(n2898), .Z(n2899) );
  NAND U3824 ( .A(n26722), .B(n2899), .Z(n2900) );
  NAND U3825 ( .A(n26723), .B(n2900), .Z(n2901) );
  NANDN U3826 ( .A(n26724), .B(n2901), .Z(n2902) );
  AND U3827 ( .A(n26725), .B(n2902), .Z(n2903) );
  OR U3828 ( .A(n26726), .B(n2903), .Z(n2904) );
  NANDN U3829 ( .A(n24401), .B(n2904), .Z(n2905) );
  NAND U3830 ( .A(n26727), .B(n2905), .Z(n2906) );
  NAND U3831 ( .A(n26728), .B(n2906), .Z(n26729) );
  NOR U3832 ( .A(n17798), .B(n17799), .Z(n26770) );
  NANDN U3833 ( .A(y[1296]), .B(x[1296]), .Z(n2907) );
  NAND U3834 ( .A(n13630), .B(n2907), .Z(n2908) );
  NAND U3835 ( .A(n7256), .B(n2908), .Z(n2909) );
  AND U3836 ( .A(n13631), .B(n2909), .Z(n24422) );
  ANDN U3837 ( .B(n13491), .A(n13490), .Z(n26782) );
  NAND U3838 ( .A(n26809), .B(n24390), .Z(n2910) );
  ANDN U3839 ( .B(n2910), .A(n26810), .Z(n2911) );
  NANDN U3840 ( .A(n2911), .B(n26811), .Z(n2912) );
  NAND U3841 ( .A(n26812), .B(n2912), .Z(n2913) );
  NAND U3842 ( .A(n26813), .B(n2913), .Z(n2914) );
  ANDN U3843 ( .B(n24389), .A(n24388), .Z(n2915) );
  NAND U3844 ( .A(n2914), .B(n2915), .Z(n2916) );
  NANDN U3845 ( .A(n26814), .B(n2916), .Z(n2917) );
  NAND U3846 ( .A(n26815), .B(n2917), .Z(n2918) );
  NAND U3847 ( .A(n26816), .B(n2918), .Z(n2919) );
  AND U3848 ( .A(n24387), .B(n2919), .Z(n2920) );
  NANDN U3849 ( .A(n2920), .B(n26817), .Z(n2921) );
  ANDN U3850 ( .B(n2921), .A(n26818), .Z(n2922) );
  NANDN U3851 ( .A(n2922), .B(n26819), .Z(n2923) );
  NAND U3852 ( .A(n26820), .B(n2923), .Z(n2924) );
  NAND U3853 ( .A(n26821), .B(n2924), .Z(n26822) );
  NOR U3854 ( .A(n13444), .B(n13445), .Z(n26862) );
  ANDN U3855 ( .B(n13436), .A(n13435), .Z(n26880) );
  NAND U3856 ( .A(n26901), .B(n26900), .Z(n2925) );
  NANDN U3857 ( .A(n26902), .B(n2925), .Z(n2926) );
  NAND U3858 ( .A(n26903), .B(n2926), .Z(n2927) );
  NANDN U3859 ( .A(n24373), .B(n2927), .Z(n2928) );
  NAND U3860 ( .A(n24372), .B(n2928), .Z(n2929) );
  ANDN U3861 ( .B(n2929), .A(n24371), .Z(n2930) );
  NANDN U3862 ( .A(n2930), .B(n24370), .Z(n2931) );
  NAND U3863 ( .A(n26904), .B(n2931), .Z(n2932) );
  NAND U3864 ( .A(n26905), .B(n2932), .Z(n2933) );
  NANDN U3865 ( .A(n26906), .B(n2933), .Z(n2934) );
  NANDN U3866 ( .A(n26907), .B(n2934), .Z(n2935) );
  ANDN U3867 ( .B(n2935), .A(n26908), .Z(n2936) );
  NANDN U3868 ( .A(n2936), .B(n26909), .Z(n2937) );
  ANDN U3869 ( .B(n2937), .A(n26910), .Z(n26912) );
  NAND U3870 ( .A(n26944), .B(n24366), .Z(n2938) );
  NAND U3871 ( .A(n26945), .B(n2938), .Z(n2939) );
  AND U3872 ( .A(n26946), .B(n2939), .Z(n2940) );
  OR U3873 ( .A(n26947), .B(n2940), .Z(n2941) );
  NAND U3874 ( .A(n26948), .B(n2941), .Z(n2942) );
  NANDN U3875 ( .A(n26949), .B(n2942), .Z(n2943) );
  NAND U3876 ( .A(n26950), .B(n2943), .Z(n2944) );
  NANDN U3877 ( .A(n26951), .B(n2944), .Z(n2945) );
  AND U3878 ( .A(n26952), .B(n2945), .Z(n2946) );
  NANDN U3879 ( .A(n2946), .B(n26953), .Z(n2947) );
  NANDN U3880 ( .A(n24365), .B(n2947), .Z(n2948) );
  NANDN U3881 ( .A(n26954), .B(n2948), .Z(n2949) );
  NAND U3882 ( .A(n26955), .B(n2949), .Z(n2950) );
  NANDN U3883 ( .A(n26956), .B(n2950), .Z(n2951) );
  AND U3884 ( .A(n26957), .B(n2951), .Z(n26959) );
  NAND U3885 ( .A(n17787), .B(n4412), .Z(n2952) );
  ANDN U3886 ( .B(n2952), .A(n17791), .Z(n26762) );
  NANDN U3887 ( .A(y[1520]), .B(x[1520]), .Z(n2953) );
  NANDN U3888 ( .A(y[1521]), .B(x[1521]), .Z(n2954) );
  AND U3889 ( .A(n2953), .B(n2954), .Z(n2955) );
  NANDN U3890 ( .A(y[1523]), .B(x[1523]), .Z(n2956) );
  NANDN U3891 ( .A(y[1522]), .B(x[1522]), .Z(n2957) );
  AND U3892 ( .A(n2956), .B(n2957), .Z(n2958) );
  NANDN U3893 ( .A(n2955), .B(n4395), .Z(n2959) );
  AND U3894 ( .A(n2958), .B(n2959), .Z(n13494) );
  NANDN U3895 ( .A(n26990), .B(n26989), .Z(n2960) );
  NAND U3896 ( .A(n26991), .B(n2960), .Z(n2961) );
  ANDN U3897 ( .B(n2961), .A(n26992), .Z(n2962) );
  OR U3898 ( .A(n26993), .B(n2962), .Z(n2963) );
  NAND U3899 ( .A(n26994), .B(n2963), .Z(n2964) );
  NANDN U3900 ( .A(n24359), .B(n2964), .Z(n2965) );
  NAND U3901 ( .A(n26995), .B(n2965), .Z(n2966) );
  NAND U3902 ( .A(n26996), .B(n2966), .Z(n2967) );
  AND U3903 ( .A(n26997), .B(n2967), .Z(n2968) );
  NANDN U3904 ( .A(n2968), .B(n26998), .Z(n2969) );
  NAND U3905 ( .A(n26999), .B(n2969), .Z(n2970) );
  NAND U3906 ( .A(n27000), .B(n2970), .Z(n2971) );
  NANDN U3907 ( .A(n27001), .B(n2971), .Z(n2972) );
  NAND U3908 ( .A(n27002), .B(n2972), .Z(n2973) );
  ANDN U3909 ( .B(n2973), .A(n27003), .Z(n2974) );
  NANDN U3910 ( .A(n2974), .B(n27004), .Z(n2975) );
  NANDN U3911 ( .A(n27005), .B(n2975), .Z(n2976) );
  NAND U3912 ( .A(n27006), .B(n2976), .Z(n27007) );
  NAND U3913 ( .A(n27036), .B(n27035), .Z(n2977) );
  NANDN U3914 ( .A(n27038), .B(n2977), .Z(n2978) );
  NAND U3915 ( .A(n27039), .B(n2978), .Z(n2979) );
  NAND U3916 ( .A(n24353), .B(n2979), .Z(n2980) );
  NANDN U3917 ( .A(n27040), .B(n2980), .Z(n2981) );
  AND U3918 ( .A(n27041), .B(n2981), .Z(n2982) );
  OR U3919 ( .A(n2982), .B(n27042), .Z(n2983) );
  NAND U3920 ( .A(n27043), .B(n2983), .Z(n2984) );
  NANDN U3921 ( .A(n27044), .B(n2984), .Z(n2985) );
  NAND U3922 ( .A(n27045), .B(n2985), .Z(n2986) );
  NANDN U3923 ( .A(n27046), .B(n2986), .Z(n2987) );
  AND U3924 ( .A(n27047), .B(n2987), .Z(n2988) );
  OR U3925 ( .A(n27048), .B(n2988), .Z(n2989) );
  NAND U3926 ( .A(n27049), .B(n2989), .Z(n2990) );
  NANDN U3927 ( .A(n27050), .B(n2990), .Z(n2991) );
  NAND U3928 ( .A(n27051), .B(n2991), .Z(n2992) );
  NANDN U3929 ( .A(n27052), .B(n2992), .Z(n2993) );
  ANDN U3930 ( .B(n2993), .A(n27053), .Z(n27056) );
  NANDN U3931 ( .A(n17929), .B(n7686), .Z(n2994) );
  AND U3932 ( .A(n17933), .B(n2994), .Z(n26837) );
  OR U3933 ( .A(n27083), .B(n27082), .Z(n2995) );
  NAND U3934 ( .A(n27085), .B(n2995), .Z(n2996) );
  NAND U3935 ( .A(n27086), .B(n2996), .Z(n2997) );
  NAND U3936 ( .A(n27087), .B(n2997), .Z(n2998) );
  NAND U3937 ( .A(n24345), .B(n2998), .Z(n2999) );
  ANDN U3938 ( .B(n2999), .A(n27088), .Z(n3000) );
  NANDN U3939 ( .A(n3000), .B(n27089), .Z(n3001) );
  NANDN U3940 ( .A(n27090), .B(n3001), .Z(n3002) );
  NAND U3941 ( .A(n27091), .B(n3002), .Z(n3003) );
  NAND U3942 ( .A(n27092), .B(n3003), .Z(n3004) );
  NANDN U3943 ( .A(n27093), .B(n3004), .Z(n3005) );
  ANDN U3944 ( .B(n3005), .A(n27094), .Z(n3006) );
  OR U3945 ( .A(n27095), .B(n3006), .Z(n3007) );
  NAND U3946 ( .A(n27096), .B(n3007), .Z(n3008) );
  NAND U3947 ( .A(n27097), .B(n3008), .Z(n3009) );
  NAND U3948 ( .A(n27098), .B(n3009), .Z(n27099) );
  NANDN U3949 ( .A(n13244), .B(n13245), .Z(n27113) );
  OR U3950 ( .A(n27168), .B(n27169), .Z(n3010) );
  NANDN U3951 ( .A(n24339), .B(n3010), .Z(n3011) );
  NAND U3952 ( .A(n27170), .B(n3011), .Z(n3012) );
  NAND U3953 ( .A(n27171), .B(n3012), .Z(n3013) );
  NANDN U3954 ( .A(n27172), .B(n3013), .Z(n3014) );
  AND U3955 ( .A(n27173), .B(n3014), .Z(n3015) );
  OR U3956 ( .A(n3015), .B(n27174), .Z(n3016) );
  NAND U3957 ( .A(n27175), .B(n3016), .Z(n3017) );
  ANDN U3958 ( .B(n3017), .A(n27176), .Z(n3018) );
  NANDN U3959 ( .A(n3018), .B(n27177), .Z(n3019) );
  NANDN U3960 ( .A(n27178), .B(n3019), .Z(n3020) );
  NAND U3961 ( .A(n27179), .B(n3020), .Z(n3021) );
  NANDN U3962 ( .A(n27180), .B(n3021), .Z(n3022) );
  NAND U3963 ( .A(n27181), .B(n3022), .Z(n3023) );
  AND U3964 ( .A(n27182), .B(n3023), .Z(n3024) );
  OR U3965 ( .A(n27183), .B(n3024), .Z(n3025) );
  NAND U3966 ( .A(n27184), .B(n3025), .Z(n3026) );
  NANDN U3967 ( .A(n27185), .B(n3026), .Z(n3027) );
  AND U3968 ( .A(n27186), .B(n3027), .Z(n27188) );
  ANDN U3969 ( .B(n13160), .A(n13159), .Z(n27213) );
  NAND U3970 ( .A(n27234), .B(n27233), .Z(n3028) );
  NANDN U3971 ( .A(n27236), .B(n3028), .Z(n3029) );
  NAND U3972 ( .A(n27237), .B(n3029), .Z(n3030) );
  NAND U3973 ( .A(n24331), .B(n3030), .Z(n3031) );
  NANDN U3974 ( .A(n27238), .B(n3031), .Z(n3032) );
  ANDN U3975 ( .B(n3032), .A(n27239), .Z(n3033) );
  OR U3976 ( .A(n24330), .B(n3033), .Z(n3034) );
  NAND U3977 ( .A(n27240), .B(n3034), .Z(n3035) );
  NAND U3978 ( .A(n27241), .B(n3035), .Z(n3036) );
  NANDN U3979 ( .A(n27242), .B(n3036), .Z(n3037) );
  NAND U3980 ( .A(n27243), .B(n3037), .Z(n3038) );
  ANDN U3981 ( .B(n3038), .A(n27244), .Z(n3039) );
  NANDN U3982 ( .A(n3039), .B(n27245), .Z(n3040) );
  NAND U3983 ( .A(n27246), .B(n3040), .Z(n3041) );
  NAND U3984 ( .A(n27247), .B(n3041), .Z(n3042) );
  NAND U3985 ( .A(n27248), .B(n3042), .Z(n27249) );
  NAND U3986 ( .A(n27278), .B(n27279), .Z(n3043) );
  NAND U3987 ( .A(n24325), .B(n3043), .Z(n3044) );
  NANDN U3988 ( .A(n24324), .B(n3044), .Z(n3045) );
  NAND U3989 ( .A(n24323), .B(n3045), .Z(n3046) );
  NAND U3990 ( .A(n27280), .B(n3046), .Z(n3047) );
  ANDN U3991 ( .B(n3047), .A(n27281), .Z(n3048) );
  NANDN U3992 ( .A(n3048), .B(n27282), .Z(n3049) );
  NANDN U3993 ( .A(n27283), .B(n3049), .Z(n3050) );
  NAND U3994 ( .A(n27284), .B(n3050), .Z(n3051) );
  NANDN U3995 ( .A(n27285), .B(n3051), .Z(n3052) );
  NANDN U3996 ( .A(n27286), .B(n3052), .Z(n3053) );
  AND U3997 ( .A(n27287), .B(n3053), .Z(n3054) );
  NANDN U3998 ( .A(n3054), .B(n27288), .Z(n3055) );
  NAND U3999 ( .A(n27289), .B(n3055), .Z(n3056) );
  NAND U4000 ( .A(n27290), .B(n3056), .Z(n3057) );
  NAND U4001 ( .A(n27291), .B(n3057), .Z(n27292) );
  NANDN U4002 ( .A(n27328), .B(n27327), .Z(n3058) );
  NAND U4003 ( .A(n27329), .B(n3058), .Z(n3059) );
  NANDN U4004 ( .A(n27330), .B(n3059), .Z(n3060) );
  NANDN U4005 ( .A(n27331), .B(n3060), .Z(n3061) );
  NAND U4006 ( .A(n27332), .B(n3061), .Z(n3062) );
  AND U4007 ( .A(n27333), .B(n3062), .Z(n3063) );
  NANDN U4008 ( .A(n3063), .B(n24316), .Z(n3064) );
  NANDN U4009 ( .A(n24315), .B(n3064), .Z(n3065) );
  NAND U4010 ( .A(n27334), .B(n3065), .Z(n3066) );
  NANDN U4011 ( .A(n27335), .B(n3066), .Z(n3067) );
  NAND U4012 ( .A(n27336), .B(n3067), .Z(n3068) );
  AND U4013 ( .A(n27337), .B(n3068), .Z(n3069) );
  OR U4014 ( .A(n3069), .B(n27338), .Z(n3070) );
  AND U4015 ( .A(n27339), .B(n3070), .Z(n3071) );
  OR U4016 ( .A(n27340), .B(n3071), .Z(n3072) );
  NAND U4017 ( .A(n27341), .B(n3072), .Z(n3073) );
  NANDN U4018 ( .A(n27342), .B(n3073), .Z(n27343) );
  NANDN U4019 ( .A(n27374), .B(n27373), .Z(n3074) );
  NAND U4020 ( .A(n27375), .B(n3074), .Z(n3075) );
  AND U4021 ( .A(n27376), .B(n3075), .Z(n3076) );
  OR U4022 ( .A(n27377), .B(n3076), .Z(n3077) );
  NAND U4023 ( .A(n27378), .B(n3077), .Z(n3078) );
  NANDN U4024 ( .A(n27379), .B(n3078), .Z(n3079) );
  NAND U4025 ( .A(n27380), .B(n3079), .Z(n3080) );
  NANDN U4026 ( .A(n27381), .B(n3080), .Z(n3081) );
  AND U4027 ( .A(n27382), .B(n3081), .Z(n3082) );
  NANDN U4028 ( .A(n3082), .B(n27383), .Z(n3083) );
  NAND U4029 ( .A(n27384), .B(n3083), .Z(n3084) );
  NAND U4030 ( .A(n27385), .B(n3084), .Z(n3085) );
  NANDN U4031 ( .A(n27386), .B(n3085), .Z(n27387) );
  NANDN U4032 ( .A(n27419), .B(n27418), .Z(n3086) );
  NAND U4033 ( .A(n27420), .B(n3086), .Z(n3087) );
  NAND U4034 ( .A(n27421), .B(n3087), .Z(n3088) );
  NANDN U4035 ( .A(n24303), .B(n3088), .Z(n3089) );
  NAND U4036 ( .A(n24302), .B(n3089), .Z(n3090) );
  ANDN U4037 ( .B(n3090), .A(n27422), .Z(n3091) );
  NANDN U4038 ( .A(n3091), .B(n27423), .Z(n3092) );
  NANDN U4039 ( .A(n24301), .B(n3092), .Z(n3093) );
  NAND U4040 ( .A(n24300), .B(n3093), .Z(n3094) );
  NAND U4041 ( .A(n27424), .B(n3094), .Z(n3095) );
  AND U4042 ( .A(n27426), .B(n3095), .Z(n3096) );
  NANDN U4043 ( .A(n27425), .B(n3096), .Z(n27427) );
  NAND U4044 ( .A(n27452), .B(n27453), .Z(n3097) );
  NANDN U4045 ( .A(n27455), .B(n3097), .Z(n3098) );
  NANDN U4046 ( .A(n27456), .B(n3098), .Z(n3099) );
  NAND U4047 ( .A(n27457), .B(n3099), .Z(n3100) );
  NANDN U4048 ( .A(n27458), .B(n3100), .Z(n3101) );
  AND U4049 ( .A(n27459), .B(n3101), .Z(n3102) );
  OR U4050 ( .A(n27460), .B(n3102), .Z(n3103) );
  NAND U4051 ( .A(n27461), .B(n3103), .Z(n3104) );
  NANDN U4052 ( .A(n24291), .B(n3104), .Z(n3105) );
  NAND U4053 ( .A(n27462), .B(n3105), .Z(n3106) );
  NAND U4054 ( .A(n27463), .B(n3106), .Z(n3107) );
  AND U4055 ( .A(n27464), .B(n3107), .Z(n3108) );
  OR U4056 ( .A(n27465), .B(n3108), .Z(n3109) );
  ANDN U4057 ( .B(n3109), .A(n27466), .Z(n3110) );
  OR U4058 ( .A(n27467), .B(n3110), .Z(n3111) );
  NAND U4059 ( .A(n27468), .B(n3111), .Z(n3112) );
  NANDN U4060 ( .A(n24290), .B(n3112), .Z(n27469) );
  AND U4061 ( .A(n8209), .B(n27192), .Z(n3113) );
  NAND U4062 ( .A(n13183), .B(n3113), .Z(n3114) );
  ANDN U4063 ( .B(n3114), .A(n13180), .Z(n3115) );
  AND U4064 ( .A(n13182), .B(n13179), .Z(n3116) );
  NANDN U4065 ( .A(n18511), .B(n3115), .Z(n3117) );
  NAND U4066 ( .A(n3116), .B(n3117), .Z(n3118) );
  AND U4067 ( .A(n13181), .B(n13177), .Z(n3119) );
  NAND U4068 ( .A(n3118), .B(n3119), .Z(n3120) );
  NAND U4069 ( .A(n27198), .B(n3120), .Z(n3121) );
  AND U4070 ( .A(n13176), .B(n27199), .Z(n3122) );
  OR U4071 ( .A(n3121), .B(n13178), .Z(n3123) );
  AND U4072 ( .A(n3122), .B(n3123), .Z(n3124) );
  NANDN U4073 ( .A(n3124), .B(n27200), .Z(n3125) );
  NAND U4074 ( .A(n27201), .B(n3125), .Z(n3126) );
  NAND U4075 ( .A(n27202), .B(n3126), .Z(n3127) );
  AND U4076 ( .A(n13172), .B(n27204), .Z(n3128) );
  NANDN U4077 ( .A(n27203), .B(n3127), .Z(n3129) );
  NAND U4078 ( .A(n3128), .B(n3129), .Z(n3130) );
  ANDN U4079 ( .B(n3130), .A(n13169), .Z(n8210) );
  NANDN U4080 ( .A(n24287), .B(n24288), .Z(n3131) );
  NAND U4081 ( .A(n27503), .B(n3131), .Z(n3132) );
  AND U4082 ( .A(n27504), .B(n3132), .Z(n3133) );
  OR U4083 ( .A(n3133), .B(n27505), .Z(n3134) );
  NAND U4084 ( .A(n27506), .B(n3134), .Z(n3135) );
  AND U4085 ( .A(n27507), .B(n3135), .Z(n3136) );
  NANDN U4086 ( .A(n3136), .B(n27508), .Z(n3137) );
  NANDN U4087 ( .A(n27509), .B(n3137), .Z(n3138) );
  NAND U4088 ( .A(n27510), .B(n3138), .Z(n3139) );
  NAND U4089 ( .A(n27511), .B(n3139), .Z(n3140) );
  NAND U4090 ( .A(n27512), .B(n3140), .Z(n3141) );
  ANDN U4091 ( .B(n3141), .A(n27513), .Z(n3142) );
  NANDN U4092 ( .A(n3142), .B(n27514), .Z(n3143) );
  ANDN U4093 ( .B(n3143), .A(n27515), .Z(n3144) );
  NANDN U4094 ( .A(n3144), .B(n27516), .Z(n3145) );
  NANDN U4095 ( .A(n27517), .B(n3145), .Z(n3146) );
  NAND U4096 ( .A(n27518), .B(n3146), .Z(n27519) );
  NANDN U4097 ( .A(y[1945]), .B(x[1945]), .Z(n3147) );
  ANDN U4098 ( .B(n3147), .A(n8304), .Z(n13110) );
  OR U4099 ( .A(n27542), .B(n27541), .Z(n3148) );
  NAND U4100 ( .A(n27543), .B(n3148), .Z(n3149) );
  ANDN U4101 ( .B(n3149), .A(n27544), .Z(n3150) );
  OR U4102 ( .A(n27545), .B(n3150), .Z(n3151) );
  NAND U4103 ( .A(n27546), .B(n3151), .Z(n3152) );
  NANDN U4104 ( .A(n27547), .B(n3152), .Z(n3153) );
  NAND U4105 ( .A(n27548), .B(n3153), .Z(n3154) );
  NANDN U4106 ( .A(n24276), .B(n3154), .Z(n3155) );
  AND U4107 ( .A(n27549), .B(n3155), .Z(n3156) );
  NANDN U4108 ( .A(n3156), .B(n27550), .Z(n3157) );
  NAND U4109 ( .A(n24275), .B(n3157), .Z(n3158) );
  NANDN U4110 ( .A(n27551), .B(n3158), .Z(n3159) );
  NAND U4111 ( .A(n27552), .B(n3159), .Z(n27553) );
  ANDN U4112 ( .B(n12852), .A(n12851), .Z(n27581) );
  NAND U4113 ( .A(n27599), .B(n27600), .Z(n3160) );
  NANDN U4114 ( .A(n27601), .B(n3160), .Z(n3161) );
  NAND U4115 ( .A(n27602), .B(n3161), .Z(n3162) );
  NAND U4116 ( .A(n27603), .B(n3162), .Z(n3163) );
  NAND U4117 ( .A(n27604), .B(n3163), .Z(n3164) );
  ANDN U4118 ( .B(n3164), .A(n24268), .Z(n3165) );
  OR U4119 ( .A(n3165), .B(n27605), .Z(n3166) );
  NAND U4120 ( .A(n27606), .B(n3166), .Z(n3167) );
  NAND U4121 ( .A(n27607), .B(n3167), .Z(n3168) );
  NAND U4122 ( .A(n27608), .B(n3168), .Z(n3169) );
  NANDN U4123 ( .A(n27609), .B(n3169), .Z(n3170) );
  AND U4124 ( .A(n27610), .B(n3170), .Z(n3171) );
  NANDN U4125 ( .A(n3171), .B(n27611), .Z(n3172) );
  AND U4126 ( .A(n27612), .B(n3172), .Z(n3173) );
  OR U4127 ( .A(n27613), .B(n3173), .Z(n3174) );
  NANDN U4128 ( .A(n27614), .B(n3174), .Z(n3175) );
  NAND U4129 ( .A(n27615), .B(n3175), .Z(n27616) );
  OR U4130 ( .A(n27648), .B(n27649), .Z(n3176) );
  NAND U4131 ( .A(n27650), .B(n3176), .Z(n3177) );
  AND U4132 ( .A(n24262), .B(n3177), .Z(n3178) );
  OR U4133 ( .A(n24261), .B(n3178), .Z(n3179) );
  NAND U4134 ( .A(n24260), .B(n3179), .Z(n3180) );
  NAND U4135 ( .A(n27651), .B(n3180), .Z(n3181) );
  NAND U4136 ( .A(n27652), .B(n3181), .Z(n3182) );
  NANDN U4137 ( .A(n24259), .B(n3182), .Z(n3183) );
  AND U4138 ( .A(n24258), .B(n3183), .Z(n3184) );
  NANDN U4139 ( .A(n3184), .B(n27653), .Z(n3185) );
  AND U4140 ( .A(n27654), .B(n3185), .Z(n3186) );
  OR U4141 ( .A(n27655), .B(n3186), .Z(n3187) );
  NAND U4142 ( .A(n27656), .B(n3187), .Z(n3188) );
  NANDN U4143 ( .A(n27657), .B(n3188), .Z(n27658) );
  NAND U4144 ( .A(n27717), .B(n27718), .Z(n3189) );
  NAND U4145 ( .A(n27720), .B(n3189), .Z(n3190) );
  NAND U4146 ( .A(n27721), .B(n3190), .Z(n3191) );
  NANDN U4147 ( .A(n27722), .B(n3191), .Z(n3192) );
  NAND U4148 ( .A(n27723), .B(n3192), .Z(n3193) );
  AND U4149 ( .A(n27724), .B(n3193), .Z(n3194) );
  NANDN U4150 ( .A(n3194), .B(n27725), .Z(n3195) );
  NANDN U4151 ( .A(n27726), .B(n3195), .Z(n3196) );
  NAND U4152 ( .A(n27727), .B(n3196), .Z(n3197) );
  NAND U4153 ( .A(n27728), .B(n3197), .Z(n3198) );
  NAND U4154 ( .A(n27729), .B(n3198), .Z(n3199) );
  ANDN U4155 ( .B(n3199), .A(n27730), .Z(n3200) );
  NANDN U4156 ( .A(n3200), .B(n27731), .Z(n3201) );
  NAND U4157 ( .A(n27732), .B(n3201), .Z(n3202) );
  NANDN U4158 ( .A(n27733), .B(n3202), .Z(n3203) );
  AND U4159 ( .A(n27734), .B(n3203), .Z(n27735) );
  NAND U4160 ( .A(n27777), .B(n27776), .Z(n3204) );
  NANDN U4161 ( .A(n27779), .B(n3204), .Z(n3205) );
  NANDN U4162 ( .A(n27780), .B(n3205), .Z(n3206) );
  NAND U4163 ( .A(n27781), .B(n3206), .Z(n3207) );
  NAND U4164 ( .A(n27782), .B(n3207), .Z(n3208) );
  ANDN U4165 ( .B(n3208), .A(n27783), .Z(n3209) );
  NAND U4166 ( .A(n27784), .B(n3209), .Z(n3210) );
  NAND U4167 ( .A(n27785), .B(n3210), .Z(n3211) );
  NANDN U4168 ( .A(n27786), .B(n3211), .Z(n3212) );
  NAND U4169 ( .A(n27788), .B(n27787), .Z(n3213) );
  NANDN U4170 ( .A(n3212), .B(n3213), .Z(n3214) );
  AND U4171 ( .A(n27789), .B(n3214), .Z(n3215) );
  OR U4172 ( .A(n27790), .B(n3215), .Z(n3216) );
  NAND U4173 ( .A(n27791), .B(n3216), .Z(n3217) );
  NANDN U4174 ( .A(n27792), .B(n3217), .Z(n3218) );
  NAND U4175 ( .A(n27793), .B(n3218), .Z(n3219) );
  ANDN U4176 ( .B(n3219), .A(n27795), .Z(n3220) );
  NANDN U4177 ( .A(n27794), .B(n3220), .Z(n27796) );
  ANDN U4178 ( .B(n8633), .A(n12953), .Z(n3221) );
  NAND U4179 ( .A(n27475), .B(n3221), .Z(n3222) );
  AND U4180 ( .A(n27476), .B(n3222), .Z(n3223) );
  OR U4181 ( .A(n12951), .B(n3223), .Z(n3224) );
  ANDN U4182 ( .B(n3224), .A(n27478), .Z(n3225) );
  ANDN U4183 ( .B(n12952), .A(n3225), .Z(n3226) );
  NAND U4184 ( .A(n27479), .B(n3226), .Z(n3227) );
  NAND U4185 ( .A(n27480), .B(n3227), .Z(n3228) );
  NANDN U4186 ( .A(n27481), .B(n3228), .Z(n3229) );
  NAND U4187 ( .A(n27482), .B(n3229), .Z(n3230) );
  AND U4188 ( .A(n12949), .B(n3230), .Z(n3231) );
  ANDN U4189 ( .B(n12948), .A(n12947), .Z(n3232) );
  NANDN U4190 ( .A(n3231), .B(n27485), .Z(n3233) );
  AND U4191 ( .A(n3232), .B(n3233), .Z(n3234) );
  OR U4192 ( .A(n19017), .B(n3234), .Z(n3235) );
  AND U4193 ( .A(n27486), .B(n3235), .Z(n3236) );
  AND U4194 ( .A(n12944), .B(n12946), .Z(n3237) );
  NANDN U4195 ( .A(n3236), .B(n12945), .Z(n3238) );
  AND U4196 ( .A(n3237), .B(n3238), .Z(n8638) );
  NAND U4197 ( .A(n27824), .B(y[2450]), .Z(n3239) );
  NANDN U4198 ( .A(x[2450]), .B(n27823), .Z(n3240) );
  NAND U4199 ( .A(n3239), .B(n3240), .Z(n3241) );
  NAND U4200 ( .A(n27825), .B(n3241), .Z(n3242) );
  NAND U4201 ( .A(n27826), .B(n3242), .Z(n3243) );
  ANDN U4202 ( .B(n3243), .A(n27827), .Z(n3244) );
  NANDN U4203 ( .A(n3244), .B(n27828), .Z(n3245) );
  NANDN U4204 ( .A(n27829), .B(n3245), .Z(n3246) );
  NAND U4205 ( .A(n27830), .B(n3246), .Z(n3247) );
  NAND U4206 ( .A(n27831), .B(n3247), .Z(n3248) );
  NAND U4207 ( .A(n27832), .B(n3248), .Z(n3249) );
  AND U4208 ( .A(n27833), .B(n3249), .Z(n3250) );
  OR U4209 ( .A(n27834), .B(n3250), .Z(n3251) );
  AND U4210 ( .A(n27835), .B(n3251), .Z(n3252) );
  ANDN U4211 ( .B(n27836), .A(n3252), .Z(n3253) );
  NANDN U4212 ( .A(n24240), .B(n24239), .Z(n3254) );
  NAND U4213 ( .A(n3253), .B(n3254), .Z(n3255) );
  NANDN U4214 ( .A(n27837), .B(n3255), .Z(n27838) );
  NAND U4215 ( .A(n27878), .B(n24237), .Z(n3256) );
  NAND U4216 ( .A(n27879), .B(n3256), .Z(n3257) );
  AND U4217 ( .A(n27880), .B(n3257), .Z(n3258) );
  NOR U4218 ( .A(n27882), .B(n3258), .Z(n3259) );
  NAND U4219 ( .A(n27881), .B(n3259), .Z(n3260) );
  AND U4220 ( .A(n27883), .B(n3260), .Z(n3261) );
  OR U4221 ( .A(n3261), .B(n27884), .Z(n3262) );
  NAND U4222 ( .A(n27885), .B(n3262), .Z(n3263) );
  ANDN U4223 ( .B(n3263), .A(n27886), .Z(n3264) );
  NANDN U4224 ( .A(n3264), .B(n27887), .Z(n3265) );
  NAND U4225 ( .A(n27888), .B(n3265), .Z(n3266) );
  NANDN U4226 ( .A(n27889), .B(n3266), .Z(n3267) );
  NAND U4227 ( .A(n27890), .B(n3267), .Z(n3268) );
  NANDN U4228 ( .A(n27891), .B(n3268), .Z(n3269) );
  AND U4229 ( .A(n27892), .B(n3269), .Z(n3270) );
  OR U4230 ( .A(n27893), .B(n3270), .Z(n3271) );
  NAND U4231 ( .A(n27894), .B(n3271), .Z(n3272) );
  NANDN U4232 ( .A(n27895), .B(n3272), .Z(n27897) );
  NOR U4233 ( .A(n12874), .B(n8756), .Z(n3273) );
  NAND U4234 ( .A(n27562), .B(n3273), .Z(n3274) );
  AND U4235 ( .A(n27563), .B(n3274), .Z(n3275) );
  OR U4236 ( .A(n8757), .B(n19171), .Z(n3276) );
  NAND U4237 ( .A(n3275), .B(n3276), .Z(n3277) );
  NANDN U4238 ( .A(n12873), .B(n3277), .Z(n3278) );
  NANDN U4239 ( .A(y[2218]), .B(n3278), .Z(n3279) );
  ANDN U4240 ( .B(n3279), .A(n19180), .Z(n3280) );
  XNOR U4241 ( .A(y[2218]), .B(n3278), .Z(n3281) );
  NAND U4242 ( .A(n3281), .B(x[2218]), .Z(n3282) );
  NAND U4243 ( .A(n3280), .B(n3282), .Z(n3283) );
  AND U4244 ( .A(n19177), .B(n27566), .Z(n3284) );
  NAND U4245 ( .A(n3283), .B(n3284), .Z(n3285) );
  NAND U4246 ( .A(n19181), .B(n3285), .Z(n3286) );
  NANDN U4247 ( .A(n3286), .B(n27567), .Z(n3287) );
  AND U4248 ( .A(n27568), .B(n3287), .Z(n3288) );
  OR U4249 ( .A(n27569), .B(n3288), .Z(n3289) );
  NAND U4250 ( .A(n12871), .B(n3289), .Z(n3290) );
  NANDN U4251 ( .A(n12869), .B(n3290), .Z(n8758) );
  NAND U4252 ( .A(n27952), .B(n27953), .Z(n3291) );
  NAND U4253 ( .A(n27954), .B(n3291), .Z(n3292) );
  AND U4254 ( .A(n27955), .B(n3292), .Z(n3293) );
  NOR U4255 ( .A(n27959), .B(n3293), .Z(n3294) );
  NANDN U4256 ( .A(n27958), .B(n27957), .Z(n3295) );
  NAND U4257 ( .A(n3294), .B(n3295), .Z(n3296) );
  NAND U4258 ( .A(n27960), .B(n3296), .Z(n3297) );
  NANDN U4259 ( .A(n27961), .B(n3297), .Z(n3298) );
  AND U4260 ( .A(n27962), .B(n3298), .Z(n3299) );
  NANDN U4261 ( .A(n3299), .B(n24225), .Z(n3300) );
  NAND U4262 ( .A(n27963), .B(n3300), .Z(n3301) );
  NANDN U4263 ( .A(n27964), .B(n3301), .Z(n3302) );
  AND U4264 ( .A(n3302), .B(n24224), .Z(n3303) );
  OR U4265 ( .A(n24222), .B(n24223), .Z(n3304) );
  AND U4266 ( .A(n3303), .B(n3304), .Z(n3305) );
  OR U4267 ( .A(n27965), .B(n3305), .Z(n3306) );
  NANDN U4268 ( .A(n27966), .B(n3306), .Z(n3307) );
  NAND U4269 ( .A(n27967), .B(n3307), .Z(n27968) );
  AND U4270 ( .A(n8861), .B(n12816), .Z(n3308) );
  NAND U4271 ( .A(n27627), .B(n3308), .Z(n3309) );
  AND U4272 ( .A(n27630), .B(n3309), .Z(n3310) );
  ANDN U4273 ( .B(n27631), .A(n3310), .Z(n3311) );
  NAND U4274 ( .A(n12813), .B(n3311), .Z(n3312) );
  ANDN U4275 ( .B(n3312), .A(n19301), .Z(n3313) );
  NOR U4276 ( .A(n27635), .B(n12812), .Z(n3314) );
  NANDN U4277 ( .A(n27632), .B(n3313), .Z(n3315) );
  NAND U4278 ( .A(n3314), .B(n3315), .Z(n3316) );
  ANDN U4279 ( .B(n27636), .A(n19300), .Z(n3317) );
  NAND U4280 ( .A(n3316), .B(n3317), .Z(n3318) );
  NAND U4281 ( .A(n27637), .B(n3318), .Z(n3319) );
  ANDN U4282 ( .B(n3319), .A(n27638), .Z(n3320) );
  ANDN U4283 ( .B(n27640), .A(n19319), .Z(n3321) );
  NANDN U4284 ( .A(n3320), .B(n27639), .Z(n3322) );
  AND U4285 ( .A(n3321), .B(n3322), .Z(n3323) );
  NANDN U4286 ( .A(n3323), .B(n27641), .Z(n3324) );
  NAND U4287 ( .A(n19318), .B(n3324), .Z(n3325) );
  NANDN U4288 ( .A(n12807), .B(n3325), .Z(n8864) );
  OR U4289 ( .A(n24207), .B(n24208), .Z(n3326) );
  AND U4290 ( .A(n24209), .B(n3326), .Z(n3327) );
  AND U4291 ( .A(n24215), .B(n27993), .Z(n3328) );
  NAND U4292 ( .A(n24216), .B(n3328), .Z(n3329) );
  NANDN U4293 ( .A(n27994), .B(n3329), .Z(n3330) );
  NANDN U4294 ( .A(n27995), .B(n3330), .Z(n3331) );
  NAND U4295 ( .A(n27996), .B(n3331), .Z(n3332) );
  AND U4296 ( .A(n24212), .B(n3332), .Z(n3333) );
  OR U4297 ( .A(n24211), .B(n3333), .Z(n3334) );
  NAND U4298 ( .A(n24210), .B(n3334), .Z(n3335) );
  NAND U4299 ( .A(n27997), .B(n3335), .Z(n3336) );
  NANDN U4300 ( .A(n27998), .B(n3336), .Z(n3337) );
  NAND U4301 ( .A(n27999), .B(n3337), .Z(n3338) );
  ANDN U4302 ( .B(n3338), .A(n28000), .Z(n3339) );
  NANDN U4303 ( .A(n3339), .B(n28001), .Z(n3340) );
  NAND U4304 ( .A(n28002), .B(n3340), .Z(n3341) );
  NAND U4305 ( .A(n3327), .B(n3341), .Z(n28004) );
  ANDN U4306 ( .B(n12526), .A(n12525), .Z(n28056) );
  ANDN U4307 ( .B(n12732), .A(n19491), .Z(n3342) );
  NANDN U4308 ( .A(n12733), .B(n9017), .Z(n3343) );
  AND U4309 ( .A(n3342), .B(n3343), .Z(n27760) );
  NANDN U4310 ( .A(n28090), .B(n28089), .Z(n3344) );
  NAND U4311 ( .A(n28091), .B(n3344), .Z(n3345) );
  NANDN U4312 ( .A(n28092), .B(n3345), .Z(n3346) );
  NAND U4313 ( .A(n28093), .B(n3346), .Z(n3347) );
  NAND U4314 ( .A(n28094), .B(n3347), .Z(n3348) );
  AND U4315 ( .A(n24198), .B(n3348), .Z(n3349) );
  OR U4316 ( .A(n24197), .B(n3349), .Z(n3350) );
  NAND U4317 ( .A(n28095), .B(n3350), .Z(n3351) );
  NAND U4318 ( .A(n28096), .B(n3351), .Z(n3352) );
  NANDN U4319 ( .A(n28097), .B(n3352), .Z(n3353) );
  NANDN U4320 ( .A(n28098), .B(n3353), .Z(n3354) );
  ANDN U4321 ( .B(n3354), .A(n28099), .Z(n3355) );
  OR U4322 ( .A(n28100), .B(n3355), .Z(n3356) );
  NANDN U4323 ( .A(n28101), .B(n3356), .Z(n3357) );
  NAND U4324 ( .A(n28102), .B(n3357), .Z(n3358) );
  NAND U4325 ( .A(n28103), .B(n3358), .Z(n28105) );
  NAND U4326 ( .A(n28129), .B(n28128), .Z(n3359) );
  NANDN U4327 ( .A(n28130), .B(n3359), .Z(n3360) );
  NAND U4328 ( .A(n28131), .B(n3360), .Z(n3361) );
  AND U4329 ( .A(n3361), .B(n28134), .Z(n3362) );
  NAND U4330 ( .A(n28133), .B(n28132), .Z(n3363) );
  AND U4331 ( .A(n3362), .B(n3363), .Z(n3364) );
  OR U4332 ( .A(n28135), .B(n3364), .Z(n3365) );
  NANDN U4333 ( .A(n28136), .B(n3365), .Z(n3366) );
  NANDN U4334 ( .A(n28137), .B(n3366), .Z(n3367) );
  AND U4335 ( .A(n3367), .B(n28138), .Z(n3368) );
  NAND U4336 ( .A(n24184), .B(n24183), .Z(n3369) );
  AND U4337 ( .A(n3368), .B(n3369), .Z(n3370) );
  NANDN U4338 ( .A(n3370), .B(n24182), .Z(n3371) );
  NANDN U4339 ( .A(n28139), .B(n3371), .Z(n3372) );
  NANDN U4340 ( .A(n28140), .B(n3372), .Z(n28141) );
  NAND U4341 ( .A(n28167), .B(n28166), .Z(n3373) );
  NANDN U4342 ( .A(n28168), .B(n3373), .Z(n3374) );
  NAND U4343 ( .A(n28169), .B(n3374), .Z(n3375) );
  NAND U4344 ( .A(n28170), .B(n3375), .Z(n3376) );
  NAND U4345 ( .A(n28171), .B(n3376), .Z(n3377) );
  AND U4346 ( .A(n28172), .B(n3377), .Z(n3378) );
  NANDN U4347 ( .A(n3378), .B(n28173), .Z(n3379) );
  NANDN U4348 ( .A(n28174), .B(n3379), .Z(n3380) );
  NAND U4349 ( .A(n28175), .B(n3380), .Z(n3381) );
  NAND U4350 ( .A(n28176), .B(n3381), .Z(n3382) );
  NANDN U4351 ( .A(n28177), .B(n3382), .Z(n3383) );
  AND U4352 ( .A(n28178), .B(n3383), .Z(n3384) );
  OR U4353 ( .A(n28179), .B(n3384), .Z(n3385) );
  ANDN U4354 ( .B(n3385), .A(n24171), .Z(n3386) );
  NANDN U4355 ( .A(n3386), .B(n24170), .Z(n3387) );
  NAND U4356 ( .A(n28180), .B(n3387), .Z(n3388) );
  NAND U4357 ( .A(n28181), .B(n3388), .Z(n28184) );
  NANDN U4358 ( .A(n12627), .B(n9245), .Z(n3389) );
  ANDN U4359 ( .B(n3389), .A(n19781), .Z(n27920) );
  NANDN U4360 ( .A(n28212), .B(n28211), .Z(n3390) );
  NAND U4361 ( .A(n28213), .B(n3390), .Z(n3391) );
  AND U4362 ( .A(n28214), .B(n3391), .Z(n3392) );
  NANDN U4363 ( .A(n3392), .B(n24161), .Z(n3393) );
  AND U4364 ( .A(n28215), .B(n3393), .Z(n3394) );
  AND U4365 ( .A(n28217), .B(n28218), .Z(n3395) );
  NANDN U4366 ( .A(n3394), .B(n28216), .Z(n3396) );
  AND U4367 ( .A(n3395), .B(n3396), .Z(n3397) );
  NANDN U4368 ( .A(n3397), .B(n28219), .Z(n3398) );
  NAND U4369 ( .A(n28220), .B(n3398), .Z(n3399) );
  NAND U4370 ( .A(n28221), .B(n3399), .Z(n3400) );
  AND U4371 ( .A(n3400), .B(n24160), .Z(n3401) );
  NANDN U4372 ( .A(n24159), .B(n24158), .Z(n3402) );
  AND U4373 ( .A(n3401), .B(n3402), .Z(n3403) );
  NANDN U4374 ( .A(n3403), .B(n28222), .Z(n3404) );
  NANDN U4375 ( .A(n24157), .B(n3404), .Z(n3405) );
  NAND U4376 ( .A(n28223), .B(n3405), .Z(n28226) );
  NANDN U4377 ( .A(n20475), .B(n20474), .Z(n3406) );
  ANDN U4378 ( .B(n3406), .A(n20476), .Z(n28295) );
  ANDN U4379 ( .B(n20505), .A(n20504), .Z(n28311) );
  NANDN U4380 ( .A(n24148), .B(n28330), .Z(n3407) );
  NAND U4381 ( .A(n28331), .B(n3407), .Z(n3408) );
  NANDN U4382 ( .A(n28332), .B(n3408), .Z(n3409) );
  NAND U4383 ( .A(n28333), .B(n3409), .Z(n3410) );
  NANDN U4384 ( .A(n28334), .B(n3410), .Z(n3411) );
  AND U4385 ( .A(n28335), .B(n3411), .Z(n3412) );
  OR U4386 ( .A(n28336), .B(n3412), .Z(n3413) );
  NAND U4387 ( .A(n28337), .B(n3413), .Z(n3414) );
  NANDN U4388 ( .A(n28338), .B(n3414), .Z(n3415) );
  NAND U4389 ( .A(n28339), .B(n3415), .Z(n3416) );
  NANDN U4390 ( .A(n28340), .B(n3416), .Z(n3417) );
  ANDN U4391 ( .B(n3417), .A(n24147), .Z(n3418) );
  NANDN U4392 ( .A(n3418), .B(n28341), .Z(n3419) );
  NAND U4393 ( .A(n28342), .B(n3419), .Z(n3420) );
  NANDN U4394 ( .A(n28343), .B(n3420), .Z(n3421) );
  NAND U4395 ( .A(n28344), .B(n3421), .Z(n3422) );
  NANDN U4396 ( .A(n28345), .B(n3422), .Z(n3423) );
  AND U4397 ( .A(n28346), .B(n3423), .Z(n28348) );
  OR U4398 ( .A(n19999), .B(n9392), .Z(n3424) );
  NAND U4399 ( .A(n28023), .B(n3424), .Z(n3425) );
  NANDN U4400 ( .A(n28026), .B(n3425), .Z(n3426) );
  NAND U4401 ( .A(n28029), .B(n3426), .Z(n3427) );
  NANDN U4402 ( .A(n28030), .B(n3427), .Z(n3428) );
  AND U4403 ( .A(n28031), .B(n3428), .Z(n3429) );
  AND U4404 ( .A(n12543), .B(n24206), .Z(n3430) );
  OR U4405 ( .A(n28032), .B(n3429), .Z(n3431) );
  AND U4406 ( .A(n3430), .B(n3431), .Z(n3432) );
  NOR U4407 ( .A(n28035), .B(n12544), .Z(n3433) );
  NANDN U4408 ( .A(n3432), .B(n3433), .Z(n3434) );
  AND U4409 ( .A(n12542), .B(n3434), .Z(n3435) );
  AND U4410 ( .A(n12541), .B(n3435), .Z(n3436) );
  NOR U4411 ( .A(n28039), .B(n24203), .Z(n3437) );
  NANDN U4412 ( .A(n3436), .B(n24204), .Z(n3438) );
  AND U4413 ( .A(n3437), .B(n3438), .Z(n3439) );
  NANDN U4414 ( .A(n3439), .B(n24205), .Z(n3440) );
  NAND U4415 ( .A(n28037), .B(n3440), .Z(n3441) );
  NAND U4416 ( .A(n24202), .B(n3441), .Z(n9394) );
  NANDN U4417 ( .A(n28375), .B(n28374), .Z(n3442) );
  NAND U4418 ( .A(n28377), .B(n3442), .Z(n3443) );
  NAND U4419 ( .A(n28378), .B(n3443), .Z(n3444) );
  NAND U4420 ( .A(n28379), .B(n3444), .Z(n3445) );
  NAND U4421 ( .A(n28380), .B(n3445), .Z(n3446) );
  ANDN U4422 ( .B(n3446), .A(n24139), .Z(n3447) );
  NANDN U4423 ( .A(n3447), .B(n28381), .Z(n3448) );
  NAND U4424 ( .A(n28382), .B(n3448), .Z(n3449) );
  NAND U4425 ( .A(n28383), .B(n3449), .Z(n3450) );
  NANDN U4426 ( .A(n28384), .B(n3450), .Z(n3451) );
  NAND U4427 ( .A(n28385), .B(n3451), .Z(n3452) );
  ANDN U4428 ( .B(n3452), .A(n28386), .Z(n3453) );
  OR U4429 ( .A(n24138), .B(n3453), .Z(n3454) );
  NAND U4430 ( .A(n24137), .B(n3454), .Z(n3455) );
  NANDN U4431 ( .A(n28387), .B(n3455), .Z(n3456) );
  NANDN U4432 ( .A(n28388), .B(n3456), .Z(n28389) );
  ANDN U4433 ( .B(n28412), .A(n28413), .Z(n3457) );
  NANDN U4434 ( .A(n28414), .B(n28415), .Z(n3458) );
  NAND U4435 ( .A(n3457), .B(n3458), .Z(n3459) );
  NANDN U4436 ( .A(n28416), .B(n3459), .Z(n3460) );
  NAND U4437 ( .A(n28417), .B(n3460), .Z(n3461) );
  ANDN U4438 ( .B(n3461), .A(n28418), .Z(n3462) );
  OR U4439 ( .A(n28419), .B(n3462), .Z(n3463) );
  NAND U4440 ( .A(n28420), .B(n3463), .Z(n3464) );
  NAND U4441 ( .A(n28421), .B(n3464), .Z(n3465) );
  NAND U4442 ( .A(n28422), .B(n3465), .Z(n3466) );
  NAND U4443 ( .A(n24126), .B(n3466), .Z(n3467) );
  ANDN U4444 ( .B(n3467), .A(n24125), .Z(n3468) );
  NANDN U4445 ( .A(n3468), .B(n24124), .Z(n3469) );
  NANDN U4446 ( .A(n24123), .B(n3469), .Z(n3470) );
  NAND U4447 ( .A(n28423), .B(n3470), .Z(n28424) );
  NAND U4448 ( .A(n28457), .B(n28456), .Z(n3471) );
  NAND U4449 ( .A(n28458), .B(n3471), .Z(n3472) );
  ANDN U4450 ( .B(n3472), .A(n24114), .Z(n3473) );
  OR U4451 ( .A(n28459), .B(n3473), .Z(n3474) );
  NAND U4452 ( .A(n28460), .B(n3474), .Z(n3475) );
  NANDN U4453 ( .A(n28461), .B(n3475), .Z(n3476) );
  AND U4454 ( .A(n28463), .B(n28462), .Z(n3477) );
  NAND U4455 ( .A(n3476), .B(n3477), .Z(n3478) );
  NANDN U4456 ( .A(n28464), .B(n3478), .Z(n3479) );
  NAND U4457 ( .A(n28465), .B(n3479), .Z(n3480) );
  NAND U4458 ( .A(n28466), .B(n3480), .Z(n3481) );
  ANDN U4459 ( .B(n3481), .A(n28467), .Z(n3482) );
  NANDN U4460 ( .A(n3482), .B(n28468), .Z(n3483) );
  AND U4461 ( .A(n28469), .B(n3483), .Z(n3484) );
  NANDN U4462 ( .A(n3484), .B(n28470), .Z(n3485) );
  NAND U4463 ( .A(n28471), .B(n3485), .Z(n3486) );
  NAND U4464 ( .A(n28472), .B(n3486), .Z(n28473) );
  NANDN U4465 ( .A(n24107), .B(n24106), .Z(n3487) );
  ANDN U4466 ( .B(n3487), .A(n24108), .Z(n3488) );
  NAND U4467 ( .A(n28501), .B(n28502), .Z(n3489) );
  NAND U4468 ( .A(n3488), .B(n3489), .Z(n3490) );
  NAND U4469 ( .A(n28503), .B(n3490), .Z(n3491) );
  NAND U4470 ( .A(n28504), .B(n3491), .Z(n3492) );
  NAND U4471 ( .A(n28505), .B(n3492), .Z(n3493) );
  AND U4472 ( .A(n24105), .B(n3493), .Z(n3494) );
  NOR U4473 ( .A(n28506), .B(n3494), .Z(n3495) );
  NAND U4474 ( .A(n24104), .B(n3495), .Z(n3496) );
  AND U4475 ( .A(n28507), .B(n3496), .Z(n3497) );
  NANDN U4476 ( .A(n3497), .B(n28508), .Z(n3498) );
  NANDN U4477 ( .A(n28509), .B(n3498), .Z(n3499) );
  NAND U4478 ( .A(n28510), .B(n3499), .Z(n3500) );
  NANDN U4479 ( .A(n28511), .B(n3500), .Z(n28512) );
  NANDN U4480 ( .A(n21004), .B(n21003), .Z(n3501) );
  AND U4481 ( .A(n21005), .B(n3501), .Z(n28552) );
  NANDN U4482 ( .A(n12383), .B(n9702), .Z(n3502) );
  AND U4483 ( .A(n20434), .B(n3502), .Z(n28251) );
  NAND U4484 ( .A(n28575), .B(n28576), .Z(n3503) );
  NANDN U4485 ( .A(n28577), .B(n3503), .Z(n3504) );
  NAND U4486 ( .A(n28578), .B(n3504), .Z(n3505) );
  NAND U4487 ( .A(n28579), .B(n3505), .Z(n3506) );
  NANDN U4488 ( .A(n24093), .B(n3506), .Z(n3507) );
  AND U4489 ( .A(n24092), .B(n3507), .Z(n3508) );
  OR U4490 ( .A(n3508), .B(n28580), .Z(n3509) );
  NAND U4491 ( .A(n28581), .B(n3509), .Z(n3510) );
  ANDN U4492 ( .B(n3510), .A(n28582), .Z(n3511) );
  NANDN U4493 ( .A(n3511), .B(n28583), .Z(n3512) );
  ANDN U4494 ( .B(n3512), .A(n28584), .Z(n3513) );
  NANDN U4495 ( .A(n3513), .B(n24091), .Z(n3514) );
  NANDN U4496 ( .A(n28585), .B(n3514), .Z(n3515) );
  NAND U4497 ( .A(n28586), .B(n3515), .Z(n28587) );
  NANDN U4498 ( .A(n28615), .B(n28614), .Z(n3516) );
  NAND U4499 ( .A(n28616), .B(n3516), .Z(n3517) );
  AND U4500 ( .A(n28617), .B(n3517), .Z(n3518) );
  OR U4501 ( .A(n24085), .B(n3518), .Z(n3519) );
  NAND U4502 ( .A(n28618), .B(n3519), .Z(n3520) );
  NANDN U4503 ( .A(n28619), .B(n3520), .Z(n3521) );
  NAND U4504 ( .A(n28620), .B(n3521), .Z(n3522) );
  NANDN U4505 ( .A(n28621), .B(n3522), .Z(n3523) );
  AND U4506 ( .A(n28622), .B(n3523), .Z(n3524) );
  OR U4507 ( .A(n3524), .B(n28623), .Z(n3525) );
  NAND U4508 ( .A(n28624), .B(n3525), .Z(n3526) );
  ANDN U4509 ( .B(n3526), .A(n28625), .Z(n3527) );
  NANDN U4510 ( .A(n3527), .B(n28626), .Z(n3528) );
  NANDN U4511 ( .A(n24084), .B(n3528), .Z(n3529) );
  NAND U4512 ( .A(n24083), .B(n3529), .Z(n3530) );
  NAND U4513 ( .A(n28627), .B(n3530), .Z(n28630) );
  NAND U4514 ( .A(n28654), .B(n24075), .Z(n3531) );
  NANDN U4515 ( .A(n28655), .B(n3531), .Z(n3532) );
  NAND U4516 ( .A(n28656), .B(n3532), .Z(n3533) );
  NANDN U4517 ( .A(n24074), .B(n3533), .Z(n3534) );
  NAND U4518 ( .A(n24073), .B(n3534), .Z(n3535) );
  ANDN U4519 ( .B(n3535), .A(n28657), .Z(n3536) );
  NANDN U4520 ( .A(n3536), .B(n28658), .Z(n3537) );
  NANDN U4521 ( .A(n28659), .B(n3537), .Z(n3538) );
  NAND U4522 ( .A(n28660), .B(n3538), .Z(n3539) );
  NAND U4523 ( .A(n28661), .B(n3539), .Z(n3540) );
  NANDN U4524 ( .A(n28662), .B(n3540), .Z(n3541) );
  AND U4525 ( .A(n28663), .B(n3541), .Z(n3542) );
  OR U4526 ( .A(n3542), .B(n28664), .Z(n3543) );
  NAND U4527 ( .A(n28665), .B(n3543), .Z(n3544) );
  NANDN U4528 ( .A(n28666), .B(n3544), .Z(n28667) );
  NANDN U4529 ( .A(n28685), .B(n28684), .Z(n3545) );
  NANDN U4530 ( .A(n28686), .B(n3545), .Z(n3546) );
  AND U4531 ( .A(n28687), .B(n3546), .Z(n3547) );
  OR U4532 ( .A(n3547), .B(n28688), .Z(n3548) );
  NAND U4533 ( .A(n28689), .B(n3548), .Z(n3549) );
  NANDN U4534 ( .A(n28690), .B(n3549), .Z(n3550) );
  NAND U4535 ( .A(n24061), .B(n3550), .Z(n3551) );
  NANDN U4536 ( .A(n28691), .B(n3551), .Z(n3552) );
  AND U4537 ( .A(n28692), .B(n3552), .Z(n3553) );
  NANDN U4538 ( .A(n3553), .B(n28693), .Z(n3554) );
  ANDN U4539 ( .B(n3554), .A(n28694), .Z(n3555) );
  NANDN U4540 ( .A(n3555), .B(n24060), .Z(n3556) );
  NANDN U4541 ( .A(n28695), .B(n3556), .Z(n3557) );
  NAND U4542 ( .A(n28696), .B(n3557), .Z(n28697) );
  NANDN U4543 ( .A(n28720), .B(n28719), .Z(n3558) );
  NANDN U4544 ( .A(n28721), .B(n3558), .Z(n3559) );
  AND U4545 ( .A(n28722), .B(n3559), .Z(n3560) );
  OR U4546 ( .A(n3560), .B(n28723), .Z(n3561) );
  NAND U4547 ( .A(n28724), .B(n3561), .Z(n3562) );
  ANDN U4548 ( .B(n3562), .A(n28725), .Z(n3563) );
  NANDN U4549 ( .A(n3563), .B(n24051), .Z(n3564) );
  NAND U4550 ( .A(n28726), .B(n3564), .Z(n3565) );
  NANDN U4551 ( .A(n28727), .B(n3565), .Z(n3566) );
  NAND U4552 ( .A(n28728), .B(n3566), .Z(n3567) );
  NANDN U4553 ( .A(n28729), .B(n3567), .Z(n3568) );
  AND U4554 ( .A(n28730), .B(n3568), .Z(n3569) );
  OR U4555 ( .A(n28731), .B(n3569), .Z(n3570) );
  NAND U4556 ( .A(n28732), .B(n3570), .Z(n3571) );
  NANDN U4557 ( .A(n24050), .B(n3571), .Z(n3572) );
  NAND U4558 ( .A(n24049), .B(n3572), .Z(n28735) );
  NAND U4559 ( .A(n20952), .B(n10065), .Z(n3573) );
  ANDN U4560 ( .B(n3573), .A(n20958), .Z(n28530) );
  NAND U4561 ( .A(n28759), .B(n28758), .Z(n3574) );
  NAND U4562 ( .A(n28760), .B(n3574), .Z(n3575) );
  ANDN U4563 ( .B(n3575), .A(n24040), .Z(n3576) );
  NANDN U4564 ( .A(n3576), .B(n28761), .Z(n3577) );
  NANDN U4565 ( .A(n28762), .B(n3577), .Z(n3578) );
  NAND U4566 ( .A(n28763), .B(n3578), .Z(n3579) );
  NAND U4567 ( .A(n28764), .B(n3579), .Z(n3580) );
  NANDN U4568 ( .A(n24039), .B(n3580), .Z(n3581) );
  AND U4569 ( .A(n24038), .B(n3581), .Z(n3582) );
  OR U4570 ( .A(n3582), .B(n28765), .Z(n3583) );
  NAND U4571 ( .A(n28766), .B(n3583), .Z(n3584) );
  ANDN U4572 ( .B(n3584), .A(n28767), .Z(n3585) );
  NANDN U4573 ( .A(n3585), .B(n28768), .Z(n3586) );
  NANDN U4574 ( .A(n28769), .B(n3586), .Z(n3587) );
  NAND U4575 ( .A(n24037), .B(n3587), .Z(n28772) );
  NAND U4576 ( .A(n28792), .B(n28791), .Z(n3588) );
  NANDN U4577 ( .A(n28794), .B(n3588), .Z(n3589) );
  ANDN U4578 ( .B(n3589), .A(n24027), .Z(n3590) );
  NANDN U4579 ( .A(n3590), .B(n24026), .Z(n3591) );
  ANDN U4580 ( .B(n3591), .A(n28795), .Z(n3592) );
  ANDN U4581 ( .B(n24025), .A(n24024), .Z(n3593) );
  NANDN U4582 ( .A(n3592), .B(n28796), .Z(n3594) );
  AND U4583 ( .A(n3593), .B(n3594), .Z(n3595) );
  NOR U4584 ( .A(n28798), .B(n28799), .Z(n3596) );
  NANDN U4585 ( .A(n3595), .B(n28797), .Z(n3597) );
  AND U4586 ( .A(n3596), .B(n3597), .Z(n3598) );
  OR U4587 ( .A(n28800), .B(n3598), .Z(n3599) );
  NAND U4588 ( .A(n28801), .B(n3599), .Z(n3600) );
  NANDN U4589 ( .A(n24023), .B(n3600), .Z(n28802) );
  ANDN U4590 ( .B(n24014), .A(n24013), .Z(n3601) );
  NAND U4591 ( .A(n28827), .B(n28826), .Z(n3602) );
  AND U4592 ( .A(n3601), .B(n3602), .Z(n3603) );
  ANDN U4593 ( .B(n28829), .A(n28830), .Z(n3604) );
  OR U4594 ( .A(n28828), .B(n3603), .Z(n3605) );
  AND U4595 ( .A(n3604), .B(n3605), .Z(n3606) );
  OR U4596 ( .A(n28831), .B(n3606), .Z(n3607) );
  NAND U4597 ( .A(n28832), .B(n3607), .Z(n3608) );
  NANDN U4598 ( .A(n24012), .B(n3608), .Z(n3609) );
  AND U4599 ( .A(n28833), .B(n3609), .Z(n3610) );
  AND U4600 ( .A(n24010), .B(n24009), .Z(n3611) );
  OR U4601 ( .A(n24011), .B(n3610), .Z(n3612) );
  AND U4602 ( .A(n3611), .B(n3612), .Z(n3613) );
  OR U4603 ( .A(n28834), .B(n3613), .Z(n3614) );
  NAND U4604 ( .A(n28835), .B(n3614), .Z(n3615) );
  NANDN U4605 ( .A(n28836), .B(n3615), .Z(n28837) );
  NANDN U4606 ( .A(n24000), .B(n28857), .Z(n3616) );
  NAND U4607 ( .A(n28858), .B(n3616), .Z(n3617) );
  NANDN U4608 ( .A(n28859), .B(n3617), .Z(n3618) );
  NAND U4609 ( .A(n28860), .B(n3618), .Z(n3619) );
  NANDN U4610 ( .A(n23999), .B(n3619), .Z(n3620) );
  AND U4611 ( .A(n23998), .B(n3620), .Z(n3621) );
  OR U4612 ( .A(n28861), .B(n3621), .Z(n3622) );
  NAND U4613 ( .A(n28862), .B(n3622), .Z(n3623) );
  NANDN U4614 ( .A(n28863), .B(n3623), .Z(n3624) );
  NAND U4615 ( .A(n28864), .B(n3624), .Z(n3625) );
  NANDN U4616 ( .A(n28865), .B(n3625), .Z(n3626) );
  AND U4617 ( .A(n28866), .B(n3626), .Z(n3627) );
  OR U4618 ( .A(n3627), .B(n28867), .Z(n3628) );
  AND U4619 ( .A(n28868), .B(n3628), .Z(n28870) );
  NAND U4620 ( .A(n28893), .B(n23990), .Z(n3629) );
  NAND U4621 ( .A(n28894), .B(n3629), .Z(n3630) );
  NANDN U4622 ( .A(n28895), .B(n3630), .Z(n3631) );
  NAND U4623 ( .A(n28896), .B(n3631), .Z(n3632) );
  NANDN U4624 ( .A(n28897), .B(n3632), .Z(n3633) );
  AND U4625 ( .A(n28898), .B(n3633), .Z(n3634) );
  OR U4626 ( .A(n3634), .B(n28899), .Z(n3635) );
  NAND U4627 ( .A(n28900), .B(n3635), .Z(n3636) );
  AND U4628 ( .A(n28901), .B(n3636), .Z(n3637) );
  AND U4629 ( .A(n28903), .B(n28902), .Z(n3638) );
  OR U4630 ( .A(n23989), .B(n3637), .Z(n3639) );
  AND U4631 ( .A(n3638), .B(n3639), .Z(n3640) );
  NANDN U4632 ( .A(n3640), .B(n28904), .Z(n3641) );
  NAND U4633 ( .A(n28905), .B(n3641), .Z(n3642) );
  NANDN U4634 ( .A(n28906), .B(n3642), .Z(n28907) );
  ANDN U4635 ( .B(n28930), .A(n28931), .Z(n3643) );
  NAND U4636 ( .A(n23980), .B(n28929), .Z(n3644) );
  AND U4637 ( .A(n3643), .B(n3644), .Z(n3645) );
  OR U4638 ( .A(n23979), .B(n3645), .Z(n3646) );
  NAND U4639 ( .A(n23978), .B(n3646), .Z(n3647) );
  NAND U4640 ( .A(n28932), .B(n3647), .Z(n3648) );
  AND U4641 ( .A(n28934), .B(n28933), .Z(n3649) );
  NAND U4642 ( .A(n3648), .B(n3649), .Z(n3650) );
  NAND U4643 ( .A(n23977), .B(n3650), .Z(n3651) );
  AND U4644 ( .A(n28935), .B(n28936), .Z(n3652) );
  NAND U4645 ( .A(n3651), .B(n3652), .Z(n3653) );
  NANDN U4646 ( .A(n28937), .B(n3653), .Z(n3654) );
  AND U4647 ( .A(n28938), .B(n28939), .Z(n3655) );
  NAND U4648 ( .A(n3654), .B(n3655), .Z(n3656) );
  NAND U4649 ( .A(n28940), .B(n3656), .Z(n28941) );
  NAND U4650 ( .A(n28975), .B(n28974), .Z(n3657) );
  NAND U4651 ( .A(n28977), .B(n3657), .Z(n3658) );
  AND U4652 ( .A(n28978), .B(n3658), .Z(n3659) );
  OR U4653 ( .A(n28979), .B(n3659), .Z(n3660) );
  NAND U4654 ( .A(n28980), .B(n3660), .Z(n3661) );
  NANDN U4655 ( .A(n23971), .B(n3661), .Z(n3662) );
  NAND U4656 ( .A(n23970), .B(n3662), .Z(n3663) );
  NANDN U4657 ( .A(n28981), .B(n3663), .Z(n3664) );
  AND U4658 ( .A(n28982), .B(n3664), .Z(n3665) );
  OR U4659 ( .A(n28983), .B(n3665), .Z(n3666) );
  AND U4660 ( .A(n28984), .B(n3666), .Z(n3667) );
  OR U4661 ( .A(n28985), .B(n3667), .Z(n3668) );
  NANDN U4662 ( .A(n28986), .B(n3668), .Z(n3669) );
  NAND U4663 ( .A(n28987), .B(n3669), .Z(n28988) );
  NAND U4664 ( .A(n29017), .B(n29016), .Z(n3670) );
  AND U4665 ( .A(n29019), .B(n3670), .Z(n3671) );
  NOR U4666 ( .A(n23963), .B(n3671), .Z(n3672) );
  NAND U4667 ( .A(n23962), .B(n3672), .Z(n3673) );
  NANDN U4668 ( .A(n29020), .B(n3673), .Z(n3674) );
  AND U4669 ( .A(n29022), .B(n29021), .Z(n3675) );
  NAND U4670 ( .A(n3674), .B(n3675), .Z(n3676) );
  NANDN U4671 ( .A(n29023), .B(n3676), .Z(n3677) );
  AND U4672 ( .A(n29025), .B(n29024), .Z(n3678) );
  NAND U4673 ( .A(n3677), .B(n3678), .Z(n3679) );
  NANDN U4674 ( .A(n29026), .B(n3679), .Z(n3680) );
  NAND U4675 ( .A(n29027), .B(n3680), .Z(n3681) );
  NANDN U4676 ( .A(n29028), .B(n3681), .Z(n3682) );
  AND U4677 ( .A(n29029), .B(n3682), .Z(n3683) );
  OR U4678 ( .A(n29030), .B(n3683), .Z(n3684) );
  NAND U4679 ( .A(n29031), .B(n3684), .Z(n3685) );
  NANDN U4680 ( .A(n29032), .B(n3685), .Z(n29033) );
  NAND U4681 ( .A(n29068), .B(n29067), .Z(n3686) );
  NAND U4682 ( .A(n29069), .B(n3686), .Z(n3687) );
  ANDN U4683 ( .B(n3687), .A(n23958), .Z(n3688) );
  NANDN U4684 ( .A(n3688), .B(n23957), .Z(n3689) );
  NAND U4685 ( .A(n29070), .B(n3689), .Z(n3690) );
  NANDN U4686 ( .A(n29071), .B(n3690), .Z(n3691) );
  AND U4687 ( .A(n23956), .B(n23955), .Z(n3692) );
  NAND U4688 ( .A(n3691), .B(n3692), .Z(n3693) );
  NANDN U4689 ( .A(n29072), .B(n3693), .Z(n3694) );
  NAND U4690 ( .A(n29073), .B(n3694), .Z(n3695) );
  NANDN U4691 ( .A(n29074), .B(n3695), .Z(n3696) );
  AND U4692 ( .A(n29075), .B(n3696), .Z(n3697) );
  NANDN U4693 ( .A(n3697), .B(n29076), .Z(n3698) );
  NANDN U4694 ( .A(n23954), .B(n3698), .Z(n3699) );
  NAND U4695 ( .A(n29077), .B(n3699), .Z(n29078) );
  NAND U4696 ( .A(n29106), .B(n29107), .Z(n3700) );
  NAND U4697 ( .A(n29108), .B(n3700), .Z(n3701) );
  NANDN U4698 ( .A(n23946), .B(n3701), .Z(n3702) );
  NAND U4699 ( .A(n23945), .B(n3702), .Z(n3703) );
  NANDN U4700 ( .A(n29109), .B(n3703), .Z(n3704) );
  AND U4701 ( .A(n29110), .B(n3704), .Z(n3705) );
  OR U4702 ( .A(n29111), .B(n3705), .Z(n3706) );
  AND U4703 ( .A(n29112), .B(n3706), .Z(n3707) );
  OR U4704 ( .A(n23944), .B(n3707), .Z(n3708) );
  NAND U4705 ( .A(n29113), .B(n3708), .Z(n3709) );
  NAND U4706 ( .A(n29114), .B(n3709), .Z(n3710) );
  AND U4707 ( .A(n29115), .B(n29116), .Z(n3711) );
  NAND U4708 ( .A(n3710), .B(n3711), .Z(n3712) );
  NANDN U4709 ( .A(n29117), .B(n3712), .Z(n29118) );
  NAND U4710 ( .A(n29149), .B(n29148), .Z(n3713) );
  NANDN U4711 ( .A(n29150), .B(n3713), .Z(n3714) );
  AND U4712 ( .A(n29151), .B(n3714), .Z(n3715) );
  OR U4713 ( .A(n3715), .B(n29152), .Z(n3716) );
  NAND U4714 ( .A(n29153), .B(n3716), .Z(n3717) );
  NANDN U4715 ( .A(n29154), .B(n3717), .Z(n3718) );
  NAND U4716 ( .A(n29155), .B(n3718), .Z(n3719) );
  NANDN U4717 ( .A(n29156), .B(n3719), .Z(n3720) );
  AND U4718 ( .A(n29157), .B(n3720), .Z(n3721) );
  OR U4719 ( .A(n3721), .B(n29158), .Z(n3722) );
  NAND U4720 ( .A(n29159), .B(n3722), .Z(n3723) );
  NAND U4721 ( .A(n23939), .B(n3723), .Z(n3724) );
  NANDN U4722 ( .A(n29160), .B(n3724), .Z(n3725) );
  NAND U4723 ( .A(n29161), .B(n3725), .Z(n3726) );
  ANDN U4724 ( .B(n3726), .A(n29162), .Z(n3727) );
  NANDN U4725 ( .A(n3727), .B(n29163), .Z(n3728) );
  NANDN U4726 ( .A(n29164), .B(n3728), .Z(n3729) );
  NAND U4727 ( .A(n29165), .B(n3729), .Z(n29166) );
  NANDN U4728 ( .A(n29185), .B(n29184), .Z(n3730) );
  AND U4729 ( .A(n29187), .B(n3730), .Z(n3731) );
  ANDN U4730 ( .B(n29189), .A(n3731), .Z(n3732) );
  NAND U4731 ( .A(n29188), .B(n3732), .Z(n3733) );
  NANDN U4732 ( .A(n29190), .B(n3733), .Z(n3734) );
  NAND U4733 ( .A(n29191), .B(n3734), .Z(n3735) );
  NANDN U4734 ( .A(n23928), .B(n3735), .Z(n3736) );
  AND U4735 ( .A(n23927), .B(n3736), .Z(n3737) );
  OR U4736 ( .A(n29192), .B(n3737), .Z(n3738) );
  NAND U4737 ( .A(n29193), .B(n3738), .Z(n3739) );
  NANDN U4738 ( .A(n29194), .B(n3739), .Z(n3740) );
  NAND U4739 ( .A(n29195), .B(n3740), .Z(n29196) );
  NAND U4740 ( .A(n29233), .B(n29232), .Z(n3741) );
  NANDN U4741 ( .A(n23921), .B(n3741), .Z(n3742) );
  AND U4742 ( .A(n29234), .B(n3742), .Z(n3743) );
  NANDN U4743 ( .A(n29235), .B(n3743), .Z(n3744) );
  NANDN U4744 ( .A(n29236), .B(n3744), .Z(n3745) );
  AND U4745 ( .A(n29237), .B(n3745), .Z(n3746) );
  NAND U4746 ( .A(n29238), .B(n3746), .Z(n3747) );
  NANDN U4747 ( .A(n29239), .B(n3747), .Z(n3748) );
  NAND U4748 ( .A(n29240), .B(n3748), .Z(n3749) );
  NANDN U4749 ( .A(n3749), .B(n29241), .Z(n3750) );
  NANDN U4750 ( .A(n29242), .B(n3750), .Z(n3751) );
  NAND U4751 ( .A(n29243), .B(n3751), .Z(n3752) );
  AND U4752 ( .A(n29245), .B(n29246), .Z(n3753) );
  NANDN U4753 ( .A(n29244), .B(n3752), .Z(n3754) );
  NAND U4754 ( .A(n3753), .B(n3754), .Z(n3755) );
  AND U4755 ( .A(n29249), .B(n29248), .Z(n3756) );
  NANDN U4756 ( .A(n29247), .B(n3755), .Z(n3757) );
  NAND U4757 ( .A(n3756), .B(n3757), .Z(n3758) );
  NANDN U4758 ( .A(n29250), .B(n3758), .Z(n29251) );
  NAND U4759 ( .A(n29277), .B(n29278), .Z(n3759) );
  ANDN U4760 ( .B(n3759), .A(n29279), .Z(n3760) );
  NOR U4761 ( .A(n29281), .B(n3760), .Z(n3761) );
  NAND U4762 ( .A(n29280), .B(n3761), .Z(n3762) );
  NANDN U4763 ( .A(n29282), .B(n3762), .Z(n3763) );
  ANDN U4764 ( .B(n23910), .A(n23909), .Z(n3764) );
  NAND U4765 ( .A(n3763), .B(n3764), .Z(n3765) );
  NANDN U4766 ( .A(n29283), .B(n3765), .Z(n3766) );
  NAND U4767 ( .A(n29284), .B(n3766), .Z(n3767) );
  NANDN U4768 ( .A(n29285), .B(n3767), .Z(n3768) );
  AND U4769 ( .A(n29286), .B(n3768), .Z(n3769) );
  AND U4770 ( .A(n23908), .B(n23907), .Z(n3770) );
  OR U4771 ( .A(n29287), .B(n3769), .Z(n3771) );
  AND U4772 ( .A(n3770), .B(n3771), .Z(n3772) );
  OR U4773 ( .A(n29288), .B(n3772), .Z(n3773) );
  AND U4774 ( .A(n29289), .B(n3773), .Z(n3774) );
  OR U4775 ( .A(n29290), .B(n3774), .Z(n3775) );
  NAND U4776 ( .A(n29291), .B(n3775), .Z(n3776) );
  NANDN U4777 ( .A(n29292), .B(n3776), .Z(n29293) );
  NANDN U4778 ( .A(n29320), .B(n29319), .Z(n3777) );
  NANDN U4779 ( .A(n29321), .B(n3777), .Z(n3778) );
  NAND U4780 ( .A(n29322), .B(n3778), .Z(n3779) );
  NANDN U4781 ( .A(n23900), .B(n3779), .Z(n3780) );
  NAND U4782 ( .A(n23899), .B(n3780), .Z(n3781) );
  AND U4783 ( .A(n29323), .B(n3781), .Z(n3782) );
  ANDN U4784 ( .B(n29324), .A(n3782), .Z(n3783) );
  NAND U4785 ( .A(n29325), .B(n3783), .Z(n3784) );
  ANDN U4786 ( .B(n3784), .A(n29326), .Z(n3785) );
  NOR U4787 ( .A(n23898), .B(n3785), .Z(n3786) );
  NAND U4788 ( .A(n29327), .B(n3786), .Z(n3787) );
  ANDN U4789 ( .B(n3787), .A(n29328), .Z(n3788) );
  NANDN U4790 ( .A(n3788), .B(n29329), .Z(n3789) );
  NANDN U4791 ( .A(n29330), .B(n3789), .Z(n3790) );
  NAND U4792 ( .A(n29331), .B(n3790), .Z(n29332) );
  NAND U4793 ( .A(n29366), .B(n29365), .Z(n3791) );
  NAND U4794 ( .A(n29367), .B(n3791), .Z(n3792) );
  ANDN U4795 ( .B(n3792), .A(n29368), .Z(n3793) );
  ANDN U4796 ( .B(n23894), .A(n3793), .Z(n3794) );
  NAND U4797 ( .A(n23893), .B(n3794), .Z(n3795) );
  ANDN U4798 ( .B(n3795), .A(n29369), .Z(n3796) );
  ANDN U4799 ( .B(n29371), .A(n3796), .Z(n3797) );
  NAND U4800 ( .A(n29370), .B(n3797), .Z(n3798) );
  ANDN U4801 ( .B(n3798), .A(n29372), .Z(n3799) );
  NANDN U4802 ( .A(n3799), .B(n29373), .Z(n3800) );
  NANDN U4803 ( .A(n23892), .B(n3800), .Z(n3801) );
  NAND U4804 ( .A(n23891), .B(n3801), .Z(n29376) );
  NANDN U4805 ( .A(n29406), .B(n29405), .Z(n3802) );
  NAND U4806 ( .A(n29408), .B(n3802), .Z(n3803) );
  AND U4807 ( .A(n29409), .B(n3803), .Z(n3804) );
  OR U4808 ( .A(n3804), .B(n29410), .Z(n3805) );
  NAND U4809 ( .A(n29411), .B(n3805), .Z(n3806) );
  NANDN U4810 ( .A(n29412), .B(n3806), .Z(n3807) );
  NAND U4811 ( .A(n29413), .B(n3807), .Z(n3808) );
  NAND U4812 ( .A(n23885), .B(n3808), .Z(n3809) );
  ANDN U4813 ( .B(n3809), .A(n29414), .Z(n3810) );
  NANDN U4814 ( .A(n3810), .B(n29415), .Z(n3811) );
  ANDN U4815 ( .B(n3811), .A(n29416), .Z(n3812) );
  NANDN U4816 ( .A(n3812), .B(n29417), .Z(n3813) );
  NANDN U4817 ( .A(n23884), .B(n3813), .Z(n3814) );
  NAND U4818 ( .A(n23883), .B(n3814), .Z(n29420) );
  NAND U4819 ( .A(n29443), .B(n29444), .Z(n3815) );
  NANDN U4820 ( .A(n29445), .B(n3815), .Z(n3816) );
  AND U4821 ( .A(n29446), .B(n3816), .Z(n3817) );
  OR U4822 ( .A(n29447), .B(n3817), .Z(n3818) );
  NAND U4823 ( .A(n29448), .B(n3818), .Z(n3819) );
  NAND U4824 ( .A(n29449), .B(n3819), .Z(n3820) );
  OR U4825 ( .A(n3820), .B(n29450), .Z(n3821) );
  NANDN U4826 ( .A(n29451), .B(n3821), .Z(n3822) );
  NAND U4827 ( .A(n29452), .B(n3822), .Z(n3823) );
  AND U4828 ( .A(n29454), .B(n29455), .Z(n3824) );
  NANDN U4829 ( .A(n29453), .B(n3823), .Z(n3825) );
  NAND U4830 ( .A(n3824), .B(n3825), .Z(n3826) );
  NANDN U4831 ( .A(n29456), .B(n3826), .Z(n3827) );
  NAND U4832 ( .A(n29457), .B(n3827), .Z(n29458) );
  NAND U4833 ( .A(n29476), .B(n29475), .Z(n3828) );
  NAND U4834 ( .A(n29477), .B(n3828), .Z(n3829) );
  ANDN U4835 ( .B(n3829), .A(n29478), .Z(n3830) );
  NANDN U4836 ( .A(n3830), .B(n29479), .Z(n3831) );
  NANDN U4837 ( .A(n23866), .B(n3831), .Z(n3832) );
  NAND U4838 ( .A(n23865), .B(n3832), .Z(n3833) );
  NANDN U4839 ( .A(n29480), .B(n3833), .Z(n3834) );
  NAND U4840 ( .A(n29481), .B(n3834), .Z(n3835) );
  ANDN U4841 ( .B(n3835), .A(n23864), .Z(n3836) );
  NANDN U4842 ( .A(n3836), .B(n23863), .Z(n3837) );
  AND U4843 ( .A(n29482), .B(n3837), .Z(n29484) );
  ANDN U4844 ( .B(n11275), .A(n29486), .Z(n3838) );
  NAND U4845 ( .A(n11212), .B(n29485), .Z(n3839) );
  AND U4846 ( .A(n3838), .B(n3839), .Z(n3840) );
  OR U4847 ( .A(n29488), .B(n3840), .Z(n3841) );
  NAND U4848 ( .A(n29489), .B(n3841), .Z(n3842) );
  NAND U4849 ( .A(n29490), .B(n3842), .Z(n3843) );
  ANDN U4850 ( .B(n11270), .A(n11271), .Z(n3844) );
  NAND U4851 ( .A(n3843), .B(n3844), .Z(n3845) );
  NAND U4852 ( .A(n29491), .B(n3845), .Z(n3846) );
  ANDN U4853 ( .B(n3846), .A(n11268), .Z(n3847) );
  XNOR U4854 ( .A(x[4060]), .B(y[4060]), .Z(n3848) );
  AND U4855 ( .A(n3847), .B(n3848), .Z(n3849) );
  ANDN U4856 ( .B(n23788), .A(n11265), .Z(n3850) );
  NANDN U4857 ( .A(n3849), .B(n29494), .Z(n3851) );
  AND U4858 ( .A(n3850), .B(n3851), .Z(n3852) );
  NANDN U4859 ( .A(n3852), .B(n29497), .Z(n3853) );
  NANDN U4860 ( .A(n29500), .B(n3853), .Z(n3854) );
  NAND U4861 ( .A(n29501), .B(n3854), .Z(n3855) );
  NANDN U4862 ( .A(n23860), .B(n3855), .Z(n11215) );
  AND U4863 ( .A(e), .B(n29531), .Z(n3856) );
  NAND U4864 ( .A(n29521), .B(n29520), .Z(n3857) );
  NAND U4865 ( .A(n29522), .B(n3857), .Z(n3858) );
  AND U4866 ( .A(n29523), .B(n3858), .Z(n3859) );
  ANDN U4867 ( .B(n23851), .A(n3859), .Z(n3860) );
  NAND U4868 ( .A(n23852), .B(n3860), .Z(n3861) );
  AND U4869 ( .A(n29524), .B(n3861), .Z(n3862) );
  NANDN U4870 ( .A(n3862), .B(n29525), .Z(n3863) );
  AND U4871 ( .A(n29526), .B(n3863), .Z(n3864) );
  OR U4872 ( .A(n29528), .B(n29527), .Z(n3865) );
  AND U4873 ( .A(n3864), .B(n3865), .Z(n3866) );
  NANDN U4874 ( .A(n29529), .B(n29530), .Z(n3867) );
  NANDN U4875 ( .A(n3866), .B(n23850), .Z(n3868) );
  NAND U4876 ( .A(n3867), .B(n3868), .Z(n3869) );
  NAND U4877 ( .A(n3869), .B(n3856), .Z(n3870) );
  NANDN U4878 ( .A(n3856), .B(g), .Z(n3871) );
  NAND U4879 ( .A(n3870), .B(n3871), .Z(n4) );
  IV U4880 ( .A(ebreg), .Z(e) );
  NANDN U4881 ( .A(x[4090]), .B(y[4090]), .Z(n3873) );
  NANDN U4882 ( .A(x[4089]), .B(y[4089]), .Z(n3872) );
  AND U4883 ( .A(n3873), .B(n3872), .Z(n3876) );
  NANDN U4884 ( .A(x[4092]), .B(y[4092]), .Z(n3875) );
  NANDN U4885 ( .A(x[4091]), .B(y[4091]), .Z(n3874) );
  NAND U4886 ( .A(n3875), .B(n3874), .Z(n29528) );
  ANDN U4887 ( .B(n3876), .A(n29528), .Z(n29525) );
  NANDN U4888 ( .A(x[4084]), .B(y[4084]), .Z(n3903) );
  NANDN U4889 ( .A(y[4095]), .B(x[4095]), .Z(n3878) );
  NANDN U4890 ( .A(y[4094]), .B(x[4094]), .Z(n3877) );
  AND U4891 ( .A(n3878), .B(n3877), .Z(n29529) );
  AND U4892 ( .A(n3903), .B(n29529), .Z(n3882) );
  NANDN U4893 ( .A(y[4090]), .B(x[4090]), .Z(n3880) );
  NANDN U4894 ( .A(y[4091]), .B(x[4091]), .Z(n3879) );
  AND U4895 ( .A(n3880), .B(n3879), .Z(n29527) );
  NANDN U4896 ( .A(x[4088]), .B(y[4088]), .Z(n23852) );
  AND U4897 ( .A(n29527), .B(n23852), .Z(n3881) );
  AND U4898 ( .A(n3882), .B(n3881), .Z(n3883) );
  AND U4899 ( .A(n29525), .B(n3883), .Z(n3902) );
  NANDN U4900 ( .A(y[4093]), .B(x[4093]), .Z(n3885) );
  NANDN U4901 ( .A(y[4092]), .B(x[4092]), .Z(n3884) );
  AND U4902 ( .A(n3885), .B(n3884), .Z(n29526) );
  NANDN U4903 ( .A(x[4086]), .B(y[4086]), .Z(n3887) );
  NANDN U4904 ( .A(x[4085]), .B(y[4085]), .Z(n3886) );
  AND U4905 ( .A(n3887), .B(n3886), .Z(n29522) );
  AND U4906 ( .A(n29526), .B(n29522), .Z(n3893) );
  NANDN U4907 ( .A(y[4089]), .B(x[4089]), .Z(n3889) );
  NANDN U4908 ( .A(y[4088]), .B(x[4088]), .Z(n3888) );
  AND U4909 ( .A(n3889), .B(n3888), .Z(n29524) );
  NANDN U4910 ( .A(y[4087]), .B(x[4087]), .Z(n3891) );
  NANDN U4911 ( .A(y[4086]), .B(x[4086]), .Z(n3890) );
  AND U4912 ( .A(n3891), .B(n3890), .Z(n29523) );
  AND U4913 ( .A(n29524), .B(n29523), .Z(n3892) );
  AND U4914 ( .A(n3893), .B(n3892), .Z(n3894) );
  NANDN U4915 ( .A(x[4087]), .B(y[4087]), .Z(n23851) );
  AND U4916 ( .A(n3894), .B(n23851), .Z(n3900) );
  NANDN U4917 ( .A(y[4084]), .B(x[4084]), .Z(n11244) );
  NANDN U4918 ( .A(y[4085]), .B(x[4085]), .Z(n3895) );
  AND U4919 ( .A(n11244), .B(n3895), .Z(n29521) );
  NANDN U4920 ( .A(x[4094]), .B(y[4094]), .Z(n3897) );
  NANDN U4921 ( .A(x[4093]), .B(y[4093]), .Z(n3896) );
  AND U4922 ( .A(n3897), .B(n3896), .Z(n3898) );
  NANDN U4923 ( .A(x[4095]), .B(y[4095]), .Z(n29530) );
  AND U4924 ( .A(n3898), .B(n29530), .Z(n23850) );
  AND U4925 ( .A(n29521), .B(n23850), .Z(n3899) );
  AND U4926 ( .A(n3900), .B(n3899), .Z(n3901) );
  AND U4927 ( .A(n3902), .B(n3901), .Z(n11242) );
  NANDN U4928 ( .A(x[4083]), .B(y[4083]), .Z(n11245) );
  AND U4929 ( .A(n11245), .B(n3903), .Z(n29519) );
  NANDN U4930 ( .A(y[4082]), .B(x[4082]), .Z(n23841) );
  NANDN U4931 ( .A(y[4083]), .B(x[4083]), .Z(n11243) );
  NAND U4932 ( .A(n23841), .B(n11243), .Z(n29518) );
  NANDN U4933 ( .A(x[4081]), .B(y[4081]), .Z(n11247) );
  NANDN U4934 ( .A(x[4082]), .B(y[4082]), .Z(n11246) );
  AND U4935 ( .A(n11247), .B(n11246), .Z(n23853) );
  XNOR U4936 ( .A(x[4078]), .B(y[4078]), .Z(n23829) );
  NANDN U4937 ( .A(y[4076]), .B(x[4076]), .Z(n3904) );
  NANDN U4938 ( .A(y[4077]), .B(x[4077]), .Z(n23830) );
  NAND U4939 ( .A(n3904), .B(n23830), .Z(n29513) );
  NANDN U4940 ( .A(x[4075]), .B(y[4075]), .Z(n23855) );
  XNOR U4941 ( .A(x[4076]), .B(y[4076]), .Z(n11252) );
  NANDN U4942 ( .A(x[4074]), .B(y[4074]), .Z(n11253) );
  ANDN U4943 ( .B(y[4073]), .A(x[4073]), .Z(n23818) );
  ANDN U4944 ( .B(n11253), .A(n23818), .Z(n29510) );
  XNOR U4945 ( .A(x[4072]), .B(y[4072]), .Z(n11257) );
  NANDN U4946 ( .A(y[4070]), .B(x[4070]), .Z(n3905) );
  NANDN U4947 ( .A(y[4071]), .B(x[4071]), .Z(n11256) );
  NAND U4948 ( .A(n3905), .B(n11256), .Z(n29505) );
  XNOR U4949 ( .A(x[4070]), .B(y[4070]), .Z(n11260) );
  NANDN U4950 ( .A(x[4065]), .B(y[4065]), .Z(n11262) );
  NANDN U4951 ( .A(x[4066]), .B(y[4066]), .Z(n11261) );
  NAND U4952 ( .A(n11262), .B(n11261), .Z(n23860) );
  NANDN U4953 ( .A(y[4064]), .B(x[4064]), .Z(n23794) );
  ANDN U4954 ( .B(x[4065]), .A(y[4065]), .Z(n23802) );
  ANDN U4955 ( .B(n23794), .A(n23802), .Z(n29501) );
  ANDN U4956 ( .B(y[4059]), .A(x[4059]), .Z(n11268) );
  NANDN U4957 ( .A(y[4058]), .B(x[4058]), .Z(n3906) );
  NANDN U4958 ( .A(y[4059]), .B(x[4059]), .Z(n11266) );
  AND U4959 ( .A(n3906), .B(n11266), .Z(n29491) );
  XNOR U4960 ( .A(x[4058]), .B(y[4058]), .Z(n11270) );
  ANDN U4961 ( .B(y[4057]), .A(x[4057]), .Z(n11271) );
  ANDN U4962 ( .B(y[4055]), .A(x[4055]), .Z(n23772) );
  ANDN U4963 ( .B(y[4056]), .A(x[4056]), .Z(n23777) );
  NOR U4964 ( .A(n23772), .B(n23777), .Z(n29489) );
  NANDN U4965 ( .A(y[4054]), .B(x[4054]), .Z(n3907) );
  NANDN U4966 ( .A(y[4055]), .B(x[4055]), .Z(n11273) );
  NAND U4967 ( .A(n3907), .B(n11273), .Z(n29488) );
  XNOR U4968 ( .A(x[4054]), .B(y[4054]), .Z(n11275) );
  ANDN U4969 ( .B(y[4053]), .A(x[4053]), .Z(n29486) );
  ANDN U4970 ( .B(y[4051]), .A(x[4051]), .Z(n11276) );
  NANDN U4971 ( .A(x[4049]), .B(y[4049]), .Z(n11278) );
  NANDN U4972 ( .A(x[4050]), .B(y[4050]), .Z(n11277) );
  NAND U4973 ( .A(n11278), .B(n11277), .Z(n23864) );
  NANDN U4974 ( .A(y[4048]), .B(x[4048]), .Z(n23752) );
  NANDN U4975 ( .A(y[4049]), .B(x[4049]), .Z(n23759) );
  AND U4976 ( .A(n23752), .B(n23759), .Z(n29481) );
  ANDN U4977 ( .B(y[4045]), .A(x[4045]), .Z(n23742) );
  NANDN U4978 ( .A(x[4046]), .B(y[4046]), .Z(n11281) );
  NANDN U4979 ( .A(n23742), .B(n11281), .Z(n23866) );
  NANDN U4980 ( .A(y[4044]), .B(x[4044]), .Z(n23738) );
  NANDN U4981 ( .A(y[4045]), .B(x[4045]), .Z(n23747) );
  AND U4982 ( .A(n23738), .B(n23747), .Z(n29479) );
  NANDN U4983 ( .A(x[4039]), .B(y[4039]), .Z(n11286) );
  NANDN U4984 ( .A(x[4040]), .B(y[4040]), .Z(n11285) );
  NAND U4985 ( .A(n11286), .B(n11285), .Z(n23868) );
  NANDN U4986 ( .A(y[4038]), .B(x[4038]), .Z(n23719) );
  NANDN U4987 ( .A(y[4039]), .B(x[4039]), .Z(n23726) );
  AND U4988 ( .A(n23719), .B(n23726), .Z(n29473) );
  NANDN U4989 ( .A(x[4035]), .B(y[4035]), .Z(n11290) );
  NANDN U4990 ( .A(x[4036]), .B(y[4036]), .Z(n11289) );
  NAND U4991 ( .A(n11290), .B(n11289), .Z(n29471) );
  NANDN U4992 ( .A(y[4032]), .B(x[4032]), .Z(n11292) );
  NANDN U4993 ( .A(y[4033]), .B(x[4033]), .Z(n23708) );
  NAND U4994 ( .A(n11292), .B(n23708), .Z(n23871) );
  NANDN U4995 ( .A(x[4031]), .B(y[4031]), .Z(n23698) );
  NANDN U4996 ( .A(x[4032]), .B(y[4032]), .Z(n23705) );
  AND U4997 ( .A(n23698), .B(n23705), .Z(n29469) );
  NANDN U4998 ( .A(y[4026]), .B(x[4026]), .Z(n11300) );
  NANDN U4999 ( .A(y[4027]), .B(x[4027]), .Z(n11297) );
  NAND U5000 ( .A(n11300), .B(n11297), .Z(n23873) );
  NANDN U5001 ( .A(x[4025]), .B(y[4025]), .Z(n23682) );
  NANDN U5002 ( .A(x[4026]), .B(y[4026]), .Z(n11299) );
  AND U5003 ( .A(n23682), .B(n11299), .Z(n29463) );
  XNOR U5004 ( .A(x[4024]), .B(y[4024]), .Z(n11302) );
  NANDN U5005 ( .A(x[4023]), .B(y[4023]), .Z(n29460) );
  AND U5006 ( .A(n11302), .B(n29460), .Z(n11197) );
  NANDN U5007 ( .A(y[4020]), .B(x[4020]), .Z(n23669) );
  NANDN U5008 ( .A(y[4021]), .B(x[4021]), .Z(n11306) );
  NAND U5009 ( .A(n23669), .B(n11306), .Z(n23875) );
  NANDN U5010 ( .A(x[4019]), .B(y[4019]), .Z(n11307) );
  NANDN U5011 ( .A(x[4020]), .B(y[4020]), .Z(n23673) );
  AND U5012 ( .A(n11307), .B(n23673), .Z(n29457) );
  XNOR U5013 ( .A(x[4018]), .B(y[4018]), .Z(n23663) );
  NANDN U5014 ( .A(x[4017]), .B(y[4017]), .Z(n29454) );
  AND U5015 ( .A(n23663), .B(n29454), .Z(n11189) );
  NANDN U5016 ( .A(x[4016]), .B(y[4016]), .Z(n11308) );
  ANDN U5017 ( .B(y[4015]), .A(x[4015]), .Z(n23655) );
  ANDN U5018 ( .B(n11308), .A(n23655), .Z(n29452) );
  NANDN U5019 ( .A(y[4014]), .B(x[4014]), .Z(n3908) );
  NANDN U5020 ( .A(y[4015]), .B(x[4015]), .Z(n23658) );
  NAND U5021 ( .A(n3908), .B(n23658), .Z(n29451) );
  NANDN U5022 ( .A(x[4013]), .B(y[4013]), .Z(n29449) );
  XNOR U5023 ( .A(x[4014]), .B(y[4014]), .Z(n11310) );
  NANDN U5024 ( .A(y[4012]), .B(x[4012]), .Z(n11312) );
  NANDN U5025 ( .A(y[4013]), .B(x[4013]), .Z(n11309) );
  AND U5026 ( .A(n11312), .B(n11309), .Z(n29448) );
  NANDN U5027 ( .A(x[4011]), .B(y[4011]), .Z(n11314) );
  NANDN U5028 ( .A(x[4012]), .B(y[4012]), .Z(n11311) );
  NAND U5029 ( .A(n11314), .B(n11311), .Z(n29447) );
  NANDN U5030 ( .A(y[4010]), .B(x[4010]), .Z(n23641) );
  NANDN U5031 ( .A(y[4011]), .B(x[4011]), .Z(n11313) );
  AND U5032 ( .A(n23641), .B(n11313), .Z(n29446) );
  NANDN U5033 ( .A(x[4009]), .B(y[4009]), .Z(n11316) );
  NANDN U5034 ( .A(x[4010]), .B(y[4010]), .Z(n11315) );
  NAND U5035 ( .A(n11316), .B(n11315), .Z(n29445) );
  NANDN U5036 ( .A(y[4008]), .B(x[4008]), .Z(n3909) );
  NANDN U5037 ( .A(y[4009]), .B(x[4009]), .Z(n23642) );
  AND U5038 ( .A(n3909), .B(n23642), .Z(n29444) );
  NANDN U5039 ( .A(x[4005]), .B(y[4005]), .Z(n11319) );
  NANDN U5040 ( .A(x[4006]), .B(y[4006]), .Z(n11318) );
  NAND U5041 ( .A(n11319), .B(n11318), .Z(n23878) );
  NANDN U5042 ( .A(y[4004]), .B(x[4004]), .Z(n23623) );
  NANDN U5043 ( .A(y[4005]), .B(x[4005]), .Z(n23630) );
  AND U5044 ( .A(n23623), .B(n23630), .Z(n29441) );
  NANDN U5045 ( .A(y[4002]), .B(x[4002]), .Z(n23617) );
  NANDN U5046 ( .A(y[4003]), .B(x[4003]), .Z(n23624) );
  AND U5047 ( .A(n23617), .B(n23624), .Z(n29439) );
  NANDN U5048 ( .A(x[4001]), .B(y[4001]), .Z(n11323) );
  NANDN U5049 ( .A(x[4002]), .B(y[4002]), .Z(n11322) );
  NAND U5050 ( .A(n11323), .B(n11322), .Z(n29438) );
  NANDN U5051 ( .A(y[3998]), .B(x[3998]), .Z(n11325) );
  NANDN U5052 ( .A(y[3999]), .B(x[3999]), .Z(n23612) );
  NAND U5053 ( .A(n11325), .B(n23612), .Z(n29435) );
  NANDN U5054 ( .A(x[3998]), .B(y[3998]), .Z(n23608) );
  ANDN U5055 ( .B(y[3997]), .A(x[3997]), .Z(n23602) );
  ANDN U5056 ( .B(n23608), .A(n23602), .Z(n29434) );
  ANDN U5057 ( .B(y[3995]), .A(x[3995]), .Z(n23597) );
  ANDN U5058 ( .B(y[3996]), .A(x[3996]), .Z(n23603) );
  NOR U5059 ( .A(n23597), .B(n23603), .Z(n29431) );
  XNOR U5060 ( .A(x[3994]), .B(y[3994]), .Z(n11330) );
  XNOR U5061 ( .A(x[3992]), .B(y[3992]), .Z(n11333) );
  NANDN U5062 ( .A(y[3990]), .B(x[3990]), .Z(n3910) );
  NANDN U5063 ( .A(y[3991]), .B(x[3991]), .Z(n11332) );
  NAND U5064 ( .A(n3910), .B(n11332), .Z(n29426) );
  XNOR U5065 ( .A(x[3990]), .B(y[3990]), .Z(n23585) );
  ANDN U5066 ( .B(y[3989]), .A(x[3989]), .Z(n11334) );
  XNOR U5067 ( .A(x[3988]), .B(y[3988]), .Z(n23579) );
  NANDN U5068 ( .A(x[3987]), .B(y[3987]), .Z(n29423) );
  AND U5069 ( .A(n23579), .B(n29423), .Z(n11150) );
  NANDN U5070 ( .A(y[3984]), .B(x[3984]), .Z(n11338) );
  NANDN U5071 ( .A(y[3985]), .B(x[3985]), .Z(n23574) );
  NAND U5072 ( .A(n11338), .B(n23574), .Z(n23884) );
  NANDN U5073 ( .A(x[3983]), .B(y[3983]), .Z(n11340) );
  NANDN U5074 ( .A(x[3984]), .B(y[3984]), .Z(n11337) );
  AND U5075 ( .A(n11340), .B(n11337), .Z(n29417) );
  NANDN U5076 ( .A(x[3981]), .B(y[3981]), .Z(n11342) );
  NANDN U5077 ( .A(x[3982]), .B(y[3982]), .Z(n11341) );
  AND U5078 ( .A(n11342), .B(n11341), .Z(n29415) );
  ANDN U5079 ( .B(x[3981]), .A(y[3981]), .Z(n23563) );
  NANDN U5080 ( .A(y[3980]), .B(x[3980]), .Z(n23556) );
  NANDN U5081 ( .A(n23563), .B(n23556), .Z(n29414) );
  NANDN U5082 ( .A(y[3978]), .B(x[3978]), .Z(n23550) );
  NANDN U5083 ( .A(y[3979]), .B(x[3979]), .Z(n23557) );
  AND U5084 ( .A(n23550), .B(n23557), .Z(n29413) );
  NANDN U5085 ( .A(x[3977]), .B(y[3977]), .Z(n23547) );
  NANDN U5086 ( .A(x[3978]), .B(y[3978]), .Z(n11345) );
  NAND U5087 ( .A(n23547), .B(n11345), .Z(n29412) );
  NANDN U5088 ( .A(y[3976]), .B(x[3976]), .Z(n11346) );
  NANDN U5089 ( .A(y[3977]), .B(x[3977]), .Z(n23551) );
  AND U5090 ( .A(n11346), .B(n23551), .Z(n29411) );
  NANDN U5091 ( .A(x[3975]), .B(y[3975]), .Z(n23541) );
  NANDN U5092 ( .A(x[3976]), .B(y[3976]), .Z(n23548) );
  NAND U5093 ( .A(n23541), .B(n23548), .Z(n29410) );
  NANDN U5094 ( .A(y[3974]), .B(x[3974]), .Z(n11348) );
  NANDN U5095 ( .A(y[3975]), .B(x[3975]), .Z(n11347) );
  AND U5096 ( .A(n11348), .B(n11347), .Z(n29409) );
  NANDN U5097 ( .A(x[3971]), .B(y[3971]), .Z(n11352) );
  NANDN U5098 ( .A(x[3972]), .B(y[3972]), .Z(n23536) );
  NAND U5099 ( .A(n11352), .B(n23536), .Z(n23887) );
  NANDN U5100 ( .A(y[3970]), .B(x[3970]), .Z(n11354) );
  NANDN U5101 ( .A(y[3971]), .B(x[3971]), .Z(n11351) );
  AND U5102 ( .A(n11354), .B(n11351), .Z(n29404) );
  NANDN U5103 ( .A(y[3966]), .B(x[3966]), .Z(n11359) );
  ANDN U5104 ( .B(x[3967]), .A(y[3967]), .Z(n23522) );
  ANDN U5105 ( .B(n11359), .A(n23522), .Z(n29399) );
  NANDN U5106 ( .A(x[3965]), .B(y[3965]), .Z(n11360) );
  NANDN U5107 ( .A(x[3966]), .B(y[3966]), .Z(n11357) );
  NAND U5108 ( .A(n11360), .B(n11357), .Z(n29398) );
  NANDN U5109 ( .A(y[3964]), .B(x[3964]), .Z(n11362) );
  NANDN U5110 ( .A(y[3965]), .B(x[3965]), .Z(n11358) );
  AND U5111 ( .A(n11362), .B(n11358), .Z(n29397) );
  NANDN U5112 ( .A(x[3963]), .B(y[3963]), .Z(n23509) );
  NANDN U5113 ( .A(x[3964]), .B(y[3964]), .Z(n11361) );
  NAND U5114 ( .A(n23509), .B(n11361), .Z(n29396) );
  NANDN U5115 ( .A(y[3962]), .B(x[3962]), .Z(n11364) );
  NANDN U5116 ( .A(y[3963]), .B(x[3963]), .Z(n11363) );
  AND U5117 ( .A(n11364), .B(n11363), .Z(n29395) );
  NANDN U5118 ( .A(x[3961]), .B(y[3961]), .Z(n23503) );
  NANDN U5119 ( .A(x[3962]), .B(y[3962]), .Z(n23510) );
  NAND U5120 ( .A(n23503), .B(n23510), .Z(n29394) );
  NANDN U5121 ( .A(y[3958]), .B(x[3958]), .Z(n23494) );
  NANDN U5122 ( .A(y[3959]), .B(x[3959]), .Z(n23501) );
  NAND U5123 ( .A(n23494), .B(n23501), .Z(n29391) );
  NANDN U5124 ( .A(x[3957]), .B(y[3957]), .Z(n11368) );
  NANDN U5125 ( .A(x[3958]), .B(y[3958]), .Z(n11367) );
  AND U5126 ( .A(n11368), .B(n11367), .Z(n29390) );
  NANDN U5127 ( .A(y[3956]), .B(x[3956]), .Z(n23488) );
  NANDN U5128 ( .A(y[3957]), .B(x[3957]), .Z(n23495) );
  NAND U5129 ( .A(n23488), .B(n23495), .Z(n29389) );
  NANDN U5130 ( .A(x[3955]), .B(y[3955]), .Z(n11370) );
  NANDN U5131 ( .A(x[3956]), .B(y[3956]), .Z(n11369) );
  AND U5132 ( .A(n11370), .B(n11369), .Z(n29388) );
  NANDN U5133 ( .A(x[3953]), .B(y[3953]), .Z(n11374) );
  NANDN U5134 ( .A(x[3954]), .B(y[3954]), .Z(n11371) );
  AND U5135 ( .A(n11374), .B(n11371), .Z(n29386) );
  NANDN U5136 ( .A(y[3952]), .B(x[3952]), .Z(n23480) );
  NANDN U5137 ( .A(y[3953]), .B(x[3953]), .Z(n11373) );
  NAND U5138 ( .A(n23480), .B(n11373), .Z(n29385) );
  NANDN U5139 ( .A(x[3951]), .B(y[3951]), .Z(n11376) );
  NANDN U5140 ( .A(x[3952]), .B(y[3952]), .Z(n11375) );
  AND U5141 ( .A(n11376), .B(n11375), .Z(n29384) );
  ANDN U5142 ( .B(x[3951]), .A(y[3951]), .Z(n23478) );
  NANDN U5143 ( .A(y[3950]), .B(x[3950]), .Z(n23471) );
  NANDN U5144 ( .A(n23478), .B(n23471), .Z(n29383) );
  NANDN U5145 ( .A(x[3949]), .B(y[3949]), .Z(n11378) );
  NANDN U5146 ( .A(x[3950]), .B(y[3950]), .Z(n11377) );
  AND U5147 ( .A(n11378), .B(n11377), .Z(n29382) );
  NANDN U5148 ( .A(y[3948]), .B(x[3948]), .Z(n3911) );
  NANDN U5149 ( .A(y[3949]), .B(x[3949]), .Z(n23472) );
  NAND U5150 ( .A(n3911), .B(n23472), .Z(n29381) );
  XNOR U5151 ( .A(x[3948]), .B(y[3948]), .Z(n23466) );
  NANDN U5152 ( .A(y[3946]), .B(x[3946]), .Z(n23459) );
  NANDN U5153 ( .A(y[3947]), .B(x[3947]), .Z(n23465) );
  NAND U5154 ( .A(n23459), .B(n23465), .Z(n29380) );
  NANDN U5155 ( .A(x[3945]), .B(y[3945]), .Z(n11380) );
  NANDN U5156 ( .A(x[3946]), .B(y[3946]), .Z(n11379) );
  AND U5157 ( .A(n11380), .B(n11379), .Z(n29379) );
  NANDN U5158 ( .A(y[3942]), .B(x[3942]), .Z(n11382) );
  NANDN U5159 ( .A(y[3943]), .B(x[3943]), .Z(n23454) );
  NAND U5160 ( .A(n11382), .B(n23454), .Z(n29374) );
  NANDN U5161 ( .A(x[3941]), .B(y[3941]), .Z(n11384) );
  NANDN U5162 ( .A(x[3942]), .B(y[3942]), .Z(n23450) );
  AND U5163 ( .A(n11384), .B(n23450), .Z(n23891) );
  XNOR U5164 ( .A(x[3938]), .B(y[3938]), .Z(n11390) );
  XNOR U5165 ( .A(x[3936]), .B(y[3936]), .Z(n23434) );
  NANDN U5166 ( .A(y[3934]), .B(x[3934]), .Z(n23427) );
  NANDN U5167 ( .A(y[3935]), .B(x[3935]), .Z(n23433) );
  NAND U5168 ( .A(n23427), .B(n23433), .Z(n29368) );
  NANDN U5169 ( .A(x[3933]), .B(y[3933]), .Z(n23423) );
  NANDN U5170 ( .A(x[3934]), .B(y[3934]), .Z(n11391) );
  AND U5171 ( .A(n23423), .B(n11391), .Z(n29367) );
  NANDN U5172 ( .A(y[3930]), .B(x[3930]), .Z(n11396) );
  NANDN U5173 ( .A(y[3931]), .B(x[3931]), .Z(n11393) );
  NAND U5174 ( .A(n11396), .B(n11393), .Z(n29363) );
  NANDN U5175 ( .A(x[3929]), .B(y[3929]), .Z(n11398) );
  NANDN U5176 ( .A(x[3930]), .B(y[3930]), .Z(n11395) );
  AND U5177 ( .A(n11398), .B(n11395), .Z(n23895) );
  NANDN U5178 ( .A(x[3925]), .B(y[3925]), .Z(n11404) );
  NANDN U5179 ( .A(x[3926]), .B(y[3926]), .Z(n11400) );
  AND U5180 ( .A(n11404), .B(n11400), .Z(n29360) );
  NANDN U5181 ( .A(y[3924]), .B(x[3924]), .Z(n11406) );
  NANDN U5182 ( .A(y[3925]), .B(x[3925]), .Z(n11403) );
  NAND U5183 ( .A(n11406), .B(n11403), .Z(n29359) );
  NANDN U5184 ( .A(x[3923]), .B(y[3923]), .Z(n11408) );
  NANDN U5185 ( .A(x[3924]), .B(y[3924]), .Z(n11405) );
  AND U5186 ( .A(n11408), .B(n11405), .Z(n29358) );
  NANDN U5187 ( .A(y[3922]), .B(x[3922]), .Z(n3912) );
  NANDN U5188 ( .A(y[3923]), .B(x[3923]), .Z(n11407) );
  NAND U5189 ( .A(n3912), .B(n11407), .Z(n29357) );
  NANDN U5190 ( .A(x[3921]), .B(y[3921]), .Z(n29355) );
  XNOR U5191 ( .A(x[3922]), .B(y[3922]), .Z(n11410) );
  AND U5192 ( .A(n29355), .B(n11410), .Z(n11075) );
  NANDN U5193 ( .A(y[3920]), .B(x[3920]), .Z(n3913) );
  NANDN U5194 ( .A(y[3921]), .B(x[3921]), .Z(n11409) );
  NAND U5195 ( .A(n3913), .B(n11409), .Z(n29354) );
  XNOR U5196 ( .A(x[3920]), .B(y[3920]), .Z(n23394) );
  NANDN U5197 ( .A(y[3918]), .B(x[3918]), .Z(n23387) );
  NANDN U5198 ( .A(y[3919]), .B(x[3919]), .Z(n23393) );
  NAND U5199 ( .A(n23387), .B(n23393), .Z(n29350) );
  NANDN U5200 ( .A(x[3917]), .B(y[3917]), .Z(n11412) );
  NANDN U5201 ( .A(x[3918]), .B(y[3918]), .Z(n11411) );
  AND U5202 ( .A(n11412), .B(n11411), .Z(n29349) );
  NANDN U5203 ( .A(y[3916]), .B(x[3916]), .Z(n23381) );
  NANDN U5204 ( .A(y[3917]), .B(x[3917]), .Z(n23388) );
  NAND U5205 ( .A(n23381), .B(n23388), .Z(n29348) );
  NANDN U5206 ( .A(x[3915]), .B(y[3915]), .Z(n11414) );
  NANDN U5207 ( .A(x[3916]), .B(y[3916]), .Z(n11413) );
  AND U5208 ( .A(n11414), .B(n11413), .Z(n29347) );
  NANDN U5209 ( .A(x[3914]), .B(y[3914]), .Z(n11415) );
  ANDN U5210 ( .B(y[3913]), .A(x[3913]), .Z(n23374) );
  ANDN U5211 ( .B(n11415), .A(n23374), .Z(n29345) );
  NANDN U5212 ( .A(y[3912]), .B(x[3912]), .Z(n11418) );
  NANDN U5213 ( .A(y[3913]), .B(x[3913]), .Z(n11417) );
  NAND U5214 ( .A(n11418), .B(n11417), .Z(n29344) );
  ANDN U5215 ( .B(y[3911]), .A(x[3911]), .Z(n23369) );
  ANDN U5216 ( .B(y[3912]), .A(x[3912]), .Z(n23375) );
  NOR U5217 ( .A(n23369), .B(n23375), .Z(n29343) );
  NANDN U5218 ( .A(y[3910]), .B(x[3910]), .Z(n3914) );
  NANDN U5219 ( .A(y[3911]), .B(x[3911]), .Z(n11419) );
  NAND U5220 ( .A(n3914), .B(n11419), .Z(n29342) );
  XNOR U5221 ( .A(x[3910]), .B(y[3910]), .Z(n11421) );
  NANDN U5222 ( .A(x[3909]), .B(y[3909]), .Z(n29340) );
  AND U5223 ( .A(n11421), .B(n29340), .Z(n11061) );
  NANDN U5224 ( .A(x[3907]), .B(y[3907]), .Z(n23358) );
  NANDN U5225 ( .A(x[3908]), .B(y[3908]), .Z(n11422) );
  AND U5226 ( .A(n23358), .B(n11422), .Z(n29338) );
  NANDN U5227 ( .A(y[3906]), .B(x[3906]), .Z(n11425) );
  NANDN U5228 ( .A(y[3907]), .B(x[3907]), .Z(n11424) );
  NAND U5229 ( .A(n11425), .B(n11424), .Z(n29337) );
  NANDN U5230 ( .A(x[3905]), .B(y[3905]), .Z(n23352) );
  NANDN U5231 ( .A(x[3906]), .B(y[3906]), .Z(n23359) );
  AND U5232 ( .A(n23352), .B(n23359), .Z(n29336) );
  NANDN U5233 ( .A(y[3904]), .B(x[3904]), .Z(n11427) );
  NANDN U5234 ( .A(y[3905]), .B(x[3905]), .Z(n11426) );
  NAND U5235 ( .A(n11427), .B(n11426), .Z(n29335) );
  NANDN U5236 ( .A(x[3903]), .B(y[3903]), .Z(n23346) );
  NANDN U5237 ( .A(x[3904]), .B(y[3904]), .Z(n23353) );
  AND U5238 ( .A(n23346), .B(n23353), .Z(n29334) );
  NANDN U5239 ( .A(x[3901]), .B(y[3901]), .Z(n23340) );
  NANDN U5240 ( .A(x[3902]), .B(y[3902]), .Z(n23347) );
  AND U5241 ( .A(n23340), .B(n23347), .Z(n29331) );
  NANDN U5242 ( .A(y[3900]), .B(x[3900]), .Z(n11431) );
  NANDN U5243 ( .A(y[3901]), .B(x[3901]), .Z(n11430) );
  NAND U5244 ( .A(n11431), .B(n11430), .Z(n29330) );
  NANDN U5245 ( .A(x[3900]), .B(y[3900]), .Z(n23341) );
  ANDN U5246 ( .B(y[3899]), .A(x[3899]), .Z(n23336) );
  ANDN U5247 ( .B(n23341), .A(n23336), .Z(n29329) );
  NANDN U5248 ( .A(y[3898]), .B(x[3898]), .Z(n3915) );
  NANDN U5249 ( .A(y[3899]), .B(x[3899]), .Z(n11432) );
  NAND U5250 ( .A(n3915), .B(n11432), .Z(n29328) );
  NANDN U5251 ( .A(x[3897]), .B(y[3897]), .Z(n29327) );
  XNOR U5252 ( .A(x[3898]), .B(y[3898]), .Z(n23333) );
  AND U5253 ( .A(n29327), .B(n23333), .Z(n11048) );
  NANDN U5254 ( .A(y[3896]), .B(x[3896]), .Z(n3916) );
  NANDN U5255 ( .A(y[3897]), .B(x[3897]), .Z(n23332) );
  NAND U5256 ( .A(n3916), .B(n23332), .Z(n29326) );
  XNOR U5257 ( .A(x[3896]), .B(y[3896]), .Z(n23326) );
  NANDN U5258 ( .A(y[3894]), .B(x[3894]), .Z(n11434) );
  NANDN U5259 ( .A(y[3895]), .B(x[3895]), .Z(n23327) );
  AND U5260 ( .A(n11434), .B(n23327), .Z(n29323) );
  NANDN U5261 ( .A(x[3893]), .B(y[3893]), .Z(n11437) );
  NANDN U5262 ( .A(x[3894]), .B(y[3894]), .Z(n11433) );
  AND U5263 ( .A(n11437), .B(n11433), .Z(n23899) );
  XNOR U5264 ( .A(x[3890]), .B(y[3890]), .Z(n23312) );
  NANDN U5265 ( .A(y[3888]), .B(x[3888]), .Z(n11441) );
  NANDN U5266 ( .A(y[3889]), .B(x[3889]), .Z(n23311) );
  NAND U5267 ( .A(n11441), .B(n23311), .Z(n29316) );
  NANDN U5268 ( .A(x[3885]), .B(y[3885]), .Z(n23297) );
  NANDN U5269 ( .A(x[3886]), .B(y[3886]), .Z(n23304) );
  NAND U5270 ( .A(n23297), .B(n23304), .Z(n29313) );
  NANDN U5271 ( .A(y[3884]), .B(x[3884]), .Z(n11445) );
  NANDN U5272 ( .A(y[3885]), .B(x[3885]), .Z(n11444) );
  AND U5273 ( .A(n11445), .B(n11444), .Z(n23901) );
  NANDN U5274 ( .A(x[3879]), .B(y[3879]), .Z(n23282) );
  NANDN U5275 ( .A(x[3880]), .B(y[3880]), .Z(n11450) );
  AND U5276 ( .A(n23282), .B(n11450), .Z(n29310) );
  XNOR U5277 ( .A(x[3878]), .B(y[3878]), .Z(n23280) );
  NANDN U5278 ( .A(y[3876]), .B(x[3876]), .Z(n11455) );
  ANDN U5279 ( .B(x[3877]), .A(y[3877]), .Z(n23279) );
  ANDN U5280 ( .B(n11455), .A(n23279), .Z(n29305) );
  NANDN U5281 ( .A(y[3874]), .B(x[3874]), .Z(n11458) );
  NANDN U5282 ( .A(y[3875]), .B(x[3875]), .Z(n11454) );
  AND U5283 ( .A(n11458), .B(n11454), .Z(n29304) );
  NANDN U5284 ( .A(x[3873]), .B(y[3873]), .Z(n11460) );
  NANDN U5285 ( .A(x[3874]), .B(y[3874]), .Z(n11457) );
  NAND U5286 ( .A(n11460), .B(n11457), .Z(n29303) );
  NANDN U5287 ( .A(y[3872]), .B(x[3872]), .Z(n11462) );
  NANDN U5288 ( .A(y[3873]), .B(x[3873]), .Z(n11459) );
  AND U5289 ( .A(n11462), .B(n11459), .Z(n29302) );
  NANDN U5290 ( .A(x[3871]), .B(y[3871]), .Z(n23265) );
  NANDN U5291 ( .A(x[3872]), .B(y[3872]), .Z(n11461) );
  NAND U5292 ( .A(n23265), .B(n11461), .Z(n29301) );
  NANDN U5293 ( .A(y[3870]), .B(x[3870]), .Z(n11464) );
  NANDN U5294 ( .A(y[3871]), .B(x[3871]), .Z(n11463) );
  AND U5295 ( .A(n11464), .B(n11463), .Z(n29300) );
  ANDN U5296 ( .B(y[3870]), .A(x[3870]), .Z(n23263) );
  NANDN U5297 ( .A(x[3869]), .B(y[3869]), .Z(n23256) );
  NANDN U5298 ( .A(n23263), .B(n23256), .Z(n29299) );
  NANDN U5299 ( .A(y[3868]), .B(x[3868]), .Z(n11466) );
  NANDN U5300 ( .A(y[3869]), .B(x[3869]), .Z(n11465) );
  AND U5301 ( .A(n11466), .B(n11465), .Z(n29298) );
  NANDN U5302 ( .A(x[3867]), .B(y[3867]), .Z(n23250) );
  NANDN U5303 ( .A(x[3868]), .B(y[3868]), .Z(n23257) );
  AND U5304 ( .A(n23250), .B(n23257), .Z(n29297) );
  NANDN U5305 ( .A(y[3866]), .B(x[3866]), .Z(n11468) );
  NANDN U5306 ( .A(y[3867]), .B(x[3867]), .Z(n11467) );
  NAND U5307 ( .A(n11468), .B(n11467), .Z(n23906) );
  NANDN U5308 ( .A(x[3865]), .B(y[3865]), .Z(n23244) );
  NANDN U5309 ( .A(x[3866]), .B(y[3866]), .Z(n23251) );
  AND U5310 ( .A(n23244), .B(n23251), .Z(n29296) );
  NANDN U5311 ( .A(x[3863]), .B(y[3863]), .Z(n23238) );
  NANDN U5312 ( .A(x[3864]), .B(y[3864]), .Z(n23245) );
  AND U5313 ( .A(n23238), .B(n23245), .Z(n29294) );
  NANDN U5314 ( .A(x[3861]), .B(y[3861]), .Z(n11472) );
  NANDN U5315 ( .A(x[3862]), .B(y[3862]), .Z(n23239) );
  AND U5316 ( .A(n11472), .B(n23239), .Z(n29291) );
  NANDN U5317 ( .A(y[3860]), .B(x[3860]), .Z(n11474) );
  NANDN U5318 ( .A(y[3861]), .B(x[3861]), .Z(n23235) );
  NAND U5319 ( .A(n11474), .B(n23235), .Z(n29290) );
  NANDN U5320 ( .A(x[3859]), .B(y[3859]), .Z(n23227) );
  NANDN U5321 ( .A(x[3860]), .B(y[3860]), .Z(n11473) );
  AND U5322 ( .A(n23227), .B(n11473), .Z(n29289) );
  NANDN U5323 ( .A(y[3858]), .B(x[3858]), .Z(n3917) );
  NANDN U5324 ( .A(y[3859]), .B(x[3859]), .Z(n11475) );
  NAND U5325 ( .A(n3917), .B(n11475), .Z(n29288) );
  NANDN U5326 ( .A(x[3857]), .B(y[3857]), .Z(n23907) );
  XNOR U5327 ( .A(x[3858]), .B(y[3858]), .Z(n23225) );
  AND U5328 ( .A(n23907), .B(n23225), .Z(n11000) );
  ANDN U5329 ( .B(x[3857]), .A(y[3857]), .Z(n23224) );
  NANDN U5330 ( .A(y[3856]), .B(x[3856]), .Z(n23218) );
  NANDN U5331 ( .A(n23224), .B(n23218), .Z(n29287) );
  NANDN U5332 ( .A(x[3855]), .B(y[3855]), .Z(n11477) );
  NANDN U5333 ( .A(x[3856]), .B(y[3856]), .Z(n11476) );
  AND U5334 ( .A(n11477), .B(n11476), .Z(n29286) );
  NANDN U5335 ( .A(y[3854]), .B(x[3854]), .Z(n23212) );
  NANDN U5336 ( .A(y[3855]), .B(x[3855]), .Z(n23219) );
  NAND U5337 ( .A(n23212), .B(n23219), .Z(n29285) );
  NANDN U5338 ( .A(x[3853]), .B(y[3853]), .Z(n11479) );
  NANDN U5339 ( .A(x[3854]), .B(y[3854]), .Z(n11478) );
  AND U5340 ( .A(n11479), .B(n11478), .Z(n29284) );
  NANDN U5341 ( .A(y[3852]), .B(x[3852]), .Z(n3918) );
  NANDN U5342 ( .A(y[3853]), .B(x[3853]), .Z(n23213) );
  NAND U5343 ( .A(n3918), .B(n23213), .Z(n29283) );
  XNOR U5344 ( .A(x[3852]), .B(y[3852]), .Z(n23206) );
  ANDN U5345 ( .B(y[3851]), .A(x[3851]), .Z(n23909) );
  ANDN U5346 ( .B(n23206), .A(n23909), .Z(n10993) );
  NANDN U5347 ( .A(y[3850]), .B(x[3850]), .Z(n3919) );
  NANDN U5348 ( .A(y[3851]), .B(x[3851]), .Z(n23207) );
  NAND U5349 ( .A(n3919), .B(n23207), .Z(n29282) );
  XNOR U5350 ( .A(x[3850]), .B(y[3850]), .Z(n11481) );
  NANDN U5351 ( .A(y[3848]), .B(x[3848]), .Z(n11483) );
  NANDN U5352 ( .A(y[3849]), .B(x[3849]), .Z(n11480) );
  NAND U5353 ( .A(n11483), .B(n11480), .Z(n29279) );
  NANDN U5354 ( .A(x[3847]), .B(y[3847]), .Z(n11485) );
  NANDN U5355 ( .A(x[3848]), .B(y[3848]), .Z(n11482) );
  AND U5356 ( .A(n11485), .B(n11482), .Z(n29278) );
  NANDN U5357 ( .A(y[3846]), .B(x[3846]), .Z(n3920) );
  NANDN U5358 ( .A(y[3847]), .B(x[3847]), .Z(n11484) );
  NAND U5359 ( .A(n3920), .B(n11484), .Z(n29276) );
  NANDN U5360 ( .A(x[3845]), .B(y[3845]), .Z(n23911) );
  XNOR U5361 ( .A(x[3846]), .B(y[3846]), .Z(n23192) );
  AND U5362 ( .A(n23911), .B(n23192), .Z(n10985) );
  NANDN U5363 ( .A(y[3844]), .B(x[3844]), .Z(n3921) );
  NANDN U5364 ( .A(y[3845]), .B(x[3845]), .Z(n23191) );
  NAND U5365 ( .A(n3921), .B(n23191), .Z(n29275) );
  XNOR U5366 ( .A(x[3844]), .B(y[3844]), .Z(n11487) );
  NANDN U5367 ( .A(y[3842]), .B(x[3842]), .Z(n11488) );
  NANDN U5368 ( .A(y[3843]), .B(x[3843]), .Z(n11486) );
  NAND U5369 ( .A(n11488), .B(n11486), .Z(n29272) );
  NANDN U5370 ( .A(x[3841]), .B(y[3841]), .Z(n23179) );
  NANDN U5371 ( .A(x[3842]), .B(y[3842]), .Z(n23185) );
  AND U5372 ( .A(n23179), .B(n23185), .Z(n29271) );
  NANDN U5373 ( .A(y[3836]), .B(x[3836]), .Z(n3922) );
  NANDN U5374 ( .A(y[3837]), .B(x[3837]), .Z(n11495) );
  NAND U5375 ( .A(n3922), .B(n11495), .Z(n29269) );
  XNOR U5376 ( .A(x[3836]), .B(y[3836]), .Z(n23166) );
  NANDN U5377 ( .A(x[3835]), .B(y[3835]), .Z(n29266) );
  AND U5378 ( .A(n23166), .B(n29266), .Z(n10973) );
  XNOR U5379 ( .A(x[3832]), .B(y[3832]), .Z(n23156) );
  XNOR U5380 ( .A(x[3830]), .B(y[3830]), .Z(n23150) );
  NANDN U5381 ( .A(y[3828]), .B(x[3828]), .Z(n3923) );
  NANDN U5382 ( .A(y[3829]), .B(x[3829]), .Z(n23151) );
  AND U5383 ( .A(n3923), .B(n23151), .Z(n29258) );
  XNOR U5384 ( .A(x[3828]), .B(y[3828]), .Z(n11501) );
  NANDN U5385 ( .A(x[3827]), .B(y[3827]), .Z(n23920) );
  AND U5386 ( .A(n11501), .B(n23920), .Z(n10960) );
  NANDN U5387 ( .A(y[3826]), .B(x[3826]), .Z(n11503) );
  NANDN U5388 ( .A(y[3827]), .B(x[3827]), .Z(n11500) );
  NAND U5389 ( .A(n11503), .B(n11500), .Z(n29257) );
  NANDN U5390 ( .A(x[3825]), .B(y[3825]), .Z(n11505) );
  NANDN U5391 ( .A(x[3826]), .B(y[3826]), .Z(n11502) );
  AND U5392 ( .A(n11505), .B(n11502), .Z(n29256) );
  NANDN U5393 ( .A(x[3823]), .B(y[3823]), .Z(n11507) );
  NANDN U5394 ( .A(x[3824]), .B(y[3824]), .Z(n11506) );
  AND U5395 ( .A(n11507), .B(n11506), .Z(n29254) );
  NANDN U5396 ( .A(y[3822]), .B(x[3822]), .Z(n23129) );
  NANDN U5397 ( .A(y[3823]), .B(x[3823]), .Z(n23136) );
  NAND U5398 ( .A(n23129), .B(n23136), .Z(n29253) );
  NANDN U5399 ( .A(x[3821]), .B(y[3821]), .Z(n11509) );
  NANDN U5400 ( .A(x[3822]), .B(y[3822]), .Z(n11508) );
  AND U5401 ( .A(n11509), .B(n11508), .Z(n29252) );
  NANDN U5402 ( .A(y[3820]), .B(x[3820]), .Z(n3924) );
  NANDN U5403 ( .A(y[3821]), .B(x[3821]), .Z(n23130) );
  NAND U5404 ( .A(n3924), .B(n23130), .Z(n29250) );
  NANDN U5405 ( .A(x[3819]), .B(y[3819]), .Z(n29248) );
  XNOR U5406 ( .A(x[3820]), .B(y[3820]), .Z(n11511) );
  AND U5407 ( .A(n29248), .B(n11511), .Z(n10951) );
  NANDN U5408 ( .A(y[3818]), .B(x[3818]), .Z(n3925) );
  NANDN U5409 ( .A(y[3819]), .B(x[3819]), .Z(n11510) );
  NAND U5410 ( .A(n3925), .B(n11510), .Z(n29247) );
  XNOR U5411 ( .A(x[3818]), .B(y[3818]), .Z(n11513) );
  NANDN U5412 ( .A(y[3816]), .B(x[3816]), .Z(n11514) );
  NANDN U5413 ( .A(y[3817]), .B(x[3817]), .Z(n11512) );
  NAND U5414 ( .A(n11514), .B(n11512), .Z(n29244) );
  NANDN U5415 ( .A(x[3815]), .B(y[3815]), .Z(n23113) );
  NANDN U5416 ( .A(x[3816]), .B(y[3816]), .Z(n23119) );
  AND U5417 ( .A(n23113), .B(n23119), .Z(n29243) );
  NANDN U5418 ( .A(y[3814]), .B(x[3814]), .Z(n3926) );
  NANDN U5419 ( .A(y[3815]), .B(x[3815]), .Z(n11515) );
  NAND U5420 ( .A(n3926), .B(n11515), .Z(n29242) );
  XNOR U5421 ( .A(x[3814]), .B(y[3814]), .Z(n11517) );
  NANDN U5422 ( .A(x[3813]), .B(y[3813]), .Z(n29240) );
  AND U5423 ( .A(n11517), .B(n29240), .Z(n10943) );
  NANDN U5424 ( .A(y[3812]), .B(x[3812]), .Z(n3927) );
  NANDN U5425 ( .A(y[3813]), .B(x[3813]), .Z(n11516) );
  NAND U5426 ( .A(n3927), .B(n11516), .Z(n29239) );
  XNOR U5427 ( .A(x[3812]), .B(y[3812]), .Z(n23106) );
  NANDN U5428 ( .A(x[3811]), .B(y[3811]), .Z(n29237) );
  XNOR U5429 ( .A(x[3810]), .B(y[3810]), .Z(n23100) );
  NANDN U5430 ( .A(y[3808]), .B(x[3808]), .Z(n3928) );
  NANDN U5431 ( .A(y[3809]), .B(x[3809]), .Z(n23101) );
  NAND U5432 ( .A(n3928), .B(n23101), .Z(n23921) );
  XNOR U5433 ( .A(x[3808]), .B(y[3808]), .Z(n11519) );
  ANDN U5434 ( .B(y[3807]), .A(x[3807]), .Z(n11520) );
  XNOR U5435 ( .A(x[3806]), .B(y[3806]), .Z(n11522) );
  NANDN U5436 ( .A(x[3805]), .B(y[3805]), .Z(n29229) );
  AND U5437 ( .A(n11522), .B(n29229), .Z(n10929) );
  NANDN U5438 ( .A(x[3803]), .B(y[3803]), .Z(n11524) );
  NANDN U5439 ( .A(x[3804]), .B(y[3804]), .Z(n11523) );
  AND U5440 ( .A(n11524), .B(n11523), .Z(n29227) );
  NANDN U5441 ( .A(y[3802]), .B(x[3802]), .Z(n23079) );
  NANDN U5442 ( .A(y[3803]), .B(x[3803]), .Z(n23086) );
  NAND U5443 ( .A(n23079), .B(n23086), .Z(n29226) );
  NANDN U5444 ( .A(x[3801]), .B(y[3801]), .Z(n11526) );
  NANDN U5445 ( .A(x[3802]), .B(y[3802]), .Z(n11525) );
  AND U5446 ( .A(n11526), .B(n11525), .Z(n29225) );
  NANDN U5447 ( .A(y[3800]), .B(x[3800]), .Z(n23073) );
  NANDN U5448 ( .A(y[3801]), .B(x[3801]), .Z(n23080) );
  NAND U5449 ( .A(n23073), .B(n23080), .Z(n29224) );
  NANDN U5450 ( .A(x[3799]), .B(y[3799]), .Z(n23069) );
  NANDN U5451 ( .A(x[3800]), .B(y[3800]), .Z(n11527) );
  AND U5452 ( .A(n23069), .B(n11527), .Z(n29223) );
  NANDN U5453 ( .A(x[3798]), .B(y[3798]), .Z(n23070) );
  ANDN U5454 ( .B(y[3797]), .A(x[3797]), .Z(n23064) );
  ANDN U5455 ( .B(n23070), .A(n23064), .Z(n29221) );
  NANDN U5456 ( .A(y[3796]), .B(x[3796]), .Z(n11530) );
  NANDN U5457 ( .A(y[3797]), .B(x[3797]), .Z(n11529) );
  NAND U5458 ( .A(n11530), .B(n11529), .Z(n29220) );
  ANDN U5459 ( .B(y[3795]), .A(x[3795]), .Z(n23059) );
  ANDN U5460 ( .B(y[3796]), .A(x[3796]), .Z(n23065) );
  NOR U5461 ( .A(n23059), .B(n23065), .Z(n29219) );
  NANDN U5462 ( .A(y[3794]), .B(x[3794]), .Z(n3929) );
  NANDN U5463 ( .A(y[3795]), .B(x[3795]), .Z(n11531) );
  NAND U5464 ( .A(n3929), .B(n11531), .Z(n29218) );
  XNOR U5465 ( .A(x[3794]), .B(y[3794]), .Z(n11533) );
  ANDN U5466 ( .B(y[3793]), .A(x[3793]), .Z(n29217) );
  ANDN U5467 ( .B(n11533), .A(n29217), .Z(n10916) );
  NANDN U5468 ( .A(y[3792]), .B(x[3792]), .Z(n3930) );
  NANDN U5469 ( .A(y[3793]), .B(x[3793]), .Z(n11532) );
  NAND U5470 ( .A(n3930), .B(n11532), .Z(n29216) );
  XNOR U5471 ( .A(x[3792]), .B(y[3792]), .Z(n11535) );
  NANDN U5472 ( .A(y[3790]), .B(x[3790]), .Z(n23047) );
  NANDN U5473 ( .A(y[3791]), .B(x[3791]), .Z(n11534) );
  NAND U5474 ( .A(n23047), .B(n11534), .Z(n29211) );
  NANDN U5475 ( .A(x[3789]), .B(y[3789]), .Z(n11537) );
  NANDN U5476 ( .A(x[3790]), .B(y[3790]), .Z(n11536) );
  AND U5477 ( .A(n11537), .B(n11536), .Z(n29210) );
  NANDN U5478 ( .A(y[3788]), .B(x[3788]), .Z(n3931) );
  NANDN U5479 ( .A(y[3789]), .B(x[3789]), .Z(n23048) );
  NAND U5480 ( .A(n3931), .B(n23048), .Z(n29209) );
  XNOR U5481 ( .A(x[3788]), .B(y[3788]), .Z(n23041) );
  NANDN U5482 ( .A(x[3787]), .B(y[3787]), .Z(n29207) );
  AND U5483 ( .A(n23041), .B(n29207), .Z(n10908) );
  NANDN U5484 ( .A(x[3786]), .B(y[3786]), .Z(n11538) );
  ANDN U5485 ( .B(y[3785]), .A(x[3785]), .Z(n23031) );
  ANDN U5486 ( .B(n11538), .A(n23031), .Z(n29205) );
  NANDN U5487 ( .A(y[3784]), .B(x[3784]), .Z(n23027) );
  NANDN U5488 ( .A(y[3785]), .B(x[3785]), .Z(n23036) );
  NAND U5489 ( .A(n23027), .B(n23036), .Z(n29204) );
  NANDN U5490 ( .A(x[3783]), .B(y[3783]), .Z(n11539) );
  ANDN U5491 ( .B(y[3784]), .A(x[3784]), .Z(n23033) );
  ANDN U5492 ( .B(n11539), .A(n23033), .Z(n29203) );
  NANDN U5493 ( .A(y[3782]), .B(x[3782]), .Z(n23020) );
  NANDN U5494 ( .A(y[3783]), .B(x[3783]), .Z(n23029) );
  NAND U5495 ( .A(n23020), .B(n23029), .Z(n29202) );
  NANDN U5496 ( .A(x[3781]), .B(y[3781]), .Z(n11541) );
  NANDN U5497 ( .A(x[3782]), .B(y[3782]), .Z(n11540) );
  AND U5498 ( .A(n11541), .B(n11540), .Z(n29201) );
  XNOR U5499 ( .A(x[3780]), .B(y[3780]), .Z(n23015) );
  NANDN U5500 ( .A(y[3778]), .B(x[3778]), .Z(n23008) );
  NANDN U5501 ( .A(y[3779]), .B(x[3779]), .Z(n23014) );
  AND U5502 ( .A(n23008), .B(n23014), .Z(n29197) );
  NANDN U5503 ( .A(x[3777]), .B(y[3777]), .Z(n23005) );
  NANDN U5504 ( .A(x[3778]), .B(y[3778]), .Z(n11542) );
  AND U5505 ( .A(n23005), .B(n11542), .Z(n23925) );
  NANDN U5506 ( .A(y[3772]), .B(x[3772]), .Z(n11547) );
  NANDN U5507 ( .A(y[3773]), .B(x[3773]), .Z(n11546) );
  NAND U5508 ( .A(n11547), .B(n11546), .Z(n29192) );
  NANDN U5509 ( .A(x[3771]), .B(y[3771]), .Z(n11549) );
  NANDN U5510 ( .A(x[3772]), .B(y[3772]), .Z(n22994) );
  AND U5511 ( .A(n11549), .B(n22994), .Z(n23927) );
  NANDN U5512 ( .A(y[3768]), .B(x[3768]), .Z(n3932) );
  NANDN U5513 ( .A(y[3769]), .B(x[3769]), .Z(n11552) );
  NAND U5514 ( .A(n3932), .B(n11552), .Z(n29190) );
  XNOR U5515 ( .A(x[3768]), .B(y[3768]), .Z(n11553) );
  NANDN U5516 ( .A(y[3766]), .B(x[3766]), .Z(n11556) );
  NANDN U5517 ( .A(y[3767]), .B(x[3767]), .Z(n11554) );
  NAND U5518 ( .A(n11556), .B(n11554), .Z(n29186) );
  NANDN U5519 ( .A(x[3765]), .B(y[3765]), .Z(n22973) );
  NANDN U5520 ( .A(x[3766]), .B(y[3766]), .Z(n11555) );
  AND U5521 ( .A(n22973), .B(n11555), .Z(n23929) );
  NANDN U5522 ( .A(y[3762]), .B(x[3762]), .Z(n11560) );
  NANDN U5523 ( .A(y[3763]), .B(x[3763]), .Z(n11559) );
  NAND U5524 ( .A(n11560), .B(n11559), .Z(n29182) );
  NANDN U5525 ( .A(y[3760]), .B(x[3760]), .Z(n11562) );
  NANDN U5526 ( .A(y[3761]), .B(x[3761]), .Z(n11561) );
  AND U5527 ( .A(n11562), .B(n11561), .Z(n29181) );
  NANDN U5528 ( .A(x[3759]), .B(y[3759]), .Z(n22955) );
  NANDN U5529 ( .A(x[3760]), .B(y[3760]), .Z(n22962) );
  NAND U5530 ( .A(n22955), .B(n22962), .Z(n29180) );
  NANDN U5531 ( .A(y[3758]), .B(x[3758]), .Z(n11564) );
  NANDN U5532 ( .A(y[3759]), .B(x[3759]), .Z(n11563) );
  AND U5533 ( .A(n11564), .B(n11563), .Z(n23932) );
  NANDN U5534 ( .A(x[3753]), .B(y[3753]), .Z(n22937) );
  NANDN U5535 ( .A(x[3754]), .B(y[3754]), .Z(n22944) );
  NAND U5536 ( .A(n22937), .B(n22944), .Z(n29174) );
  NANDN U5537 ( .A(y[3752]), .B(x[3752]), .Z(n22934) );
  NANDN U5538 ( .A(y[3753]), .B(x[3753]), .Z(n11569) );
  AND U5539 ( .A(n22934), .B(n11569), .Z(n23934) );
  NANDN U5540 ( .A(x[3748]), .B(y[3748]), .Z(n11572) );
  ANDN U5541 ( .B(y[3747]), .A(x[3747]), .Z(n22920) );
  ANDN U5542 ( .B(n11572), .A(n22920), .Z(n29171) );
  XNOR U5543 ( .A(x[3746]), .B(y[3746]), .Z(n11574) );
  NANDN U5544 ( .A(y[3744]), .B(x[3744]), .Z(n11576) );
  NANDN U5545 ( .A(y[3745]), .B(x[3745]), .Z(n11573) );
  AND U5546 ( .A(n11576), .B(n11573), .Z(n29167) );
  NANDN U5547 ( .A(y[3742]), .B(x[3742]), .Z(n22906) );
  NANDN U5548 ( .A(y[3743]), .B(x[3743]), .Z(n11577) );
  AND U5549 ( .A(n22906), .B(n11577), .Z(n29165) );
  NANDN U5550 ( .A(x[3741]), .B(y[3741]), .Z(n11580) );
  NANDN U5551 ( .A(x[3742]), .B(y[3742]), .Z(n11579) );
  NAND U5552 ( .A(n11580), .B(n11579), .Z(n29164) );
  NANDN U5553 ( .A(y[3740]), .B(x[3740]), .Z(n22900) );
  NANDN U5554 ( .A(y[3741]), .B(x[3741]), .Z(n22907) );
  AND U5555 ( .A(n22900), .B(n22907), .Z(n29163) );
  NANDN U5556 ( .A(x[3739]), .B(y[3739]), .Z(n11582) );
  NANDN U5557 ( .A(x[3740]), .B(y[3740]), .Z(n11581) );
  NAND U5558 ( .A(n11582), .B(n11581), .Z(n29162) );
  NANDN U5559 ( .A(y[3738]), .B(x[3738]), .Z(n22894) );
  NANDN U5560 ( .A(y[3739]), .B(x[3739]), .Z(n22901) );
  AND U5561 ( .A(n22894), .B(n22901), .Z(n29161) );
  NANDN U5562 ( .A(x[3737]), .B(y[3737]), .Z(n22891) );
  NANDN U5563 ( .A(x[3738]), .B(y[3738]), .Z(n11583) );
  NAND U5564 ( .A(n22891), .B(n11583), .Z(n29160) );
  NANDN U5565 ( .A(x[3735]), .B(y[3735]), .Z(n22885) );
  NANDN U5566 ( .A(x[3736]), .B(y[3736]), .Z(n22892) );
  AND U5567 ( .A(n22885), .B(n22892), .Z(n29159) );
  NANDN U5568 ( .A(y[3734]), .B(x[3734]), .Z(n11586) );
  NANDN U5569 ( .A(y[3735]), .B(x[3735]), .Z(n11585) );
  NAND U5570 ( .A(n11586), .B(n11585), .Z(n29158) );
  NANDN U5571 ( .A(x[3733]), .B(y[3733]), .Z(n22879) );
  NANDN U5572 ( .A(x[3734]), .B(y[3734]), .Z(n22886) );
  AND U5573 ( .A(n22879), .B(n22886), .Z(n29157) );
  NANDN U5574 ( .A(y[3732]), .B(x[3732]), .Z(n11588) );
  NANDN U5575 ( .A(y[3733]), .B(x[3733]), .Z(n11587) );
  NAND U5576 ( .A(n11588), .B(n11587), .Z(n29156) );
  NANDN U5577 ( .A(x[3731]), .B(y[3731]), .Z(n22873) );
  NANDN U5578 ( .A(x[3732]), .B(y[3732]), .Z(n22880) );
  AND U5579 ( .A(n22873), .B(n22880), .Z(n29155) );
  NANDN U5580 ( .A(x[3729]), .B(y[3729]), .Z(n11592) );
  NANDN U5581 ( .A(x[3730]), .B(y[3730]), .Z(n22874) );
  AND U5582 ( .A(n11592), .B(n22874), .Z(n29153) );
  NANDN U5583 ( .A(y[3728]), .B(x[3728]), .Z(n11594) );
  NANDN U5584 ( .A(y[3729]), .B(x[3729]), .Z(n11591) );
  NAND U5585 ( .A(n11594), .B(n11591), .Z(n29152) );
  NANDN U5586 ( .A(x[3727]), .B(y[3727]), .Z(n22863) );
  NANDN U5587 ( .A(x[3728]), .B(y[3728]), .Z(n11593) );
  AND U5588 ( .A(n22863), .B(n11593), .Z(n29151) );
  NANDN U5589 ( .A(y[3726]), .B(x[3726]), .Z(n3933) );
  NANDN U5590 ( .A(y[3727]), .B(x[3727]), .Z(n11595) );
  NAND U5591 ( .A(n3933), .B(n11595), .Z(n29150) );
  XNOR U5592 ( .A(x[3726]), .B(y[3726]), .Z(n22860) );
  NANDN U5593 ( .A(x[3725]), .B(y[3725]), .Z(n29147) );
  AND U5594 ( .A(n22860), .B(n29147), .Z(n10838) );
  NANDN U5595 ( .A(x[3723]), .B(y[3723]), .Z(n11599) );
  NANDN U5596 ( .A(x[3724]), .B(y[3724]), .Z(n11596) );
  AND U5597 ( .A(n11599), .B(n11596), .Z(n29145) );
  NANDN U5598 ( .A(y[3722]), .B(x[3722]), .Z(n11601) );
  NANDN U5599 ( .A(y[3723]), .B(x[3723]), .Z(n11597) );
  NAND U5600 ( .A(n11601), .B(n11597), .Z(n29144) );
  NANDN U5601 ( .A(x[3721]), .B(y[3721]), .Z(n11603) );
  NANDN U5602 ( .A(x[3722]), .B(y[3722]), .Z(n11600) );
  AND U5603 ( .A(n11603), .B(n11600), .Z(n29143) );
  XNOR U5604 ( .A(x[3720]), .B(y[3720]), .Z(n22846) );
  NANDN U5605 ( .A(x[3719]), .B(y[3719]), .Z(n29140) );
  AND U5606 ( .A(n22846), .B(n29140), .Z(n10830) );
  NANDN U5607 ( .A(x[3717]), .B(y[3717]), .Z(n11605) );
  NANDN U5608 ( .A(x[3718]), .B(y[3718]), .Z(n11604) );
  AND U5609 ( .A(n11605), .B(n11604), .Z(n29138) );
  NANDN U5610 ( .A(y[3716]), .B(x[3716]), .Z(n11607) );
  NANDN U5611 ( .A(y[3717]), .B(x[3717]), .Z(n22841) );
  NAND U5612 ( .A(n11607), .B(n22841), .Z(n29137) );
  NANDN U5613 ( .A(x[3715]), .B(y[3715]), .Z(n11609) );
  NANDN U5614 ( .A(x[3716]), .B(y[3716]), .Z(n11606) );
  AND U5615 ( .A(n11609), .B(n11606), .Z(n23940) );
  NANDN U5616 ( .A(y[3710]), .B(x[3710]), .Z(n22817) );
  NANDN U5617 ( .A(y[3711]), .B(x[3711]), .Z(n22824) );
  NAND U5618 ( .A(n22817), .B(n22824), .Z(n29132) );
  NANDN U5619 ( .A(x[3709]), .B(y[3709]), .Z(n11615) );
  NANDN U5620 ( .A(x[3710]), .B(y[3710]), .Z(n11614) );
  AND U5621 ( .A(n11615), .B(n11614), .Z(n29131) );
  NANDN U5622 ( .A(y[3708]), .B(x[3708]), .Z(n22811) );
  NANDN U5623 ( .A(y[3709]), .B(x[3709]), .Z(n22818) );
  NAND U5624 ( .A(n22811), .B(n22818), .Z(n29130) );
  NANDN U5625 ( .A(x[3707]), .B(y[3707]), .Z(n11617) );
  NANDN U5626 ( .A(x[3708]), .B(y[3708]), .Z(n11616) );
  AND U5627 ( .A(n11617), .B(n11616), .Z(n29129) );
  NANDN U5628 ( .A(y[3706]), .B(x[3706]), .Z(n22805) );
  NANDN U5629 ( .A(y[3707]), .B(x[3707]), .Z(n22812) );
  NAND U5630 ( .A(n22805), .B(n22812), .Z(n29128) );
  XNOR U5631 ( .A(x[3704]), .B(y[3704]), .Z(n22800) );
  ANDN U5632 ( .B(y[3703]), .A(x[3703]), .Z(n11620) );
  ANDN U5633 ( .B(n22800), .A(n11620), .Z(n10812) );
  NANDN U5634 ( .A(x[3701]), .B(y[3701]), .Z(n11622) );
  NANDN U5635 ( .A(x[3702]), .B(y[3702]), .Z(n11621) );
  AND U5636 ( .A(n11622), .B(n11621), .Z(n29123) );
  NANDN U5637 ( .A(y[3700]), .B(x[3700]), .Z(n22787) );
  NANDN U5638 ( .A(y[3701]), .B(x[3701]), .Z(n22794) );
  NAND U5639 ( .A(n22787), .B(n22794), .Z(n29122) );
  NANDN U5640 ( .A(x[3699]), .B(y[3699]), .Z(n11624) );
  NANDN U5641 ( .A(x[3700]), .B(y[3700]), .Z(n11623) );
  AND U5642 ( .A(n11624), .B(n11623), .Z(n29121) );
  NANDN U5643 ( .A(y[3698]), .B(x[3698]), .Z(n22781) );
  NANDN U5644 ( .A(y[3699]), .B(x[3699]), .Z(n22788) );
  NAND U5645 ( .A(n22781), .B(n22788), .Z(n29120) );
  NANDN U5646 ( .A(x[3697]), .B(y[3697]), .Z(n11626) );
  NANDN U5647 ( .A(x[3698]), .B(y[3698]), .Z(n11625) );
  AND U5648 ( .A(n11626), .B(n11625), .Z(n29119) );
  XNOR U5649 ( .A(x[3696]), .B(y[3696]), .Z(n22776) );
  NANDN U5650 ( .A(y[3694]), .B(x[3694]), .Z(n11628) );
  NANDN U5651 ( .A(y[3695]), .B(x[3695]), .Z(n22775) );
  AND U5652 ( .A(n11628), .B(n22775), .Z(n29114) );
  NANDN U5653 ( .A(x[3694]), .B(y[3694]), .Z(n11627) );
  ANDN U5654 ( .B(y[3693]), .A(x[3693]), .Z(n22768) );
  ANDN U5655 ( .B(n11627), .A(n22768), .Z(n29113) );
  NANDN U5656 ( .A(x[3691]), .B(y[3691]), .Z(n22762) );
  ANDN U5657 ( .B(y[3692]), .A(x[3692]), .Z(n22769) );
  ANDN U5658 ( .B(n22762), .A(n22769), .Z(n29112) );
  NANDN U5659 ( .A(x[3689]), .B(y[3689]), .Z(n22756) );
  ANDN U5660 ( .B(y[3690]), .A(x[3690]), .Z(n22763) );
  ANDN U5661 ( .B(n22756), .A(n22763), .Z(n29110) );
  NANDN U5662 ( .A(y[3688]), .B(x[3688]), .Z(n11634) );
  NANDN U5663 ( .A(y[3689]), .B(x[3689]), .Z(n11633) );
  NAND U5664 ( .A(n11634), .B(n11633), .Z(n29109) );
  NANDN U5665 ( .A(x[3687]), .B(y[3687]), .Z(n11636) );
  NANDN U5666 ( .A(x[3688]), .B(y[3688]), .Z(n22757) );
  AND U5667 ( .A(n11636), .B(n22757), .Z(n23945) );
  NANDN U5668 ( .A(y[3684]), .B(x[3684]), .Z(n3934) );
  NANDN U5669 ( .A(y[3685]), .B(x[3685]), .Z(n11639) );
  NAND U5670 ( .A(n3934), .B(n11639), .Z(n29105) );
  NANDN U5671 ( .A(x[3683]), .B(y[3683]), .Z(n29103) );
  XNOR U5672 ( .A(x[3684]), .B(y[3684]), .Z(n22743) );
  NANDN U5673 ( .A(y[3682]), .B(x[3682]), .Z(n3935) );
  NANDN U5674 ( .A(y[3683]), .B(x[3683]), .Z(n22742) );
  NAND U5675 ( .A(n3935), .B(n22742), .Z(n29102) );
  XNOR U5676 ( .A(x[3682]), .B(y[3682]), .Z(n22737) );
  NANDN U5677 ( .A(x[3681]), .B(y[3681]), .Z(n23947) );
  AND U5678 ( .A(n22737), .B(n23947), .Z(n10786) );
  NANDN U5679 ( .A(y[3680]), .B(x[3680]), .Z(n22731) );
  NANDN U5680 ( .A(y[3681]), .B(x[3681]), .Z(n22738) );
  NAND U5681 ( .A(n22731), .B(n22738), .Z(n29101) );
  NANDN U5682 ( .A(x[3679]), .B(y[3679]), .Z(n11641) );
  NANDN U5683 ( .A(x[3680]), .B(y[3680]), .Z(n11640) );
  AND U5684 ( .A(n11641), .B(n11640), .Z(n29100) );
  NANDN U5685 ( .A(x[3677]), .B(y[3677]), .Z(n11643) );
  NANDN U5686 ( .A(x[3678]), .B(y[3678]), .Z(n11642) );
  AND U5687 ( .A(n11643), .B(n11642), .Z(n29098) );
  NANDN U5688 ( .A(y[3676]), .B(x[3676]), .Z(n11645) );
  NANDN U5689 ( .A(y[3677]), .B(x[3677]), .Z(n22726) );
  NAND U5690 ( .A(n11645), .B(n22726), .Z(n29097) );
  NANDN U5691 ( .A(x[3676]), .B(y[3676]), .Z(n11644) );
  ANDN U5692 ( .B(y[3675]), .A(x[3675]), .Z(n22719) );
  ANDN U5693 ( .B(n11644), .A(n22719), .Z(n29096) );
  NANDN U5694 ( .A(y[3674]), .B(x[3674]), .Z(n3936) );
  NANDN U5695 ( .A(y[3675]), .B(x[3675]), .Z(n11646) );
  NAND U5696 ( .A(n3936), .B(n11646), .Z(n29095) );
  XNOR U5697 ( .A(x[3674]), .B(y[3674]), .Z(n22714) );
  ANDN U5698 ( .B(y[3673]), .A(x[3673]), .Z(n29093) );
  ANDN U5699 ( .B(n22714), .A(n29093), .Z(n10777) );
  NANDN U5700 ( .A(y[3672]), .B(x[3672]), .Z(n11647) );
  NANDN U5701 ( .A(y[3673]), .B(x[3673]), .Z(n22715) );
  NAND U5702 ( .A(n11647), .B(n22715), .Z(n29092) );
  ANDN U5703 ( .B(y[3671]), .A(x[3671]), .Z(n22706) );
  ANDN U5704 ( .B(y[3672]), .A(x[3672]), .Z(n22712) );
  NOR U5705 ( .A(n22706), .B(n22712), .Z(n29091) );
  NANDN U5706 ( .A(y[3670]), .B(x[3670]), .Z(n3937) );
  NANDN U5707 ( .A(y[3671]), .B(x[3671]), .Z(n11648) );
  NAND U5708 ( .A(n3937), .B(n11648), .Z(n29090) );
  XNOR U5709 ( .A(x[3670]), .B(y[3670]), .Z(n11650) );
  ANDN U5710 ( .B(y[3669]), .A(x[3669]), .Z(n22700) );
  XNOR U5711 ( .A(x[3668]), .B(y[3668]), .Z(n11652) );
  NANDN U5712 ( .A(x[3667]), .B(y[3667]), .Z(n29086) );
  AND U5713 ( .A(n11652), .B(n29086), .Z(n10768) );
  ANDN U5714 ( .B(x[3664]), .A(y[3664]), .Z(n22689) );
  ANDN U5715 ( .B(x[3665]), .A(y[3665]), .Z(n22693) );
  OR U5716 ( .A(n22689), .B(n22693), .Z(n29083) );
  NANDN U5717 ( .A(y[3662]), .B(x[3662]), .Z(n3938) );
  ANDN U5718 ( .B(x[3663]), .A(y[3663]), .Z(n11655) );
  ANDN U5719 ( .B(n3938), .A(n11655), .Z(n29081) );
  NANDN U5720 ( .A(x[3661]), .B(y[3661]), .Z(n22681) );
  NANDN U5721 ( .A(x[3662]), .B(y[3662]), .Z(n11654) );
  NAND U5722 ( .A(n22681), .B(n11654), .Z(n29080) );
  NANDN U5723 ( .A(y[3660]), .B(x[3660]), .Z(n11659) );
  NANDN U5724 ( .A(y[3661]), .B(x[3661]), .Z(n11658) );
  AND U5725 ( .A(n11659), .B(n11658), .Z(n23952) );
  NANDN U5726 ( .A(x[3657]), .B(y[3657]), .Z(n22669) );
  NANDN U5727 ( .A(x[3658]), .B(y[3658]), .Z(n22676) );
  NAND U5728 ( .A(n22669), .B(n22676), .Z(n23954) );
  NANDN U5729 ( .A(x[3655]), .B(y[3655]), .Z(n22663) );
  NANDN U5730 ( .A(x[3656]), .B(y[3656]), .Z(n22670) );
  AND U5731 ( .A(n22663), .B(n22670), .Z(n29075) );
  NANDN U5732 ( .A(y[3654]), .B(x[3654]), .Z(n11665) );
  NANDN U5733 ( .A(y[3655]), .B(x[3655]), .Z(n11664) );
  NAND U5734 ( .A(n11665), .B(n11664), .Z(n29074) );
  NANDN U5735 ( .A(x[3653]), .B(y[3653]), .Z(n22657) );
  NANDN U5736 ( .A(x[3654]), .B(y[3654]), .Z(n22664) );
  AND U5737 ( .A(n22657), .B(n22664), .Z(n29073) );
  NANDN U5738 ( .A(y[3652]), .B(x[3652]), .Z(n3939) );
  NANDN U5739 ( .A(y[3653]), .B(x[3653]), .Z(n11666) );
  NAND U5740 ( .A(n3939), .B(n11666), .Z(n29072) );
  XNOR U5741 ( .A(x[3652]), .B(y[3652]), .Z(n22655) );
  ANDN U5742 ( .B(x[3651]), .A(y[3651]), .Z(n22654) );
  NANDN U5743 ( .A(y[3650]), .B(x[3650]), .Z(n11669) );
  NANDN U5744 ( .A(n22654), .B(n11669), .Z(n29071) );
  NANDN U5745 ( .A(x[3645]), .B(y[3645]), .Z(n22635) );
  NANDN U5746 ( .A(x[3646]), .B(y[3646]), .Z(n22642) );
  NAND U5747 ( .A(n22635), .B(n22642), .Z(n29066) );
  NANDN U5748 ( .A(y[3644]), .B(x[3644]), .Z(n11676) );
  NANDN U5749 ( .A(y[3645]), .B(x[3645]), .Z(n11675) );
  AND U5750 ( .A(n11676), .B(n11675), .Z(n23959) );
  NANDN U5751 ( .A(x[3641]), .B(y[3641]), .Z(n22623) );
  NANDN U5752 ( .A(x[3642]), .B(y[3642]), .Z(n22630) );
  NAND U5753 ( .A(n22623), .B(n22630), .Z(n29064) );
  NANDN U5754 ( .A(x[3639]), .B(y[3639]), .Z(n22617) );
  NANDN U5755 ( .A(x[3640]), .B(y[3640]), .Z(n22624) );
  AND U5756 ( .A(n22617), .B(n22624), .Z(n29062) );
  NANDN U5757 ( .A(y[3638]), .B(x[3638]), .Z(n22613) );
  NANDN U5758 ( .A(y[3639]), .B(x[3639]), .Z(n11681) );
  NAND U5759 ( .A(n22613), .B(n11681), .Z(n29061) );
  NANDN U5760 ( .A(x[3637]), .B(y[3637]), .Z(n22610) );
  NANDN U5761 ( .A(x[3638]), .B(y[3638]), .Z(n22618) );
  AND U5762 ( .A(n22610), .B(n22618), .Z(n29060) );
  NANDN U5763 ( .A(y[3636]), .B(x[3636]), .Z(n11682) );
  NANDN U5764 ( .A(y[3637]), .B(x[3637]), .Z(n22614) );
  NAND U5765 ( .A(n11682), .B(n22614), .Z(n29059) );
  NANDN U5766 ( .A(x[3635]), .B(y[3635]), .Z(n11684) );
  NANDN U5767 ( .A(x[3636]), .B(y[3636]), .Z(n22612) );
  AND U5768 ( .A(n11684), .B(n22612), .Z(n29058) );
  XNOR U5769 ( .A(x[3634]), .B(y[3634]), .Z(n22602) );
  XNOR U5770 ( .A(x[3632]), .B(y[3632]), .Z(n22596) );
  NANDN U5771 ( .A(y[3630]), .B(x[3630]), .Z(n11686) );
  NANDN U5772 ( .A(y[3631]), .B(x[3631]), .Z(n22597) );
  NAND U5773 ( .A(n11686), .B(n22597), .Z(n29049) );
  NANDN U5774 ( .A(x[3629]), .B(y[3629]), .Z(n11688) );
  NANDN U5775 ( .A(x[3630]), .B(y[3630]), .Z(n11685) );
  AND U5776 ( .A(n11688), .B(n11685), .Z(n29048) );
  NANDN U5777 ( .A(y[3628]), .B(x[3628]), .Z(n3940) );
  NANDN U5778 ( .A(y[3629]), .B(x[3629]), .Z(n11687) );
  NAND U5779 ( .A(n3940), .B(n11687), .Z(n29047) );
  XNOR U5780 ( .A(x[3628]), .B(y[3628]), .Z(n11690) );
  NANDN U5781 ( .A(x[3627]), .B(y[3627]), .Z(n29045) );
  AND U5782 ( .A(n11690), .B(n29045), .Z(n10720) );
  NANDN U5783 ( .A(x[3626]), .B(y[3626]), .Z(n11691) );
  ANDN U5784 ( .B(y[3625]), .A(x[3625]), .Z(n22580) );
  ANDN U5785 ( .B(n11691), .A(n22580), .Z(n29043) );
  NANDN U5786 ( .A(y[3624]), .B(x[3624]), .Z(n11694) );
  NANDN U5787 ( .A(y[3625]), .B(x[3625]), .Z(n11693) );
  NAND U5788 ( .A(n11694), .B(n11693), .Z(n29042) );
  ANDN U5789 ( .B(y[3623]), .A(x[3623]), .Z(n22575) );
  ANDN U5790 ( .B(y[3624]), .A(x[3624]), .Z(n22581) );
  NOR U5791 ( .A(n22575), .B(n22581), .Z(n29041) );
  NANDN U5792 ( .A(y[3622]), .B(x[3622]), .Z(n3941) );
  NANDN U5793 ( .A(y[3623]), .B(x[3623]), .Z(n11695) );
  NAND U5794 ( .A(n3941), .B(n11695), .Z(n29040) );
  XNOR U5795 ( .A(x[3622]), .B(y[3622]), .Z(n11697) );
  ANDN U5796 ( .B(y[3621]), .A(x[3621]), .Z(n29038) );
  ANDN U5797 ( .B(n11697), .A(n29038), .Z(n10713) );
  NANDN U5798 ( .A(y[3620]), .B(x[3620]), .Z(n3942) );
  NANDN U5799 ( .A(y[3621]), .B(x[3621]), .Z(n11696) );
  NAND U5800 ( .A(n3942), .B(n11696), .Z(n29037) );
  XNOR U5801 ( .A(x[3620]), .B(y[3620]), .Z(n11699) );
  NANDN U5802 ( .A(y[3618]), .B(x[3618]), .Z(n11701) );
  NANDN U5803 ( .A(y[3619]), .B(x[3619]), .Z(n11698) );
  NAND U5804 ( .A(n11701), .B(n11698), .Z(n29035) );
  NANDN U5805 ( .A(x[3617]), .B(y[3617]), .Z(n11703) );
  NANDN U5806 ( .A(x[3618]), .B(y[3618]), .Z(n11700) );
  AND U5807 ( .A(n11703), .B(n11700), .Z(n29034) );
  NANDN U5808 ( .A(y[3616]), .B(x[3616]), .Z(n11705) );
  NANDN U5809 ( .A(y[3617]), .B(x[3617]), .Z(n11702) );
  NAND U5810 ( .A(n11705), .B(n11702), .Z(n29032) );
  NANDN U5811 ( .A(x[3615]), .B(y[3615]), .Z(n11707) );
  NANDN U5812 ( .A(x[3616]), .B(y[3616]), .Z(n11704) );
  AND U5813 ( .A(n11707), .B(n11704), .Z(n29031) );
  NANDN U5814 ( .A(x[3613]), .B(y[3613]), .Z(n11711) );
  NANDN U5815 ( .A(x[3614]), .B(y[3614]), .Z(n11708) );
  AND U5816 ( .A(n11711), .B(n11708), .Z(n29029) );
  NANDN U5817 ( .A(y[3612]), .B(x[3612]), .Z(n22551) );
  NANDN U5818 ( .A(y[3613]), .B(x[3613]), .Z(n11710) );
  NAND U5819 ( .A(n22551), .B(n11710), .Z(n29028) );
  NANDN U5820 ( .A(x[3611]), .B(y[3611]), .Z(n11713) );
  NANDN U5821 ( .A(x[3612]), .B(y[3612]), .Z(n11712) );
  AND U5822 ( .A(n11713), .B(n11712), .Z(n29027) );
  ANDN U5823 ( .B(x[3611]), .A(y[3611]), .Z(n22553) );
  NANDN U5824 ( .A(y[3610]), .B(x[3610]), .Z(n3943) );
  NANDN U5825 ( .A(n22553), .B(n3943), .Z(n29026) );
  XNOR U5826 ( .A(x[3610]), .B(y[3610]), .Z(n22545) );
  NANDN U5827 ( .A(x[3609]), .B(y[3609]), .Z(n29024) );
  AND U5828 ( .A(n22545), .B(n29024), .Z(n10699) );
  XNOR U5829 ( .A(x[3608]), .B(y[3608]), .Z(n11715) );
  XNOR U5830 ( .A(x[3606]), .B(y[3606]), .Z(n11717) );
  NANDN U5831 ( .A(y[3604]), .B(x[3604]), .Z(n3944) );
  NANDN U5832 ( .A(y[3605]), .B(x[3605]), .Z(n11716) );
  NAND U5833 ( .A(n3944), .B(n11716), .Z(n29018) );
  XNOR U5834 ( .A(x[3604]), .B(y[3604]), .Z(n11719) );
  ANDN U5835 ( .B(y[3603]), .A(x[3603]), .Z(n29015) );
  ANDN U5836 ( .B(n11719), .A(n29015), .Z(n10688) );
  NANDN U5837 ( .A(y[3602]), .B(x[3602]), .Z(n11720) );
  NANDN U5838 ( .A(y[3603]), .B(x[3603]), .Z(n11718) );
  NAND U5839 ( .A(n11720), .B(n11718), .Z(n29014) );
  NANDN U5840 ( .A(x[3601]), .B(y[3601]), .Z(n22524) );
  ANDN U5841 ( .B(y[3602]), .A(x[3602]), .Z(n22530) );
  ANDN U5842 ( .B(n22524), .A(n22530), .Z(n29013) );
  XNOR U5843 ( .A(x[3600]), .B(y[3600]), .Z(n11723) );
  NANDN U5844 ( .A(y[3598]), .B(x[3598]), .Z(n11724) );
  NANDN U5845 ( .A(y[3599]), .B(x[3599]), .Z(n11722) );
  NAND U5846 ( .A(n11724), .B(n11722), .Z(n29011) );
  NANDN U5847 ( .A(x[3595]), .B(y[3595]), .Z(n22507) );
  NANDN U5848 ( .A(x[3596]), .B(y[3596]), .Z(n22514) );
  NAND U5849 ( .A(n22507), .B(n22514), .Z(n23967) );
  NANDN U5850 ( .A(y[3594]), .B(x[3594]), .Z(n11728) );
  NANDN U5851 ( .A(y[3595]), .B(x[3595]), .Z(n11727) );
  AND U5852 ( .A(n11728), .B(n11727), .Z(n29009) );
  NANDN U5853 ( .A(x[3591]), .B(y[3591]), .Z(n22495) );
  NANDN U5854 ( .A(x[3592]), .B(y[3592]), .Z(n22502) );
  NAND U5855 ( .A(n22495), .B(n22502), .Z(n23969) );
  NANDN U5856 ( .A(x[3589]), .B(y[3589]), .Z(n22489) );
  NANDN U5857 ( .A(x[3590]), .B(y[3590]), .Z(n22496) );
  AND U5858 ( .A(n22489), .B(n22496), .Z(n29004) );
  NANDN U5859 ( .A(y[3588]), .B(x[3588]), .Z(n11734) );
  NANDN U5860 ( .A(y[3589]), .B(x[3589]), .Z(n11733) );
  NAND U5861 ( .A(n11734), .B(n11733), .Z(n29003) );
  NANDN U5862 ( .A(x[3587]), .B(y[3587]), .Z(n22483) );
  NANDN U5863 ( .A(x[3588]), .B(y[3588]), .Z(n22490) );
  AND U5864 ( .A(n22483), .B(n22490), .Z(n29002) );
  NANDN U5865 ( .A(y[3586]), .B(x[3586]), .Z(n22479) );
  NANDN U5866 ( .A(y[3587]), .B(x[3587]), .Z(n11735) );
  NAND U5867 ( .A(n22479), .B(n11735), .Z(n29001) );
  NANDN U5868 ( .A(x[3585]), .B(y[3585]), .Z(n22478) );
  NANDN U5869 ( .A(x[3586]), .B(y[3586]), .Z(n22484) );
  AND U5870 ( .A(n22478), .B(n22484), .Z(n29000) );
  NANDN U5871 ( .A(x[3583]), .B(y[3583]), .Z(n22469) );
  ANDN U5872 ( .B(y[3584]), .A(x[3584]), .Z(n22476) );
  ANDN U5873 ( .B(n22469), .A(n22476), .Z(n28998) );
  NANDN U5874 ( .A(y[3582]), .B(x[3582]), .Z(n11738) );
  NANDN U5875 ( .A(y[3583]), .B(x[3583]), .Z(n11737) );
  NAND U5876 ( .A(n11738), .B(n11737), .Z(n28997) );
  NANDN U5877 ( .A(x[3581]), .B(y[3581]), .Z(n22463) );
  NANDN U5878 ( .A(x[3582]), .B(y[3582]), .Z(n22470) );
  AND U5879 ( .A(n22463), .B(n22470), .Z(n28996) );
  NANDN U5880 ( .A(y[3580]), .B(x[3580]), .Z(n11740) );
  NANDN U5881 ( .A(y[3581]), .B(x[3581]), .Z(n11739) );
  NAND U5882 ( .A(n11740), .B(n11739), .Z(n28995) );
  NANDN U5883 ( .A(x[3579]), .B(y[3579]), .Z(n22457) );
  NANDN U5884 ( .A(x[3580]), .B(y[3580]), .Z(n22464) );
  AND U5885 ( .A(n22457), .B(n22464), .Z(n28994) );
  NANDN U5886 ( .A(y[3578]), .B(x[3578]), .Z(n22453) );
  NANDN U5887 ( .A(y[3579]), .B(x[3579]), .Z(n11741) );
  NAND U5888 ( .A(n22453), .B(n11741), .Z(n28993) );
  NANDN U5889 ( .A(y[3577]), .B(x[3577]), .Z(n22454) );
  ANDN U5890 ( .B(x[3576]), .A(y[3576]), .Z(n22448) );
  ANDN U5891 ( .B(n22454), .A(n22448), .Z(n28991) );
  NANDN U5892 ( .A(x[3575]), .B(y[3575]), .Z(n22446) );
  NANDN U5893 ( .A(x[3576]), .B(y[3576]), .Z(n22452) );
  NAND U5894 ( .A(n22446), .B(n22452), .Z(n28990) );
  NANDN U5895 ( .A(y[3575]), .B(x[3575]), .Z(n3946) );
  NANDN U5896 ( .A(y[3574]), .B(x[3574]), .Z(n3945) );
  AND U5897 ( .A(n3946), .B(n3945), .Z(n28989) );
  ANDN U5898 ( .B(y[3572]), .A(x[3572]), .Z(n11743) );
  NANDN U5899 ( .A(x[3571]), .B(y[3571]), .Z(n11744) );
  NANDN U5900 ( .A(n11743), .B(n11744), .Z(n28985) );
  NANDN U5901 ( .A(y[3570]), .B(x[3570]), .Z(n22432) );
  ANDN U5902 ( .B(x[3571]), .A(y[3571]), .Z(n22440) );
  ANDN U5903 ( .B(n22432), .A(n22440), .Z(n28984) );
  NANDN U5904 ( .A(x[3569]), .B(y[3569]), .Z(n11746) );
  NANDN U5905 ( .A(x[3570]), .B(y[3570]), .Z(n11745) );
  NAND U5906 ( .A(n11746), .B(n11745), .Z(n28983) );
  NANDN U5907 ( .A(y[3568]), .B(x[3568]), .Z(n22426) );
  NANDN U5908 ( .A(y[3569]), .B(x[3569]), .Z(n22433) );
  AND U5909 ( .A(n22426), .B(n22433), .Z(n28982) );
  NANDN U5910 ( .A(x[3565]), .B(y[3565]), .Z(n11750) );
  NANDN U5911 ( .A(x[3566]), .B(y[3566]), .Z(n22423) );
  NAND U5912 ( .A(n11750), .B(n22423), .Z(n23971) );
  NANDN U5913 ( .A(y[3564]), .B(x[3564]), .Z(n11752) );
  NANDN U5914 ( .A(y[3565]), .B(x[3565]), .Z(n11749) );
  AND U5915 ( .A(n11752), .B(n11749), .Z(n28980) );
  NANDN U5916 ( .A(x[3561]), .B(y[3561]), .Z(n3948) );
  NANDN U5917 ( .A(x[3562]), .B(y[3562]), .Z(n3947) );
  NAND U5918 ( .A(n3948), .B(n3947), .Z(n28976) );
  NANDN U5919 ( .A(y[3559]), .B(x[3559]), .Z(n3950) );
  NANDN U5920 ( .A(y[3558]), .B(x[3558]), .Z(n3949) );
  AND U5921 ( .A(n3950), .B(n3949), .Z(n28972) );
  NANDN U5922 ( .A(x[3557]), .B(y[3557]), .Z(n3952) );
  NANDN U5923 ( .A(x[3558]), .B(y[3558]), .Z(n3951) );
  AND U5924 ( .A(n3952), .B(n3951), .Z(n28971) );
  NANDN U5925 ( .A(y[3556]), .B(x[3556]), .Z(n3953) );
  ANDN U5926 ( .B(x[3557]), .A(y[3557]), .Z(n22401) );
  ANDN U5927 ( .B(n3953), .A(n22401), .Z(n28970) );
  NANDN U5928 ( .A(x[3556]), .B(y[3556]), .Z(n3954) );
  NANDN U5929 ( .A(x[3555]), .B(y[3555]), .Z(n11755) );
  NAND U5930 ( .A(n3954), .B(n11755), .Z(n28969) );
  NANDN U5931 ( .A(y[3554]), .B(x[3554]), .Z(n22394) );
  NANDN U5932 ( .A(y[3555]), .B(x[3555]), .Z(n22400) );
  AND U5933 ( .A(n22394), .B(n22400), .Z(n28968) );
  NANDN U5934 ( .A(y[3552]), .B(x[3552]), .Z(n22388) );
  NANDN U5935 ( .A(y[3553]), .B(x[3553]), .Z(n22395) );
  AND U5936 ( .A(n22388), .B(n22395), .Z(n28966) );
  NANDN U5937 ( .A(x[3551]), .B(y[3551]), .Z(n11759) );
  NANDN U5938 ( .A(x[3552]), .B(y[3552]), .Z(n11758) );
  NAND U5939 ( .A(n11759), .B(n11758), .Z(n28965) );
  NANDN U5940 ( .A(y[3550]), .B(x[3550]), .Z(n11761) );
  NANDN U5941 ( .A(y[3551]), .B(x[3551]), .Z(n22389) );
  AND U5942 ( .A(n11761), .B(n22389), .Z(n28964) );
  NANDN U5943 ( .A(x[3549]), .B(y[3549]), .Z(n11763) );
  NANDN U5944 ( .A(x[3550]), .B(y[3550]), .Z(n11760) );
  NAND U5945 ( .A(n11763), .B(n11760), .Z(n28963) );
  NANDN U5946 ( .A(y[3548]), .B(x[3548]), .Z(n22380) );
  NANDN U5947 ( .A(y[3549]), .B(x[3549]), .Z(n11762) );
  AND U5948 ( .A(n22380), .B(n11762), .Z(n28962) );
  NANDN U5949 ( .A(x[3547]), .B(y[3547]), .Z(n11765) );
  NANDN U5950 ( .A(x[3548]), .B(y[3548]), .Z(n11764) );
  NAND U5951 ( .A(n11765), .B(n11764), .Z(n28961) );
  NANDN U5952 ( .A(y[3546]), .B(x[3546]), .Z(n22371) );
  ANDN U5953 ( .B(x[3547]), .A(y[3547]), .Z(n22378) );
  ANDN U5954 ( .B(n22371), .A(n22378), .Z(n28960) );
  NANDN U5955 ( .A(x[3545]), .B(y[3545]), .Z(n11767) );
  NANDN U5956 ( .A(x[3546]), .B(y[3546]), .Z(n11766) );
  AND U5957 ( .A(n11767), .B(n11766), .Z(n23972) );
  NANDN U5958 ( .A(y[3544]), .B(x[3544]), .Z(n22365) );
  NANDN U5959 ( .A(y[3545]), .B(x[3545]), .Z(n22372) );
  NAND U5960 ( .A(n22365), .B(n22372), .Z(n28959) );
  NANDN U5961 ( .A(x[3543]), .B(y[3543]), .Z(n11769) );
  NANDN U5962 ( .A(x[3544]), .B(y[3544]), .Z(n11768) );
  AND U5963 ( .A(n11769), .B(n11768), .Z(n28958) );
  NANDN U5964 ( .A(y[3542]), .B(x[3542]), .Z(n22359) );
  NANDN U5965 ( .A(y[3543]), .B(x[3543]), .Z(n22366) );
  NAND U5966 ( .A(n22359), .B(n22366), .Z(n28957) );
  NANDN U5967 ( .A(x[3541]), .B(y[3541]), .Z(n11771) );
  NANDN U5968 ( .A(x[3542]), .B(y[3542]), .Z(n11770) );
  AND U5969 ( .A(n11771), .B(n11770), .Z(n28955) );
  NANDN U5970 ( .A(x[3539]), .B(y[3539]), .Z(n11773) );
  NANDN U5971 ( .A(x[3540]), .B(y[3540]), .Z(n11772) );
  AND U5972 ( .A(n11773), .B(n11772), .Z(n28953) );
  NANDN U5973 ( .A(y[3538]), .B(x[3538]), .Z(n11775) );
  NANDN U5974 ( .A(y[3539]), .B(x[3539]), .Z(n22354) );
  NAND U5975 ( .A(n11775), .B(n22354), .Z(n28952) );
  NANDN U5976 ( .A(x[3538]), .B(y[3538]), .Z(n11774) );
  ANDN U5977 ( .B(y[3537]), .A(x[3537]), .Z(n22346) );
  ANDN U5978 ( .B(n11774), .A(n22346), .Z(n28951) );
  NANDN U5979 ( .A(y[3536]), .B(x[3536]), .Z(n11777) );
  NANDN U5980 ( .A(y[3537]), .B(x[3537]), .Z(n11776) );
  NAND U5981 ( .A(n11777), .B(n11776), .Z(n28950) );
  ANDN U5982 ( .B(y[3535]), .A(x[3535]), .Z(n22341) );
  ANDN U5983 ( .B(y[3536]), .A(x[3536]), .Z(n22347) );
  NOR U5984 ( .A(n22341), .B(n22347), .Z(n28949) );
  XNOR U5985 ( .A(x[3534]), .B(y[3534]), .Z(n11780) );
  NANDN U5986 ( .A(y[3532]), .B(x[3532]), .Z(n11782) );
  NANDN U5987 ( .A(y[3533]), .B(x[3533]), .Z(n11779) );
  NAND U5988 ( .A(n11782), .B(n11779), .Z(n28947) );
  NANDN U5989 ( .A(x[3531]), .B(y[3531]), .Z(n22331) );
  NANDN U5990 ( .A(x[3532]), .B(y[3532]), .Z(n11781) );
  AND U5991 ( .A(n22331), .B(n11781), .Z(n28946) );
  NANDN U5992 ( .A(y[3530]), .B(x[3530]), .Z(n3955) );
  NANDN U5993 ( .A(y[3531]), .B(x[3531]), .Z(n11783) );
  NAND U5994 ( .A(n3955), .B(n11783), .Z(n28945) );
  NANDN U5995 ( .A(y[3528]), .B(x[3528]), .Z(n3956) );
  NANDN U5996 ( .A(y[3529]), .B(x[3529]), .Z(n11784) );
  AND U5997 ( .A(n3956), .B(n11784), .Z(n28942) );
  XNOR U5998 ( .A(x[3528]), .B(y[3528]), .Z(n22324) );
  NANDN U5999 ( .A(y[3526]), .B(x[3526]), .Z(n3957) );
  NANDN U6000 ( .A(y[3527]), .B(x[3527]), .Z(n22325) );
  AND U6001 ( .A(n3957), .B(n22325), .Z(n28940) );
  ANDN U6002 ( .B(y[3525]), .A(x[3525]), .Z(n11787) );
  XNOR U6003 ( .A(x[3526]), .B(y[3526]), .Z(n22318) );
  NANDN U6004 ( .A(y[3524]), .B(x[3524]), .Z(n3958) );
  NANDN U6005 ( .A(y[3525]), .B(x[3525]), .Z(n22319) );
  NAND U6006 ( .A(n3958), .B(n22319), .Z(n28937) );
  XNOR U6007 ( .A(x[3524]), .B(y[3524]), .Z(n11789) );
  ANDN U6008 ( .B(y[3523]), .A(x[3523]), .Z(n11790) );
  XNOR U6009 ( .A(x[3522]), .B(y[3522]), .Z(n11792) );
  ANDN U6010 ( .B(y[3521]), .A(x[3521]), .Z(n22305) );
  ANDN U6011 ( .B(n11792), .A(n22305), .Z(n10589) );
  NANDN U6012 ( .A(y[3518]), .B(x[3518]), .Z(n3959) );
  NANDN U6013 ( .A(y[3519]), .B(x[3519]), .Z(n11794) );
  NAND U6014 ( .A(n3959), .B(n11794), .Z(n23979) );
  XNOR U6015 ( .A(x[3518]), .B(y[3518]), .Z(n11796) );
  NANDN U6016 ( .A(x[3517]), .B(y[3517]), .Z(n28930) );
  NANDN U6017 ( .A(x[3515]), .B(y[3515]), .Z(n22291) );
  NANDN U6018 ( .A(x[3516]), .B(y[3516]), .Z(n22296) );
  AND U6019 ( .A(n22291), .B(n22296), .Z(n28928) );
  XNOR U6020 ( .A(x[3514]), .B(y[3514]), .Z(n11800) );
  NANDN U6021 ( .A(y[3512]), .B(x[3512]), .Z(n11803) );
  NANDN U6022 ( .A(y[3513]), .B(x[3513]), .Z(n11799) );
  NAND U6023 ( .A(n11803), .B(n11799), .Z(n28926) );
  NANDN U6024 ( .A(x[3509]), .B(y[3509]), .Z(n22276) );
  NANDN U6025 ( .A(x[3510]), .B(y[3510]), .Z(n11805) );
  NAND U6026 ( .A(n22276), .B(n11805), .Z(n23984) );
  NANDN U6027 ( .A(y[3508]), .B(x[3508]), .Z(n11808) );
  NANDN U6028 ( .A(y[3509]), .B(x[3509]), .Z(n11807) );
  AND U6029 ( .A(n11808), .B(n11807), .Z(n28924) );
  NANDN U6030 ( .A(y[3504]), .B(x[3504]), .Z(n11812) );
  NANDN U6031 ( .A(y[3505]), .B(x[3505]), .Z(n11811) );
  AND U6032 ( .A(n11812), .B(n11811), .Z(n28921) );
  NANDN U6033 ( .A(x[3503]), .B(y[3503]), .Z(n22258) );
  NANDN U6034 ( .A(x[3504]), .B(y[3504]), .Z(n22265) );
  NAND U6035 ( .A(n22258), .B(n22265), .Z(n28920) );
  NANDN U6036 ( .A(y[3502]), .B(x[3502]), .Z(n11814) );
  NANDN U6037 ( .A(y[3503]), .B(x[3503]), .Z(n11813) );
  AND U6038 ( .A(n11814), .B(n11813), .Z(n28918) );
  NANDN U6039 ( .A(x[3501]), .B(y[3501]), .Z(n22252) );
  NANDN U6040 ( .A(x[3502]), .B(y[3502]), .Z(n22259) );
  NAND U6041 ( .A(n22252), .B(n22259), .Z(n28917) );
  NANDN U6042 ( .A(y[3500]), .B(x[3500]), .Z(n11816) );
  NANDN U6043 ( .A(y[3501]), .B(x[3501]), .Z(n11815) );
  AND U6044 ( .A(n11816), .B(n11815), .Z(n28916) );
  NANDN U6045 ( .A(x[3499]), .B(y[3499]), .Z(n22246) );
  NANDN U6046 ( .A(x[3500]), .B(y[3500]), .Z(n22253) );
  NAND U6047 ( .A(n22246), .B(n22253), .Z(n28915) );
  NANDN U6048 ( .A(y[3496]), .B(x[3496]), .Z(n11820) );
  NANDN U6049 ( .A(y[3497]), .B(x[3497]), .Z(n11819) );
  NAND U6050 ( .A(n11820), .B(n11819), .Z(n23987) );
  NANDN U6051 ( .A(x[3495]), .B(y[3495]), .Z(n22234) );
  NANDN U6052 ( .A(x[3496]), .B(y[3496]), .Z(n22241) );
  AND U6053 ( .A(n22234), .B(n22241), .Z(n28913) );
  NANDN U6054 ( .A(x[3491]), .B(y[3491]), .Z(n22222) );
  NANDN U6055 ( .A(x[3492]), .B(y[3492]), .Z(n22229) );
  AND U6056 ( .A(n22222), .B(n22229), .Z(n28910) );
  NANDN U6057 ( .A(y[3490]), .B(x[3490]), .Z(n22218) );
  NANDN U6058 ( .A(y[3491]), .B(x[3491]), .Z(n11825) );
  NAND U6059 ( .A(n22218), .B(n11825), .Z(n28909) );
  NANDN U6060 ( .A(x[3489]), .B(y[3489]), .Z(n22215) );
  NANDN U6061 ( .A(x[3490]), .B(y[3490]), .Z(n22223) );
  AND U6062 ( .A(n22215), .B(n22223), .Z(n28908) );
  NANDN U6063 ( .A(y[3488]), .B(x[3488]), .Z(n11826) );
  NANDN U6064 ( .A(y[3489]), .B(x[3489]), .Z(n22219) );
  NAND U6065 ( .A(n11826), .B(n22219), .Z(n28906) );
  NANDN U6066 ( .A(x[3487]), .B(y[3487]), .Z(n11828) );
  NANDN U6067 ( .A(x[3488]), .B(y[3488]), .Z(n22217) );
  AND U6068 ( .A(n11828), .B(n22217), .Z(n28905) );
  NANDN U6069 ( .A(x[3485]), .B(y[3485]), .Z(n28902) );
  XNOR U6070 ( .A(x[3486]), .B(y[3486]), .Z(n22207) );
  ANDN U6071 ( .B(x[3485]), .A(y[3485]), .Z(n22209) );
  NANDN U6072 ( .A(y[3484]), .B(x[3484]), .Z(n22201) );
  NANDN U6073 ( .A(n22209), .B(n22201), .Z(n23989) );
  NANDN U6074 ( .A(x[3483]), .B(y[3483]), .Z(n11830) );
  NANDN U6075 ( .A(x[3484]), .B(y[3484]), .Z(n11829) );
  AND U6076 ( .A(n11830), .B(n11829), .Z(n28901) );
  NANDN U6077 ( .A(y[3482]), .B(x[3482]), .Z(n11832) );
  NANDN U6078 ( .A(y[3483]), .B(x[3483]), .Z(n22202) );
  AND U6079 ( .A(n11832), .B(n22202), .Z(n28900) );
  NANDN U6080 ( .A(x[3481]), .B(y[3481]), .Z(n11834) );
  NANDN U6081 ( .A(x[3482]), .B(y[3482]), .Z(n11831) );
  NAND U6082 ( .A(n11834), .B(n11831), .Z(n28899) );
  NANDN U6083 ( .A(y[3480]), .B(x[3480]), .Z(n11836) );
  NANDN U6084 ( .A(y[3481]), .B(x[3481]), .Z(n11833) );
  AND U6085 ( .A(n11836), .B(n11833), .Z(n28898) );
  NANDN U6086 ( .A(x[3479]), .B(y[3479]), .Z(n22189) );
  NANDN U6087 ( .A(x[3480]), .B(y[3480]), .Z(n11835) );
  NAND U6088 ( .A(n22189), .B(n11835), .Z(n28897) );
  NANDN U6089 ( .A(y[3478]), .B(x[3478]), .Z(n11838) );
  NANDN U6090 ( .A(y[3479]), .B(x[3479]), .Z(n11837) );
  AND U6091 ( .A(n11838), .B(n11837), .Z(n28896) );
  ANDN U6092 ( .B(y[3478]), .A(x[3478]), .Z(n22191) );
  NANDN U6093 ( .A(x[3477]), .B(y[3477]), .Z(n22183) );
  NANDN U6094 ( .A(n22191), .B(n22183), .Z(n28895) );
  NANDN U6095 ( .A(y[3474]), .B(x[3474]), .Z(n11842) );
  NANDN U6096 ( .A(y[3475]), .B(x[3475]), .Z(n11841) );
  NAND U6097 ( .A(n11842), .B(n11841), .Z(n23991) );
  NANDN U6098 ( .A(x[3473]), .B(y[3473]), .Z(n22171) );
  NANDN U6099 ( .A(x[3474]), .B(y[3474]), .Z(n22178) );
  AND U6100 ( .A(n22171), .B(n22178), .Z(n28892) );
  XNOR U6101 ( .A(x[3470]), .B(y[3470]), .Z(n22163) );
  ANDN U6102 ( .B(x[3469]), .A(y[3469]), .Z(n22162) );
  NANDN U6103 ( .A(y[3468]), .B(x[3468]), .Z(n11848) );
  NANDN U6104 ( .A(n22162), .B(n11848), .Z(n23993) );
  NANDN U6105 ( .A(y[3466]), .B(x[3466]), .Z(n11851) );
  NANDN U6106 ( .A(y[3467]), .B(x[3467]), .Z(n11847) );
  AND U6107 ( .A(n11851), .B(n11847), .Z(n28886) );
  NANDN U6108 ( .A(x[3465]), .B(y[3465]), .Z(n22149) );
  NANDN U6109 ( .A(x[3466]), .B(y[3466]), .Z(n11850) );
  NAND U6110 ( .A(n22149), .B(n11850), .Z(n28885) );
  NANDN U6111 ( .A(y[3464]), .B(x[3464]), .Z(n11853) );
  NANDN U6112 ( .A(y[3465]), .B(x[3465]), .Z(n11852) );
  AND U6113 ( .A(n11853), .B(n11852), .Z(n28883) );
  NANDN U6114 ( .A(x[3463]), .B(y[3463]), .Z(n22143) );
  NANDN U6115 ( .A(x[3464]), .B(y[3464]), .Z(n22150) );
  NAND U6116 ( .A(n22143), .B(n22150), .Z(n28882) );
  NANDN U6117 ( .A(y[3462]), .B(x[3462]), .Z(n11855) );
  NANDN U6118 ( .A(y[3463]), .B(x[3463]), .Z(n11854) );
  AND U6119 ( .A(n11855), .B(n11854), .Z(n28881) );
  NANDN U6120 ( .A(x[3461]), .B(y[3461]), .Z(n11857) );
  NANDN U6121 ( .A(x[3462]), .B(y[3462]), .Z(n22144) );
  NAND U6122 ( .A(n11857), .B(n22144), .Z(n28880) );
  NANDN U6123 ( .A(x[3460]), .B(y[3460]), .Z(n11858) );
  ANDN U6124 ( .B(y[3459]), .A(x[3459]), .Z(n22136) );
  ANDN U6125 ( .B(n11858), .A(n22136), .Z(n28878) );
  NANDN U6126 ( .A(y[3458]), .B(x[3458]), .Z(n3961) );
  NANDN U6127 ( .A(y[3459]), .B(x[3459]), .Z(n3960) );
  NAND U6128 ( .A(n3961), .B(n3960), .Z(n11859) );
  NANDN U6129 ( .A(x[3458]), .B(y[3458]), .Z(n3963) );
  NANDN U6130 ( .A(x[3457]), .B(y[3457]), .Z(n3962) );
  AND U6131 ( .A(n3963), .B(n3962), .Z(n11860) );
  ANDN U6132 ( .B(y[3455]), .A(x[3455]), .Z(n22124) );
  ANDN U6133 ( .B(y[3456]), .A(x[3456]), .Z(n22131) );
  NOR U6134 ( .A(n22124), .B(n22131), .Z(n28874) );
  NANDN U6135 ( .A(y[3454]), .B(x[3454]), .Z(n11863) );
  NANDN U6136 ( .A(y[3455]), .B(x[3455]), .Z(n11862) );
  NAND U6137 ( .A(n11863), .B(n11862), .Z(n23994) );
  NANDN U6138 ( .A(x[3453]), .B(y[3453]), .Z(n11865) );
  ANDN U6139 ( .B(y[3454]), .A(x[3454]), .Z(n22125) );
  ANDN U6140 ( .B(n11865), .A(n22125), .Z(n28873) );
  NANDN U6141 ( .A(x[3451]), .B(y[3451]), .Z(n22114) );
  NANDN U6142 ( .A(x[3452]), .B(y[3452]), .Z(n11866) );
  AND U6143 ( .A(n22114), .B(n11866), .Z(n28872) );
  XNOR U6144 ( .A(x[3450]), .B(y[3450]), .Z(n22111) );
  NANDN U6145 ( .A(x[3447]), .B(y[3447]), .Z(n11872) );
  NANDN U6146 ( .A(x[3448]), .B(y[3448]), .Z(n11869) );
  AND U6147 ( .A(n11872), .B(n11869), .Z(n28868) );
  NANDN U6148 ( .A(y[3446]), .B(x[3446]), .Z(n11874) );
  NANDN U6149 ( .A(y[3447]), .B(x[3447]), .Z(n11870) );
  NAND U6150 ( .A(n11874), .B(n11870), .Z(n28867) );
  NANDN U6151 ( .A(x[3445]), .B(y[3445]), .Z(n22098) );
  NANDN U6152 ( .A(x[3446]), .B(y[3446]), .Z(n11873) );
  AND U6153 ( .A(n22098), .B(n11873), .Z(n28866) );
  NANDN U6154 ( .A(y[3444]), .B(x[3444]), .Z(n11876) );
  NANDN U6155 ( .A(y[3445]), .B(x[3445]), .Z(n11875) );
  NAND U6156 ( .A(n11876), .B(n11875), .Z(n28865) );
  NANDN U6157 ( .A(x[3443]), .B(y[3443]), .Z(n22092) );
  NANDN U6158 ( .A(x[3444]), .B(y[3444]), .Z(n22099) );
  AND U6159 ( .A(n22092), .B(n22099), .Z(n28864) );
  NANDN U6160 ( .A(y[3442]), .B(x[3442]), .Z(n22089) );
  NANDN U6161 ( .A(y[3443]), .B(x[3443]), .Z(n11877) );
  NAND U6162 ( .A(n22089), .B(n11877), .Z(n28863) );
  NANDN U6163 ( .A(x[3441]), .B(y[3441]), .Z(n11878) );
  NANDN U6164 ( .A(x[3442]), .B(y[3442]), .Z(n22093) );
  AND U6165 ( .A(n11878), .B(n22093), .Z(n28862) );
  NANDN U6166 ( .A(y[3436]), .B(x[3436]), .Z(n22071) );
  NANDN U6167 ( .A(y[3437]), .B(x[3437]), .Z(n22078) );
  NAND U6168 ( .A(n22071), .B(n22078), .Z(n28859) );
  NANDN U6169 ( .A(x[3436]), .B(y[3436]), .Z(n11883) );
  ANDN U6170 ( .B(y[3435]), .A(x[3435]), .Z(n22069) );
  ANDN U6171 ( .B(n11883), .A(n22069), .Z(n28858) );
  XNOR U6172 ( .A(x[3434]), .B(y[3434]), .Z(n11885) );
  NANDN U6173 ( .A(x[3433]), .B(y[3433]), .Z(n24001) );
  AND U6174 ( .A(n11885), .B(n24001), .Z(n10489) );
  NANDN U6175 ( .A(y[3430]), .B(x[3430]), .Z(n22055) );
  NANDN U6176 ( .A(y[3431]), .B(x[3431]), .Z(n11888) );
  NAND U6177 ( .A(n22055), .B(n11888), .Z(n28854) );
  NANDN U6178 ( .A(x[3429]), .B(y[3429]), .Z(n11891) );
  NANDN U6179 ( .A(x[3430]), .B(y[3430]), .Z(n11890) );
  AND U6180 ( .A(n11891), .B(n11890), .Z(n24003) );
  NANDN U6181 ( .A(y[3428]), .B(x[3428]), .Z(n22049) );
  NANDN U6182 ( .A(y[3429]), .B(x[3429]), .Z(n22056) );
  NAND U6183 ( .A(n22049), .B(n22056), .Z(n28853) );
  NANDN U6184 ( .A(x[3427]), .B(y[3427]), .Z(n11893) );
  NANDN U6185 ( .A(x[3428]), .B(y[3428]), .Z(n11892) );
  AND U6186 ( .A(n11893), .B(n11892), .Z(n28852) );
  NANDN U6187 ( .A(y[3426]), .B(x[3426]), .Z(n22043) );
  NANDN U6188 ( .A(y[3427]), .B(x[3427]), .Z(n22050) );
  NAND U6189 ( .A(n22043), .B(n22050), .Z(n28851) );
  NANDN U6190 ( .A(x[3423]), .B(y[3423]), .Z(n11897) );
  NANDN U6191 ( .A(x[3424]), .B(y[3424]), .Z(n11896) );
  NAND U6192 ( .A(n11897), .B(n11896), .Z(n28849) );
  NANDN U6193 ( .A(y[3422]), .B(x[3422]), .Z(n22031) );
  NANDN U6194 ( .A(y[3423]), .B(x[3423]), .Z(n22038) );
  AND U6195 ( .A(n22031), .B(n22038), .Z(n28848) );
  NANDN U6196 ( .A(x[3421]), .B(y[3421]), .Z(n11899) );
  NANDN U6197 ( .A(x[3422]), .B(y[3422]), .Z(n11898) );
  NAND U6198 ( .A(n11899), .B(n11898), .Z(n28847) );
  NANDN U6199 ( .A(y[3420]), .B(x[3420]), .Z(n22025) );
  NANDN U6200 ( .A(y[3421]), .B(x[3421]), .Z(n22032) );
  AND U6201 ( .A(n22025), .B(n22032), .Z(n28845) );
  NANDN U6202 ( .A(x[3417]), .B(y[3417]), .Z(n11903) );
  NANDN U6203 ( .A(x[3418]), .B(y[3418]), .Z(n11902) );
  NAND U6204 ( .A(n11903), .B(n11902), .Z(n24006) );
  NANDN U6205 ( .A(y[3416]), .B(x[3416]), .Z(n22013) );
  NANDN U6206 ( .A(y[3417]), .B(x[3417]), .Z(n22020) );
  AND U6207 ( .A(n22013), .B(n22020), .Z(n28843) );
  NANDN U6208 ( .A(x[3413]), .B(y[3413]), .Z(n11907) );
  NANDN U6209 ( .A(x[3414]), .B(y[3414]), .Z(n11906) );
  NAND U6210 ( .A(n11907), .B(n11906), .Z(n28841) );
  NANDN U6211 ( .A(y[3410]), .B(x[3410]), .Z(n21995) );
  NANDN U6212 ( .A(y[3411]), .B(x[3411]), .Z(n22002) );
  NAND U6213 ( .A(n21995), .B(n22002), .Z(n28838) );
  NANDN U6214 ( .A(x[3409]), .B(y[3409]), .Z(n11911) );
  NANDN U6215 ( .A(x[3410]), .B(y[3410]), .Z(n11910) );
  AND U6216 ( .A(n11911), .B(n11910), .Z(n24008) );
  NANDN U6217 ( .A(y[3408]), .B(x[3408]), .Z(n21989) );
  NANDN U6218 ( .A(y[3409]), .B(x[3409]), .Z(n21996) );
  NAND U6219 ( .A(n21989), .B(n21996), .Z(n28836) );
  NANDN U6220 ( .A(x[3407]), .B(y[3407]), .Z(n11913) );
  NANDN U6221 ( .A(x[3408]), .B(y[3408]), .Z(n11912) );
  AND U6222 ( .A(n11913), .B(n11912), .Z(n28835) );
  XNOR U6223 ( .A(x[3406]), .B(y[3406]), .Z(n21984) );
  NANDN U6224 ( .A(y[3404]), .B(x[3404]), .Z(n11915) );
  NANDN U6225 ( .A(y[3405]), .B(x[3405]), .Z(n21983) );
  NAND U6226 ( .A(n11915), .B(n21983), .Z(n24011) );
  NANDN U6227 ( .A(x[3404]), .B(y[3404]), .Z(n11914) );
  ANDN U6228 ( .B(y[3403]), .A(x[3403]), .Z(n21976) );
  ANDN U6229 ( .B(n11914), .A(n21976), .Z(n28833) );
  ANDN U6230 ( .B(y[3401]), .A(x[3401]), .Z(n21971) );
  ANDN U6231 ( .B(y[3402]), .A(x[3402]), .Z(n21977) );
  NOR U6232 ( .A(n21971), .B(n21977), .Z(n28832) );
  XNOR U6233 ( .A(x[3400]), .B(y[3400]), .Z(n11920) );
  NANDN U6234 ( .A(y[3398]), .B(x[3398]), .Z(n3964) );
  NANDN U6235 ( .A(y[3399]), .B(x[3399]), .Z(n11919) );
  NAND U6236 ( .A(n3964), .B(n11919), .Z(n28828) );
  XNOR U6237 ( .A(x[3398]), .B(y[3398]), .Z(n21964) );
  ANDN U6238 ( .B(x[3396]), .A(y[3396]), .Z(n21957) );
  ANDN U6239 ( .B(x[3397]), .A(y[3397]), .Z(n21963) );
  OR U6240 ( .A(n21957), .B(n21963), .Z(n24015) );
  NANDN U6241 ( .A(x[3395]), .B(y[3395]), .Z(n21955) );
  NANDN U6242 ( .A(x[3396]), .B(y[3396]), .Z(n11921) );
  AND U6243 ( .A(n21955), .B(n11921), .Z(n24016) );
  NANDN U6244 ( .A(y[3392]), .B(x[3392]), .Z(n3966) );
  NANDN U6245 ( .A(y[3393]), .B(x[3393]), .Z(n3965) );
  NAND U6246 ( .A(n3966), .B(n3965), .Z(n28824) );
  NANDN U6247 ( .A(x[3392]), .B(y[3392]), .Z(n3968) );
  NANDN U6248 ( .A(x[3391]), .B(y[3391]), .Z(n3967) );
  AND U6249 ( .A(n3968), .B(n3967), .Z(n28823) );
  ANDN U6250 ( .B(x[3389]), .A(y[3389]), .Z(n21946) );
  NANDN U6251 ( .A(y[3388]), .B(x[3388]), .Z(n11922) );
  NANDN U6252 ( .A(n21946), .B(n11922), .Z(n24019) );
  NANDN U6253 ( .A(x[3388]), .B(y[3388]), .Z(n21944) );
  NANDN U6254 ( .A(x[3387]), .B(y[3387]), .Z(n11924) );
  AND U6255 ( .A(n21944), .B(n11924), .Z(n28821) );
  NANDN U6256 ( .A(y[3384]), .B(x[3384]), .Z(n21929) );
  NANDN U6257 ( .A(y[3385]), .B(x[3385]), .Z(n21936) );
  NAND U6258 ( .A(n21929), .B(n21936), .Z(n28816) );
  NANDN U6259 ( .A(x[3383]), .B(y[3383]), .Z(n11928) );
  NANDN U6260 ( .A(x[3384]), .B(y[3384]), .Z(n11927) );
  AND U6261 ( .A(n11928), .B(n11927), .Z(n28815) );
  NANDN U6262 ( .A(y[3382]), .B(x[3382]), .Z(n21923) );
  NANDN U6263 ( .A(y[3383]), .B(x[3383]), .Z(n21930) );
  AND U6264 ( .A(n21923), .B(n21930), .Z(n28814) );
  NANDN U6265 ( .A(x[3381]), .B(y[3381]), .Z(n11930) );
  NANDN U6266 ( .A(x[3382]), .B(y[3382]), .Z(n11929) );
  NAND U6267 ( .A(n11930), .B(n11929), .Z(n28813) );
  NANDN U6268 ( .A(y[3380]), .B(x[3380]), .Z(n21917) );
  NANDN U6269 ( .A(y[3381]), .B(x[3381]), .Z(n21924) );
  AND U6270 ( .A(n21917), .B(n21924), .Z(n24021) );
  NANDN U6271 ( .A(x[3379]), .B(y[3379]), .Z(n11932) );
  NANDN U6272 ( .A(x[3380]), .B(y[3380]), .Z(n11931) );
  NAND U6273 ( .A(n11932), .B(n11931), .Z(n28812) );
  NANDN U6274 ( .A(y[3378]), .B(x[3378]), .Z(n21911) );
  NANDN U6275 ( .A(y[3379]), .B(x[3379]), .Z(n21918) );
  AND U6276 ( .A(n21911), .B(n21918), .Z(n28811) );
  NANDN U6277 ( .A(x[3377]), .B(y[3377]), .Z(n11934) );
  NANDN U6278 ( .A(x[3378]), .B(y[3378]), .Z(n11933) );
  NAND U6279 ( .A(n11934), .B(n11933), .Z(n28810) );
  NANDN U6280 ( .A(y[3374]), .B(x[3374]), .Z(n21899) );
  NANDN U6281 ( .A(y[3375]), .B(x[3375]), .Z(n21906) );
  NAND U6282 ( .A(n21899), .B(n21906), .Z(n28808) );
  NANDN U6283 ( .A(x[3373]), .B(y[3373]), .Z(n11938) );
  NANDN U6284 ( .A(x[3374]), .B(y[3374]), .Z(n11937) );
  AND U6285 ( .A(n11938), .B(n11937), .Z(n28807) );
  NANDN U6286 ( .A(y[3372]), .B(x[3372]), .Z(n21893) );
  NANDN U6287 ( .A(y[3373]), .B(x[3373]), .Z(n21900) );
  NAND U6288 ( .A(n21893), .B(n21900), .Z(n28806) );
  NANDN U6289 ( .A(x[3371]), .B(y[3371]), .Z(n21889) );
  NANDN U6290 ( .A(x[3372]), .B(y[3372]), .Z(n11939) );
  AND U6291 ( .A(n21889), .B(n11939), .Z(n28805) );
  NANDN U6292 ( .A(x[3370]), .B(y[3370]), .Z(n21890) );
  ANDN U6293 ( .B(y[3369]), .A(x[3369]), .Z(n21884) );
  ANDN U6294 ( .B(n21890), .A(n21884), .Z(n28803) );
  NANDN U6295 ( .A(y[3368]), .B(x[3368]), .Z(n11942) );
  NANDN U6296 ( .A(y[3369]), .B(x[3369]), .Z(n11941) );
  NAND U6297 ( .A(n11942), .B(n11941), .Z(n24023) );
  ANDN U6298 ( .B(y[3367]), .A(x[3367]), .Z(n21879) );
  ANDN U6299 ( .B(y[3368]), .A(x[3368]), .Z(n21885) );
  NOR U6300 ( .A(n21879), .B(n21885), .Z(n28801) );
  XNOR U6301 ( .A(x[3366]), .B(y[3366]), .Z(n11945) );
  ANDN U6302 ( .B(y[3365]), .A(x[3365]), .Z(n28798) );
  ANDN U6303 ( .B(n11945), .A(n28798), .Z(n10408) );
  NANDN U6304 ( .A(y[3362]), .B(x[3362]), .Z(n11949) );
  NANDN U6305 ( .A(y[3363]), .B(x[3363]), .Z(n11946) );
  AND U6306 ( .A(n11949), .B(n11946), .Z(n28796) );
  NANDN U6307 ( .A(x[3357]), .B(y[3357]), .Z(n21852) );
  NANDN U6308 ( .A(x[3358]), .B(y[3358]), .Z(n21859) );
  NAND U6309 ( .A(n21852), .B(n21859), .Z(n28790) );
  NANDN U6310 ( .A(y[3356]), .B(x[3356]), .Z(n21848) );
  NANDN U6311 ( .A(y[3357]), .B(x[3357]), .Z(n11954) );
  AND U6312 ( .A(n21848), .B(n11954), .Z(n24028) );
  NANDN U6313 ( .A(x[3355]), .B(y[3355]), .Z(n11955) );
  NANDN U6314 ( .A(x[3356]), .B(y[3356]), .Z(n21853) );
  NAND U6315 ( .A(n11955), .B(n21853), .Z(n28789) );
  NANDN U6316 ( .A(y[3355]), .B(x[3355]), .Z(n21849) );
  ANDN U6317 ( .B(x[3354]), .A(y[3354]), .Z(n21845) );
  ANDN U6318 ( .B(n21849), .A(n21845), .Z(n28788) );
  NANDN U6319 ( .A(x[3353]), .B(y[3353]), .Z(n21843) );
  NANDN U6320 ( .A(x[3354]), .B(y[3354]), .Z(n11956) );
  NAND U6321 ( .A(n21843), .B(n11956), .Z(n28787) );
  ANDN U6322 ( .B(x[3351]), .A(y[3351]), .Z(n21837) );
  NANDN U6323 ( .A(y[3350]), .B(x[3350]), .Z(n3969) );
  NANDN U6324 ( .A(n21837), .B(n3969), .Z(n11957) );
  NANDN U6325 ( .A(x[3349]), .B(y[3349]), .Z(n11960) );
  NANDN U6326 ( .A(x[3350]), .B(y[3350]), .Z(n21836) );
  AND U6327 ( .A(n11960), .B(n21836), .Z(n24030) );
  NANDN U6328 ( .A(y[3346]), .B(x[3346]), .Z(n21824) );
  NANDN U6329 ( .A(y[3347]), .B(x[3347]), .Z(n11962) );
  NAND U6330 ( .A(n21824), .B(n11962), .Z(n28783) );
  NANDN U6331 ( .A(x[3345]), .B(y[3345]), .Z(n11965) );
  NANDN U6332 ( .A(x[3346]), .B(y[3346]), .Z(n11964) );
  AND U6333 ( .A(n11965), .B(n11964), .Z(n24032) );
  NANDN U6334 ( .A(y[3344]), .B(x[3344]), .Z(n21818) );
  NANDN U6335 ( .A(y[3345]), .B(x[3345]), .Z(n21825) );
  NAND U6336 ( .A(n21818), .B(n21825), .Z(n28782) );
  NANDN U6337 ( .A(x[3343]), .B(y[3343]), .Z(n11967) );
  NANDN U6338 ( .A(x[3344]), .B(y[3344]), .Z(n11966) );
  AND U6339 ( .A(n11967), .B(n11966), .Z(n28780) );
  NANDN U6340 ( .A(x[3341]), .B(y[3341]), .Z(n11969) );
  NANDN U6341 ( .A(x[3342]), .B(y[3342]), .Z(n11968) );
  AND U6342 ( .A(n11969), .B(n11968), .Z(n28778) );
  NANDN U6343 ( .A(y[3340]), .B(x[3340]), .Z(n21806) );
  NANDN U6344 ( .A(y[3341]), .B(x[3341]), .Z(n21813) );
  NAND U6345 ( .A(n21806), .B(n21813), .Z(n28777) );
  NANDN U6346 ( .A(x[3339]), .B(y[3339]), .Z(n11971) );
  NANDN U6347 ( .A(x[3340]), .B(y[3340]), .Z(n11970) );
  AND U6348 ( .A(n11971), .B(n11970), .Z(n24033) );
  NANDN U6349 ( .A(y[3336]), .B(x[3336]), .Z(n21795) );
  NANDN U6350 ( .A(y[3337]), .B(x[3337]), .Z(n21801) );
  NAND U6351 ( .A(n21795), .B(n21801), .Z(n28775) );
  NANDN U6352 ( .A(y[3334]), .B(x[3334]), .Z(n21786) );
  ANDN U6353 ( .B(x[3335]), .A(y[3335]), .Z(n21793) );
  ANDN U6354 ( .B(n21786), .A(n21793), .Z(n28774) );
  NANDN U6355 ( .A(x[3333]), .B(y[3333]), .Z(n11975) );
  NANDN U6356 ( .A(x[3334]), .B(y[3334]), .Z(n11974) );
  NAND U6357 ( .A(n11975), .B(n11974), .Z(n24036) );
  NANDN U6358 ( .A(y[3332]), .B(x[3332]), .Z(n21780) );
  NANDN U6359 ( .A(y[3333]), .B(x[3333]), .Z(n21787) );
  AND U6360 ( .A(n21780), .B(n21787), .Z(n28773) );
  NANDN U6361 ( .A(y[3328]), .B(x[3328]), .Z(n21768) );
  NANDN U6362 ( .A(y[3329]), .B(x[3329]), .Z(n21775) );
  AND U6363 ( .A(n21768), .B(n21775), .Z(n28768) );
  NANDN U6364 ( .A(x[3327]), .B(y[3327]), .Z(n11981) );
  NANDN U6365 ( .A(x[3328]), .B(y[3328]), .Z(n11980) );
  NAND U6366 ( .A(n11981), .B(n11980), .Z(n28767) );
  NANDN U6367 ( .A(y[3326]), .B(x[3326]), .Z(n21762) );
  NANDN U6368 ( .A(y[3327]), .B(x[3327]), .Z(n21769) );
  AND U6369 ( .A(n21762), .B(n21769), .Z(n28766) );
  NANDN U6370 ( .A(x[3325]), .B(y[3325]), .Z(n11983) );
  NANDN U6371 ( .A(x[3326]), .B(y[3326]), .Z(n11982) );
  NAND U6372 ( .A(n11983), .B(n11982), .Z(n28765) );
  NANDN U6373 ( .A(x[3323]), .B(y[3323]), .Z(n21752) );
  NANDN U6374 ( .A(x[3324]), .B(y[3324]), .Z(n11984) );
  NAND U6375 ( .A(n21752), .B(n11984), .Z(n24039) );
  NANDN U6376 ( .A(x[3321]), .B(y[3321]), .Z(n11985) );
  NANDN U6377 ( .A(x[3322]), .B(y[3322]), .Z(n21753) );
  AND U6378 ( .A(n11985), .B(n21753), .Z(n28763) );
  NANDN U6379 ( .A(y[3320]), .B(x[3320]), .Z(n11987) );
  NANDN U6380 ( .A(y[3321]), .B(x[3321]), .Z(n21751) );
  NAND U6381 ( .A(n11987), .B(n21751), .Z(n28762) );
  NANDN U6382 ( .A(x[3320]), .B(y[3320]), .Z(n11986) );
  ANDN U6383 ( .B(y[3319]), .A(x[3319]), .Z(n21741) );
  ANDN U6384 ( .B(n11986), .A(n21741), .Z(n28761) );
  ANDN U6385 ( .B(y[3317]), .A(x[3317]), .Z(n21736) );
  ANDN U6386 ( .B(y[3318]), .A(x[3318]), .Z(n21742) );
  NOR U6387 ( .A(n21736), .B(n21742), .Z(n28760) );
  XNOR U6388 ( .A(x[3316]), .B(y[3316]), .Z(n11992) );
  NANDN U6389 ( .A(y[3314]), .B(x[3314]), .Z(n21730) );
  NANDN U6390 ( .A(y[3315]), .B(x[3315]), .Z(n11991) );
  NAND U6391 ( .A(n21730), .B(n11991), .Z(n28754) );
  ANDN U6392 ( .B(y[3312]), .A(x[3312]), .Z(n21724) );
  NANDN U6393 ( .A(x[3311]), .B(y[3311]), .Z(n21717) );
  NANDN U6394 ( .A(n21724), .B(n21717), .Z(n28751) );
  NANDN U6395 ( .A(y[3310]), .B(x[3310]), .Z(n11995) );
  NANDN U6396 ( .A(y[3311]), .B(x[3311]), .Z(n11994) );
  AND U6397 ( .A(n11995), .B(n11994), .Z(n24041) );
  NANDN U6398 ( .A(x[3309]), .B(y[3309]), .Z(n21711) );
  NANDN U6399 ( .A(x[3310]), .B(y[3310]), .Z(n21718) );
  NAND U6400 ( .A(n21711), .B(n21718), .Z(n28750) );
  NANDN U6401 ( .A(y[3308]), .B(x[3308]), .Z(n21707) );
  NANDN U6402 ( .A(y[3309]), .B(x[3309]), .Z(n11996) );
  AND U6403 ( .A(n21707), .B(n11996), .Z(n28749) );
  NANDN U6404 ( .A(x[3307]), .B(y[3307]), .Z(n11997) );
  NANDN U6405 ( .A(x[3308]), .B(y[3308]), .Z(n21712) );
  NAND U6406 ( .A(n11997), .B(n21712), .Z(n28748) );
  NANDN U6407 ( .A(y[3304]), .B(x[3304]), .Z(n12003) );
  NANDN U6408 ( .A(y[3305]), .B(x[3305]), .Z(n12000) );
  NAND U6409 ( .A(n12003), .B(n12000), .Z(n28746) );
  NANDN U6410 ( .A(x[3303]), .B(y[3303]), .Z(n21696) );
  NANDN U6411 ( .A(x[3304]), .B(y[3304]), .Z(n12002) );
  AND U6412 ( .A(n21696), .B(n12002), .Z(n28745) );
  NANDN U6413 ( .A(y[3302]), .B(x[3302]), .Z(n3970) );
  NANDN U6414 ( .A(y[3303]), .B(x[3303]), .Z(n12004) );
  NAND U6415 ( .A(n3970), .B(n12004), .Z(n28744) );
  XNOR U6416 ( .A(x[3302]), .B(y[3302]), .Z(n21693) );
  NANDN U6417 ( .A(x[3301]), .B(y[3301]), .Z(n24043) );
  AND U6418 ( .A(n21693), .B(n24043), .Z(n10334) );
  NANDN U6419 ( .A(y[3298]), .B(x[3298]), .Z(n12010) );
  NANDN U6420 ( .A(y[3299]), .B(x[3299]), .Z(n12006) );
  NAND U6421 ( .A(n12010), .B(n12006), .Z(n24047) );
  NANDN U6422 ( .A(x[3297]), .B(y[3297]), .Z(n21680) );
  NANDN U6423 ( .A(x[3298]), .B(y[3298]), .Z(n12009) );
  AND U6424 ( .A(n21680), .B(n12009), .Z(n28742) );
  NANDN U6425 ( .A(x[3293]), .B(y[3293]), .Z(n21668) );
  NANDN U6426 ( .A(x[3294]), .B(y[3294]), .Z(n21675) );
  AND U6427 ( .A(n21668), .B(n21675), .Z(n28739) );
  NANDN U6428 ( .A(y[3292]), .B(x[3292]), .Z(n21665) );
  NANDN U6429 ( .A(y[3293]), .B(x[3293]), .Z(n12015) );
  NAND U6430 ( .A(n21665), .B(n12015), .Z(n28738) );
  NANDN U6431 ( .A(x[3291]), .B(y[3291]), .Z(n12016) );
  NANDN U6432 ( .A(x[3292]), .B(y[3292]), .Z(n21669) );
  AND U6433 ( .A(n12016), .B(n21669), .Z(n28737) );
  NANDN U6434 ( .A(y[3290]), .B(x[3290]), .Z(n3971) );
  NANDN U6435 ( .A(y[3291]), .B(x[3291]), .Z(n21666) );
  NAND U6436 ( .A(n3971), .B(n21666), .Z(n28736) );
  XNOR U6437 ( .A(x[3290]), .B(y[3290]), .Z(n21659) );
  NANDN U6438 ( .A(x[3289]), .B(y[3289]), .Z(n24049) );
  AND U6439 ( .A(n21659), .B(n24049), .Z(n10321) );
  NANDN U6440 ( .A(x[3288]), .B(y[3288]), .Z(n12017) );
  ANDN U6441 ( .B(y[3287]), .A(x[3287]), .Z(n21649) );
  ANDN U6442 ( .B(n12017), .A(n21649), .Z(n28732) );
  NANDN U6443 ( .A(y[3286]), .B(x[3286]), .Z(n21645) );
  NANDN U6444 ( .A(y[3287]), .B(x[3287]), .Z(n21654) );
  NAND U6445 ( .A(n21645), .B(n21654), .Z(n28731) );
  NANDN U6446 ( .A(x[3285]), .B(y[3285]), .Z(n12018) );
  ANDN U6447 ( .B(y[3286]), .A(x[3286]), .Z(n21651) );
  ANDN U6448 ( .B(n12018), .A(n21651), .Z(n28730) );
  NANDN U6449 ( .A(y[3284]), .B(x[3284]), .Z(n21638) );
  NANDN U6450 ( .A(y[3285]), .B(x[3285]), .Z(n21647) );
  NAND U6451 ( .A(n21638), .B(n21647), .Z(n28729) );
  NANDN U6452 ( .A(x[3283]), .B(y[3283]), .Z(n12020) );
  NANDN U6453 ( .A(x[3284]), .B(y[3284]), .Z(n12019) );
  AND U6454 ( .A(n12020), .B(n12019), .Z(n28728) );
  NANDN U6455 ( .A(y[3282]), .B(x[3282]), .Z(n21632) );
  NANDN U6456 ( .A(y[3283]), .B(x[3283]), .Z(n21639) );
  NAND U6457 ( .A(n21632), .B(n21639), .Z(n28727) );
  NANDN U6458 ( .A(x[3279]), .B(y[3279]), .Z(n21622) );
  NANDN U6459 ( .A(x[3280]), .B(y[3280]), .Z(n12023) );
  NAND U6460 ( .A(n21622), .B(n12023), .Z(n28725) );
  NANDN U6461 ( .A(y[3278]), .B(x[3278]), .Z(n21621) );
  NANDN U6462 ( .A(y[3279]), .B(x[3279]), .Z(n21627) );
  AND U6463 ( .A(n21621), .B(n21627), .Z(n28724) );
  NANDN U6464 ( .A(x[3277]), .B(y[3277]), .Z(n12024) );
  NANDN U6465 ( .A(x[3278]), .B(y[3278]), .Z(n21623) );
  NAND U6466 ( .A(n12024), .B(n21623), .Z(n28723) );
  NANDN U6467 ( .A(y[3276]), .B(x[3276]), .Z(n21612) );
  ANDN U6468 ( .B(x[3277]), .A(y[3277]), .Z(n21619) );
  ANDN U6469 ( .B(n21612), .A(n21619), .Z(n28722) );
  NANDN U6470 ( .A(x[3273]), .B(y[3273]), .Z(n12028) );
  NANDN U6471 ( .A(x[3274]), .B(y[3274]), .Z(n12027) );
  NAND U6472 ( .A(n12028), .B(n12027), .Z(n24053) );
  NANDN U6473 ( .A(y[3272]), .B(x[3272]), .Z(n21600) );
  NANDN U6474 ( .A(y[3273]), .B(x[3273]), .Z(n21607) );
  AND U6475 ( .A(n21600), .B(n21607), .Z(n28718) );
  NANDN U6476 ( .A(x[3269]), .B(y[3269]), .Z(n12032) );
  NANDN U6477 ( .A(x[3270]), .B(y[3270]), .Z(n12031) );
  NAND U6478 ( .A(n12032), .B(n12031), .Z(n28716) );
  NANDN U6479 ( .A(y[3266]), .B(x[3266]), .Z(n21582) );
  NANDN U6480 ( .A(y[3267]), .B(x[3267]), .Z(n21589) );
  NAND U6481 ( .A(n21582), .B(n21589), .Z(n28713) );
  NANDN U6482 ( .A(x[3265]), .B(y[3265]), .Z(n12036) );
  NANDN U6483 ( .A(x[3266]), .B(y[3266]), .Z(n12035) );
  AND U6484 ( .A(n12036), .B(n12035), .Z(n24055) );
  NANDN U6485 ( .A(y[3264]), .B(x[3264]), .Z(n21576) );
  NANDN U6486 ( .A(y[3265]), .B(x[3265]), .Z(n21583) );
  NAND U6487 ( .A(n21576), .B(n21583), .Z(n28712) );
  NANDN U6488 ( .A(x[3263]), .B(y[3263]), .Z(n12038) );
  NANDN U6489 ( .A(x[3264]), .B(y[3264]), .Z(n12037) );
  AND U6490 ( .A(n12038), .B(n12037), .Z(n28711) );
  NANDN U6491 ( .A(x[3261]), .B(y[3261]), .Z(n12040) );
  NANDN U6492 ( .A(x[3262]), .B(y[3262]), .Z(n12039) );
  AND U6493 ( .A(n12040), .B(n12039), .Z(n28709) );
  NANDN U6494 ( .A(y[3260]), .B(x[3260]), .Z(n21564) );
  NANDN U6495 ( .A(y[3261]), .B(x[3261]), .Z(n21571) );
  NAND U6496 ( .A(n21564), .B(n21571), .Z(n28707) );
  NANDN U6497 ( .A(x[3259]), .B(y[3259]), .Z(n12042) );
  NANDN U6498 ( .A(x[3260]), .B(y[3260]), .Z(n12041) );
  AND U6499 ( .A(n12042), .B(n12041), .Z(n24056) );
  XNOR U6500 ( .A(x[3256]), .B(y[3256]), .Z(n21553) );
  NANDN U6501 ( .A(y[3254]), .B(x[3254]), .Z(n21546) );
  NANDN U6502 ( .A(y[3255]), .B(x[3255]), .Z(n21552) );
  NAND U6503 ( .A(n21546), .B(n21552), .Z(n28702) );
  NANDN U6504 ( .A(x[3253]), .B(y[3253]), .Z(n12046) );
  NANDN U6505 ( .A(x[3254]), .B(y[3254]), .Z(n12045) );
  AND U6506 ( .A(n12046), .B(n12045), .Z(n28701) );
  NANDN U6507 ( .A(y[3252]), .B(x[3252]), .Z(n21540) );
  NANDN U6508 ( .A(y[3253]), .B(x[3253]), .Z(n21547) );
  NAND U6509 ( .A(n21540), .B(n21547), .Z(n28700) );
  NANDN U6510 ( .A(x[3251]), .B(y[3251]), .Z(n12048) );
  NANDN U6511 ( .A(x[3252]), .B(y[3252]), .Z(n12047) );
  AND U6512 ( .A(n12048), .B(n12047), .Z(n28699) );
  NANDN U6513 ( .A(y[3248]), .B(x[3248]), .Z(n21529) );
  NANDN U6514 ( .A(y[3249]), .B(x[3249]), .Z(n21535) );
  NAND U6515 ( .A(n21529), .B(n21535), .Z(n24059) );
  NANDN U6516 ( .A(x[3247]), .B(y[3247]), .Z(n12050) );
  NANDN U6517 ( .A(x[3248]), .B(y[3248]), .Z(n21531) );
  AND U6518 ( .A(n12050), .B(n21531), .Z(n28696) );
  NANDN U6519 ( .A(y[3244]), .B(x[3244]), .Z(n21514) );
  NANDN U6520 ( .A(y[3245]), .B(x[3245]), .Z(n21521) );
  NAND U6521 ( .A(n21514), .B(n21521), .Z(n28694) );
  NANDN U6522 ( .A(x[3241]), .B(y[3241]), .Z(n12056) );
  NANDN U6523 ( .A(x[3242]), .B(y[3242]), .Z(n12055) );
  NAND U6524 ( .A(n12056), .B(n12055), .Z(n28691) );
  NANDN U6525 ( .A(y[3240]), .B(x[3240]), .Z(n21502) );
  NANDN U6526 ( .A(y[3241]), .B(x[3241]), .Z(n21509) );
  AND U6527 ( .A(n21502), .B(n21509), .Z(n24061) );
  NANDN U6528 ( .A(x[3239]), .B(y[3239]), .Z(n12058) );
  NANDN U6529 ( .A(x[3240]), .B(y[3240]), .Z(n12057) );
  NAND U6530 ( .A(n12058), .B(n12057), .Z(n28690) );
  NANDN U6531 ( .A(y[3238]), .B(x[3238]), .Z(n21496) );
  NANDN U6532 ( .A(y[3239]), .B(x[3239]), .Z(n21503) );
  AND U6533 ( .A(n21496), .B(n21503), .Z(n28689) );
  NANDN U6534 ( .A(y[3236]), .B(x[3236]), .Z(n21490) );
  NANDN U6535 ( .A(y[3237]), .B(x[3237]), .Z(n21497) );
  AND U6536 ( .A(n21490), .B(n21497), .Z(n28687) );
  NANDN U6537 ( .A(x[3235]), .B(y[3235]), .Z(n12062) );
  NANDN U6538 ( .A(x[3236]), .B(y[3236]), .Z(n12061) );
  NAND U6539 ( .A(n12062), .B(n12061), .Z(n28686) );
  NANDN U6540 ( .A(y[3234]), .B(x[3234]), .Z(n21484) );
  NANDN U6541 ( .A(y[3235]), .B(x[3235]), .Z(n21491) );
  AND U6542 ( .A(n21484), .B(n21491), .Z(n24062) );
  NANDN U6543 ( .A(x[3231]), .B(y[3231]), .Z(n12066) );
  NANDN U6544 ( .A(x[3232]), .B(y[3232]), .Z(n12065) );
  NAND U6545 ( .A(n12066), .B(n12065), .Z(n28682) );
  NANDN U6546 ( .A(y[3228]), .B(x[3228]), .Z(n21466) );
  NANDN U6547 ( .A(y[3229]), .B(x[3229]), .Z(n21473) );
  NAND U6548 ( .A(n21466), .B(n21473), .Z(n24066) );
  NANDN U6549 ( .A(x[3227]), .B(y[3227]), .Z(n12070) );
  NANDN U6550 ( .A(x[3228]), .B(y[3228]), .Z(n12069) );
  AND U6551 ( .A(n12070), .B(n12069), .Z(n28681) );
  NANDN U6552 ( .A(x[3223]), .B(y[3223]), .Z(n21451) );
  NANDN U6553 ( .A(x[3224]), .B(y[3224]), .Z(n12073) );
  AND U6554 ( .A(n21451), .B(n12073), .Z(n28678) );
  NANDN U6555 ( .A(y[3222]), .B(x[3222]), .Z(n12074) );
  NANDN U6556 ( .A(y[3223]), .B(x[3223]), .Z(n21455) );
  NAND U6557 ( .A(n12074), .B(n21455), .Z(n28676) );
  NANDN U6558 ( .A(x[3221]), .B(y[3221]), .Z(n21445) );
  NANDN U6559 ( .A(x[3222]), .B(y[3222]), .Z(n21452) );
  AND U6560 ( .A(n21445), .B(n21452), .Z(n28675) );
  NANDN U6561 ( .A(y[3220]), .B(x[3220]), .Z(n12076) );
  NANDN U6562 ( .A(y[3221]), .B(x[3221]), .Z(n12075) );
  NAND U6563 ( .A(n12076), .B(n12075), .Z(n28674) );
  NANDN U6564 ( .A(y[3218]), .B(x[3218]), .Z(n12078) );
  NANDN U6565 ( .A(y[3219]), .B(x[3219]), .Z(n12077) );
  NAND U6566 ( .A(n12078), .B(n12077), .Z(n24069) );
  NANDN U6567 ( .A(y[3216]), .B(x[3216]), .Z(n12082) );
  NANDN U6568 ( .A(y[3217]), .B(x[3217]), .Z(n12079) );
  AND U6569 ( .A(n12082), .B(n12079), .Z(n28672) );
  NANDN U6570 ( .A(x[3215]), .B(y[3215]), .Z(n21431) );
  NANDN U6571 ( .A(x[3216]), .B(y[3216]), .Z(n12081) );
  NAND U6572 ( .A(n21431), .B(n12081), .Z(n28671) );
  NANDN U6573 ( .A(y[3214]), .B(x[3214]), .Z(n12084) );
  NANDN U6574 ( .A(y[3215]), .B(x[3215]), .Z(n12083) );
  AND U6575 ( .A(n12084), .B(n12083), .Z(n24070) );
  NANDN U6576 ( .A(x[3209]), .B(y[3209]), .Z(n12088) );
  NANDN U6577 ( .A(x[3210]), .B(y[3210]), .Z(n21417) );
  NAND U6578 ( .A(n12088), .B(n21417), .Z(n28666) );
  NANDN U6579 ( .A(y[3209]), .B(x[3209]), .Z(n21413) );
  ANDN U6580 ( .B(x[3208]), .A(y[3208]), .Z(n21407) );
  ANDN U6581 ( .B(n21413), .A(n21407), .Z(n28665) );
  NANDN U6582 ( .A(x[3207]), .B(y[3207]), .Z(n12090) );
  NANDN U6583 ( .A(x[3208]), .B(y[3208]), .Z(n12089) );
  NAND U6584 ( .A(n12090), .B(n12089), .Z(n28664) );
  NANDN U6585 ( .A(y[3206]), .B(x[3206]), .Z(n21401) );
  ANDN U6586 ( .B(x[3207]), .A(y[3207]), .Z(n21408) );
  ANDN U6587 ( .B(n21401), .A(n21408), .Z(n28663) );
  NANDN U6588 ( .A(x[3205]), .B(y[3205]), .Z(n12092) );
  NANDN U6589 ( .A(x[3206]), .B(y[3206]), .Z(n12091) );
  NAND U6590 ( .A(n12092), .B(n12091), .Z(n28662) );
  NANDN U6591 ( .A(x[3203]), .B(y[3203]), .Z(n12094) );
  NANDN U6592 ( .A(x[3204]), .B(y[3204]), .Z(n12093) );
  AND U6593 ( .A(n12094), .B(n12093), .Z(n28660) );
  NANDN U6594 ( .A(y[3202]), .B(x[3202]), .Z(n21389) );
  NANDN U6595 ( .A(y[3203]), .B(x[3203]), .Z(n21396) );
  NAND U6596 ( .A(n21389), .B(n21396), .Z(n28659) );
  NANDN U6597 ( .A(x[3201]), .B(y[3201]), .Z(n12096) );
  NANDN U6598 ( .A(x[3202]), .B(y[3202]), .Z(n12095) );
  AND U6599 ( .A(n12096), .B(n12095), .Z(n28658) );
  NANDN U6600 ( .A(y[3200]), .B(x[3200]), .Z(n12098) );
  NANDN U6601 ( .A(y[3201]), .B(x[3201]), .Z(n21390) );
  NAND U6602 ( .A(n12098), .B(n21390), .Z(n28657) );
  ANDN U6603 ( .B(x[3197]), .A(y[3197]), .Z(n21379) );
  NANDN U6604 ( .A(y[3196]), .B(x[3196]), .Z(n21372) );
  NANDN U6605 ( .A(n21379), .B(n21372), .Z(n28655) );
  NANDN U6606 ( .A(x[3195]), .B(y[3195]), .Z(n12104) );
  NANDN U6607 ( .A(x[3196]), .B(y[3196]), .Z(n12103) );
  AND U6608 ( .A(n12104), .B(n12103), .Z(n24075) );
  NANDN U6609 ( .A(y[3194]), .B(x[3194]), .Z(n21366) );
  NANDN U6610 ( .A(y[3195]), .B(x[3195]), .Z(n21373) );
  NAND U6611 ( .A(n21366), .B(n21373), .Z(n28653) );
  NANDN U6612 ( .A(x[3193]), .B(y[3193]), .Z(n12106) );
  NANDN U6613 ( .A(x[3194]), .B(y[3194]), .Z(n12105) );
  AND U6614 ( .A(n12106), .B(n12105), .Z(n28652) );
  NANDN U6615 ( .A(y[3192]), .B(x[3192]), .Z(n21360) );
  NANDN U6616 ( .A(y[3193]), .B(x[3193]), .Z(n21367) );
  NAND U6617 ( .A(n21360), .B(n21367), .Z(n28651) );
  NANDN U6618 ( .A(x[3189]), .B(y[3189]), .Z(n12110) );
  NANDN U6619 ( .A(x[3190]), .B(y[3190]), .Z(n12109) );
  NAND U6620 ( .A(n12110), .B(n12109), .Z(n28649) );
  NANDN U6621 ( .A(y[3188]), .B(x[3188]), .Z(n21348) );
  NANDN U6622 ( .A(y[3189]), .B(x[3189]), .Z(n21355) );
  AND U6623 ( .A(n21348), .B(n21355), .Z(n28648) );
  NANDN U6624 ( .A(x[3187]), .B(y[3187]), .Z(n12112) );
  NANDN U6625 ( .A(x[3188]), .B(y[3188]), .Z(n12111) );
  NAND U6626 ( .A(n12112), .B(n12111), .Z(n28647) );
  NANDN U6627 ( .A(y[3186]), .B(x[3186]), .Z(n21342) );
  NANDN U6628 ( .A(y[3187]), .B(x[3187]), .Z(n21349) );
  AND U6629 ( .A(n21342), .B(n21349), .Z(n28646) );
  NANDN U6630 ( .A(x[3183]), .B(y[3183]), .Z(n12116) );
  NANDN U6631 ( .A(x[3184]), .B(y[3184]), .Z(n12115) );
  NAND U6632 ( .A(n12116), .B(n12115), .Z(n24078) );
  NANDN U6633 ( .A(y[3182]), .B(x[3182]), .Z(n21330) );
  NANDN U6634 ( .A(y[3183]), .B(x[3183]), .Z(n21337) );
  AND U6635 ( .A(n21330), .B(n21337), .Z(n28644) );
  NANDN U6636 ( .A(x[3179]), .B(y[3179]), .Z(n12120) );
  NANDN U6637 ( .A(x[3180]), .B(y[3180]), .Z(n12119) );
  NAND U6638 ( .A(n12120), .B(n12119), .Z(n28640) );
  NANDN U6639 ( .A(y[3176]), .B(x[3176]), .Z(n21312) );
  NANDN U6640 ( .A(y[3177]), .B(x[3177]), .Z(n21319) );
  NAND U6641 ( .A(n21312), .B(n21319), .Z(n28637) );
  NANDN U6642 ( .A(x[3175]), .B(y[3175]), .Z(n12124) );
  NANDN U6643 ( .A(x[3176]), .B(y[3176]), .Z(n12123) );
  AND U6644 ( .A(n12124), .B(n12123), .Z(n24080) );
  NANDN U6645 ( .A(y[3174]), .B(x[3174]), .Z(n21306) );
  NANDN U6646 ( .A(y[3175]), .B(x[3175]), .Z(n21313) );
  NAND U6647 ( .A(n21306), .B(n21313), .Z(n28636) );
  NANDN U6648 ( .A(x[3173]), .B(y[3173]), .Z(n21303) );
  NANDN U6649 ( .A(x[3174]), .B(y[3174]), .Z(n12125) );
  AND U6650 ( .A(n21303), .B(n12125), .Z(n28635) );
  NANDN U6651 ( .A(x[3171]), .B(y[3171]), .Z(n21297) );
  NANDN U6652 ( .A(x[3172]), .B(y[3172]), .Z(n21304) );
  AND U6653 ( .A(n21297), .B(n21304), .Z(n28633) );
  NANDN U6654 ( .A(y[3170]), .B(x[3170]), .Z(n12128) );
  NANDN U6655 ( .A(y[3171]), .B(x[3171]), .Z(n12127) );
  NAND U6656 ( .A(n12128), .B(n12127), .Z(n28632) );
  NANDN U6657 ( .A(x[3169]), .B(y[3169]), .Z(n21291) );
  NANDN U6658 ( .A(x[3170]), .B(y[3170]), .Z(n21298) );
  AND U6659 ( .A(n21291), .B(n21298), .Z(n24081) );
  NANDN U6660 ( .A(y[3166]), .B(x[3166]), .Z(n21281) );
  NANDN U6661 ( .A(y[3167]), .B(x[3167]), .Z(n12131) );
  NAND U6662 ( .A(n21281), .B(n12131), .Z(n28628) );
  ANDN U6663 ( .B(y[3164]), .A(x[3164]), .Z(n21276) );
  NANDN U6664 ( .A(x[3163]), .B(y[3163]), .Z(n21271) );
  NANDN U6665 ( .A(n21276), .B(n21271), .Z(n24084) );
  NANDN U6666 ( .A(y[3163]), .B(x[3163]), .Z(n12132) );
  ANDN U6667 ( .B(x[3162]), .A(y[3162]), .Z(n21267) );
  ANDN U6668 ( .B(n12132), .A(n21267), .Z(n28626) );
  ANDN U6669 ( .B(x[3160]), .A(y[3160]), .Z(n21261) );
  ANDN U6670 ( .B(x[3161]), .A(y[3161]), .Z(n21269) );
  NOR U6671 ( .A(n21261), .B(n21269), .Z(n28624) );
  ANDN U6672 ( .B(x[3158]), .A(y[3158]), .Z(n21252) );
  ANDN U6673 ( .B(x[3159]), .A(y[3159]), .Z(n21262) );
  NOR U6674 ( .A(n21252), .B(n21262), .Z(n28622) );
  NANDN U6675 ( .A(x[3157]), .B(y[3157]), .Z(n21249) );
  NANDN U6676 ( .A(x[3158]), .B(y[3158]), .Z(n21256) );
  NAND U6677 ( .A(n21249), .B(n21256), .Z(n28621) );
  ANDN U6678 ( .B(x[3156]), .A(y[3156]), .Z(n21245) );
  ANDN U6679 ( .B(x[3157]), .A(y[3157]), .Z(n21255) );
  NOR U6680 ( .A(n21245), .B(n21255), .Z(n28620) );
  NANDN U6681 ( .A(x[3155]), .B(y[3155]), .Z(n12136) );
  NANDN U6682 ( .A(x[3156]), .B(y[3156]), .Z(n21250) );
  NAND U6683 ( .A(n12136), .B(n21250), .Z(n28619) );
  ANDN U6684 ( .B(x[3154]), .A(y[3154]), .Z(n21239) );
  ANDN U6685 ( .B(x[3155]), .A(y[3155]), .Z(n21247) );
  NOR U6686 ( .A(n21239), .B(n21247), .Z(n28618) );
  NANDN U6687 ( .A(x[3153]), .B(y[3153]), .Z(n21235) );
  NANDN U6688 ( .A(x[3154]), .B(y[3154]), .Z(n12137) );
  NAND U6689 ( .A(n21235), .B(n12137), .Z(n24085) );
  NANDN U6690 ( .A(x[3151]), .B(y[3151]), .Z(n3972) );
  NANDN U6691 ( .A(x[3152]), .B(y[3152]), .Z(n21234) );
  AND U6692 ( .A(n3972), .B(n21234), .Z(n28616) );
  ANDN U6693 ( .B(x[3150]), .A(y[3150]), .Z(n21224) );
  NANDN U6694 ( .A(y[3151]), .B(x[3151]), .Z(n12139) );
  NANDN U6695 ( .A(n21224), .B(n12139), .Z(n28615) );
  NANDN U6696 ( .A(x[3150]), .B(y[3150]), .Z(n21227) );
  NANDN U6697 ( .A(x[3149]), .B(y[3149]), .Z(n3973) );
  NAND U6698 ( .A(n21227), .B(n3973), .Z(n28613) );
  NANDN U6699 ( .A(x[3147]), .B(y[3147]), .Z(n21216) );
  ANDN U6700 ( .B(y[3148]), .A(x[3148]), .Z(n21222) );
  ANDN U6701 ( .B(n21216), .A(n21222), .Z(n28611) );
  ANDN U6702 ( .B(x[3146]), .A(y[3146]), .Z(n21214) );
  NANDN U6703 ( .A(y[3147]), .B(x[3147]), .Z(n21220) );
  NANDN U6704 ( .A(n21214), .B(n21220), .Z(n24086) );
  NANDN U6705 ( .A(x[3143]), .B(y[3143]), .Z(n3975) );
  NANDN U6706 ( .A(x[3144]), .B(y[3144]), .Z(n3974) );
  AND U6707 ( .A(n3975), .B(n3974), .Z(n28608) );
  NANDN U6708 ( .A(y[3142]), .B(x[3142]), .Z(n3976) );
  ANDN U6709 ( .B(x[3143]), .A(y[3143]), .Z(n21207) );
  ANDN U6710 ( .B(n3976), .A(n21207), .Z(n28607) );
  NANDN U6711 ( .A(x[3141]), .B(y[3141]), .Z(n21201) );
  NANDN U6712 ( .A(x[3142]), .B(y[3142]), .Z(n21206) );
  NAND U6713 ( .A(n21201), .B(n21206), .Z(n28606) );
  NANDN U6714 ( .A(y[3141]), .B(x[3141]), .Z(n12140) );
  ANDN U6715 ( .B(x[3140]), .A(y[3140]), .Z(n21197) );
  ANDN U6716 ( .B(n12140), .A(n21197), .Z(n28605) );
  ANDN U6717 ( .B(y[3140]), .A(x[3140]), .Z(n21203) );
  NANDN U6718 ( .A(x[3139]), .B(y[3139]), .Z(n12141) );
  NANDN U6719 ( .A(n21203), .B(n12141), .Z(n28604) );
  ANDN U6720 ( .B(x[3138]), .A(y[3138]), .Z(n21191) );
  ANDN U6721 ( .B(x[3139]), .A(y[3139]), .Z(n21199) );
  NOR U6722 ( .A(n21191), .B(n21199), .Z(n28603) );
  NANDN U6723 ( .A(x[3137]), .B(y[3137]), .Z(n21187) );
  NANDN U6724 ( .A(x[3138]), .B(y[3138]), .Z(n12142) );
  NAND U6725 ( .A(n21187), .B(n12142), .Z(n28602) );
  ANDN U6726 ( .B(x[3136]), .A(y[3136]), .Z(n21182) );
  ANDN U6727 ( .B(x[3137]), .A(y[3137]), .Z(n21192) );
  NOR U6728 ( .A(n21182), .B(n21192), .Z(n28601) );
  ANDN U6729 ( .B(x[3134]), .A(y[3134]), .Z(n21175) );
  ANDN U6730 ( .B(x[3135]), .A(y[3135]), .Z(n21185) );
  NOR U6731 ( .A(n21175), .B(n21185), .Z(n28599) );
  NANDN U6732 ( .A(x[3133]), .B(y[3133]), .Z(n12143) );
  NANDN U6733 ( .A(x[3134]), .B(y[3134]), .Z(n21180) );
  NAND U6734 ( .A(n12143), .B(n21180), .Z(n28598) );
  ANDN U6735 ( .B(x[3132]), .A(y[3132]), .Z(n21169) );
  ANDN U6736 ( .B(x[3133]), .A(y[3133]), .Z(n21177) );
  NOR U6737 ( .A(n21169), .B(n21177), .Z(n28597) );
  NANDN U6738 ( .A(x[3131]), .B(y[3131]), .Z(n21165) );
  NANDN U6739 ( .A(x[3132]), .B(y[3132]), .Z(n12144) );
  NAND U6740 ( .A(n21165), .B(n12144), .Z(n28596) );
  ANDN U6741 ( .B(x[3130]), .A(y[3130]), .Z(n21160) );
  ANDN U6742 ( .B(x[3131]), .A(y[3131]), .Z(n21170) );
  NOR U6743 ( .A(n21160), .B(n21170), .Z(n28595) );
  ANDN U6744 ( .B(x[3128]), .A(y[3128]), .Z(n21153) );
  ANDN U6745 ( .B(x[3129]), .A(y[3129]), .Z(n21163) );
  NOR U6746 ( .A(n21153), .B(n21163), .Z(n28593) );
  NANDN U6747 ( .A(x[3127]), .B(y[3127]), .Z(n12145) );
  NANDN U6748 ( .A(x[3128]), .B(y[3128]), .Z(n21158) );
  NAND U6749 ( .A(n12145), .B(n21158), .Z(n28592) );
  ANDN U6750 ( .B(x[3126]), .A(y[3126]), .Z(n21147) );
  ANDN U6751 ( .B(x[3127]), .A(y[3127]), .Z(n21155) );
  NOR U6752 ( .A(n21147), .B(n21155), .Z(n28591) );
  ANDN U6753 ( .B(x[3124]), .A(y[3124]), .Z(n21138) );
  ANDN U6754 ( .B(x[3125]), .A(y[3125]), .Z(n21148) );
  NOR U6755 ( .A(n21138), .B(n21148), .Z(n28590) );
  NANDN U6756 ( .A(x[3123]), .B(y[3123]), .Z(n21135) );
  NANDN U6757 ( .A(x[3124]), .B(y[3124]), .Z(n21142) );
  NAND U6758 ( .A(n21135), .B(n21142), .Z(n28589) );
  ANDN U6759 ( .B(x[3120]), .A(y[3120]), .Z(n21125) );
  ANDN U6760 ( .B(x[3121]), .A(y[3121]), .Z(n21133) );
  OR U6761 ( .A(n21125), .B(n21133), .Z(n24090) );
  NANDN U6762 ( .A(x[3119]), .B(y[3119]), .Z(n21121) );
  NANDN U6763 ( .A(x[3120]), .B(y[3120]), .Z(n12148) );
  AND U6764 ( .A(n21121), .B(n12148), .Z(n28586) );
  NANDN U6765 ( .A(x[3115]), .B(y[3115]), .Z(n12149) );
  NANDN U6766 ( .A(x[3116]), .B(y[3116]), .Z(n21114) );
  AND U6767 ( .A(n12149), .B(n21114), .Z(n28583) );
  ANDN U6768 ( .B(x[3114]), .A(y[3114]), .Z(n21103) );
  ANDN U6769 ( .B(x[3115]), .A(y[3115]), .Z(n21111) );
  OR U6770 ( .A(n21103), .B(n21111), .Z(n28582) );
  NANDN U6771 ( .A(x[3113]), .B(y[3113]), .Z(n21099) );
  NANDN U6772 ( .A(x[3114]), .B(y[3114]), .Z(n12150) );
  AND U6773 ( .A(n21099), .B(n12150), .Z(n28581) );
  ANDN U6774 ( .B(x[3112]), .A(y[3112]), .Z(n21094) );
  ANDN U6775 ( .B(x[3113]), .A(y[3113]), .Z(n21104) );
  OR U6776 ( .A(n21094), .B(n21104), .Z(n28580) );
  ANDN U6777 ( .B(x[3110]), .A(y[3110]), .Z(n21087) );
  ANDN U6778 ( .B(x[3111]), .A(y[3111]), .Z(n21097) );
  OR U6779 ( .A(n21087), .B(n21097), .Z(n24093) );
  ANDN U6780 ( .B(x[3108]), .A(y[3108]), .Z(n21081) );
  ANDN U6781 ( .B(x[3109]), .A(y[3109]), .Z(n21089) );
  NOR U6782 ( .A(n21081), .B(n21089), .Z(n28578) );
  NANDN U6783 ( .A(x[3107]), .B(y[3107]), .Z(n21077) );
  NANDN U6784 ( .A(x[3108]), .B(y[3108]), .Z(n12152) );
  NAND U6785 ( .A(n21077), .B(n12152), .Z(n28577) );
  ANDN U6786 ( .B(x[3106]), .A(y[3106]), .Z(n21072) );
  ANDN U6787 ( .B(x[3107]), .A(y[3107]), .Z(n21082) );
  NOR U6788 ( .A(n21072), .B(n21082), .Z(n28576) );
  ANDN U6789 ( .B(x[3104]), .A(y[3104]), .Z(n21065) );
  ANDN U6790 ( .B(x[3105]), .A(y[3105]), .Z(n21075) );
  NOR U6791 ( .A(n21065), .B(n21075), .Z(n28574) );
  ANDN U6792 ( .B(x[3102]), .A(y[3102]), .Z(n21059) );
  ANDN U6793 ( .B(x[3103]), .A(y[3103]), .Z(n21067) );
  NOR U6794 ( .A(n21059), .B(n21067), .Z(n28572) );
  NANDN U6795 ( .A(x[3101]), .B(y[3101]), .Z(n21055) );
  NANDN U6796 ( .A(x[3102]), .B(y[3102]), .Z(n12154) );
  NAND U6797 ( .A(n21055), .B(n12154), .Z(n28571) );
  ANDN U6798 ( .B(x[3100]), .A(y[3100]), .Z(n21050) );
  ANDN U6799 ( .B(x[3101]), .A(y[3101]), .Z(n21060) );
  NOR U6800 ( .A(n21050), .B(n21060), .Z(n28570) );
  NANDN U6801 ( .A(x[3099]), .B(y[3099]), .Z(n21047) );
  NANDN U6802 ( .A(x[3100]), .B(y[3100]), .Z(n21054) );
  NAND U6803 ( .A(n21047), .B(n21054), .Z(n28569) );
  ANDN U6804 ( .B(x[3098]), .A(y[3098]), .Z(n21043) );
  ANDN U6805 ( .B(x[3099]), .A(y[3099]), .Z(n21053) );
  NOR U6806 ( .A(n21043), .B(n21053), .Z(n28568) );
  ANDN U6807 ( .B(x[3096]), .A(y[3096]), .Z(n21037) );
  ANDN U6808 ( .B(x[3097]), .A(y[3097]), .Z(n21045) );
  NOR U6809 ( .A(n21037), .B(n21045), .Z(n28566) );
  NANDN U6810 ( .A(x[3095]), .B(y[3095]), .Z(n21033) );
  NANDN U6811 ( .A(x[3096]), .B(y[3096]), .Z(n12156) );
  NAND U6812 ( .A(n21033), .B(n12156), .Z(n28565) );
  ANDN U6813 ( .B(x[3094]), .A(y[3094]), .Z(n21028) );
  ANDN U6814 ( .B(x[3095]), .A(y[3095]), .Z(n21038) );
  NOR U6815 ( .A(n21028), .B(n21038), .Z(n28564) );
  ANDN U6816 ( .B(x[3092]), .A(y[3092]), .Z(n12157) );
  ANDN U6817 ( .B(x[3093]), .A(y[3093]), .Z(n21031) );
  NOR U6818 ( .A(n12157), .B(n21031), .Z(n28562) );
  NANDN U6819 ( .A(x[3092]), .B(y[3092]), .Z(n12160) );
  NANDN U6820 ( .A(x[3091]), .B(y[3091]), .Z(n3977) );
  NAND U6821 ( .A(n12160), .B(n3977), .Z(n12161) );
  NANDN U6822 ( .A(x[3089]), .B(y[3089]), .Z(n21017) );
  NANDN U6823 ( .A(x[3090]), .B(y[3090]), .Z(n12162) );
  AND U6824 ( .A(n21017), .B(n12162), .Z(n28558) );
  ANDN U6825 ( .B(x[3088]), .A(y[3088]), .Z(n21015) );
  ANDN U6826 ( .B(x[3089]), .A(y[3089]), .Z(n21020) );
  OR U6827 ( .A(n21015), .B(n21020), .Z(n28557) );
  NANDN U6828 ( .A(x[3087]), .B(y[3087]), .Z(n3979) );
  ANDN U6829 ( .B(y[3088]), .A(x[3088]), .Z(n3978) );
  ANDN U6830 ( .B(n3979), .A(n3978), .Z(n28556) );
  NANDN U6831 ( .A(y[3086]), .B(x[3086]), .Z(n21010) );
  NANDN U6832 ( .A(y[3087]), .B(x[3087]), .Z(n3980) );
  NAND U6833 ( .A(n21010), .B(n3980), .Z(n28555) );
  NANDN U6834 ( .A(y[3084]), .B(x[3084]), .Z(n3982) );
  NANDN U6835 ( .A(y[3085]), .B(x[3085]), .Z(n3981) );
  AND U6836 ( .A(n3982), .B(n3981), .Z(n28553) );
  NANDN U6837 ( .A(y[3082]), .B(x[3082]), .Z(n3983) );
  NANDN U6838 ( .A(y[3083]), .B(x[3083]), .Z(n21003) );
  AND U6839 ( .A(n3983), .B(n21003), .Z(n28551) );
  ANDN U6840 ( .B(y[3081]), .A(x[3081]), .Z(n28550) );
  NANDN U6841 ( .A(x[3082]), .B(y[3082]), .Z(n21004) );
  NANDN U6842 ( .A(n28550), .B(n21004), .Z(n10102) );
  NANDN U6843 ( .A(y[3080]), .B(x[3080]), .Z(n20994) );
  NANDN U6844 ( .A(y[3081]), .B(x[3081]), .Z(n21001) );
  AND U6845 ( .A(n20994), .B(n21001), .Z(n28549) );
  NANDN U6846 ( .A(y[3078]), .B(x[3078]), .Z(n3984) );
  NANDN U6847 ( .A(y[3079]), .B(x[3079]), .Z(n28547) );
  AND U6848 ( .A(n3984), .B(n28547), .Z(n10098) );
  XNOR U6849 ( .A(x[3078]), .B(y[3078]), .Z(n12165) );
  ANDN U6850 ( .B(x[3077]), .A(y[3077]), .Z(n12164) );
  NANDN U6851 ( .A(x[3075]), .B(y[3075]), .Z(n12167) );
  ANDN U6852 ( .B(y[3076]), .A(x[3076]), .Z(n20989) );
  ANDN U6853 ( .B(n12167), .A(n20989), .Z(n28542) );
  NANDN U6854 ( .A(y[3074]), .B(x[3074]), .Z(n12168) );
  NANDN U6855 ( .A(y[3075]), .B(x[3075]), .Z(n20985) );
  NAND U6856 ( .A(n12168), .B(n20985), .Z(n28541) );
  NANDN U6857 ( .A(x[3073]), .B(y[3073]), .Z(n12170) );
  NANDN U6858 ( .A(x[3074]), .B(y[3074]), .Z(n12166) );
  AND U6859 ( .A(n12170), .B(n12166), .Z(n28540) );
  NANDN U6860 ( .A(x[3071]), .B(y[3071]), .Z(n12172) );
  NANDN U6861 ( .A(x[3072]), .B(y[3072]), .Z(n12171) );
  AND U6862 ( .A(n12172), .B(n12171), .Z(n28538) );
  ANDN U6863 ( .B(x[3070]), .A(y[3070]), .Z(n20970) );
  NANDN U6864 ( .A(y[3071]), .B(x[3071]), .Z(n20976) );
  NANDN U6865 ( .A(n20970), .B(n20976), .Z(n28537) );
  NANDN U6866 ( .A(x[3070]), .B(y[3070]), .Z(n28536) );
  ANDN U6867 ( .B(x[3069]), .A(y[3069]), .Z(n20971) );
  ANDN U6868 ( .B(x[3068]), .A(y[3068]), .Z(n20966) );
  NANDN U6869 ( .A(x[3069]), .B(y[3069]), .Z(n3987) );
  NAND U6870 ( .A(n20966), .B(n3987), .Z(n3985) );
  NANDN U6871 ( .A(n20971), .B(n3985), .Z(n28535) );
  NANDN U6872 ( .A(x[3068]), .B(y[3068]), .Z(n3986) );
  AND U6873 ( .A(n3987), .B(n3986), .Z(n28534) );
  NANDN U6874 ( .A(x[3067]), .B(y[3067]), .Z(n12174) );
  NANDN U6875 ( .A(y[3067]), .B(x[3067]), .Z(n24096) );
  ANDN U6876 ( .B(x[3066]), .A(y[3066]), .Z(n20963) );
  ANDN U6877 ( .B(n24096), .A(n20963), .Z(n28533) );
  NANDN U6878 ( .A(x[3065]), .B(y[3065]), .Z(n28532) );
  ANDN U6879 ( .B(y[3066]), .A(x[3066]), .Z(n12173) );
  ANDN U6880 ( .B(n28532), .A(n12173), .Z(n10081) );
  ANDN U6881 ( .B(x[3058]), .A(y[3058]), .Z(n20947) );
  ANDN U6882 ( .B(x[3059]), .A(y[3059]), .Z(n20954) );
  OR U6883 ( .A(n20947), .B(n20954), .Z(n24100) );
  NANDN U6884 ( .A(x[3057]), .B(y[3057]), .Z(n20943) );
  NANDN U6885 ( .A(x[3058]), .B(y[3058]), .Z(n12176) );
  AND U6886 ( .A(n20943), .B(n12176), .Z(n28527) );
  ANDN U6887 ( .B(x[3056]), .A(y[3056]), .Z(n12177) );
  NANDN U6888 ( .A(x[3056]), .B(y[3056]), .Z(n28525) );
  NANDN U6889 ( .A(x[3055]), .B(y[3055]), .Z(n12179) );
  NAND U6890 ( .A(n28525), .B(n12179), .Z(n28523) );
  NANDN U6891 ( .A(y[3052]), .B(x[3052]), .Z(n12182) );
  ANDN U6892 ( .B(x[3053]), .A(y[3053]), .Z(n20938) );
  ANDN U6893 ( .B(n12182), .A(n20938), .Z(n28521) );
  NANDN U6894 ( .A(y[3050]), .B(x[3050]), .Z(n12185) );
  NANDN U6895 ( .A(y[3051]), .B(x[3051]), .Z(n12181) );
  AND U6896 ( .A(n12185), .B(n12181), .Z(n28519) );
  NANDN U6897 ( .A(x[3049]), .B(y[3049]), .Z(n20922) );
  NANDN U6898 ( .A(x[3050]), .B(y[3050]), .Z(n12184) );
  NAND U6899 ( .A(n20922), .B(n12184), .Z(n28518) );
  NANDN U6900 ( .A(y[3048]), .B(x[3048]), .Z(n20918) );
  NANDN U6901 ( .A(y[3049]), .B(x[3049]), .Z(n12186) );
  AND U6902 ( .A(n20918), .B(n12186), .Z(n24102) );
  NANDN U6903 ( .A(y[3047]), .B(x[3047]), .Z(n20919) );
  ANDN U6904 ( .B(x[3046]), .A(y[3046]), .Z(n20914) );
  ANDN U6905 ( .B(n20919), .A(n20914), .Z(n28517) );
  NANDN U6906 ( .A(x[3046]), .B(y[3046]), .Z(n28513) );
  ANDN U6907 ( .B(x[3044]), .A(y[3044]), .Z(n20910) );
  ANDN U6908 ( .B(x[3045]), .A(y[3045]), .Z(n28514) );
  OR U6909 ( .A(n20910), .B(n28514), .Z(n28511) );
  NANDN U6910 ( .A(x[3043]), .B(y[3043]), .Z(n28510) );
  NANDN U6911 ( .A(y[3042]), .B(x[3042]), .Z(n3989) );
  NANDN U6912 ( .A(y[3043]), .B(x[3043]), .Z(n3988) );
  NAND U6913 ( .A(n3989), .B(n3988), .Z(n28509) );
  NANDN U6914 ( .A(x[3041]), .B(y[3041]), .Z(n3991) );
  NANDN U6915 ( .A(x[3042]), .B(y[3042]), .Z(n3990) );
  AND U6916 ( .A(n3991), .B(n3990), .Z(n28508) );
  NANDN U6917 ( .A(y[3040]), .B(x[3040]), .Z(n3993) );
  ANDN U6918 ( .B(x[3041]), .A(y[3041]), .Z(n3992) );
  ANDN U6919 ( .B(n3993), .A(n3992), .Z(n28507) );
  ANDN U6920 ( .B(y[3037]), .A(x[3037]), .Z(n12193) );
  ANDN U6921 ( .B(y[3038]), .A(x[3038]), .Z(n12190) );
  NOR U6922 ( .A(n12193), .B(n12190), .Z(n10035) );
  NANDN U6923 ( .A(x[3035]), .B(y[3035]), .Z(n20892) );
  NANDN U6924 ( .A(x[3036]), .B(y[3036]), .Z(n12194) );
  AND U6925 ( .A(n20892), .B(n12194), .Z(n28503) );
  NANDN U6926 ( .A(y[3034]), .B(x[3034]), .Z(n20888) );
  ANDN U6927 ( .B(x[3035]), .A(y[3035]), .Z(n24108) );
  ANDN U6928 ( .B(n20888), .A(n24108), .Z(n10031) );
  NANDN U6929 ( .A(y[3032]), .B(x[3032]), .Z(n28500) );
  NANDN U6930 ( .A(x[3031]), .B(y[3031]), .Z(n12198) );
  NANDN U6931 ( .A(x[3032]), .B(y[3032]), .Z(n12196) );
  NAND U6932 ( .A(n12198), .B(n12196), .Z(n28499) );
  NANDN U6933 ( .A(y[3028]), .B(x[3028]), .Z(n12204) );
  NANDN U6934 ( .A(y[3029]), .B(x[3029]), .Z(n12201) );
  NAND U6935 ( .A(n12204), .B(n12201), .Z(n28496) );
  NANDN U6936 ( .A(x[3027]), .B(y[3027]), .Z(n12206) );
  NANDN U6937 ( .A(x[3028]), .B(y[3028]), .Z(n12203) );
  AND U6938 ( .A(n12206), .B(n12203), .Z(n24109) );
  ANDN U6939 ( .B(x[3026]), .A(y[3026]), .Z(n20870) );
  NANDN U6940 ( .A(y[3027]), .B(x[3027]), .Z(n12205) );
  NANDN U6941 ( .A(n20870), .B(n12205), .Z(n28495) );
  NANDN U6942 ( .A(x[3025]), .B(y[3025]), .Z(n20868) );
  NANDN U6943 ( .A(x[3026]), .B(y[3026]), .Z(n12207) );
  AND U6944 ( .A(n20868), .B(n12207), .Z(n28494) );
  ANDN U6945 ( .B(x[3024]), .A(y[3024]), .Z(n20866) );
  ANDN U6946 ( .B(x[3025]), .A(y[3025]), .Z(n20873) );
  OR U6947 ( .A(n20866), .B(n20873), .Z(n28493) );
  NANDN U6948 ( .A(x[3024]), .B(y[3024]), .Z(n28490) );
  ANDN U6949 ( .B(x[3022]), .A(y[3022]), .Z(n20860) );
  ANDN U6950 ( .B(x[3023]), .A(y[3023]), .Z(n28491) );
  OR U6951 ( .A(n20860), .B(n28491), .Z(n28489) );
  NANDN U6952 ( .A(x[3021]), .B(y[3021]), .Z(n28488) );
  ANDN U6953 ( .B(x[3020]), .A(y[3020]), .Z(n20854) );
  ANDN U6954 ( .B(x[3021]), .A(y[3021]), .Z(n20861) );
  NOR U6955 ( .A(n20854), .B(n20861), .Z(n28487) );
  NANDN U6956 ( .A(x[3019]), .B(y[3019]), .Z(n20850) );
  NANDN U6957 ( .A(x[3020]), .B(y[3020]), .Z(n12210) );
  NAND U6958 ( .A(n20850), .B(n12210), .Z(n24110) );
  NANDN U6959 ( .A(y[3018]), .B(x[3018]), .Z(n12211) );
  ANDN U6960 ( .B(x[3019]), .A(y[3019]), .Z(n20855) );
  ANDN U6961 ( .B(n12211), .A(n20855), .Z(n28485) );
  ANDN U6962 ( .B(y[3018]), .A(x[3018]), .Z(n20849) );
  XNOR U6963 ( .A(x[3016]), .B(y[3016]), .Z(n20844) );
  NANDN U6964 ( .A(y[3015]), .B(x[3015]), .Z(n20843) );
  ANDN U6965 ( .B(x[3014]), .A(y[3014]), .Z(n12214) );
  ANDN U6966 ( .B(n20843), .A(n12214), .Z(n10003) );
  XNOR U6967 ( .A(x[3012]), .B(y[3012]), .Z(n20834) );
  NANDN U6968 ( .A(x[3011]), .B(y[3011]), .Z(n20830) );
  AND U6969 ( .A(n20834), .B(n20830), .Z(n9997) );
  ANDN U6970 ( .B(x[3010]), .A(y[3010]), .Z(n12215) );
  NANDN U6971 ( .A(x[3010]), .B(y[3010]), .Z(n20831) );
  NANDN U6972 ( .A(y[3008]), .B(x[3008]), .Z(n12219) );
  NANDN U6973 ( .A(y[3006]), .B(x[3006]), .Z(n20821) );
  ANDN U6974 ( .B(y[3005]), .A(x[3005]), .Z(n12221) );
  NANDN U6975 ( .A(x[3004]), .B(y[3004]), .Z(n12222) );
  NANDN U6976 ( .A(x[3003]), .B(y[3003]), .Z(n28468) );
  AND U6977 ( .A(n12222), .B(n28468), .Z(n9981) );
  NANDN U6978 ( .A(y[3002]), .B(x[3002]), .Z(n12224) );
  NANDN U6979 ( .A(y[3003]), .B(x[3003]), .Z(n12223) );
  NAND U6980 ( .A(n12224), .B(n12223), .Z(n28467) );
  NANDN U6981 ( .A(x[3001]), .B(y[3001]), .Z(n12225) );
  NANDN U6982 ( .A(x[2999]), .B(y[2999]), .Z(n20811) );
  NANDN U6983 ( .A(y[2999]), .B(x[2999]), .Z(n3995) );
  NANDN U6984 ( .A(y[2998]), .B(x[2998]), .Z(n3994) );
  AND U6985 ( .A(n3995), .B(n3994), .Z(n4002) );
  NANDN U6986 ( .A(x[2997]), .B(y[2997]), .Z(n3997) );
  NANDN U6987 ( .A(x[2998]), .B(y[2998]), .Z(n3996) );
  AND U6988 ( .A(n3997), .B(n3996), .Z(n4006) );
  NANDN U6989 ( .A(y[2997]), .B(x[2997]), .Z(n3999) );
  NANDN U6990 ( .A(y[2996]), .B(x[2996]), .Z(n3998) );
  NAND U6991 ( .A(n3999), .B(n3998), .Z(n4000) );
  NAND U6992 ( .A(n4006), .B(n4000), .Z(n4001) );
  NAND U6993 ( .A(n4002), .B(n4001), .Z(n20810) );
  NANDN U6994 ( .A(x[2996]), .B(y[2996]), .Z(n4004) );
  NANDN U6995 ( .A(x[2995]), .B(y[2995]), .Z(n4003) );
  AND U6996 ( .A(n4004), .B(n4003), .Z(n4005) );
  AND U6997 ( .A(n4006), .B(n4005), .Z(n12229) );
  NANDN U6998 ( .A(y[2992]), .B(x[2992]), .Z(n20798) );
  NANDN U6999 ( .A(y[2993]), .B(x[2993]), .Z(n20806) );
  NAND U7000 ( .A(n20798), .B(n20806), .Z(n24114) );
  NANDN U7001 ( .A(x[2991]), .B(y[2991]), .Z(n12230) );
  ANDN U7002 ( .B(y[2992]), .A(x[2992]), .Z(n20801) );
  ANDN U7003 ( .B(n12230), .A(n20801), .Z(n28458) );
  ANDN U7004 ( .B(x[2990]), .A(y[2990]), .Z(n12231) );
  NANDN U7005 ( .A(y[2991]), .B(x[2991]), .Z(n24118) );
  NANDN U7006 ( .A(x[2990]), .B(y[2990]), .Z(n24115) );
  NANDN U7007 ( .A(x[2989]), .B(y[2989]), .Z(n20791) );
  NAND U7008 ( .A(n24115), .B(n20791), .Z(n28455) );
  NANDN U7009 ( .A(y[2986]), .B(x[2986]), .Z(n20780) );
  ANDN U7010 ( .B(x[2987]), .A(y[2987]), .Z(n20789) );
  ANDN U7011 ( .B(n20780), .A(n20789), .Z(n28452) );
  NANDN U7012 ( .A(x[2983]), .B(y[2983]), .Z(n12238) );
  NANDN U7013 ( .A(x[2984]), .B(y[2984]), .Z(n12236) );
  NAND U7014 ( .A(n12238), .B(n12236), .Z(n24120) );
  NANDN U7015 ( .A(y[2983]), .B(x[2983]), .Z(n20775) );
  ANDN U7016 ( .B(x[2982]), .A(y[2982]), .Z(n20769) );
  ANDN U7017 ( .B(n20775), .A(n20769), .Z(n28450) );
  NANDN U7018 ( .A(x[2981]), .B(y[2981]), .Z(n20765) );
  NANDN U7019 ( .A(x[2982]), .B(y[2982]), .Z(n12237) );
  NAND U7020 ( .A(n20765), .B(n12237), .Z(n28449) );
  ANDN U7021 ( .B(x[2980]), .A(y[2980]), .Z(n20763) );
  ANDN U7022 ( .B(x[2981]), .A(y[2981]), .Z(n20770) );
  NOR U7023 ( .A(n20763), .B(n20770), .Z(n28448) );
  NANDN U7024 ( .A(x[2978]), .B(y[2978]), .Z(n12239) );
  ANDN U7025 ( .B(y[2977]), .A(x[2977]), .Z(n24121) );
  ANDN U7026 ( .B(n12239), .A(n24121), .Z(n9947) );
  NANDN U7027 ( .A(y[2974]), .B(x[2974]), .Z(n4008) );
  NANDN U7028 ( .A(y[2975]), .B(x[2975]), .Z(n4007) );
  NAND U7029 ( .A(n4008), .B(n4007), .Z(n20752) );
  NANDN U7030 ( .A(x[2974]), .B(y[2974]), .Z(n4010) );
  NANDN U7031 ( .A(x[2973]), .B(y[2973]), .Z(n4009) );
  AND U7032 ( .A(n4010), .B(n4009), .Z(n12248) );
  NANDN U7033 ( .A(x[2969]), .B(y[2969]), .Z(n12253) );
  ANDN U7034 ( .B(y[2970]), .A(x[2970]), .Z(n12252) );
  ANDN U7035 ( .B(n12253), .A(n12252), .Z(n28436) );
  ANDN U7036 ( .B(x[2968]), .A(y[2968]), .Z(n12254) );
  ANDN U7037 ( .B(x[2969]), .A(y[2969]), .Z(n28435) );
  NOR U7038 ( .A(n12254), .B(n28435), .Z(n9933) );
  NANDN U7039 ( .A(x[2965]), .B(y[2965]), .Z(n20736) );
  NANDN U7040 ( .A(x[2966]), .B(y[2966]), .Z(n12256) );
  NAND U7041 ( .A(n20736), .B(n12256), .Z(n28432) );
  NANDN U7042 ( .A(y[2964]), .B(x[2964]), .Z(n9925) );
  NANDN U7043 ( .A(x[2963]), .B(y[2963]), .Z(n28426) );
  XOR U7044 ( .A(x[2964]), .B(y[2964]), .Z(n20732) );
  ANDN U7045 ( .B(n28426), .A(n20732), .Z(n9923) );
  NANDN U7046 ( .A(x[2961]), .B(y[2961]), .Z(n4011) );
  ANDN U7047 ( .B(y[2962]), .A(x[2962]), .Z(n12260) );
  ANDN U7048 ( .B(n4011), .A(n12260), .Z(n28423) );
  ANDN U7049 ( .B(x[2960]), .A(y[2960]), .Z(n20725) );
  NANDN U7050 ( .A(y[2961]), .B(x[2961]), .Z(n12259) );
  NANDN U7051 ( .A(n20725), .B(n12259), .Z(n24123) );
  NANDN U7052 ( .A(x[2959]), .B(y[2959]), .Z(n12262) );
  NANDN U7053 ( .A(x[2960]), .B(y[2960]), .Z(n20727) );
  AND U7054 ( .A(n12262), .B(n20727), .Z(n24124) );
  NANDN U7055 ( .A(x[2957]), .B(y[2957]), .Z(n12263) );
  NANDN U7056 ( .A(x[2958]), .B(y[2958]), .Z(n24126) );
  AND U7057 ( .A(n12263), .B(n24126), .Z(n9915) );
  NANDN U7058 ( .A(y[2956]), .B(x[2956]), .Z(n28420) );
  NANDN U7059 ( .A(y[2957]), .B(x[2957]), .Z(n28422) );
  NAND U7060 ( .A(n28420), .B(n28422), .Z(n9913) );
  ANDN U7061 ( .B(x[2954]), .A(y[2954]), .Z(n20710) );
  NANDN U7062 ( .A(y[2955]), .B(x[2955]), .Z(n12265) );
  NANDN U7063 ( .A(n20710), .B(n12265), .Z(n28418) );
  NANDN U7064 ( .A(x[2953]), .B(y[2953]), .Z(n4012) );
  ANDN U7065 ( .B(y[2954]), .A(x[2954]), .Z(n12266) );
  ANDN U7066 ( .B(n4012), .A(n12266), .Z(n28417) );
  ANDN U7067 ( .B(x[2952]), .A(y[2952]), .Z(n20704) );
  NANDN U7068 ( .A(y[2953]), .B(x[2953]), .Z(n4013) );
  NANDN U7069 ( .A(n20704), .B(n4013), .Z(n28416) );
  NANDN U7070 ( .A(x[2951]), .B(y[2951]), .Z(n12267) );
  NANDN U7071 ( .A(x[2952]), .B(y[2952]), .Z(n24127) );
  AND U7072 ( .A(n12267), .B(n24127), .Z(n9906) );
  ANDN U7073 ( .B(x[2948]), .A(y[2948]), .Z(n20693) );
  ANDN U7074 ( .B(x[2949]), .A(y[2949]), .Z(n20699) );
  OR U7075 ( .A(n20693), .B(n20699), .Z(n28410) );
  NANDN U7076 ( .A(x[2947]), .B(y[2947]), .Z(n20689) );
  NANDN U7077 ( .A(x[2948]), .B(y[2948]), .Z(n12269) );
  AND U7078 ( .A(n20689), .B(n12269), .Z(n28409) );
  ANDN U7079 ( .B(x[2947]), .A(y[2947]), .Z(n24131) );
  NANDN U7080 ( .A(x[2946]), .B(y[2946]), .Z(n20691) );
  IV U7081 ( .A(n20691), .Z(n24129) );
  ANDN U7082 ( .B(y[2945]), .A(x[2945]), .Z(n20686) );
  NOR U7083 ( .A(n24129), .B(n20686), .Z(n28408) );
  ANDN U7084 ( .B(x[2944]), .A(y[2944]), .Z(n28407) );
  NANDN U7085 ( .A(x[2943]), .B(y[2943]), .Z(n4014) );
  ANDN U7086 ( .B(y[2944]), .A(x[2944]), .Z(n12273) );
  ANDN U7087 ( .B(n4014), .A(n12273), .Z(n28406) );
  NANDN U7088 ( .A(y[2942]), .B(x[2942]), .Z(n12276) );
  NANDN U7089 ( .A(y[2943]), .B(x[2943]), .Z(n12272) );
  AND U7090 ( .A(n12276), .B(n12272), .Z(n28405) );
  NANDN U7091 ( .A(x[2941]), .B(y[2941]), .Z(n12277) );
  NANDN U7092 ( .A(x[2942]), .B(y[2942]), .Z(n20680) );
  NAND U7093 ( .A(n12277), .B(n20680), .Z(n28404) );
  NANDN U7094 ( .A(y[2940]), .B(x[2940]), .Z(n12280) );
  NANDN U7095 ( .A(y[2941]), .B(x[2941]), .Z(n12275) );
  AND U7096 ( .A(n12280), .B(n12275), .Z(n28403) );
  ANDN U7097 ( .B(y[2939]), .A(x[2939]), .Z(n20671) );
  NANDN U7098 ( .A(x[2940]), .B(y[2940]), .Z(n12278) );
  NANDN U7099 ( .A(n20671), .B(n12278), .Z(n28402) );
  NANDN U7100 ( .A(y[2938]), .B(x[2938]), .Z(n12281) );
  NANDN U7101 ( .A(y[2939]), .B(x[2939]), .Z(n12279) );
  AND U7102 ( .A(n12281), .B(n12279), .Z(n24132) );
  NANDN U7103 ( .A(y[2935]), .B(x[2935]), .Z(n24134) );
  ANDN U7104 ( .B(x[2934]), .A(y[2934]), .Z(n20660) );
  ANDN U7105 ( .B(n24134), .A(n20660), .Z(n28399) );
  NANDN U7106 ( .A(x[2934]), .B(y[2934]), .Z(n12284) );
  ANDN U7107 ( .B(y[2933]), .A(x[2933]), .Z(n12285) );
  ANDN U7108 ( .B(n12284), .A(n12285), .Z(n9883) );
  NANDN U7109 ( .A(x[2931]), .B(y[2931]), .Z(n28395) );
  NANDN U7110 ( .A(x[2929]), .B(y[2929]), .Z(n20645) );
  NANDN U7111 ( .A(x[2930]), .B(y[2930]), .Z(n28393) );
  AND U7112 ( .A(n20645), .B(n28393), .Z(n9877) );
  ANDN U7113 ( .B(x[2928]), .A(y[2928]), .Z(n9875) );
  ANDN U7114 ( .B(y[2927]), .A(x[2927]), .Z(n28388) );
  ANDN U7115 ( .B(x[2924]), .A(y[2924]), .Z(n9867) );
  ANDN U7116 ( .B(x[2925]), .A(y[2925]), .Z(n24138) );
  NANDN U7117 ( .A(x[2923]), .B(y[2923]), .Z(n12292) );
  XNOR U7118 ( .A(x[2924]), .B(y[2924]), .Z(n12291) );
  NANDN U7119 ( .A(y[2923]), .B(x[2923]), .Z(n12290) );
  ANDN U7120 ( .B(x[2922]), .A(y[2922]), .Z(n20629) );
  ANDN U7121 ( .B(n12290), .A(n20629), .Z(n9862) );
  NANDN U7122 ( .A(y[2921]), .B(x[2921]), .Z(n28381) );
  NANDN U7123 ( .A(y[2919]), .B(x[2919]), .Z(n12293) );
  ANDN U7124 ( .B(x[2918]), .A(y[2918]), .Z(n12297) );
  ANDN U7125 ( .B(n12293), .A(n12297), .Z(n9855) );
  NANDN U7126 ( .A(y[2917]), .B(x[2917]), .Z(n12298) );
  NANDN U7127 ( .A(x[2916]), .B(y[2916]), .Z(n4016) );
  NANDN U7128 ( .A(x[2917]), .B(y[2917]), .Z(n4015) );
  NAND U7129 ( .A(n4016), .B(n4015), .Z(n28376) );
  NANDN U7130 ( .A(x[2915]), .B(y[2915]), .Z(n4024) );
  XNOR U7131 ( .A(x[2915]), .B(y[2915]), .Z(n4018) );
  NANDN U7132 ( .A(y[2914]), .B(x[2914]), .Z(n4017) );
  NAND U7133 ( .A(n4018), .B(n4017), .Z(n4019) );
  NAND U7134 ( .A(n4024), .B(n4019), .Z(n4021) );
  NANDN U7135 ( .A(y[2916]), .B(x[2916]), .Z(n4020) );
  AND U7136 ( .A(n4021), .B(n4020), .Z(n24140) );
  NANDN U7137 ( .A(x[2914]), .B(y[2914]), .Z(n4023) );
  NANDN U7138 ( .A(x[2913]), .B(y[2913]), .Z(n4022) );
  AND U7139 ( .A(n4023), .B(n4022), .Z(n4025) );
  AND U7140 ( .A(n4025), .B(n4024), .Z(n12302) );
  NANDN U7141 ( .A(y[2913]), .B(x[2913]), .Z(n12299) );
  NANDN U7142 ( .A(y[2912]), .B(x[2912]), .Z(n4026) );
  AND U7143 ( .A(n12299), .B(n4026), .Z(n24142) );
  ANDN U7144 ( .B(y[2910]), .A(x[2910]), .Z(n12304) );
  NANDN U7145 ( .A(y[2908]), .B(x[2908]), .Z(n20610) );
  NANDN U7146 ( .A(y[2909]), .B(x[2909]), .Z(n12306) );
  AND U7147 ( .A(n20610), .B(n12306), .Z(n28369) );
  ANDN U7148 ( .B(y[2907]), .A(x[2907]), .Z(n20607) );
  ANDN U7149 ( .B(x[2906]), .A(y[2906]), .Z(n9839) );
  XNOR U7150 ( .A(x[2906]), .B(y[2906]), .Z(n12308) );
  ANDN U7151 ( .B(x[2905]), .A(y[2905]), .Z(n12307) );
  NANDN U7152 ( .A(y[2902]), .B(x[2902]), .Z(n4027) );
  NANDN U7153 ( .A(y[2903]), .B(x[2903]), .Z(n12309) );
  AND U7154 ( .A(n4027), .B(n12309), .Z(n9831) );
  ANDN U7155 ( .B(y[2901]), .A(x[2901]), .Z(n12312) );
  NANDN U7156 ( .A(y[2901]), .B(x[2901]), .Z(n12311) );
  NANDN U7157 ( .A(x[2899]), .B(y[2899]), .Z(n20589) );
  NANDN U7158 ( .A(x[2900]), .B(y[2900]), .Z(n12313) );
  NAND U7159 ( .A(n20589), .B(n12313), .Z(n24144) );
  XNOR U7160 ( .A(x[2898]), .B(y[2898]), .Z(n12315) );
  NANDN U7161 ( .A(x[2897]), .B(y[2897]), .Z(n28352) );
  NANDN U7162 ( .A(x[2894]), .B(y[2894]), .Z(n20579) );
  ANDN U7163 ( .B(y[2893]), .A(x[2893]), .Z(n20574) );
  ANDN U7164 ( .B(n20579), .A(n20574), .Z(n28350) );
  ANDN U7165 ( .B(x[2893]), .A(y[2893]), .Z(n12317) );
  NANDN U7166 ( .A(y[2892]), .B(x[2892]), .Z(n12320) );
  NANDN U7167 ( .A(n12317), .B(n12320), .Z(n28349) );
  NANDN U7168 ( .A(x[2890]), .B(y[2890]), .Z(n12322) );
  NANDN U7169 ( .A(x[2889]), .B(y[2889]), .Z(n12323) );
  AND U7170 ( .A(n12322), .B(n12323), .Z(n9809) );
  NANDN U7171 ( .A(x[2888]), .B(y[2888]), .Z(n12324) );
  ANDN U7172 ( .B(y[2887]), .A(x[2887]), .Z(n20563) );
  ANDN U7173 ( .B(n12324), .A(n20563), .Z(n28341) );
  NANDN U7174 ( .A(y[2886]), .B(x[2886]), .Z(n20558) );
  NANDN U7175 ( .A(y[2887]), .B(x[2887]), .Z(n20565) );
  NAND U7176 ( .A(n20558), .B(n20565), .Z(n24147) );
  XNOR U7177 ( .A(x[2884]), .B(y[2884]), .Z(n12331) );
  NANDN U7178 ( .A(x[2883]), .B(y[2883]), .Z(n20553) );
  AND U7179 ( .A(n12331), .B(n20553), .Z(n9798) );
  ANDN U7180 ( .B(x[2883]), .A(y[2883]), .Z(n12330) );
  NANDN U7181 ( .A(y[2882]), .B(x[2882]), .Z(n28335) );
  NANDN U7182 ( .A(y[2881]), .B(x[2881]), .Z(n28333) );
  NANDN U7183 ( .A(y[2880]), .B(x[2880]), .Z(n4028) );
  AND U7184 ( .A(n28333), .B(n4028), .Z(n9791) );
  ANDN U7185 ( .B(y[2879]), .A(x[2879]), .Z(n24148) );
  NANDN U7186 ( .A(x[2877]), .B(y[2877]), .Z(n20539) );
  NANDN U7187 ( .A(x[2878]), .B(y[2878]), .Z(n20546) );
  AND U7188 ( .A(n20539), .B(n20546), .Z(n28328) );
  ANDN U7189 ( .B(x[2877]), .A(y[2877]), .Z(n20544) );
  NANDN U7190 ( .A(y[2876]), .B(x[2876]), .Z(n12335) );
  NANDN U7191 ( .A(n20544), .B(n12335), .Z(n28327) );
  NANDN U7192 ( .A(x[2875]), .B(y[2875]), .Z(n12336) );
  NANDN U7193 ( .A(x[2876]), .B(y[2876]), .Z(n20538) );
  NAND U7194 ( .A(n12336), .B(n20538), .Z(n28326) );
  NANDN U7195 ( .A(y[2874]), .B(x[2874]), .Z(n12338) );
  NANDN U7196 ( .A(y[2875]), .B(x[2875]), .Z(n12334) );
  AND U7197 ( .A(n12338), .B(n12334), .Z(n24149) );
  NANDN U7198 ( .A(x[2873]), .B(y[2873]), .Z(n20528) );
  NANDN U7199 ( .A(x[2874]), .B(y[2874]), .Z(n12337) );
  NAND U7200 ( .A(n20528), .B(n12337), .Z(n28325) );
  NANDN U7201 ( .A(y[2872]), .B(x[2872]), .Z(n12341) );
  NANDN U7202 ( .A(y[2873]), .B(x[2873]), .Z(n12339) );
  AND U7203 ( .A(n12341), .B(n12339), .Z(n28324) );
  ANDN U7204 ( .B(y[2871]), .A(x[2871]), .Z(n20523) );
  NANDN U7205 ( .A(x[2872]), .B(y[2872]), .Z(n20529) );
  NANDN U7206 ( .A(n20523), .B(n20529), .Z(n28323) );
  NANDN U7207 ( .A(y[2868]), .B(x[2868]), .Z(n28318) );
  NANDN U7208 ( .A(y[2869]), .B(x[2869]), .Z(n28320) );
  NAND U7209 ( .A(n28318), .B(n28320), .Z(n9775) );
  NANDN U7210 ( .A(x[2867]), .B(y[2867]), .Z(n28317) );
  NANDN U7211 ( .A(y[2866]), .B(x[2866]), .Z(n12347) );
  NANDN U7212 ( .A(y[2867]), .B(x[2867]), .Z(n12345) );
  NAND U7213 ( .A(n12347), .B(n12345), .Z(n28316) );
  NANDN U7214 ( .A(x[2866]), .B(y[2866]), .Z(n20514) );
  ANDN U7215 ( .B(y[2865]), .A(x[2865]), .Z(n20510) );
  ANDN U7216 ( .B(n20514), .A(n20510), .Z(n28315) );
  NANDN U7217 ( .A(y[2864]), .B(x[2864]), .Z(n12348) );
  NANDN U7218 ( .A(y[2865]), .B(x[2865]), .Z(n12346) );
  NAND U7219 ( .A(n12348), .B(n12346), .Z(n28314) );
  NANDN U7220 ( .A(x[2863]), .B(y[2863]), .Z(n20505) );
  ANDN U7221 ( .B(y[2864]), .A(x[2864]), .Z(n28312) );
  ANDN U7222 ( .B(n20505), .A(n28312), .Z(n9768) );
  ANDN U7223 ( .B(x[2862]), .A(y[2862]), .Z(n12349) );
  NANDN U7224 ( .A(y[2860]), .B(x[2860]), .Z(n12353) );
  ANDN U7225 ( .B(y[2859]), .A(x[2859]), .Z(n12355) );
  NANDN U7226 ( .A(y[2859]), .B(x[2859]), .Z(n12354) );
  XOR U7227 ( .A(x[2858]), .B(y[2858]), .Z(n12356) );
  ANDN U7228 ( .B(y[2854]), .A(x[2854]), .Z(n20493) );
  NANDN U7229 ( .A(x[2853]), .B(y[2853]), .Z(n12361) );
  NANDN U7230 ( .A(n20493), .B(n12361), .Z(n28302) );
  NANDN U7231 ( .A(y[2852]), .B(x[2852]), .Z(n12363) );
  NANDN U7232 ( .A(y[2853]), .B(x[2853]), .Z(n20486) );
  AND U7233 ( .A(n12363), .B(n20486), .Z(n28301) );
  NANDN U7234 ( .A(x[2851]), .B(y[2851]), .Z(n12365) );
  NANDN U7235 ( .A(x[2852]), .B(y[2852]), .Z(n12362) );
  NAND U7236 ( .A(n12365), .B(n12362), .Z(n28300) );
  NANDN U7237 ( .A(y[2850]), .B(x[2850]), .Z(n12366) );
  NANDN U7238 ( .A(y[2851]), .B(x[2851]), .Z(n12364) );
  AND U7239 ( .A(n12366), .B(n12364), .Z(n28299) );
  NANDN U7240 ( .A(x[2850]), .B(y[2850]), .Z(n28298) );
  NANDN U7241 ( .A(x[2849]), .B(y[2849]), .Z(n9741) );
  XNOR U7242 ( .A(x[2849]), .B(y[2849]), .Z(n4030) );
  NANDN U7243 ( .A(y[2848]), .B(x[2848]), .Z(n4029) );
  NAND U7244 ( .A(n4030), .B(n4029), .Z(n4031) );
  NAND U7245 ( .A(n9741), .B(n4031), .Z(n28297) );
  NANDN U7246 ( .A(y[2846]), .B(x[2846]), .Z(n4032) );
  NANDN U7247 ( .A(y[2847]), .B(x[2847]), .Z(n20474) );
  AND U7248 ( .A(n4032), .B(n20474), .Z(n28292) );
  NANDN U7249 ( .A(y[2844]), .B(x[2844]), .Z(n12368) );
  NANDN U7250 ( .A(y[2845]), .B(x[2845]), .Z(n12367) );
  NAND U7251 ( .A(n12368), .B(n12367), .Z(n28288) );
  ANDN U7252 ( .B(y[2843]), .A(x[2843]), .Z(n20464) );
  ANDN U7253 ( .B(y[2844]), .A(x[2844]), .Z(n20470) );
  NOR U7254 ( .A(n20464), .B(n20470), .Z(n28287) );
  NANDN U7255 ( .A(y[2842]), .B(x[2842]), .Z(n20460) );
  NANDN U7256 ( .A(y[2843]), .B(x[2843]), .Z(n12369) );
  NAND U7257 ( .A(n20460), .B(n12369), .Z(n28285) );
  NANDN U7258 ( .A(x[2841]), .B(y[2841]), .Z(n12370) );
  NANDN U7259 ( .A(x[2842]), .B(y[2842]), .Z(n20465) );
  AND U7260 ( .A(n12370), .B(n20465), .Z(n9732) );
  ANDN U7261 ( .B(x[2841]), .A(y[2841]), .Z(n20459) );
  NANDN U7262 ( .A(y[2840]), .B(x[2840]), .Z(n9729) );
  NANDN U7263 ( .A(x[2839]), .B(y[2839]), .Z(n28274) );
  NANDN U7264 ( .A(y[2839]), .B(x[2839]), .Z(n12373) );
  ANDN U7265 ( .B(y[2837]), .A(x[2837]), .Z(n20451) );
  NANDN U7266 ( .A(x[2838]), .B(y[2838]), .Z(n12374) );
  NANDN U7267 ( .A(n20451), .B(n12374), .Z(n28271) );
  NANDN U7268 ( .A(y[2836]), .B(x[2836]), .Z(n4033) );
  NANDN U7269 ( .A(y[2837]), .B(x[2837]), .Z(n28269) );
  AND U7270 ( .A(n4033), .B(n28269), .Z(n9722) );
  NANDN U7271 ( .A(x[2835]), .B(y[2835]), .Z(n28259) );
  NANDN U7272 ( .A(y[2835]), .B(x[2835]), .Z(n12376) );
  NANDN U7273 ( .A(x[2833]), .B(y[2833]), .Z(n20444) );
  NANDN U7274 ( .A(x[2834]), .B(y[2834]), .Z(n12377) );
  NAND U7275 ( .A(n20444), .B(n12377), .Z(n28260) );
  NANDN U7276 ( .A(y[2833]), .B(x[2833]), .Z(n12378) );
  NANDN U7277 ( .A(y[2832]), .B(x[2832]), .Z(n20440) );
  AND U7278 ( .A(n12378), .B(n20440), .Z(n9715) );
  ANDN U7279 ( .B(y[2832]), .A(x[2832]), .Z(n28255) );
  NANDN U7280 ( .A(y[2831]), .B(x[2831]), .Z(n20441) );
  ANDN U7281 ( .B(y[2829]), .A(x[2829]), .Z(n20435) );
  NANDN U7282 ( .A(x[2828]), .B(y[2828]), .Z(n20436) );
  NANDN U7283 ( .A(y[2828]), .B(x[2828]), .Z(n4035) );
  NANDN U7284 ( .A(y[2827]), .B(x[2827]), .Z(n4034) );
  AND U7285 ( .A(n4035), .B(n4034), .Z(n20434) );
  NANDN U7286 ( .A(y[2826]), .B(x[2826]), .Z(n12383) );
  NANDN U7287 ( .A(x[2827]), .B(y[2827]), .Z(n9702) );
  ANDN U7288 ( .B(y[2825]), .A(x[2825]), .Z(n4036) );
  NANDN U7289 ( .A(y[2824]), .B(x[2824]), .Z(n12384) );
  NANDN U7290 ( .A(y[2825]), .B(x[2825]), .Z(n28249) );
  AND U7291 ( .A(n12384), .B(n28249), .Z(n28247) );
  OR U7292 ( .A(n4036), .B(n28247), .Z(n9701) );
  NANDN U7293 ( .A(x[2824]), .B(y[2824]), .Z(n4037) );
  ANDN U7294 ( .B(n4037), .A(n4036), .Z(n28248) );
  NANDN U7295 ( .A(x[2823]), .B(y[2823]), .Z(n28246) );
  AND U7296 ( .A(n28248), .B(n28246), .Z(n9699) );
  NANDN U7297 ( .A(x[2822]), .B(y[2822]), .Z(n20424) );
  ANDN U7298 ( .B(y[2821]), .A(x[2821]), .Z(n20420) );
  ANDN U7299 ( .B(n20424), .A(n20420), .Z(n28244) );
  NANDN U7300 ( .A(y[2820]), .B(x[2820]), .Z(n12388) );
  NANDN U7301 ( .A(y[2821]), .B(x[2821]), .Z(n12386) );
  NAND U7302 ( .A(n12388), .B(n12386), .Z(n28243) );
  NANDN U7303 ( .A(x[2818]), .B(y[2818]), .Z(n20415) );
  ANDN U7304 ( .B(y[2817]), .A(x[2817]), .Z(n28238) );
  ANDN U7305 ( .B(n20415), .A(n28238), .Z(n9689) );
  NANDN U7306 ( .A(y[2816]), .B(x[2816]), .Z(n28237) );
  NANDN U7307 ( .A(x[2815]), .B(y[2815]), .Z(n12391) );
  ANDN U7308 ( .B(y[2816]), .A(x[2816]), .Z(n20411) );
  ANDN U7309 ( .B(n12391), .A(n20411), .Z(n28236) );
  ANDN U7310 ( .B(x[2814]), .A(y[2814]), .Z(n12392) );
  ANDN U7311 ( .B(y[2814]), .A(x[2814]), .Z(n12390) );
  NANDN U7312 ( .A(y[2813]), .B(x[2813]), .Z(n12393) );
  ANDN U7313 ( .B(y[2811]), .A(x[2811]), .Z(n28231) );
  NANDN U7314 ( .A(y[2810]), .B(x[2810]), .Z(n12395) );
  NANDN U7315 ( .A(x[2809]), .B(y[2809]), .Z(n12397) );
  NANDN U7316 ( .A(x[2810]), .B(y[2810]), .Z(n20399) );
  AND U7317 ( .A(n12397), .B(n20399), .Z(n28229) );
  NANDN U7318 ( .A(y[2808]), .B(x[2808]), .Z(n28227) );
  NANDN U7319 ( .A(x[2807]), .B(y[2807]), .Z(n20390) );
  NANDN U7320 ( .A(x[2808]), .B(y[2808]), .Z(n12398) );
  NAND U7321 ( .A(n20390), .B(n12398), .Z(n28224) );
  NANDN U7322 ( .A(y[2807]), .B(x[2807]), .Z(n12399) );
  ANDN U7323 ( .B(x[2806]), .A(y[2806]), .Z(n20386) );
  ANDN U7324 ( .B(n12399), .A(n20386), .Z(n28223) );
  NANDN U7325 ( .A(y[2804]), .B(x[2804]), .Z(n12400) );
  ANDN U7326 ( .B(x[2805]), .A(y[2805]), .Z(n20388) );
  ANDN U7327 ( .B(n12400), .A(n20388), .Z(n28222) );
  ANDN U7328 ( .B(y[2804]), .A(x[2804]), .Z(n20381) );
  NANDN U7329 ( .A(y[2803]), .B(x[2803]), .Z(n24158) );
  ANDN U7330 ( .B(x[2802]), .A(y[2802]), .Z(n20377) );
  ANDN U7331 ( .B(n24158), .A(n20377), .Z(n28221) );
  NANDN U7332 ( .A(x[2801]), .B(y[2801]), .Z(n28220) );
  ANDN U7333 ( .B(x[2801]), .A(y[2801]), .Z(n20372) );
  NANDN U7334 ( .A(y[2800]), .B(x[2800]), .Z(n4038) );
  NANDN U7335 ( .A(n20372), .B(n4038), .Z(n20367) );
  ANDN U7336 ( .B(x[2798]), .A(y[2798]), .Z(n20364) );
  ANDN U7337 ( .B(x[2799]), .A(y[2799]), .Z(n20370) );
  NOR U7338 ( .A(n20364), .B(n20370), .Z(n28216) );
  ANDN U7339 ( .B(y[2798]), .A(x[2798]), .Z(n12403) );
  NANDN U7340 ( .A(y[2797]), .B(x[2797]), .Z(n24161) );
  NANDN U7341 ( .A(y[2796]), .B(x[2796]), .Z(n9655) );
  NANDN U7342 ( .A(x[2795]), .B(y[2795]), .Z(n28210) );
  NANDN U7343 ( .A(y[2795]), .B(x[2795]), .Z(n12405) );
  ANDN U7344 ( .B(y[2794]), .A(x[2794]), .Z(n20358) );
  NANDN U7345 ( .A(x[2793]), .B(y[2793]), .Z(n12406) );
  NANDN U7346 ( .A(n20358), .B(n12406), .Z(n24162) );
  XNOR U7347 ( .A(x[2792]), .B(y[2792]), .Z(n12408) );
  ANDN U7348 ( .B(y[2790]), .A(x[2790]), .Z(n20349) );
  NANDN U7349 ( .A(x[2789]), .B(y[2789]), .Z(n12409) );
  NANDN U7350 ( .A(n20349), .B(n12409), .Z(n24166) );
  NANDN U7351 ( .A(y[2788]), .B(x[2788]), .Z(n4039) );
  NANDN U7352 ( .A(y[2789]), .B(x[2789]), .Z(n28206) );
  AND U7353 ( .A(n4039), .B(n28206), .Z(n9640) );
  ANDN U7354 ( .B(y[2787]), .A(x[2787]), .Z(n24167) );
  NANDN U7355 ( .A(x[2785]), .B(y[2785]), .Z(n12412) );
  ANDN U7356 ( .B(y[2786]), .A(x[2786]), .Z(n20341) );
  ANDN U7357 ( .B(n12412), .A(n20341), .Z(n28202) );
  NANDN U7358 ( .A(y[2784]), .B(x[2784]), .Z(n20331) );
  NANDN U7359 ( .A(y[2785]), .B(x[2785]), .Z(n20338) );
  NAND U7360 ( .A(n20331), .B(n20338), .Z(n24168) );
  NANDN U7361 ( .A(x[2783]), .B(y[2783]), .Z(n12414) );
  NANDN U7362 ( .A(x[2784]), .B(y[2784]), .Z(n12413) );
  NAND U7363 ( .A(n12414), .B(n12413), .Z(n28200) );
  NANDN U7364 ( .A(y[2782]), .B(x[2782]), .Z(n20326) );
  NANDN U7365 ( .A(y[2783]), .B(x[2783]), .Z(n20332) );
  AND U7366 ( .A(n20326), .B(n20332), .Z(n28199) );
  NANDN U7367 ( .A(x[2781]), .B(y[2781]), .Z(n20323) );
  NANDN U7368 ( .A(x[2782]), .B(y[2782]), .Z(n12415) );
  NAND U7369 ( .A(n20323), .B(n12415), .Z(n28198) );
  NANDN U7370 ( .A(y[2780]), .B(x[2780]), .Z(n20320) );
  NANDN U7371 ( .A(y[2781]), .B(x[2781]), .Z(n28196) );
  AND U7372 ( .A(n20320), .B(n28196), .Z(n28195) );
  ANDN U7373 ( .B(y[2779]), .A(x[2779]), .Z(n28194) );
  ANDN U7374 ( .B(y[2780]), .A(x[2780]), .Z(n28197) );
  NANDN U7375 ( .A(y[2778]), .B(x[2778]), .Z(n12416) );
  NANDN U7376 ( .A(y[2779]), .B(x[2779]), .Z(n20322) );
  AND U7377 ( .A(n12416), .B(n20322), .Z(n28193) );
  NANDN U7378 ( .A(x[2775]), .B(y[2775]), .Z(n4041) );
  NANDN U7379 ( .A(x[2776]), .B(y[2776]), .Z(n4040) );
  NAND U7380 ( .A(n4041), .B(n4040), .Z(n12422) );
  NANDN U7381 ( .A(y[2775]), .B(x[2775]), .Z(n12420) );
  NANDN U7382 ( .A(y[2774]), .B(x[2774]), .Z(n4042) );
  AND U7383 ( .A(n12420), .B(n4042), .Z(n28190) );
  ANDN U7384 ( .B(y[2774]), .A(x[2774]), .Z(n12421) );
  NANDN U7385 ( .A(y[2772]), .B(x[2772]), .Z(n12423) );
  NANDN U7386 ( .A(y[2773]), .B(x[2773]), .Z(n20310) );
  NAND U7387 ( .A(n12423), .B(n20310), .Z(n28188) );
  ANDN U7388 ( .B(y[2771]), .A(x[2771]), .Z(n20302) );
  ANDN U7389 ( .B(y[2772]), .A(x[2772]), .Z(n20308) );
  NOR U7390 ( .A(n20302), .B(n20308), .Z(n28187) );
  ANDN U7391 ( .B(x[2770]), .A(y[2770]), .Z(n9616) );
  XOR U7392 ( .A(x[2770]), .B(y[2770]), .Z(n12424) );
  NANDN U7393 ( .A(y[2768]), .B(x[2768]), .Z(n24170) );
  NANDN U7394 ( .A(y[2769]), .B(x[2769]), .Z(n12425) );
  NANDN U7395 ( .A(x[2767]), .B(y[2767]), .Z(n20293) );
  NANDN U7396 ( .A(x[2768]), .B(y[2768]), .Z(n12427) );
  NAND U7397 ( .A(n20293), .B(n12427), .Z(n24171) );
  ANDN U7398 ( .B(x[2766]), .A(y[2766]), .Z(n20289) );
  NANDN U7399 ( .A(y[2767]), .B(x[2767]), .Z(n12428) );
  NANDN U7400 ( .A(n20289), .B(n12428), .Z(n28179) );
  NANDN U7401 ( .A(x[2765]), .B(y[2765]), .Z(n20285) );
  ANDN U7402 ( .B(y[2766]), .A(x[2766]), .Z(n20295) );
  ANDN U7403 ( .B(n20285), .A(n20295), .Z(n28178) );
  ANDN U7404 ( .B(x[2765]), .A(y[2765]), .Z(n20291) );
  NANDN U7405 ( .A(y[2764]), .B(x[2764]), .Z(n20283) );
  NANDN U7406 ( .A(n20291), .B(n20283), .Z(n28177) );
  NANDN U7407 ( .A(x[2764]), .B(y[2764]), .Z(n20287) );
  ANDN U7408 ( .B(y[2763]), .A(x[2763]), .Z(n20281) );
  ANDN U7409 ( .B(n20287), .A(n20281), .Z(n28176) );
  NANDN U7410 ( .A(x[2760]), .B(y[2760]), .Z(n4044) );
  NANDN U7411 ( .A(x[2759]), .B(y[2759]), .Z(n4043) );
  AND U7412 ( .A(n4044), .B(n4043), .Z(n12432) );
  NANDN U7413 ( .A(y[2758]), .B(x[2758]), .Z(n4045) );
  ANDN U7414 ( .B(x[2759]), .A(y[2759]), .Z(n12429) );
  ANDN U7415 ( .B(n4045), .A(n12429), .Z(n12434) );
  NANDN U7416 ( .A(y[2754]), .B(x[2754]), .Z(n4046) );
  NANDN U7417 ( .A(y[2755]), .B(x[2755]), .Z(n20270) );
  AND U7418 ( .A(n4046), .B(n20270), .Z(n12436) );
  NANDN U7419 ( .A(y[2752]), .B(x[2752]), .Z(n9581) );
  NANDN U7420 ( .A(y[2750]), .B(x[2750]), .Z(n28164) );
  NANDN U7421 ( .A(y[2748]), .B(x[2748]), .Z(n4047) );
  NANDN U7422 ( .A(y[2749]), .B(x[2749]), .Z(n28162) );
  AND U7423 ( .A(n4047), .B(n28162), .Z(n9574) );
  NANDN U7424 ( .A(x[2747]), .B(y[2747]), .Z(n28159) );
  NANDN U7425 ( .A(x[2746]), .B(y[2746]), .Z(n12443) );
  ANDN U7426 ( .B(y[2745]), .A(x[2745]), .Z(n20253) );
  ANDN U7427 ( .B(n12443), .A(n20253), .Z(n24172) );
  ANDN U7428 ( .B(x[2745]), .A(y[2745]), .Z(n12444) );
  ANDN U7429 ( .B(x[2744]), .A(y[2744]), .Z(n4048) );
  NOR U7430 ( .A(n12444), .B(n4048), .Z(n9567) );
  XNOR U7431 ( .A(x[2744]), .B(y[2744]), .Z(n20249) );
  NANDN U7432 ( .A(y[2742]), .B(x[2742]), .Z(n28155) );
  NANDN U7433 ( .A(y[2740]), .B(x[2740]), .Z(n28151) );
  ANDN U7434 ( .B(x[2741]), .A(y[2741]), .Z(n28156) );
  ANDN U7435 ( .B(n28151), .A(n28156), .Z(n9559) );
  NANDN U7436 ( .A(x[2739]), .B(y[2739]), .Z(n24176) );
  NANDN U7437 ( .A(y[2738]), .B(x[2738]), .Z(n12449) );
  ANDN U7438 ( .B(x[2739]), .A(y[2739]), .Z(n20241) );
  ANDN U7439 ( .B(n12449), .A(n20241), .Z(n24177) );
  ANDN U7440 ( .B(y[2738]), .A(x[2738]), .Z(n12448) );
  NANDN U7441 ( .A(x[2737]), .B(y[2737]), .Z(n12451) );
  ANDN U7442 ( .B(x[2736]), .A(y[2736]), .Z(n20235) );
  NANDN U7443 ( .A(y[2737]), .B(x[2737]), .Z(n24178) );
  NANDN U7444 ( .A(n20235), .B(n24178), .Z(n28149) );
  NANDN U7445 ( .A(y[2734]), .B(x[2734]), .Z(n12452) );
  ANDN U7446 ( .B(x[2735]), .A(y[2735]), .Z(n20233) );
  ANDN U7447 ( .B(n12452), .A(n20233), .Z(n28147) );
  NANDN U7448 ( .A(x[2734]), .B(y[2734]), .Z(n28146) );
  NANDN U7449 ( .A(y[2732]), .B(x[2732]), .Z(n20224) );
  NANDN U7450 ( .A(y[2733]), .B(x[2733]), .Z(n12453) );
  NAND U7451 ( .A(n20224), .B(n12453), .Z(n24181) );
  NANDN U7452 ( .A(x[2731]), .B(y[2731]), .Z(n20220) );
  NANDN U7453 ( .A(x[2732]), .B(y[2732]), .Z(n28145) );
  AND U7454 ( .A(n20220), .B(n28145), .Z(n9545) );
  ANDN U7455 ( .B(x[2731]), .A(y[2731]), .Z(n28144) );
  NANDN U7456 ( .A(x[2730]), .B(y[2730]), .Z(n20221) );
  NANDN U7457 ( .A(y[2729]), .B(x[2729]), .Z(n12455) );
  ANDN U7458 ( .B(x[2728]), .A(y[2728]), .Z(n28139) );
  ANDN U7459 ( .B(n12455), .A(n28139), .Z(n9539) );
  ANDN U7460 ( .B(x[2726]), .A(y[2726]), .Z(n20209) );
  ANDN U7461 ( .B(x[2727]), .A(y[2727]), .Z(n20214) );
  NOR U7462 ( .A(n20209), .B(n20214), .Z(n28138) );
  NANDN U7463 ( .A(x[2725]), .B(y[2725]), .Z(n20203) );
  NANDN U7464 ( .A(x[2726]), .B(y[2726]), .Z(n24183) );
  NAND U7465 ( .A(n20203), .B(n24183), .Z(n28137) );
  NANDN U7466 ( .A(y[2725]), .B(x[2725]), .Z(n20206) );
  NANDN U7467 ( .A(x[2723]), .B(y[2723]), .Z(n20195) );
  NANDN U7468 ( .A(x[2724]), .B(y[2724]), .Z(n20204) );
  NAND U7469 ( .A(n20195), .B(n20204), .Z(n28135) );
  ANDN U7470 ( .B(x[2722]), .A(y[2722]), .Z(n12457) );
  ANDN U7471 ( .B(x[2723]), .A(y[2723]), .Z(n20199) );
  NOR U7472 ( .A(n12457), .B(n20199), .Z(n28134) );
  NANDN U7473 ( .A(y[2720]), .B(x[2720]), .Z(n12458) );
  IV U7474 ( .A(n12458), .Z(n28130) );
  ANDN U7475 ( .B(x[2721]), .A(y[2721]), .Z(n28133) );
  NOR U7476 ( .A(n28130), .B(n28133), .Z(n9529) );
  ANDN U7477 ( .B(y[2718]), .A(x[2718]), .Z(n28126) );
  NANDN U7478 ( .A(x[2717]), .B(y[2717]), .Z(n4051) );
  NANDN U7479 ( .A(y[2716]), .B(x[2716]), .Z(n20176) );
  NANDN U7480 ( .A(y[2717]), .B(x[2717]), .Z(n20180) );
  NAND U7481 ( .A(n20176), .B(n20180), .Z(n4049) );
  AND U7482 ( .A(n4051), .B(n4049), .Z(n28125) );
  NANDN U7483 ( .A(x[2716]), .B(y[2716]), .Z(n4050) );
  AND U7484 ( .A(n4051), .B(n4050), .Z(n12460) );
  NANDN U7485 ( .A(x[2715]), .B(y[2715]), .Z(n12462) );
  NAND U7486 ( .A(n12460), .B(n12462), .Z(n9523) );
  NANDN U7487 ( .A(y[2714]), .B(x[2714]), .Z(n28121) );
  NANDN U7488 ( .A(y[2715]), .B(x[2715]), .Z(n28123) );
  AND U7489 ( .A(n28121), .B(n28123), .Z(n9521) );
  ANDN U7490 ( .B(y[2713]), .A(x[2713]), .Z(n20171) );
  NANDN U7491 ( .A(y[2713]), .B(x[2713]), .Z(n4053) );
  NANDN U7492 ( .A(y[2712]), .B(x[2712]), .Z(n4052) );
  NAND U7493 ( .A(n4053), .B(n4052), .Z(n20172) );
  NANDN U7494 ( .A(x[2711]), .B(y[2711]), .Z(n4055) );
  NANDN U7495 ( .A(x[2712]), .B(y[2712]), .Z(n4054) );
  NAND U7496 ( .A(n4055), .B(n4054), .Z(n12467) );
  NANDN U7497 ( .A(y[2711]), .B(x[2711]), .Z(n12463) );
  NANDN U7498 ( .A(y[2710]), .B(x[2710]), .Z(n4056) );
  AND U7499 ( .A(n12463), .B(n4056), .Z(n12469) );
  ANDN U7500 ( .B(y[2709]), .A(x[2709]), .Z(n20167) );
  NANDN U7501 ( .A(y[2708]), .B(x[2708]), .Z(n9511) );
  XOR U7502 ( .A(x[2708]), .B(y[2708]), .Z(n12470) );
  ANDN U7503 ( .B(y[2706]), .A(x[2706]), .Z(n20164) );
  NANDN U7504 ( .A(x[2705]), .B(y[2705]), .Z(n20159) );
  NANDN U7505 ( .A(n20164), .B(n20159), .Z(n24189) );
  NANDN U7506 ( .A(y[2704]), .B(x[2704]), .Z(n9503) );
  XOR U7507 ( .A(x[2704]), .B(y[2704]), .Z(n12473) );
  NANDN U7508 ( .A(y[2701]), .B(x[2701]), .Z(n12477) );
  NANDN U7509 ( .A(y[2700]), .B(x[2700]), .Z(n4057) );
  AND U7510 ( .A(n12477), .B(n4057), .Z(n9496) );
  ANDN U7511 ( .B(y[2699]), .A(x[2699]), .Z(n12480) );
  NANDN U7512 ( .A(y[2699]), .B(x[2699]), .Z(n12479) );
  NANDN U7513 ( .A(x[2697]), .B(y[2697]), .Z(n20143) );
  NANDN U7514 ( .A(x[2698]), .B(y[2698]), .Z(n12481) );
  NAND U7515 ( .A(n20143), .B(n12481), .Z(n24196) );
  NANDN U7516 ( .A(y[2696]), .B(x[2696]), .Z(n12484) );
  ANDN U7517 ( .B(x[2697]), .A(y[2697]), .Z(n20147) );
  ANDN U7518 ( .B(n12484), .A(n20147), .Z(n28108) );
  ANDN U7519 ( .B(y[2694]), .A(x[2694]), .Z(n12485) );
  NANDN U7520 ( .A(x[2693]), .B(y[2693]), .Z(n12488) );
  ANDN U7521 ( .B(x[2692]), .A(y[2692]), .Z(n28101) );
  NANDN U7522 ( .A(y[2693]), .B(x[2693]), .Z(n28103) );
  NANDN U7523 ( .A(x[2692]), .B(y[2692]), .Z(n12489) );
  ANDN U7524 ( .B(x[2691]), .A(y[2691]), .Z(n12490) );
  NANDN U7525 ( .A(y[2690]), .B(x[2690]), .Z(n20130) );
  NANDN U7526 ( .A(n12490), .B(n20130), .Z(n28099) );
  ANDN U7527 ( .B(y[2690]), .A(x[2690]), .Z(n28098) );
  NANDN U7528 ( .A(x[2689]), .B(y[2689]), .Z(n4060) );
  NANDN U7529 ( .A(y[2689]), .B(x[2689]), .Z(n12491) );
  NANDN U7530 ( .A(y[2688]), .B(x[2688]), .Z(n4058) );
  AND U7531 ( .A(n12491), .B(n4058), .Z(n12492) );
  ANDN U7532 ( .B(n4060), .A(n12492), .Z(n28097) );
  NANDN U7533 ( .A(x[2688]), .B(y[2688]), .Z(n4059) );
  AND U7534 ( .A(n4060), .B(n4059), .Z(n28096) );
  NANDN U7535 ( .A(x[2687]), .B(y[2687]), .Z(n12493) );
  ANDN U7536 ( .B(x[2686]), .A(y[2686]), .Z(n9475) );
  NANDN U7537 ( .A(y[2687]), .B(x[2687]), .Z(n28095) );
  NANDN U7538 ( .A(x[2686]), .B(y[2686]), .Z(n12494) );
  NANDN U7539 ( .A(y[2685]), .B(x[2685]), .Z(n12496) );
  NANDN U7540 ( .A(y[2684]), .B(x[2684]), .Z(n12499) );
  AND U7541 ( .A(n12496), .B(n12499), .Z(n9470) );
  ANDN U7542 ( .B(y[2684]), .A(x[2684]), .Z(n12497) );
  NANDN U7543 ( .A(x[2683]), .B(y[2683]), .Z(n20118) );
  NANDN U7544 ( .A(y[2683]), .B(x[2683]), .Z(n12500) );
  NANDN U7545 ( .A(y[2682]), .B(x[2682]), .Z(n4061) );
  AND U7546 ( .A(n12500), .B(n4061), .Z(n9466) );
  XNOR U7547 ( .A(x[2682]), .B(y[2682]), .Z(n12502) );
  NANDN U7548 ( .A(y[2680]), .B(x[2680]), .Z(n28088) );
  ANDN U7549 ( .B(y[2679]), .A(x[2679]), .Z(n20107) );
  ANDN U7550 ( .B(y[2680]), .A(x[2680]), .Z(n20115) );
  NOR U7551 ( .A(n20107), .B(n20115), .Z(n28087) );
  NANDN U7552 ( .A(y[2678]), .B(x[2678]), .Z(n20104) );
  NANDN U7553 ( .A(y[2679]), .B(x[2679]), .Z(n20111) );
  NAND U7554 ( .A(n20104), .B(n20111), .Z(n28086) );
  ANDN U7555 ( .B(y[2677]), .A(x[2677]), .Z(n20100) );
  ANDN U7556 ( .B(y[2678]), .A(x[2678]), .Z(n20110) );
  NOR U7557 ( .A(n20100), .B(n20110), .Z(n28085) );
  NANDN U7558 ( .A(y[2676]), .B(x[2676]), .Z(n12503) );
  NANDN U7559 ( .A(y[2677]), .B(x[2677]), .Z(n20105) );
  NAND U7560 ( .A(n12503), .B(n20105), .Z(n28084) );
  ANDN U7561 ( .B(y[2675]), .A(x[2675]), .Z(n20094) );
  ANDN U7562 ( .B(y[2676]), .A(x[2676]), .Z(n20102) );
  NOR U7563 ( .A(n20094), .B(n20102), .Z(n28083) );
  NANDN U7564 ( .A(y[2674]), .B(x[2674]), .Z(n20090) );
  NANDN U7565 ( .A(y[2675]), .B(x[2675]), .Z(n12504) );
  NAND U7566 ( .A(n20090), .B(n12504), .Z(n24199) );
  ANDN U7567 ( .B(y[2674]), .A(x[2674]), .Z(n20095) );
  NANDN U7568 ( .A(x[2673]), .B(y[2673]), .Z(n12505) );
  NANDN U7569 ( .A(n20095), .B(n12505), .Z(n28082) );
  NANDN U7570 ( .A(y[2672]), .B(x[2672]), .Z(n20086) );
  NANDN U7571 ( .A(y[2673]), .B(x[2673]), .Z(n20089) );
  AND U7572 ( .A(n20086), .B(n20089), .Z(n28081) );
  NANDN U7573 ( .A(x[2671]), .B(y[2671]), .Z(n20083) );
  NANDN U7574 ( .A(x[2672]), .B(y[2672]), .Z(n12506) );
  NAND U7575 ( .A(n20083), .B(n12506), .Z(n28080) );
  NANDN U7576 ( .A(y[2671]), .B(x[2671]), .Z(n12508) );
  NANDN U7577 ( .A(y[2670]), .B(x[2670]), .Z(n4062) );
  AND U7578 ( .A(n12508), .B(n4062), .Z(n28078) );
  ANDN U7579 ( .B(x[2669]), .A(y[2669]), .Z(n20081) );
  NANDN U7580 ( .A(y[2668]), .B(x[2668]), .Z(n12510) );
  NANDN U7581 ( .A(n20081), .B(n12510), .Z(n28076) );
  ANDN U7582 ( .B(y[2667]), .A(x[2667]), .Z(n20071) );
  ANDN U7583 ( .B(y[2668]), .A(x[2668]), .Z(n20078) );
  NOR U7584 ( .A(n20071), .B(n20078), .Z(n28075) );
  NANDN U7585 ( .A(x[2665]), .B(y[2665]), .Z(n12512) );
  NANDN U7586 ( .A(x[2666]), .B(y[2666]), .Z(n20072) );
  AND U7587 ( .A(n12512), .B(n20072), .Z(n9445) );
  ANDN U7588 ( .B(x[2664]), .A(y[2664]), .Z(n9443) );
  NANDN U7589 ( .A(y[2665]), .B(x[2665]), .Z(n28071) );
  NANDN U7590 ( .A(y[2662]), .B(x[2662]), .Z(n28067) );
  NANDN U7591 ( .A(y[2661]), .B(x[2661]), .Z(n28065) );
  NANDN U7592 ( .A(y[2660]), .B(x[2660]), .Z(n4063) );
  AND U7593 ( .A(n28065), .B(n4063), .Z(n9435) );
  XNOR U7594 ( .A(x[2660]), .B(y[2660]), .Z(n12519) );
  NANDN U7595 ( .A(x[2657]), .B(y[2657]), .Z(n12520) );
  ANDN U7596 ( .B(y[2658]), .A(x[2658]), .Z(n20056) );
  ANDN U7597 ( .B(n12520), .A(n20056), .Z(n28061) );
  ANDN U7598 ( .B(x[2657]), .A(y[2657]), .Z(n20052) );
  NANDN U7599 ( .A(x[2653]), .B(y[2653]), .Z(n12528) );
  ANDN U7600 ( .B(x[2652]), .A(y[2652]), .Z(n28053) );
  NANDN U7601 ( .A(x[2645]), .B(y[2645]), .Z(n4065) );
  NANDN U7602 ( .A(x[2646]), .B(y[2646]), .Z(n4064) );
  NAND U7603 ( .A(n4065), .B(n4064), .Z(n12535) );
  NANDN U7604 ( .A(y[2644]), .B(x[2644]), .Z(n4066) );
  NANDN U7605 ( .A(y[2645]), .B(x[2645]), .Z(n12533) );
  AND U7606 ( .A(n4066), .B(n12533), .Z(n12537) );
  ANDN U7607 ( .B(y[2644]), .A(x[2644]), .Z(n12534) );
  NANDN U7608 ( .A(x[2643]), .B(y[2643]), .Z(n12539) );
  NANDN U7609 ( .A(y[2643]), .B(x[2643]), .Z(n12536) );
  NANDN U7610 ( .A(y[2642]), .B(x[2642]), .Z(n4067) );
  AND U7611 ( .A(n12536), .B(n4067), .Z(n9399) );
  ANDN U7612 ( .B(y[2642]), .A(x[2642]), .Z(n12538) );
  ANDN U7613 ( .B(x[2640]), .A(y[2640]), .Z(n28042) );
  ANDN U7614 ( .B(x[2641]), .A(y[2641]), .Z(n20034) );
  NOR U7615 ( .A(n28042), .B(n20034), .Z(n9395) );
  ANDN U7616 ( .B(x[2638]), .A(y[2638]), .Z(n20023) );
  ANDN U7617 ( .B(x[2639]), .A(y[2639]), .Z(n20029) );
  NOR U7618 ( .A(n20023), .B(n20029), .Z(n28037) );
  NANDN U7619 ( .A(x[2637]), .B(y[2637]), .Z(n20021) );
  NANDN U7620 ( .A(x[2638]), .B(y[2638]), .Z(n28038) );
  AND U7621 ( .A(n20021), .B(n28038), .Z(n24205) );
  NANDN U7622 ( .A(x[2636]), .B(y[2636]), .Z(n20019) );
  ANDN U7623 ( .B(y[2635]), .A(x[2635]), .Z(n20015) );
  ANDN U7624 ( .B(n20019), .A(n20015), .Z(n24204) );
  NANDN U7625 ( .A(y[2634]), .B(x[2634]), .Z(n12542) );
  ANDN U7626 ( .B(y[2633]), .A(x[2633]), .Z(n12544) );
  NANDN U7627 ( .A(y[2630]), .B(x[2630]), .Z(n20005) );
  NANDN U7628 ( .A(y[2631]), .B(x[2631]), .Z(n4068) );
  AND U7629 ( .A(n20005), .B(n4068), .Z(n28031) );
  NANDN U7630 ( .A(x[2629]), .B(y[2629]), .Z(n4070) );
  NANDN U7631 ( .A(x[2630]), .B(y[2630]), .Z(n4069) );
  NAND U7632 ( .A(n4070), .B(n4069), .Z(n28030) );
  NANDN U7633 ( .A(y[2629]), .B(x[2629]), .Z(n4072) );
  NANDN U7634 ( .A(y[2628]), .B(x[2628]), .Z(n4071) );
  AND U7635 ( .A(n4072), .B(n4071), .Z(n28029) );
  NANDN U7636 ( .A(x[2627]), .B(y[2627]), .Z(n4074) );
  NANDN U7637 ( .A(x[2628]), .B(y[2628]), .Z(n4073) );
  NAND U7638 ( .A(n4074), .B(n4073), .Z(n28026) );
  NANDN U7639 ( .A(y[2626]), .B(x[2626]), .Z(n4075) );
  ANDN U7640 ( .B(x[2627]), .A(y[2627]), .Z(n28025) );
  ANDN U7641 ( .B(n4075), .A(n28025), .Z(n28023) );
  NANDN U7642 ( .A(x[2625]), .B(y[2625]), .Z(n28021) );
  NANDN U7643 ( .A(x[2626]), .B(y[2626]), .Z(n28024) );
  NAND U7644 ( .A(n28021), .B(n28024), .Z(n19999) );
  NANDN U7645 ( .A(y[2625]), .B(x[2625]), .Z(n19997) );
  NANDN U7646 ( .A(y[2624]), .B(x[2624]), .Z(n4076) );
  AND U7647 ( .A(n19997), .B(n4076), .Z(n28020) );
  NANDN U7648 ( .A(y[2622]), .B(x[2622]), .Z(n19985) );
  NANDN U7649 ( .A(y[2623]), .B(x[2623]), .Z(n19991) );
  AND U7650 ( .A(n19985), .B(n19991), .Z(n28018) );
  ANDN U7651 ( .B(y[2622]), .A(x[2622]), .Z(n28017) );
  NANDN U7652 ( .A(x[2621]), .B(y[2621]), .Z(n12546) );
  ANDN U7653 ( .B(x[2620]), .A(y[2620]), .Z(n28014) );
  NANDN U7654 ( .A(y[2621]), .B(x[2621]), .Z(n28016) );
  NANDN U7655 ( .A(x[2620]), .B(y[2620]), .Z(n12547) );
  ANDN U7656 ( .B(x[2618]), .A(y[2618]), .Z(n12549) );
  ANDN U7657 ( .B(x[2619]), .A(y[2619]), .Z(n19981) );
  OR U7658 ( .A(n12549), .B(n19981), .Z(n28012) );
  NANDN U7659 ( .A(x[2618]), .B(y[2618]), .Z(n19977) );
  ANDN U7660 ( .B(y[2617]), .A(x[2617]), .Z(n19973) );
  ANDN U7661 ( .B(n19977), .A(n19973), .Z(n28011) );
  ANDN U7662 ( .B(x[2616]), .A(y[2616]), .Z(n9380) );
  XOR U7663 ( .A(x[2616]), .B(y[2616]), .Z(n12550) );
  NANDN U7664 ( .A(y[2614]), .B(x[2614]), .Z(n28005) );
  NANDN U7665 ( .A(y[2615]), .B(x[2615]), .Z(n12551) );
  ANDN U7666 ( .B(y[2613]), .A(x[2613]), .Z(n19965) );
  NANDN U7667 ( .A(x[2614]), .B(y[2614]), .Z(n12553) );
  NANDN U7668 ( .A(n19965), .B(n12553), .Z(n28006) );
  NANDN U7669 ( .A(y[2612]), .B(x[2612]), .Z(n12555) );
  NANDN U7670 ( .A(x[2611]), .B(y[2611]), .Z(n12557) );
  NANDN U7671 ( .A(x[2612]), .B(y[2612]), .Z(n19966) );
  AND U7672 ( .A(n12557), .B(n19966), .Z(n28002) );
  NANDN U7673 ( .A(y[2610]), .B(x[2610]), .Z(n28001) );
  NANDN U7674 ( .A(x[2609]), .B(y[2609]), .Z(n19956) );
  NANDN U7675 ( .A(x[2610]), .B(y[2610]), .Z(n12558) );
  NAND U7676 ( .A(n19956), .B(n12558), .Z(n28000) );
  NANDN U7677 ( .A(y[2609]), .B(x[2609]), .Z(n12559) );
  ANDN U7678 ( .B(x[2608]), .A(y[2608]), .Z(n19952) );
  ANDN U7679 ( .B(n12559), .A(n19952), .Z(n27999) );
  ANDN U7680 ( .B(y[2608]), .A(x[2608]), .Z(n19958) );
  NANDN U7681 ( .A(x[2607]), .B(y[2607]), .Z(n19948) );
  NANDN U7682 ( .A(n19958), .B(n19948), .Z(n27998) );
  ANDN U7683 ( .B(x[2606]), .A(y[2606]), .Z(n12560) );
  ANDN U7684 ( .B(x[2607]), .A(y[2607]), .Z(n19954) );
  NOR U7685 ( .A(n12560), .B(n19954), .Z(n27997) );
  ANDN U7686 ( .B(x[2604]), .A(y[2604]), .Z(n19941) );
  NANDN U7687 ( .A(y[2603]), .B(x[2603]), .Z(n19939) );
  NANDN U7688 ( .A(y[2602]), .B(x[2602]), .Z(n4077) );
  AND U7689 ( .A(n19939), .B(n4077), .Z(n4080) );
  NANDN U7690 ( .A(x[2602]), .B(y[2602]), .Z(n19937) );
  ANDN U7691 ( .B(y[2601]), .A(x[2601]), .Z(n19929) );
  ANDN U7692 ( .B(n19937), .A(n19929), .Z(n4081) );
  NANDN U7693 ( .A(y[2600]), .B(x[2600]), .Z(n19925) );
  NANDN U7694 ( .A(y[2601]), .B(x[2601]), .Z(n19933) );
  NAND U7695 ( .A(n19925), .B(n19933), .Z(n4078) );
  NAND U7696 ( .A(n4081), .B(n4078), .Z(n4079) );
  NAND U7697 ( .A(n4080), .B(n4079), .Z(n27994) );
  NANDN U7698 ( .A(x[2599]), .B(y[2599]), .Z(n12562) );
  ANDN U7699 ( .B(y[2600]), .A(x[2600]), .Z(n19931) );
  ANDN U7700 ( .B(n4081), .A(n19931), .Z(n24216) );
  NANDN U7701 ( .A(y[2599]), .B(x[2599]), .Z(n24213) );
  NANDN U7702 ( .A(y[2598]), .B(x[2598]), .Z(n12563) );
  NAND U7703 ( .A(n24213), .B(n12563), .Z(n27992) );
  ANDN U7704 ( .B(y[2596]), .A(x[2596]), .Z(n19919) );
  NANDN U7705 ( .A(x[2595]), .B(y[2595]), .Z(n12566) );
  NANDN U7706 ( .A(n19919), .B(n12566), .Z(n27989) );
  NANDN U7707 ( .A(y[2593]), .B(x[2593]), .Z(n12568) );
  NANDN U7708 ( .A(y[2592]), .B(x[2592]), .Z(n24217) );
  AND U7709 ( .A(n12568), .B(n24217), .Z(n9345) );
  NANDN U7710 ( .A(x[2591]), .B(y[2591]), .Z(n12570) );
  ANDN U7711 ( .B(y[2592]), .A(x[2592]), .Z(n19909) );
  ANDN U7712 ( .B(n12570), .A(n19909), .Z(n27984) );
  NANDN U7713 ( .A(y[2590]), .B(x[2590]), .Z(n12571) );
  NANDN U7714 ( .A(y[2591]), .B(x[2591]), .Z(n19905) );
  NAND U7715 ( .A(n12571), .B(n19905), .Z(n27983) );
  NANDN U7716 ( .A(x[2589]), .B(y[2589]), .Z(n12573) );
  NANDN U7717 ( .A(x[2590]), .B(y[2590]), .Z(n12569) );
  AND U7718 ( .A(n12573), .B(n12569), .Z(n27982) );
  NANDN U7719 ( .A(y[2588]), .B(x[2588]), .Z(n19895) );
  NANDN U7720 ( .A(y[2589]), .B(x[2589]), .Z(n12572) );
  NAND U7721 ( .A(n19895), .B(n12572), .Z(n27981) );
  NANDN U7722 ( .A(y[2586]), .B(x[2586]), .Z(n19889) );
  NANDN U7723 ( .A(y[2587]), .B(x[2587]), .Z(n19896) );
  NAND U7724 ( .A(n19889), .B(n19896), .Z(n24219) );
  NANDN U7725 ( .A(x[2585]), .B(y[2585]), .Z(n19885) );
  NANDN U7726 ( .A(x[2586]), .B(y[2586]), .Z(n12576) );
  NAND U7727 ( .A(n19885), .B(n12576), .Z(n27979) );
  NANDN U7728 ( .A(y[2584]), .B(x[2584]), .Z(n19883) );
  NANDN U7729 ( .A(y[2585]), .B(x[2585]), .Z(n19890) );
  AND U7730 ( .A(n19883), .B(n19890), .Z(n27978) );
  ANDN U7731 ( .B(y[2583]), .A(x[2583]), .Z(n19881) );
  NANDN U7732 ( .A(x[2584]), .B(y[2584]), .Z(n19886) );
  NANDN U7733 ( .A(n19881), .B(n19886), .Z(n27977) );
  NANDN U7734 ( .A(y[2582]), .B(x[2582]), .Z(n19879) );
  NANDN U7735 ( .A(y[2583]), .B(x[2583]), .Z(n27976) );
  AND U7736 ( .A(n19879), .B(n27976), .Z(n9334) );
  ANDN U7737 ( .B(y[2582]), .A(x[2582]), .Z(n19877) );
  NANDN U7738 ( .A(y[2579]), .B(x[2579]), .Z(n12578) );
  NANDN U7739 ( .A(y[2578]), .B(x[2578]), .Z(n4082) );
  AND U7740 ( .A(n12578), .B(n4082), .Z(n12581) );
  NANDN U7741 ( .A(x[2578]), .B(y[2578]), .Z(n12577) );
  NANDN U7742 ( .A(x[2577]), .B(y[2577]), .Z(n12582) );
  ANDN U7743 ( .B(x[2577]), .A(y[2577]), .Z(n12580) );
  XNOR U7744 ( .A(x[2576]), .B(y[2576]), .Z(n12585) );
  NANDN U7745 ( .A(x[2575]), .B(y[2575]), .Z(n12586) );
  ANDN U7746 ( .B(x[2574]), .A(y[2574]), .Z(n12588) );
  NANDN U7747 ( .A(x[2574]), .B(y[2574]), .Z(n12587) );
  NANDN U7748 ( .A(y[2572]), .B(x[2572]), .Z(n19862) );
  NANDN U7749 ( .A(y[2573]), .B(x[2573]), .Z(n27967) );
  AND U7750 ( .A(n19862), .B(n27967), .Z(n9312) );
  ANDN U7751 ( .B(y[2571]), .A(x[2571]), .Z(n12589) );
  ANDN U7752 ( .B(x[2570]), .A(y[2570]), .Z(n24222) );
  NANDN U7753 ( .A(x[2569]), .B(y[2569]), .Z(n24223) );
  ANDN U7754 ( .B(y[2567]), .A(x[2567]), .Z(n12592) );
  NANDN U7755 ( .A(y[2566]), .B(x[2566]), .Z(n12594) );
  ANDN U7756 ( .B(y[2565]), .A(x[2565]), .Z(n12596) );
  NANDN U7757 ( .A(y[2564]), .B(x[2564]), .Z(n12599) );
  ANDN U7758 ( .B(x[2562]), .A(y[2562]), .Z(n27957) );
  NANDN U7759 ( .A(x[2561]), .B(y[2561]), .Z(n12601) );
  NANDN U7760 ( .A(y[2560]), .B(x[2560]), .Z(n12603) );
  NANDN U7761 ( .A(y[2561]), .B(x[2561]), .Z(n27954) );
  NAND U7762 ( .A(n12603), .B(n27954), .Z(n9288) );
  NANDN U7763 ( .A(x[2559]), .B(y[2559]), .Z(n27950) );
  ANDN U7764 ( .B(x[2558]), .A(y[2558]), .Z(n19837) );
  ANDN U7765 ( .B(x[2559]), .A(y[2559]), .Z(n19843) );
  OR U7766 ( .A(n19837), .B(n19843), .Z(n27949) );
  NANDN U7767 ( .A(x[2557]), .B(y[2557]), .Z(n19833) );
  NANDN U7768 ( .A(x[2558]), .B(y[2558]), .Z(n12604) );
  AND U7769 ( .A(n19833), .B(n12604), .Z(n27948) );
  ANDN U7770 ( .B(x[2557]), .A(y[2557]), .Z(n19838) );
  NANDN U7771 ( .A(y[2556]), .B(x[2556]), .Z(n12605) );
  NANDN U7772 ( .A(n19838), .B(n12605), .Z(n27947) );
  NANDN U7773 ( .A(x[2555]), .B(y[2555]), .Z(n12606) );
  NANDN U7774 ( .A(x[2556]), .B(y[2556]), .Z(n27946) );
  AND U7775 ( .A(n12606), .B(n27946), .Z(n9281) );
  ANDN U7776 ( .B(x[2554]), .A(y[2554]), .Z(n9279) );
  NANDN U7777 ( .A(y[2551]), .B(x[2551]), .Z(n12611) );
  NANDN U7778 ( .A(y[2550]), .B(x[2550]), .Z(n19820) );
  AND U7779 ( .A(n12611), .B(n19820), .Z(n9271) );
  ANDN U7780 ( .B(y[2550]), .A(x[2550]), .Z(n12612) );
  NANDN U7781 ( .A(y[2549]), .B(x[2549]), .Z(n19821) );
  NANDN U7782 ( .A(y[2548]), .B(x[2548]), .Z(n12615) );
  AND U7783 ( .A(n19821), .B(n12615), .Z(n9267) );
  ANDN U7784 ( .B(y[2546]), .A(x[2546]), .Z(n19814) );
  NANDN U7785 ( .A(x[2545]), .B(y[2545]), .Z(n12616) );
  NANDN U7786 ( .A(n19814), .B(n12616), .Z(n27932) );
  NANDN U7787 ( .A(y[2544]), .B(x[2544]), .Z(n12618) );
  NANDN U7788 ( .A(y[2545]), .B(x[2545]), .Z(n19807) );
  NAND U7789 ( .A(n12618), .B(n19807), .Z(n27931) );
  NANDN U7790 ( .A(x[2543]), .B(y[2543]), .Z(n12620) );
  NANDN U7791 ( .A(x[2544]), .B(y[2544]), .Z(n12617) );
  AND U7792 ( .A(n12620), .B(n12617), .Z(n27930) );
  NANDN U7793 ( .A(y[2542]), .B(x[2542]), .Z(n12621) );
  NANDN U7794 ( .A(y[2543]), .B(x[2543]), .Z(n12619) );
  NAND U7795 ( .A(n12621), .B(n12619), .Z(n27929) );
  NANDN U7796 ( .A(x[2542]), .B(y[2542]), .Z(n27928) );
  NANDN U7797 ( .A(x[2539]), .B(y[2539]), .Z(n12623) );
  NANDN U7798 ( .A(x[2541]), .B(y[2541]), .Z(n9256) );
  NANDN U7799 ( .A(x[2540]), .B(y[2540]), .Z(n4083) );
  AND U7800 ( .A(n9256), .B(n4083), .Z(n27927) );
  AND U7801 ( .A(n12623), .B(n27927), .Z(n9255) );
  NANDN U7802 ( .A(y[2539]), .B(x[2539]), .Z(n12626) );
  NANDN U7803 ( .A(y[2538]), .B(x[2538]), .Z(n4084) );
  NAND U7804 ( .A(n12626), .B(n4084), .Z(n27926) );
  NANDN U7805 ( .A(x[2537]), .B(y[2537]), .Z(n27925) );
  NANDN U7806 ( .A(x[2535]), .B(y[2535]), .Z(n19783) );
  NANDN U7807 ( .A(x[2536]), .B(y[2536]), .Z(n19789) );
  AND U7808 ( .A(n19783), .B(n19789), .Z(n27923) );
  ANDN U7809 ( .B(x[2534]), .A(y[2534]), .Z(n19779) );
  ANDN U7810 ( .B(x[2535]), .A(y[2535]), .Z(n19788) );
  OR U7811 ( .A(n19779), .B(n19788), .Z(n27922) );
  NANDN U7812 ( .A(x[2534]), .B(y[2534]), .Z(n24229) );
  NANDN U7813 ( .A(y[2530]), .B(x[2530]), .Z(n12631) );
  NANDN U7814 ( .A(y[2531]), .B(x[2531]), .Z(n12628) );
  NAND U7815 ( .A(n12631), .B(n12628), .Z(n27918) );
  NANDN U7816 ( .A(x[2529]), .B(y[2529]), .Z(n12633) );
  NANDN U7817 ( .A(x[2530]), .B(y[2530]), .Z(n12630) );
  AND U7818 ( .A(n12633), .B(n12630), .Z(n27917) );
  ANDN U7819 ( .B(x[2528]), .A(y[2528]), .Z(n19767) );
  NANDN U7820 ( .A(y[2529]), .B(x[2529]), .Z(n12632) );
  NANDN U7821 ( .A(n19767), .B(n12632), .Z(n27916) );
  NANDN U7822 ( .A(x[2528]), .B(y[2528]), .Z(n27915) );
  ANDN U7823 ( .B(y[2527]), .A(x[2527]), .Z(n27914) );
  ANDN U7824 ( .B(n27915), .A(n27914), .Z(n9239) );
  ANDN U7825 ( .B(x[2526]), .A(y[2526]), .Z(n12634) );
  NANDN U7826 ( .A(y[2525]), .B(x[2525]), .Z(n12635) );
  NANDN U7827 ( .A(y[2524]), .B(x[2524]), .Z(n4085) );
  AND U7828 ( .A(n12635), .B(n4085), .Z(n9234) );
  ANDN U7829 ( .B(y[2523]), .A(x[2523]), .Z(n24234) );
  NANDN U7830 ( .A(y[2523]), .B(x[2523]), .Z(n12638) );
  NANDN U7831 ( .A(y[2522]), .B(x[2522]), .Z(n24235) );
  AND U7832 ( .A(n12638), .B(n24235), .Z(n9230) );
  NANDN U7833 ( .A(y[2516]), .B(x[2516]), .Z(n4086) );
  NANDN U7834 ( .A(y[2517]), .B(x[2517]), .Z(n12641) );
  AND U7835 ( .A(n4086), .B(n12641), .Z(n27906) );
  ANDN U7836 ( .B(x[2515]), .A(y[2515]), .Z(n19744) );
  NANDN U7837 ( .A(y[2514]), .B(x[2514]), .Z(n12645) );
  NANDN U7838 ( .A(n19744), .B(n12645), .Z(n27904) );
  ANDN U7839 ( .B(y[2513]), .A(x[2513]), .Z(n19735) );
  ANDN U7840 ( .B(y[2514]), .A(x[2514]), .Z(n19741) );
  NOR U7841 ( .A(n19735), .B(n19741), .Z(n27903) );
  NANDN U7842 ( .A(y[2512]), .B(x[2512]), .Z(n12646) );
  NANDN U7843 ( .A(y[2513]), .B(x[2513]), .Z(n12644) );
  NAND U7844 ( .A(n12646), .B(n12644), .Z(n27902) );
  NANDN U7845 ( .A(x[2511]), .B(y[2511]), .Z(n19729) );
  ANDN U7846 ( .B(y[2512]), .A(x[2512]), .Z(n27901) );
  ANDN U7847 ( .B(n19729), .A(n27901), .Z(n9211) );
  NANDN U7848 ( .A(y[2511]), .B(x[2511]), .Z(n27900) );
  NANDN U7849 ( .A(x[2510]), .B(y[2510]), .Z(n19730) );
  ANDN U7850 ( .B(x[2508]), .A(y[2508]), .Z(n19721) );
  NANDN U7851 ( .A(y[2509]), .B(x[2509]), .Z(n12647) );
  NANDN U7852 ( .A(n19721), .B(n12647), .Z(n27895) );
  NANDN U7853 ( .A(x[2507]), .B(y[2507]), .Z(n19717) );
  NANDN U7854 ( .A(x[2508]), .B(y[2508]), .Z(n19725) );
  AND U7855 ( .A(n19717), .B(n19725), .Z(n27894) );
  ANDN U7856 ( .B(x[2506]), .A(y[2506]), .Z(n12648) );
  NANDN U7857 ( .A(x[2505]), .B(y[2505]), .Z(n27890) );
  NANDN U7858 ( .A(x[2506]), .B(y[2506]), .Z(n27892) );
  NAND U7859 ( .A(n27890), .B(n27892), .Z(n9201) );
  NANDN U7860 ( .A(y[2505]), .B(x[2505]), .Z(n12649) );
  ANDN U7861 ( .B(x[2504]), .A(y[2504]), .Z(n27889) );
  ANDN U7862 ( .B(n12649), .A(n27889), .Z(n9199) );
  NANDN U7863 ( .A(y[2502]), .B(x[2502]), .Z(n4088) );
  ANDN U7864 ( .B(x[2503]), .A(y[2503]), .Z(n4087) );
  ANDN U7865 ( .B(n4088), .A(n4087), .Z(n27887) );
  NANDN U7866 ( .A(y[2501]), .B(x[2501]), .Z(n19707) );
  NANDN U7867 ( .A(y[2500]), .B(x[2500]), .Z(n4089) );
  AND U7868 ( .A(n19707), .B(n4089), .Z(n27885) );
  ANDN U7869 ( .B(y[2499]), .A(x[2499]), .Z(n19700) );
  ANDN U7870 ( .B(y[2500]), .A(x[2500]), .Z(n19705) );
  OR U7871 ( .A(n19700), .B(n19705), .Z(n27884) );
  NANDN U7872 ( .A(y[2499]), .B(x[2499]), .Z(n19702) );
  NANDN U7873 ( .A(x[2497]), .B(y[2497]), .Z(n4098) );
  XNOR U7874 ( .A(x[2497]), .B(y[2497]), .Z(n4091) );
  NANDN U7875 ( .A(y[2496]), .B(x[2496]), .Z(n4090) );
  NAND U7876 ( .A(n4091), .B(n4090), .Z(n4092) );
  NAND U7877 ( .A(n4098), .B(n4092), .Z(n4094) );
  NANDN U7878 ( .A(y[2498]), .B(x[2498]), .Z(n4093) );
  AND U7879 ( .A(n4094), .B(n4093), .Z(n19696) );
  NANDN U7880 ( .A(x[2498]), .B(y[2498]), .Z(n19698) );
  NANDN U7881 ( .A(n19696), .B(n19698), .Z(n4095) );
  AND U7882 ( .A(n19702), .B(n4095), .Z(n27883) );
  NANDN U7883 ( .A(x[2496]), .B(y[2496]), .Z(n4097) );
  NANDN U7884 ( .A(x[2495]), .B(y[2495]), .Z(n4096) );
  AND U7885 ( .A(n4097), .B(n4096), .Z(n4099) );
  NAND U7886 ( .A(n4099), .B(n4098), .Z(n19694) );
  ANDN U7887 ( .B(n19698), .A(n19694), .Z(n27881) );
  NANDN U7888 ( .A(y[2495]), .B(x[2495]), .Z(n12650) );
  NANDN U7889 ( .A(y[2494]), .B(x[2494]), .Z(n4100) );
  NAND U7890 ( .A(n12650), .B(n4100), .Z(n12652) );
  NANDN U7891 ( .A(x[2492]), .B(y[2492]), .Z(n27877) );
  NANDN U7892 ( .A(x[2491]), .B(y[2491]), .Z(n27876) );
  NAND U7893 ( .A(n27877), .B(n27876), .Z(n9183) );
  NANDN U7894 ( .A(y[2491]), .B(x[2491]), .Z(n12656) );
  ANDN U7895 ( .B(x[2490]), .A(y[2490]), .Z(n19681) );
  ANDN U7896 ( .B(n12656), .A(n19681), .Z(n27875) );
  ANDN U7897 ( .B(y[2489]), .A(x[2489]), .Z(n12657) );
  NANDN U7898 ( .A(x[2490]), .B(y[2490]), .Z(n27874) );
  NANDN U7899 ( .A(x[2488]), .B(y[2488]), .Z(n12658) );
  ANDN U7900 ( .B(y[2487]), .A(x[2487]), .Z(n12660) );
  ANDN U7901 ( .B(n12658), .A(n12660), .Z(n9176) );
  NANDN U7902 ( .A(x[2485]), .B(y[2485]), .Z(n19669) );
  NANDN U7903 ( .A(x[2486]), .B(y[2486]), .Z(n12661) );
  AND U7904 ( .A(n19669), .B(n12661), .Z(n27868) );
  ANDN U7905 ( .B(x[2485]), .A(y[2485]), .Z(n27867) );
  NANDN U7906 ( .A(x[2484]), .B(y[2484]), .Z(n27866) );
  NANDN U7907 ( .A(y[2482]), .B(x[2482]), .Z(n27862) );
  NANDN U7908 ( .A(x[2482]), .B(y[2482]), .Z(n12665) );
  ANDN U7909 ( .B(x[2481]), .A(y[2481]), .Z(n12666) );
  NANDN U7910 ( .A(x[2480]), .B(y[2480]), .Z(n27859) );
  NANDN U7911 ( .A(y[2479]), .B(x[2479]), .Z(n4102) );
  NANDN U7912 ( .A(y[2480]), .B(x[2480]), .Z(n4101) );
  NAND U7913 ( .A(n4102), .B(n4101), .Z(n27858) );
  NANDN U7914 ( .A(x[2479]), .B(y[2479]), .Z(n4104) );
  NANDN U7915 ( .A(x[2478]), .B(y[2478]), .Z(n4103) );
  AND U7916 ( .A(n4104), .B(n4103), .Z(n27856) );
  NANDN U7917 ( .A(x[2477]), .B(y[2477]), .Z(n4106) );
  NANDN U7918 ( .A(x[2476]), .B(y[2476]), .Z(n4105) );
  AND U7919 ( .A(n4106), .B(n4105), .Z(n27854) );
  NANDN U7920 ( .A(y[2475]), .B(x[2475]), .Z(n4108) );
  ANDN U7921 ( .B(x[2476]), .A(y[2476]), .Z(n4107) );
  ANDN U7922 ( .B(n4108), .A(n4107), .Z(n4112) );
  XNOR U7923 ( .A(x[2475]), .B(y[2475]), .Z(n4110) );
  ANDN U7924 ( .B(x[2474]), .A(y[2474]), .Z(n4109) );
  NAND U7925 ( .A(n4110), .B(n4109), .Z(n4111) );
  NAND U7926 ( .A(n4112), .B(n4111), .Z(n27853) );
  NANDN U7927 ( .A(y[2472]), .B(x[2472]), .Z(n4113) );
  NANDN U7928 ( .A(y[2473]), .B(x[2473]), .Z(n12667) );
  AND U7929 ( .A(n4113), .B(n12667), .Z(n27851) );
  NANDN U7930 ( .A(y[2471]), .B(x[2471]), .Z(n12670) );
  ANDN U7931 ( .B(x[2470]), .A(y[2470]), .Z(n19652) );
  ANDN U7932 ( .B(n12670), .A(n19652), .Z(n27850) );
  ANDN U7933 ( .B(x[2464]), .A(y[2464]), .Z(n19640) );
  ANDN U7934 ( .B(x[2465]), .A(y[2465]), .Z(n19644) );
  NOR U7935 ( .A(n19640), .B(n19644), .Z(n27841) );
  NANDN U7936 ( .A(x[2463]), .B(y[2463]), .Z(n12679) );
  NANDN U7937 ( .A(x[2464]), .B(y[2464]), .Z(n19642) );
  NAND U7938 ( .A(n12679), .B(n19642), .Z(n24238) );
  NANDN U7939 ( .A(x[2461]), .B(y[2461]), .Z(n27836) );
  NANDN U7940 ( .A(x[2462]), .B(y[2462]), .Z(n27839) );
  NAND U7941 ( .A(n27836), .B(n27839), .Z(n9130) );
  NANDN U7942 ( .A(x[2460]), .B(y[2460]), .Z(n19633) );
  ANDN U7943 ( .B(y[2459]), .A(x[2459]), .Z(n19628) );
  ANDN U7944 ( .B(n19633), .A(n19628), .Z(n24240) );
  NANDN U7945 ( .A(y[2459]), .B(x[2459]), .Z(n12682) );
  NANDN U7946 ( .A(y[2458]), .B(x[2458]), .Z(n12684) );
  AND U7947 ( .A(n12682), .B(n12684), .Z(n9125) );
  NANDN U7948 ( .A(x[2457]), .B(y[2457]), .Z(n27832) );
  ANDN U7949 ( .B(x[2456]), .A(y[2456]), .Z(n12686) );
  NANDN U7950 ( .A(x[2456]), .B(y[2456]), .Z(n12685) );
  ANDN U7951 ( .B(y[2455]), .A(x[2455]), .Z(n19619) );
  ANDN U7952 ( .B(n12685), .A(n19619), .Z(n27830) );
  NANDN U7953 ( .A(y[2454]), .B(x[2454]), .Z(n12688) );
  NANDN U7954 ( .A(y[2455]), .B(x[2455]), .Z(n12687) );
  NAND U7955 ( .A(n12688), .B(n12687), .Z(n27829) );
  ANDN U7956 ( .B(y[2453]), .A(x[2453]), .Z(n19613) );
  ANDN U7957 ( .B(y[2454]), .A(x[2454]), .Z(n19620) );
  NOR U7958 ( .A(n19613), .B(n19620), .Z(n27828) );
  NANDN U7959 ( .A(x[2451]), .B(y[2451]), .Z(n12691) );
  ANDN U7960 ( .B(y[2452]), .A(x[2452]), .Z(n19614) );
  ANDN U7961 ( .B(n12691), .A(n19614), .Z(n27826) );
  NANDN U7962 ( .A(y[2450]), .B(x[2450]), .Z(n19606) );
  NANDN U7963 ( .A(y[2451]), .B(x[2451]), .Z(n27825) );
  NAND U7964 ( .A(n19606), .B(n27825), .Z(n9114) );
  NANDN U7965 ( .A(x[2449]), .B(y[2449]), .Z(n19603) );
  NANDN U7966 ( .A(x[2450]), .B(y[2450]), .Z(n12690) );
  NANDN U7967 ( .A(y[2449]), .B(x[2449]), .Z(n4115) );
  NANDN U7968 ( .A(y[2448]), .B(x[2448]), .Z(n4114) );
  NAND U7969 ( .A(n4115), .B(n4114), .Z(n19601) );
  NANDN U7970 ( .A(x[2448]), .B(y[2448]), .Z(n4117) );
  NANDN U7971 ( .A(x[2447]), .B(y[2447]), .Z(n4116) );
  AND U7972 ( .A(n4117), .B(n4116), .Z(n19599) );
  NANDN U7973 ( .A(y[2447]), .B(x[2447]), .Z(n19598) );
  NANDN U7974 ( .A(y[2446]), .B(x[2446]), .Z(n4118) );
  AND U7975 ( .A(n19598), .B(n4118), .Z(n9106) );
  NANDN U7976 ( .A(y[2445]), .B(x[2445]), .Z(n4119) );
  AND U7977 ( .A(n9106), .B(n4119), .Z(n27819) );
  NANDN U7978 ( .A(x[2444]), .B(y[2444]), .Z(n19594) );
  ANDN U7979 ( .B(y[2443]), .A(x[2443]), .Z(n19587) );
  NANDN U7980 ( .A(y[2444]), .B(x[2444]), .Z(n4120) );
  NAND U7981 ( .A(n19587), .B(n4120), .Z(n24241) );
  AND U7982 ( .A(n19594), .B(n24241), .Z(n9103) );
  XNOR U7983 ( .A(y[2444]), .B(x[2444]), .Z(n4122) );
  NANDN U7984 ( .A(y[2443]), .B(x[2443]), .Z(n4121) );
  AND U7985 ( .A(n4122), .B(n4121), .Z(n19592) );
  NANDN U7986 ( .A(y[2442]), .B(x[2442]), .Z(n19585) );
  NAND U7987 ( .A(n19592), .B(n19585), .Z(n24242) );
  ANDN U7988 ( .B(y[2441]), .A(x[2441]), .Z(n19583) );
  ANDN U7989 ( .B(y[2442]), .A(x[2442]), .Z(n19590) );
  NOR U7990 ( .A(n19583), .B(n19590), .Z(n27817) );
  NANDN U7991 ( .A(y[2440]), .B(x[2440]), .Z(n12694) );
  NANDN U7992 ( .A(y[2441]), .B(x[2441]), .Z(n24244) );
  NAND U7993 ( .A(n12694), .B(n24244), .Z(n9099) );
  NANDN U7994 ( .A(x[2439]), .B(y[2439]), .Z(n4123) );
  NANDN U7995 ( .A(x[2440]), .B(y[2440]), .Z(n12692) );
  AND U7996 ( .A(n4123), .B(n12692), .Z(n12696) );
  NANDN U7997 ( .A(x[2437]), .B(y[2437]), .Z(n12700) );
  NANDN U7998 ( .A(x[2436]), .B(y[2436]), .Z(n12699) );
  NANDN U7999 ( .A(y[2435]), .B(x[2435]), .Z(n4125) );
  NANDN U8000 ( .A(y[2436]), .B(x[2436]), .Z(n4124) );
  NAND U8001 ( .A(n4125), .B(n4124), .Z(n12701) );
  NANDN U8002 ( .A(y[2433]), .B(x[2433]), .Z(n4126) );
  ANDN U8003 ( .B(x[2434]), .A(y[2434]), .Z(n9084) );
  ANDN U8004 ( .B(n4126), .A(n9084), .Z(n12705) );
  NANDN U8005 ( .A(y[2432]), .B(x[2432]), .Z(n4127) );
  AND U8006 ( .A(n12705), .B(n4127), .Z(n27811) );
  ANDN U8007 ( .B(y[2432]), .A(x[2432]), .Z(n12704) );
  ANDN U8008 ( .B(y[2431]), .A(x[2431]), .Z(n27810) );
  NANDN U8009 ( .A(y[2430]), .B(x[2430]), .Z(n12709) );
  NANDN U8010 ( .A(y[2431]), .B(x[2431]), .Z(n12706) );
  AND U8011 ( .A(n12709), .B(n12706), .Z(n27809) );
  ANDN U8012 ( .B(y[2429]), .A(x[2429]), .Z(n12710) );
  ANDN U8013 ( .B(x[2428]), .A(y[2428]), .Z(n12712) );
  NANDN U8014 ( .A(x[2427]), .B(y[2427]), .Z(n12714) );
  NANDN U8015 ( .A(x[2428]), .B(y[2428]), .Z(n12711) );
  NANDN U8016 ( .A(y[2426]), .B(x[2426]), .Z(n12715) );
  NANDN U8017 ( .A(y[2427]), .B(x[2427]), .Z(n12713) );
  NAND U8018 ( .A(n12715), .B(n12713), .Z(n27802) );
  ANDN U8019 ( .B(y[2426]), .A(x[2426]), .Z(n19565) );
  NANDN U8020 ( .A(x[2425]), .B(y[2425]), .Z(n4129) );
  NANDN U8021 ( .A(x[2424]), .B(y[2424]), .Z(n4128) );
  NAND U8022 ( .A(n4129), .B(n4128), .Z(n19561) );
  NANDN U8023 ( .A(y[2425]), .B(x[2425]), .Z(n12716) );
  NAND U8024 ( .A(n19561), .B(n12716), .Z(n4130) );
  NANDN U8025 ( .A(n19565), .B(n4130), .Z(n24245) );
  NANDN U8026 ( .A(y[2424]), .B(x[2424]), .Z(n4132) );
  NANDN U8027 ( .A(y[2423]), .B(x[2423]), .Z(n4131) );
  AND U8028 ( .A(n4132), .B(n4131), .Z(n19554) );
  AND U8029 ( .A(n19554), .B(n12716), .Z(n27801) );
  ANDN U8030 ( .B(y[2423]), .A(x[2423]), .Z(n9066) );
  NANDN U8031 ( .A(y[2422]), .B(x[2422]), .Z(n19555) );
  OR U8032 ( .A(n9066), .B(n19555), .Z(n4133) );
  AND U8033 ( .A(n27801), .B(n4133), .Z(n9071) );
  NANDN U8034 ( .A(y[2420]), .B(x[2420]), .Z(n27799) );
  NANDN U8035 ( .A(y[2421]), .B(x[2421]), .Z(n19556) );
  AND U8036 ( .A(n27799), .B(n19556), .Z(n9065) );
  NANDN U8037 ( .A(x[2420]), .B(y[2420]), .Z(n4135) );
  NANDN U8038 ( .A(x[2419]), .B(y[2419]), .Z(n4134) );
  NAND U8039 ( .A(n4135), .B(n4134), .Z(n27798) );
  NANDN U8040 ( .A(y[2418]), .B(x[2418]), .Z(n4136) );
  NANDN U8041 ( .A(y[2419]), .B(x[2419]), .Z(n24247) );
  AND U8042 ( .A(n4136), .B(n24247), .Z(n4140) );
  ANDN U8043 ( .B(y[2417]), .A(x[2417]), .Z(n27795) );
  ANDN U8044 ( .B(y[2418]), .A(x[2418]), .Z(n24248) );
  OR U8045 ( .A(n27795), .B(n24248), .Z(n4137) );
  NAND U8046 ( .A(n4140), .B(n4137), .Z(n4138) );
  NANDN U8047 ( .A(n27798), .B(n4138), .Z(n19549) );
  NANDN U8048 ( .A(y[2417]), .B(x[2417]), .Z(n4139) );
  AND U8049 ( .A(n4140), .B(n4139), .Z(n27797) );
  ANDN U8050 ( .B(y[2416]), .A(x[2416]), .Z(n27794) );
  NANDN U8051 ( .A(y[2416]), .B(x[2416]), .Z(n4142) );
  NANDN U8052 ( .A(y[2415]), .B(x[2415]), .Z(n4141) );
  AND U8053 ( .A(n4142), .B(n4141), .Z(n27793) );
  NANDN U8054 ( .A(x[2414]), .B(y[2414]), .Z(n4144) );
  NANDN U8055 ( .A(x[2415]), .B(y[2415]), .Z(n4143) );
  NAND U8056 ( .A(n4144), .B(n4143), .Z(n27792) );
  NANDN U8057 ( .A(y[2414]), .B(x[2414]), .Z(n4146) );
  NANDN U8058 ( .A(y[2413]), .B(x[2413]), .Z(n4145) );
  AND U8059 ( .A(n4146), .B(n4145), .Z(n27791) );
  NANDN U8060 ( .A(x[2412]), .B(y[2412]), .Z(n4148) );
  NANDN U8061 ( .A(x[2413]), .B(y[2413]), .Z(n4147) );
  NAND U8062 ( .A(n4148), .B(n4147), .Z(n27790) );
  NANDN U8063 ( .A(y[2412]), .B(x[2412]), .Z(n4150) );
  NANDN U8064 ( .A(y[2411]), .B(x[2411]), .Z(n4149) );
  AND U8065 ( .A(n4150), .B(n4149), .Z(n27789) );
  NANDN U8066 ( .A(x[2410]), .B(y[2410]), .Z(n4152) );
  NANDN U8067 ( .A(x[2411]), .B(y[2411]), .Z(n4151) );
  NAND U8068 ( .A(n4152), .B(n4151), .Z(n27786) );
  NANDN U8069 ( .A(y[2410]), .B(x[2410]), .Z(n27787) );
  NANDN U8070 ( .A(y[2409]), .B(x[2409]), .Z(n4153) );
  AND U8071 ( .A(n27787), .B(n4153), .Z(n4157) );
  ANDN U8072 ( .B(y[2408]), .A(x[2408]), .Z(n27783) );
  ANDN U8073 ( .B(y[2409]), .A(x[2409]), .Z(n27788) );
  OR U8074 ( .A(n27783), .B(n27788), .Z(n4154) );
  NAND U8075 ( .A(n4157), .B(n4154), .Z(n4155) );
  NANDN U8076 ( .A(n27786), .B(n4155), .Z(n19541) );
  NANDN U8077 ( .A(y[2408]), .B(x[2408]), .Z(n4156) );
  AND U8078 ( .A(n4157), .B(n4156), .Z(n27785) );
  NANDN U8079 ( .A(y[2406]), .B(x[2406]), .Z(n4158) );
  ANDN U8080 ( .B(x[2407]), .A(y[2407]), .Z(n12718) );
  ANDN U8081 ( .B(n4158), .A(n12718), .Z(n27782) );
  NANDN U8082 ( .A(y[2405]), .B(x[2405]), .Z(n4160) );
  NANDN U8083 ( .A(y[2404]), .B(x[2404]), .Z(n4159) );
  NAND U8084 ( .A(n4160), .B(n4159), .Z(n19535) );
  NANDN U8085 ( .A(x[2404]), .B(y[2404]), .Z(n12720) );
  NANDN U8086 ( .A(x[2403]), .B(y[2403]), .Z(n4161) );
  AND U8087 ( .A(n12720), .B(n4161), .Z(n9046) );
  ANDN U8088 ( .B(x[2402]), .A(y[2402]), .Z(n19529) );
  ANDN U8089 ( .B(x[2403]), .A(y[2403]), .Z(n12721) );
  OR U8090 ( .A(n19529), .B(n12721), .Z(n4162) );
  NAND U8091 ( .A(n9046), .B(n4162), .Z(n4163) );
  NANDN U8092 ( .A(n19535), .B(n4163), .Z(n27780) );
  NANDN U8093 ( .A(x[2401]), .B(y[2401]), .Z(n12722) );
  ANDN U8094 ( .B(x[2401]), .A(y[2401]), .Z(n27775) );
  NANDN U8095 ( .A(y[2400]), .B(x[2400]), .Z(n9040) );
  XNOR U8096 ( .A(y[2400]), .B(x[2400]), .Z(n4165) );
  NANDN U8097 ( .A(x[2399]), .B(y[2399]), .Z(n4164) );
  NAND U8098 ( .A(n4165), .B(n4164), .Z(n4166) );
  NAND U8099 ( .A(n9040), .B(n4166), .Z(n12723) );
  NANDN U8100 ( .A(y[2396]), .B(x[2396]), .Z(n4168) );
  NANDN U8101 ( .A(y[2397]), .B(x[2397]), .Z(n4167) );
  NAND U8102 ( .A(n4168), .B(n4167), .Z(n19523) );
  NANDN U8103 ( .A(x[2395]), .B(y[2395]), .Z(n4169) );
  ANDN U8104 ( .B(y[2396]), .A(x[2396]), .Z(n19517) );
  ANDN U8105 ( .B(n4169), .A(n19517), .Z(n27771) );
  ANDN U8106 ( .B(x[2394]), .A(y[2394]), .Z(n19513) );
  NANDN U8107 ( .A(y[2395]), .B(x[2395]), .Z(n4170) );
  NANDN U8108 ( .A(n19513), .B(n4170), .Z(n27770) );
  NANDN U8109 ( .A(x[2393]), .B(y[2393]), .Z(n19510) );
  NANDN U8110 ( .A(x[2394]), .B(y[2394]), .Z(n19516) );
  AND U8111 ( .A(n19510), .B(n19516), .Z(n27769) );
  ANDN U8112 ( .B(x[2393]), .A(y[2393]), .Z(n27768) );
  ANDN U8113 ( .B(y[2390]), .A(x[2390]), .Z(n19506) );
  NANDN U8114 ( .A(x[2389]), .B(y[2389]), .Z(n12725) );
  NANDN U8115 ( .A(n19506), .B(n12725), .Z(n27766) );
  NANDN U8116 ( .A(y[2388]), .B(x[2388]), .Z(n12727) );
  NANDN U8117 ( .A(y[2389]), .B(x[2389]), .Z(n19502) );
  AND U8118 ( .A(n12727), .B(n19502), .Z(n27765) );
  NANDN U8119 ( .A(x[2387]), .B(y[2387]), .Z(n12729) );
  NANDN U8120 ( .A(x[2388]), .B(y[2388]), .Z(n12726) );
  NAND U8121 ( .A(n12729), .B(n12726), .Z(n27763) );
  NANDN U8122 ( .A(y[2386]), .B(x[2386]), .Z(n12731) );
  NANDN U8123 ( .A(y[2387]), .B(x[2387]), .Z(n12728) );
  AND U8124 ( .A(n12731), .B(n12728), .Z(n27762) );
  NANDN U8125 ( .A(x[2386]), .B(y[2386]), .Z(n12730) );
  NANDN U8126 ( .A(x[2385]), .B(y[2385]), .Z(n4172) );
  NANDN U8127 ( .A(x[2384]), .B(y[2384]), .Z(n4171) );
  AND U8128 ( .A(n4172), .B(n4171), .Z(n19493) );
  NANDN U8129 ( .A(y[2385]), .B(x[2385]), .Z(n12732) );
  NANDN U8130 ( .A(n19493), .B(n12732), .Z(n4173) );
  AND U8131 ( .A(n12730), .B(n4173), .Z(n27761) );
  NANDN U8132 ( .A(x[2382]), .B(y[2382]), .Z(n4174) );
  NANDN U8133 ( .A(x[2383]), .B(y[2383]), .Z(n9017) );
  AND U8134 ( .A(n4174), .B(n9017), .Z(n27759) );
  NANDN U8135 ( .A(x[2380]), .B(y[2380]), .Z(n4175) );
  NANDN U8136 ( .A(x[2381]), .B(y[2381]), .Z(n9012) );
  AND U8137 ( .A(n4175), .B(n9012), .Z(n27757) );
  NANDN U8138 ( .A(x[2379]), .B(y[2379]), .Z(n19480) );
  ANDN U8139 ( .B(x[2378]), .A(y[2378]), .Z(n12735) );
  NANDN U8140 ( .A(y[2377]), .B(x[2377]), .Z(n12736) );
  NANDN U8141 ( .A(y[2376]), .B(x[2376]), .Z(n27752) );
  NANDN U8142 ( .A(y[2374]), .B(x[2374]), .Z(n12738) );
  NANDN U8143 ( .A(y[2375]), .B(x[2375]), .Z(n27750) );
  AND U8144 ( .A(n12738), .B(n27750), .Z(n9002) );
  NANDN U8145 ( .A(x[2374]), .B(y[2374]), .Z(n27749) );
  NANDN U8146 ( .A(y[2373]), .B(x[2373]), .Z(n12739) );
  ANDN U8147 ( .B(y[2371]), .A(x[2371]), .Z(n19464) );
  ANDN U8148 ( .B(y[2372]), .A(x[2372]), .Z(n19468) );
  OR U8149 ( .A(n19464), .B(n19468), .Z(n27745) );
  NANDN U8150 ( .A(y[2370]), .B(x[2370]), .Z(n12740) );
  NANDN U8151 ( .A(y[2371]), .B(x[2371]), .Z(n27743) );
  AND U8152 ( .A(n12740), .B(n27743), .Z(n8995) );
  ANDN U8153 ( .B(y[2370]), .A(x[2370]), .Z(n24253) );
  NANDN U8154 ( .A(y[2369]), .B(x[2369]), .Z(n12741) );
  NANDN U8155 ( .A(x[2368]), .B(y[2368]), .Z(n12743) );
  NANDN U8156 ( .A(x[2367]), .B(y[2367]), .Z(n19457) );
  AND U8157 ( .A(n12743), .B(n19457), .Z(n8989) );
  ANDN U8158 ( .B(x[2367]), .A(y[2367]), .Z(n12744) );
  ANDN U8159 ( .B(y[2365]), .A(x[2365]), .Z(n27738) );
  NANDN U8160 ( .A(y[2365]), .B(x[2365]), .Z(n12746) );
  ANDN U8161 ( .B(x[2364]), .A(y[2364]), .Z(n19449) );
  ANDN U8162 ( .B(n12746), .A(n19449), .Z(n27737) );
  NANDN U8163 ( .A(x[2363]), .B(y[2363]), .Z(n19447) );
  NANDN U8164 ( .A(x[2364]), .B(y[2364]), .Z(n19452) );
  NAND U8165 ( .A(n19447), .B(n19452), .Z(n27736) );
  ANDN U8166 ( .B(x[2362]), .A(y[2362]), .Z(n19445) );
  ANDN U8167 ( .B(x[2363]), .A(y[2363]), .Z(n24255) );
  NOR U8168 ( .A(n19445), .B(n24255), .Z(n8981) );
  NANDN U8169 ( .A(y[2356]), .B(x[2356]), .Z(n4176) );
  NANDN U8170 ( .A(y[2357]), .B(x[2357]), .Z(n27729) );
  AND U8171 ( .A(n4176), .B(n27729), .Z(n8966) );
  XNOR U8172 ( .A(x[2356]), .B(y[2356]), .Z(n12749) );
  ANDN U8173 ( .B(y[2353]), .A(x[2353]), .Z(n19425) );
  ANDN U8174 ( .B(y[2354]), .A(x[2354]), .Z(n19429) );
  NOR U8175 ( .A(n19425), .B(n19429), .Z(n27724) );
  NANDN U8176 ( .A(y[2353]), .B(x[2353]), .Z(n27723) );
  ANDN U8177 ( .B(x[2350]), .A(y[2350]), .Z(n12752) );
  NANDN U8178 ( .A(x[2350]), .B(y[2350]), .Z(n19421) );
  NANDN U8179 ( .A(y[2349]), .B(x[2349]), .Z(n12753) );
  ANDN U8180 ( .B(x[2348]), .A(y[2348]), .Z(n12756) );
  ANDN U8181 ( .B(n12753), .A(n12756), .Z(n8951) );
  ANDN U8182 ( .B(y[2347]), .A(x[2347]), .Z(n12758) );
  NANDN U8183 ( .A(x[2345]), .B(y[2345]), .Z(n12762) );
  NANDN U8184 ( .A(x[2343]), .B(y[2343]), .Z(n12767) );
  ANDN U8185 ( .B(y[2341]), .A(x[2341]), .Z(n12770) );
  ANDN U8186 ( .B(y[2339]), .A(x[2339]), .Z(n19402) );
  ANDN U8187 ( .B(x[2338]), .A(y[2338]), .Z(n12773) );
  ANDN U8188 ( .B(x[2339]), .A(y[2339]), .Z(n19407) );
  NOR U8189 ( .A(n12773), .B(n19407), .Z(n27693) );
  NANDN U8190 ( .A(x[2338]), .B(y[2338]), .Z(n19403) );
  ANDN U8191 ( .B(y[2337]), .A(x[2337]), .Z(n19397) );
  ANDN U8192 ( .B(n19403), .A(n19397), .Z(n27692) );
  ANDN U8193 ( .B(x[2337]), .A(y[2337]), .Z(n12772) );
  NANDN U8194 ( .A(y[2336]), .B(x[2336]), .Z(n12775) );
  NANDN U8195 ( .A(n12772), .B(n12775), .Z(n27690) );
  NANDN U8196 ( .A(x[2336]), .B(y[2336]), .Z(n19398) );
  ANDN U8197 ( .B(x[2334]), .A(y[2334]), .Z(n12778) );
  NANDN U8198 ( .A(y[2332]), .B(x[2332]), .Z(n27675) );
  NANDN U8199 ( .A(x[2331]), .B(y[2331]), .Z(n19385) );
  ANDN U8200 ( .B(y[2332]), .A(x[2332]), .Z(n19390) );
  ANDN U8201 ( .B(n19385), .A(n19390), .Z(n27676) );
  ANDN U8202 ( .B(x[2331]), .A(y[2331]), .Z(n12780) );
  XNOR U8203 ( .A(x[2330]), .B(y[2330]), .Z(n12782) );
  NANDN U8204 ( .A(y[2329]), .B(x[2329]), .Z(n12781) );
  ANDN U8205 ( .B(x[2328]), .A(y[2328]), .Z(n27669) );
  ANDN U8206 ( .B(n12781), .A(n27669), .Z(n8914) );
  NANDN U8207 ( .A(y[2327]), .B(x[2327]), .Z(n4178) );
  NANDN U8208 ( .A(y[2326]), .B(x[2326]), .Z(n4177) );
  AND U8209 ( .A(n4178), .B(n4177), .Z(n19376) );
  NANDN U8210 ( .A(x[2326]), .B(y[2326]), .Z(n19375) );
  NANDN U8211 ( .A(x[2325]), .B(y[2325]), .Z(n4179) );
  NAND U8212 ( .A(n19375), .B(n4179), .Z(n12783) );
  NANDN U8213 ( .A(y[2324]), .B(x[2324]), .Z(n27667) );
  NANDN U8214 ( .A(x[2323]), .B(y[2323]), .Z(n12786) );
  NANDN U8215 ( .A(x[2324]), .B(y[2324]), .Z(n12784) );
  NAND U8216 ( .A(n12786), .B(n12784), .Z(n27666) );
  NANDN U8217 ( .A(y[2322]), .B(x[2322]), .Z(n12789) );
  NANDN U8218 ( .A(y[2323]), .B(x[2323]), .Z(n12785) );
  AND U8219 ( .A(n12789), .B(n12785), .Z(n27665) );
  NANDN U8220 ( .A(x[2321]), .B(y[2321]), .Z(n19365) );
  NANDN U8221 ( .A(x[2322]), .B(y[2322]), .Z(n12787) );
  NAND U8222 ( .A(n19365), .B(n12787), .Z(n27664) );
  NANDN U8223 ( .A(y[2321]), .B(x[2321]), .Z(n12788) );
  ANDN U8224 ( .B(x[2320]), .A(y[2320]), .Z(n19363) );
  ANDN U8225 ( .B(n12788), .A(n19363), .Z(n27663) );
  ANDN U8226 ( .B(y[2317]), .A(x[2317]), .Z(n27660) );
  NANDN U8227 ( .A(y[2316]), .B(x[2316]), .Z(n4180) );
  ANDN U8228 ( .B(x[2317]), .A(y[2317]), .Z(n19356) );
  ANDN U8229 ( .B(n4180), .A(n19356), .Z(n27659) );
  ANDN U8230 ( .B(y[2315]), .A(x[2315]), .Z(n19349) );
  NANDN U8231 ( .A(x[2316]), .B(y[2316]), .Z(n19355) );
  NANDN U8232 ( .A(n19349), .B(n19355), .Z(n27657) );
  NANDN U8233 ( .A(y[2314]), .B(x[2314]), .Z(n19347) );
  ANDN U8234 ( .B(x[2315]), .A(y[2315]), .Z(n19352) );
  ANDN U8235 ( .B(n19347), .A(n19352), .Z(n27656) );
  ANDN U8236 ( .B(y[2314]), .A(x[2314]), .Z(n27655) );
  ANDN U8237 ( .B(y[2312]), .A(x[2312]), .Z(n19344) );
  NANDN U8238 ( .A(y[2312]), .B(x[2312]), .Z(n4182) );
  NANDN U8239 ( .A(y[2311]), .B(x[2311]), .Z(n4181) );
  AND U8240 ( .A(n4182), .B(n4181), .Z(n24258) );
  NANDN U8241 ( .A(x[2305]), .B(y[2305]), .Z(n12797) );
  NANDN U8242 ( .A(x[2306]), .B(y[2306]), .Z(n12794) );
  NAND U8243 ( .A(n12797), .B(n12794), .Z(n24261) );
  NANDN U8244 ( .A(y[2305]), .B(x[2305]), .Z(n24262) );
  NANDN U8245 ( .A(y[2304]), .B(x[2304]), .Z(n12798) );
  ANDN U8246 ( .B(y[2304]), .A(x[2304]), .Z(n12796) );
  NANDN U8247 ( .A(y[2303]), .B(x[2303]), .Z(n12799) );
  NANDN U8248 ( .A(y[2302]), .B(x[2302]), .Z(n12802) );
  AND U8249 ( .A(n12799), .B(n12802), .Z(n8871) );
  NANDN U8250 ( .A(x[2302]), .B(y[2302]), .Z(n12801) );
  NANDN U8251 ( .A(x[2301]), .B(y[2301]), .Z(n12805) );
  NANDN U8252 ( .A(y[2300]), .B(x[2300]), .Z(n12809) );
  NANDN U8253 ( .A(x[2300]), .B(y[2300]), .Z(n12804) );
  ANDN U8254 ( .B(y[2299]), .A(x[2299]), .Z(n12806) );
  ANDN U8255 ( .B(n12804), .A(n12806), .Z(n8865) );
  NANDN U8256 ( .A(x[2298]), .B(y[2298]), .Z(n4184) );
  NANDN U8257 ( .A(x[2297]), .B(y[2297]), .Z(n4183) );
  AND U8258 ( .A(n4184), .B(n4183), .Z(n19318) );
  NANDN U8259 ( .A(y[2296]), .B(x[2296]), .Z(n4185) );
  NANDN U8260 ( .A(y[2297]), .B(x[2297]), .Z(n19320) );
  AND U8261 ( .A(n4185), .B(n19320), .Z(n27641) );
  NANDN U8262 ( .A(y[2295]), .B(x[2295]), .Z(n19314) );
  ANDN U8263 ( .B(x[2294]), .A(y[2294]), .Z(n19309) );
  ANDN U8264 ( .B(n19314), .A(n19309), .Z(n27639) );
  NANDN U8265 ( .A(x[2293]), .B(y[2293]), .Z(n12811) );
  NANDN U8266 ( .A(x[2294]), .B(y[2294]), .Z(n12810) );
  NAND U8267 ( .A(n12811), .B(n12810), .Z(n27638) );
  NANDN U8268 ( .A(y[2292]), .B(x[2292]), .Z(n19304) );
  ANDN U8269 ( .B(x[2293]), .A(y[2293]), .Z(n19310) );
  ANDN U8270 ( .B(n19304), .A(n19310), .Z(n27637) );
  ANDN U8271 ( .B(y[2291]), .A(x[2291]), .Z(n19300) );
  NANDN U8272 ( .A(x[2292]), .B(y[2292]), .Z(n27636) );
  ANDN U8273 ( .B(x[2290]), .A(y[2290]), .Z(n12812) );
  ANDN U8274 ( .B(x[2291]), .A(y[2291]), .Z(n27635) );
  ANDN U8275 ( .B(y[2290]), .A(x[2290]), .Z(n19301) );
  NANDN U8276 ( .A(x[2287]), .B(y[2287]), .Z(n12814) );
  ANDN U8277 ( .B(y[2288]), .A(x[2288]), .Z(n19297) );
  ANDN U8278 ( .B(n12814), .A(n19297), .Z(n27630) );
  NANDN U8279 ( .A(x[2286]), .B(y[2286]), .Z(n27626) );
  NANDN U8280 ( .A(x[2285]), .B(y[2285]), .Z(n19289) );
  AND U8281 ( .A(n27626), .B(n19289), .Z(n8860) );
  ANDN U8282 ( .B(x[2285]), .A(y[2285]), .Z(n12815) );
  NANDN U8283 ( .A(y[2284]), .B(x[2284]), .Z(n27622) );
  NANDN U8284 ( .A(x[2283]), .B(y[2283]), .Z(n27623) );
  NANDN U8285 ( .A(y[2282]), .B(x[2282]), .Z(n19281) );
  NANDN U8286 ( .A(y[2281]), .B(x[2281]), .Z(n19282) );
  NANDN U8287 ( .A(y[2280]), .B(x[2280]), .Z(n12819) );
  AND U8288 ( .A(n19282), .B(n12819), .Z(n8851) );
  NANDN U8289 ( .A(y[2278]), .B(x[2278]), .Z(n19273) );
  ANDN U8290 ( .B(x[2279]), .A(y[2279]), .Z(n19277) );
  ANDN U8291 ( .B(n19273), .A(n19277), .Z(n27619) );
  NANDN U8292 ( .A(x[2277]), .B(y[2277]), .Z(n4187) );
  NANDN U8293 ( .A(x[2278]), .B(y[2278]), .Z(n4186) );
  NAND U8294 ( .A(n4187), .B(n4186), .Z(n27618) );
  NANDN U8295 ( .A(y[2277]), .B(x[2277]), .Z(n4189) );
  NANDN U8296 ( .A(y[2276]), .B(x[2276]), .Z(n4188) );
  AND U8297 ( .A(n4189), .B(n4188), .Z(n24267) );
  NANDN U8298 ( .A(x[2274]), .B(y[2274]), .Z(n19267) );
  ANDN U8299 ( .B(y[2273]), .A(x[2273]), .Z(n27614) );
  ANDN U8300 ( .B(n19267), .A(n27614), .Z(n8840) );
  NANDN U8301 ( .A(y[2273]), .B(x[2273]), .Z(n4191) );
  NANDN U8302 ( .A(y[2272]), .B(x[2272]), .Z(n4190) );
  AND U8303 ( .A(n4191), .B(n4190), .Z(n12823) );
  NANDN U8304 ( .A(x[2271]), .B(y[2271]), .Z(n4192) );
  ANDN U8305 ( .B(y[2272]), .A(x[2272]), .Z(n12821) );
  ANDN U8306 ( .B(n4192), .A(n12821), .Z(n4196) );
  NANDN U8307 ( .A(y[2270]), .B(x[2270]), .Z(n12824) );
  NANDN U8308 ( .A(y[2271]), .B(x[2271]), .Z(n12820) );
  NAND U8309 ( .A(n12824), .B(n12820), .Z(n4193) );
  NAND U8310 ( .A(n4196), .B(n4193), .Z(n4194) );
  NAND U8311 ( .A(n12823), .B(n4194), .Z(n27613) );
  NANDN U8312 ( .A(x[2270]), .B(y[2270]), .Z(n4195) );
  AND U8313 ( .A(n4196), .B(n4195), .Z(n27612) );
  NANDN U8314 ( .A(x[2268]), .B(y[2268]), .Z(n4198) );
  NANDN U8315 ( .A(x[2269]), .B(y[2269]), .Z(n4197) );
  AND U8316 ( .A(n4198), .B(n4197), .Z(n27610) );
  XNOR U8317 ( .A(x[2268]), .B(y[2268]), .Z(n4199) );
  NANDN U8318 ( .A(y[2267]), .B(x[2267]), .Z(n12826) );
  AND U8319 ( .A(n4199), .B(n12826), .Z(n4201) );
  NANDN U8320 ( .A(y[2266]), .B(x[2266]), .Z(n12827) );
  NANDN U8321 ( .A(x[2267]), .B(y[2267]), .Z(n4203) );
  NANDN U8322 ( .A(n12827), .B(n4203), .Z(n4200) );
  NAND U8323 ( .A(n4201), .B(n4200), .Z(n27609) );
  NANDN U8324 ( .A(x[2266]), .B(y[2266]), .Z(n4202) );
  AND U8325 ( .A(n4203), .B(n4202), .Z(n27608) );
  NANDN U8326 ( .A(y[2265]), .B(x[2265]), .Z(n27607) );
  NANDN U8327 ( .A(x[2265]), .B(y[2265]), .Z(n4205) );
  NANDN U8328 ( .A(x[2264]), .B(y[2264]), .Z(n4204) );
  AND U8329 ( .A(n4205), .B(n4204), .Z(n27606) );
  NANDN U8330 ( .A(y[2264]), .B(x[2264]), .Z(n4207) );
  NANDN U8331 ( .A(y[2263]), .B(x[2263]), .Z(n4206) );
  AND U8332 ( .A(n4207), .B(n4206), .Z(n12828) );
  NANDN U8333 ( .A(x[2263]), .B(y[2263]), .Z(n4209) );
  NANDN U8334 ( .A(x[2262]), .B(y[2262]), .Z(n4208) );
  AND U8335 ( .A(n4209), .B(n4208), .Z(n19249) );
  NANDN U8336 ( .A(x[2261]), .B(y[2261]), .Z(n12830) );
  NANDN U8337 ( .A(y[2262]), .B(x[2262]), .Z(n8826) );
  NANDN U8338 ( .A(n12830), .B(n8826), .Z(n4210) );
  NAND U8339 ( .A(n19249), .B(n4210), .Z(n24268) );
  NANDN U8340 ( .A(y[2260]), .B(x[2260]), .Z(n12831) );
  NANDN U8341 ( .A(x[2259]), .B(y[2259]), .Z(n12834) );
  NANDN U8342 ( .A(y[2258]), .B(x[2258]), .Z(n12835) );
  ANDN U8343 ( .B(y[2257]), .A(x[2257]), .Z(n12837) );
  NANDN U8344 ( .A(y[2257]), .B(x[2257]), .Z(n12836) );
  NANDN U8345 ( .A(x[2255]), .B(y[2255]), .Z(n19237) );
  NANDN U8346 ( .A(x[2256]), .B(y[2256]), .Z(n12838) );
  NAND U8347 ( .A(n19237), .B(n12838), .Z(n8816) );
  NANDN U8348 ( .A(y[2254]), .B(x[2254]), .Z(n4212) );
  NANDN U8349 ( .A(y[2255]), .B(x[2255]), .Z(n4211) );
  NAND U8350 ( .A(n4212), .B(n4211), .Z(n12839) );
  NANDN U8351 ( .A(y[2252]), .B(x[2252]), .Z(n4213) );
  NANDN U8352 ( .A(y[2253]), .B(x[2253]), .Z(n19239) );
  AND U8353 ( .A(n4213), .B(n19239), .Z(n27596) );
  NANDN U8354 ( .A(y[2250]), .B(x[2250]), .Z(n4214) );
  ANDN U8355 ( .B(x[2251]), .A(y[2251]), .Z(n12842) );
  ANDN U8356 ( .B(n4214), .A(n12842), .Z(n27594) );
  ANDN U8357 ( .B(y[2249]), .A(x[2249]), .Z(n19229) );
  NANDN U8358 ( .A(x[2250]), .B(y[2250]), .Z(n12841) );
  NANDN U8359 ( .A(n19229), .B(n12841), .Z(n27593) );
  NANDN U8360 ( .A(y[2248]), .B(x[2248]), .Z(n19224) );
  NANDN U8361 ( .A(y[2249]), .B(x[2249]), .Z(n19231) );
  AND U8362 ( .A(n19224), .B(n19231), .Z(n24270) );
  ANDN U8363 ( .B(y[2247]), .A(x[2247]), .Z(n12845) );
  ANDN U8364 ( .B(x[2246]), .A(y[2246]), .Z(n12847) );
  NANDN U8365 ( .A(x[2245]), .B(y[2245]), .Z(n19219) );
  ANDN U8366 ( .B(x[2244]), .A(y[2244]), .Z(n19217) );
  NANDN U8367 ( .A(x[2243]), .B(y[2243]), .Z(n4216) );
  NANDN U8368 ( .A(x[2244]), .B(y[2244]), .Z(n4215) );
  NAND U8369 ( .A(n4216), .B(n4215), .Z(n19216) );
  ANDN U8370 ( .B(x[2240]), .A(y[2240]), .Z(n8786) );
  NANDN U8371 ( .A(y[2239]), .B(x[2239]), .Z(n4217) );
  NANDN U8372 ( .A(n8786), .B(n4217), .Z(n19212) );
  IV U8373 ( .A(n19212), .Z(n27584) );
  NANDN U8374 ( .A(y[2238]), .B(x[2238]), .Z(n19206) );
  ANDN U8375 ( .B(y[2237]), .A(x[2237]), .Z(n12851) );
  NANDN U8376 ( .A(y[2236]), .B(x[2236]), .Z(n19202) );
  ANDN U8377 ( .B(y[2235]), .A(x[2235]), .Z(n12853) );
  NANDN U8378 ( .A(y[2235]), .B(x[2235]), .Z(n19203) );
  NANDN U8379 ( .A(x[2234]), .B(y[2234]), .Z(n12854) );
  ANDN U8380 ( .B(y[2233]), .A(x[2233]), .Z(n12858) );
  ANDN U8381 ( .B(n12854), .A(n12858), .Z(n8771) );
  NANDN U8382 ( .A(x[2232]), .B(y[2232]), .Z(n4219) );
  NANDN U8383 ( .A(x[2231]), .B(y[2231]), .Z(n4218) );
  AND U8384 ( .A(n4219), .B(n4218), .Z(n12859) );
  NANDN U8385 ( .A(y[2230]), .B(x[2230]), .Z(n4220) );
  NANDN U8386 ( .A(y[2231]), .B(x[2231]), .Z(n12860) );
  AND U8387 ( .A(n4220), .B(n12860), .Z(n27576) );
  NANDN U8388 ( .A(x[2229]), .B(y[2229]), .Z(n24271) );
  ANDN U8389 ( .B(x[2228]), .A(y[2228]), .Z(n12863) );
  NANDN U8390 ( .A(y[2229]), .B(x[2229]), .Z(n12867) );
  NANDN U8391 ( .A(n12863), .B(n12867), .Z(n24272) );
  NANDN U8392 ( .A(x[2228]), .B(y[2228]), .Z(n12862) );
  NANDN U8393 ( .A(x[2227]), .B(y[2227]), .Z(n4221) );
  AND U8394 ( .A(n12862), .B(n4221), .Z(n27575) );
  NANDN U8395 ( .A(x[2225]), .B(y[2225]), .Z(n12870) );
  NANDN U8396 ( .A(x[2226]), .B(y[2226]), .Z(n24273) );
  AND U8397 ( .A(n12870), .B(n24273), .Z(n8759) );
  NANDN U8398 ( .A(x[2224]), .B(y[2224]), .Z(n12871) );
  NANDN U8399 ( .A(y[2223]), .B(x[2223]), .Z(n4223) );
  NANDN U8400 ( .A(y[2224]), .B(x[2224]), .Z(n4222) );
  NAND U8401 ( .A(n4223), .B(n4222), .Z(n27569) );
  NANDN U8402 ( .A(x[2223]), .B(y[2223]), .Z(n4225) );
  NANDN U8403 ( .A(x[2222]), .B(y[2222]), .Z(n4224) );
  AND U8404 ( .A(n4225), .B(n4224), .Z(n19187) );
  NANDN U8405 ( .A(x[2221]), .B(y[2221]), .Z(n12872) );
  NANDN U8406 ( .A(y[2222]), .B(x[2222]), .Z(n4226) );
  NANDN U8407 ( .A(y[2221]), .B(x[2221]), .Z(n4227) );
  AND U8408 ( .A(n4227), .B(n4226), .Z(n27567) );
  NANDN U8409 ( .A(y[2220]), .B(x[2220]), .Z(n19181) );
  ANDN U8410 ( .B(x[2217]), .A(y[2217]), .Z(n12873) );
  NANDN U8411 ( .A(x[2216]), .B(y[2216]), .Z(n4229) );
  NANDN U8412 ( .A(x[2217]), .B(y[2217]), .Z(n4228) );
  AND U8413 ( .A(n4229), .B(n4228), .Z(n27563) );
  NANDN U8414 ( .A(y[2215]), .B(x[2215]), .Z(n4230) );
  XOR U8415 ( .A(x[2216]), .B(y[2216]), .Z(n8757) );
  ANDN U8416 ( .B(n4230), .A(n8757), .Z(n27562) );
  ANDN U8417 ( .B(x[2214]), .A(y[2214]), .Z(n12874) );
  NANDN U8418 ( .A(x[2213]), .B(y[2213]), .Z(n12877) );
  ANDN U8419 ( .B(x[2212]), .A(y[2212]), .Z(n12879) );
  NANDN U8420 ( .A(x[2209]), .B(y[2209]), .Z(n4232) );
  NANDN U8421 ( .A(x[2210]), .B(y[2210]), .Z(n4231) );
  NAND U8422 ( .A(n4232), .B(n4231), .Z(n12880) );
  NANDN U8423 ( .A(x[2207]), .B(y[2207]), .Z(n27555) );
  NANDN U8424 ( .A(x[2206]), .B(y[2206]), .Z(n12885) );
  NANDN U8425 ( .A(x[2204]), .B(y[2204]), .Z(n4234) );
  NANDN U8426 ( .A(x[2205]), .B(y[2205]), .Z(n4233) );
  AND U8427 ( .A(n4234), .B(n4233), .Z(n24275) );
  NANDN U8428 ( .A(y[2202]), .B(x[2202]), .Z(n12888) );
  ANDN U8429 ( .B(x[2204]), .A(y[2204]), .Z(n8736) );
  NANDN U8430 ( .A(y[2203]), .B(x[2203]), .Z(n4235) );
  NANDN U8431 ( .A(n8736), .B(n4235), .Z(n19158) );
  IV U8432 ( .A(n19158), .Z(n27550) );
  AND U8433 ( .A(n12888), .B(n27550), .Z(n8734) );
  ANDN U8434 ( .B(y[2202]), .A(x[2202]), .Z(n12886) );
  NANDN U8435 ( .A(x[2201]), .B(y[2201]), .Z(n12893) );
  NANDN U8436 ( .A(x[2200]), .B(y[2200]), .Z(n4237) );
  NANDN U8437 ( .A(x[2199]), .B(y[2199]), .Z(n4236) );
  NAND U8438 ( .A(n4237), .B(n4236), .Z(n12891) );
  NANDN U8439 ( .A(y[2199]), .B(x[2199]), .Z(n4239) );
  NANDN U8440 ( .A(y[2198]), .B(x[2198]), .Z(n4238) );
  NAND U8441 ( .A(n4239), .B(n4238), .Z(n19153) );
  NANDN U8442 ( .A(y[2194]), .B(x[2194]), .Z(n19138) );
  ANDN U8443 ( .B(x[2195]), .A(y[2195]), .Z(n19146) );
  ANDN U8444 ( .B(n19138), .A(n19146), .Z(n27543) );
  NANDN U8445 ( .A(x[2193]), .B(y[2193]), .Z(n12896) );
  NANDN U8446 ( .A(x[2194]), .B(y[2194]), .Z(n12895) );
  NAND U8447 ( .A(n12896), .B(n12895), .Z(n27542) );
  NANDN U8448 ( .A(y[2192]), .B(x[2192]), .Z(n19132) );
  NANDN U8449 ( .A(y[2193]), .B(x[2193]), .Z(n19139) );
  NAND U8450 ( .A(n19132), .B(n19139), .Z(n27540) );
  NANDN U8451 ( .A(x[2191]), .B(y[2191]), .Z(n12899) );
  NANDN U8452 ( .A(x[2192]), .B(y[2192]), .Z(n12897) );
  AND U8453 ( .A(n12899), .B(n12897), .Z(n24277) );
  NANDN U8454 ( .A(y[2190]), .B(x[2190]), .Z(n19127) );
  NANDN U8455 ( .A(y[2191]), .B(x[2191]), .Z(n19133) );
  NAND U8456 ( .A(n19127), .B(n19133), .Z(n27539) );
  NANDN U8457 ( .A(x[2190]), .B(y[2190]), .Z(n12898) );
  ANDN U8458 ( .B(y[2189]), .A(x[2189]), .Z(n19124) );
  ANDN U8459 ( .B(n12898), .A(n19124), .Z(n27538) );
  ANDN U8460 ( .B(x[2189]), .A(y[2189]), .Z(n19129) );
  NANDN U8461 ( .A(y[2188]), .B(x[2188]), .Z(n12900) );
  NANDN U8462 ( .A(n19129), .B(n12900), .Z(n27537) );
  NANDN U8463 ( .A(y[2186]), .B(x[2186]), .Z(n12902) );
  NANDN U8464 ( .A(y[2187]), .B(x[2187]), .Z(n24278) );
  AND U8465 ( .A(n12902), .B(n24278), .Z(n27536) );
  ANDN U8466 ( .B(y[2185]), .A(x[2185]), .Z(n12903) );
  NANDN U8467 ( .A(y[2184]), .B(x[2184]), .Z(n19110) );
  NANDN U8468 ( .A(y[2185]), .B(x[2185]), .Z(n12901) );
  AND U8469 ( .A(n19110), .B(n12901), .Z(n24281) );
  NANDN U8470 ( .A(x[2184]), .B(y[2184]), .Z(n27534) );
  NANDN U8471 ( .A(x[2183]), .B(y[2183]), .Z(n19112) );
  NAND U8472 ( .A(n27534), .B(n19112), .Z(n8708) );
  XNOR U8473 ( .A(y[2180]), .B(x[2180]), .Z(n12909) );
  NANDN U8474 ( .A(y[2178]), .B(x[2178]), .Z(n19100) );
  NANDN U8475 ( .A(y[2179]), .B(x[2179]), .Z(n12908) );
  AND U8476 ( .A(n19100), .B(n12908), .Z(n24282) );
  ANDN U8477 ( .B(y[2177]), .A(x[2177]), .Z(n19098) );
  NANDN U8478 ( .A(x[2178]), .B(y[2178]), .Z(n12911) );
  NANDN U8479 ( .A(n19098), .B(n12911), .Z(n24283) );
  NANDN U8480 ( .A(x[2175]), .B(y[2175]), .Z(n27524) );
  NANDN U8481 ( .A(x[2176]), .B(y[2176]), .Z(n12912) );
  AND U8482 ( .A(n27524), .B(n12912), .Z(n8692) );
  ANDN U8483 ( .B(x[2174]), .A(y[2174]), .Z(n19088) );
  ANDN U8484 ( .B(y[2173]), .A(x[2173]), .Z(n19087) );
  ANDN U8485 ( .B(y[2174]), .A(x[2174]), .Z(n19094) );
  NOR U8486 ( .A(n19087), .B(n19094), .Z(n27522) );
  ANDN U8487 ( .B(x[2173]), .A(y[2173]), .Z(n19091) );
  NANDN U8488 ( .A(y[2172]), .B(x[2172]), .Z(n12915) );
  NANDN U8489 ( .A(n19091), .B(n12915), .Z(n24284) );
  NANDN U8490 ( .A(x[2171]), .B(y[2171]), .Z(n19078) );
  ANDN U8491 ( .B(y[2172]), .A(x[2172]), .Z(n19084) );
  ANDN U8492 ( .B(n19078), .A(n19084), .Z(n27521) );
  ANDN U8493 ( .B(x[2166]), .A(y[2166]), .Z(n19066) );
  NANDN U8494 ( .A(y[2167]), .B(x[2167]), .Z(n12920) );
  NANDN U8495 ( .A(n19066), .B(n12920), .Z(n27517) );
  NANDN U8496 ( .A(x[2163]), .B(y[2163]), .Z(n27512) );
  ANDN U8497 ( .B(y[2164]), .A(x[2164]), .Z(n12922) );
  ANDN U8498 ( .B(n27512), .A(n12922), .Z(n8676) );
  NANDN U8499 ( .A(x[2162]), .B(y[2162]), .Z(n12924) );
  NANDN U8500 ( .A(x[2161]), .B(y[2161]), .Z(n4240) );
  AND U8501 ( .A(n12924), .B(n4240), .Z(n8670) );
  NANDN U8502 ( .A(x[2160]), .B(y[2160]), .Z(n4241) );
  AND U8503 ( .A(n8670), .B(n4241), .Z(n27510) );
  ANDN U8504 ( .B(x[2159]), .A(y[2159]), .Z(n27509) );
  NANDN U8505 ( .A(x[2158]), .B(y[2158]), .Z(n4243) );
  NANDN U8506 ( .A(x[2159]), .B(y[2159]), .Z(n4242) );
  AND U8507 ( .A(n4243), .B(n4242), .Z(n27508) );
  NANDN U8508 ( .A(x[2157]), .B(y[2157]), .Z(n27506) );
  ANDN U8509 ( .B(x[2156]), .A(y[2156]), .Z(n19047) );
  NANDN U8510 ( .A(y[2157]), .B(x[2157]), .Z(n12926) );
  NANDN U8511 ( .A(n19047), .B(n12926), .Z(n27505) );
  NANDN U8512 ( .A(x[2155]), .B(y[2155]), .Z(n19044) );
  NANDN U8513 ( .A(x[2156]), .B(y[2156]), .Z(n12927) );
  AND U8514 ( .A(n19044), .B(n12927), .Z(n27504) );
  ANDN U8515 ( .B(x[2155]), .A(y[2155]), .Z(n27502) );
  NANDN U8516 ( .A(y[2154]), .B(x[2154]), .Z(n12929) );
  NANDN U8517 ( .A(n27502), .B(n12929), .Z(n8661) );
  NANDN U8518 ( .A(x[2154]), .B(y[2154]), .Z(n24288) );
  ANDN U8519 ( .B(y[2153]), .A(x[2153]), .Z(n19041) );
  ANDN U8520 ( .B(n24288), .A(n19041), .Z(n27501) );
  ANDN U8521 ( .B(x[2152]), .A(y[2152]), .Z(n12931) );
  ANDN U8522 ( .B(y[2151]), .A(x[2151]), .Z(n19034) );
  ANDN U8523 ( .B(y[2152]), .A(x[2152]), .Z(n19039) );
  NOR U8524 ( .A(n19034), .B(n19039), .Z(n27499) );
  ANDN U8525 ( .B(x[2151]), .A(y[2151]), .Z(n12930) );
  NANDN U8526 ( .A(y[2150]), .B(x[2150]), .Z(n12932) );
  ANDN U8527 ( .B(y[2149]), .A(x[2149]), .Z(n19029) );
  NANDN U8528 ( .A(y[2148]), .B(x[2148]), .Z(n19026) );
  ANDN U8529 ( .B(y[2147]), .A(x[2147]), .Z(n12934) );
  NANDN U8530 ( .A(y[2147]), .B(x[2147]), .Z(n19027) );
  NANDN U8531 ( .A(x[2145]), .B(y[2145]), .Z(n12939) );
  ANDN U8532 ( .B(y[2146]), .A(x[2146]), .Z(n12935) );
  ANDN U8533 ( .B(n12939), .A(n12935), .Z(n8645) );
  NANDN U8534 ( .A(x[2144]), .B(y[2144]), .Z(n4245) );
  NANDN U8535 ( .A(x[2143]), .B(y[2143]), .Z(n4244) );
  AND U8536 ( .A(n4245), .B(n4244), .Z(n12940) );
  NANDN U8537 ( .A(y[2142]), .B(x[2142]), .Z(n4246) );
  NANDN U8538 ( .A(y[2143]), .B(x[2143]), .Z(n12942) );
  AND U8539 ( .A(n4246), .B(n12942), .Z(n12943) );
  NANDN U8540 ( .A(y[2140]), .B(x[2140]), .Z(n12946) );
  NANDN U8541 ( .A(x[2140]), .B(y[2140]), .Z(n12945) );
  NANDN U8542 ( .A(x[2138]), .B(y[2138]), .Z(n27484) );
  NANDN U8543 ( .A(x[2139]), .B(y[2139]), .Z(n27488) );
  NAND U8544 ( .A(n27484), .B(n27488), .Z(n19017) );
  ANDN U8545 ( .B(y[2133]), .A(x[2133]), .Z(n19001) );
  ANDN U8546 ( .B(y[2134]), .A(x[2134]), .Z(n19007) );
  NOR U8547 ( .A(n19001), .B(n19007), .Z(n27480) );
  NANDN U8548 ( .A(y[2132]), .B(x[2132]), .Z(n12952) );
  NANDN U8549 ( .A(y[2133]), .B(x[2133]), .Z(n27479) );
  ANDN U8550 ( .B(y[2132]), .A(x[2132]), .Z(n27478) );
  ANDN U8551 ( .B(x[2131]), .A(y[2131]), .Z(n12951) );
  NANDN U8552 ( .A(y[2130]), .B(x[2130]), .Z(n8634) );
  ANDN U8553 ( .B(y[2129]), .A(x[2129]), .Z(n18995) );
  NANDN U8554 ( .A(x[2131]), .B(y[2131]), .Z(n4248) );
  NANDN U8555 ( .A(x[2130]), .B(y[2130]), .Z(n4247) );
  NAND U8556 ( .A(n4248), .B(n4247), .Z(n18998) );
  ANDN U8557 ( .B(x[2128]), .A(y[2128]), .Z(n12953) );
  NANDN U8558 ( .A(x[2127]), .B(y[2127]), .Z(n12955) );
  ANDN U8559 ( .B(x[2126]), .A(y[2126]), .Z(n12957) );
  NANDN U8560 ( .A(x[2125]), .B(y[2125]), .Z(n18987) );
  NANDN U8561 ( .A(y[2124]), .B(x[2124]), .Z(n27468) );
  NANDN U8562 ( .A(x[2121]), .B(y[2121]), .Z(n12961) );
  ANDN U8563 ( .B(y[2122]), .A(x[2122]), .Z(n27465) );
  ANDN U8564 ( .B(n12961), .A(n27465), .Z(n8621) );
  NANDN U8565 ( .A(y[2121]), .B(x[2121]), .Z(n27464) );
  ANDN U8566 ( .B(y[2118]), .A(x[2118]), .Z(n27460) );
  NANDN U8567 ( .A(y[2117]), .B(x[2117]), .Z(n18971) );
  NANDN U8568 ( .A(y[2116]), .B(x[2116]), .Z(n12963) );
  NANDN U8569 ( .A(x[2117]), .B(y[2117]), .Z(n4250) );
  NANDN U8570 ( .A(x[2116]), .B(y[2116]), .Z(n4249) );
  NAND U8571 ( .A(n4250), .B(n4249), .Z(n27458) );
  NANDN U8572 ( .A(x[2115]), .B(y[2115]), .Z(n12964) );
  NANDN U8573 ( .A(y[2114]), .B(x[2114]), .Z(n27454) );
  NANDN U8574 ( .A(y[2115]), .B(x[2115]), .Z(n27457) );
  NAND U8575 ( .A(n27454), .B(n27457), .Z(n8610) );
  NANDN U8576 ( .A(x[2114]), .B(y[2114]), .Z(n12965) );
  NANDN U8577 ( .A(x[2113]), .B(y[2113]), .Z(n27453) );
  AND U8578 ( .A(n12965), .B(n27453), .Z(n8608) );
  NANDN U8579 ( .A(y[2112]), .B(x[2112]), .Z(n12968) );
  NANDN U8580 ( .A(y[2113]), .B(x[2113]), .Z(n12966) );
  NAND U8581 ( .A(n12968), .B(n12966), .Z(n27451) );
  NANDN U8582 ( .A(x[2112]), .B(y[2112]), .Z(n18962) );
  ANDN U8583 ( .B(y[2111]), .A(x[2111]), .Z(n18957) );
  ANDN U8584 ( .B(n18962), .A(n18957), .Z(n27450) );
  ANDN U8585 ( .B(x[2110]), .A(y[2110]), .Z(n12969) );
  NANDN U8586 ( .A(x[2109]), .B(y[2109]), .Z(n12972) );
  NANDN U8587 ( .A(x[2110]), .B(y[2110]), .Z(n18958) );
  AND U8588 ( .A(n12972), .B(n18958), .Z(n27448) );
  NANDN U8589 ( .A(y[2109]), .B(x[2109]), .Z(n12970) );
  NANDN U8590 ( .A(y[2108]), .B(x[2108]), .Z(n27447) );
  ANDN U8591 ( .B(y[2107]), .A(x[2107]), .Z(n18949) );
  NANDN U8592 ( .A(x[2108]), .B(y[2108]), .Z(n12971) );
  NANDN U8593 ( .A(n18949), .B(n12971), .Z(n27446) );
  NANDN U8594 ( .A(y[2107]), .B(x[2107]), .Z(n27445) );
  NANDN U8595 ( .A(y[2106]), .B(x[2106]), .Z(n12973) );
  AND U8596 ( .A(n27445), .B(n12973), .Z(n8598) );
  NANDN U8597 ( .A(x[2106]), .B(y[2106]), .Z(n27444) );
  NANDN U8598 ( .A(y[2105]), .B(x[2105]), .Z(n12974) );
  ANDN U8599 ( .B(y[2103]), .A(x[2103]), .Z(n12975) );
  ANDN U8600 ( .B(y[2101]), .A(x[2101]), .Z(n12977) );
  NANDN U8601 ( .A(y[2101]), .B(x[2101]), .Z(n12980) );
  NANDN U8602 ( .A(y[2100]), .B(x[2100]), .Z(n4251) );
  AND U8603 ( .A(n12980), .B(n4251), .Z(n18936) );
  ANDN U8604 ( .B(y[2100]), .A(x[2100]), .Z(n12978) );
  NANDN U8605 ( .A(x[2099]), .B(y[2099]), .Z(n12982) );
  ANDN U8606 ( .B(y[2097]), .A(x[2097]), .Z(n24297) );
  NANDN U8607 ( .A(y[2096]), .B(x[2096]), .Z(n18926) );
  NANDN U8608 ( .A(y[2097]), .B(x[2097]), .Z(n12983) );
  AND U8609 ( .A(n18926), .B(n12983), .Z(n27435) );
  ANDN U8610 ( .B(y[2095]), .A(x[2095]), .Z(n18923) );
  ANDN U8611 ( .B(y[2096]), .A(x[2096]), .Z(n18929) );
  OR U8612 ( .A(n18923), .B(n18929), .Z(n27434) );
  NANDN U8613 ( .A(y[2094]), .B(x[2094]), .Z(n18919) );
  NANDN U8614 ( .A(y[2095]), .B(x[2095]), .Z(n18927) );
  AND U8615 ( .A(n18919), .B(n18927), .Z(n24298) );
  ANDN U8616 ( .B(y[2094]), .A(x[2094]), .Z(n24299) );
  NANDN U8617 ( .A(x[2092]), .B(y[2092]), .Z(n12985) );
  NANDN U8618 ( .A(x[2091]), .B(y[2091]), .Z(n27430) );
  AND U8619 ( .A(n12985), .B(n27430), .Z(n8572) );
  ANDN U8620 ( .B(x[2090]), .A(y[2090]), .Z(n12989) );
  NANDN U8621 ( .A(x[2090]), .B(y[2090]), .Z(n12988) );
  ANDN U8622 ( .B(y[2089]), .A(x[2089]), .Z(n18912) );
  ANDN U8623 ( .B(n12988), .A(n18912), .Z(n27428) );
  ANDN U8624 ( .B(x[2089]), .A(y[2089]), .Z(n12990) );
  ANDN U8625 ( .B(x[2074]), .A(y[2074]), .Z(n13002) );
  ANDN U8626 ( .B(x[2075]), .A(y[2075]), .Z(n18892) );
  OR U8627 ( .A(n13002), .B(n18892), .Z(n27414) );
  NANDN U8628 ( .A(x[2074]), .B(y[2074]), .Z(n18888) );
  ANDN U8629 ( .B(y[2073]), .A(x[2073]), .Z(n18884) );
  ANDN U8630 ( .B(n18888), .A(n18884), .Z(n27413) );
  ANDN U8631 ( .B(x[2073]), .A(y[2073]), .Z(n13001) );
  NANDN U8632 ( .A(y[2072]), .B(x[2072]), .Z(n13003) );
  NANDN U8633 ( .A(n13001), .B(n13003), .Z(n27412) );
  NANDN U8634 ( .A(x[2071]), .B(y[2071]), .Z(n18878) );
  ANDN U8635 ( .B(y[2072]), .A(x[2072]), .Z(n27411) );
  ANDN U8636 ( .B(n18878), .A(n27411), .Z(n8531) );
  ANDN U8637 ( .B(x[2070]), .A(y[2070]), .Z(n8529) );
  ANDN U8638 ( .B(y[2069]), .A(x[2069]), .Z(n27408) );
  NANDN U8639 ( .A(y[2069]), .B(x[2069]), .Z(n13005) );
  ANDN U8640 ( .B(y[2067]), .A(x[2067]), .Z(n18871) );
  ANDN U8641 ( .B(y[2068]), .A(x[2068]), .Z(n18876) );
  OR U8642 ( .A(n18871), .B(n18876), .Z(n24305) );
  NANDN U8643 ( .A(y[2067]), .B(x[2067]), .Z(n13006) );
  NANDN U8644 ( .A(y[2066]), .B(x[2066]), .Z(n4252) );
  AND U8645 ( .A(n13006), .B(n4252), .Z(n8521) );
  NANDN U8646 ( .A(x[2065]), .B(y[2065]), .Z(n27401) );
  ANDN U8647 ( .B(x[2062]), .A(y[2062]), .Z(n13012) );
  NANDN U8648 ( .A(x[2061]), .B(y[2061]), .Z(n18860) );
  ANDN U8649 ( .B(x[2060]), .A(y[2060]), .Z(n13014) );
  NANDN U8650 ( .A(x[2059]), .B(y[2059]), .Z(n13016) );
  NANDN U8651 ( .A(y[2058]), .B(x[2058]), .Z(n27394) );
  NANDN U8652 ( .A(x[2057]), .B(y[2057]), .Z(n24309) );
  NANDN U8653 ( .A(y[2056]), .B(x[2056]), .Z(n13020) );
  NANDN U8654 ( .A(y[2057]), .B(x[2057]), .Z(n13018) );
  NAND U8655 ( .A(n13020), .B(n13018), .Z(n24308) );
  NANDN U8656 ( .A(x[2055]), .B(y[2055]), .Z(n18850) );
  NANDN U8657 ( .A(y[2054]), .B(x[2054]), .Z(n27391) );
  NANDN U8658 ( .A(x[2051]), .B(y[2051]), .Z(n18839) );
  NANDN U8659 ( .A(x[2052]), .B(y[2052]), .Z(n18846) );
  AND U8660 ( .A(n18839), .B(n18846), .Z(n27388) );
  ANDN U8661 ( .B(x[2051]), .A(y[2051]), .Z(n18844) );
  NANDN U8662 ( .A(y[2050]), .B(x[2050]), .Z(n13022) );
  NANDN U8663 ( .A(n18844), .B(n13022), .Z(n27386) );
  NANDN U8664 ( .A(x[2050]), .B(y[2050]), .Z(n27385) );
  NANDN U8665 ( .A(y[2049]), .B(x[2049]), .Z(n27384) );
  NANDN U8666 ( .A(y[2048]), .B(x[2048]), .Z(n27382) );
  AND U8667 ( .A(n27384), .B(n27382), .Z(n8490) );
  ANDN U8668 ( .B(y[2047]), .A(x[2047]), .Z(n27381) );
  NANDN U8669 ( .A(y[2046]), .B(x[2046]), .Z(n13025) );
  NANDN U8670 ( .A(y[2047]), .B(x[2047]), .Z(n18833) );
  AND U8671 ( .A(n13025), .B(n18833), .Z(n27380) );
  XOR U8672 ( .A(x[2044]), .B(y[2044]), .Z(n13026) );
  NANDN U8673 ( .A(x[2039]), .B(y[2039]), .Z(n27369) );
  XNOR U8674 ( .A(x[2040]), .B(y[2040]), .Z(n13031) );
  AND U8675 ( .A(n27369), .B(n13031), .Z(n8473) );
  NANDN U8676 ( .A(y[2038]), .B(x[2038]), .Z(n27368) );
  NANDN U8677 ( .A(x[2038]), .B(y[2038]), .Z(n13032) );
  ANDN U8678 ( .B(y[2037]), .A(x[2037]), .Z(n18807) );
  ANDN U8679 ( .B(n13032), .A(n18807), .Z(n27367) );
  ANDN U8680 ( .B(y[2035]), .A(x[2035]), .Z(n18802) );
  ANDN U8681 ( .B(y[2036]), .A(x[2036]), .Z(n18810) );
  NOR U8682 ( .A(n18802), .B(n18810), .Z(n27366) );
  NANDN U8683 ( .A(x[2029]), .B(y[2029]), .Z(n4253) );
  ANDN U8684 ( .B(y[2030]), .A(x[2030]), .Z(n13037) );
  ANDN U8685 ( .B(n4253), .A(n13037), .Z(n27359) );
  NANDN U8686 ( .A(y[2028]), .B(x[2028]), .Z(n13041) );
  NANDN U8687 ( .A(y[2029]), .B(x[2029]), .Z(n13036) );
  NAND U8688 ( .A(n13041), .B(n13036), .Z(n27358) );
  NANDN U8689 ( .A(x[2027]), .B(y[2027]), .Z(n13044) );
  NANDN U8690 ( .A(x[2028]), .B(y[2028]), .Z(n13040) );
  NAND U8691 ( .A(n13044), .B(n13040), .Z(n27357) );
  NANDN U8692 ( .A(y[2027]), .B(x[2027]), .Z(n13042) );
  ANDN U8693 ( .B(x[2026]), .A(y[2026]), .Z(n18784) );
  ANDN U8694 ( .B(n13042), .A(n18784), .Z(n27356) );
  ANDN U8695 ( .B(x[2024]), .A(y[2024]), .Z(n18778) );
  ANDN U8696 ( .B(x[2025]), .A(y[2025]), .Z(n18785) );
  NOR U8697 ( .A(n18778), .B(n18785), .Z(n27355) );
  NANDN U8698 ( .A(x[2023]), .B(y[2023]), .Z(n18775) );
  NANDN U8699 ( .A(x[2024]), .B(y[2024]), .Z(n13046) );
  NAND U8700 ( .A(n18775), .B(n13046), .Z(n27354) );
  XOR U8701 ( .A(x[2022]), .B(y[2022]), .Z(n13047) );
  NANDN U8702 ( .A(x[2019]), .B(y[2019]), .Z(n13053) );
  NANDN U8703 ( .A(x[2020]), .B(y[2020]), .Z(n13050) );
  NAND U8704 ( .A(n13053), .B(n13050), .Z(n27350) );
  NANDN U8705 ( .A(y[2018]), .B(x[2018]), .Z(n13054) );
  ANDN U8706 ( .B(y[2017]), .A(x[2017]), .Z(n13056) );
  NANDN U8707 ( .A(y[2016]), .B(x[2016]), .Z(n13058) );
  ANDN U8708 ( .B(y[2015]), .A(x[2015]), .Z(n13060) );
  NANDN U8709 ( .A(y[2015]), .B(x[2015]), .Z(n13059) );
  NANDN U8710 ( .A(x[2014]), .B(y[2014]), .Z(n13061) );
  NANDN U8711 ( .A(x[2013]), .B(y[2013]), .Z(n27339) );
  NAND U8712 ( .A(n13061), .B(n27339), .Z(n8428) );
  NANDN U8713 ( .A(y[2012]), .B(x[2012]), .Z(n4255) );
  NANDN U8714 ( .A(y[2013]), .B(x[2013]), .Z(n4254) );
  AND U8715 ( .A(n4255), .B(n4254), .Z(n13062) );
  NANDN U8716 ( .A(y[2010]), .B(x[2010]), .Z(n4256) );
  ANDN U8717 ( .B(x[2011]), .A(y[2011]), .Z(n18757) );
  ANDN U8718 ( .B(n4256), .A(n18757), .Z(n27336) );
  NANDN U8719 ( .A(y[2008]), .B(x[2008]), .Z(n4258) );
  NANDN U8720 ( .A(y[2009]), .B(x[2009]), .Z(n4257) );
  AND U8721 ( .A(n4258), .B(n4257), .Z(n27334) );
  ANDN U8722 ( .B(y[2004]), .A(x[2004]), .Z(n13064) );
  NANDN U8723 ( .A(x[2001]), .B(y[2001]), .Z(n18740) );
  ANDN U8724 ( .B(y[2002]), .A(x[2002]), .Z(n18746) );
  ANDN U8725 ( .B(n18740), .A(n18746), .Z(n27329) );
  NANDN U8726 ( .A(x[1999]), .B(y[1999]), .Z(n13069) );
  ANDN U8727 ( .B(y[2000]), .A(x[2000]), .Z(n27325) );
  ANDN U8728 ( .B(n13069), .A(n27325), .Z(n24319) );
  ANDN U8729 ( .B(x[1999]), .A(y[1999]), .Z(n27324) );
  NANDN U8730 ( .A(x[1997]), .B(y[1997]), .Z(n13071) );
  NANDN U8731 ( .A(x[1998]), .B(y[1998]), .Z(n13068) );
  NAND U8732 ( .A(n13071), .B(n13068), .Z(n24317) );
  ANDN U8733 ( .B(x[1997]), .A(y[1997]), .Z(n13070) );
  NANDN U8734 ( .A(y[1996]), .B(x[1996]), .Z(n13073) );
  NANDN U8735 ( .A(x[1996]), .B(y[1996]), .Z(n27322) );
  NANDN U8736 ( .A(x[1995]), .B(y[1995]), .Z(n13075) );
  AND U8737 ( .A(n27322), .B(n13075), .Z(n8396) );
  NANDN U8738 ( .A(y[1994]), .B(x[1994]), .Z(n13076) );
  ANDN U8739 ( .B(y[1993]), .A(x[1993]), .Z(n13078) );
  NANDN U8740 ( .A(y[1990]), .B(x[1990]), .Z(n13081) );
  ANDN U8741 ( .B(x[1991]), .A(y[1991]), .Z(n18724) );
  ANDN U8742 ( .B(n13081), .A(n18724), .Z(n27315) );
  ANDN U8743 ( .B(y[1990]), .A(x[1990]), .Z(n18719) );
  NANDN U8744 ( .A(x[1989]), .B(y[1989]), .Z(n13082) );
  NANDN U8745 ( .A(y[1989]), .B(x[1989]), .Z(n27313) );
  NANDN U8746 ( .A(x[1988]), .B(y[1988]), .Z(n13083) );
  ANDN U8747 ( .B(x[1986]), .A(y[1986]), .Z(n27309) );
  ANDN U8748 ( .B(y[1983]), .A(x[1983]), .Z(n18703) );
  ANDN U8749 ( .B(y[1984]), .A(x[1984]), .Z(n18710) );
  NOR U8750 ( .A(n18703), .B(n18710), .Z(n27305) );
  ANDN U8751 ( .B(x[1983]), .A(y[1983]), .Z(n18704) );
  NANDN U8752 ( .A(x[1979]), .B(y[1979]), .Z(n13094) );
  NANDN U8753 ( .A(y[1978]), .B(x[1978]), .Z(n27298) );
  NANDN U8754 ( .A(y[1977]), .B(x[1977]), .Z(n18693) );
  ANDN U8755 ( .B(x[1976]), .A(y[1976]), .Z(n18689) );
  ANDN U8756 ( .B(n18693), .A(n18689), .Z(n27296) );
  NANDN U8757 ( .A(y[1968]), .B(x[1968]), .Z(n4259) );
  NANDN U8758 ( .A(y[1969]), .B(x[1969]), .Z(n13097) );
  AND U8759 ( .A(n4259), .B(n13097), .Z(n27289) );
  ANDN U8760 ( .B(y[1967]), .A(x[1967]), .Z(n18677) );
  NANDN U8761 ( .A(y[1966]), .B(x[1966]), .Z(n4260) );
  NANDN U8762 ( .A(y[1967]), .B(x[1967]), .Z(n18675) );
  AND U8763 ( .A(n4260), .B(n18675), .Z(n27287) );
  ANDN U8764 ( .B(y[1965]), .A(x[1965]), .Z(n27286) );
  ANDN U8765 ( .B(x[1964]), .A(y[1964]), .Z(n18668) );
  NANDN U8766 ( .A(y[1965]), .B(x[1965]), .Z(n13100) );
  NANDN U8767 ( .A(n18668), .B(n13100), .Z(n27285) );
  NANDN U8768 ( .A(x[1963]), .B(y[1963]), .Z(n18664) );
  NANDN U8769 ( .A(x[1964]), .B(y[1964]), .Z(n18671) );
  AND U8770 ( .A(n18664), .B(n18671), .Z(n27284) );
  ANDN U8771 ( .B(x[1963]), .A(y[1963]), .Z(n27283) );
  NANDN U8772 ( .A(x[1962]), .B(y[1962]), .Z(n27282) );
  NANDN U8773 ( .A(y[1961]), .B(x[1961]), .Z(n4262) );
  NANDN U8774 ( .A(y[1962]), .B(x[1962]), .Z(n4261) );
  NAND U8775 ( .A(n4262), .B(n4261), .Z(n27281) );
  NANDN U8776 ( .A(x[1961]), .B(y[1961]), .Z(n4264) );
  NANDN U8777 ( .A(x[1960]), .B(y[1960]), .Z(n4263) );
  AND U8778 ( .A(n4264), .B(n4263), .Z(n27280) );
  NANDN U8779 ( .A(y[1960]), .B(x[1960]), .Z(n4266) );
  NANDN U8780 ( .A(y[1959]), .B(x[1959]), .Z(n4265) );
  AND U8781 ( .A(n4266), .B(n4265), .Z(n24323) );
  NANDN U8782 ( .A(x[1958]), .B(y[1958]), .Z(n4268) );
  NANDN U8783 ( .A(x[1959]), .B(y[1959]), .Z(n4267) );
  NAND U8784 ( .A(n4268), .B(n4267), .Z(n24324) );
  NANDN U8785 ( .A(y[1958]), .B(x[1958]), .Z(n4270) );
  NANDN U8786 ( .A(y[1957]), .B(x[1957]), .Z(n4269) );
  AND U8787 ( .A(n4270), .B(n4269), .Z(n24325) );
  ANDN U8788 ( .B(y[1953]), .A(x[1953]), .Z(n18654) );
  ANDN U8789 ( .B(y[1954]), .A(x[1954]), .Z(n13102) );
  OR U8790 ( .A(n18654), .B(n13102), .Z(n27276) );
  NANDN U8791 ( .A(y[1953]), .B(x[1953]), .Z(n27275) );
  ANDN U8792 ( .B(y[1952]), .A(x[1952]), .Z(n27274) );
  NANDN U8793 ( .A(y[1951]), .B(x[1951]), .Z(n4272) );
  NANDN U8794 ( .A(y[1952]), .B(x[1952]), .Z(n4271) );
  AND U8795 ( .A(n4272), .B(n4271), .Z(n24327) );
  NANDN U8796 ( .A(y[1950]), .B(x[1950]), .Z(n4274) );
  NANDN U8797 ( .A(y[1949]), .B(x[1949]), .Z(n4273) );
  AND U8798 ( .A(n4274), .B(n4273), .Z(n27272) );
  NANDN U8799 ( .A(x[1948]), .B(y[1948]), .Z(n4276) );
  NANDN U8800 ( .A(x[1949]), .B(y[1949]), .Z(n4275) );
  NAND U8801 ( .A(n4276), .B(n4275), .Z(n27271) );
  NANDN U8802 ( .A(y[1948]), .B(x[1948]), .Z(n4278) );
  NANDN U8803 ( .A(y[1947]), .B(x[1947]), .Z(n4277) );
  AND U8804 ( .A(n4278), .B(n4277), .Z(n27270) );
  ANDN U8805 ( .B(x[1946]), .A(y[1946]), .Z(n8304) );
  NANDN U8806 ( .A(y[1944]), .B(x[1944]), .Z(n4279) );
  AND U8807 ( .A(n13110), .B(n4279), .Z(n27268) );
  ANDN U8808 ( .B(y[1944]), .A(x[1944]), .Z(n13109) );
  ANDN U8809 ( .B(y[1943]), .A(x[1943]), .Z(n27267) );
  NOR U8810 ( .A(n13109), .B(n27267), .Z(n8302) );
  ANDN U8811 ( .B(y[1941]), .A(x[1941]), .Z(n18634) );
  ANDN U8812 ( .B(y[1942]), .A(x[1942]), .Z(n18640) );
  NOR U8813 ( .A(n18634), .B(n18640), .Z(n27264) );
  NANDN U8814 ( .A(y[1940]), .B(x[1940]), .Z(n13112) );
  NANDN U8815 ( .A(y[1941]), .B(x[1941]), .Z(n27263) );
  NAND U8816 ( .A(n13112), .B(n27263), .Z(n8298) );
  NANDN U8817 ( .A(x[1939]), .B(y[1939]), .Z(n13113) );
  NANDN U8818 ( .A(x[1940]), .B(y[1940]), .Z(n18635) );
  AND U8819 ( .A(n13113), .B(n18635), .Z(n8296) );
  ANDN U8820 ( .B(x[1938]), .A(y[1938]), .Z(n13115) );
  NANDN U8821 ( .A(y[1936]), .B(x[1936]), .Z(n13120) );
  ANDN U8822 ( .B(x[1934]), .A(y[1934]), .Z(n13123) );
  ANDN U8823 ( .B(x[1932]), .A(y[1932]), .Z(n18618) );
  NANDN U8824 ( .A(x[1931]), .B(y[1931]), .Z(n13125) );
  ANDN U8825 ( .B(y[1932]), .A(x[1932]), .Z(n18623) );
  ANDN U8826 ( .B(n13125), .A(n18623), .Z(n27252) );
  NANDN U8827 ( .A(y[1930]), .B(x[1930]), .Z(n13127) );
  NANDN U8828 ( .A(y[1931]), .B(x[1931]), .Z(n18619) );
  NAND U8829 ( .A(n13127), .B(n18619), .Z(n24328) );
  NANDN U8830 ( .A(x[1929]), .B(y[1929]), .Z(n13129) );
  NANDN U8831 ( .A(x[1930]), .B(y[1930]), .Z(n13126) );
  AND U8832 ( .A(n13129), .B(n13126), .Z(n27251) );
  NANDN U8833 ( .A(x[1927]), .B(y[1927]), .Z(n13132) );
  NANDN U8834 ( .A(x[1928]), .B(y[1928]), .Z(n24329) );
  AND U8835 ( .A(n13132), .B(n24329), .Z(n8276) );
  ANDN U8836 ( .B(x[1926]), .A(y[1926]), .Z(n13133) );
  NANDN U8837 ( .A(y[1927]), .B(x[1927]), .Z(n27248) );
  NANDN U8838 ( .A(y[1924]), .B(x[1924]), .Z(n18604) );
  ANDN U8839 ( .B(x[1920]), .A(y[1920]), .Z(n13140) );
  ANDN U8840 ( .B(x[1921]), .A(y[1921]), .Z(n18600) );
  NOR U8841 ( .A(n13140), .B(n18600), .Z(n27240) );
  ANDN U8842 ( .B(y[1919]), .A(x[1919]), .Z(n18591) );
  NANDN U8843 ( .A(x[1920]), .B(y[1920]), .Z(n18596) );
  NANDN U8844 ( .A(n18591), .B(n18596), .Z(n24330) );
  ANDN U8845 ( .B(y[1917]), .A(x[1917]), .Z(n18586) );
  ANDN U8846 ( .B(y[1916]), .A(x[1916]), .Z(n18587) );
  NANDN U8847 ( .A(y[1916]), .B(x[1916]), .Z(n4281) );
  NANDN U8848 ( .A(y[1915]), .B(x[1915]), .Z(n4280) );
  AND U8849 ( .A(n4281), .B(n4280), .Z(n27235) );
  NANDN U8850 ( .A(y[1914]), .B(x[1914]), .Z(n13146) );
  NANDN U8851 ( .A(x[1914]), .B(y[1914]), .Z(n13144) );
  NANDN U8852 ( .A(x[1913]), .B(y[1913]), .Z(n18581) );
  AND U8853 ( .A(n13144), .B(n18581), .Z(n8251) );
  ANDN U8854 ( .B(x[1913]), .A(y[1913]), .Z(n13145) );
  NANDN U8855 ( .A(y[1912]), .B(x[1912]), .Z(n18577) );
  ANDN U8856 ( .B(y[1911]), .A(x[1911]), .Z(n27229) );
  NANDN U8857 ( .A(y[1910]), .B(x[1910]), .Z(n13147) );
  NANDN U8858 ( .A(y[1911]), .B(x[1911]), .Z(n18578) );
  NANDN U8859 ( .A(x[1909]), .B(y[1909]), .Z(n18568) );
  NANDN U8860 ( .A(x[1910]), .B(y[1910]), .Z(n18575) );
  NAND U8861 ( .A(n18568), .B(n18575), .Z(n27227) );
  ANDN U8862 ( .B(x[1908]), .A(y[1908]), .Z(n13149) );
  ANDN U8863 ( .B(x[1909]), .A(y[1909]), .Z(n18573) );
  OR U8864 ( .A(n13149), .B(n18573), .Z(n27226) );
  NANDN U8865 ( .A(x[1908]), .B(y[1908]), .Z(n18567) );
  ANDN U8866 ( .B(y[1907]), .A(x[1907]), .Z(n18562) );
  ANDN U8867 ( .B(n18567), .A(n18562), .Z(n27225) );
  NANDN U8868 ( .A(x[1905]), .B(y[1905]), .Z(n13152) );
  NANDN U8869 ( .A(x[1906]), .B(y[1906]), .Z(n18563) );
  AND U8870 ( .A(n13152), .B(n18563), .Z(n8239) );
  ANDN U8871 ( .B(x[1905]), .A(y[1905]), .Z(n13150) );
  NANDN U8872 ( .A(x[1904]), .B(y[1904]), .Z(n13153) );
  NANDN U8873 ( .A(y[1902]), .B(x[1902]), .Z(n24336) );
  NANDN U8874 ( .A(y[1903]), .B(x[1903]), .Z(n24334) );
  NAND U8875 ( .A(n24336), .B(n24334), .Z(n13154) );
  NANDN U8876 ( .A(x[1902]), .B(y[1902]), .Z(n18550) );
  NANDN U8877 ( .A(x[1901]), .B(y[1901]), .Z(n18551) );
  AND U8878 ( .A(n18550), .B(n18551), .Z(n8232) );
  NANDN U8879 ( .A(x[1900]), .B(y[1900]), .Z(n18552) );
  ANDN U8880 ( .B(y[1899]), .A(x[1899]), .Z(n27217) );
  ANDN U8881 ( .B(n18552), .A(n27217), .Z(n8229) );
  ANDN U8882 ( .B(x[1898]), .A(y[1898]), .Z(n18543) );
  NANDN U8883 ( .A(y[1899]), .B(x[1899]), .Z(n13158) );
  NANDN U8884 ( .A(n18543), .B(n13158), .Z(n27216) );
  NANDN U8885 ( .A(x[1898]), .B(y[1898]), .Z(n27215) );
  NANDN U8886 ( .A(y[1894]), .B(x[1894]), .Z(n13165) );
  NANDN U8887 ( .A(x[1893]), .B(y[1893]), .Z(n13167) );
  NANDN U8888 ( .A(y[1893]), .B(x[1893]), .Z(n13166) );
  NANDN U8889 ( .A(y[1892]), .B(x[1892]), .Z(n18534) );
  NAND U8890 ( .A(n13166), .B(n18534), .Z(n8216) );
  NANDN U8891 ( .A(x[1891]), .B(y[1891]), .Z(n13170) );
  NANDN U8892 ( .A(y[1890]), .B(x[1890]), .Z(n13171) );
  NANDN U8893 ( .A(x[1889]), .B(y[1889]), .Z(n27205) );
  NANDN U8894 ( .A(y[1888]), .B(x[1888]), .Z(n27204) );
  NANDN U8895 ( .A(y[1886]), .B(x[1886]), .Z(n13174) );
  NANDN U8896 ( .A(y[1887]), .B(x[1887]), .Z(n13173) );
  AND U8897 ( .A(n13174), .B(n13173), .Z(n27202) );
  NANDN U8898 ( .A(x[1886]), .B(y[1886]), .Z(n27201) );
  NANDN U8899 ( .A(y[1885]), .B(x[1885]), .Z(n13175) );
  NANDN U8900 ( .A(y[1884]), .B(x[1884]), .Z(n18519) );
  NANDN U8901 ( .A(x[1885]), .B(y[1885]), .Z(n4282) );
  NANDN U8902 ( .A(x[1884]), .B(y[1884]), .Z(n4283) );
  AND U8903 ( .A(n4283), .B(n4282), .Z(n27199) );
  NANDN U8904 ( .A(x[1883]), .B(y[1883]), .Z(n13176) );
  ANDN U8905 ( .B(x[1882]), .A(y[1882]), .Z(n13178) );
  NANDN U8906 ( .A(x[1881]), .B(y[1881]), .Z(n13181) );
  NANDN U8907 ( .A(y[1880]), .B(x[1880]), .Z(n13182) );
  ANDN U8908 ( .B(y[1879]), .A(x[1879]), .Z(n18511) );
  ANDN U8909 ( .B(y[1877]), .A(x[1877]), .Z(n13185) );
  NANDN U8910 ( .A(y[1877]), .B(x[1877]), .Z(n13184) );
  ANDN U8911 ( .B(x[1876]), .A(y[1876]), .Z(n18504) );
  ANDN U8912 ( .B(n13184), .A(n18504), .Z(n27190) );
  NANDN U8913 ( .A(x[1871]), .B(y[1871]), .Z(n13194) );
  NANDN U8914 ( .A(y[1871]), .B(x[1871]), .Z(n13192) );
  NANDN U8915 ( .A(y[1870]), .B(x[1870]), .Z(n13196) );
  AND U8916 ( .A(n13192), .B(n13196), .Z(n8196) );
  ANDN U8917 ( .B(y[1870]), .A(x[1870]), .Z(n13193) );
  NANDN U8918 ( .A(x[1869]), .B(y[1869]), .Z(n13198) );
  NANDN U8919 ( .A(y[1869]), .B(x[1869]), .Z(n13195) );
  ANDN U8920 ( .B(x[1868]), .A(y[1868]), .Z(n13199) );
  ANDN U8921 ( .B(n13195), .A(n13199), .Z(n8192) );
  ANDN U8922 ( .B(y[1867]), .A(x[1867]), .Z(n27178) );
  NANDN U8923 ( .A(y[1867]), .B(x[1867]), .Z(n13200) );
  ANDN U8924 ( .B(y[1865]), .A(x[1865]), .Z(n18482) );
  ANDN U8925 ( .B(y[1866]), .A(x[1866]), .Z(n18490) );
  OR U8926 ( .A(n18482), .B(n18490), .Z(n27176) );
  NANDN U8927 ( .A(y[1864]), .B(x[1864]), .Z(n18479) );
  NANDN U8928 ( .A(y[1865]), .B(x[1865]), .Z(n18486) );
  AND U8929 ( .A(n18479), .B(n18486), .Z(n27175) );
  ANDN U8930 ( .B(y[1863]), .A(x[1863]), .Z(n18476) );
  ANDN U8931 ( .B(y[1864]), .A(x[1864]), .Z(n18485) );
  OR U8932 ( .A(n18476), .B(n18485), .Z(n27174) );
  NANDN U8933 ( .A(y[1862]), .B(x[1862]), .Z(n18473) );
  NANDN U8934 ( .A(y[1863]), .B(x[1863]), .Z(n18480) );
  AND U8935 ( .A(n18473), .B(n18480), .Z(n27173) );
  ANDN U8936 ( .B(y[1862]), .A(x[1862]), .Z(n27172) );
  NANDN U8937 ( .A(y[1860]), .B(x[1860]), .Z(n13203) );
  NANDN U8938 ( .A(x[1859]), .B(y[1859]), .Z(n13206) );
  NANDN U8939 ( .A(y[1858]), .B(x[1858]), .Z(n13207) );
  NANDN U8940 ( .A(x[1857]), .B(y[1857]), .Z(n13210) );
  NANDN U8941 ( .A(y[1856]), .B(x[1856]), .Z(n27163) );
  NANDN U8942 ( .A(x[1855]), .B(y[1855]), .Z(n27160) );
  NANDN U8943 ( .A(y[1855]), .B(x[1855]), .Z(n13211) );
  ANDN U8944 ( .B(x[1854]), .A(y[1854]), .Z(n18461) );
  ANDN U8945 ( .B(n13211), .A(n18461), .Z(n27159) );
  NANDN U8946 ( .A(x[1853]), .B(y[1853]), .Z(n18457) );
  NANDN U8947 ( .A(x[1854]), .B(y[1854]), .Z(n13212) );
  NAND U8948 ( .A(n18457), .B(n13212), .Z(n27156) );
  NANDN U8949 ( .A(x[1849]), .B(y[1849]), .Z(n13220) );
  NANDN U8950 ( .A(y[1849]), .B(x[1849]), .Z(n13218) );
  NANDN U8951 ( .A(y[1848]), .B(x[1848]), .Z(n18450) );
  AND U8952 ( .A(n13218), .B(n18450), .Z(n8158) );
  NANDN U8953 ( .A(x[1847]), .B(y[1847]), .Z(n13222) );
  NANDN U8954 ( .A(y[1847]), .B(x[1847]), .Z(n18451) );
  NANDN U8955 ( .A(y[1846]), .B(x[1846]), .Z(n13223) );
  AND U8956 ( .A(n18451), .B(n13223), .Z(n8154) );
  ANDN U8957 ( .B(y[1846]), .A(x[1846]), .Z(n13221) );
  NANDN U8958 ( .A(x[1845]), .B(y[1845]), .Z(n27136) );
  ANDN U8959 ( .B(x[1844]), .A(y[1844]), .Z(n27135) );
  NANDN U8960 ( .A(x[1843]), .B(y[1843]), .Z(n13225) );
  NANDN U8961 ( .A(x[1844]), .B(y[1844]), .Z(n18446) );
  AND U8962 ( .A(n13225), .B(n18446), .Z(n27133) );
  ANDN U8963 ( .B(x[1842]), .A(y[1842]), .Z(n18439) );
  ANDN U8964 ( .B(x[1843]), .A(y[1843]), .Z(n18444) );
  OR U8965 ( .A(n18439), .B(n18444), .Z(n27131) );
  NANDN U8966 ( .A(x[1842]), .B(y[1842]), .Z(n27129) );
  NANDN U8967 ( .A(x[1841]), .B(y[1841]), .Z(n4286) );
  NANDN U8968 ( .A(y[1840]), .B(x[1840]), .Z(n4284) );
  ANDN U8969 ( .B(x[1841]), .A(y[1841]), .Z(n18435) );
  ANDN U8970 ( .B(n4284), .A(n18435), .Z(n13226) );
  ANDN U8971 ( .B(n4286), .A(n13226), .Z(n27127) );
  NANDN U8972 ( .A(x[1840]), .B(y[1840]), .Z(n4285) );
  NAND U8973 ( .A(n4286), .B(n4285), .Z(n18434) );
  ANDN U8974 ( .B(y[1837]), .A(x[1837]), .Z(n13231) );
  NANDN U8975 ( .A(y[1836]), .B(x[1836]), .Z(n13234) );
  ANDN U8976 ( .B(x[1834]), .A(y[1834]), .Z(n13237) );
  ANDN U8977 ( .B(x[1832]), .A(y[1832]), .Z(n18421) );
  NANDN U8978 ( .A(y[1833]), .B(x[1833]), .Z(n13238) );
  NANDN U8979 ( .A(n18421), .B(n13238), .Z(n27118) );
  NANDN U8980 ( .A(x[1831]), .B(y[1831]), .Z(n18417) );
  NANDN U8981 ( .A(x[1832]), .B(y[1832]), .Z(n18423) );
  AND U8982 ( .A(n18417), .B(n18423), .Z(n27117) );
  ANDN U8983 ( .B(x[1830]), .A(y[1830]), .Z(n13242) );
  NANDN U8984 ( .A(x[1829]), .B(y[1829]), .Z(n13245) );
  NANDN U8985 ( .A(y[1828]), .B(x[1828]), .Z(n13246) );
  ANDN U8986 ( .B(y[1827]), .A(x[1827]), .Z(n13248) );
  NANDN U8987 ( .A(y[1827]), .B(x[1827]), .Z(n13247) );
  ANDN U8988 ( .B(y[1825]), .A(x[1825]), .Z(n13250) );
  NANDN U8989 ( .A(y[1824]), .B(x[1824]), .Z(n13253) );
  NANDN U8990 ( .A(y[1822]), .B(x[1822]), .Z(n27105) );
  ANDN U8991 ( .B(x[1823]), .A(y[1823]), .Z(n13252) );
  ANDN U8992 ( .B(n27105), .A(n13252), .Z(n8112) );
  NANDN U8993 ( .A(x[1819]), .B(y[1819]), .Z(n4288) );
  NANDN U8994 ( .A(x[1820]), .B(y[1820]), .Z(n4287) );
  NAND U8995 ( .A(n4288), .B(n4287), .Z(n27102) );
  NANDN U8996 ( .A(y[1819]), .B(x[1819]), .Z(n4290) );
  NANDN U8997 ( .A(y[1818]), .B(x[1818]), .Z(n4289) );
  AND U8998 ( .A(n4290), .B(n4289), .Z(n24342) );
  ANDN U8999 ( .B(y[1818]), .A(x[1818]), .Z(n24343) );
  NANDN U9000 ( .A(x[1817]), .B(y[1817]), .Z(n13255) );
  ANDN U9001 ( .B(x[1817]), .A(y[1817]), .Z(n13254) );
  NANDN U9002 ( .A(x[1816]), .B(y[1816]), .Z(n13256) );
  NANDN U9003 ( .A(y[1815]), .B(x[1815]), .Z(n13258) );
  NANDN U9004 ( .A(y[1814]), .B(x[1814]), .Z(n18391) );
  AND U9005 ( .A(n13258), .B(n18391), .Z(n8098) );
  ANDN U9006 ( .B(y[1814]), .A(x[1814]), .Z(n13259) );
  NANDN U9007 ( .A(x[1813]), .B(y[1813]), .Z(n18387) );
  ANDN U9008 ( .B(x[1812]), .A(y[1812]), .Z(n27095) );
  ANDN U9009 ( .B(y[1809]), .A(x[1809]), .Z(n18375) );
  ANDN U9010 ( .B(y[1810]), .A(x[1810]), .Z(n18381) );
  NOR U9011 ( .A(n18375), .B(n18381), .Z(n27092) );
  ANDN U9012 ( .B(x[1809]), .A(y[1809]), .Z(n18376) );
  NANDN U9013 ( .A(y[1807]), .B(x[1807]), .Z(n13262) );
  NANDN U9014 ( .A(y[1806]), .B(x[1806]), .Z(n13265) );
  NAND U9015 ( .A(n13262), .B(n13265), .Z(n8084) );
  ANDN U9016 ( .B(y[1805]), .A(x[1805]), .Z(n18366) );
  NANDN U9017 ( .A(y[1805]), .B(x[1805]), .Z(n13266) );
  NANDN U9018 ( .A(x[1803]), .B(y[1803]), .Z(n13269) );
  ANDN U9019 ( .B(x[1802]), .A(y[1802]), .Z(n27083) );
  NANDN U9020 ( .A(x[1802]), .B(y[1802]), .Z(n13270) );
  NANDN U9021 ( .A(x[1800]), .B(y[1800]), .Z(n4292) );
  NANDN U9022 ( .A(x[1799]), .B(y[1799]), .Z(n4291) );
  AND U9023 ( .A(n4292), .B(n4291), .Z(n27079) );
  NANDN U9024 ( .A(y[1799]), .B(x[1799]), .Z(n24346) );
  NANDN U9025 ( .A(y[1798]), .B(x[1798]), .Z(n27076) );
  NAND U9026 ( .A(n24346), .B(n27076), .Z(n18359) );
  NANDN U9027 ( .A(x[1797]), .B(y[1797]), .Z(n13271) );
  NANDN U9028 ( .A(y[1796]), .B(x[1796]), .Z(n13274) );
  NANDN U9029 ( .A(x[1795]), .B(y[1795]), .Z(n13275) );
  NANDN U9030 ( .A(x[1793]), .B(y[1793]), .Z(n13279) );
  NANDN U9031 ( .A(x[1791]), .B(y[1791]), .Z(n13283) );
  NANDN U9032 ( .A(y[1790]), .B(x[1790]), .Z(n27069) );
  NANDN U9033 ( .A(x[1790]), .B(y[1790]), .Z(n13284) );
  ANDN U9034 ( .B(x[1789]), .A(y[1789]), .Z(n18348) );
  NANDN U9035 ( .A(y[1788]), .B(x[1788]), .Z(n13285) );
  NANDN U9036 ( .A(n18348), .B(n13285), .Z(n27067) );
  NANDN U9037 ( .A(x[1788]), .B(y[1788]), .Z(n27066) );
  NANDN U9038 ( .A(x[1787]), .B(y[1787]), .Z(n13286) );
  AND U9039 ( .A(n27066), .B(n13286), .Z(n8048) );
  NANDN U9040 ( .A(y[1787]), .B(x[1787]), .Z(n27064) );
  NANDN U9041 ( .A(x[1786]), .B(y[1786]), .Z(n13287) );
  NANDN U9042 ( .A(y[1785]), .B(x[1785]), .Z(n13289) );
  NANDN U9043 ( .A(y[1784]), .B(x[1784]), .Z(n13292) );
  AND U9044 ( .A(n13289), .B(n13292), .Z(n8042) );
  ANDN U9045 ( .B(y[1784]), .A(x[1784]), .Z(n13290) );
  NANDN U9046 ( .A(x[1783]), .B(y[1783]), .Z(n18335) );
  NANDN U9047 ( .A(y[1782]), .B(x[1782]), .Z(n18332) );
  NANDN U9048 ( .A(x[1782]), .B(y[1782]), .Z(n18336) );
  NANDN U9049 ( .A(x[1781]), .B(y[1781]), .Z(n18329) );
  NAND U9050 ( .A(n18336), .B(n18329), .Z(n8036) );
  NANDN U9051 ( .A(y[1780]), .B(x[1780]), .Z(n13295) );
  ANDN U9052 ( .B(x[1778]), .A(y[1778]), .Z(n13296) );
  NANDN U9053 ( .A(x[1777]), .B(y[1777]), .Z(n13298) );
  NANDN U9054 ( .A(x[1778]), .B(y[1778]), .Z(n18326) );
  AND U9055 ( .A(n13298), .B(n18326), .Z(n24351) );
  NANDN U9056 ( .A(y[1776]), .B(x[1776]), .Z(n18319) );
  NANDN U9057 ( .A(y[1777]), .B(x[1777]), .Z(n13297) );
  NAND U9058 ( .A(n18319), .B(n13297), .Z(n24352) );
  NANDN U9059 ( .A(x[1775]), .B(y[1775]), .Z(n18317) );
  NANDN U9060 ( .A(x[1776]), .B(y[1776]), .Z(n13299) );
  AND U9061 ( .A(n18317), .B(n13299), .Z(n27054) );
  NANDN U9062 ( .A(x[1773]), .B(y[1773]), .Z(n13302) );
  NANDN U9063 ( .A(x[1774]), .B(y[1774]), .Z(n13300) );
  AND U9064 ( .A(n13302), .B(n13300), .Z(n8023) );
  ANDN U9065 ( .B(x[1773]), .A(y[1773]), .Z(n18310) );
  NANDN U9066 ( .A(y[1772]), .B(x[1772]), .Z(n8020) );
  NANDN U9067 ( .A(x[1771]), .B(y[1771]), .Z(n13306) );
  NANDN U9068 ( .A(y[1771]), .B(x[1771]), .Z(n13304) );
  ANDN U9069 ( .B(y[1769]), .A(x[1769]), .Z(n13309) );
  NANDN U9070 ( .A(y[1768]), .B(x[1768]), .Z(n27045) );
  ANDN U9071 ( .B(y[1767]), .A(x[1767]), .Z(n27044) );
  NANDN U9072 ( .A(y[1766]), .B(x[1766]), .Z(n18298) );
  NANDN U9073 ( .A(y[1767]), .B(x[1767]), .Z(n13311) );
  AND U9074 ( .A(n18298), .B(n13311), .Z(n27043) );
  ANDN U9075 ( .B(y[1765]), .A(x[1765]), .Z(n18295) );
  ANDN U9076 ( .B(y[1766]), .A(x[1766]), .Z(n18300) );
  OR U9077 ( .A(n18295), .B(n18300), .Z(n27042) );
  NANDN U9078 ( .A(y[1765]), .B(x[1765]), .Z(n27041) );
  ANDN U9079 ( .B(y[1763]), .A(x[1763]), .Z(n18290) );
  NANDN U9080 ( .A(y[1762]), .B(x[1762]), .Z(n18287) );
  NANDN U9081 ( .A(y[1760]), .B(x[1760]), .Z(n13316) );
  ANDN U9082 ( .B(y[1759]), .A(x[1759]), .Z(n18282) );
  NANDN U9083 ( .A(y[1759]), .B(x[1759]), .Z(n13317) );
  NANDN U9084 ( .A(x[1758]), .B(y[1758]), .Z(n18283) );
  ANDN U9085 ( .B(y[1757]), .A(x[1757]), .Z(n27032) );
  ANDN U9086 ( .B(n18283), .A(n27032), .Z(n7992) );
  ANDN U9087 ( .B(x[1756]), .A(y[1756]), .Z(n27031) );
  NANDN U9088 ( .A(x[1755]), .B(y[1755]), .Z(n18272) );
  NANDN U9089 ( .A(x[1756]), .B(y[1756]), .Z(n18279) );
  AND U9090 ( .A(n18272), .B(n18279), .Z(n27030) );
  ANDN U9091 ( .B(x[1755]), .A(y[1755]), .Z(n18277) );
  NANDN U9092 ( .A(y[1754]), .B(x[1754]), .Z(n13320) );
  NANDN U9093 ( .A(n18277), .B(n13320), .Z(n27029) );
  NANDN U9094 ( .A(x[1754]), .B(y[1754]), .Z(n27027) );
  NANDN U9095 ( .A(y[1753]), .B(x[1753]), .Z(n27026) );
  NANDN U9096 ( .A(x[1753]), .B(y[1753]), .Z(n27028) );
  NANDN U9097 ( .A(x[1752]), .B(y[1752]), .Z(n27025) );
  AND U9098 ( .A(n27028), .B(n27025), .Z(n18269) );
  NANDN U9099 ( .A(y[1751]), .B(x[1751]), .Z(n4294) );
  NANDN U9100 ( .A(y[1752]), .B(x[1752]), .Z(n4293) );
  NAND U9101 ( .A(n4294), .B(n4293), .Z(n27024) );
  NANDN U9102 ( .A(x[1751]), .B(y[1751]), .Z(n4296) );
  NANDN U9103 ( .A(x[1750]), .B(y[1750]), .Z(n4295) );
  AND U9104 ( .A(n4296), .B(n4295), .Z(n27023) );
  NANDN U9105 ( .A(x[1749]), .B(y[1749]), .Z(n4298) );
  NANDN U9106 ( .A(x[1748]), .B(y[1748]), .Z(n4297) );
  AND U9107 ( .A(n4298), .B(n4297), .Z(n24355) );
  NANDN U9108 ( .A(y[1746]), .B(x[1746]), .Z(n27017) );
  NANDN U9109 ( .A(y[1745]), .B(x[1745]), .Z(n13323) );
  ANDN U9110 ( .B(x[1744]), .A(y[1744]), .Z(n18256) );
  ANDN U9111 ( .B(n13323), .A(n18256), .Z(n27015) );
  NANDN U9112 ( .A(x[1743]), .B(y[1743]), .Z(n18252) );
  NANDN U9113 ( .A(x[1744]), .B(y[1744]), .Z(n13324) );
  NAND U9114 ( .A(n18252), .B(n13324), .Z(n27014) );
  ANDN U9115 ( .B(x[1743]), .A(y[1743]), .Z(n24356) );
  ANDN U9116 ( .B(x[1740]), .A(y[1740]), .Z(n18247) );
  NANDN U9117 ( .A(x[1739]), .B(y[1739]), .Z(n18244) );
  ANDN U9118 ( .B(x[1738]), .A(y[1738]), .Z(n27009) );
  NANDN U9119 ( .A(x[1737]), .B(y[1737]), .Z(n18238) );
  XNOR U9120 ( .A(x[1738]), .B(y[1738]), .Z(n18241) );
  ANDN U9121 ( .B(x[1737]), .A(y[1737]), .Z(n18242) );
  IV U9122 ( .A(n18242), .Z(n27010) );
  ANDN U9123 ( .B(x[1736]), .A(y[1736]), .Z(n13329) );
  ANDN U9124 ( .B(n27010), .A(n13329), .Z(n7956) );
  ANDN U9125 ( .B(y[1735]), .A(x[1735]), .Z(n27005) );
  NANDN U9126 ( .A(y[1735]), .B(x[1735]), .Z(n13330) );
  ANDN U9127 ( .B(y[1734]), .A(x[1734]), .Z(n18234) );
  NANDN U9128 ( .A(x[1733]), .B(y[1733]), .Z(n13331) );
  NANDN U9129 ( .A(n18234), .B(n13331), .Z(n27003) );
  NANDN U9130 ( .A(y[1732]), .B(x[1732]), .Z(n13333) );
  NANDN U9131 ( .A(y[1733]), .B(x[1733]), .Z(n18230) );
  AND U9132 ( .A(n13333), .B(n18230), .Z(n27002) );
  NANDN U9133 ( .A(x[1731]), .B(y[1731]), .Z(n13335) );
  NANDN U9134 ( .A(x[1732]), .B(y[1732]), .Z(n13332) );
  NAND U9135 ( .A(n13335), .B(n13332), .Z(n27001) );
  NANDN U9136 ( .A(y[1730]), .B(x[1730]), .Z(n13337) );
  NANDN U9137 ( .A(y[1731]), .B(x[1731]), .Z(n13334) );
  AND U9138 ( .A(n13337), .B(n13334), .Z(n27000) );
  ANDN U9139 ( .B(y[1729]), .A(x[1729]), .Z(n13338) );
  ANDN U9140 ( .B(x[1729]), .A(y[1729]), .Z(n13336) );
  NANDN U9141 ( .A(y[1727]), .B(x[1727]), .Z(n13341) );
  NANDN U9142 ( .A(y[1726]), .B(x[1726]), .Z(n18216) );
  AND U9143 ( .A(n13341), .B(n18216), .Z(n7940) );
  NANDN U9144 ( .A(x[1725]), .B(y[1725]), .Z(n26994) );
  NANDN U9145 ( .A(y[1725]), .B(x[1725]), .Z(n18217) );
  ANDN U9146 ( .B(y[1723]), .A(x[1723]), .Z(n18208) );
  NANDN U9147 ( .A(x[1724]), .B(y[1724]), .Z(n13344) );
  NANDN U9148 ( .A(n18208), .B(n13344), .Z(n26992) );
  NANDN U9149 ( .A(y[1722]), .B(x[1722]), .Z(n13345) );
  NANDN U9150 ( .A(y[1723]), .B(x[1723]), .Z(n18212) );
  AND U9151 ( .A(n13345), .B(n18212), .Z(n26991) );
  ANDN U9152 ( .B(y[1721]), .A(x[1721]), .Z(n18203) );
  ANDN U9153 ( .B(y[1722]), .A(x[1722]), .Z(n18210) );
  OR U9154 ( .A(n18203), .B(n18210), .Z(n26990) );
  NANDN U9155 ( .A(y[1720]), .B(x[1720]), .Z(n13347) );
  NANDN U9156 ( .A(y[1721]), .B(x[1721]), .Z(n26988) );
  AND U9157 ( .A(n13347), .B(n26988), .Z(n7931) );
  ANDN U9158 ( .B(y[1720]), .A(x[1720]), .Z(n26987) );
  NANDN U9159 ( .A(x[1719]), .B(y[1719]), .Z(n13348) );
  ANDN U9160 ( .B(x[1718]), .A(y[1718]), .Z(n13350) );
  NANDN U9161 ( .A(x[1718]), .B(y[1718]), .Z(n13349) );
  ANDN U9162 ( .B(x[1716]), .A(y[1716]), .Z(n18195) );
  NANDN U9163 ( .A(x[1715]), .B(y[1715]), .Z(n4300) );
  NANDN U9164 ( .A(x[1716]), .B(y[1716]), .Z(n4299) );
  AND U9165 ( .A(n4300), .B(n4299), .Z(n18193) );
  NANDN U9166 ( .A(y[1714]), .B(x[1714]), .Z(n4302) );
  NANDN U9167 ( .A(y[1715]), .B(x[1715]), .Z(n4301) );
  NAND U9168 ( .A(n4302), .B(n4301), .Z(n18191) );
  NANDN U9169 ( .A(x[1714]), .B(y[1714]), .Z(n4304) );
  NANDN U9170 ( .A(x[1713]), .B(y[1713]), .Z(n4303) );
  AND U9171 ( .A(n4304), .B(n4303), .Z(n13352) );
  NANDN U9172 ( .A(y[1711]), .B(x[1711]), .Z(n4308) );
  NANDN U9173 ( .A(x[1710]), .B(y[1710]), .Z(n13355) );
  NANDN U9174 ( .A(x[1709]), .B(y[1709]), .Z(n4305) );
  AND U9175 ( .A(n13355), .B(n4305), .Z(n7910) );
  ANDN U9176 ( .B(x[1708]), .A(y[1708]), .Z(n18178) );
  NANDN U9177 ( .A(y[1709]), .B(x[1709]), .Z(n13354) );
  NANDN U9178 ( .A(n18178), .B(n13354), .Z(n4306) );
  NAND U9179 ( .A(n7910), .B(n4306), .Z(n4307) );
  AND U9180 ( .A(n4308), .B(n4307), .Z(n4309) );
  NANDN U9181 ( .A(y[1710]), .B(x[1710]), .Z(n13353) );
  NAND U9182 ( .A(n4309), .B(n13353), .Z(n24361) );
  NANDN U9183 ( .A(x[1707]), .B(y[1707]), .Z(n13357) );
  NANDN U9184 ( .A(y[1706]), .B(x[1706]), .Z(n13360) );
  NANDN U9185 ( .A(x[1705]), .B(y[1705]), .Z(n13361) );
  ANDN U9186 ( .B(x[1704]), .A(y[1704]), .Z(n13363) );
  NANDN U9187 ( .A(x[1703]), .B(y[1703]), .Z(n13366) );
  ANDN U9188 ( .B(y[1702]), .A(x[1702]), .Z(n13365) );
  NANDN U9189 ( .A(y[1701]), .B(x[1701]), .Z(n13368) );
  NANDN U9190 ( .A(y[1698]), .B(x[1698]), .Z(n13369) );
  NANDN U9191 ( .A(y[1700]), .B(x[1700]), .Z(n7894) );
  NANDN U9192 ( .A(y[1699]), .B(x[1699]), .Z(n4310) );
  AND U9193 ( .A(n7894), .B(n4310), .Z(n26969) );
  AND U9194 ( .A(n13369), .B(n26969), .Z(n7891) );
  NANDN U9195 ( .A(x[1697]), .B(y[1697]), .Z(n18161) );
  NANDN U9196 ( .A(x[1698]), .B(y[1698]), .Z(n26968) );
  NAND U9197 ( .A(n18161), .B(n26968), .Z(n7889) );
  NANDN U9198 ( .A(y[1696]), .B(x[1696]), .Z(n26964) );
  NANDN U9199 ( .A(y[1694]), .B(x[1694]), .Z(n26960) );
  NANDN U9200 ( .A(y[1695]), .B(x[1695]), .Z(n26963) );
  AND U9201 ( .A(n26960), .B(n26963), .Z(n18157) );
  ANDN U9202 ( .B(x[1692]), .A(y[1692]), .Z(n13375) );
  NANDN U9203 ( .A(x[1691]), .B(y[1691]), .Z(n13377) );
  ANDN U9204 ( .B(x[1690]), .A(y[1690]), .Z(n18149) );
  NANDN U9205 ( .A(y[1689]), .B(x[1689]), .Z(n4312) );
  NANDN U9206 ( .A(y[1688]), .B(x[1688]), .Z(n4311) );
  AND U9207 ( .A(n4312), .B(n4311), .Z(n18145) );
  NANDN U9208 ( .A(x[1687]), .B(y[1687]), .Z(n4313) );
  ANDN U9209 ( .B(y[1688]), .A(x[1688]), .Z(n18143) );
  ANDN U9210 ( .B(n4313), .A(n18143), .Z(n4317) );
  ANDN U9211 ( .B(x[1686]), .A(y[1686]), .Z(n18138) );
  NANDN U9212 ( .A(y[1687]), .B(x[1687]), .Z(n18142) );
  NANDN U9213 ( .A(n18138), .B(n18142), .Z(n4314) );
  NAND U9214 ( .A(n4317), .B(n4314), .Z(n4315) );
  NAND U9215 ( .A(n18145), .B(n4315), .Z(n24365) );
  NANDN U9216 ( .A(x[1686]), .B(y[1686]), .Z(n4316) );
  AND U9217 ( .A(n4317), .B(n4316), .Z(n26953) );
  NANDN U9218 ( .A(x[1685]), .B(y[1685]), .Z(n13380) );
  ANDN U9219 ( .B(x[1685]), .A(y[1685]), .Z(n18137) );
  NANDN U9220 ( .A(x[1684]), .B(y[1684]), .Z(n13381) );
  NANDN U9221 ( .A(y[1682]), .B(x[1682]), .Z(n13386) );
  NANDN U9222 ( .A(x[1682]), .B(y[1682]), .Z(n13385) );
  NANDN U9223 ( .A(x[1681]), .B(y[1681]), .Z(n13388) );
  NAND U9224 ( .A(n13385), .B(n13388), .Z(n7864) );
  NANDN U9225 ( .A(y[1681]), .B(x[1681]), .Z(n13387) );
  NANDN U9226 ( .A(y[1680]), .B(x[1680]), .Z(n26946) );
  AND U9227 ( .A(n13387), .B(n26946), .Z(n7862) );
  ANDN U9228 ( .B(y[1679]), .A(x[1679]), .Z(n13392) );
  NANDN U9229 ( .A(y[1678]), .B(x[1678]), .Z(n13394) );
  NANDN U9230 ( .A(y[1679]), .B(x[1679]), .Z(n13390) );
  AND U9231 ( .A(n13394), .B(n13390), .Z(n24366) );
  NANDN U9232 ( .A(y[1677]), .B(x[1677]), .Z(n26942) );
  NANDN U9233 ( .A(x[1677]), .B(y[1677]), .Z(n4319) );
  NANDN U9234 ( .A(x[1676]), .B(y[1676]), .Z(n4318) );
  NAND U9235 ( .A(n4319), .B(n4318), .Z(n26941) );
  NANDN U9236 ( .A(y[1676]), .B(x[1676]), .Z(n4321) );
  NANDN U9237 ( .A(y[1675]), .B(x[1675]), .Z(n4320) );
  AND U9238 ( .A(n4321), .B(n4320), .Z(n26940) );
  NANDN U9239 ( .A(y[1670]), .B(x[1670]), .Z(n13401) );
  ANDN U9240 ( .B(y[1669]), .A(x[1669]), .Z(n13402) );
  NANDN U9241 ( .A(x[1668]), .B(y[1668]), .Z(n13403) );
  ANDN U9242 ( .B(y[1667]), .A(x[1667]), .Z(n18111) );
  ANDN U9243 ( .B(n13403), .A(n18111), .Z(n26932) );
  NANDN U9244 ( .A(x[1665]), .B(y[1665]), .Z(n7830) );
  NANDN U9245 ( .A(x[1664]), .B(y[1664]), .Z(n4322) );
  AND U9246 ( .A(n7830), .B(n4322), .Z(n26927) );
  NANDN U9247 ( .A(x[1663]), .B(y[1663]), .Z(n13405) );
  ANDN U9248 ( .B(y[1661]), .A(x[1661]), .Z(n13408) );
  NANDN U9249 ( .A(y[1660]), .B(x[1660]), .Z(n13410) );
  ANDN U9250 ( .B(y[1659]), .A(x[1659]), .Z(n13412) );
  NANDN U9251 ( .A(y[1658]), .B(x[1658]), .Z(n24368) );
  NANDN U9252 ( .A(y[1659]), .B(x[1659]), .Z(n13411) );
  ANDN U9253 ( .B(y[1658]), .A(x[1658]), .Z(n13413) );
  NANDN U9254 ( .A(x[1655]), .B(y[1655]), .Z(n13415) );
  ANDN U9255 ( .B(y[1656]), .A(x[1656]), .Z(n26918) );
  ANDN U9256 ( .B(n13415), .A(n26918), .Z(n7814) );
  NANDN U9257 ( .A(y[1655]), .B(x[1655]), .Z(n26917) );
  NANDN U9258 ( .A(y[1652]), .B(x[1652]), .Z(n13421) );
  ANDN U9259 ( .B(x[1650]), .A(y[1650]), .Z(n13422) );
  NANDN U9260 ( .A(x[1649]), .B(y[1649]), .Z(n13424) );
  NANDN U9261 ( .A(y[1648]), .B(x[1648]), .Z(n26909) );
  NANDN U9262 ( .A(x[1645]), .B(y[1645]), .Z(n18070) );
  ANDN U9263 ( .B(y[1646]), .A(x[1646]), .Z(n26906) );
  ANDN U9264 ( .B(n18070), .A(n26906), .Z(n7795) );
  NANDN U9265 ( .A(y[1645]), .B(x[1645]), .Z(n26905) );
  NANDN U9266 ( .A(y[1644]), .B(x[1644]), .Z(n18066) );
  NAND U9267 ( .A(n26905), .B(n18066), .Z(n7793) );
  ANDN U9268 ( .B(y[1643]), .A(x[1643]), .Z(n24371) );
  NANDN U9269 ( .A(y[1643]), .B(x[1643]), .Z(n18067) );
  ANDN U9270 ( .B(y[1641]), .A(x[1641]), .Z(n18059) );
  ANDN U9271 ( .B(y[1642]), .A(x[1642]), .Z(n18064) );
  OR U9272 ( .A(n18059), .B(n18064), .Z(n24373) );
  NANDN U9273 ( .A(y[1640]), .B(x[1640]), .Z(n18057) );
  NANDN U9274 ( .A(y[1641]), .B(x[1641]), .Z(n18060) );
  AND U9275 ( .A(n18057), .B(n18060), .Z(n26903) );
  ANDN U9276 ( .B(y[1640]), .A(x[1640]), .Z(n18055) );
  ANDN U9277 ( .B(y[1639]), .A(x[1639]), .Z(n18050) );
  OR U9278 ( .A(n18055), .B(n18050), .Z(n26902) );
  NANDN U9279 ( .A(y[1639]), .B(x[1639]), .Z(n18053) );
  NANDN U9280 ( .A(y[1638]), .B(x[1638]), .Z(n18046) );
  AND U9281 ( .A(n18053), .B(n18046), .Z(n26901) );
  ANDN U9282 ( .B(y[1638]), .A(x[1638]), .Z(n26899) );
  NANDN U9283 ( .A(x[1637]), .B(y[1637]), .Z(n13428) );
  NANDN U9284 ( .A(y[1636]), .B(x[1636]), .Z(n26896) );
  NANDN U9285 ( .A(y[1637]), .B(x[1637]), .Z(n26898) );
  AND U9286 ( .A(n26896), .B(n26898), .Z(n7781) );
  ANDN U9287 ( .B(y[1635]), .A(x[1635]), .Z(n26895) );
  NANDN U9288 ( .A(y[1635]), .B(x[1635]), .Z(n13429) );
  ANDN U9289 ( .B(x[1634]), .A(y[1634]), .Z(n18037) );
  ANDN U9290 ( .B(n13429), .A(n18037), .Z(n26894) );
  NANDN U9291 ( .A(x[1633]), .B(y[1633]), .Z(n18033) );
  NANDN U9292 ( .A(x[1634]), .B(y[1634]), .Z(n18041) );
  NAND U9293 ( .A(n18033), .B(n18041), .Z(n26893) );
  ANDN U9294 ( .B(x[1632]), .A(y[1632]), .Z(n18028) );
  ANDN U9295 ( .B(x[1633]), .A(y[1633]), .Z(n18039) );
  NOR U9296 ( .A(n18028), .B(n18039), .Z(n26892) );
  ANDN U9297 ( .B(x[1630]), .A(y[1630]), .Z(n18024) );
  ANDN U9298 ( .B(x[1631]), .A(y[1631]), .Z(n18031) );
  NOR U9299 ( .A(n18024), .B(n18031), .Z(n26890) );
  ANDN U9300 ( .B(y[1629]), .A(x[1629]), .Z(n18018) );
  NANDN U9301 ( .A(x[1630]), .B(y[1630]), .Z(n26888) );
  NANDN U9302 ( .A(y[1629]), .B(x[1629]), .Z(n18021) );
  NANDN U9303 ( .A(y[1628]), .B(x[1628]), .Z(n4323) );
  AND U9304 ( .A(n18021), .B(n4323), .Z(n26887) );
  ANDN U9305 ( .B(y[1627]), .A(x[1627]), .Z(n13431) );
  NANDN U9306 ( .A(y[1626]), .B(x[1626]), .Z(n13433) );
  NANDN U9307 ( .A(y[1627]), .B(x[1627]), .Z(n13430) );
  AND U9308 ( .A(n13433), .B(n13430), .Z(n24374) );
  ANDN U9309 ( .B(y[1624]), .A(x[1624]), .Z(n26881) );
  NANDN U9310 ( .A(y[1622]), .B(x[1622]), .Z(n13438) );
  NANDN U9311 ( .A(x[1622]), .B(y[1622]), .Z(n13436) );
  NANDN U9312 ( .A(x[1621]), .B(y[1621]), .Z(n18001) );
  AND U9313 ( .A(n13436), .B(n18001), .Z(n7760) );
  ANDN U9314 ( .B(x[1621]), .A(y[1621]), .Z(n13437) );
  NANDN U9315 ( .A(y[1620]), .B(x[1620]), .Z(n13440) );
  NANDN U9316 ( .A(x[1620]), .B(y[1620]), .Z(n18002) );
  ANDN U9317 ( .B(y[1619]), .A(x[1619]), .Z(n26877) );
  ANDN U9318 ( .B(n18002), .A(n26877), .Z(n7756) );
  ANDN U9319 ( .B(x[1619]), .A(y[1619]), .Z(n13439) );
  ANDN U9320 ( .B(y[1617]), .A(x[1617]), .Z(n17991) );
  ANDN U9321 ( .B(y[1618]), .A(x[1618]), .Z(n17998) );
  OR U9322 ( .A(n17991), .B(n17998), .Z(n24379) );
  NANDN U9323 ( .A(y[1616]), .B(x[1616]), .Z(n17989) );
  NANDN U9324 ( .A(y[1617]), .B(x[1617]), .Z(n17994) );
  AND U9325 ( .A(n17989), .B(n17994), .Z(n24380) );
  ANDN U9326 ( .B(y[1615]), .A(x[1615]), .Z(n13441) );
  ANDN U9327 ( .B(x[1614]), .A(y[1614]), .Z(n26873) );
  NANDN U9328 ( .A(x[1613]), .B(y[1613]), .Z(n26872) );
  NANDN U9329 ( .A(x[1612]), .B(y[1612]), .Z(n26869) );
  ANDN U9330 ( .B(x[1611]), .A(y[1611]), .Z(n26868) );
  NANDN U9331 ( .A(x[1610]), .B(y[1610]), .Z(n4325) );
  NANDN U9332 ( .A(x[1611]), .B(y[1611]), .Z(n4324) );
  AND U9333 ( .A(n4325), .B(n4324), .Z(n26867) );
  ANDN U9334 ( .B(x[1610]), .A(y[1610]), .Z(n26866) );
  ANDN U9335 ( .B(y[1609]), .A(x[1609]), .Z(n26865) );
  NANDN U9336 ( .A(y[1608]), .B(x[1608]), .Z(n17971) );
  ANDN U9337 ( .B(x[1609]), .A(y[1609]), .Z(n13443) );
  ANDN U9338 ( .B(n17971), .A(n13443), .Z(n26864) );
  ANDN U9339 ( .B(y[1608]), .A(x[1608]), .Z(n24381) );
  NANDN U9340 ( .A(y[1606]), .B(x[1606]), .Z(n13446) );
  ANDN U9341 ( .B(y[1606]), .A(x[1606]), .Z(n13445) );
  NANDN U9342 ( .A(x[1605]), .B(y[1605]), .Z(n7729) );
  XNOR U9343 ( .A(x[1605]), .B(y[1605]), .Z(n4327) );
  NANDN U9344 ( .A(y[1604]), .B(x[1604]), .Z(n4326) );
  NAND U9345 ( .A(n4327), .B(n4326), .Z(n4328) );
  NAND U9346 ( .A(n7729), .B(n4328), .Z(n13447) );
  NANDN U9347 ( .A(y[1603]), .B(x[1603]), .Z(n17966) );
  NANDN U9348 ( .A(y[1602]), .B(x[1602]), .Z(n4329) );
  AND U9349 ( .A(n17966), .B(n4329), .Z(n26859) );
  NANDN U9350 ( .A(x[1600]), .B(y[1600]), .Z(n4331) );
  NANDN U9351 ( .A(x[1599]), .B(y[1599]), .Z(n4330) );
  AND U9352 ( .A(n4331), .B(n4330), .Z(n17960) );
  NANDN U9353 ( .A(x[1598]), .B(y[1598]), .Z(n17959) );
  NANDN U9354 ( .A(x[1597]), .B(y[1597]), .Z(n26854) );
  AND U9355 ( .A(n17959), .B(n26854), .Z(n7717) );
  NANDN U9356 ( .A(y[1597]), .B(x[1597]), .Z(n4333) );
  NANDN U9357 ( .A(y[1596]), .B(x[1596]), .Z(n4332) );
  NAND U9358 ( .A(n4333), .B(n4332), .Z(n26852) );
  NANDN U9359 ( .A(x[1596]), .B(y[1596]), .Z(n4335) );
  NANDN U9360 ( .A(x[1595]), .B(y[1595]), .Z(n4334) );
  AND U9361 ( .A(n4335), .B(n4334), .Z(n26851) );
  ANDN U9362 ( .B(x[1595]), .A(y[1595]), .Z(n17953) );
  ANDN U9363 ( .B(x[1594]), .A(y[1594]), .Z(n17949) );
  OR U9364 ( .A(n17953), .B(n17949), .Z(n26850) );
  ANDN U9365 ( .B(y[1593]), .A(x[1593]), .Z(n13450) );
  NANDN U9366 ( .A(y[1593]), .B(x[1593]), .Z(n13449) );
  NANDN U9367 ( .A(x[1592]), .B(y[1592]), .Z(n13451) );
  ANDN U9368 ( .B(y[1591]), .A(x[1591]), .Z(n7705) );
  NANDN U9369 ( .A(y[1590]), .B(x[1590]), .Z(n26844) );
  OR U9370 ( .A(n7705), .B(n26844), .Z(n4338) );
  NANDN U9371 ( .A(y[1592]), .B(x[1592]), .Z(n4337) );
  NANDN U9372 ( .A(y[1591]), .B(x[1591]), .Z(n4336) );
  AND U9373 ( .A(n4337), .B(n4336), .Z(n24382) );
  AND U9374 ( .A(n4338), .B(n24382), .Z(n17944) );
  NANDN U9375 ( .A(y[1588]), .B(x[1588]), .Z(n13454) );
  NANDN U9376 ( .A(y[1587]), .B(x[1587]), .Z(n13455) );
  NANDN U9377 ( .A(x[1586]), .B(y[1586]), .Z(n4340) );
  NANDN U9378 ( .A(x[1587]), .B(y[1587]), .Z(n4339) );
  AND U9379 ( .A(n4340), .B(n4339), .Z(n26842) );
  NANDN U9380 ( .A(y[1586]), .B(x[1586]), .Z(n4342) );
  NANDN U9381 ( .A(y[1585]), .B(x[1585]), .Z(n4341) );
  AND U9382 ( .A(n4342), .B(n4341), .Z(n26841) );
  NANDN U9383 ( .A(x[1584]), .B(y[1584]), .Z(n4344) );
  NANDN U9384 ( .A(x[1585]), .B(y[1585]), .Z(n4343) );
  NAND U9385 ( .A(n4344), .B(n4343), .Z(n26840) );
  NANDN U9386 ( .A(x[1583]), .B(y[1583]), .Z(n7694) );
  XNOR U9387 ( .A(x[1583]), .B(y[1583]), .Z(n4346) );
  NANDN U9388 ( .A(y[1582]), .B(x[1582]), .Z(n4345) );
  NAND U9389 ( .A(n4346), .B(n4345), .Z(n4347) );
  NAND U9390 ( .A(n7694), .B(n4347), .Z(n4349) );
  NANDN U9391 ( .A(y[1584]), .B(x[1584]), .Z(n4348) );
  AND U9392 ( .A(n4349), .B(n4348), .Z(n26839) );
  NANDN U9393 ( .A(y[1581]), .B(x[1581]), .Z(n13458) );
  NANDN U9394 ( .A(y[1580]), .B(x[1580]), .Z(n4350) );
  AND U9395 ( .A(n13458), .B(n4350), .Z(n26835) );
  NANDN U9396 ( .A(x[1581]), .B(y[1581]), .Z(n4352) );
  NANDN U9397 ( .A(n26835), .B(n4352), .Z(n7692) );
  NANDN U9398 ( .A(x[1580]), .B(y[1580]), .Z(n4351) );
  NAND U9399 ( .A(n4352), .B(n4351), .Z(n13457) );
  NANDN U9400 ( .A(y[1579]), .B(x[1579]), .Z(n17933) );
  NANDN U9401 ( .A(y[1578]), .B(x[1578]), .Z(n17929) );
  NANDN U9402 ( .A(x[1579]), .B(y[1579]), .Z(n7686) );
  ANDN U9403 ( .B(y[1577]), .A(x[1577]), .Z(n13459) );
  NANDN U9404 ( .A(y[1577]), .B(x[1577]), .Z(n13462) );
  NANDN U9405 ( .A(y[1576]), .B(x[1576]), .Z(n4353) );
  AND U9406 ( .A(n13462), .B(n4353), .Z(n26832) );
  ANDN U9407 ( .B(y[1576]), .A(x[1576]), .Z(n13460) );
  ANDN U9408 ( .B(y[1573]), .A(x[1573]), .Z(n17915) );
  ANDN U9409 ( .B(y[1574]), .A(x[1574]), .Z(n17922) );
  NOR U9410 ( .A(n17915), .B(n17922), .Z(n26829) );
  NANDN U9411 ( .A(y[1572]), .B(x[1572]), .Z(n17913) );
  NANDN U9412 ( .A(y[1573]), .B(x[1573]), .Z(n17920) );
  NAND U9413 ( .A(n17913), .B(n17920), .Z(n26828) );
  NANDN U9414 ( .A(y[1571]), .B(x[1571]), .Z(n4362) );
  XNOR U9415 ( .A(y[1571]), .B(x[1571]), .Z(n4355) );
  NANDN U9416 ( .A(x[1570]), .B(y[1570]), .Z(n4354) );
  NAND U9417 ( .A(n4355), .B(n4354), .Z(n4356) );
  AND U9418 ( .A(n4362), .B(n4356), .Z(n17911) );
  ANDN U9419 ( .B(y[1572]), .A(x[1572]), .Z(n17917) );
  NOR U9420 ( .A(n17911), .B(n17917), .Z(n26827) );
  NANDN U9421 ( .A(y[1568]), .B(x[1568]), .Z(n4357) );
  NANDN U9422 ( .A(x[1569]), .B(n4357), .Z(n4360) );
  XNOR U9423 ( .A(x[1569]), .B(n4357), .Z(n4358) );
  NAND U9424 ( .A(n4358), .B(y[1569]), .Z(n4359) );
  NAND U9425 ( .A(n4360), .B(n4359), .Z(n4361) );
  AND U9426 ( .A(n4362), .B(n4361), .Z(n4364) );
  NANDN U9427 ( .A(y[1570]), .B(x[1570]), .Z(n4363) );
  AND U9428 ( .A(n4364), .B(n4363), .Z(n24384) );
  NANDN U9429 ( .A(x[1568]), .B(y[1568]), .Z(n4366) );
  NANDN U9430 ( .A(x[1567]), .B(y[1567]), .Z(n4365) );
  AND U9431 ( .A(n4366), .B(n4365), .Z(n4368) );
  NANDN U9432 ( .A(x[1569]), .B(y[1569]), .Z(n4367) );
  NAND U9433 ( .A(n4368), .B(n4367), .Z(n13465) );
  NANDN U9434 ( .A(y[1566]), .B(x[1566]), .Z(n4369) );
  NANDN U9435 ( .A(y[1567]), .B(x[1567]), .Z(n13463) );
  AND U9436 ( .A(n4369), .B(n13463), .Z(n13467) );
  ANDN U9437 ( .B(y[1565]), .A(x[1565]), .Z(n13469) );
  NANDN U9438 ( .A(y[1565]), .B(x[1565]), .Z(n13466) );
  ANDN U9439 ( .B(y[1563]), .A(x[1563]), .Z(n13470) );
  NANDN U9440 ( .A(y[1562]), .B(x[1562]), .Z(n26820) );
  ANDN U9441 ( .B(y[1562]), .A(x[1562]), .Z(n13471) );
  NANDN U9442 ( .A(x[1561]), .B(y[1561]), .Z(n26819) );
  NANDN U9443 ( .A(x[1560]), .B(y[1560]), .Z(n26817) );
  NANDN U9444 ( .A(x[1559]), .B(y[1559]), .Z(n17893) );
  AND U9445 ( .A(n26817), .B(n17893), .Z(n7663) );
  ANDN U9446 ( .B(x[1558]), .A(y[1558]), .Z(n13473) );
  ANDN U9447 ( .B(y[1558]), .A(x[1558]), .Z(n17892) );
  NANDN U9448 ( .A(x[1557]), .B(y[1557]), .Z(n13475) );
  XNOR U9449 ( .A(y[1556]), .B(x[1556]), .Z(n17887) );
  NANDN U9450 ( .A(x[1555]), .B(y[1555]), .Z(n13478) );
  AND U9451 ( .A(n17887), .B(n13478), .Z(n7655) );
  ANDN U9452 ( .B(x[1554]), .A(y[1554]), .Z(n17883) );
  NANDN U9453 ( .A(y[1555]), .B(x[1555]), .Z(n24389) );
  ANDN U9454 ( .B(y[1553]), .A(x[1553]), .Z(n13479) );
  ANDN U9455 ( .B(x[1552]), .A(y[1552]), .Z(n26810) );
  NANDN U9456 ( .A(y[1553]), .B(x[1553]), .Z(n17884) );
  NANDN U9457 ( .A(x[1552]), .B(y[1552]), .Z(n13480) );
  ANDN U9458 ( .B(x[1549]), .A(y[1549]), .Z(n17875) );
  NANDN U9459 ( .A(y[1548]), .B(x[1548]), .Z(n17866) );
  NANDN U9460 ( .A(n17875), .B(n17866), .Z(n26807) );
  ANDN U9461 ( .B(x[1546]), .A(y[1546]), .Z(n26804) );
  NANDN U9462 ( .A(y[1547]), .B(x[1547]), .Z(n26805) );
  NANDN U9463 ( .A(n26804), .B(n26805), .Z(n7640) );
  NANDN U9464 ( .A(x[1546]), .B(y[1546]), .Z(n17864) );
  NANDN U9465 ( .A(x[1545]), .B(y[1545]), .Z(n4371) );
  NANDN U9466 ( .A(y[1544]), .B(x[1544]), .Z(n13482) );
  NANDN U9467 ( .A(y[1545]), .B(x[1545]), .Z(n17861) );
  NAND U9468 ( .A(n13482), .B(n17861), .Z(n7635) );
  AND U9469 ( .A(n4371), .B(n7635), .Z(n26803) );
  NANDN U9470 ( .A(x[1544]), .B(y[1544]), .Z(n4370) );
  AND U9471 ( .A(n4371), .B(n4370), .Z(n17858) );
  NANDN U9472 ( .A(x[1543]), .B(y[1543]), .Z(n13483) );
  NAND U9473 ( .A(n17858), .B(n13483), .Z(n4372) );
  NANDN U9474 ( .A(n26803), .B(n4372), .Z(n4373) );
  AND U9475 ( .A(n17864), .B(n4373), .Z(n7638) );
  ANDN U9476 ( .B(x[1543]), .A(y[1543]), .Z(n13481) );
  NANDN U9477 ( .A(x[1542]), .B(y[1542]), .Z(n13484) );
  ANDN U9478 ( .B(x[1540]), .A(y[1540]), .Z(n26797) );
  NANDN U9479 ( .A(x[1539]), .B(y[1539]), .Z(n4375) );
  NANDN U9480 ( .A(x[1540]), .B(y[1540]), .Z(n4374) );
  AND U9481 ( .A(n4375), .B(n4374), .Z(n26795) );
  NANDN U9482 ( .A(y[1538]), .B(x[1538]), .Z(n4377) );
  NANDN U9483 ( .A(y[1539]), .B(x[1539]), .Z(n4376) );
  NAND U9484 ( .A(n4377), .B(n4376), .Z(n26794) );
  NANDN U9485 ( .A(y[1537]), .B(x[1537]), .Z(n4385) );
  XNOR U9486 ( .A(y[1537]), .B(x[1537]), .Z(n4379) );
  NANDN U9487 ( .A(x[1536]), .B(y[1536]), .Z(n4378) );
  NAND U9488 ( .A(n4379), .B(n4378), .Z(n4380) );
  NAND U9489 ( .A(n4385), .B(n4380), .Z(n4382) );
  NANDN U9490 ( .A(x[1538]), .B(y[1538]), .Z(n4381) );
  AND U9491 ( .A(n4382), .B(n4381), .Z(n26793) );
  NANDN U9492 ( .A(y[1536]), .B(x[1536]), .Z(n4384) );
  NANDN U9493 ( .A(y[1535]), .B(x[1535]), .Z(n4383) );
  AND U9494 ( .A(n4384), .B(n4383), .Z(n4386) );
  NAND U9495 ( .A(n4386), .B(n4385), .Z(n17848) );
  ANDN U9496 ( .B(x[1534]), .A(y[1534]), .Z(n17844) );
  NANDN U9497 ( .A(x[1535]), .B(y[1535]), .Z(n4389) );
  NAND U9498 ( .A(n17844), .B(n4389), .Z(n4387) );
  NANDN U9499 ( .A(n17848), .B(n4387), .Z(n26792) );
  NANDN U9500 ( .A(x[1533]), .B(y[1533]), .Z(n13487) );
  NANDN U9501 ( .A(x[1534]), .B(y[1534]), .Z(n4388) );
  AND U9502 ( .A(n4389), .B(n4388), .Z(n26791) );
  ANDN U9503 ( .B(x[1533]), .A(y[1533]), .Z(n26790) );
  NANDN U9504 ( .A(y[1532]), .B(x[1532]), .Z(n26789) );
  NANDN U9505 ( .A(n26790), .B(n26789), .Z(n7622) );
  NANDN U9506 ( .A(x[1531]), .B(y[1531]), .Z(n17837) );
  ANDN U9507 ( .B(x[1531]), .A(y[1531]), .Z(n17841) );
  NANDN U9508 ( .A(y[1530]), .B(x[1530]), .Z(n17832) );
  NANDN U9509 ( .A(n17841), .B(n17832), .Z(n24394) );
  ANDN U9510 ( .B(y[1529]), .A(x[1529]), .Z(n17828) );
  ANDN U9511 ( .B(y[1530]), .A(x[1530]), .Z(n17836) );
  NOR U9512 ( .A(n17828), .B(n17836), .Z(n26787) );
  NANDN U9513 ( .A(x[1527]), .B(y[1527]), .Z(n17823) );
  NANDN U9514 ( .A(x[1528]), .B(y[1528]), .Z(n13489) );
  AND U9515 ( .A(n17823), .B(n13489), .Z(n7615) );
  ANDN U9516 ( .B(x[1526]), .A(y[1526]), .Z(n13490) );
  NANDN U9517 ( .A(y[1527]), .B(x[1527]), .Z(n26784) );
  NANDN U9518 ( .A(y[1524]), .B(x[1524]), .Z(n13495) );
  ANDN U9519 ( .B(y[1523]), .A(x[1523]), .Z(n13498) );
  NANDN U9520 ( .A(x[1522]), .B(y[1522]), .Z(n4391) );
  NANDN U9521 ( .A(x[1521]), .B(y[1521]), .Z(n4390) );
  AND U9522 ( .A(n4391), .B(n4390), .Z(n4395) );
  NANDN U9523 ( .A(x[1520]), .B(y[1520]), .Z(n4393) );
  NANDN U9524 ( .A(x[1519]), .B(y[1519]), .Z(n4392) );
  AND U9525 ( .A(n4393), .B(n4392), .Z(n4394) );
  NAND U9526 ( .A(n4395), .B(n4394), .Z(n13499) );
  NANDN U9527 ( .A(y[1519]), .B(x[1519]), .Z(n13497) );
  NANDN U9528 ( .A(y[1518]), .B(x[1518]), .Z(n4396) );
  AND U9529 ( .A(n13497), .B(n4396), .Z(n26777) );
  NANDN U9530 ( .A(x[1518]), .B(y[1518]), .Z(n13496) );
  NANDN U9531 ( .A(y[1516]), .B(x[1516]), .Z(n17810) );
  NANDN U9532 ( .A(y[1517]), .B(x[1517]), .Z(n13500) );
  NAND U9533 ( .A(n17810), .B(n13500), .Z(n24395) );
  NANDN U9534 ( .A(y[1514]), .B(x[1514]), .Z(n26772) );
  NANDN U9535 ( .A(y[1515]), .B(x[1515]), .Z(n26774) );
  AND U9536 ( .A(n26772), .B(n26774), .Z(n7597) );
  ANDN U9537 ( .B(y[1511]), .A(x[1511]), .Z(n17798) );
  NANDN U9538 ( .A(y[1510]), .B(x[1510]), .Z(n17797) );
  NANDN U9539 ( .A(y[1511]), .B(x[1511]), .Z(n26769) );
  AND U9540 ( .A(n17797), .B(n26769), .Z(n26768) );
  ANDN U9541 ( .B(y[1510]), .A(x[1510]), .Z(n17799) );
  NANDN U9542 ( .A(y[1508]), .B(x[1508]), .Z(n4398) );
  NANDN U9543 ( .A(y[1509]), .B(x[1509]), .Z(n4397) );
  AND U9544 ( .A(n4398), .B(n4397), .Z(n4405) );
  NANDN U9545 ( .A(y[1506]), .B(x[1506]), .Z(n4400) );
  NANDN U9546 ( .A(y[1507]), .B(x[1507]), .Z(n4399) );
  AND U9547 ( .A(n4400), .B(n4399), .Z(n4403) );
  NANDN U9548 ( .A(x[1507]), .B(y[1507]), .Z(n4402) );
  NANDN U9549 ( .A(x[1508]), .B(y[1508]), .Z(n4401) );
  AND U9550 ( .A(n4402), .B(n4401), .Z(n4409) );
  NANDN U9551 ( .A(n4403), .B(n4409), .Z(n4404) );
  AND U9552 ( .A(n4405), .B(n4404), .Z(n26766) );
  NANDN U9553 ( .A(x[1506]), .B(y[1506]), .Z(n4407) );
  NANDN U9554 ( .A(x[1505]), .B(y[1505]), .Z(n4406) );
  AND U9555 ( .A(n4407), .B(n4406), .Z(n4408) );
  AND U9556 ( .A(n4409), .B(n4408), .Z(n13504) );
  NANDN U9557 ( .A(y[1503]), .B(x[1503]), .Z(n4412) );
  ANDN U9558 ( .B(y[1502]), .A(x[1502]), .Z(n17787) );
  NANDN U9559 ( .A(x[1504]), .B(y[1504]), .Z(n4411) );
  NANDN U9560 ( .A(x[1503]), .B(y[1503]), .Z(n4410) );
  NAND U9561 ( .A(n4411), .B(n4410), .Z(n17791) );
  NANDN U9562 ( .A(y[1502]), .B(x[1502]), .Z(n4413) );
  AND U9563 ( .A(n4413), .B(n4412), .Z(n17789) );
  NANDN U9564 ( .A(y[1501]), .B(x[1501]), .Z(n13506) );
  NANDN U9565 ( .A(y[1500]), .B(x[1500]), .Z(n4414) );
  AND U9566 ( .A(n13506), .B(n4414), .Z(n17783) );
  NANDN U9567 ( .A(x[1501]), .B(y[1501]), .Z(n4417) );
  NANDN U9568 ( .A(n17783), .B(n4417), .Z(n4415) );
  NAND U9569 ( .A(n17789), .B(n4415), .Z(n24398) );
  NANDN U9570 ( .A(x[1500]), .B(y[1500]), .Z(n4416) );
  AND U9571 ( .A(n4417), .B(n4416), .Z(n26761) );
  ANDN U9572 ( .B(x[1499]), .A(y[1499]), .Z(n26760) );
  NANDN U9573 ( .A(y[1498]), .B(x[1498]), .Z(n13508) );
  IV U9574 ( .A(n13508), .Z(n26759) );
  OR U9575 ( .A(n26760), .B(n26759), .Z(n7578) );
  NANDN U9576 ( .A(x[1497]), .B(y[1497]), .Z(n26758) );
  ANDN U9577 ( .B(x[1496]), .A(y[1496]), .Z(n17773) );
  NANDN U9578 ( .A(y[1497]), .B(x[1497]), .Z(n13507) );
  NANDN U9579 ( .A(n17773), .B(n13507), .Z(n26757) );
  NANDN U9580 ( .A(x[1496]), .B(y[1496]), .Z(n26756) );
  NANDN U9581 ( .A(x[1495]), .B(y[1495]), .Z(n7570) );
  NANDN U9582 ( .A(x[1494]), .B(y[1494]), .Z(n4418) );
  AND U9583 ( .A(n7570), .B(n4418), .Z(n26754) );
  NANDN U9584 ( .A(x[1493]), .B(y[1493]), .Z(n4420) );
  NANDN U9585 ( .A(x[1492]), .B(y[1492]), .Z(n4419) );
  AND U9586 ( .A(n4420), .B(n4419), .Z(n26752) );
  ANDN U9587 ( .B(y[1489]), .A(x[1489]), .Z(n13511) );
  NANDN U9588 ( .A(y[1490]), .B(x[1490]), .Z(n4424) );
  NAND U9589 ( .A(n13511), .B(n4424), .Z(n7562) );
  NANDN U9590 ( .A(x[1490]), .B(y[1490]), .Z(n4422) );
  NANDN U9591 ( .A(x[1491]), .B(y[1491]), .Z(n4421) );
  NAND U9592 ( .A(n4422), .B(n4421), .Z(n13514) );
  NANDN U9593 ( .A(y[1489]), .B(x[1489]), .Z(n4423) );
  AND U9594 ( .A(n4424), .B(n4423), .Z(n13513) );
  NANDN U9595 ( .A(y[1488]), .B(x[1488]), .Z(n4425) );
  AND U9596 ( .A(n13513), .B(n4425), .Z(n17764) );
  NANDN U9597 ( .A(x[1488]), .B(y[1488]), .Z(n13512) );
  NANDN U9598 ( .A(x[1487]), .B(y[1487]), .Z(n26747) );
  NANDN U9599 ( .A(y[1487]), .B(x[1487]), .Z(n4427) );
  NANDN U9600 ( .A(y[1486]), .B(x[1486]), .Z(n4426) );
  NAND U9601 ( .A(n4427), .B(n4426), .Z(n26746) );
  NANDN U9602 ( .A(x[1486]), .B(y[1486]), .Z(n4429) );
  NANDN U9603 ( .A(x[1485]), .B(y[1485]), .Z(n4428) );
  AND U9604 ( .A(n4429), .B(n4428), .Z(n26745) );
  NANDN U9605 ( .A(x[1484]), .B(y[1484]), .Z(n13515) );
  ANDN U9606 ( .B(y[1483]), .A(x[1483]), .Z(n17755) );
  ANDN U9607 ( .B(n13515), .A(n17755), .Z(n26743) );
  ANDN U9608 ( .B(x[1483]), .A(y[1483]), .Z(n17759) );
  NANDN U9609 ( .A(y[1482]), .B(x[1482]), .Z(n17751) );
  NANDN U9610 ( .A(n17759), .B(n17751), .Z(n26742) );
  NANDN U9611 ( .A(y[1481]), .B(x[1481]), .Z(n26741) );
  NANDN U9612 ( .A(y[1478]), .B(x[1478]), .Z(n17743) );
  NANDN U9613 ( .A(y[1479]), .B(x[1479]), .Z(n17747) );
  AND U9614 ( .A(n17743), .B(n17747), .Z(n26737) );
  ANDN U9615 ( .B(y[1478]), .A(x[1478]), .Z(n26736) );
  ANDN U9616 ( .B(x[1477]), .A(y[1477]), .Z(n26735) );
  NANDN U9617 ( .A(x[1475]), .B(y[1475]), .Z(n4437) );
  XNOR U9618 ( .A(x[1475]), .B(y[1475]), .Z(n4431) );
  NANDN U9619 ( .A(y[1474]), .B(x[1474]), .Z(n4430) );
  NAND U9620 ( .A(n4431), .B(n4430), .Z(n4432) );
  NAND U9621 ( .A(n4437), .B(n4432), .Z(n4434) );
  NANDN U9622 ( .A(y[1476]), .B(x[1476]), .Z(n4433) );
  AND U9623 ( .A(n4434), .B(n4433), .Z(n26733) );
  NANDN U9624 ( .A(x[1474]), .B(y[1474]), .Z(n4436) );
  NANDN U9625 ( .A(x[1473]), .B(y[1473]), .Z(n4435) );
  AND U9626 ( .A(n4436), .B(n4435), .Z(n4438) );
  NAND U9627 ( .A(n4438), .B(n4437), .Z(n13522) );
  NANDN U9628 ( .A(y[1472]), .B(x[1472]), .Z(n4439) );
  ANDN U9629 ( .B(x[1473]), .A(y[1473]), .Z(n13521) );
  ANDN U9630 ( .B(n4439), .A(n13521), .Z(n26731) );
  ANDN U9631 ( .B(y[1472]), .A(x[1472]), .Z(n13520) );
  ANDN U9632 ( .B(y[1471]), .A(x[1471]), .Z(n26730) );
  NOR U9633 ( .A(n13520), .B(n26730), .Z(n7536) );
  ANDN U9634 ( .B(y[1469]), .A(x[1469]), .Z(n17724) );
  ANDN U9635 ( .B(y[1470]), .A(x[1470]), .Z(n17732) );
  NOR U9636 ( .A(n17724), .B(n17732), .Z(n26727) );
  NANDN U9637 ( .A(y[1468]), .B(x[1468]), .Z(n17722) );
  NANDN U9638 ( .A(y[1469]), .B(x[1469]), .Z(n17727) );
  NAND U9639 ( .A(n17722), .B(n17727), .Z(n24401) );
  NANDN U9640 ( .A(y[1467]), .B(x[1467]), .Z(n26725) );
  ANDN U9641 ( .B(y[1464]), .A(x[1464]), .Z(n17714) );
  NANDN U9642 ( .A(x[1463]), .B(y[1463]), .Z(n13527) );
  ANDN U9643 ( .B(x[1463]), .A(y[1463]), .Z(n13525) );
  NANDN U9644 ( .A(x[1462]), .B(y[1462]), .Z(n13528) );
  NANDN U9645 ( .A(y[1461]), .B(x[1461]), .Z(n13530) );
  NANDN U9646 ( .A(y[1460]), .B(x[1460]), .Z(n13534) );
  AND U9647 ( .A(n13530), .B(n13534), .Z(n7518) );
  NANDN U9648 ( .A(x[1459]), .B(y[1459]), .Z(n26716) );
  ANDN U9649 ( .B(x[1458]), .A(y[1458]), .Z(n26714) );
  NANDN U9650 ( .A(x[1457]), .B(y[1457]), .Z(n17703) );
  NANDN U9651 ( .A(x[1458]), .B(y[1458]), .Z(n13535) );
  AND U9652 ( .A(n17703), .B(n13535), .Z(n26713) );
  NANDN U9653 ( .A(y[1456]), .B(x[1456]), .Z(n4441) );
  NANDN U9654 ( .A(y[1457]), .B(x[1457]), .Z(n4440) );
  NAND U9655 ( .A(n4441), .B(n4440), .Z(n26712) );
  NANDN U9656 ( .A(x[1456]), .B(y[1456]), .Z(n4443) );
  NANDN U9657 ( .A(x[1455]), .B(y[1455]), .Z(n4442) );
  AND U9658 ( .A(n4443), .B(n4442), .Z(n26711) );
  NANDN U9659 ( .A(y[1454]), .B(x[1454]), .Z(n4445) );
  NANDN U9660 ( .A(y[1455]), .B(x[1455]), .Z(n4444) );
  NAND U9661 ( .A(n4445), .B(n4444), .Z(n26710) );
  NANDN U9662 ( .A(x[1454]), .B(y[1454]), .Z(n4447) );
  NANDN U9663 ( .A(x[1453]), .B(y[1453]), .Z(n4446) );
  AND U9664 ( .A(n4447), .B(n4446), .Z(n26709) );
  NANDN U9665 ( .A(y[1452]), .B(x[1452]), .Z(n4449) );
  NANDN U9666 ( .A(y[1453]), .B(x[1453]), .Z(n4448) );
  NAND U9667 ( .A(n4449), .B(n4448), .Z(n26708) );
  NANDN U9668 ( .A(x[1452]), .B(y[1452]), .Z(n4451) );
  NANDN U9669 ( .A(x[1451]), .B(y[1451]), .Z(n4450) );
  AND U9670 ( .A(n4451), .B(n4450), .Z(n26707) );
  NANDN U9671 ( .A(y[1450]), .B(x[1450]), .Z(n4453) );
  NANDN U9672 ( .A(y[1451]), .B(x[1451]), .Z(n4452) );
  NAND U9673 ( .A(n4453), .B(n4452), .Z(n26706) );
  NANDN U9674 ( .A(x[1450]), .B(y[1450]), .Z(n4455) );
  NANDN U9675 ( .A(x[1449]), .B(y[1449]), .Z(n4454) );
  AND U9676 ( .A(n4455), .B(n4454), .Z(n13538) );
  ANDN U9677 ( .B(x[1449]), .A(y[1449]), .Z(n13537) );
  NANDN U9678 ( .A(y[1448]), .B(x[1448]), .Z(n4456) );
  NANDN U9679 ( .A(n13537), .B(n4456), .Z(n26704) );
  ANDN U9680 ( .B(x[1446]), .A(y[1446]), .Z(n17684) );
  ANDN U9681 ( .B(x[1447]), .A(y[1447]), .Z(n17693) );
  NOR U9682 ( .A(n17684), .B(n17693), .Z(n26702) );
  NANDN U9683 ( .A(x[1445]), .B(y[1445]), .Z(n17682) );
  NANDN U9684 ( .A(x[1446]), .B(y[1446]), .Z(n17689) );
  NAND U9685 ( .A(n17682), .B(n17689), .Z(n26701) );
  ANDN U9686 ( .B(x[1444]), .A(y[1444]), .Z(n17681) );
  ANDN U9687 ( .B(x[1445]), .A(y[1445]), .Z(n17687) );
  NOR U9688 ( .A(n17681), .B(n17687), .Z(n26700) );
  NANDN U9689 ( .A(x[1443]), .B(y[1443]), .Z(n4458) );
  NANDN U9690 ( .A(x[1444]), .B(y[1444]), .Z(n4457) );
  NAND U9691 ( .A(n4458), .B(n4457), .Z(n13541) );
  NANDN U9692 ( .A(y[1442]), .B(x[1442]), .Z(n4459) );
  ANDN U9693 ( .B(x[1443]), .A(y[1443]), .Z(n13540) );
  ANDN U9694 ( .B(n4459), .A(n13540), .Z(n7494) );
  ANDN U9695 ( .B(y[1442]), .A(x[1442]), .Z(n13539) );
  NANDN U9696 ( .A(x[1441]), .B(y[1441]), .Z(n13543) );
  NANDN U9697 ( .A(n13539), .B(n13543), .Z(n4460) );
  NAND U9698 ( .A(n7494), .B(n4460), .Z(n4461) );
  NANDN U9699 ( .A(n13541), .B(n4461), .Z(n7497) );
  ANDN U9700 ( .B(y[1432]), .A(x[1432]), .Z(n4462) );
  NAND U9701 ( .A(n4462), .B(y[1433]), .Z(n4465) );
  XOR U9702 ( .A(n4462), .B(y[1433]), .Z(n4463) );
  NANDN U9703 ( .A(x[1433]), .B(n4463), .Z(n4464) );
  AND U9704 ( .A(n4465), .B(n4464), .Z(n26690) );
  NANDN U9705 ( .A(y[1432]), .B(x[1432]), .Z(n4467) );
  NANDN U9706 ( .A(y[1431]), .B(x[1431]), .Z(n4466) );
  AND U9707 ( .A(n4467), .B(n4466), .Z(n4469) );
  NANDN U9708 ( .A(y[1433]), .B(x[1433]), .Z(n4468) );
  NAND U9709 ( .A(n4469), .B(n4468), .Z(n26689) );
  NANDN U9710 ( .A(y[1428]), .B(x[1428]), .Z(n17665) );
  NANDN U9711 ( .A(x[1426]), .B(y[1426]), .Z(n17662) );
  NANDN U9712 ( .A(y[1426]), .B(x[1426]), .Z(n4471) );
  NANDN U9713 ( .A(y[1425]), .B(x[1425]), .Z(n4470) );
  NAND U9714 ( .A(n4471), .B(n4470), .Z(n17659) );
  ANDN U9715 ( .B(x[1424]), .A(y[1424]), .Z(n17653) );
  NANDN U9716 ( .A(x[1425]), .B(y[1425]), .Z(n4474) );
  NAND U9717 ( .A(n17653), .B(n4474), .Z(n4472) );
  NANDN U9718 ( .A(n17659), .B(n4472), .Z(n26683) );
  NANDN U9719 ( .A(x[1424]), .B(y[1424]), .Z(n4473) );
  AND U9720 ( .A(n4474), .B(n4473), .Z(n17658) );
  NANDN U9721 ( .A(x[1423]), .B(y[1423]), .Z(n17650) );
  AND U9722 ( .A(n17658), .B(n17650), .Z(n24404) );
  NANDN U9723 ( .A(y[1422]), .B(x[1422]), .Z(n17647) );
  ANDN U9724 ( .B(x[1423]), .A(y[1423]), .Z(n17656) );
  ANDN U9725 ( .B(n17647), .A(n17656), .Z(n26682) );
  ANDN U9726 ( .B(y[1421]), .A(x[1421]), .Z(n17645) );
  NANDN U9727 ( .A(x[1422]), .B(y[1422]), .Z(n17651) );
  NANDN U9728 ( .A(n17645), .B(n17651), .Z(n26681) );
  NANDN U9729 ( .A(y[1420]), .B(x[1420]), .Z(n26677) );
  ANDN U9730 ( .B(x[1421]), .A(y[1421]), .Z(n26679) );
  ANDN U9731 ( .B(n26677), .A(n26679), .Z(n7450) );
  ANDN U9732 ( .B(y[1420]), .A(x[1420]), .Z(n26678) );
  NANDN U9733 ( .A(y[1418]), .B(x[1418]), .Z(n17634) );
  NANDN U9734 ( .A(y[1419]), .B(x[1419]), .Z(n17640) );
  AND U9735 ( .A(n17634), .B(n17640), .Z(n26675) );
  ANDN U9736 ( .B(y[1417]), .A(x[1417]), .Z(n17631) );
  ANDN U9737 ( .B(y[1418]), .A(x[1418]), .Z(n17637) );
  OR U9738 ( .A(n17631), .B(n17637), .Z(n26674) );
  NANDN U9739 ( .A(y[1416]), .B(x[1416]), .Z(n17627) );
  NANDN U9740 ( .A(y[1417]), .B(x[1417]), .Z(n17635) );
  AND U9741 ( .A(n17627), .B(n17635), .Z(n26673) );
  NANDN U9742 ( .A(y[1414]), .B(x[1414]), .Z(n26669) );
  NANDN U9743 ( .A(y[1415]), .B(x[1415]), .Z(n26671) );
  AND U9744 ( .A(n26669), .B(n26671), .Z(n7441) );
  NANDN U9745 ( .A(y[1412]), .B(x[1412]), .Z(n17618) );
  NANDN U9746 ( .A(y[1413]), .B(x[1413]), .Z(n17623) );
  NAND U9747 ( .A(n17618), .B(n17623), .Z(n24406) );
  NANDN U9748 ( .A(x[1411]), .B(y[1411]), .Z(n13549) );
  NANDN U9749 ( .A(y[1410]), .B(x[1410]), .Z(n26665) );
  NANDN U9750 ( .A(y[1411]), .B(x[1411]), .Z(n26667) );
  NAND U9751 ( .A(n26665), .B(n26667), .Z(n7434) );
  NANDN U9752 ( .A(x[1409]), .B(y[1409]), .Z(n17613) );
  NANDN U9753 ( .A(y[1408]), .B(x[1408]), .Z(n17609) );
  NANDN U9754 ( .A(y[1409]), .B(x[1409]), .Z(n13551) );
  NAND U9755 ( .A(n17609), .B(n13551), .Z(n24407) );
  NANDN U9756 ( .A(x[1408]), .B(y[1408]), .Z(n13552) );
  NANDN U9757 ( .A(y[1406]), .B(x[1406]), .Z(n26659) );
  NANDN U9758 ( .A(y[1407]), .B(x[1407]), .Z(n26661) );
  NAND U9759 ( .A(n26659), .B(n26661), .Z(n7427) );
  ANDN U9760 ( .B(y[1405]), .A(x[1405]), .Z(n26658) );
  NANDN U9761 ( .A(y[1404]), .B(x[1404]), .Z(n17603) );
  NANDN U9762 ( .A(y[1405]), .B(x[1405]), .Z(n17605) );
  NAND U9763 ( .A(n17603), .B(n17605), .Z(n26657) );
  NANDN U9764 ( .A(x[1404]), .B(y[1404]), .Z(n4476) );
  NANDN U9765 ( .A(x[1403]), .B(y[1403]), .Z(n4475) );
  AND U9766 ( .A(n4476), .B(n4475), .Z(n26656) );
  NANDN U9767 ( .A(x[1401]), .B(y[1401]), .Z(n17595) );
  NANDN U9768 ( .A(x[1402]), .B(y[1402]), .Z(n13555) );
  AND U9769 ( .A(n17595), .B(n13555), .Z(n26654) );
  ANDN U9770 ( .B(x[1400]), .A(y[1400]), .Z(n17592) );
  ANDN U9771 ( .B(x[1401]), .A(y[1401]), .Z(n17599) );
  OR U9772 ( .A(n17592), .B(n17599), .Z(n26653) );
  NANDN U9773 ( .A(x[1400]), .B(y[1400]), .Z(n26652) );
  ANDN U9774 ( .B(x[1399]), .A(y[1399]), .Z(n26651) );
  ANDN U9775 ( .B(x[1398]), .A(y[1398]), .Z(n7414) );
  NANDN U9776 ( .A(x[1397]), .B(y[1397]), .Z(n13562) );
  XNOR U9777 ( .A(x[1398]), .B(y[1398]), .Z(n13561) );
  NANDN U9778 ( .A(y[1396]), .B(x[1396]), .Z(n13565) );
  NANDN U9779 ( .A(x[1396]), .B(y[1396]), .Z(n13563) );
  ANDN U9780 ( .B(x[1394]), .A(y[1394]), .Z(n26645) );
  NANDN U9781 ( .A(x[1393]), .B(y[1393]), .Z(n17578) );
  NANDN U9782 ( .A(x[1394]), .B(y[1394]), .Z(n17585) );
  AND U9783 ( .A(n17578), .B(n17585), .Z(n26643) );
  ANDN U9784 ( .B(x[1392]), .A(y[1392]), .Z(n17577) );
  ANDN U9785 ( .B(x[1393]), .A(y[1393]), .Z(n17582) );
  OR U9786 ( .A(n17577), .B(n17582), .Z(n26641) );
  NANDN U9787 ( .A(x[1391]), .B(y[1391]), .Z(n13567) );
  NANDN U9788 ( .A(x[1392]), .B(y[1392]), .Z(n26639) );
  AND U9789 ( .A(n13567), .B(n26639), .Z(n7402) );
  ANDN U9790 ( .B(x[1391]), .A(y[1391]), .Z(n26637) );
  NANDN U9791 ( .A(y[1388]), .B(x[1388]), .Z(n13571) );
  NANDN U9792 ( .A(y[1389]), .B(x[1389]), .Z(n13569) );
  AND U9793 ( .A(n13571), .B(n13569), .Z(n26629) );
  NANDN U9794 ( .A(x[1387]), .B(y[1387]), .Z(n17566) );
  NANDN U9795 ( .A(x[1388]), .B(y[1388]), .Z(n13570) );
  NAND U9796 ( .A(n17566), .B(n13570), .Z(n26627) );
  ANDN U9797 ( .B(x[1386]), .A(y[1386]), .Z(n17564) );
  NANDN U9798 ( .A(y[1387]), .B(x[1387]), .Z(n13572) );
  NANDN U9799 ( .A(n17564), .B(n13572), .Z(n26625) );
  NANDN U9800 ( .A(x[1386]), .B(y[1386]), .Z(n26623) );
  ANDN U9801 ( .B(x[1385]), .A(y[1385]), .Z(n26621) );
  NANDN U9802 ( .A(x[1384]), .B(y[1384]), .Z(n4478) );
  NANDN U9803 ( .A(x[1385]), .B(y[1385]), .Z(n4477) );
  AND U9804 ( .A(n4478), .B(n4477), .Z(n26619) );
  ANDN U9805 ( .B(x[1384]), .A(y[1384]), .Z(n26617) );
  NANDN U9806 ( .A(x[1383]), .B(y[1383]), .Z(n26614) );
  NANDN U9807 ( .A(y[1383]), .B(x[1383]), .Z(n4480) );
  NANDN U9808 ( .A(y[1382]), .B(x[1382]), .Z(n4479) );
  NAND U9809 ( .A(n4480), .B(n4479), .Z(n26613) );
  ANDN U9810 ( .B(x[1381]), .A(y[1381]), .Z(n17556) );
  ANDN U9811 ( .B(x[1380]), .A(y[1380]), .Z(n17550) );
  NOR U9812 ( .A(n17556), .B(n17550), .Z(n26608) );
  NANDN U9813 ( .A(y[1376]), .B(x[1376]), .Z(n4481) );
  NANDN U9814 ( .A(y[1377]), .B(x[1377]), .Z(n13575) );
  AND U9815 ( .A(n4481), .B(n13575), .Z(n13578) );
  NANDN U9816 ( .A(x[1375]), .B(y[1375]), .Z(n26600) );
  NANDN U9817 ( .A(x[1376]), .B(y[1376]), .Z(n13576) );
  NAND U9818 ( .A(n26600), .B(n13576), .Z(n7374) );
  NANDN U9819 ( .A(y[1375]), .B(x[1375]), .Z(n13577) );
  XNOR U9820 ( .A(x[1374]), .B(y[1374]), .Z(n17543) );
  NANDN U9821 ( .A(y[1372]), .B(x[1372]), .Z(n17540) );
  ANDN U9822 ( .B(x[1370]), .A(y[1370]), .Z(n13583) );
  ANDN U9823 ( .B(x[1371]), .A(y[1371]), .Z(n17539) );
  NOR U9824 ( .A(n13583), .B(n17539), .Z(n26594) );
  ANDN U9825 ( .B(y[1369]), .A(x[1369]), .Z(n17530) );
  NANDN U9826 ( .A(x[1370]), .B(y[1370]), .Z(n17535) );
  NANDN U9827 ( .A(n17530), .B(n17535), .Z(n24408) );
  ANDN U9828 ( .B(x[1369]), .A(y[1369]), .Z(n13582) );
  NANDN U9829 ( .A(y[1368]), .B(x[1368]), .Z(n17526) );
  NANDN U9830 ( .A(n13582), .B(n17526), .Z(n26593) );
  ANDN U9831 ( .B(y[1368]), .A(x[1368]), .Z(n26592) );
  NANDN U9832 ( .A(y[1367]), .B(x[1367]), .Z(n26591) );
  ANDN U9833 ( .B(x[1366]), .A(y[1366]), .Z(n13586) );
  ANDN U9834 ( .B(n26591), .A(n13586), .Z(n7359) );
  ANDN U9835 ( .B(y[1365]), .A(x[1365]), .Z(n17521) );
  NANDN U9836 ( .A(y[1365]), .B(x[1365]), .Z(n13587) );
  ANDN U9837 ( .B(y[1363]), .A(x[1363]), .Z(n26585) );
  NANDN U9838 ( .A(y[1360]), .B(x[1360]), .Z(n17506) );
  NANDN U9839 ( .A(y[1361]), .B(x[1361]), .Z(n13588) );
  AND U9840 ( .A(n17506), .B(n13588), .Z(n26583) );
  NANDN U9841 ( .A(y[1358]), .B(x[1358]), .Z(n26579) );
  NANDN U9842 ( .A(y[1359]), .B(x[1359]), .Z(n26581) );
  NAND U9843 ( .A(n26579), .B(n26581), .Z(n7345) );
  NANDN U9844 ( .A(x[1357]), .B(y[1357]), .Z(n26577) );
  NANDN U9845 ( .A(y[1356]), .B(x[1356]), .Z(n13592) );
  NANDN U9846 ( .A(y[1357]), .B(x[1357]), .Z(n17502) );
  NAND U9847 ( .A(n13592), .B(n17502), .Z(n26578) );
  NANDN U9848 ( .A(x[1355]), .B(y[1355]), .Z(n13593) );
  NANDN U9849 ( .A(y[1354]), .B(x[1354]), .Z(n13595) );
  NANDN U9850 ( .A(y[1355]), .B(x[1355]), .Z(n24411) );
  NAND U9851 ( .A(n13595), .B(n24411), .Z(n26573) );
  NANDN U9852 ( .A(x[1353]), .B(y[1353]), .Z(n13597) );
  NANDN U9853 ( .A(y[1353]), .B(x[1353]), .Z(n13596) );
  ANDN U9854 ( .B(x[1352]), .A(y[1352]), .Z(n17491) );
  ANDN U9855 ( .B(n13596), .A(n17491), .Z(n26571) );
  NANDN U9856 ( .A(x[1351]), .B(y[1351]), .Z(n17487) );
  ANDN U9857 ( .B(y[1352]), .A(x[1352]), .Z(n13598) );
  ANDN U9858 ( .B(n17487), .A(n13598), .Z(n26570) );
  ANDN U9859 ( .B(x[1350]), .A(y[1350]), .Z(n17482) );
  ANDN U9860 ( .B(x[1351]), .A(y[1351]), .Z(n17492) );
  OR U9861 ( .A(n17482), .B(n17492), .Z(n24412) );
  NANDN U9862 ( .A(x[1349]), .B(y[1349]), .Z(n17479) );
  NANDN U9863 ( .A(x[1350]), .B(y[1350]), .Z(n17486) );
  AND U9864 ( .A(n17479), .B(n17486), .Z(n26569) );
  ANDN U9865 ( .B(x[1348]), .A(y[1348]), .Z(n17475) );
  ANDN U9866 ( .B(x[1349]), .A(y[1349]), .Z(n17485) );
  OR U9867 ( .A(n17475), .B(n17485), .Z(n26568) );
  NANDN U9868 ( .A(x[1347]), .B(y[1347]), .Z(n17471) );
  NANDN U9869 ( .A(x[1348]), .B(y[1348]), .Z(n17480) );
  AND U9870 ( .A(n17471), .B(n17480), .Z(n26567) );
  ANDN U9871 ( .B(x[1347]), .A(y[1347]), .Z(n17477) );
  NANDN U9872 ( .A(y[1346]), .B(x[1346]), .Z(n13599) );
  NANDN U9873 ( .A(n17477), .B(n13599), .Z(n26566) );
  NANDN U9874 ( .A(y[1345]), .B(x[1345]), .Z(n13600) );
  NANDN U9875 ( .A(y[1344]), .B(x[1344]), .Z(n17464) );
  NANDN U9876 ( .A(x[1345]), .B(y[1345]), .Z(n4484) );
  NANDN U9877 ( .A(n17464), .B(n4484), .Z(n4482) );
  NAND U9878 ( .A(n13600), .B(n4482), .Z(n24413) );
  NANDN U9879 ( .A(x[1344]), .B(y[1344]), .Z(n4483) );
  AND U9880 ( .A(n4484), .B(n4483), .Z(n17468) );
  ANDN U9881 ( .B(y[1343]), .A(x[1343]), .Z(n17460) );
  ANDN U9882 ( .B(n17468), .A(n17460), .Z(n26564) );
  ANDN U9883 ( .B(x[1343]), .A(y[1343]), .Z(n17466) );
  NANDN U9884 ( .A(y[1342]), .B(x[1342]), .Z(n17456) );
  NANDN U9885 ( .A(n17466), .B(n17456), .Z(n26563) );
  NANDN U9886 ( .A(x[1341]), .B(y[1341]), .Z(n13602) );
  ANDN U9887 ( .B(y[1342]), .A(x[1342]), .Z(n17462) );
  ANDN U9888 ( .B(n13602), .A(n17462), .Z(n26562) );
  ANDN U9889 ( .B(x[1340]), .A(y[1340]), .Z(n17450) );
  NANDN U9890 ( .A(y[1341]), .B(x[1341]), .Z(n17455) );
  NANDN U9891 ( .A(n17450), .B(n17455), .Z(n26561) );
  NANDN U9892 ( .A(x[1340]), .B(y[1340]), .Z(n13601) );
  NANDN U9893 ( .A(x[1339]), .B(y[1339]), .Z(n4486) );
  NANDN U9894 ( .A(x[1338]), .B(y[1338]), .Z(n4485) );
  AND U9895 ( .A(n4486), .B(n4485), .Z(n17448) );
  NANDN U9896 ( .A(y[1339]), .B(x[1339]), .Z(n4490) );
  IV U9897 ( .A(n4490), .Z(n17451) );
  OR U9898 ( .A(n17448), .B(n17451), .Z(n4487) );
  AND U9899 ( .A(n13601), .B(n4487), .Z(n26560) );
  NANDN U9900 ( .A(y[1338]), .B(x[1338]), .Z(n4489) );
  NANDN U9901 ( .A(y[1337]), .B(x[1337]), .Z(n4488) );
  NAND U9902 ( .A(n4489), .B(n4488), .Z(n17446) );
  ANDN U9903 ( .B(n4490), .A(n17446), .Z(n26559) );
  NANDN U9904 ( .A(x[1336]), .B(y[1336]), .Z(n4492) );
  NANDN U9905 ( .A(x[1337]), .B(y[1337]), .Z(n4491) );
  NAND U9906 ( .A(n4492), .B(n4491), .Z(n17443) );
  NANDN U9907 ( .A(y[1336]), .B(x[1336]), .Z(n4494) );
  NANDN U9908 ( .A(y[1335]), .B(x[1335]), .Z(n4493) );
  AND U9909 ( .A(n4494), .B(n4493), .Z(n13603) );
  NANDN U9910 ( .A(y[1332]), .B(x[1332]), .Z(n13605) );
  ANDN U9911 ( .B(y[1330]), .A(x[1330]), .Z(n13606) );
  NANDN U9912 ( .A(y[1330]), .B(x[1330]), .Z(n4496) );
  NANDN U9913 ( .A(y[1329]), .B(x[1329]), .Z(n4495) );
  AND U9914 ( .A(n4496), .B(n4495), .Z(n26550) );
  NANDN U9915 ( .A(x[1329]), .B(y[1329]), .Z(n4498) );
  NANDN U9916 ( .A(x[1328]), .B(y[1328]), .Z(n4497) );
  AND U9917 ( .A(n4498), .B(n4497), .Z(n26549) );
  NANDN U9918 ( .A(y[1328]), .B(x[1328]), .Z(n4500) );
  NANDN U9919 ( .A(y[1327]), .B(x[1327]), .Z(n4499) );
  NAND U9920 ( .A(n4500), .B(n4499), .Z(n17432) );
  ANDN U9921 ( .B(x[1326]), .A(y[1326]), .Z(n17428) );
  NANDN U9922 ( .A(x[1327]), .B(y[1327]), .Z(n4503) );
  NAND U9923 ( .A(n17428), .B(n4503), .Z(n4501) );
  NANDN U9924 ( .A(n17432), .B(n4501), .Z(n24414) );
  NANDN U9925 ( .A(x[1325]), .B(y[1325]), .Z(n13607) );
  NANDN U9926 ( .A(x[1326]), .B(y[1326]), .Z(n4502) );
  AND U9927 ( .A(n4503), .B(n4502), .Z(n26548) );
  NANDN U9928 ( .A(y[1324]), .B(x[1324]), .Z(n26547) );
  NANDN U9929 ( .A(y[1325]), .B(x[1325]), .Z(n24415) );
  NAND U9930 ( .A(n26547), .B(n24415), .Z(n7298) );
  ANDN U9931 ( .B(y[1323]), .A(x[1323]), .Z(n26545) );
  ANDN U9932 ( .B(x[1322]), .A(y[1322]), .Z(n17419) );
  NANDN U9933 ( .A(y[1323]), .B(x[1323]), .Z(n17424) );
  NANDN U9934 ( .A(n17419), .B(n17424), .Z(n26544) );
  NANDN U9935 ( .A(x[1321]), .B(y[1321]), .Z(n17415) );
  ANDN U9936 ( .B(y[1322]), .A(x[1322]), .Z(n13609) );
  ANDN U9937 ( .B(n17415), .A(n13609), .Z(n26543) );
  ANDN U9938 ( .B(x[1320]), .A(y[1320]), .Z(n17413) );
  ANDN U9939 ( .B(x[1321]), .A(y[1321]), .Z(n17420) );
  OR U9940 ( .A(n17413), .B(n17420), .Z(n26542) );
  NANDN U9941 ( .A(x[1319]), .B(y[1319]), .Z(n17411) );
  NANDN U9942 ( .A(x[1320]), .B(y[1320]), .Z(n17414) );
  AND U9943 ( .A(n17411), .B(n17414), .Z(n26541) );
  NANDN U9944 ( .A(y[1318]), .B(x[1318]), .Z(n4505) );
  NANDN U9945 ( .A(y[1319]), .B(x[1319]), .Z(n4504) );
  NAND U9946 ( .A(n4505), .B(n4504), .Z(n26540) );
  ANDN U9947 ( .B(y[1317]), .A(x[1317]), .Z(n13611) );
  NANDN U9948 ( .A(y[1316]), .B(x[1316]), .Z(n4506) );
  NANDN U9949 ( .A(y[1317]), .B(x[1317]), .Z(n13610) );
  AND U9950 ( .A(n4506), .B(n13610), .Z(n26538) );
  ANDN U9951 ( .B(y[1315]), .A(x[1315]), .Z(n26537) );
  NANDN U9952 ( .A(y[1314]), .B(x[1314]), .Z(n13614) );
  ANDN U9953 ( .B(x[1315]), .A(y[1315]), .Z(n17407) );
  ANDN U9954 ( .B(n13614), .A(n17407), .Z(n26536) );
  NANDN U9955 ( .A(y[1311]), .B(x[1311]), .Z(n26535) );
  NANDN U9956 ( .A(y[1310]), .B(x[1310]), .Z(n26533) );
  AND U9957 ( .A(n26535), .B(n26533), .Z(n7279) );
  ANDN U9958 ( .B(y[1310]), .A(x[1310]), .Z(n13616) );
  ANDN U9959 ( .B(x[1307]), .A(y[1307]), .Z(n13620) );
  NANDN U9960 ( .A(x[1306]), .B(y[1306]), .Z(n4508) );
  NANDN U9961 ( .A(x[1307]), .B(y[1307]), .Z(n4507) );
  AND U9962 ( .A(n4508), .B(n4507), .Z(n24420) );
  NANDN U9963 ( .A(y[1306]), .B(x[1306]), .Z(n4510) );
  NANDN U9964 ( .A(y[1305]), .B(x[1305]), .Z(n4509) );
  NAND U9965 ( .A(n4510), .B(n4509), .Z(n17382) );
  ANDN U9966 ( .B(x[1304]), .A(y[1304]), .Z(n17378) );
  NANDN U9967 ( .A(x[1305]), .B(y[1305]), .Z(n7268) );
  NAND U9968 ( .A(n17378), .B(n7268), .Z(n4511) );
  NANDN U9969 ( .A(n17382), .B(n4511), .Z(n24421) );
  NANDN U9970 ( .A(x[1303]), .B(y[1303]), .Z(n13621) );
  ANDN U9971 ( .B(x[1302]), .A(y[1302]), .Z(n13623) );
  NANDN U9972 ( .A(x[1301]), .B(y[1301]), .Z(n13626) );
  NANDN U9973 ( .A(y[1300]), .B(x[1300]), .Z(n13627) );
  ANDN U9974 ( .B(y[1299]), .A(x[1299]), .Z(n13629) );
  NANDN U9975 ( .A(y[1299]), .B(x[1299]), .Z(n13628) );
  ANDN U9976 ( .B(x[1292]), .A(y[1292]), .Z(n13637) );
  NANDN U9977 ( .A(x[1292]), .B(y[1292]), .Z(n13636) );
  ANDN U9978 ( .B(x[1290]), .A(y[1290]), .Z(n13643) );
  NANDN U9979 ( .A(y[1287]), .B(x[1287]), .Z(n13646) );
  NANDN U9980 ( .A(y[1286]), .B(x[1286]), .Z(n4512) );
  NAND U9981 ( .A(n13646), .B(n4512), .Z(n26509) );
  NANDN U9982 ( .A(x[1285]), .B(y[1285]), .Z(n13648) );
  XNOR U9983 ( .A(y[1286]), .B(x[1286]), .Z(n13647) );
  NANDN U9984 ( .A(x[1283]), .B(y[1283]), .Z(n17344) );
  ANDN U9985 ( .B(y[1284]), .A(x[1284]), .Z(n13649) );
  ANDN U9986 ( .B(n17344), .A(n13649), .Z(n26507) );
  ANDN U9987 ( .B(x[1282]), .A(y[1282]), .Z(n17339) );
  ANDN U9988 ( .B(x[1283]), .A(y[1283]), .Z(n17349) );
  OR U9989 ( .A(n17339), .B(n17349), .Z(n24425) );
  NANDN U9990 ( .A(x[1281]), .B(y[1281]), .Z(n17336) );
  NANDN U9991 ( .A(x[1282]), .B(y[1282]), .Z(n17343) );
  AND U9992 ( .A(n17336), .B(n17343), .Z(n26506) );
  ANDN U9993 ( .B(x[1280]), .A(y[1280]), .Z(n17332) );
  ANDN U9994 ( .B(x[1281]), .A(y[1281]), .Z(n17342) );
  OR U9995 ( .A(n17332), .B(n17342), .Z(n26505) );
  NANDN U9996 ( .A(x[1279]), .B(y[1279]), .Z(n17328) );
  NANDN U9997 ( .A(x[1280]), .B(y[1280]), .Z(n17337) );
  AND U9998 ( .A(n17328), .B(n17337), .Z(n26504) );
  ANDN U9999 ( .B(x[1278]), .A(y[1278]), .Z(n17327) );
  ANDN U10000 ( .B(x[1279]), .A(y[1279]), .Z(n17334) );
  OR U10001 ( .A(n17327), .B(n17334), .Z(n26502) );
  NANDN U10002 ( .A(x[1277]), .B(y[1277]), .Z(n13651) );
  NANDN U10003 ( .A(x[1278]), .B(y[1278]), .Z(n26501) );
  AND U10004 ( .A(n13651), .B(n26501), .Z(n7222) );
  ANDN U10005 ( .B(x[1277]), .A(y[1277]), .Z(n26500) );
  NANDN U10006 ( .A(y[1276]), .B(x[1276]), .Z(n13652) );
  ANDN U10007 ( .B(y[1275]), .A(x[1275]), .Z(n13654) );
  NANDN U10008 ( .A(y[1275]), .B(x[1275]), .Z(n13653) );
  NANDN U10009 ( .A(x[1273]), .B(y[1273]), .Z(n4513) );
  ANDN U10010 ( .B(y[1274]), .A(x[1274]), .Z(n17317) );
  ANDN U10011 ( .B(n4513), .A(n17317), .Z(n7213) );
  NANDN U10012 ( .A(x[1272]), .B(y[1272]), .Z(n4514) );
  NAND U10013 ( .A(n7213), .B(n4514), .Z(n17314) );
  NANDN U10014 ( .A(y[1271]), .B(x[1271]), .Z(n24426) );
  XNOR U10015 ( .A(x[1270]), .B(y[1270]), .Z(n7204) );
  NANDN U10016 ( .A(y[1269]), .B(x[1269]), .Z(n4515) );
  AND U10017 ( .A(n7204), .B(n4515), .Z(n17307) );
  NANDN U10018 ( .A(y[1268]), .B(x[1268]), .Z(n13657) );
  ANDN U10019 ( .B(y[1267]), .A(x[1267]), .Z(n13659) );
  NANDN U10020 ( .A(y[1267]), .B(x[1267]), .Z(n13658) );
  NANDN U10021 ( .A(x[1265]), .B(y[1265]), .Z(n17295) );
  NANDN U10022 ( .A(x[1266]), .B(y[1266]), .Z(n17303) );
  NAND U10023 ( .A(n17295), .B(n17303), .Z(n24427) );
  NANDN U10024 ( .A(y[1264]), .B(x[1264]), .Z(n13661) );
  ANDN U10025 ( .B(x[1265]), .A(y[1265]), .Z(n17299) );
  ANDN U10026 ( .B(n13661), .A(n17299), .Z(n26488) );
  NANDN U10027 ( .A(y[1262]), .B(x[1262]), .Z(n17286) );
  NANDN U10028 ( .A(y[1263]), .B(x[1263]), .Z(n13660) );
  AND U10029 ( .A(n17286), .B(n13660), .Z(n26486) );
  NANDN U10030 ( .A(y[1260]), .B(x[1260]), .Z(n17282) );
  NANDN U10031 ( .A(y[1261]), .B(x[1261]), .Z(n24430) );
  AND U10032 ( .A(n17282), .B(n24430), .Z(n26485) );
  NANDN U10033 ( .A(x[1259]), .B(y[1259]), .Z(n26484) );
  NANDN U10034 ( .A(y[1258]), .B(x[1258]), .Z(n17277) );
  NANDN U10035 ( .A(y[1259]), .B(x[1259]), .Z(n17281) );
  NAND U10036 ( .A(n17277), .B(n17281), .Z(n26483) );
  ANDN U10037 ( .B(y[1258]), .A(x[1258]), .Z(n26482) );
  NANDN U10038 ( .A(y[1255]), .B(x[1255]), .Z(n13668) );
  NANDN U10039 ( .A(x[1253]), .B(y[1253]), .Z(n4517) );
  NANDN U10040 ( .A(x[1254]), .B(y[1254]), .Z(n4516) );
  NAND U10041 ( .A(n4517), .B(n4516), .Z(n7175) );
  NANDN U10042 ( .A(y[1252]), .B(x[1252]), .Z(n4519) );
  NANDN U10043 ( .A(y[1253]), .B(x[1253]), .Z(n4518) );
  AND U10044 ( .A(n4519), .B(n4518), .Z(n4520) );
  OR U10045 ( .A(n7175), .B(n4520), .Z(n4522) );
  NANDN U10046 ( .A(y[1254]), .B(x[1254]), .Z(n4521) );
  AND U10047 ( .A(n4522), .B(n4521), .Z(n24434) );
  AND U10048 ( .A(n13668), .B(n24434), .Z(n7181) );
  NANDN U10049 ( .A(y[1250]), .B(x[1250]), .Z(n4524) );
  NANDN U10050 ( .A(y[1249]), .B(x[1249]), .Z(n4523) );
  AND U10051 ( .A(n4524), .B(n4523), .Z(n4526) );
  NANDN U10052 ( .A(y[1251]), .B(x[1251]), .Z(n4525) );
  AND U10053 ( .A(n4526), .B(n4525), .Z(n17270) );
  ANDN U10054 ( .B(y[1249]), .A(x[1249]), .Z(n7166) );
  NANDN U10055 ( .A(y[1248]), .B(x[1248]), .Z(n17266) );
  OR U10056 ( .A(n7166), .B(n17266), .Z(n4527) );
  AND U10057 ( .A(n17270), .B(n4527), .Z(n26477) );
  NANDN U10058 ( .A(y[1246]), .B(x[1246]), .Z(n26473) );
  NANDN U10059 ( .A(y[1247]), .B(x[1247]), .Z(n26475) );
  AND U10060 ( .A(n26473), .B(n26475), .Z(n7165) );
  NANDN U10061 ( .A(y[1244]), .B(x[1244]), .Z(n17255) );
  NANDN U10062 ( .A(y[1245]), .B(x[1245]), .Z(n13669) );
  NAND U10063 ( .A(n17255), .B(n13669), .Z(n26471) );
  ANDN U10064 ( .B(y[1244]), .A(x[1244]), .Z(n26470) );
  ANDN U10065 ( .B(x[1242]), .A(y[1242]), .Z(n17249) );
  NANDN U10066 ( .A(x[1239]), .B(y[1239]), .Z(n13673) );
  NANDN U10067 ( .A(x[1240]), .B(y[1240]), .Z(n13672) );
  AND U10068 ( .A(n13673), .B(n13672), .Z(n7153) );
  ANDN U10069 ( .B(x[1238]), .A(y[1238]), .Z(n13675) );
  NANDN U10070 ( .A(x[1238]), .B(y[1238]), .Z(n13674) );
  NANDN U10071 ( .A(x[1237]), .B(y[1237]), .Z(n13677) );
  AND U10072 ( .A(n13674), .B(n13677), .Z(n7149) );
  NANDN U10073 ( .A(y[1236]), .B(x[1236]), .Z(n13680) );
  NANDN U10074 ( .A(x[1236]), .B(y[1236]), .Z(n13678) );
  ANDN U10075 ( .B(x[1234]), .A(y[1234]), .Z(n26457) );
  NANDN U10076 ( .A(x[1233]), .B(y[1233]), .Z(n17233) );
  NANDN U10077 ( .A(x[1234]), .B(y[1234]), .Z(n13681) );
  AND U10078 ( .A(n17233), .B(n13681), .Z(n26456) );
  ANDN U10079 ( .B(x[1233]), .A(y[1233]), .Z(n17236) );
  NANDN U10080 ( .A(y[1232]), .B(x[1232]), .Z(n4528) );
  NANDN U10081 ( .A(n17236), .B(n4528), .Z(n26455) );
  NANDN U10082 ( .A(x[1231]), .B(y[1231]), .Z(n26454) );
  ANDN U10083 ( .B(x[1231]), .A(y[1231]), .Z(n13683) );
  NANDN U10084 ( .A(y[1230]), .B(x[1230]), .Z(n17224) );
  NANDN U10085 ( .A(n13683), .B(n17224), .Z(n26452) );
  ANDN U10086 ( .B(y[1229]), .A(x[1229]), .Z(n17219) );
  ANDN U10087 ( .B(y[1230]), .A(x[1230]), .Z(n17228) );
  NOR U10088 ( .A(n17219), .B(n17228), .Z(n26451) );
  NANDN U10089 ( .A(x[1227]), .B(y[1227]), .Z(n4530) );
  NANDN U10090 ( .A(x[1226]), .B(y[1226]), .Z(n4529) );
  NAND U10091 ( .A(n4530), .B(n4529), .Z(n17213) );
  NANDN U10092 ( .A(y[1227]), .B(x[1227]), .Z(n17217) );
  NAND U10093 ( .A(n17213), .B(n17217), .Z(n4531) );
  ANDN U10094 ( .B(y[1228]), .A(x[1228]), .Z(n17222) );
  ANDN U10095 ( .B(n4531), .A(n17222), .Z(n26450) );
  NANDN U10096 ( .A(y[1225]), .B(x[1225]), .Z(n4533) );
  NANDN U10097 ( .A(y[1226]), .B(x[1226]), .Z(n4532) );
  AND U10098 ( .A(n4533), .B(n4532), .Z(n17212) );
  NANDN U10099 ( .A(y[1224]), .B(x[1224]), .Z(n13684) );
  NANDN U10100 ( .A(x[1225]), .B(y[1225]), .Z(n7130) );
  NANDN U10101 ( .A(n13684), .B(n7130), .Z(n4534) );
  AND U10102 ( .A(n4534), .B(n17217), .Z(n4535) );
  NAND U10103 ( .A(n17212), .B(n4535), .Z(n26449) );
  NANDN U10104 ( .A(x[1223]), .B(y[1223]), .Z(n13686) );
  NANDN U10105 ( .A(y[1222]), .B(x[1222]), .Z(n26443) );
  NANDN U10106 ( .A(y[1223]), .B(x[1223]), .Z(n26447) );
  NAND U10107 ( .A(n26443), .B(n26447), .Z(n7128) );
  NANDN U10108 ( .A(y[1220]), .B(x[1220]), .Z(n13688) );
  NANDN U10109 ( .A(y[1221]), .B(x[1221]), .Z(n13687) );
  AND U10110 ( .A(n13688), .B(n13687), .Z(n26440) );
  ANDN U10111 ( .B(y[1219]), .A(x[1219]), .Z(n13689) );
  NANDN U10112 ( .A(y[1219]), .B(x[1219]), .Z(n26436) );
  ANDN U10113 ( .B(x[1218]), .A(y[1218]), .Z(n26432) );
  ANDN U10114 ( .B(n26436), .A(n26432), .Z(n7121) );
  NANDN U10115 ( .A(x[1217]), .B(y[1217]), .Z(n26430) );
  NANDN U10116 ( .A(y[1216]), .B(x[1216]), .Z(n4537) );
  NANDN U10117 ( .A(y[1217]), .B(x[1217]), .Z(n4536) );
  AND U10118 ( .A(n4537), .B(n4536), .Z(n17196) );
  NANDN U10119 ( .A(x[1215]), .B(y[1215]), .Z(n4539) );
  NANDN U10120 ( .A(x[1216]), .B(y[1216]), .Z(n4538) );
  NAND U10121 ( .A(n4539), .B(n4538), .Z(n17194) );
  NANDN U10122 ( .A(y[1215]), .B(x[1215]), .Z(n4541) );
  NANDN U10123 ( .A(y[1214]), .B(x[1214]), .Z(n4540) );
  AND U10124 ( .A(n4541), .B(n4540), .Z(n17192) );
  NANDN U10125 ( .A(x[1214]), .B(y[1214]), .Z(n17191) );
  NANDN U10126 ( .A(x[1213]), .B(y[1213]), .Z(n4542) );
  AND U10127 ( .A(n17191), .B(n4542), .Z(n26422) );
  ANDN U10128 ( .B(x[1212]), .A(y[1212]), .Z(n17180) );
  NANDN U10129 ( .A(y[1213]), .B(x[1213]), .Z(n17189) );
  NANDN U10130 ( .A(n17180), .B(n17189), .Z(n26420) );
  NANDN U10131 ( .A(x[1211]), .B(y[1211]), .Z(n17177) );
  NANDN U10132 ( .A(x[1212]), .B(y[1212]), .Z(n17184) );
  AND U10133 ( .A(n17177), .B(n17184), .Z(n26418) );
  ANDN U10134 ( .B(x[1210]), .A(y[1210]), .Z(n17173) );
  ANDN U10135 ( .B(x[1211]), .A(y[1211]), .Z(n17183) );
  OR U10136 ( .A(n17173), .B(n17183), .Z(n26416) );
  NANDN U10137 ( .A(x[1209]), .B(y[1209]), .Z(n17169) );
  NANDN U10138 ( .A(x[1210]), .B(y[1210]), .Z(n17178) );
  AND U10139 ( .A(n17169), .B(n17178), .Z(n26414) );
  ANDN U10140 ( .B(x[1208]), .A(y[1208]), .Z(n13691) );
  ANDN U10141 ( .B(x[1209]), .A(y[1209]), .Z(n17175) );
  OR U10142 ( .A(n13691), .B(n17175), .Z(n26412) );
  NANDN U10143 ( .A(x[1207]), .B(y[1207]), .Z(n17164) );
  ANDN U10144 ( .B(x[1206]), .A(y[1206]), .Z(n7106) );
  ANDN U10145 ( .B(x[1207]), .A(y[1207]), .Z(n26408) );
  NANDN U10146 ( .A(x[1205]), .B(y[1205]), .Z(n13695) );
  XNOR U10147 ( .A(x[1206]), .B(y[1206]), .Z(n13693) );
  NANDN U10148 ( .A(y[1205]), .B(x[1205]), .Z(n13692) );
  ANDN U10149 ( .B(x[1204]), .A(y[1204]), .Z(n13696) );
  ANDN U10150 ( .B(n13692), .A(n13696), .Z(n7101) );
  ANDN U10151 ( .B(y[1203]), .A(x[1203]), .Z(n17157) );
  NANDN U10152 ( .A(y[1203]), .B(x[1203]), .Z(n13697) );
  NANDN U10153 ( .A(x[1201]), .B(y[1201]), .Z(n17152) );
  NANDN U10154 ( .A(x[1202]), .B(y[1202]), .Z(n17158) );
  NAND U10155 ( .A(n17152), .B(n17158), .Z(n24438) );
  ANDN U10156 ( .B(x[1200]), .A(y[1200]), .Z(n17148) );
  ANDN U10157 ( .B(x[1201]), .A(y[1201]), .Z(n17154) );
  NOR U10158 ( .A(n17148), .B(n17154), .Z(n26399) );
  ANDN U10159 ( .B(y[1200]), .A(x[1200]), .Z(n13699) );
  NANDN U10160 ( .A(y[1198]), .B(x[1198]), .Z(n17144) );
  NANDN U10161 ( .A(y[1199]), .B(x[1199]), .Z(n24439) );
  AND U10162 ( .A(n17144), .B(n24439), .Z(n26398) );
  ANDN U10163 ( .B(y[1198]), .A(x[1198]), .Z(n13701) );
  NANDN U10164 ( .A(y[1196]), .B(x[1196]), .Z(n17139) );
  NANDN U10165 ( .A(y[1197]), .B(x[1197]), .Z(n17143) );
  AND U10166 ( .A(n17139), .B(n17143), .Z(n24442) );
  NANDN U10167 ( .A(x[1195]), .B(y[1195]), .Z(n4544) );
  NANDN U10168 ( .A(x[1194]), .B(y[1194]), .Z(n4543) );
  NAND U10169 ( .A(n4544), .B(n4543), .Z(n26394) );
  NANDN U10170 ( .A(x[1193]), .B(y[1193]), .Z(n4552) );
  XNOR U10171 ( .A(x[1193]), .B(y[1193]), .Z(n4546) );
  NANDN U10172 ( .A(y[1192]), .B(x[1192]), .Z(n4545) );
  NAND U10173 ( .A(n4546), .B(n4545), .Z(n4547) );
  NAND U10174 ( .A(n4552), .B(n4547), .Z(n4549) );
  NANDN U10175 ( .A(y[1194]), .B(x[1194]), .Z(n4548) );
  AND U10176 ( .A(n4549), .B(n4548), .Z(n24444) );
  NANDN U10177 ( .A(x[1192]), .B(y[1192]), .Z(n4551) );
  NANDN U10178 ( .A(x[1191]), .B(y[1191]), .Z(n4550) );
  AND U10179 ( .A(n4551), .B(n4550), .Z(n4553) );
  NAND U10180 ( .A(n4553), .B(n4552), .Z(n13706) );
  NANDN U10181 ( .A(y[1190]), .B(x[1190]), .Z(n4554) );
  ANDN U10182 ( .B(x[1191]), .A(y[1191]), .Z(n13705) );
  ANDN U10183 ( .B(n4554), .A(n13705), .Z(n26390) );
  NANDN U10184 ( .A(x[1189]), .B(y[1189]), .Z(n13707) );
  NANDN U10185 ( .A(y[1188]), .B(x[1188]), .Z(n17128) );
  NANDN U10186 ( .A(y[1189]), .B(x[1189]), .Z(n17133) );
  NAND U10187 ( .A(n17128), .B(n17133), .Z(n26388) );
  NANDN U10188 ( .A(x[1187]), .B(y[1187]), .Z(n17126) );
  ANDN U10189 ( .B(y[1188]), .A(x[1188]), .Z(n17131) );
  ANDN U10190 ( .B(n17126), .A(n17131), .Z(n26387) );
  NANDN U10191 ( .A(y[1187]), .B(x[1187]), .Z(n4556) );
  NANDN U10192 ( .A(y[1186]), .B(x[1186]), .Z(n4555) );
  AND U10193 ( .A(n4556), .B(n4555), .Z(n13708) );
  NANDN U10194 ( .A(x[1185]), .B(y[1185]), .Z(n4558) );
  NANDN U10195 ( .A(x[1186]), .B(y[1186]), .Z(n4557) );
  NAND U10196 ( .A(n4558), .B(n4557), .Z(n13711) );
  NANDN U10197 ( .A(y[1184]), .B(x[1184]), .Z(n4559) );
  NANDN U10198 ( .A(y[1185]), .B(x[1185]), .Z(n13709) );
  AND U10199 ( .A(n4559), .B(n13709), .Z(n26384) );
  NANDN U10200 ( .A(x[1183]), .B(y[1183]), .Z(n26383) );
  ANDN U10201 ( .B(x[1182]), .A(y[1182]), .Z(n17113) );
  ANDN U10202 ( .B(x[1183]), .A(y[1183]), .Z(n17121) );
  NOR U10203 ( .A(n17113), .B(n17121), .Z(n26382) );
  NANDN U10204 ( .A(x[1181]), .B(y[1181]), .Z(n17110) );
  NANDN U10205 ( .A(x[1182]), .B(y[1182]), .Z(n17118) );
  NAND U10206 ( .A(n17110), .B(n17118), .Z(n26381) );
  ANDN U10207 ( .B(x[1180]), .A(y[1180]), .Z(n17106) );
  ANDN U10208 ( .B(x[1181]), .A(y[1181]), .Z(n17116) );
  NOR U10209 ( .A(n17106), .B(n17116), .Z(n26380) );
  NANDN U10210 ( .A(x[1180]), .B(y[1180]), .Z(n17111) );
  NANDN U10211 ( .A(x[1178]), .B(y[1178]), .Z(n4561) );
  NANDN U10212 ( .A(x[1179]), .B(y[1179]), .Z(n4560) );
  AND U10213 ( .A(n4561), .B(n4560), .Z(n17104) );
  NANDN U10214 ( .A(y[1179]), .B(x[1179]), .Z(n4563) );
  IV U10215 ( .A(n4563), .Z(n17107) );
  OR U10216 ( .A(n17104), .B(n17107), .Z(n4562) );
  NAND U10217 ( .A(n17111), .B(n4562), .Z(n24445) );
  NANDN U10218 ( .A(y[1178]), .B(x[1178]), .Z(n17102) );
  AND U10219 ( .A(n17102), .B(n4563), .Z(n4566) );
  NANDN U10220 ( .A(y[1177]), .B(x[1177]), .Z(n13712) );
  NANDN U10221 ( .A(y[1176]), .B(x[1176]), .Z(n4564) );
  AND U10222 ( .A(n13712), .B(n4564), .Z(n13713) );
  ANDN U10223 ( .B(y[1177]), .A(x[1177]), .Z(n7064) );
  OR U10224 ( .A(n13713), .B(n7064), .Z(n4565) );
  AND U10225 ( .A(n4566), .B(n4565), .Z(n26379) );
  ANDN U10226 ( .B(y[1175]), .A(x[1175]), .Z(n13714) );
  NANDN U10227 ( .A(x[1173]), .B(y[1173]), .Z(n13718) );
  NANDN U10228 ( .A(y[1173]), .B(x[1173]), .Z(n13717) );
  NANDN U10229 ( .A(x[1172]), .B(y[1172]), .Z(n13719) );
  ANDN U10230 ( .B(y[1171]), .A(x[1171]), .Z(n13722) );
  ANDN U10231 ( .B(n13719), .A(n13722), .Z(n7057) );
  ANDN U10232 ( .B(x[1170]), .A(y[1170]), .Z(n13724) );
  NANDN U10233 ( .A(x[1170]), .B(y[1170]), .Z(n13723) );
  ANDN U10234 ( .B(x[1168]), .A(y[1168]), .Z(n13728) );
  NANDN U10235 ( .A(y[1167]), .B(x[1167]), .Z(n4568) );
  NANDN U10236 ( .A(y[1166]), .B(x[1166]), .Z(n4567) );
  NAND U10237 ( .A(n4568), .B(n4567), .Z(n17085) );
  NANDN U10238 ( .A(x[1166]), .B(y[1166]), .Z(n4570) );
  NANDN U10239 ( .A(x[1165]), .B(y[1165]), .Z(n4569) );
  AND U10240 ( .A(n4570), .B(n4569), .Z(n13732) );
  NANDN U10241 ( .A(y[1165]), .B(x[1165]), .Z(n13729) );
  NANDN U10242 ( .A(y[1164]), .B(x[1164]), .Z(n4571) );
  NAND U10243 ( .A(n13729), .B(n4571), .Z(n26365) );
  ANDN U10244 ( .B(x[1162]), .A(y[1162]), .Z(n17074) );
  ANDN U10245 ( .B(x[1163]), .A(y[1163]), .Z(n17082) );
  NOR U10246 ( .A(n17074), .B(n17082), .Z(n26363) );
  ANDN U10247 ( .B(x[1160]), .A(y[1160]), .Z(n17068) );
  ANDN U10248 ( .B(x[1161]), .A(y[1161]), .Z(n17077) );
  NOR U10249 ( .A(n17068), .B(n17077), .Z(n26361) );
  ANDN U10250 ( .B(y[1160]), .A(x[1160]), .Z(n13733) );
  NANDN U10251 ( .A(y[1158]), .B(x[1158]), .Z(n26355) );
  ANDN U10252 ( .B(y[1158]), .A(x[1158]), .Z(n13735) );
  NANDN U10253 ( .A(y[1157]), .B(x[1157]), .Z(n17063) );
  NANDN U10254 ( .A(y[1156]), .B(x[1156]), .Z(n13736) );
  NANDN U10255 ( .A(x[1157]), .B(y[1157]), .Z(n4572) );
  NANDN U10256 ( .A(x[1156]), .B(y[1156]), .Z(n4573) );
  AND U10257 ( .A(n4573), .B(n4572), .Z(n17062) );
  ANDN U10258 ( .B(y[1155]), .A(x[1155]), .Z(n17057) );
  ANDN U10259 ( .B(n17062), .A(n17057), .Z(n26353) );
  NANDN U10260 ( .A(y[1154]), .B(x[1154]), .Z(n17053) );
  NANDN U10261 ( .A(y[1155]), .B(x[1155]), .Z(n13737) );
  NAND U10262 ( .A(n17053), .B(n13737), .Z(n26352) );
  ANDN U10263 ( .B(y[1154]), .A(x[1154]), .Z(n26351) );
  ANDN U10264 ( .B(x[1152]), .A(y[1152]), .Z(n13740) );
  NANDN U10265 ( .A(x[1149]), .B(y[1149]), .Z(n17041) );
  NANDN U10266 ( .A(x[1150]), .B(y[1150]), .Z(n17049) );
  NAND U10267 ( .A(n17041), .B(n17049), .Z(n26346) );
  NANDN U10268 ( .A(y[1148]), .B(x[1148]), .Z(n17039) );
  ANDN U10269 ( .B(x[1149]), .A(y[1149]), .Z(n17045) );
  ANDN U10270 ( .B(n17039), .A(n17045), .Z(n26345) );
  NANDN U10271 ( .A(y[1145]), .B(x[1145]), .Z(n13746) );
  NANDN U10272 ( .A(y[1144]), .B(x[1144]), .Z(n4574) );
  AND U10273 ( .A(n13746), .B(n4574), .Z(n13748) );
  NANDN U10274 ( .A(x[1143]), .B(y[1143]), .Z(n17030) );
  ANDN U10275 ( .B(x[1143]), .A(y[1143]), .Z(n13747) );
  ANDN U10276 ( .B(x[1142]), .A(y[1142]), .Z(n4575) );
  NOR U10277 ( .A(n13747), .B(n4575), .Z(n7013) );
  NANDN U10278 ( .A(x[1141]), .B(y[1141]), .Z(n13750) );
  NANDN U10279 ( .A(y[1141]), .B(x[1141]), .Z(n17027) );
  NANDN U10280 ( .A(x[1139]), .B(y[1139]), .Z(n13754) );
  NANDN U10281 ( .A(y[1138]), .B(x[1138]), .Z(n13756) );
  NANDN U10282 ( .A(x[1137]), .B(y[1137]), .Z(n7001) );
  NANDN U10283 ( .A(x[1136]), .B(y[1136]), .Z(n4576) );
  NAND U10284 ( .A(n7001), .B(n4576), .Z(n17021) );
  ANDN U10285 ( .B(y[1135]), .A(x[1135]), .Z(n17015) );
  NOR U10286 ( .A(n17021), .B(n17015), .Z(n26336) );
  NANDN U10287 ( .A(y[1134]), .B(x[1134]), .Z(n26334) );
  NANDN U10288 ( .A(y[1135]), .B(x[1135]), .Z(n24453) );
  NAND U10289 ( .A(n26334), .B(n24453), .Z(n6998) );
  ANDN U10290 ( .B(y[1130]), .A(x[1130]), .Z(n26329) );
  NANDN U10291 ( .A(y[1128]), .B(x[1128]), .Z(n16993) );
  ANDN U10292 ( .B(y[1127]), .A(x[1127]), .Z(n24458) );
  NANDN U10293 ( .A(y[1126]), .B(x[1126]), .Z(n26327) );
  NANDN U10294 ( .A(y[1127]), .B(x[1127]), .Z(n16994) );
  ANDN U10295 ( .B(y[1125]), .A(x[1125]), .Z(n16985) );
  ANDN U10296 ( .B(y[1126]), .A(x[1126]), .Z(n16992) );
  OR U10297 ( .A(n16985), .B(n16992), .Z(n26326) );
  NANDN U10298 ( .A(y[1124]), .B(x[1124]), .Z(n16981) );
  NANDN U10299 ( .A(y[1125]), .B(x[1125]), .Z(n13759) );
  NAND U10300 ( .A(n16981), .B(n13759), .Z(n26325) );
  NANDN U10301 ( .A(x[1124]), .B(y[1124]), .Z(n16986) );
  ANDN U10302 ( .B(x[1122]), .A(y[1122]), .Z(n13764) );
  NANDN U10303 ( .A(y[1121]), .B(x[1121]), .Z(n4578) );
  NANDN U10304 ( .A(y[1120]), .B(x[1120]), .Z(n4577) );
  NAND U10305 ( .A(n4578), .B(n4577), .Z(n13763) );
  NANDN U10306 ( .A(x[1120]), .B(y[1120]), .Z(n4580) );
  NANDN U10307 ( .A(x[1119]), .B(y[1119]), .Z(n4579) );
  AND U10308 ( .A(n4580), .B(n4579), .Z(n13765) );
  NANDN U10309 ( .A(y[1119]), .B(x[1119]), .Z(n13767) );
  NANDN U10310 ( .A(y[1118]), .B(x[1118]), .Z(n4581) );
  NAND U10311 ( .A(n13767), .B(n4581), .Z(n13769) );
  NANDN U10312 ( .A(x[1117]), .B(y[1117]), .Z(n26316) );
  NANDN U10313 ( .A(y[1116]), .B(x[1116]), .Z(n13772) );
  NANDN U10314 ( .A(y[1117]), .B(x[1117]), .Z(n13770) );
  NAND U10315 ( .A(n13772), .B(n13770), .Z(n26317) );
  NANDN U10316 ( .A(x[1115]), .B(y[1115]), .Z(n16969) );
  NANDN U10317 ( .A(y[1114]), .B(x[1114]), .Z(n26312) );
  NANDN U10318 ( .A(x[1113]), .B(y[1113]), .Z(n26311) );
  NANDN U10319 ( .A(y[1112]), .B(x[1112]), .Z(n13775) );
  NANDN U10320 ( .A(y[1113]), .B(x[1113]), .Z(n13773) );
  NAND U10321 ( .A(n13775), .B(n13773), .Z(n26310) );
  NANDN U10322 ( .A(x[1111]), .B(y[1111]), .Z(n13777) );
  NANDN U10323 ( .A(x[1110]), .B(y[1110]), .Z(n13776) );
  ANDN U10324 ( .B(x[1109]), .A(y[1109]), .Z(n13778) );
  NANDN U10325 ( .A(x[1109]), .B(y[1109]), .Z(n4583) );
  NANDN U10326 ( .A(x[1108]), .B(y[1108]), .Z(n4582) );
  AND U10327 ( .A(n4583), .B(n4582), .Z(n26306) );
  NANDN U10328 ( .A(y[1107]), .B(x[1107]), .Z(n4585) );
  ANDN U10329 ( .B(x[1108]), .A(y[1108]), .Z(n4584) );
  ANDN U10330 ( .B(n4585), .A(n4584), .Z(n4589) );
  XNOR U10331 ( .A(x[1107]), .B(y[1107]), .Z(n4587) );
  ANDN U10332 ( .B(x[1106]), .A(y[1106]), .Z(n4586) );
  NAND U10333 ( .A(n4587), .B(n4586), .Z(n4588) );
  NAND U10334 ( .A(n4589), .B(n4588), .Z(n26303) );
  NANDN U10335 ( .A(x[1106]), .B(y[1106]), .Z(n4591) );
  NANDN U10336 ( .A(x[1105]), .B(y[1105]), .Z(n4590) );
  AND U10337 ( .A(n4591), .B(n4590), .Z(n4593) );
  NANDN U10338 ( .A(x[1107]), .B(y[1107]), .Z(n4592) );
  AND U10339 ( .A(n4593), .B(n4592), .Z(n26302) );
  ANDN U10340 ( .B(y[1101]), .A(x[1101]), .Z(n4598) );
  ANDN U10341 ( .B(x[1100]), .A(y[1100]), .Z(n13785) );
  NANDN U10342 ( .A(n4598), .B(n13785), .Z(n4597) );
  NANDN U10343 ( .A(y[1102]), .B(x[1102]), .Z(n4595) );
  NANDN U10344 ( .A(y[1101]), .B(x[1101]), .Z(n4594) );
  AND U10345 ( .A(n4595), .B(n4594), .Z(n4596) );
  NANDN U10346 ( .A(y[1103]), .B(x[1103]), .Z(n6949) );
  NAND U10347 ( .A(n4596), .B(n6949), .Z(n16955) );
  ANDN U10348 ( .B(n4597), .A(n16955), .Z(n26300) );
  NANDN U10349 ( .A(x[1099]), .B(y[1099]), .Z(n4603) );
  NANDN U10350 ( .A(x[1098]), .B(y[1098]), .Z(n4599) );
  AND U10351 ( .A(n4603), .B(n4599), .Z(n13783) );
  NANDN U10352 ( .A(x[1097]), .B(y[1097]), .Z(n4600) );
  AND U10353 ( .A(n13783), .B(n4600), .Z(n4607) );
  ANDN U10354 ( .B(x[1096]), .A(y[1096]), .Z(n16947) );
  ANDN U10355 ( .B(x[1097]), .A(y[1097]), .Z(n13781) );
  OR U10356 ( .A(n16947), .B(n13781), .Z(n4601) );
  AND U10357 ( .A(n4607), .B(n4601), .Z(n4605) );
  ANDN U10358 ( .B(x[1099]), .A(y[1099]), .Z(n16949) );
  ANDN U10359 ( .B(x[1098]), .A(y[1098]), .Z(n13780) );
  OR U10360 ( .A(n16949), .B(n13780), .Z(n4602) );
  NAND U10361 ( .A(n4603), .B(n4602), .Z(n4604) );
  NANDN U10362 ( .A(n4605), .B(n4604), .Z(n26298) );
  NANDN U10363 ( .A(x[1095]), .B(y[1095]), .Z(n13787) );
  NANDN U10364 ( .A(x[1096]), .B(y[1096]), .Z(n4606) );
  AND U10365 ( .A(n4607), .B(n4606), .Z(n26297) );
  NANDN U10366 ( .A(x[1091]), .B(y[1091]), .Z(n4609) );
  NANDN U10367 ( .A(x[1092]), .B(y[1092]), .Z(n4608) );
  NAND U10368 ( .A(n4609), .B(n4608), .Z(n13791) );
  NANDN U10369 ( .A(y[1090]), .B(x[1090]), .Z(n4610) );
  NANDN U10370 ( .A(y[1091]), .B(x[1091]), .Z(n13793) );
  AND U10371 ( .A(n4610), .B(n13793), .Z(n26292) );
  NANDN U10372 ( .A(x[1089]), .B(y[1089]), .Z(n24461) );
  ANDN U10373 ( .B(x[1089]), .A(y[1089]), .Z(n16936) );
  NANDN U10374 ( .A(y[1088]), .B(x[1088]), .Z(n4611) );
  NANDN U10375 ( .A(n16936), .B(n4611), .Z(n13795) );
  NANDN U10376 ( .A(x[1087]), .B(y[1087]), .Z(n26289) );
  ANDN U10377 ( .B(x[1086]), .A(y[1086]), .Z(n16929) );
  NANDN U10378 ( .A(y[1087]), .B(x[1087]), .Z(n13796) );
  NANDN U10379 ( .A(n16929), .B(n13796), .Z(n26288) );
  NANDN U10380 ( .A(x[1085]), .B(y[1085]), .Z(n16925) );
  NANDN U10381 ( .A(x[1086]), .B(y[1086]), .Z(n13797) );
  AND U10382 ( .A(n16925), .B(n13797), .Z(n26287) );
  ANDN U10383 ( .B(x[1085]), .A(y[1085]), .Z(n16930) );
  NANDN U10384 ( .A(y[1084]), .B(x[1084]), .Z(n16923) );
  NANDN U10385 ( .A(n16930), .B(n16923), .Z(n26286) );
  NANDN U10386 ( .A(x[1084]), .B(y[1084]), .Z(n16927) );
  ANDN U10387 ( .B(y[1083]), .A(x[1083]), .Z(n16921) );
  ANDN U10388 ( .B(n16927), .A(n16921), .Z(n24463) );
  NANDN U10389 ( .A(y[1083]), .B(x[1083]), .Z(n13799) );
  NANDN U10390 ( .A(y[1082]), .B(x[1082]), .Z(n4612) );
  NAND U10391 ( .A(n13799), .B(n4612), .Z(n13800) );
  NANDN U10392 ( .A(x[1081]), .B(y[1081]), .Z(n13802) );
  NANDN U10393 ( .A(y[1081]), .B(x[1081]), .Z(n13803) );
  NANDN U10394 ( .A(y[1080]), .B(x[1080]), .Z(n4613) );
  AND U10395 ( .A(n13803), .B(n4613), .Z(n6933) );
  NANDN U10396 ( .A(x[1080]), .B(y[1080]), .Z(n13801) );
  NANDN U10397 ( .A(x[1079]), .B(y[1079]), .Z(n13804) );
  NAND U10398 ( .A(n13801), .B(n13804), .Z(n4614) );
  NAND U10399 ( .A(n6933), .B(n4614), .Z(n4615) );
  NANDN U10400 ( .A(x[1082]), .B(y[1082]), .Z(n13798) );
  AND U10401 ( .A(n4615), .B(n13798), .Z(n6936) );
  NANDN U10402 ( .A(y[1078]), .B(x[1078]), .Z(n13806) );
  NANDN U10403 ( .A(x[1078]), .B(y[1078]), .Z(n13805) );
  NANDN U10404 ( .A(y[1077]), .B(x[1077]), .Z(n13807) );
  ANDN U10405 ( .B(x[1076]), .A(y[1076]), .Z(n13810) );
  ANDN U10406 ( .B(n13807), .A(n13810), .Z(n6928) );
  ANDN U10407 ( .B(y[1075]), .A(x[1075]), .Z(n13812) );
  NANDN U10408 ( .A(y[1075]), .B(x[1075]), .Z(n13811) );
  NANDN U10409 ( .A(x[1073]), .B(y[1073]), .Z(n16902) );
  NANDN U10410 ( .A(x[1074]), .B(y[1074]), .Z(n16910) );
  NAND U10411 ( .A(n16902), .B(n16910), .Z(n24466) );
  ANDN U10412 ( .B(x[1072]), .A(y[1072]), .Z(n16900) );
  ANDN U10413 ( .B(x[1073]), .A(y[1073]), .Z(n16906) );
  NOR U10414 ( .A(n16900), .B(n16906), .Z(n26277) );
  NANDN U10415 ( .A(x[1069]), .B(y[1069]), .Z(n4617) );
  NANDN U10416 ( .A(x[1070]), .B(y[1070]), .Z(n4616) );
  NAND U10417 ( .A(n4617), .B(n4616), .Z(n13815) );
  NANDN U10418 ( .A(y[1069]), .B(x[1069]), .Z(n13813) );
  NANDN U10419 ( .A(y[1068]), .B(x[1068]), .Z(n4618) );
  AND U10420 ( .A(n13813), .B(n4618), .Z(n26272) );
  ANDN U10421 ( .B(y[1067]), .A(x[1067]), .Z(n24468) );
  NANDN U10422 ( .A(y[1066]), .B(x[1066]), .Z(n16890) );
  NANDN U10423 ( .A(y[1067]), .B(x[1067]), .Z(n16892) );
  AND U10424 ( .A(n16890), .B(n16892), .Z(n24469) );
  NANDN U10425 ( .A(x[1065]), .B(y[1065]), .Z(n4620) );
  NANDN U10426 ( .A(x[1066]), .B(y[1066]), .Z(n4619) );
  NAND U10427 ( .A(n4620), .B(n4619), .Z(n13818) );
  NANDN U10428 ( .A(y[1064]), .B(x[1064]), .Z(n4621) );
  NANDN U10429 ( .A(y[1065]), .B(x[1065]), .Z(n13816) );
  AND U10430 ( .A(n4621), .B(n13816), .Z(n26270) );
  ANDN U10431 ( .B(y[1063]), .A(x[1063]), .Z(n13819) );
  ANDN U10432 ( .B(x[1062]), .A(y[1062]), .Z(n16879) );
  ANDN U10433 ( .B(x[1063]), .A(y[1063]), .Z(n16887) );
  NOR U10434 ( .A(n16879), .B(n16887), .Z(n26268) );
  NANDN U10435 ( .A(x[1061]), .B(y[1061]), .Z(n16875) );
  NANDN U10436 ( .A(x[1062]), .B(y[1062]), .Z(n16883) );
  NAND U10437 ( .A(n16875), .B(n16883), .Z(n26267) );
  ANDN U10438 ( .B(x[1060]), .A(y[1060]), .Z(n16874) );
  ANDN U10439 ( .B(x[1061]), .A(y[1061]), .Z(n16881) );
  NOR U10440 ( .A(n16874), .B(n16881), .Z(n26266) );
  NANDN U10441 ( .A(x[1060]), .B(y[1060]), .Z(n26265) );
  ANDN U10442 ( .B(x[1058]), .A(y[1058]), .Z(n26262) );
  ANDN U10443 ( .B(x[1059]), .A(y[1059]), .Z(n26264) );
  NOR U10444 ( .A(n26262), .B(n26264), .Z(n6902) );
  ANDN U10445 ( .B(y[1057]), .A(x[1057]), .Z(n13822) );
  ANDN U10446 ( .B(x[1056]), .A(y[1056]), .Z(n16861) );
  ANDN U10447 ( .B(x[1057]), .A(y[1057]), .Z(n16870) );
  NOR U10448 ( .A(n16861), .B(n16870), .Z(n26260) );
  NANDN U10449 ( .A(y[1054]), .B(x[1054]), .Z(n13825) );
  ANDN U10450 ( .B(x[1055]), .A(y[1055]), .Z(n16862) );
  ANDN U10451 ( .B(n13825), .A(n16862), .Z(n26258) );
  ANDN U10452 ( .B(y[1053]), .A(x[1053]), .Z(n16855) );
  NANDN U10453 ( .A(x[1054]), .B(y[1054]), .Z(n13824) );
  NANDN U10454 ( .A(n16855), .B(n13824), .Z(n26257) );
  NANDN U10455 ( .A(y[1052]), .B(x[1052]), .Z(n16851) );
  NANDN U10456 ( .A(y[1053]), .B(x[1053]), .Z(n13826) );
  NAND U10457 ( .A(n16851), .B(n13826), .Z(n26256) );
  ANDN U10458 ( .B(y[1052]), .A(x[1052]), .Z(n26255) );
  NANDN U10459 ( .A(y[1050]), .B(x[1050]), .Z(n26253) );
  NANDN U10460 ( .A(y[1051]), .B(x[1051]), .Z(n24471) );
  NAND U10461 ( .A(n26253), .B(n24471), .Z(n6891) );
  ANDN U10462 ( .B(y[1048]), .A(x[1048]), .Z(n26250) );
  NANDN U10463 ( .A(y[1046]), .B(x[1046]), .Z(n13832) );
  ANDN U10464 ( .B(y[1045]), .A(x[1045]), .Z(n13834) );
  NANDN U10465 ( .A(y[1044]), .B(x[1044]), .Z(n13836) );
  ANDN U10466 ( .B(y[1043]), .A(x[1043]), .Z(n13838) );
  NANDN U10467 ( .A(y[1043]), .B(x[1043]), .Z(n13837) );
  NANDN U10468 ( .A(y[1037]), .B(x[1037]), .Z(n4623) );
  NANDN U10469 ( .A(y[1036]), .B(x[1036]), .Z(n4622) );
  AND U10470 ( .A(n4623), .B(n4622), .Z(n26240) );
  NANDN U10471 ( .A(x[1035]), .B(y[1035]), .Z(n4625) );
  ANDN U10472 ( .B(y[1036]), .A(x[1036]), .Z(n4624) );
  ANDN U10473 ( .B(n4625), .A(n4624), .Z(n4629) );
  XNOR U10474 ( .A(y[1035]), .B(x[1035]), .Z(n4627) );
  ANDN U10475 ( .B(y[1034]), .A(x[1034]), .Z(n4626) );
  NAND U10476 ( .A(n4627), .B(n4626), .Z(n4628) );
  NAND U10477 ( .A(n4629), .B(n4628), .Z(n26239) );
  NANDN U10478 ( .A(y[1034]), .B(x[1034]), .Z(n4631) );
  NANDN U10479 ( .A(y[1033]), .B(x[1033]), .Z(n4630) );
  AND U10480 ( .A(n4631), .B(n4630), .Z(n4633) );
  NANDN U10481 ( .A(y[1035]), .B(x[1035]), .Z(n4632) );
  AND U10482 ( .A(n4633), .B(n4632), .Z(n26238) );
  NANDN U10483 ( .A(x[1032]), .B(y[1032]), .Z(n4635) );
  NANDN U10484 ( .A(x[1033]), .B(y[1033]), .Z(n4634) );
  NAND U10485 ( .A(n4635), .B(n4634), .Z(n26237) );
  NANDN U10486 ( .A(y[1032]), .B(x[1032]), .Z(n4637) );
  NANDN U10487 ( .A(y[1031]), .B(x[1031]), .Z(n4636) );
  AND U10488 ( .A(n4637), .B(n4636), .Z(n16828) );
  NANDN U10489 ( .A(y[1030]), .B(x[1030]), .Z(n16823) );
  NANDN U10490 ( .A(x[1031]), .B(y[1031]), .Z(n6850) );
  NANDN U10491 ( .A(y[1029]), .B(x[1029]), .Z(n16822) );
  NANDN U10492 ( .A(y[1028]), .B(x[1028]), .Z(n16817) );
  NANDN U10493 ( .A(x[1029]), .B(y[1029]), .Z(n4638) );
  ANDN U10494 ( .B(y[1027]), .A(x[1027]), .Z(n16812) );
  NANDN U10495 ( .A(x[1028]), .B(y[1028]), .Z(n4639) );
  AND U10496 ( .A(n4639), .B(n4638), .Z(n16821) );
  NANDN U10497 ( .A(n16812), .B(n16821), .Z(n26233) );
  NANDN U10498 ( .A(y[1026]), .B(x[1026]), .Z(n16809) );
  NANDN U10499 ( .A(y[1027]), .B(x[1027]), .Z(n16816) );
  AND U10500 ( .A(n16809), .B(n16816), .Z(n26232) );
  ANDN U10501 ( .B(y[1026]), .A(x[1026]), .Z(n16815) );
  NANDN U10502 ( .A(x[1024]), .B(y[1024]), .Z(n4641) );
  NANDN U10503 ( .A(x[1025]), .B(y[1025]), .Z(n4640) );
  NAND U10504 ( .A(n4641), .B(n4640), .Z(n16807) );
  NANDN U10505 ( .A(y[1025]), .B(x[1025]), .Z(n16810) );
  NAND U10506 ( .A(n16807), .B(n16810), .Z(n4642) );
  NANDN U10507 ( .A(n16815), .B(n4642), .Z(n26229) );
  NANDN U10508 ( .A(y[1024]), .B(x[1024]), .Z(n4644) );
  NANDN U10509 ( .A(y[1023]), .B(x[1023]), .Z(n4643) );
  AND U10510 ( .A(n4644), .B(n4643), .Z(n16805) );
  NANDN U10511 ( .A(y[1022]), .B(x[1022]), .Z(n16800) );
  NANDN U10512 ( .A(x[1023]), .B(y[1023]), .Z(n4645) );
  NANDN U10513 ( .A(x[1021]), .B(y[1021]), .Z(n13843) );
  NANDN U10514 ( .A(x[1022]), .B(y[1022]), .Z(n4646) );
  AND U10515 ( .A(n4646), .B(n4645), .Z(n26227) );
  ANDN U10516 ( .B(x[1020]), .A(y[1020]), .Z(n13844) );
  NANDN U10517 ( .A(y[1021]), .B(x[1021]), .Z(n26226) );
  ANDN U10518 ( .B(y[1019]), .A(x[1019]), .Z(n13846) );
  NANDN U10519 ( .A(y[1019]), .B(x[1019]), .Z(n13845) );
  NANDN U10520 ( .A(x[1018]), .B(y[1018]), .Z(n4648) );
  NANDN U10521 ( .A(x[1017]), .B(y[1017]), .Z(n4647) );
  NAND U10522 ( .A(n4648), .B(n4647), .Z(n13847) );
  NANDN U10523 ( .A(y[1016]), .B(x[1016]), .Z(n4649) );
  NANDN U10524 ( .A(y[1017]), .B(x[1017]), .Z(n13849) );
  AND U10525 ( .A(n4649), .B(n13849), .Z(n13851) );
  ANDN U10526 ( .B(y[1016]), .A(x[1016]), .Z(n13848) );
  NANDN U10527 ( .A(x[1015]), .B(y[1015]), .Z(n16793) );
  ANDN U10528 ( .B(x[1014]), .A(y[1014]), .Z(n13853) );
  NANDN U10529 ( .A(x[1014]), .B(y[1014]), .Z(n16794) );
  NANDN U10530 ( .A(y[1012]), .B(x[1012]), .Z(n26220) );
  NANDN U10531 ( .A(x[1010]), .B(y[1010]), .Z(n26219) );
  ANDN U10532 ( .B(y[1009]), .A(x[1009]), .Z(n26218) );
  ANDN U10533 ( .B(n26219), .A(n26218), .Z(n6823) );
  NANDN U10534 ( .A(y[1008]), .B(x[1008]), .Z(n16779) );
  NANDN U10535 ( .A(y[1009]), .B(x[1009]), .Z(n13857) );
  NAND U10536 ( .A(n16779), .B(n13857), .Z(n26217) );
  NANDN U10537 ( .A(x[1007]), .B(y[1007]), .Z(n13860) );
  ANDN U10538 ( .B(y[1008]), .A(x[1008]), .Z(n26215) );
  ANDN U10539 ( .B(n13860), .A(n26215), .Z(n6820) );
  ANDN U10540 ( .B(x[1006]), .A(y[1006]), .Z(n13861) );
  NANDN U10541 ( .A(y[1007]), .B(x[1007]), .Z(n26214) );
  NANDN U10542 ( .A(x[1005]), .B(y[1005]), .Z(n13863) );
  NANDN U10543 ( .A(y[1005]), .B(x[1005]), .Z(n13862) );
  NANDN U10544 ( .A(x[1004]), .B(y[1004]), .Z(n13864) );
  ANDN U10545 ( .B(y[1003]), .A(x[1003]), .Z(n13867) );
  ANDN U10546 ( .B(n13864), .A(n13867), .Z(n6812) );
  ANDN U10547 ( .B(x[1002]), .A(y[1002]), .Z(n16771) );
  NANDN U10548 ( .A(x[1002]), .B(y[1002]), .Z(n13868) );
  ANDN U10549 ( .B(x[1000]), .A(y[1000]), .Z(n24480) );
  ANDN U10550 ( .B(x[997]), .A(y[997]), .Z(n16761) );
  NANDN U10551 ( .A(y[996]), .B(x[996]), .Z(n16750) );
  NANDN U10552 ( .A(n16761), .B(n16750), .Z(n26205) );
  NANDN U10553 ( .A(y[995]), .B(x[995]), .Z(n16751) );
  NANDN U10554 ( .A(x[993]), .B(y[993]), .Z(n4657) );
  XNOR U10555 ( .A(x[993]), .B(y[993]), .Z(n4651) );
  NANDN U10556 ( .A(y[992]), .B(x[992]), .Z(n4650) );
  NAND U10557 ( .A(n4651), .B(n4650), .Z(n4652) );
  NAND U10558 ( .A(n4657), .B(n4652), .Z(n4654) );
  NANDN U10559 ( .A(y[994]), .B(x[994]), .Z(n4653) );
  NAND U10560 ( .A(n4654), .B(n4653), .Z(n16747) );
  ANDN U10561 ( .B(n16751), .A(n16747), .Z(n26202) );
  NANDN U10562 ( .A(x[992]), .B(y[992]), .Z(n4656) );
  NANDN U10563 ( .A(x[991]), .B(y[991]), .Z(n4655) );
  AND U10564 ( .A(n4656), .B(n4655), .Z(n4658) );
  NAND U10565 ( .A(n4658), .B(n4657), .Z(n13871) );
  NANDN U10566 ( .A(y[990]), .B(x[990]), .Z(n4659) );
  NANDN U10567 ( .A(y[991]), .B(x[991]), .Z(n13869) );
  AND U10568 ( .A(n4659), .B(n13869), .Z(n26200) );
  NANDN U10569 ( .A(y[988]), .B(x[988]), .Z(n16736) );
  ANDN U10570 ( .B(x[989]), .A(y[989]), .Z(n16744) );
  ANDN U10571 ( .B(n16736), .A(n16744), .Z(n26198) );
  ANDN U10572 ( .B(y[987]), .A(x[987]), .Z(n16732) );
  NANDN U10573 ( .A(x[988]), .B(y[988]), .Z(n16740) );
  NANDN U10574 ( .A(n16732), .B(n16740), .Z(n24482) );
  ANDN U10575 ( .B(x[987]), .A(y[987]), .Z(n16738) );
  NANDN U10576 ( .A(y[986]), .B(x[986]), .Z(n16728) );
  NANDN U10577 ( .A(n16738), .B(n16728), .Z(n26197) );
  ANDN U10578 ( .B(y[985]), .A(x[985]), .Z(n16724) );
  ANDN U10579 ( .B(y[986]), .A(x[986]), .Z(n16734) );
  NOR U10580 ( .A(n16724), .B(n16734), .Z(n26196) );
  NANDN U10581 ( .A(y[984]), .B(x[984]), .Z(n16722) );
  NANDN U10582 ( .A(y[985]), .B(x[985]), .Z(n16727) );
  NAND U10583 ( .A(n16722), .B(n16727), .Z(n26195) );
  NANDN U10584 ( .A(x[983]), .B(y[983]), .Z(n13873) );
  ANDN U10585 ( .B(y[984]), .A(x[984]), .Z(n26194) );
  ANDN U10586 ( .B(n13873), .A(n26194), .Z(n6786) );
  ANDN U10587 ( .B(x[982]), .A(y[982]), .Z(n6784) );
  ANDN U10588 ( .B(y[981]), .A(x[981]), .Z(n13876) );
  NANDN U10589 ( .A(y[981]), .B(x[981]), .Z(n13875) );
  ANDN U10590 ( .B(y[980]), .A(x[980]), .Z(n13877) );
  NANDN U10591 ( .A(y[978]), .B(x[978]), .Z(n16710) );
  NANDN U10592 ( .A(x[978]), .B(y[978]), .Z(n16715) );
  NANDN U10593 ( .A(y[977]), .B(x[977]), .Z(n16711) );
  NANDN U10594 ( .A(y[976]), .B(x[976]), .Z(n16707) );
  NANDN U10595 ( .A(x[977]), .B(y[977]), .Z(n4663) );
  NANDN U10596 ( .A(y[979]), .B(x[979]), .Z(n13879) );
  NANDN U10597 ( .A(y[975]), .B(x[975]), .Z(n4667) );
  XNOR U10598 ( .A(y[975]), .B(x[975]), .Z(n4661) );
  NANDN U10599 ( .A(x[974]), .B(y[974]), .Z(n4660) );
  NAND U10600 ( .A(n4661), .B(n4660), .Z(n4662) );
  AND U10601 ( .A(n4667), .B(n4662), .Z(n16705) );
  ANDN U10602 ( .B(n16715), .A(n16705), .Z(n4665) );
  NANDN U10603 ( .A(x[976]), .B(y[976]), .Z(n4664) );
  AND U10604 ( .A(n4664), .B(n4663), .Z(n16709) );
  AND U10605 ( .A(n4665), .B(n16709), .Z(n26186) );
  NANDN U10606 ( .A(y[974]), .B(x[974]), .Z(n4666) );
  AND U10607 ( .A(n4667), .B(n4666), .Z(n16703) );
  NANDN U10608 ( .A(y[973]), .B(x[973]), .Z(n13880) );
  NANDN U10609 ( .A(y[972]), .B(x[972]), .Z(n4668) );
  AND U10610 ( .A(n13880), .B(n4668), .Z(n13881) );
  NANDN U10611 ( .A(x[973]), .B(y[973]), .Z(n4669) );
  NANDN U10612 ( .A(x[972]), .B(y[972]), .Z(n4670) );
  AND U10613 ( .A(n4670), .B(n4669), .Z(n26184) );
  NANDN U10614 ( .A(y[971]), .B(x[971]), .Z(n26183) );
  ANDN U10615 ( .B(y[969]), .A(x[969]), .Z(n13882) );
  NANDN U10616 ( .A(y[969]), .B(x[969]), .Z(n16693) );
  NANDN U10617 ( .A(x[967]), .B(y[967]), .Z(n13886) );
  ANDN U10618 ( .B(y[968]), .A(x[968]), .Z(n13883) );
  ANDN U10619 ( .B(n13886), .A(n13883), .Z(n6763) );
  NANDN U10620 ( .A(y[966]), .B(x[966]), .Z(n13889) );
  NANDN U10621 ( .A(x[966]), .B(y[966]), .Z(n13887) );
  NANDN U10622 ( .A(y[964]), .B(x[964]), .Z(n13893) );
  NANDN U10623 ( .A(x[963]), .B(y[963]), .Z(n26175) );
  ANDN U10624 ( .B(x[962]), .A(y[962]), .Z(n26174) );
  NANDN U10625 ( .A(x[962]), .B(y[962]), .Z(n16684) );
  ANDN U10626 ( .B(y[961]), .A(x[961]), .Z(n16677) );
  ANDN U10627 ( .B(n16684), .A(n16677), .Z(n26173) );
  NANDN U10628 ( .A(y[960]), .B(x[960]), .Z(n16673) );
  NANDN U10629 ( .A(y[961]), .B(x[961]), .Z(n16681) );
  NAND U10630 ( .A(n16673), .B(n16681), .Z(n26172) );
  ANDN U10631 ( .B(y[959]), .A(x[959]), .Z(n16669) );
  ANDN U10632 ( .B(y[960]), .A(x[960]), .Z(n16679) );
  NOR U10633 ( .A(n16669), .B(n16679), .Z(n26171) );
  NANDN U10634 ( .A(y[958]), .B(x[958]), .Z(n16667) );
  NANDN U10635 ( .A(y[959]), .B(x[959]), .Z(n16672) );
  NAND U10636 ( .A(n16667), .B(n16672), .Z(n26169) );
  NANDN U10637 ( .A(y[957]), .B(x[957]), .Z(n26167) );
  NANDN U10638 ( .A(x[956]), .B(y[956]), .Z(n16664) );
  ANDN U10639 ( .B(x[954]), .A(y[954]), .Z(n13898) );
  NANDN U10640 ( .A(x[953]), .B(y[953]), .Z(n13901) );
  NANDN U10641 ( .A(y[953]), .B(x[953]), .Z(n13899) );
  NANDN U10642 ( .A(y[952]), .B(x[952]), .Z(n13902) );
  NANDN U10643 ( .A(x[951]), .B(y[951]), .Z(n13904) );
  NANDN U10644 ( .A(y[951]), .B(x[951]), .Z(n13903) );
  NANDN U10645 ( .A(x[950]), .B(y[950]), .Z(n13905) );
  ANDN U10646 ( .B(y[949]), .A(x[949]), .Z(n13908) );
  ANDN U10647 ( .B(n13905), .A(n13908), .Z(n6731) );
  ANDN U10648 ( .B(x[948]), .A(y[948]), .Z(n13910) );
  NANDN U10649 ( .A(x[948]), .B(y[948]), .Z(n13909) );
  ANDN U10650 ( .B(x[946]), .A(y[946]), .Z(n13914) );
  NANDN U10651 ( .A(x[945]), .B(y[945]), .Z(n13916) );
  ANDN U10652 ( .B(x[944]), .A(y[944]), .Z(n13918) );
  NANDN U10653 ( .A(x[944]), .B(y[944]), .Z(n13917) );
  NANDN U10654 ( .A(y[942]), .B(x[942]), .Z(n16643) );
  NANDN U10655 ( .A(y[943]), .B(x[943]), .Z(n13919) );
  NAND U10656 ( .A(n16643), .B(n13919), .Z(n24486) );
  NANDN U10657 ( .A(x[942]), .B(y[942]), .Z(n13920) );
  NANDN U10658 ( .A(x[941]), .B(y[941]), .Z(n6712) );
  NANDN U10659 ( .A(y[940]), .B(x[940]), .Z(n26146) );
  NANDN U10660 ( .A(y[941]), .B(x[941]), .Z(n26148) );
  NAND U10661 ( .A(n26146), .B(n26148), .Z(n4671) );
  AND U10662 ( .A(n6712), .B(n4671), .Z(n6715) );
  NANDN U10663 ( .A(x[939]), .B(y[939]), .Z(n6708) );
  NANDN U10664 ( .A(y[938]), .B(x[938]), .Z(n13922) );
  NANDN U10665 ( .A(y[939]), .B(x[939]), .Z(n16639) );
  NAND U10666 ( .A(n13922), .B(n16639), .Z(n4672) );
  AND U10667 ( .A(n6708), .B(n4672), .Z(n26145) );
  NANDN U10668 ( .A(y[936]), .B(x[936]), .Z(n16630) );
  NANDN U10669 ( .A(y[937]), .B(x[937]), .Z(n13923) );
  AND U10670 ( .A(n16630), .B(n13923), .Z(n26143) );
  ANDN U10671 ( .B(y[936]), .A(x[936]), .Z(n26142) );
  NANDN U10672 ( .A(y[934]), .B(x[934]), .Z(n13926) );
  NANDN U10673 ( .A(x[933]), .B(y[933]), .Z(n13929) );
  NANDN U10674 ( .A(y[933]), .B(x[933]), .Z(n13927) );
  ANDN U10675 ( .B(y[931]), .A(x[931]), .Z(n26137) );
  NANDN U10676 ( .A(y[931]), .B(x[931]), .Z(n16623) );
  NANDN U10677 ( .A(y[930]), .B(x[930]), .Z(n4673) );
  AND U10678 ( .A(n16623), .B(n4673), .Z(n26136) );
  NANDN U10679 ( .A(x[925]), .B(y[925]), .Z(n13931) );
  NANDN U10680 ( .A(y[924]), .B(x[924]), .Z(n4674) );
  NANDN U10681 ( .A(y[925]), .B(x[925]), .Z(n13932) );
  AND U10682 ( .A(n4674), .B(n13932), .Z(n26132) );
  NANDN U10683 ( .A(x[923]), .B(y[923]), .Z(n26131) );
  NANDN U10684 ( .A(x[919]), .B(y[919]), .Z(n13934) );
  NANDN U10685 ( .A(x[921]), .B(y[921]), .Z(n6675) );
  NANDN U10686 ( .A(x[920]), .B(y[920]), .Z(n4675) );
  AND U10687 ( .A(n6675), .B(n4675), .Z(n24491) );
  AND U10688 ( .A(n13934), .B(n24491), .Z(n6674) );
  ANDN U10689 ( .B(x[918]), .A(y[918]), .Z(n13936) );
  NANDN U10690 ( .A(x[918]), .B(y[918]), .Z(n13935) );
  NANDN U10691 ( .A(x[917]), .B(y[917]), .Z(n13938) );
  AND U10692 ( .A(n13935), .B(n13938), .Z(n6670) );
  ANDN U10693 ( .B(x[916]), .A(y[916]), .Z(n13940) );
  NANDN U10694 ( .A(x[916]), .B(y[916]), .Z(n13939) );
  ANDN U10695 ( .B(x[914]), .A(y[914]), .Z(n26119) );
  NANDN U10696 ( .A(x[913]), .B(y[913]), .Z(n16584) );
  NANDN U10697 ( .A(x[914]), .B(y[914]), .Z(n16591) );
  AND U10698 ( .A(n16584), .B(n16591), .Z(n24492) );
  ANDN U10699 ( .B(x[913]), .A(y[913]), .Z(n16588) );
  NANDN U10700 ( .A(y[912]), .B(x[912]), .Z(n13943) );
  NANDN U10701 ( .A(n16588), .B(n13943), .Z(n24493) );
  NANDN U10702 ( .A(x[911]), .B(y[911]), .Z(n13945) );
  NANDN U10703 ( .A(x[912]), .B(y[912]), .Z(n16583) );
  AND U10704 ( .A(n13945), .B(n16583), .Z(n24494) );
  NANDN U10705 ( .A(x[909]), .B(y[909]), .Z(n16575) );
  NANDN U10706 ( .A(x[910]), .B(y[910]), .Z(n13946) );
  AND U10707 ( .A(n16575), .B(n13946), .Z(n26118) );
  ANDN U10708 ( .B(x[908]), .A(y[908]), .Z(n16573) );
  NANDN U10709 ( .A(y[909]), .B(x[909]), .Z(n13948) );
  NANDN U10710 ( .A(n16573), .B(n13948), .Z(n26117) );
  NANDN U10711 ( .A(x[908]), .B(y[908]), .Z(n26116) );
  ANDN U10712 ( .B(x[907]), .A(y[907]), .Z(n26115) );
  NANDN U10713 ( .A(x[906]), .B(y[906]), .Z(n13950) );
  NANDN U10714 ( .A(y[905]), .B(x[905]), .Z(n13952) );
  ANDN U10715 ( .B(x[904]), .A(y[904]), .Z(n13955) );
  ANDN U10716 ( .B(n13952), .A(n13955), .Z(n6650) );
  ANDN U10717 ( .B(y[903]), .A(x[903]), .Z(n16564) );
  NANDN U10718 ( .A(y[903]), .B(x[903]), .Z(n13956) );
  ANDN U10719 ( .B(y[901]), .A(x[901]), .Z(n13957) );
  NANDN U10720 ( .A(y[900]), .B(x[900]), .Z(n13960) );
  ANDN U10721 ( .B(y[900]), .A(x[900]), .Z(n13958) );
  NANDN U10722 ( .A(x[899]), .B(y[899]), .Z(n26104) );
  NANDN U10723 ( .A(y[898]), .B(x[898]), .Z(n26105) );
  NANDN U10724 ( .A(x[897]), .B(y[897]), .Z(n13965) );
  NANDN U10725 ( .A(y[896]), .B(x[896]), .Z(n16553) );
  NANDN U10726 ( .A(y[897]), .B(x[897]), .Z(n13962) );
  NAND U10727 ( .A(n16553), .B(n13962), .Z(n26102) );
  NANDN U10728 ( .A(x[895]), .B(y[895]), .Z(n13967) );
  NANDN U10729 ( .A(y[894]), .B(x[894]), .Z(n26100) );
  NANDN U10730 ( .A(y[895]), .B(x[895]), .Z(n24497) );
  NAND U10731 ( .A(n26100), .B(n24497), .Z(n6631) );
  NANDN U10732 ( .A(x[893]), .B(y[893]), .Z(n26099) );
  NANDN U10733 ( .A(y[892]), .B(x[892]), .Z(n16544) );
  NANDN U10734 ( .A(y[893]), .B(x[893]), .Z(n16549) );
  NAND U10735 ( .A(n16544), .B(n16549), .Z(n26098) );
  NANDN U10736 ( .A(x[891]), .B(y[891]), .Z(n13970) );
  NANDN U10737 ( .A(y[890]), .B(x[890]), .Z(n26093) );
  ANDN U10738 ( .B(y[888]), .A(x[888]), .Z(n13972) );
  NANDN U10739 ( .A(x[887]), .B(y[887]), .Z(n13973) );
  NANDN U10740 ( .A(y[887]), .B(x[887]), .Z(n26090) );
  NANDN U10741 ( .A(x[886]), .B(y[886]), .Z(n13974) );
  NANDN U10742 ( .A(y[885]), .B(x[885]), .Z(n13976) );
  NANDN U10743 ( .A(y[884]), .B(x[884]), .Z(n13978) );
  AND U10744 ( .A(n13976), .B(n13978), .Z(n6613) );
  ANDN U10745 ( .B(y[883]), .A(x[883]), .Z(n26086) );
  ANDN U10746 ( .B(y[881]), .A(x[881]), .Z(n16521) );
  ANDN U10747 ( .B(y[882]), .A(x[882]), .Z(n16528) );
  NOR U10748 ( .A(n16521), .B(n16528), .Z(n26084) );
  NANDN U10749 ( .A(y[880]), .B(x[880]), .Z(n16517) );
  NANDN U10750 ( .A(y[881]), .B(x[881]), .Z(n13979) );
  NAND U10751 ( .A(n16517), .B(n13979), .Z(n26083) );
  ANDN U10752 ( .B(y[879]), .A(x[879]), .Z(n16512) );
  ANDN U10753 ( .B(y[880]), .A(x[880]), .Z(n16522) );
  OR U10754 ( .A(n16512), .B(n16522), .Z(n24502) );
  NANDN U10755 ( .A(y[878]), .B(x[878]), .Z(n16509) );
  NANDN U10756 ( .A(y[879]), .B(x[879]), .Z(n16516) );
  AND U10757 ( .A(n16509), .B(n16516), .Z(n26082) );
  NANDN U10758 ( .A(y[875]), .B(x[875]), .Z(n24504) );
  NANDN U10759 ( .A(y[874]), .B(x[874]), .Z(n26076) );
  AND U10760 ( .A(n24504), .B(n26076), .Z(n6599) );
  ANDN U10761 ( .B(y[873]), .A(x[873]), .Z(n13982) );
  NANDN U10762 ( .A(y[872]), .B(x[872]), .Z(n13984) );
  NANDN U10763 ( .A(y[873]), .B(x[873]), .Z(n13981) );
  AND U10764 ( .A(n13984), .B(n13981), .Z(n24505) );
  ANDN U10765 ( .B(y[871]), .A(x[871]), .Z(n13985) );
  NANDN U10766 ( .A(y[870]), .B(x[870]), .Z(n6592) );
  XOR U10767 ( .A(x[870]), .B(y[870]), .Z(n13986) );
  NANDN U10768 ( .A(y[868]), .B(x[868]), .Z(n13991) );
  NANDN U10769 ( .A(x[867]), .B(y[867]), .Z(n13993) );
  NANDN U10770 ( .A(y[867]), .B(x[867]), .Z(n13990) );
  ANDN U10771 ( .B(y[865]), .A(x[865]), .Z(n26066) );
  NANDN U10772 ( .A(y[864]), .B(x[864]), .Z(n16479) );
  NANDN U10773 ( .A(y[865]), .B(x[865]), .Z(n16485) );
  AND U10774 ( .A(n16479), .B(n16485), .Z(n26064) );
  ANDN U10775 ( .B(y[863]), .A(x[863]), .Z(n16477) );
  ANDN U10776 ( .B(y[864]), .A(x[864]), .Z(n16482) );
  OR U10777 ( .A(n16477), .B(n16482), .Z(n26063) );
  NANDN U10778 ( .A(y[862]), .B(x[862]), .Z(n13995) );
  NANDN U10779 ( .A(y[863]), .B(x[863]), .Z(n16480) );
  AND U10780 ( .A(n13995), .B(n16480), .Z(n26062) );
  ANDN U10781 ( .B(y[861]), .A(x[861]), .Z(n16469) );
  ANDN U10782 ( .B(y[862]), .A(x[862]), .Z(n16474) );
  NOR U10783 ( .A(n16469), .B(n16474), .Z(n26061) );
  NANDN U10784 ( .A(y[860]), .B(x[860]), .Z(n16465) );
  NANDN U10785 ( .A(y[861]), .B(x[861]), .Z(n13994) );
  NAND U10786 ( .A(n16465), .B(n13994), .Z(n24506) );
  ANDN U10787 ( .B(y[859]), .A(x[859]), .Z(n16460) );
  ANDN U10788 ( .B(y[860]), .A(x[860]), .Z(n16470) );
  NOR U10789 ( .A(n16460), .B(n16470), .Z(n26060) );
  ANDN U10790 ( .B(y[857]), .A(x[857]), .Z(n16454) );
  ANDN U10791 ( .B(y[858]), .A(x[858]), .Z(n16463) );
  NOR U10792 ( .A(n16454), .B(n16463), .Z(n26059) );
  NANDN U10793 ( .A(y[856]), .B(x[856]), .Z(n26056) );
  NANDN U10794 ( .A(y[857]), .B(x[857]), .Z(n26058) );
  NAND U10795 ( .A(n26056), .B(n26058), .Z(n6571) );
  NANDN U10796 ( .A(x[854]), .B(y[854]), .Z(n13998) );
  NANDN U10797 ( .A(x[853]), .B(y[853]), .Z(n14003) );
  AND U10798 ( .A(n13998), .B(n14003), .Z(n6565) );
  NANDN U10799 ( .A(y[853]), .B(x[853]), .Z(n14001) );
  NANDN U10800 ( .A(y[852]), .B(x[852]), .Z(n14004) );
  ANDN U10801 ( .B(y[851]), .A(x[851]), .Z(n26050) );
  NANDN U10802 ( .A(y[851]), .B(x[851]), .Z(n14005) );
  ANDN U10803 ( .B(y[850]), .A(x[850]), .Z(n14006) );
  NANDN U10804 ( .A(x[849]), .B(y[849]), .Z(n16444) );
  NANDN U10805 ( .A(n14006), .B(n16444), .Z(n26047) );
  NANDN U10806 ( .A(y[849]), .B(x[849]), .Z(n4677) );
  NANDN U10807 ( .A(y[848]), .B(x[848]), .Z(n4676) );
  NAND U10808 ( .A(n4677), .B(n4676), .Z(n26046) );
  NANDN U10809 ( .A(y[846]), .B(x[846]), .Z(n4678) );
  NANDN U10810 ( .A(y[847]), .B(x[847]), .Z(n14007) );
  AND U10811 ( .A(n4678), .B(n14007), .Z(n26044) );
  ANDN U10812 ( .B(x[844]), .A(y[844]), .Z(n16435) );
  ANDN U10813 ( .B(x[845]), .A(y[845]), .Z(n16440) );
  OR U10814 ( .A(n16435), .B(n16440), .Z(n24509) );
  NANDN U10815 ( .A(x[843]), .B(y[843]), .Z(n14011) );
  ANDN U10816 ( .B(x[843]), .A(y[843]), .Z(n26042) );
  NANDN U10817 ( .A(y[842]), .B(x[842]), .Z(n26040) );
  NANDN U10818 ( .A(n26042), .B(n26040), .Z(n6546) );
  ANDN U10819 ( .B(x[840]), .A(y[840]), .Z(n16425) );
  ANDN U10820 ( .B(x[841]), .A(y[841]), .Z(n16431) );
  NOR U10821 ( .A(n16425), .B(n16431), .Z(n26038) );
  NANDN U10822 ( .A(x[839]), .B(y[839]), .Z(n4680) );
  NANDN U10823 ( .A(x[838]), .B(y[838]), .Z(n4679) );
  NAND U10824 ( .A(n4680), .B(n4679), .Z(n16421) );
  NANDN U10825 ( .A(x[837]), .B(y[837]), .Z(n4682) );
  NANDN U10826 ( .A(x[836]), .B(y[836]), .Z(n4681) );
  AND U10827 ( .A(n4682), .B(n4681), .Z(n26033) );
  NANDN U10828 ( .A(y[835]), .B(x[835]), .Z(n4684) );
  NANDN U10829 ( .A(y[836]), .B(x[836]), .Z(n4683) );
  NAND U10830 ( .A(n4684), .B(n4683), .Z(n26031) );
  NANDN U10831 ( .A(x[835]), .B(y[835]), .Z(n14015) );
  NANDN U10832 ( .A(y[834]), .B(x[834]), .Z(n14017) );
  XNOR U10833 ( .A(x[834]), .B(y[834]), .Z(n6531) );
  NANDN U10834 ( .A(x[833]), .B(y[833]), .Z(n14018) );
  NANDN U10835 ( .A(x[832]), .B(y[832]), .Z(n14019) );
  NANDN U10836 ( .A(x[831]), .B(y[831]), .Z(n26021) );
  AND U10837 ( .A(n14019), .B(n26021), .Z(n6526) );
  ANDN U10838 ( .B(x[830]), .A(y[830]), .Z(n16410) );
  ANDN U10839 ( .B(x[831]), .A(y[831]), .Z(n16414) );
  OR U10840 ( .A(n16410), .B(n16414), .Z(n26019) );
  NANDN U10841 ( .A(x[830]), .B(y[830]), .Z(n4686) );
  NANDN U10842 ( .A(x[829]), .B(y[829]), .Z(n4685) );
  AND U10843 ( .A(n4686), .B(n4685), .Z(n26017) );
  NANDN U10844 ( .A(y[828]), .B(x[828]), .Z(n4687) );
  ANDN U10845 ( .B(x[829]), .A(y[829]), .Z(n16402) );
  ANDN U10846 ( .B(n4687), .A(n16402), .Z(n26015) );
  NANDN U10847 ( .A(x[827]), .B(y[827]), .Z(n16398) );
  NANDN U10848 ( .A(x[828]), .B(y[828]), .Z(n4688) );
  AND U10849 ( .A(n16398), .B(n4688), .Z(n26012) );
  NANDN U10850 ( .A(y[826]), .B(x[826]), .Z(n16394) );
  NANDN U10851 ( .A(y[827]), .B(x[827]), .Z(n26011) );
  NAND U10852 ( .A(n16394), .B(n26011), .Z(n6520) );
  NANDN U10853 ( .A(x[826]), .B(y[826]), .Z(n26009) );
  ANDN U10854 ( .B(x[824]), .A(y[824]), .Z(n16391) );
  ANDN U10855 ( .B(x[825]), .A(y[825]), .Z(n16397) );
  OR U10856 ( .A(n16391), .B(n16397), .Z(n26003) );
  NANDN U10857 ( .A(x[823]), .B(y[823]), .Z(n14020) );
  NANDN U10858 ( .A(y[822]), .B(x[822]), .Z(n14023) );
  NANDN U10859 ( .A(x[821]), .B(y[821]), .Z(n14025) );
  ANDN U10860 ( .B(x[820]), .A(y[820]), .Z(n14026) );
  NANDN U10861 ( .A(x[820]), .B(y[820]), .Z(n14024) );
  NANDN U10862 ( .A(y[819]), .B(x[819]), .Z(n14027) );
  NANDN U10863 ( .A(y[818]), .B(x[818]), .Z(n14031) );
  AND U10864 ( .A(n14027), .B(n14031), .Z(n6505) );
  ANDN U10865 ( .B(y[818]), .A(x[818]), .Z(n14028) );
  NANDN U10866 ( .A(x[817]), .B(y[817]), .Z(n14032) );
  NANDN U10867 ( .A(y[816]), .B(x[816]), .Z(n14034) );
  NANDN U10868 ( .A(x[816]), .B(y[816]), .Z(n14033) );
  NANDN U10869 ( .A(y[815]), .B(x[815]), .Z(n14035) );
  ANDN U10870 ( .B(x[814]), .A(y[814]), .Z(n14038) );
  ANDN U10871 ( .B(n14035), .A(n14038), .Z(n6497) );
  ANDN U10872 ( .B(y[813]), .A(x[813]), .Z(n14040) );
  NANDN U10873 ( .A(y[813]), .B(x[813]), .Z(n14039) );
  ANDN U10874 ( .B(y[811]), .A(x[811]), .Z(n14043) );
  NANDN U10875 ( .A(y[811]), .B(x[811]), .Z(n14042) );
  NANDN U10876 ( .A(y[810]), .B(x[810]), .Z(n6487) );
  NANDN U10877 ( .A(x[810]), .B(y[810]), .Z(n14044) );
  NANDN U10878 ( .A(x[809]), .B(y[809]), .Z(n14048) );
  ANDN U10879 ( .B(x[809]), .A(y[809]), .Z(n14046) );
  ANDN U10880 ( .B(x[808]), .A(y[808]), .Z(n14049) );
  NANDN U10881 ( .A(x[808]), .B(y[808]), .Z(n14047) );
  NANDN U10882 ( .A(y[807]), .B(x[807]), .Z(n14050) );
  ANDN U10883 ( .B(x[806]), .A(y[806]), .Z(n14055) );
  ANDN U10884 ( .B(n14050), .A(n14055), .Z(n6479) );
  NANDN U10885 ( .A(x[805]), .B(y[805]), .Z(n14060) );
  NANDN U10886 ( .A(y[805]), .B(x[805]), .Z(n14056) );
  ANDN U10887 ( .B(y[803]), .A(x[803]), .Z(n14063) );
  NANDN U10888 ( .A(y[802]), .B(x[802]), .Z(n14067) );
  ANDN U10889 ( .B(y[801]), .A(x[801]), .Z(n14068) );
  NANDN U10890 ( .A(y[801]), .B(x[801]), .Z(n14066) );
  NANDN U10891 ( .A(x[800]), .B(y[800]), .Z(n14069) );
  ANDN U10892 ( .B(y[799]), .A(x[799]), .Z(n14072) );
  ANDN U10893 ( .B(n14069), .A(n14072), .Z(n6464) );
  ANDN U10894 ( .B(x[798]), .A(y[798]), .Z(n14074) );
  NANDN U10895 ( .A(x[798]), .B(y[798]), .Z(n14073) );
  NANDN U10896 ( .A(y[796]), .B(x[796]), .Z(n14079) );
  ANDN U10897 ( .B(x[795]), .A(y[795]), .Z(n14078) );
  NANDN U10898 ( .A(x[795]), .B(y[795]), .Z(n4690) );
  NANDN U10899 ( .A(x[794]), .B(y[794]), .Z(n4689) );
  AND U10900 ( .A(n4690), .B(n4689), .Z(n25946) );
  NANDN U10901 ( .A(y[794]), .B(x[794]), .Z(n4692) );
  NANDN U10902 ( .A(y[793]), .B(x[793]), .Z(n4691) );
  AND U10903 ( .A(n4692), .B(n4691), .Z(n14080) );
  NANDN U10904 ( .A(x[792]), .B(y[792]), .Z(n4694) );
  NANDN U10905 ( .A(x[793]), .B(y[793]), .Z(n4693) );
  NAND U10906 ( .A(n4694), .B(n4693), .Z(n14081) );
  NANDN U10907 ( .A(y[792]), .B(x[792]), .Z(n4696) );
  NANDN U10908 ( .A(y[791]), .B(x[791]), .Z(n4695) );
  AND U10909 ( .A(n4696), .B(n4695), .Z(n14082) );
  NANDN U10910 ( .A(x[788]), .B(y[788]), .Z(n4698) );
  NANDN U10911 ( .A(x[789]), .B(y[789]), .Z(n4697) );
  NAND U10912 ( .A(n4698), .B(n4697), .Z(n16352) );
  NANDN U10913 ( .A(y[788]), .B(x[788]), .Z(n4700) );
  NANDN U10914 ( .A(y[787]), .B(x[787]), .Z(n4699) );
  AND U10915 ( .A(n4700), .B(n4699), .Z(n14084) );
  NANDN U10916 ( .A(x[786]), .B(y[786]), .Z(n14086) );
  ANDN U10917 ( .B(y[787]), .A(x[787]), .Z(n14085) );
  ANDN U10918 ( .B(n14086), .A(n14085), .Z(n6442) );
  XNOR U10919 ( .A(y[786]), .B(x[786]), .Z(n6440) );
  NANDN U10920 ( .A(y[785]), .B(x[785]), .Z(n14087) );
  NANDN U10921 ( .A(x[784]), .B(y[784]), .Z(n4702) );
  NANDN U10922 ( .A(x[785]), .B(y[785]), .Z(n4701) );
  NAND U10923 ( .A(n4702), .B(n4701), .Z(n14089) );
  ANDN U10924 ( .B(x[781]), .A(y[781]), .Z(n14090) );
  NANDN U10925 ( .A(x[780]), .B(y[780]), .Z(n4704) );
  NANDN U10926 ( .A(x[781]), .B(y[781]), .Z(n4703) );
  NAND U10927 ( .A(n4704), .B(n4703), .Z(n24510) );
  NANDN U10928 ( .A(y[780]), .B(x[780]), .Z(n4706) );
  NANDN U10929 ( .A(y[779]), .B(x[779]), .Z(n4705) );
  AND U10930 ( .A(n4706), .B(n4705), .Z(n24511) );
  NANDN U10931 ( .A(y[774]), .B(x[774]), .Z(n14092) );
  NANDN U10932 ( .A(x[773]), .B(y[773]), .Z(n14094) );
  XNOR U10933 ( .A(y[773]), .B(x[773]), .Z(n6407) );
  NANDN U10934 ( .A(y[772]), .B(x[772]), .Z(n14096) );
  ANDN U10935 ( .B(y[771]), .A(x[771]), .Z(n14097) );
  NANDN U10936 ( .A(y[771]), .B(x[771]), .Z(n14095) );
  ANDN U10937 ( .B(y[769]), .A(x[769]), .Z(n16330) );
  NANDN U10938 ( .A(y[768]), .B(x[768]), .Z(n14102) );
  ANDN U10939 ( .B(y[768]), .A(x[768]), .Z(n16329) );
  NANDN U10940 ( .A(x[767]), .B(y[767]), .Z(n14103) );
  ANDN U10941 ( .B(x[766]), .A(y[766]), .Z(n14105) );
  NANDN U10942 ( .A(x[766]), .B(y[766]), .Z(n14104) );
  NANDN U10943 ( .A(y[765]), .B(x[765]), .Z(n14106) );
  ANDN U10944 ( .B(x[764]), .A(y[764]), .Z(n14109) );
  ANDN U10945 ( .B(n14106), .A(n14109), .Z(n6390) );
  ANDN U10946 ( .B(y[763]), .A(x[763]), .Z(n16320) );
  NANDN U10947 ( .A(y[763]), .B(x[763]), .Z(n14110) );
  ANDN U10948 ( .B(y[761]), .A(x[761]), .Z(n14111) );
  NANDN U10949 ( .A(y[760]), .B(x[760]), .Z(n6381) );
  ANDN U10950 ( .B(y[760]), .A(x[760]), .Z(n14112) );
  NANDN U10951 ( .A(x[759]), .B(y[759]), .Z(n14117) );
  NANDN U10952 ( .A(y[758]), .B(x[758]), .Z(n14120) );
  NANDN U10953 ( .A(x[758]), .B(y[758]), .Z(n14118) );
  ANDN U10954 ( .B(x[756]), .A(y[756]), .Z(n6373) );
  NANDN U10955 ( .A(x[755]), .B(y[755]), .Z(n14125) );
  ANDN U10956 ( .B(x[755]), .A(y[755]), .Z(n14121) );
  NANDN U10957 ( .A(y[754]), .B(x[754]), .Z(n6367) );
  ANDN U10958 ( .B(y[753]), .A(x[753]), .Z(n14128) );
  NANDN U10959 ( .A(y[753]), .B(x[753]), .Z(n14127) );
  ANDN U10960 ( .B(y[751]), .A(x[751]), .Z(n16302) );
  NANDN U10961 ( .A(y[750]), .B(x[750]), .Z(n6357) );
  ANDN U10962 ( .B(y[749]), .A(x[749]), .Z(n14132) );
  NANDN U10963 ( .A(y[749]), .B(x[749]), .Z(n16300) );
  NANDN U10964 ( .A(x[747]), .B(y[747]), .Z(n14136) );
  XNOR U10965 ( .A(x[748]), .B(y[748]), .Z(n14134) );
  AND U10966 ( .A(n14136), .B(n14134), .Z(n6350) );
  ANDN U10967 ( .B(x[747]), .A(y[747]), .Z(n14133) );
  NANDN U10968 ( .A(y[746]), .B(x[746]), .Z(n14137) );
  ANDN U10969 ( .B(y[745]), .A(x[745]), .Z(n16292) );
  NANDN U10970 ( .A(y[745]), .B(x[745]), .Z(n14138) );
  NANDN U10971 ( .A(x[744]), .B(y[744]), .Z(n16293) );
  ANDN U10972 ( .B(y[743]), .A(x[743]), .Z(n14141) );
  ANDN U10973 ( .B(n16293), .A(n14141), .Z(n6342) );
  ANDN U10974 ( .B(x[742]), .A(y[742]), .Z(n6339) );
  NANDN U10975 ( .A(x[742]), .B(y[742]), .Z(n14143) );
  ANDN U10976 ( .B(x[740]), .A(y[740]), .Z(n6335) );
  NANDN U10977 ( .A(x[739]), .B(y[739]), .Z(n16285) );
  ANDN U10978 ( .B(x[738]), .A(y[738]), .Z(n14152) );
  NANDN U10979 ( .A(x[738]), .B(y[738]), .Z(n16284) );
  NANDN U10980 ( .A(y[737]), .B(x[737]), .Z(n14153) );
  ANDN U10981 ( .B(x[736]), .A(y[736]), .Z(n4707) );
  ANDN U10982 ( .B(n14153), .A(n4707), .Z(n6326) );
  ANDN U10983 ( .B(y[735]), .A(x[735]), .Z(n14158) );
  NANDN U10984 ( .A(y[735]), .B(x[735]), .Z(n14156) );
  ANDN U10985 ( .B(y[733]), .A(x[733]), .Z(n16276) );
  NANDN U10986 ( .A(y[732]), .B(x[732]), .Z(n6316) );
  ANDN U10987 ( .B(y[731]), .A(x[731]), .Z(n14162) );
  NANDN U10988 ( .A(y[731]), .B(x[731]), .Z(n16274) );
  NANDN U10989 ( .A(x[730]), .B(y[730]), .Z(n14163) );
  NANDN U10990 ( .A(x[729]), .B(y[729]), .Z(n14168) );
  AND U10991 ( .A(n14163), .B(n14168), .Z(n6310) );
  ANDN U10992 ( .B(x[729]), .A(y[729]), .Z(n14164) );
  NANDN U10993 ( .A(y[728]), .B(x[728]), .Z(n14170) );
  ANDN U10994 ( .B(y[727]), .A(x[727]), .Z(n16266) );
  NANDN U10995 ( .A(y[727]), .B(x[727]), .Z(n14169) );
  NANDN U10996 ( .A(x[726]), .B(y[726]), .Z(n16267) );
  ANDN U10997 ( .B(y[725]), .A(x[725]), .Z(n14174) );
  ANDN U10998 ( .B(n16267), .A(n14174), .Z(n6302) );
  ANDN U10999 ( .B(x[724]), .A(y[724]), .Z(n14176) );
  NANDN U11000 ( .A(x[724]), .B(y[724]), .Z(n14175) );
  NANDN U11001 ( .A(y[723]), .B(x[723]), .Z(n14177) );
  ANDN U11002 ( .B(x[722]), .A(y[722]), .Z(n4708) );
  ANDN U11003 ( .B(n14177), .A(n4708), .Z(n6296) );
  ANDN U11004 ( .B(y[721]), .A(x[721]), .Z(n16258) );
  NANDN U11005 ( .A(y[721]), .B(x[721]), .Z(n14180) );
  ANDN U11006 ( .B(y[719]), .A(x[719]), .Z(n14183) );
  NANDN U11007 ( .A(y[718]), .B(x[718]), .Z(n14185) );
  ANDN U11008 ( .B(y[717]), .A(x[717]), .Z(n14187) );
  NANDN U11009 ( .A(y[717]), .B(x[717]), .Z(n14186) );
  NANDN U11010 ( .A(x[716]), .B(y[716]), .Z(n14188) );
  NANDN U11011 ( .A(x[715]), .B(y[715]), .Z(n16248) );
  AND U11012 ( .A(n14188), .B(n16248), .Z(n6282) );
  ANDN U11013 ( .B(x[715]), .A(y[715]), .Z(n14189) );
  NANDN U11014 ( .A(y[714]), .B(x[714]), .Z(n6279) );
  ANDN U11015 ( .B(y[714]), .A(x[714]), .Z(n16247) );
  NANDN U11016 ( .A(y[713]), .B(x[713]), .Z(n16245) );
  NANDN U11017 ( .A(y[712]), .B(x[712]), .Z(n4709) );
  AND U11018 ( .A(n16245), .B(n4709), .Z(n6275) );
  XNOR U11019 ( .A(x[712]), .B(y[712]), .Z(n14193) );
  NANDN U11020 ( .A(y[710]), .B(x[710]), .Z(n14197) );
  NANDN U11021 ( .A(x[707]), .B(y[707]), .Z(n14200) );
  NANDN U11022 ( .A(y[706]), .B(x[706]), .Z(n14204) );
  NANDN U11023 ( .A(x[706]), .B(y[706]), .Z(n14201) );
  ANDN U11024 ( .B(x[705]), .A(y[705]), .Z(n14202) );
  ANDN U11025 ( .B(x[704]), .A(y[704]), .Z(n4710) );
  NOR U11026 ( .A(n14202), .B(n4710), .Z(n6259) );
  ANDN U11027 ( .B(y[703]), .A(x[703]), .Z(n16228) );
  NANDN U11028 ( .A(y[703]), .B(x[703]), .Z(n14209) );
  ANDN U11029 ( .B(y[701]), .A(x[701]), .Z(n14210) );
  NANDN U11030 ( .A(y[700]), .B(x[700]), .Z(n14213) );
  ANDN U11031 ( .B(y[699]), .A(x[699]), .Z(n14215) );
  NANDN U11032 ( .A(y[699]), .B(x[699]), .Z(n14214) );
  NANDN U11033 ( .A(x[698]), .B(y[698]), .Z(n14217) );
  NANDN U11034 ( .A(x[697]), .B(y[697]), .Z(n16219) );
  NAND U11035 ( .A(n14217), .B(n16219), .Z(n6244) );
  NANDN U11036 ( .A(y[697]), .B(x[697]), .Z(n14219) );
  NANDN U11037 ( .A(y[696]), .B(x[696]), .Z(n16216) );
  AND U11038 ( .A(n14219), .B(n16216), .Z(n6242) );
  NANDN U11039 ( .A(x[695]), .B(y[695]), .Z(n14221) );
  NANDN U11040 ( .A(y[694]), .B(x[694]), .Z(n14222) );
  ANDN U11041 ( .B(y[693]), .A(x[693]), .Z(n14224) );
  NANDN U11042 ( .A(y[693]), .B(x[693]), .Z(n14223) );
  ANDN U11043 ( .B(y[691]), .A(x[691]), .Z(n16208) );
  IV U11044 ( .A(n16208), .Z(n25859) );
  ANDN U11045 ( .B(y[692]), .A(x[692]), .Z(n14225) );
  ANDN U11046 ( .B(n25859), .A(n14225), .Z(n6232) );
  ANDN U11047 ( .B(y[689]), .A(x[689]), .Z(n16201) );
  ANDN U11048 ( .B(y[690]), .A(x[690]), .Z(n16205) );
  NOR U11049 ( .A(n16201), .B(n16205), .Z(n25858) );
  NANDN U11050 ( .A(y[689]), .B(x[689]), .Z(n25857) );
  NANDN U11051 ( .A(x[687]), .B(y[687]), .Z(n14228) );
  ANDN U11052 ( .B(x[686]), .A(y[686]), .Z(n6224) );
  NANDN U11053 ( .A(x[685]), .B(y[685]), .Z(n14230) );
  ANDN U11054 ( .B(x[684]), .A(y[684]), .Z(n6218) );
  NANDN U11055 ( .A(x[684]), .B(y[684]), .Z(n14231) );
  NANDN U11056 ( .A(y[682]), .B(x[682]), .Z(n4711) );
  NANDN U11057 ( .A(y[683]), .B(x[683]), .Z(n14232) );
  AND U11058 ( .A(n4711), .B(n14232), .Z(n6214) );
  ANDN U11059 ( .B(y[682]), .A(x[682]), .Z(n14233) );
  NANDN U11060 ( .A(x[681]), .B(y[681]), .Z(n14237) );
  ANDN U11061 ( .B(x[681]), .A(y[681]), .Z(n14236) );
  ANDN U11062 ( .B(x[680]), .A(y[680]), .Z(n14239) );
  NANDN U11063 ( .A(x[680]), .B(y[680]), .Z(n14238) );
  ANDN U11064 ( .B(x[678]), .A(y[678]), .Z(n6206) );
  NANDN U11065 ( .A(x[677]), .B(y[677]), .Z(n14245) );
  NANDN U11066 ( .A(x[676]), .B(y[676]), .Z(n14246) );
  NANDN U11067 ( .A(x[675]), .B(y[675]), .Z(n14249) );
  AND U11068 ( .A(n14246), .B(n14249), .Z(n6198) );
  NANDN U11069 ( .A(y[674]), .B(x[674]), .Z(n14252) );
  NANDN U11070 ( .A(x[674]), .B(y[674]), .Z(n14250) );
  ANDN U11071 ( .B(x[672]), .A(y[672]), .Z(n6192) );
  NANDN U11072 ( .A(x[671]), .B(y[671]), .Z(n14257) );
  NANDN U11073 ( .A(x[670]), .B(y[670]), .Z(n14258) );
  NANDN U11074 ( .A(x[669]), .B(y[669]), .Z(n14261) );
  AND U11075 ( .A(n14258), .B(n14261), .Z(n6185) );
  NANDN U11076 ( .A(y[668]), .B(x[668]), .Z(n14264) );
  NANDN U11077 ( .A(x[668]), .B(y[668]), .Z(n14262) );
  NANDN U11078 ( .A(y[666]), .B(x[666]), .Z(n14268) );
  ANDN U11079 ( .B(x[665]), .A(y[665]), .Z(n14267) );
  NANDN U11080 ( .A(x[665]), .B(y[665]), .Z(n4713) );
  NANDN U11081 ( .A(x[664]), .B(y[664]), .Z(n4712) );
  AND U11082 ( .A(n4713), .B(n4712), .Z(n25816) );
  NANDN U11083 ( .A(x[663]), .B(y[663]), .Z(n14270) );
  NANDN U11084 ( .A(y[662]), .B(x[662]), .Z(n14272) );
  XNOR U11085 ( .A(x[662]), .B(y[662]), .Z(n6169) );
  NANDN U11086 ( .A(x[661]), .B(y[661]), .Z(n14273) );
  ANDN U11087 ( .B(x[660]), .A(y[660]), .Z(n6165) );
  NANDN U11088 ( .A(x[660]), .B(y[660]), .Z(n14274) );
  ANDN U11089 ( .B(x[658]), .A(y[658]), .Z(n14279) );
  NANDN U11090 ( .A(x[657]), .B(y[657]), .Z(n14281) );
  NANDN U11091 ( .A(x[656]), .B(y[656]), .Z(n14282) );
  NANDN U11092 ( .A(x[655]), .B(y[655]), .Z(n14286) );
  AND U11093 ( .A(n14282), .B(n14286), .Z(n6155) );
  NANDN U11094 ( .A(y[654]), .B(x[654]), .Z(n14288) );
  NANDN U11095 ( .A(x[654]), .B(y[654]), .Z(n14285) );
  ANDN U11096 ( .B(x[653]), .A(y[653]), .Z(n14287) );
  XNOR U11097 ( .A(x[652]), .B(y[652]), .Z(n14292) );
  NANDN U11098 ( .A(x[651]), .B(y[651]), .Z(n14293) );
  NANDN U11099 ( .A(x[649]), .B(y[649]), .Z(n14297) );
  XNOR U11100 ( .A(x[650]), .B(y[650]), .Z(n14296) );
  AND U11101 ( .A(n14297), .B(n14296), .Z(n6141) );
  ANDN U11102 ( .B(x[648]), .A(y[648]), .Z(n6138) );
  XNOR U11103 ( .A(x[648]), .B(y[648]), .Z(n14300) );
  NANDN U11104 ( .A(x[647]), .B(y[647]), .Z(n14302) );
  NANDN U11105 ( .A(y[646]), .B(x[646]), .Z(n14303) );
  NANDN U11106 ( .A(x[645]), .B(y[645]), .Z(n14306) );
  NANDN U11107 ( .A(x[644]), .B(y[644]), .Z(n14305) );
  NANDN U11108 ( .A(x[643]), .B(y[643]), .Z(n14309) );
  AND U11109 ( .A(n14305), .B(n14309), .Z(n6128) );
  ANDN U11110 ( .B(x[642]), .A(y[642]), .Z(n14311) );
  NANDN U11111 ( .A(x[642]), .B(y[642]), .Z(n14310) );
  ANDN U11112 ( .B(x[640]), .A(y[640]), .Z(n14315) );
  NANDN U11113 ( .A(x[639]), .B(y[639]), .Z(n14317) );
  NANDN U11114 ( .A(x[638]), .B(y[638]), .Z(n14318) );
  NANDN U11115 ( .A(x[637]), .B(y[637]), .Z(n14322) );
  AND U11116 ( .A(n14318), .B(n14322), .Z(n6115) );
  ANDN U11117 ( .B(x[636]), .A(y[636]), .Z(n14323) );
  NANDN U11118 ( .A(x[636]), .B(y[636]), .Z(n14321) );
  ANDN U11119 ( .B(x[634]), .A(y[634]), .Z(n14327) );
  NANDN U11120 ( .A(x[633]), .B(y[633]), .Z(n14329) );
  NANDN U11121 ( .A(x[632]), .B(y[632]), .Z(n14330) );
  NANDN U11122 ( .A(x[631]), .B(y[631]), .Z(n14333) );
  AND U11123 ( .A(n14330), .B(n14333), .Z(n6103) );
  NANDN U11124 ( .A(y[630]), .B(x[630]), .Z(n14336) );
  NANDN U11125 ( .A(x[630]), .B(y[630]), .Z(n14334) );
  ANDN U11126 ( .B(x[628]), .A(y[628]), .Z(n14339) );
  NANDN U11127 ( .A(x[627]), .B(y[627]), .Z(n14341) );
  NANDN U11128 ( .A(x[626]), .B(y[626]), .Z(n14342) );
  NANDN U11129 ( .A(x[625]), .B(y[625]), .Z(n14345) );
  AND U11130 ( .A(n14342), .B(n14345), .Z(n6090) );
  ANDN U11131 ( .B(x[624]), .A(y[624]), .Z(n6087) );
  NANDN U11132 ( .A(x[623]), .B(y[623]), .Z(n14349) );
  XNOR U11133 ( .A(x[624]), .B(y[624]), .Z(n14348) );
  ANDN U11134 ( .B(x[622]), .A(y[622]), .Z(n14351) );
  NANDN U11135 ( .A(x[621]), .B(y[621]), .Z(n14353) );
  NANDN U11136 ( .A(x[620]), .B(y[620]), .Z(n14354) );
  NANDN U11137 ( .A(x[619]), .B(y[619]), .Z(n14357) );
  AND U11138 ( .A(n14354), .B(n14357), .Z(n6077) );
  ANDN U11139 ( .B(x[618]), .A(y[618]), .Z(n14359) );
  NANDN U11140 ( .A(x[618]), .B(y[618]), .Z(n14358) );
  NANDN U11141 ( .A(y[616]), .B(x[616]), .Z(n14364) );
  NANDN U11142 ( .A(x[615]), .B(y[615]), .Z(n14365) );
  NANDN U11143 ( .A(x[614]), .B(y[614]), .Z(n14366) );
  NANDN U11144 ( .A(x[613]), .B(y[613]), .Z(n14369) );
  AND U11145 ( .A(n14366), .B(n14369), .Z(n6064) );
  ANDN U11146 ( .B(x[612]), .A(y[612]), .Z(n6061) );
  NANDN U11147 ( .A(x[612]), .B(y[612]), .Z(n14370) );
  NANDN U11148 ( .A(y[610]), .B(x[610]), .Z(n14376) );
  NANDN U11149 ( .A(x[609]), .B(y[609]), .Z(n14378) );
  NANDN U11150 ( .A(x[608]), .B(y[608]), .Z(n14377) );
  NANDN U11151 ( .A(x[607]), .B(y[607]), .Z(n14382) );
  AND U11152 ( .A(n14377), .B(n14382), .Z(n6051) );
  NANDN U11153 ( .A(y[606]), .B(x[606]), .Z(n14384) );
  NANDN U11154 ( .A(x[606]), .B(y[606]), .Z(n14381) );
  NANDN U11155 ( .A(y[604]), .B(x[604]), .Z(n14388) );
  NANDN U11156 ( .A(x[603]), .B(y[603]), .Z(n14389) );
  NANDN U11157 ( .A(x[602]), .B(y[602]), .Z(n14390) );
  NANDN U11158 ( .A(x[601]), .B(y[601]), .Z(n14394) );
  AND U11159 ( .A(n14390), .B(n14394), .Z(n6039) );
  NANDN U11160 ( .A(y[600]), .B(x[600]), .Z(n14396) );
  NANDN U11161 ( .A(x[600]), .B(y[600]), .Z(n14393) );
  NANDN U11162 ( .A(x[599]), .B(y[599]), .Z(n14398) );
  NANDN U11163 ( .A(y[598]), .B(x[598]), .Z(n14400) );
  XNOR U11164 ( .A(x[598]), .B(y[598]), .Z(n6031) );
  NANDN U11165 ( .A(x[597]), .B(y[597]), .Z(n14401) );
  NANDN U11166 ( .A(x[596]), .B(y[596]), .Z(n14402) );
  ANDN U11167 ( .B(x[595]), .A(y[595]), .Z(n14403) );
  NANDN U11168 ( .A(x[594]), .B(y[594]), .Z(n4715) );
  NANDN U11169 ( .A(x[595]), .B(y[595]), .Z(n4714) );
  AND U11170 ( .A(n4715), .B(n4714), .Z(n25676) );
  NANDN U11171 ( .A(y[594]), .B(x[594]), .Z(n4716) );
  NANDN U11172 ( .A(y[593]), .B(x[593]), .Z(n14405) );
  NAND U11173 ( .A(n4716), .B(n14405), .Z(n6023) );
  NANDN U11174 ( .A(x[593]), .B(y[593]), .Z(n4718) );
  NANDN U11175 ( .A(x[592]), .B(y[592]), .Z(n4717) );
  AND U11176 ( .A(n4718), .B(n4717), .Z(n25672) );
  NANDN U11177 ( .A(x[591]), .B(y[591]), .Z(n14408) );
  NANDN U11178 ( .A(y[590]), .B(x[590]), .Z(n14410) );
  XNOR U11179 ( .A(x[590]), .B(y[590]), .Z(n6015) );
  NANDN U11180 ( .A(x[589]), .B(y[589]), .Z(n14411) );
  NANDN U11181 ( .A(x[588]), .B(y[588]), .Z(n14412) );
  NANDN U11182 ( .A(x[587]), .B(y[587]), .Z(n14415) );
  AND U11183 ( .A(n14412), .B(n14415), .Z(n6009) );
  ANDN U11184 ( .B(x[586]), .A(y[586]), .Z(n14417) );
  NANDN U11185 ( .A(x[586]), .B(y[586]), .Z(n14416) );
  ANDN U11186 ( .B(x[584]), .A(y[584]), .Z(n6003) );
  NANDN U11187 ( .A(x[583]), .B(y[583]), .Z(n14423) );
  NANDN U11188 ( .A(x[582]), .B(y[582]), .Z(n14424) );
  NANDN U11189 ( .A(x[581]), .B(y[581]), .Z(n14427) );
  AND U11190 ( .A(n14424), .B(n14427), .Z(n5995) );
  ANDN U11191 ( .B(x[580]), .A(y[580]), .Z(n16087) );
  NANDN U11192 ( .A(x[579]), .B(y[579]), .Z(n14429) );
  ANDN U11193 ( .B(x[578]), .A(y[578]), .Z(n5989) );
  ANDN U11194 ( .B(x[577]), .A(y[577]), .Z(n14432) );
  NANDN U11195 ( .A(x[577]), .B(y[577]), .Z(n4720) );
  NANDN U11196 ( .A(x[576]), .B(y[576]), .Z(n4719) );
  AND U11197 ( .A(n4720), .B(n4719), .Z(n25643) );
  NANDN U11198 ( .A(x[575]), .B(y[575]), .Z(n14434) );
  NANDN U11199 ( .A(y[574]), .B(x[574]), .Z(n14435) );
  XNOR U11200 ( .A(x[574]), .B(y[574]), .Z(n5978) );
  NANDN U11201 ( .A(x[573]), .B(y[573]), .Z(n14438) );
  NANDN U11202 ( .A(x[572]), .B(y[572]), .Z(n14437) );
  NANDN U11203 ( .A(x[571]), .B(y[571]), .Z(n14442) );
  AND U11204 ( .A(n14437), .B(n14442), .Z(n5973) );
  NANDN U11205 ( .A(y[570]), .B(x[570]), .Z(n14444) );
  NANDN U11206 ( .A(x[570]), .B(y[570]), .Z(n14441) );
  ANDN U11207 ( .B(x[568]), .A(y[568]), .Z(n16074) );
  NANDN U11208 ( .A(x[566]), .B(y[566]), .Z(n14448) );
  NANDN U11209 ( .A(x[565]), .B(y[565]), .Z(n14451) );
  AND U11210 ( .A(n14448), .B(n14451), .Z(n5960) );
  ANDN U11211 ( .B(x[564]), .A(y[564]), .Z(n14453) );
  NANDN U11212 ( .A(x[564]), .B(y[564]), .Z(n14452) );
  NANDN U11213 ( .A(y[562]), .B(x[562]), .Z(n14458) );
  NANDN U11214 ( .A(x[561]), .B(y[561]), .Z(n14459) );
  NANDN U11215 ( .A(x[560]), .B(y[560]), .Z(n14460) );
  ANDN U11216 ( .B(x[559]), .A(y[559]), .Z(n14462) );
  ANDN U11217 ( .B(x[558]), .A(y[558]), .Z(n5944) );
  NANDN U11218 ( .A(x[557]), .B(y[557]), .Z(n14468) );
  XNOR U11219 ( .A(x[558]), .B(y[558]), .Z(n14466) );
  ANDN U11220 ( .B(x[556]), .A(y[556]), .Z(n14469) );
  NANDN U11221 ( .A(x[555]), .B(y[555]), .Z(n14471) );
  NANDN U11222 ( .A(y[555]), .B(x[555]), .Z(n14470) );
  NANDN U11223 ( .A(y[554]), .B(x[554]), .Z(n4721) );
  NAND U11224 ( .A(n14470), .B(n4721), .Z(n5936) );
  NANDN U11225 ( .A(x[553]), .B(y[553]), .Z(n14475) );
  NANDN U11226 ( .A(x[552]), .B(y[552]), .Z(n14476) );
  NANDN U11227 ( .A(x[551]), .B(y[551]), .Z(n14480) );
  AND U11228 ( .A(n14476), .B(n14480), .Z(n5929) );
  NANDN U11229 ( .A(y[550]), .B(x[550]), .Z(n14482) );
  NANDN U11230 ( .A(x[550]), .B(y[550]), .Z(n14479) );
  ANDN U11231 ( .B(x[548]), .A(y[548]), .Z(n14485) );
  NANDN U11232 ( .A(x[547]), .B(y[547]), .Z(n14487) );
  NANDN U11233 ( .A(x[546]), .B(y[546]), .Z(n14488) );
  NANDN U11234 ( .A(x[545]), .B(y[545]), .Z(n14491) );
  AND U11235 ( .A(n14488), .B(n14491), .Z(n5917) );
  ANDN U11236 ( .B(x[544]), .A(y[544]), .Z(n14493) );
  NANDN U11237 ( .A(x[544]), .B(y[544]), .Z(n14492) );
  ANDN U11238 ( .B(x[542]), .A(y[542]), .Z(n5911) );
  NANDN U11239 ( .A(x[541]), .B(y[541]), .Z(n14499) );
  NANDN U11240 ( .A(x[540]), .B(y[540]), .Z(n14500) );
  NANDN U11241 ( .A(x[539]), .B(y[539]), .Z(n14503) );
  AND U11242 ( .A(n14500), .B(n14503), .Z(n5904) );
  ANDN U11243 ( .B(x[538]), .A(y[538]), .Z(n14505) );
  NANDN U11244 ( .A(x[538]), .B(y[538]), .Z(n14504) );
  NANDN U11245 ( .A(y[536]), .B(x[536]), .Z(n14510) );
  NANDN U11246 ( .A(x[535]), .B(y[535]), .Z(n14511) );
  NANDN U11247 ( .A(x[533]), .B(y[533]), .Z(n14515) );
  XNOR U11248 ( .A(x[534]), .B(y[534]), .Z(n14514) );
  AND U11249 ( .A(n14515), .B(n14514), .Z(n5891) );
  NANDN U11250 ( .A(y[532]), .B(x[532]), .Z(n14518) );
  NANDN U11251 ( .A(x[532]), .B(y[532]), .Z(n14516) );
  ANDN U11252 ( .B(x[530]), .A(y[530]), .Z(n14521) );
  NANDN U11253 ( .A(x[529]), .B(y[529]), .Z(n14523) );
  NANDN U11254 ( .A(x[528]), .B(y[528]), .Z(n14524) );
  NANDN U11255 ( .A(x[527]), .B(y[527]), .Z(n14527) );
  AND U11256 ( .A(n14524), .B(n14527), .Z(n5878) );
  NANDN U11257 ( .A(y[526]), .B(x[526]), .Z(n14530) );
  NANDN U11258 ( .A(x[526]), .B(y[526]), .Z(n14528) );
  ANDN U11259 ( .B(x[524]), .A(y[524]), .Z(n14533) );
  NANDN U11260 ( .A(x[523]), .B(y[523]), .Z(n14535) );
  NANDN U11261 ( .A(x[522]), .B(y[522]), .Z(n14536) );
  NANDN U11262 ( .A(x[521]), .B(y[521]), .Z(n14540) );
  AND U11263 ( .A(n14536), .B(n14540), .Z(n5865) );
  NANDN U11264 ( .A(y[520]), .B(x[520]), .Z(n14542) );
  NANDN U11265 ( .A(x[520]), .B(y[520]), .Z(n14539) );
  ANDN U11266 ( .B(x[518]), .A(y[518]), .Z(n5859) );
  NANDN U11267 ( .A(x[517]), .B(y[517]), .Z(n14547) );
  NANDN U11268 ( .A(x[516]), .B(y[516]), .Z(n14548) );
  NANDN U11269 ( .A(x[515]), .B(y[515]), .Z(n14552) );
  AND U11270 ( .A(n14548), .B(n14552), .Z(n5852) );
  NANDN U11271 ( .A(y[514]), .B(x[514]), .Z(n14554) );
  NANDN U11272 ( .A(x[514]), .B(y[514]), .Z(n14551) );
  NANDN U11273 ( .A(y[512]), .B(x[512]), .Z(n14558) );
  NANDN U11274 ( .A(x[511]), .B(y[511]), .Z(n14559) );
  NANDN U11275 ( .A(x[510]), .B(y[510]), .Z(n14560) );
  NANDN U11276 ( .A(x[509]), .B(y[509]), .Z(n14563) );
  AND U11277 ( .A(n14560), .B(n14563), .Z(n5839) );
  ANDN U11278 ( .B(x[508]), .A(y[508]), .Z(n16012) );
  NANDN U11279 ( .A(x[507]), .B(y[507]), .Z(n14565) );
  ANDN U11280 ( .B(x[506]), .A(y[506]), .Z(n14567) );
  NANDN U11281 ( .A(x[505]), .B(y[505]), .Z(n14569) );
  NANDN U11282 ( .A(x[504]), .B(y[504]), .Z(n14570) );
  NANDN U11283 ( .A(x[503]), .B(y[503]), .Z(n14574) );
  AND U11284 ( .A(n14570), .B(n14574), .Z(n5827) );
  NANDN U11285 ( .A(y[502]), .B(x[502]), .Z(n14576) );
  NANDN U11286 ( .A(x[502]), .B(y[502]), .Z(n14573) );
  ANDN U11287 ( .B(x[500]), .A(y[500]), .Z(n14579) );
  NANDN U11288 ( .A(x[499]), .B(y[499]), .Z(n14581) );
  NANDN U11289 ( .A(x[498]), .B(y[498]), .Z(n14582) );
  NANDN U11290 ( .A(x[497]), .B(y[497]), .Z(n14585) );
  AND U11291 ( .A(n14582), .B(n14585), .Z(n5815) );
  ANDN U11292 ( .B(x[496]), .A(y[496]), .Z(n14587) );
  NANDN U11293 ( .A(x[496]), .B(y[496]), .Z(n14586) );
  NANDN U11294 ( .A(y[494]), .B(x[494]), .Z(n14592) );
  NANDN U11295 ( .A(x[493]), .B(y[493]), .Z(n14594) );
  NANDN U11296 ( .A(x[492]), .B(y[492]), .Z(n14593) );
  NANDN U11297 ( .A(x[491]), .B(y[491]), .Z(n14597) );
  AND U11298 ( .A(n14593), .B(n14597), .Z(n5803) );
  NANDN U11299 ( .A(y[490]), .B(x[490]), .Z(n14600) );
  NANDN U11300 ( .A(x[490]), .B(y[490]), .Z(n14598) );
  NANDN U11301 ( .A(y[488]), .B(x[488]), .Z(n14605) );
  NANDN U11302 ( .A(x[487]), .B(y[487]), .Z(n14606) );
  NANDN U11303 ( .A(x[486]), .B(y[486]), .Z(n14607) );
  NANDN U11304 ( .A(x[485]), .B(y[485]), .Z(n14610) );
  AND U11305 ( .A(n14607), .B(n14610), .Z(n5790) );
  ANDN U11306 ( .B(x[484]), .A(y[484]), .Z(n14612) );
  NANDN U11307 ( .A(x[484]), .B(y[484]), .Z(n14611) );
  ANDN U11308 ( .B(x[482]), .A(y[482]), .Z(n14616) );
  NANDN U11309 ( .A(x[481]), .B(y[481]), .Z(n14619) );
  NANDN U11310 ( .A(x[480]), .B(y[480]), .Z(n14618) );
  NANDN U11311 ( .A(x[479]), .B(y[479]), .Z(n14623) );
  AND U11312 ( .A(n14618), .B(n14623), .Z(n5778) );
  ANDN U11313 ( .B(x[478]), .A(y[478]), .Z(n14624) );
  NANDN U11314 ( .A(x[478]), .B(y[478]), .Z(n14622) );
  NANDN U11315 ( .A(y[476]), .B(x[476]), .Z(n14629) );
  NANDN U11316 ( .A(x[475]), .B(y[475]), .Z(n14631) );
  NANDN U11317 ( .A(x[474]), .B(y[474]), .Z(n14630) );
  NANDN U11318 ( .A(x[473]), .B(y[473]), .Z(n14634) );
  AND U11319 ( .A(n14630), .B(n14634), .Z(n5766) );
  ANDN U11320 ( .B(x[472]), .A(y[472]), .Z(n14636) );
  NANDN U11321 ( .A(x[472]), .B(y[472]), .Z(n14635) );
  ANDN U11322 ( .B(x[470]), .A(y[470]), .Z(n14640) );
  NANDN U11323 ( .A(x[469]), .B(y[469]), .Z(n14642) );
  NANDN U11324 ( .A(x[468]), .B(y[468]), .Z(n14643) );
  NANDN U11325 ( .A(x[467]), .B(y[467]), .Z(n14647) );
  AND U11326 ( .A(n14643), .B(n14647), .Z(n5754) );
  NANDN U11327 ( .A(y[466]), .B(x[466]), .Z(n14649) );
  NANDN U11328 ( .A(x[466]), .B(y[466]), .Z(n14646) );
  ANDN U11329 ( .B(x[464]), .A(y[464]), .Z(n5748) );
  NANDN U11330 ( .A(x[463]), .B(y[463]), .Z(n14654) );
  NANDN U11331 ( .A(x[462]), .B(y[462]), .Z(n14655) );
  NANDN U11332 ( .A(x[461]), .B(y[461]), .Z(n14658) );
  AND U11333 ( .A(n14655), .B(n14658), .Z(n5741) );
  ANDN U11334 ( .B(x[460]), .A(y[460]), .Z(n14660) );
  NANDN U11335 ( .A(x[460]), .B(y[460]), .Z(n14659) );
  NANDN U11336 ( .A(y[458]), .B(x[458]), .Z(n14665) );
  NANDN U11337 ( .A(x[457]), .B(y[457]), .Z(n14666) );
  NANDN U11338 ( .A(x[456]), .B(y[456]), .Z(n14667) );
  NANDN U11339 ( .A(x[455]), .B(y[455]), .Z(n14671) );
  AND U11340 ( .A(n14667), .B(n14671), .Z(n5728) );
  NANDN U11341 ( .A(y[454]), .B(x[454]), .Z(n14673) );
  NANDN U11342 ( .A(x[454]), .B(y[454]), .Z(n14670) );
  NANDN U11343 ( .A(y[452]), .B(x[452]), .Z(n14677) );
  NANDN U11344 ( .A(x[451]), .B(y[451]), .Z(n14678) );
  NANDN U11345 ( .A(x[450]), .B(y[450]), .Z(n14679) );
  NANDN U11346 ( .A(x[449]), .B(y[449]), .Z(n14683) );
  AND U11347 ( .A(n14679), .B(n14683), .Z(n5715) );
  NANDN U11348 ( .A(y[448]), .B(x[448]), .Z(n14685) );
  NANDN U11349 ( .A(x[448]), .B(y[448]), .Z(n14682) );
  ANDN U11350 ( .B(x[446]), .A(y[446]), .Z(n14688) );
  NANDN U11351 ( .A(x[445]), .B(y[445]), .Z(n14690) );
  NANDN U11352 ( .A(x[444]), .B(y[444]), .Z(n14691) );
  NANDN U11353 ( .A(x[443]), .B(y[443]), .Z(n14694) );
  AND U11354 ( .A(n14691), .B(n14694), .Z(n5703) );
  NANDN U11355 ( .A(x[442]), .B(y[442]), .Z(n14695) );
  ANDN U11356 ( .B(x[442]), .A(y[442]), .Z(n14696) );
  ANDN U11357 ( .B(x[440]), .A(y[440]), .Z(n14700) );
  NANDN U11358 ( .A(x[439]), .B(y[439]), .Z(n14702) );
  NANDN U11359 ( .A(x[438]), .B(y[438]), .Z(n14703) );
  NANDN U11360 ( .A(x[437]), .B(y[437]), .Z(n14706) );
  AND U11361 ( .A(n14703), .B(n14706), .Z(n5690) );
  ANDN U11362 ( .B(x[436]), .A(y[436]), .Z(n14708) );
  NANDN U11363 ( .A(x[436]), .B(y[436]), .Z(n14707) );
  ANDN U11364 ( .B(x[434]), .A(y[434]), .Z(n5684) );
  NANDN U11365 ( .A(x[433]), .B(y[433]), .Z(n14714) );
  ANDN U11366 ( .B(x[433]), .A(y[433]), .Z(n14713) );
  NANDN U11367 ( .A(y[431]), .B(x[431]), .Z(n4723) );
  NANDN U11368 ( .A(y[432]), .B(x[432]), .Z(n4722) );
  NAND U11369 ( .A(n4723), .B(n4722), .Z(n25381) );
  NANDN U11370 ( .A(x[431]), .B(y[431]), .Z(n4725) );
  NANDN U11371 ( .A(x[430]), .B(y[430]), .Z(n4724) );
  AND U11372 ( .A(n4725), .B(n4724), .Z(n25379) );
  NANDN U11373 ( .A(x[429]), .B(y[429]), .Z(n14716) );
  ANDN U11374 ( .B(x[428]), .A(y[428]), .Z(n5671) );
  NANDN U11375 ( .A(x[427]), .B(y[427]), .Z(n14720) );
  NANDN U11376 ( .A(x[426]), .B(y[426]), .Z(n14721) );
  NANDN U11377 ( .A(x[425]), .B(y[425]), .Z(n14724) );
  AND U11378 ( .A(n14721), .B(n14724), .Z(n5664) );
  NANDN U11379 ( .A(y[424]), .B(x[424]), .Z(n14727) );
  NANDN U11380 ( .A(x[424]), .B(y[424]), .Z(n14725) );
  NANDN U11381 ( .A(y[422]), .B(x[422]), .Z(n14731) );
  ANDN U11382 ( .B(x[421]), .A(y[421]), .Z(n14730) );
  NANDN U11383 ( .A(x[421]), .B(y[421]), .Z(n4727) );
  NANDN U11384 ( .A(x[420]), .B(y[420]), .Z(n4726) );
  AND U11385 ( .A(n4727), .B(n4726), .Z(n25359) );
  NANDN U11386 ( .A(x[419]), .B(y[419]), .Z(n14733) );
  NANDN U11387 ( .A(y[418]), .B(x[418]), .Z(n14735) );
  XNOR U11388 ( .A(x[418]), .B(y[418]), .Z(n5648) );
  NANDN U11389 ( .A(x[417]), .B(y[417]), .Z(n14736) );
  ANDN U11390 ( .B(x[416]), .A(y[416]), .Z(n5645) );
  NANDN U11391 ( .A(x[415]), .B(y[415]), .Z(n14740) );
  NANDN U11392 ( .A(x[414]), .B(y[414]), .Z(n14741) );
  NANDN U11393 ( .A(x[413]), .B(y[413]), .Z(n14744) );
  AND U11394 ( .A(n14741), .B(n14744), .Z(n5638) );
  ANDN U11395 ( .B(x[412]), .A(y[412]), .Z(n14746) );
  NANDN U11396 ( .A(x[412]), .B(y[412]), .Z(n14745) );
  ANDN U11397 ( .B(x[410]), .A(y[410]), .Z(n5632) );
  NANDN U11398 ( .A(x[409]), .B(y[409]), .Z(n14753) );
  NANDN U11399 ( .A(x[408]), .B(y[408]), .Z(n14752) );
  NANDN U11400 ( .A(x[407]), .B(y[407]), .Z(n14756) );
  AND U11401 ( .A(n14752), .B(n14756), .Z(n5625) );
  ANDN U11402 ( .B(x[406]), .A(y[406]), .Z(n14758) );
  NANDN U11403 ( .A(x[406]), .B(y[406]), .Z(n14757) );
  ANDN U11404 ( .B(x[404]), .A(y[404]), .Z(n14762) );
  NANDN U11405 ( .A(x[403]), .B(y[403]), .Z(n14764) );
  NANDN U11406 ( .A(x[402]), .B(y[402]), .Z(n14765) );
  ANDN U11407 ( .B(x[401]), .A(y[401]), .Z(n14767) );
  NANDN U11408 ( .A(x[401]), .B(y[401]), .Z(n4729) );
  NANDN U11409 ( .A(x[400]), .B(y[400]), .Z(n4728) );
  AND U11410 ( .A(n4729), .B(n4728), .Z(n25319) );
  NANDN U11411 ( .A(y[399]), .B(x[399]), .Z(n4731) );
  NANDN U11412 ( .A(y[400]), .B(x[400]), .Z(n4730) );
  NAND U11413 ( .A(n4731), .B(n4730), .Z(n25317) );
  NANDN U11414 ( .A(x[399]), .B(y[399]), .Z(n4733) );
  NANDN U11415 ( .A(x[398]), .B(y[398]), .Z(n4732) );
  AND U11416 ( .A(n4733), .B(n4732), .Z(n25315) );
  NANDN U11417 ( .A(y[397]), .B(x[397]), .Z(n4735) );
  NANDN U11418 ( .A(y[398]), .B(x[398]), .Z(n4734) );
  NAND U11419 ( .A(n4735), .B(n4734), .Z(n25313) );
  NANDN U11420 ( .A(x[397]), .B(y[397]), .Z(n4737) );
  NANDN U11421 ( .A(x[396]), .B(y[396]), .Z(n4736) );
  AND U11422 ( .A(n4737), .B(n4736), .Z(n25311) );
  NANDN U11423 ( .A(y[395]), .B(x[395]), .Z(n4739) );
  NANDN U11424 ( .A(y[396]), .B(x[396]), .Z(n4738) );
  NAND U11425 ( .A(n4739), .B(n4738), .Z(n25309) );
  NANDN U11426 ( .A(x[395]), .B(y[395]), .Z(n4741) );
  NANDN U11427 ( .A(x[394]), .B(y[394]), .Z(n4740) );
  AND U11428 ( .A(n4741), .B(n4740), .Z(n25307) );
  NANDN U11429 ( .A(y[393]), .B(x[393]), .Z(n4743) );
  NANDN U11430 ( .A(y[394]), .B(x[394]), .Z(n4742) );
  NAND U11431 ( .A(n4743), .B(n4742), .Z(n25305) );
  NANDN U11432 ( .A(x[393]), .B(y[393]), .Z(n4745) );
  NANDN U11433 ( .A(x[392]), .B(y[392]), .Z(n4744) );
  AND U11434 ( .A(n4745), .B(n4744), .Z(n25303) );
  NANDN U11435 ( .A(x[391]), .B(y[391]), .Z(n14769) );
  NANDN U11436 ( .A(y[390]), .B(x[390]), .Z(n14771) );
  XNOR U11437 ( .A(x[390]), .B(y[390]), .Z(n5596) );
  NANDN U11438 ( .A(x[389]), .B(y[389]), .Z(n14773) );
  NANDN U11439 ( .A(y[388]), .B(x[388]), .Z(n14775) );
  NANDN U11440 ( .A(x[387]), .B(y[387]), .Z(n14776) );
  NANDN U11441 ( .A(x[386]), .B(y[386]), .Z(n14777) );
  NANDN U11442 ( .A(x[385]), .B(y[385]), .Z(n14781) );
  AND U11443 ( .A(n14777), .B(n14781), .Z(n5587) );
  NANDN U11444 ( .A(y[384]), .B(x[384]), .Z(n14783) );
  NANDN U11445 ( .A(x[384]), .B(y[384]), .Z(n14780) );
  ANDN U11446 ( .B(x[382]), .A(y[382]), .Z(n14786) );
  NANDN U11447 ( .A(x[381]), .B(y[381]), .Z(n14789) );
  NANDN U11448 ( .A(x[380]), .B(y[380]), .Z(n14788) );
  NANDN U11449 ( .A(x[379]), .B(y[379]), .Z(n14793) );
  AND U11450 ( .A(n14788), .B(n14793), .Z(n5575) );
  NANDN U11451 ( .A(y[378]), .B(x[378]), .Z(n14795) );
  NANDN U11452 ( .A(x[378]), .B(y[378]), .Z(n14792) );
  NANDN U11453 ( .A(y[376]), .B(x[376]), .Z(n14798) );
  NANDN U11454 ( .A(x[375]), .B(y[375]), .Z(n14801) );
  NANDN U11455 ( .A(x[374]), .B(y[374]), .Z(n14800) );
  NANDN U11456 ( .A(x[373]), .B(y[373]), .Z(n14804) );
  AND U11457 ( .A(n14800), .B(n14804), .Z(n5563) );
  ANDN U11458 ( .B(x[372]), .A(y[372]), .Z(n14806) );
  NANDN U11459 ( .A(x[372]), .B(y[372]), .Z(n14805) );
  ANDN U11460 ( .B(x[370]), .A(y[370]), .Z(n14810) );
  NANDN U11461 ( .A(x[369]), .B(y[369]), .Z(n14812) );
  NANDN U11462 ( .A(x[368]), .B(y[368]), .Z(n14813) );
  NANDN U11463 ( .A(x[367]), .B(y[367]), .Z(n14816) );
  AND U11464 ( .A(n14813), .B(n14816), .Z(n5550) );
  ANDN U11465 ( .B(x[366]), .A(y[366]), .Z(n14818) );
  NANDN U11466 ( .A(x[366]), .B(y[366]), .Z(n14817) );
  ANDN U11467 ( .B(x[364]), .A(y[364]), .Z(n14822) );
  NANDN U11468 ( .A(x[363]), .B(y[363]), .Z(n14824) );
  NANDN U11469 ( .A(x[362]), .B(y[362]), .Z(n14825) );
  NANDN U11470 ( .A(x[361]), .B(y[361]), .Z(n14828) );
  AND U11471 ( .A(n14825), .B(n14828), .Z(n5537) );
  ANDN U11472 ( .B(x[360]), .A(y[360]), .Z(n5534) );
  NANDN U11473 ( .A(x[360]), .B(y[360]), .Z(n14829) );
  ANDN U11474 ( .B(x[358]), .A(y[358]), .Z(n14834) );
  NANDN U11475 ( .A(x[357]), .B(y[357]), .Z(n14837) );
  NANDN U11476 ( .A(x[356]), .B(y[356]), .Z(n14836) );
  NANDN U11477 ( .A(x[355]), .B(y[355]), .Z(n14840) );
  AND U11478 ( .A(n14836), .B(n14840), .Z(n5524) );
  ANDN U11479 ( .B(x[354]), .A(y[354]), .Z(n5521) );
  NANDN U11480 ( .A(x[354]), .B(y[354]), .Z(n14841) );
  NANDN U11481 ( .A(y[352]), .B(x[352]), .Z(n15854) );
  NANDN U11482 ( .A(x[350]), .B(y[350]), .Z(n15851) );
  NANDN U11483 ( .A(x[349]), .B(y[349]), .Z(n14848) );
  AND U11484 ( .A(n15851), .B(n14848), .Z(n5511) );
  NANDN U11485 ( .A(y[348]), .B(x[348]), .Z(n14851) );
  NANDN U11486 ( .A(x[348]), .B(y[348]), .Z(n14849) );
  NANDN U11487 ( .A(y[346]), .B(x[346]), .Z(n14855) );
  NANDN U11488 ( .A(x[345]), .B(y[345]), .Z(n14857) );
  NANDN U11489 ( .A(x[344]), .B(y[344]), .Z(n14856) );
  NANDN U11490 ( .A(x[343]), .B(y[343]), .Z(n14860) );
  AND U11491 ( .A(n14856), .B(n14860), .Z(n5499) );
  NANDN U11492 ( .A(y[342]), .B(x[342]), .Z(n14863) );
  NANDN U11493 ( .A(x[342]), .B(y[342]), .Z(n14861) );
  NANDN U11494 ( .A(x[341]), .B(y[341]), .Z(n4747) );
  NANDN U11495 ( .A(x[340]), .B(y[340]), .Z(n4746) );
  AND U11496 ( .A(n4747), .B(n4746), .Z(n25215) );
  NANDN U11497 ( .A(y[339]), .B(x[339]), .Z(n4749) );
  NANDN U11498 ( .A(y[340]), .B(x[340]), .Z(n4748) );
  NAND U11499 ( .A(n4749), .B(n4748), .Z(n25213) );
  NANDN U11500 ( .A(x[339]), .B(y[339]), .Z(n4751) );
  NANDN U11501 ( .A(x[338]), .B(y[338]), .Z(n4750) );
  AND U11502 ( .A(n4751), .B(n4750), .Z(n25211) );
  NANDN U11503 ( .A(y[336]), .B(x[336]), .Z(n14867) );
  ANDN U11504 ( .B(y[335]), .A(x[335]), .Z(n14868) );
  NANDN U11505 ( .A(y[334]), .B(x[334]), .Z(n14870) );
  NANDN U11506 ( .A(y[333]), .B(x[333]), .Z(n14871) );
  NANDN U11507 ( .A(y[332]), .B(x[332]), .Z(n14874) );
  AND U11508 ( .A(n14871), .B(n14874), .Z(n5478) );
  ANDN U11509 ( .B(y[331]), .A(x[331]), .Z(n14876) );
  NANDN U11510 ( .A(y[331]), .B(x[331]), .Z(n14875) );
  ANDN U11511 ( .B(y[329]), .A(x[329]), .Z(n14880) );
  NANDN U11512 ( .A(y[328]), .B(x[328]), .Z(n14882) );
  NANDN U11513 ( .A(y[327]), .B(x[327]), .Z(n14883) );
  NANDN U11514 ( .A(y[326]), .B(x[326]), .Z(n14887) );
  AND U11515 ( .A(n14883), .B(n14887), .Z(n5466) );
  ANDN U11516 ( .B(y[325]), .A(x[325]), .Z(n14888) );
  NANDN U11517 ( .A(y[325]), .B(x[325]), .Z(n14886) );
  XOR U11518 ( .A(x[324]), .B(y[324]), .Z(n14889) );
  NANDN U11519 ( .A(y[322]), .B(x[322]), .Z(n14893) );
  NANDN U11520 ( .A(y[321]), .B(x[321]), .Z(n14894) );
  NANDN U11521 ( .A(y[320]), .B(x[320]), .Z(n4752) );
  AND U11522 ( .A(n14894), .B(n4752), .Z(n5453) );
  ANDN U11523 ( .B(y[319]), .A(x[319]), .Z(n14898) );
  NANDN U11524 ( .A(y[319]), .B(x[319]), .Z(n14897) );
  XOR U11525 ( .A(x[318]), .B(y[318]), .Z(n14899) );
  NANDN U11526 ( .A(y[316]), .B(x[316]), .Z(n14903) );
  NANDN U11527 ( .A(y[315]), .B(x[315]), .Z(n14904) );
  NANDN U11528 ( .A(y[314]), .B(x[314]), .Z(n14907) );
  AND U11529 ( .A(n14904), .B(n14907), .Z(n5440) );
  ANDN U11530 ( .B(y[313]), .A(x[313]), .Z(n14909) );
  NANDN U11531 ( .A(y[313]), .B(x[313]), .Z(n14908) );
  NANDN U11532 ( .A(x[311]), .B(y[311]), .Z(n14915) );
  NANDN U11533 ( .A(y[310]), .B(x[310]), .Z(n14916) );
  NANDN U11534 ( .A(y[309]), .B(x[309]), .Z(n14917) );
  NANDN U11535 ( .A(y[308]), .B(x[308]), .Z(n4753) );
  AND U11536 ( .A(n14917), .B(n4753), .Z(n5428) );
  ANDN U11537 ( .B(y[307]), .A(x[307]), .Z(n14923) );
  NANDN U11538 ( .A(y[307]), .B(x[307]), .Z(n14920) );
  ANDN U11539 ( .B(y[305]), .A(x[305]), .Z(n14927) );
  NANDN U11540 ( .A(y[305]), .B(x[305]), .Z(n14926) );
  NANDN U11541 ( .A(y[304]), .B(x[304]), .Z(n14929) );
  NANDN U11542 ( .A(y[303]), .B(x[303]), .Z(n14930) );
  NANDN U11543 ( .A(y[302]), .B(x[302]), .Z(n4754) );
  AND U11544 ( .A(n14930), .B(n4754), .Z(n5415) );
  NANDN U11545 ( .A(x[301]), .B(y[301]), .Z(n14935) );
  NANDN U11546 ( .A(y[301]), .B(x[301]), .Z(n14933) );
  NANDN U11547 ( .A(x[299]), .B(y[299]), .Z(n14939) );
  NANDN U11548 ( .A(y[298]), .B(x[298]), .Z(n14940) );
  NANDN U11549 ( .A(y[297]), .B(x[297]), .Z(n14941) );
  NANDN U11550 ( .A(y[296]), .B(x[296]), .Z(n4755) );
  AND U11551 ( .A(n14941), .B(n4755), .Z(n5403) );
  NANDN U11552 ( .A(x[295]), .B(y[295]), .Z(n14946) );
  NANDN U11553 ( .A(y[295]), .B(x[295]), .Z(n14944) );
  NANDN U11554 ( .A(x[293]), .B(y[293]), .Z(n14950) );
  NANDN U11555 ( .A(y[292]), .B(x[292]), .Z(n14952) );
  NANDN U11556 ( .A(y[291]), .B(x[291]), .Z(n14951) );
  NANDN U11557 ( .A(y[290]), .B(x[290]), .Z(n14955) );
  AND U11558 ( .A(n14951), .B(n14955), .Z(n5391) );
  ANDN U11559 ( .B(y[289]), .A(x[289]), .Z(n14957) );
  NANDN U11560 ( .A(y[289]), .B(x[289]), .Z(n14956) );
  ANDN U11561 ( .B(y[287]), .A(x[287]), .Z(n14962) );
  NANDN U11562 ( .A(y[287]), .B(x[287]), .Z(n14959) );
  NANDN U11563 ( .A(y[286]), .B(x[286]), .Z(n14966) );
  NANDN U11564 ( .A(y[285]), .B(x[285]), .Z(n14965) );
  NANDN U11565 ( .A(y[284]), .B(x[284]), .Z(n14970) );
  AND U11566 ( .A(n14965), .B(n14970), .Z(n5378) );
  ANDN U11567 ( .B(y[283]), .A(x[283]), .Z(n14971) );
  NANDN U11568 ( .A(y[283]), .B(x[283]), .Z(n14969) );
  ANDN U11569 ( .B(y[281]), .A(x[281]), .Z(n14975) );
  NANDN U11570 ( .A(y[280]), .B(x[280]), .Z(n14978) );
  NANDN U11571 ( .A(y[279]), .B(x[279]), .Z(n14977) );
  NANDN U11572 ( .A(y[278]), .B(x[278]), .Z(n4756) );
  AND U11573 ( .A(n14977), .B(n4756), .Z(n5366) );
  NANDN U11574 ( .A(x[277]), .B(y[277]), .Z(n14983) );
  NANDN U11575 ( .A(y[277]), .B(x[277]), .Z(n14981) );
  ANDN U11576 ( .B(y[275]), .A(x[275]), .Z(n14986) );
  NANDN U11577 ( .A(y[274]), .B(x[274]), .Z(n14989) );
  NANDN U11578 ( .A(y[273]), .B(x[273]), .Z(n14988) );
  NANDN U11579 ( .A(y[272]), .B(x[272]), .Z(n14993) );
  AND U11580 ( .A(n14988), .B(n14993), .Z(n5354) );
  NANDN U11581 ( .A(y[271]), .B(x[271]), .Z(n14992) );
  NANDN U11582 ( .A(x[270]), .B(y[270]), .Z(n4758) );
  NANDN U11583 ( .A(x[271]), .B(y[271]), .Z(n4757) );
  NAND U11584 ( .A(n4758), .B(n4757), .Z(n14994) );
  NANDN U11585 ( .A(y[270]), .B(x[270]), .Z(n4760) );
  NANDN U11586 ( .A(y[269]), .B(x[269]), .Z(n4759) );
  AND U11587 ( .A(n4760), .B(n4759), .Z(n15768) );
  NANDN U11588 ( .A(x[268]), .B(y[268]), .Z(n4762) );
  NANDN U11589 ( .A(x[269]), .B(y[269]), .Z(n4761) );
  NAND U11590 ( .A(n4762), .B(n4761), .Z(n15766) );
  NANDN U11591 ( .A(y[268]), .B(x[268]), .Z(n4764) );
  NANDN U11592 ( .A(y[267]), .B(x[267]), .Z(n4763) );
  AND U11593 ( .A(n4764), .B(n4763), .Z(n14995) );
  NANDN U11594 ( .A(x[264]), .B(y[264]), .Z(n4766) );
  NANDN U11595 ( .A(x[265]), .B(y[265]), .Z(n4765) );
  NAND U11596 ( .A(n4766), .B(n4765), .Z(n14998) );
  NANDN U11597 ( .A(y[264]), .B(x[264]), .Z(n4768) );
  NANDN U11598 ( .A(y[263]), .B(x[263]), .Z(n4767) );
  AND U11599 ( .A(n4768), .B(n4767), .Z(n15760) );
  ANDN U11600 ( .B(y[261]), .A(x[261]), .Z(n15002) );
  NANDN U11601 ( .A(y[261]), .B(x[261]), .Z(n15000) );
  ANDN U11602 ( .B(y[259]), .A(x[259]), .Z(n15005) );
  NANDN U11603 ( .A(y[259]), .B(x[259]), .Z(n15004) );
  NANDN U11604 ( .A(y[258]), .B(x[258]), .Z(n15008) );
  NANDN U11605 ( .A(y[257]), .B(x[257]), .Z(n15007) );
  NANDN U11606 ( .A(y[256]), .B(x[256]), .Z(n15012) );
  AND U11607 ( .A(n15007), .B(n15012), .Z(n5323) );
  ANDN U11608 ( .B(y[255]), .A(x[255]), .Z(n15013) );
  NANDN U11609 ( .A(y[255]), .B(x[255]), .Z(n15011) );
  ANDN U11610 ( .B(y[253]), .A(x[253]), .Z(n15016) );
  NANDN U11611 ( .A(y[253]), .B(x[253]), .Z(n15015) );
  NANDN U11612 ( .A(y[252]), .B(x[252]), .Z(n15019) );
  NANDN U11613 ( .A(y[251]), .B(x[251]), .Z(n15018) );
  NANDN U11614 ( .A(y[250]), .B(x[250]), .Z(n15023) );
  AND U11615 ( .A(n15018), .B(n15023), .Z(n5310) );
  NANDN U11616 ( .A(x[249]), .B(y[249]), .Z(n15025) );
  NANDN U11617 ( .A(y[249]), .B(x[249]), .Z(n15022) );
  NANDN U11618 ( .A(x[247]), .B(y[247]), .Z(n15029) );
  NANDN U11619 ( .A(y[246]), .B(x[246]), .Z(n15031) );
  NANDN U11620 ( .A(y[245]), .B(x[245]), .Z(n15030) );
  NANDN U11621 ( .A(y[244]), .B(x[244]), .Z(n15034) );
  AND U11622 ( .A(n15030), .B(n15034), .Z(n5298) );
  ANDN U11623 ( .B(y[243]), .A(x[243]), .Z(n15036) );
  NANDN U11624 ( .A(y[243]), .B(x[243]), .Z(n15035) );
  NANDN U11625 ( .A(x[241]), .B(y[241]), .Z(n15040) );
  NANDN U11626 ( .A(y[241]), .B(x[241]), .Z(n15038) );
  NANDN U11627 ( .A(y[240]), .B(x[240]), .Z(n15041) );
  NANDN U11628 ( .A(y[239]), .B(x[239]), .Z(n15042) );
  NANDN U11629 ( .A(y[238]), .B(x[238]), .Z(n15046) );
  AND U11630 ( .A(n15042), .B(n15046), .Z(n5285) );
  ANDN U11631 ( .B(y[237]), .A(x[237]), .Z(n15047) );
  NANDN U11632 ( .A(y[237]), .B(x[237]), .Z(n15045) );
  ANDN U11633 ( .B(y[235]), .A(x[235]), .Z(n15051) );
  NANDN U11634 ( .A(y[234]), .B(x[234]), .Z(n15054) );
  NANDN U11635 ( .A(y[233]), .B(x[233]), .Z(n15053) );
  NANDN U11636 ( .A(y[232]), .B(x[232]), .Z(n15057) );
  AND U11637 ( .A(n15053), .B(n15057), .Z(n5273) );
  ANDN U11638 ( .B(y[231]), .A(x[231]), .Z(n15059) );
  NANDN U11639 ( .A(y[231]), .B(x[231]), .Z(n15058) );
  ANDN U11640 ( .B(y[229]), .A(x[229]), .Z(n15062) );
  NANDN U11641 ( .A(y[229]), .B(x[229]), .Z(n15061) );
  NANDN U11642 ( .A(y[228]), .B(x[228]), .Z(n15064) );
  NANDN U11643 ( .A(y[227]), .B(x[227]), .Z(n15065) );
  NANDN U11644 ( .A(y[226]), .B(x[226]), .Z(n15070) );
  AND U11645 ( .A(n15065), .B(n15070), .Z(n5260) );
  NANDN U11646 ( .A(x[225]), .B(y[225]), .Z(n15072) );
  NANDN U11647 ( .A(y[225]), .B(x[225]), .Z(n15069) );
  NANDN U11648 ( .A(x[223]), .B(y[223]), .Z(n15076) );
  NANDN U11649 ( .A(y[222]), .B(x[222]), .Z(n15078) );
  NANDN U11650 ( .A(y[221]), .B(x[221]), .Z(n15077) );
  NANDN U11651 ( .A(y[220]), .B(x[220]), .Z(n15082) );
  AND U11652 ( .A(n15077), .B(n15082), .Z(n5248) );
  ANDN U11653 ( .B(y[219]), .A(x[219]), .Z(n15083) );
  NANDN U11654 ( .A(y[219]), .B(x[219]), .Z(n15081) );
  ANDN U11655 ( .B(y[217]), .A(x[217]), .Z(n15087) );
  NANDN U11656 ( .A(y[216]), .B(x[216]), .Z(n15089) );
  NANDN U11657 ( .A(y[215]), .B(x[215]), .Z(n15090) );
  NANDN U11658 ( .A(y[214]), .B(x[214]), .Z(n15093) );
  AND U11659 ( .A(n15090), .B(n15093), .Z(n5236) );
  ANDN U11660 ( .B(y[213]), .A(x[213]), .Z(n15095) );
  NANDN U11661 ( .A(y[213]), .B(x[213]), .Z(n15094) );
  ANDN U11662 ( .B(y[211]), .A(x[211]), .Z(n15099) );
  NANDN U11663 ( .A(y[210]), .B(x[210]), .Z(n5227) );
  NANDN U11664 ( .A(y[208]), .B(x[208]), .Z(n15105) );
  NANDN U11665 ( .A(y[209]), .B(x[209]), .Z(n15101) );
  AND U11666 ( .A(n15105), .B(n15101), .Z(n5223) );
  NANDN U11667 ( .A(x[207]), .B(y[207]), .Z(n15108) );
  NANDN U11668 ( .A(y[207]), .B(x[207]), .Z(n15104) );
  ANDN U11669 ( .B(y[205]), .A(x[205]), .Z(n15111) );
  NANDN U11670 ( .A(y[204]), .B(x[204]), .Z(n15113) );
  NANDN U11671 ( .A(y[203]), .B(x[203]), .Z(n15114) );
  NANDN U11672 ( .A(y[202]), .B(x[202]), .Z(n15117) );
  AND U11673 ( .A(n15114), .B(n15117), .Z(n5211) );
  ANDN U11674 ( .B(y[201]), .A(x[201]), .Z(n15119) );
  NANDN U11675 ( .A(y[201]), .B(x[201]), .Z(n15118) );
  ANDN U11676 ( .B(y[199]), .A(x[199]), .Z(n15123) );
  NANDN U11677 ( .A(y[198]), .B(x[198]), .Z(n5202) );
  NANDN U11678 ( .A(y[196]), .B(x[196]), .Z(n15129) );
  NANDN U11679 ( .A(y[197]), .B(x[197]), .Z(n15125) );
  AND U11680 ( .A(n15129), .B(n15125), .Z(n5198) );
  ANDN U11681 ( .B(y[195]), .A(x[195]), .Z(n15130) );
  NANDN U11682 ( .A(y[195]), .B(x[195]), .Z(n15128) );
  ANDN U11683 ( .B(y[193]), .A(x[193]), .Z(n15134) );
  NANDN U11684 ( .A(y[192]), .B(x[192]), .Z(n15136) );
  NANDN U11685 ( .A(y[191]), .B(x[191]), .Z(n15137) );
  NANDN U11686 ( .A(y[190]), .B(x[190]), .Z(n15141) );
  AND U11687 ( .A(n15137), .B(n15141), .Z(n5186) );
  NANDN U11688 ( .A(x[189]), .B(y[189]), .Z(n15143) );
  NANDN U11689 ( .A(y[189]), .B(x[189]), .Z(n15140) );
  NANDN U11690 ( .A(x[187]), .B(y[187]), .Z(n15148) );
  NANDN U11691 ( .A(y[186]), .B(x[186]), .Z(n15149) );
  NANDN U11692 ( .A(y[185]), .B(x[185]), .Z(n15150) );
  NANDN U11693 ( .A(y[184]), .B(x[184]), .Z(n15153) );
  AND U11694 ( .A(n15150), .B(n15153), .Z(n5174) );
  ANDN U11695 ( .B(y[183]), .A(x[183]), .Z(n15155) );
  NANDN U11696 ( .A(y[183]), .B(x[183]), .Z(n15154) );
  ANDN U11697 ( .B(y[181]), .A(x[181]), .Z(n15158) );
  NANDN U11698 ( .A(y[181]), .B(x[181]), .Z(n15157) );
  NANDN U11699 ( .A(y[180]), .B(x[180]), .Z(n5164) );
  NANDN U11700 ( .A(y[178]), .B(x[178]), .Z(n15164) );
  NANDN U11701 ( .A(y[179]), .B(x[179]), .Z(n15160) );
  AND U11702 ( .A(n15164), .B(n15160), .Z(n5160) );
  ANDN U11703 ( .B(y[177]), .A(x[177]), .Z(n15165) );
  NANDN U11704 ( .A(y[177]), .B(x[177]), .Z(n15163) );
  ANDN U11705 ( .B(y[175]), .A(x[175]), .Z(n15170) );
  NANDN U11706 ( .A(y[175]), .B(x[175]), .Z(n15167) );
  NANDN U11707 ( .A(y[174]), .B(x[174]), .Z(n5150) );
  NANDN U11708 ( .A(y[172]), .B(x[172]), .Z(n15179) );
  NANDN U11709 ( .A(y[173]), .B(x[173]), .Z(n15173) );
  AND U11710 ( .A(n15179), .B(n15173), .Z(n5146) );
  ANDN U11711 ( .B(y[171]), .A(x[171]), .Z(n15181) );
  NANDN U11712 ( .A(y[171]), .B(x[171]), .Z(n15180) );
  XOR U11713 ( .A(x[170]), .B(y[170]), .Z(n15182) );
  NANDN U11714 ( .A(y[168]), .B(x[168]), .Z(n15186) );
  NANDN U11715 ( .A(y[167]), .B(x[167]), .Z(n15187) );
  NANDN U11716 ( .A(y[166]), .B(x[166]), .Z(n15191) );
  AND U11717 ( .A(n15187), .B(n15191), .Z(n5133) );
  ANDN U11718 ( .B(y[165]), .A(x[165]), .Z(n15193) );
  NANDN U11719 ( .A(y[165]), .B(x[165]), .Z(n15192) );
  ANDN U11720 ( .B(y[163]), .A(x[163]), .Z(n15197) );
  NANDN U11721 ( .A(y[162]), .B(x[162]), .Z(n15200) );
  NANDN U11722 ( .A(y[161]), .B(x[161]), .Z(n15199) );
  NANDN U11723 ( .A(y[160]), .B(x[160]), .Z(n15204) );
  AND U11724 ( .A(n15199), .B(n15204), .Z(n5121) );
  NANDN U11725 ( .A(x[159]), .B(y[159]), .Z(n15206) );
  NANDN U11726 ( .A(y[159]), .B(x[159]), .Z(n15203) );
  NANDN U11727 ( .A(x[157]), .B(y[157]), .Z(n15210) );
  NANDN U11728 ( .A(y[156]), .B(x[156]), .Z(n15211) );
  NANDN U11729 ( .A(y[155]), .B(x[155]), .Z(n15212) );
  NANDN U11730 ( .A(y[154]), .B(x[154]), .Z(n15216) );
  AND U11731 ( .A(n15212), .B(n15216), .Z(n5109) );
  ANDN U11732 ( .B(y[153]), .A(x[153]), .Z(n15217) );
  NANDN U11733 ( .A(y[153]), .B(x[153]), .Z(n15215) );
  ANDN U11734 ( .B(y[151]), .A(x[151]), .Z(n15221) );
  NANDN U11735 ( .A(y[150]), .B(x[150]), .Z(n5100) );
  NANDN U11736 ( .A(y[148]), .B(x[148]), .Z(n15227) );
  NANDN U11737 ( .A(y[149]), .B(x[149]), .Z(n15223) );
  AND U11738 ( .A(n15227), .B(n15223), .Z(n5096) );
  ANDN U11739 ( .B(y[147]), .A(x[147]), .Z(n15228) );
  NANDN U11740 ( .A(y[147]), .B(x[147]), .Z(n15226) );
  ANDN U11741 ( .B(y[145]), .A(x[145]), .Z(n15231) );
  NANDN U11742 ( .A(y[145]), .B(x[145]), .Z(n15230) );
  NANDN U11743 ( .A(x[144]), .B(y[144]), .Z(n15232) );
  NANDN U11744 ( .A(y[144]), .B(x[144]), .Z(n4770) );
  NANDN U11745 ( .A(y[143]), .B(x[143]), .Z(n4769) );
  AND U11746 ( .A(n4770), .B(n4769), .Z(n15639) );
  NANDN U11747 ( .A(y[142]), .B(x[142]), .Z(n15234) );
  NANDN U11748 ( .A(x[141]), .B(y[141]), .Z(n15236) );
  XNOR U11749 ( .A(y[141]), .B(x[141]), .Z(n5079) );
  NANDN U11750 ( .A(y[140]), .B(x[140]), .Z(n15237) );
  NANDN U11751 ( .A(y[139]), .B(x[139]), .Z(n15238) );
  NANDN U11752 ( .A(y[138]), .B(x[138]), .Z(n15242) );
  AND U11753 ( .A(n15238), .B(n15242), .Z(n5074) );
  ANDN U11754 ( .B(y[137]), .A(x[137]), .Z(n15243) );
  NANDN U11755 ( .A(y[137]), .B(x[137]), .Z(n15241) );
  NANDN U11756 ( .A(x[135]), .B(y[135]), .Z(n15248) );
  NANDN U11757 ( .A(y[134]), .B(x[134]), .Z(n15249) );
  NANDN U11758 ( .A(y[133]), .B(x[133]), .Z(n15250) );
  NANDN U11759 ( .A(y[132]), .B(x[132]), .Z(n15254) );
  AND U11760 ( .A(n15250), .B(n15254), .Z(n5062) );
  ANDN U11761 ( .B(y[131]), .A(x[131]), .Z(n15255) );
  NANDN U11762 ( .A(y[131]), .B(x[131]), .Z(n15253) );
  ANDN U11763 ( .B(y[129]), .A(x[129]), .Z(n15259) );
  NANDN U11764 ( .A(y[128]), .B(x[128]), .Z(n5053) );
  NANDN U11765 ( .A(y[126]), .B(x[126]), .Z(n15264) );
  NANDN U11766 ( .A(y[127]), .B(x[127]), .Z(n15261) );
  AND U11767 ( .A(n15264), .B(n15261), .Z(n5049) );
  ANDN U11768 ( .B(y[125]), .A(x[125]), .Z(n15266) );
  NANDN U11769 ( .A(y[125]), .B(x[125]), .Z(n15265) );
  NANDN U11770 ( .A(x[123]), .B(y[123]), .Z(n15271) );
  NANDN U11771 ( .A(y[122]), .B(x[122]), .Z(n15272) );
  NANDN U11772 ( .A(y[121]), .B(x[121]), .Z(n15273) );
  NANDN U11773 ( .A(y[120]), .B(x[120]), .Z(n15276) );
  AND U11774 ( .A(n15273), .B(n15276), .Z(n5037) );
  NANDN U11775 ( .A(x[119]), .B(y[119]), .Z(n15279) );
  NANDN U11776 ( .A(y[119]), .B(x[119]), .Z(n15277) );
  ANDN U11777 ( .B(y[117]), .A(x[117]), .Z(n15282) );
  NANDN U11778 ( .A(y[116]), .B(x[116]), .Z(n15284) );
  NANDN U11779 ( .A(y[115]), .B(x[115]), .Z(n15285) );
  NANDN U11780 ( .A(y[114]), .B(x[114]), .Z(n4771) );
  AND U11781 ( .A(n15285), .B(n4771), .Z(n5025) );
  ANDN U11782 ( .B(y[113]), .A(x[113]), .Z(n15291) );
  NANDN U11783 ( .A(y[113]), .B(x[113]), .Z(n15288) );
  NANDN U11784 ( .A(x[111]), .B(y[111]), .Z(n15297) );
  NANDN U11785 ( .A(y[110]), .B(x[110]), .Z(n15299) );
  NANDN U11786 ( .A(y[109]), .B(x[109]), .Z(n15298) );
  NANDN U11787 ( .A(y[108]), .B(x[108]), .Z(n15302) );
  AND U11788 ( .A(n15298), .B(n15302), .Z(n5013) );
  NANDN U11789 ( .A(x[107]), .B(y[107]), .Z(n15305) );
  NANDN U11790 ( .A(y[107]), .B(x[107]), .Z(n15303) );
  NANDN U11791 ( .A(x[105]), .B(y[105]), .Z(n15309) );
  NANDN U11792 ( .A(y[104]), .B(x[104]), .Z(n15310) );
  NANDN U11793 ( .A(y[103]), .B(x[103]), .Z(n15311) );
  NANDN U11794 ( .A(x[102]), .B(y[102]), .Z(n15313) );
  NANDN U11795 ( .A(y[102]), .B(x[102]), .Z(n4773) );
  NANDN U11796 ( .A(y[101]), .B(x[101]), .Z(n4772) );
  AND U11797 ( .A(n4773), .B(n4772), .Z(n15595) );
  NANDN U11798 ( .A(x[99]), .B(y[99]), .Z(n15317) );
  NANDN U11799 ( .A(y[98]), .B(x[98]), .Z(n15319) );
  NANDN U11800 ( .A(x[97]), .B(y[97]), .Z(n15320) );
  NANDN U11801 ( .A(x[95]), .B(y[95]), .Z(n15325) );
  XNOR U11802 ( .A(x[96]), .B(y[96]), .Z(n15323) );
  AND U11803 ( .A(n15325), .B(n15323), .Z(n4985) );
  ANDN U11804 ( .B(x[94]), .A(y[94]), .Z(n15326) );
  NANDN U11805 ( .A(x[94]), .B(y[94]), .Z(n15324) );
  NANDN U11806 ( .A(y[92]), .B(x[92]), .Z(n15330) );
  NANDN U11807 ( .A(x[91]), .B(y[91]), .Z(n15332) );
  NANDN U11808 ( .A(x[90]), .B(y[90]), .Z(n15333) );
  NANDN U11809 ( .A(x[89]), .B(y[89]), .Z(n15337) );
  AND U11810 ( .A(n15333), .B(n15337), .Z(n4973) );
  NANDN U11811 ( .A(y[88]), .B(x[88]), .Z(n15339) );
  NANDN U11812 ( .A(x[88]), .B(y[88]), .Z(n15336) );
  NANDN U11813 ( .A(y[86]), .B(x[86]), .Z(n15343) );
  NANDN U11814 ( .A(x[85]), .B(y[85]), .Z(n15344) );
  NANDN U11815 ( .A(x[84]), .B(y[84]), .Z(n15345) );
  NANDN U11816 ( .A(x[83]), .B(y[83]), .Z(n15348) );
  AND U11817 ( .A(n15345), .B(n15348), .Z(n4960) );
  NANDN U11818 ( .A(y[82]), .B(x[82]), .Z(n15351) );
  NANDN U11819 ( .A(x[82]), .B(y[82]), .Z(n15349) );
  ANDN U11820 ( .B(x[80]), .A(y[80]), .Z(n4954) );
  ANDN U11821 ( .B(x[79]), .A(y[79]), .Z(n15355) );
  NANDN U11822 ( .A(x[79]), .B(y[79]), .Z(n4775) );
  NANDN U11823 ( .A(x[78]), .B(y[78]), .Z(n4774) );
  AND U11824 ( .A(n4775), .B(n4774), .Z(n24691) );
  NANDN U11825 ( .A(x[77]), .B(y[77]), .Z(n15357) );
  NANDN U11826 ( .A(y[76]), .B(x[76]), .Z(n15359) );
  XNOR U11827 ( .A(x[76]), .B(y[76]), .Z(n4943) );
  NANDN U11828 ( .A(x[75]), .B(y[75]), .Z(n15360) );
  NANDN U11829 ( .A(x[74]), .B(y[74]), .Z(n15361) );
  NANDN U11830 ( .A(x[73]), .B(y[73]), .Z(n15364) );
  AND U11831 ( .A(n15361), .B(n15364), .Z(n4938) );
  NANDN U11832 ( .A(x[72]), .B(y[72]), .Z(n15365) );
  NANDN U11833 ( .A(y[71]), .B(x[71]), .Z(n4777) );
  NANDN U11834 ( .A(y[72]), .B(x[72]), .Z(n4776) );
  NAND U11835 ( .A(n4777), .B(n4776), .Z(n24677) );
  NANDN U11836 ( .A(x[71]), .B(y[71]), .Z(n4779) );
  NANDN U11837 ( .A(x[70]), .B(y[70]), .Z(n4778) );
  AND U11838 ( .A(n4779), .B(n4778), .Z(n24675) );
  NANDN U11839 ( .A(y[68]), .B(x[68]), .Z(n15370) );
  NANDN U11840 ( .A(x[68]), .B(y[68]), .Z(n15367) );
  NANDN U11841 ( .A(y[66]), .B(x[66]), .Z(n15374) );
  ANDN U11842 ( .B(x[65]), .A(y[65]), .Z(n15373) );
  NANDN U11843 ( .A(x[65]), .B(y[65]), .Z(n4781) );
  NANDN U11844 ( .A(x[64]), .B(y[64]), .Z(n4780) );
  AND U11845 ( .A(n4781), .B(n4780), .Z(n24663) );
  NANDN U11846 ( .A(y[63]), .B(x[63]), .Z(n4783) );
  NANDN U11847 ( .A(y[64]), .B(x[64]), .Z(n4782) );
  NAND U11848 ( .A(n4783), .B(n4782), .Z(n24661) );
  NANDN U11849 ( .A(x[63]), .B(y[63]), .Z(n4785) );
  NANDN U11850 ( .A(x[62]), .B(y[62]), .Z(n4784) );
  AND U11851 ( .A(n4785), .B(n4784), .Z(n24659) );
  NANDN U11852 ( .A(y[61]), .B(x[61]), .Z(n4787) );
  NANDN U11853 ( .A(y[62]), .B(x[62]), .Z(n4786) );
  NAND U11854 ( .A(n4787), .B(n4786), .Z(n24657) );
  NANDN U11855 ( .A(x[61]), .B(y[61]), .Z(n15376) );
  NANDN U11856 ( .A(y[60]), .B(x[60]), .Z(n15378) );
  XNOR U11857 ( .A(x[60]), .B(y[60]), .Z(n4914) );
  NANDN U11858 ( .A(x[59]), .B(y[59]), .Z(n15379) );
  ANDN U11859 ( .B(x[58]), .A(y[58]), .Z(n15381) );
  NANDN U11860 ( .A(x[58]), .B(y[58]), .Z(n15380) );
  ANDN U11861 ( .B(x[56]), .A(y[56]), .Z(n15385) );
  NANDN U11862 ( .A(x[55]), .B(y[55]), .Z(n15387) );
  NANDN U11863 ( .A(x[54]), .B(y[54]), .Z(n15388) );
  NANDN U11864 ( .A(x[53]), .B(y[53]), .Z(n15392) );
  AND U11865 ( .A(n15388), .B(n15392), .Z(n4900) );
  NANDN U11866 ( .A(y[52]), .B(x[52]), .Z(n15394) );
  NANDN U11867 ( .A(x[52]), .B(y[52]), .Z(n15391) );
  ANDN U11868 ( .B(x[50]), .A(y[50]), .Z(n15397) );
  NANDN U11869 ( .A(x[49]), .B(y[49]), .Z(n15399) );
  NANDN U11870 ( .A(x[48]), .B(y[48]), .Z(n15400) );
  NANDN U11871 ( .A(x[47]), .B(y[47]), .Z(n15403) );
  AND U11872 ( .A(n15400), .B(n15403), .Z(n4888) );
  ANDN U11873 ( .B(x[46]), .A(y[46]), .Z(n15405) );
  NANDN U11874 ( .A(x[46]), .B(y[46]), .Z(n15404) );
  NANDN U11875 ( .A(y[44]), .B(x[44]), .Z(n15410) );
  NANDN U11876 ( .A(x[43]), .B(y[43]), .Z(n15412) );
  NANDN U11877 ( .A(x[42]), .B(y[42]), .Z(n15411) );
  NANDN U11878 ( .A(x[41]), .B(y[41]), .Z(n15416) );
  AND U11879 ( .A(n15411), .B(n15416), .Z(n4876) );
  NANDN U11880 ( .A(y[40]), .B(x[40]), .Z(n15418) );
  NANDN U11881 ( .A(x[40]), .B(y[40]), .Z(n15415) );
  ANDN U11882 ( .B(x[38]), .A(y[38]), .Z(n4870) );
  ANDN U11883 ( .B(x[37]), .A(y[37]), .Z(n15422) );
  NANDN U11884 ( .A(x[37]), .B(y[37]), .Z(n15423) );
  ANDN U11885 ( .B(x[36]), .A(y[36]), .Z(n4864) );
  NANDN U11886 ( .A(x[35]), .B(y[35]), .Z(n15428) );
  XNOR U11887 ( .A(x[36]), .B(y[36]), .Z(n15426) );
  AND U11888 ( .A(n15428), .B(n15426), .Z(n4862) );
  NANDN U11889 ( .A(y[34]), .B(x[34]), .Z(n15430) );
  NANDN U11890 ( .A(x[34]), .B(y[34]), .Z(n15427) );
  ANDN U11891 ( .B(x[32]), .A(y[32]), .Z(n4856) );
  NANDN U11892 ( .A(x[31]), .B(y[31]), .Z(n15435) );
  NANDN U11893 ( .A(x[29]), .B(y[29]), .Z(n15439) );
  XNOR U11894 ( .A(x[30]), .B(y[30]), .Z(n15438) );
  AND U11895 ( .A(n15439), .B(n15438), .Z(n4848) );
  NANDN U11896 ( .A(y[28]), .B(x[28]), .Z(n15442) );
  NANDN U11897 ( .A(x[28]), .B(y[28]), .Z(n15440) );
  ANDN U11898 ( .B(x[26]), .A(y[26]), .Z(n4842) );
  NANDN U11899 ( .A(x[25]), .B(y[25]), .Z(n15448) );
  NANDN U11900 ( .A(x[24]), .B(y[24]), .Z(n15447) );
  NANDN U11901 ( .A(x[23]), .B(y[23]), .Z(n15452) );
  AND U11902 ( .A(n15447), .B(n15452), .Z(n4835) );
  ANDN U11903 ( .B(x[22]), .A(y[22]), .Z(n15453) );
  NANDN U11904 ( .A(x[22]), .B(y[22]), .Z(n15451) );
  NANDN U11905 ( .A(y[20]), .B(x[20]), .Z(n15458) );
  NANDN U11906 ( .A(x[19]), .B(y[19]), .Z(n15460) );
  NANDN U11907 ( .A(x[18]), .B(y[18]), .Z(n15459) );
  NANDN U11908 ( .A(x[17]), .B(y[17]), .Z(n15464) );
  AND U11909 ( .A(n15459), .B(n15464), .Z(n4823) );
  ANDN U11910 ( .B(x[16]), .A(y[16]), .Z(n15465) );
  NANDN U11911 ( .A(x[16]), .B(y[16]), .Z(n15463) );
  ANDN U11912 ( .B(x[14]), .A(y[14]), .Z(n15469) );
  NANDN U11913 ( .A(x[13]), .B(y[13]), .Z(n15472) );
  NANDN U11914 ( .A(x[12]), .B(y[12]), .Z(n15471) );
  NANDN U11915 ( .A(x[11]), .B(y[11]), .Z(n15476) );
  AND U11916 ( .A(n15471), .B(n15476), .Z(n4811) );
  NANDN U11917 ( .A(y[10]), .B(x[10]), .Z(n15478) );
  NANDN U11918 ( .A(x[10]), .B(y[10]), .Z(n15475) );
  NANDN U11919 ( .A(y[8]), .B(x[8]), .Z(n15481) );
  NANDN U11920 ( .A(x[7]), .B(y[7]), .Z(n15483) );
  NANDN U11921 ( .A(x[6]), .B(y[6]), .Z(n15484) );
  NANDN U11922 ( .A(x[5]), .B(y[5]), .Z(n15488) );
  AND U11923 ( .A(n15484), .B(n15488), .Z(n4799) );
  NANDN U11924 ( .A(y[4]), .B(x[4]), .Z(n15490) );
  NANDN U11925 ( .A(x[4]), .B(y[4]), .Z(n15487) );
  NANDN U11926 ( .A(x[3]), .B(y[3]), .Z(n4789) );
  NANDN U11927 ( .A(x[2]), .B(y[2]), .Z(n4788) );
  AND U11928 ( .A(n4789), .B(n4788), .Z(n15496) );
  NANDN U11929 ( .A(y[1]), .B(x[1]), .Z(n4791) );
  NANDN U11930 ( .A(y[2]), .B(x[2]), .Z(n4790) );
  NAND U11931 ( .A(n4791), .B(n4790), .Z(n15494) );
  NANDN U11932 ( .A(x[1]), .B(y[1]), .Z(n15492) );
  ANDN U11933 ( .B(n15492), .A(y[0]), .Z(n4792) );
  NAND U11934 ( .A(x[0]), .B(n4792), .Z(n4793) );
  NANDN U11935 ( .A(n15494), .B(n4793), .Z(n4794) );
  AND U11936 ( .A(n15496), .B(n4794), .Z(n24540) );
  ANDN U11937 ( .B(x[3]), .A(y[3]), .Z(n15489) );
  OR U11938 ( .A(n24540), .B(n15489), .Z(n4795) );
  NAND U11939 ( .A(n15487), .B(n4795), .Z(n4796) );
  NAND U11940 ( .A(n15490), .B(n4796), .Z(n4797) );
  NANDN U11941 ( .A(y[5]), .B(x[5]), .Z(n15486) );
  NANDN U11942 ( .A(n4797), .B(n15486), .Z(n4798) );
  AND U11943 ( .A(n4799), .B(n4798), .Z(n4801) );
  NANDN U11944 ( .A(y[7]), .B(x[7]), .Z(n15482) );
  ANDN U11945 ( .B(x[6]), .A(y[6]), .Z(n15485) );
  ANDN U11946 ( .B(n15482), .A(n15485), .Z(n4800) );
  NANDN U11947 ( .A(n4801), .B(n4800), .Z(n4802) );
  AND U11948 ( .A(n15483), .B(n4802), .Z(n4803) );
  NANDN U11949 ( .A(x[8]), .B(y[8]), .Z(n15480) );
  NAND U11950 ( .A(n4803), .B(n15480), .Z(n4804) );
  ANDN U11951 ( .B(x[9]), .A(y[9]), .Z(n15477) );
  ANDN U11952 ( .B(n4804), .A(n15477), .Z(n4805) );
  NAND U11953 ( .A(n15481), .B(n4805), .Z(n4806) );
  NANDN U11954 ( .A(x[9]), .B(y[9]), .Z(n15479) );
  AND U11955 ( .A(n4806), .B(n15479), .Z(n4807) );
  NAND U11956 ( .A(n15475), .B(n4807), .Z(n4808) );
  NAND U11957 ( .A(n15478), .B(n4808), .Z(n4809) );
  ANDN U11958 ( .B(x[11]), .A(y[11]), .Z(n15473) );
  OR U11959 ( .A(n4809), .B(n15473), .Z(n4810) );
  AND U11960 ( .A(n4811), .B(n4810), .Z(n4813) );
  NANDN U11961 ( .A(y[13]), .B(x[13]), .Z(n15470) );
  NANDN U11962 ( .A(y[12]), .B(x[12]), .Z(n15474) );
  AND U11963 ( .A(n15470), .B(n15474), .Z(n4812) );
  NANDN U11964 ( .A(n4813), .B(n4812), .Z(n4814) );
  AND U11965 ( .A(n15472), .B(n4814), .Z(n4815) );
  NANDN U11966 ( .A(x[14]), .B(y[14]), .Z(n15467) );
  NAND U11967 ( .A(n4815), .B(n15467), .Z(n4816) );
  NANDN U11968 ( .A(y[15]), .B(x[15]), .Z(n15466) );
  AND U11969 ( .A(n4816), .B(n15466), .Z(n4817) );
  NANDN U11970 ( .A(n15469), .B(n4817), .Z(n4818) );
  NANDN U11971 ( .A(x[15]), .B(y[15]), .Z(n15468) );
  AND U11972 ( .A(n4818), .B(n15468), .Z(n4819) );
  NAND U11973 ( .A(n15463), .B(n4819), .Z(n4820) );
  NANDN U11974 ( .A(n15465), .B(n4820), .Z(n4821) );
  ANDN U11975 ( .B(x[17]), .A(y[17]), .Z(n15461) );
  OR U11976 ( .A(n4821), .B(n15461), .Z(n4822) );
  AND U11977 ( .A(n4823), .B(n4822), .Z(n4825) );
  NANDN U11978 ( .A(y[18]), .B(x[18]), .Z(n15462) );
  ANDN U11979 ( .B(x[19]), .A(y[19]), .Z(n15457) );
  ANDN U11980 ( .B(n15462), .A(n15457), .Z(n4824) );
  NANDN U11981 ( .A(n4825), .B(n4824), .Z(n4826) );
  AND U11982 ( .A(n15460), .B(n4826), .Z(n4827) );
  NANDN U11983 ( .A(x[20]), .B(y[20]), .Z(n15456) );
  NAND U11984 ( .A(n4827), .B(n15456), .Z(n4828) );
  NANDN U11985 ( .A(y[21]), .B(x[21]), .Z(n15454) );
  AND U11986 ( .A(n4828), .B(n15454), .Z(n4829) );
  NAND U11987 ( .A(n15458), .B(n4829), .Z(n4830) );
  NANDN U11988 ( .A(x[21]), .B(y[21]), .Z(n15455) );
  AND U11989 ( .A(n4830), .B(n15455), .Z(n4831) );
  NAND U11990 ( .A(n15451), .B(n4831), .Z(n4832) );
  NANDN U11991 ( .A(n15453), .B(n4832), .Z(n4833) );
  ANDN U11992 ( .B(x[23]), .A(y[23]), .Z(n15449) );
  OR U11993 ( .A(n4833), .B(n15449), .Z(n4834) );
  AND U11994 ( .A(n4835), .B(n4834), .Z(n4837) );
  NANDN U11995 ( .A(y[24]), .B(x[24]), .Z(n15450) );
  ANDN U11996 ( .B(x[25]), .A(y[25]), .Z(n15446) );
  ANDN U11997 ( .B(n15450), .A(n15446), .Z(n4836) );
  NANDN U11998 ( .A(n4837), .B(n4836), .Z(n4838) );
  AND U11999 ( .A(n15448), .B(n4838), .Z(n4839) );
  NANDN U12000 ( .A(x[26]), .B(y[26]), .Z(n15444) );
  NAND U12001 ( .A(n4839), .B(n15444), .Z(n4840) );
  ANDN U12002 ( .B(x[27]), .A(y[27]), .Z(n15441) );
  ANDN U12003 ( .B(n4840), .A(n15441), .Z(n4841) );
  NANDN U12004 ( .A(n4842), .B(n4841), .Z(n4843) );
  NANDN U12005 ( .A(x[27]), .B(y[27]), .Z(n15443) );
  AND U12006 ( .A(n4843), .B(n15443), .Z(n4844) );
  NAND U12007 ( .A(n15440), .B(n4844), .Z(n4845) );
  NAND U12008 ( .A(n15442), .B(n4845), .Z(n4846) );
  ANDN U12009 ( .B(x[29]), .A(y[29]), .Z(n15437) );
  OR U12010 ( .A(n4846), .B(n15437), .Z(n4847) );
  AND U12011 ( .A(n4848), .B(n4847), .Z(n4851) );
  ANDN U12012 ( .B(x[31]), .A(y[31]), .Z(n15434) );
  ANDN U12013 ( .B(x[30]), .A(y[30]), .Z(n4849) );
  NOR U12014 ( .A(n15434), .B(n4849), .Z(n4850) );
  NANDN U12015 ( .A(n4851), .B(n4850), .Z(n4852) );
  AND U12016 ( .A(n15435), .B(n4852), .Z(n4853) );
  NANDN U12017 ( .A(x[32]), .B(y[32]), .Z(n15432) );
  NAND U12018 ( .A(n4853), .B(n15432), .Z(n4854) );
  ANDN U12019 ( .B(x[33]), .A(y[33]), .Z(n15429) );
  ANDN U12020 ( .B(n4854), .A(n15429), .Z(n4855) );
  NANDN U12021 ( .A(n4856), .B(n4855), .Z(n4857) );
  NANDN U12022 ( .A(x[33]), .B(y[33]), .Z(n15431) );
  AND U12023 ( .A(n4857), .B(n15431), .Z(n4858) );
  NAND U12024 ( .A(n15427), .B(n4858), .Z(n4859) );
  NAND U12025 ( .A(n15430), .B(n4859), .Z(n4860) );
  ANDN U12026 ( .B(x[35]), .A(y[35]), .Z(n15425) );
  OR U12027 ( .A(n4860), .B(n15425), .Z(n4861) );
  AND U12028 ( .A(n4862), .B(n4861), .Z(n4863) );
  OR U12029 ( .A(n4864), .B(n4863), .Z(n4865) );
  NAND U12030 ( .A(n15423), .B(n4865), .Z(n4866) );
  NANDN U12031 ( .A(n15422), .B(n4866), .Z(n4867) );
  NANDN U12032 ( .A(x[38]), .B(y[38]), .Z(n15420) );
  NAND U12033 ( .A(n4867), .B(n15420), .Z(n4868) );
  ANDN U12034 ( .B(x[39]), .A(y[39]), .Z(n15417) );
  ANDN U12035 ( .B(n4868), .A(n15417), .Z(n4869) );
  NANDN U12036 ( .A(n4870), .B(n4869), .Z(n4871) );
  NANDN U12037 ( .A(x[39]), .B(y[39]), .Z(n15419) );
  AND U12038 ( .A(n4871), .B(n15419), .Z(n4872) );
  NAND U12039 ( .A(n15415), .B(n4872), .Z(n4873) );
  NAND U12040 ( .A(n15418), .B(n4873), .Z(n4874) );
  ANDN U12041 ( .B(x[41]), .A(y[41]), .Z(n15413) );
  OR U12042 ( .A(n4874), .B(n15413), .Z(n4875) );
  AND U12043 ( .A(n4876), .B(n4875), .Z(n4878) );
  NANDN U12044 ( .A(y[42]), .B(x[42]), .Z(n15414) );
  ANDN U12045 ( .B(x[43]), .A(y[43]), .Z(n15409) );
  ANDN U12046 ( .B(n15414), .A(n15409), .Z(n4877) );
  NANDN U12047 ( .A(n4878), .B(n4877), .Z(n4879) );
  AND U12048 ( .A(n15412), .B(n4879), .Z(n4880) );
  NANDN U12049 ( .A(x[44]), .B(y[44]), .Z(n15408) );
  NAND U12050 ( .A(n4880), .B(n15408), .Z(n4881) );
  NANDN U12051 ( .A(y[45]), .B(x[45]), .Z(n15406) );
  AND U12052 ( .A(n4881), .B(n15406), .Z(n4882) );
  NAND U12053 ( .A(n15410), .B(n4882), .Z(n4883) );
  NANDN U12054 ( .A(x[45]), .B(y[45]), .Z(n15407) );
  AND U12055 ( .A(n4883), .B(n15407), .Z(n4884) );
  NAND U12056 ( .A(n15404), .B(n4884), .Z(n4885) );
  NANDN U12057 ( .A(n15405), .B(n4885), .Z(n4886) );
  NANDN U12058 ( .A(y[47]), .B(x[47]), .Z(n15402) );
  NANDN U12059 ( .A(n4886), .B(n15402), .Z(n4887) );
  AND U12060 ( .A(n4888), .B(n4887), .Z(n4890) );
  NANDN U12061 ( .A(y[49]), .B(x[49]), .Z(n15398) );
  ANDN U12062 ( .B(x[48]), .A(y[48]), .Z(n15401) );
  ANDN U12063 ( .B(n15398), .A(n15401), .Z(n4889) );
  NANDN U12064 ( .A(n4890), .B(n4889), .Z(n4891) );
  AND U12065 ( .A(n15399), .B(n4891), .Z(n4892) );
  NANDN U12066 ( .A(x[50]), .B(y[50]), .Z(n15396) );
  NAND U12067 ( .A(n4892), .B(n15396), .Z(n4893) );
  ANDN U12068 ( .B(x[51]), .A(y[51]), .Z(n15393) );
  ANDN U12069 ( .B(n4893), .A(n15393), .Z(n4894) );
  NANDN U12070 ( .A(n15397), .B(n4894), .Z(n4895) );
  NANDN U12071 ( .A(x[51]), .B(y[51]), .Z(n15395) );
  AND U12072 ( .A(n4895), .B(n15395), .Z(n4896) );
  NAND U12073 ( .A(n15391), .B(n4896), .Z(n4897) );
  NAND U12074 ( .A(n15394), .B(n4897), .Z(n4898) );
  ANDN U12075 ( .B(x[53]), .A(y[53]), .Z(n15390) );
  OR U12076 ( .A(n4898), .B(n15390), .Z(n4899) );
  AND U12077 ( .A(n4900), .B(n4899), .Z(n4903) );
  NANDN U12078 ( .A(y[55]), .B(x[55]), .Z(n15386) );
  ANDN U12079 ( .B(x[54]), .A(y[54]), .Z(n4901) );
  ANDN U12080 ( .B(n15386), .A(n4901), .Z(n4902) );
  NANDN U12081 ( .A(n4903), .B(n4902), .Z(n4904) );
  AND U12082 ( .A(n15387), .B(n4904), .Z(n4905) );
  NANDN U12083 ( .A(x[56]), .B(y[56]), .Z(n15384) );
  NAND U12084 ( .A(n4905), .B(n15384), .Z(n4906) );
  NANDN U12085 ( .A(y[57]), .B(x[57]), .Z(n15382) );
  AND U12086 ( .A(n4906), .B(n15382), .Z(n4907) );
  NANDN U12087 ( .A(n15385), .B(n4907), .Z(n4908) );
  NANDN U12088 ( .A(x[57]), .B(y[57]), .Z(n15383) );
  AND U12089 ( .A(n4908), .B(n15383), .Z(n4909) );
  NAND U12090 ( .A(n15380), .B(n4909), .Z(n4910) );
  NANDN U12091 ( .A(n15381), .B(n4910), .Z(n4911) );
  ANDN U12092 ( .B(x[59]), .A(y[59]), .Z(n15377) );
  OR U12093 ( .A(n4911), .B(n15377), .Z(n4912) );
  AND U12094 ( .A(n15379), .B(n4912), .Z(n4913) );
  NAND U12095 ( .A(n4914), .B(n4913), .Z(n4915) );
  NAND U12096 ( .A(n15378), .B(n4915), .Z(n4916) );
  AND U12097 ( .A(n15376), .B(n4916), .Z(n4917) );
  OR U12098 ( .A(n24657), .B(n4917), .Z(n4918) );
  AND U12099 ( .A(n24659), .B(n4918), .Z(n4919) );
  OR U12100 ( .A(n24661), .B(n4919), .Z(n4920) );
  NAND U12101 ( .A(n24663), .B(n4920), .Z(n4921) );
  NANDN U12102 ( .A(n15373), .B(n4921), .Z(n4922) );
  NANDN U12103 ( .A(x[66]), .B(y[66]), .Z(n15371) );
  NAND U12104 ( .A(n4922), .B(n15371), .Z(n4923) );
  ANDN U12105 ( .B(x[67]), .A(y[67]), .Z(n15369) );
  ANDN U12106 ( .B(n4923), .A(n15369), .Z(n4924) );
  NAND U12107 ( .A(n15374), .B(n4924), .Z(n4925) );
  NANDN U12108 ( .A(x[67]), .B(y[67]), .Z(n15372) );
  AND U12109 ( .A(n4925), .B(n15372), .Z(n4926) );
  NAND U12110 ( .A(n15367), .B(n4926), .Z(n4927) );
  NAND U12111 ( .A(n15370), .B(n4927), .Z(n4929) );
  NANDN U12112 ( .A(y[69]), .B(n4929), .Z(n4928) );
  ANDN U12113 ( .B(x[70]), .A(y[70]), .Z(n15366) );
  ANDN U12114 ( .B(n4928), .A(n15366), .Z(n4932) );
  XNOR U12115 ( .A(n4929), .B(y[69]), .Z(n4930) );
  NAND U12116 ( .A(n4930), .B(x[69]), .Z(n4931) );
  NAND U12117 ( .A(n4932), .B(n4931), .Z(n4933) );
  NAND U12118 ( .A(n24675), .B(n4933), .Z(n4934) );
  NANDN U12119 ( .A(n24677), .B(n4934), .Z(n4935) );
  AND U12120 ( .A(n15365), .B(n4935), .Z(n4936) );
  ANDN U12121 ( .B(x[73]), .A(y[73]), .Z(n15362) );
  OR U12122 ( .A(n4936), .B(n15362), .Z(n4937) );
  AND U12123 ( .A(n4938), .B(n4937), .Z(n4940) );
  NANDN U12124 ( .A(y[74]), .B(x[74]), .Z(n15363) );
  ANDN U12125 ( .B(x[75]), .A(y[75]), .Z(n15358) );
  ANDN U12126 ( .B(n15363), .A(n15358), .Z(n4939) );
  NANDN U12127 ( .A(n4940), .B(n4939), .Z(n4941) );
  AND U12128 ( .A(n15360), .B(n4941), .Z(n4942) );
  NAND U12129 ( .A(n4943), .B(n4942), .Z(n4944) );
  NAND U12130 ( .A(n15359), .B(n4944), .Z(n4945) );
  AND U12131 ( .A(n15357), .B(n4945), .Z(n4948) );
  NANDN U12132 ( .A(y[77]), .B(x[77]), .Z(n4947) );
  NANDN U12133 ( .A(y[78]), .B(x[78]), .Z(n4946) );
  NAND U12134 ( .A(n4947), .B(n4946), .Z(n24689) );
  OR U12135 ( .A(n4948), .B(n24689), .Z(n4949) );
  NAND U12136 ( .A(n24691), .B(n4949), .Z(n4950) );
  NANDN U12137 ( .A(n15355), .B(n4950), .Z(n4951) );
  NANDN U12138 ( .A(x[80]), .B(y[80]), .Z(n15353) );
  NAND U12139 ( .A(n4951), .B(n15353), .Z(n4952) );
  ANDN U12140 ( .B(x[81]), .A(y[81]), .Z(n15350) );
  ANDN U12141 ( .B(n4952), .A(n15350), .Z(n4953) );
  NANDN U12142 ( .A(n4954), .B(n4953), .Z(n4955) );
  NANDN U12143 ( .A(x[81]), .B(y[81]), .Z(n15352) );
  AND U12144 ( .A(n4955), .B(n15352), .Z(n4956) );
  NAND U12145 ( .A(n15349), .B(n4956), .Z(n4957) );
  NAND U12146 ( .A(n15351), .B(n4957), .Z(n4958) );
  ANDN U12147 ( .B(x[83]), .A(y[83]), .Z(n15347) );
  OR U12148 ( .A(n4958), .B(n15347), .Z(n4959) );
  AND U12149 ( .A(n4960), .B(n4959), .Z(n4963) );
  ANDN U12150 ( .B(x[85]), .A(y[85]), .Z(n15342) );
  ANDN U12151 ( .B(x[84]), .A(y[84]), .Z(n4961) );
  NOR U12152 ( .A(n15342), .B(n4961), .Z(n4962) );
  NANDN U12153 ( .A(n4963), .B(n4962), .Z(n4964) );
  AND U12154 ( .A(n15344), .B(n4964), .Z(n4965) );
  NANDN U12155 ( .A(x[86]), .B(y[86]), .Z(n15340) );
  NAND U12156 ( .A(n4965), .B(n15340), .Z(n4966) );
  ANDN U12157 ( .B(x[87]), .A(y[87]), .Z(n15338) );
  ANDN U12158 ( .B(n4966), .A(n15338), .Z(n4967) );
  NAND U12159 ( .A(n15343), .B(n4967), .Z(n4968) );
  NANDN U12160 ( .A(x[87]), .B(y[87]), .Z(n15341) );
  AND U12161 ( .A(n4968), .B(n15341), .Z(n4969) );
  NAND U12162 ( .A(n15336), .B(n4969), .Z(n4970) );
  NAND U12163 ( .A(n15339), .B(n4970), .Z(n4971) );
  NANDN U12164 ( .A(y[89]), .B(x[89]), .Z(n15335) );
  NANDN U12165 ( .A(n4971), .B(n15335), .Z(n4972) );
  AND U12166 ( .A(n4973), .B(n4972), .Z(n4975) );
  NANDN U12167 ( .A(y[91]), .B(x[91]), .Z(n15331) );
  ANDN U12168 ( .B(x[90]), .A(y[90]), .Z(n15334) );
  ANDN U12169 ( .B(n15331), .A(n15334), .Z(n4974) );
  NANDN U12170 ( .A(n4975), .B(n4974), .Z(n4976) );
  AND U12171 ( .A(n15332), .B(n4976), .Z(n4977) );
  NANDN U12172 ( .A(x[92]), .B(y[92]), .Z(n15329) );
  NAND U12173 ( .A(n4977), .B(n15329), .Z(n4978) );
  NANDN U12174 ( .A(y[93]), .B(x[93]), .Z(n15327) );
  AND U12175 ( .A(n4978), .B(n15327), .Z(n4979) );
  NAND U12176 ( .A(n15330), .B(n4979), .Z(n4980) );
  NANDN U12177 ( .A(x[93]), .B(y[93]), .Z(n15328) );
  AND U12178 ( .A(n4980), .B(n15328), .Z(n4981) );
  NAND U12179 ( .A(n15324), .B(n4981), .Z(n4982) );
  NANDN U12180 ( .A(n15326), .B(n4982), .Z(n4983) );
  ANDN U12181 ( .B(x[95]), .A(y[95]), .Z(n15322) );
  OR U12182 ( .A(n4983), .B(n15322), .Z(n4984) );
  AND U12183 ( .A(n4985), .B(n4984), .Z(n4988) );
  ANDN U12184 ( .B(x[97]), .A(y[97]), .Z(n15318) );
  ANDN U12185 ( .B(x[96]), .A(y[96]), .Z(n4986) );
  NOR U12186 ( .A(n15318), .B(n4986), .Z(n4987) );
  NANDN U12187 ( .A(n4988), .B(n4987), .Z(n4989) );
  AND U12188 ( .A(n15320), .B(n4989), .Z(n4990) );
  NANDN U12189 ( .A(x[98]), .B(y[98]), .Z(n15316) );
  NAND U12190 ( .A(n4990), .B(n15316), .Z(n4991) );
  ANDN U12191 ( .B(x[99]), .A(y[99]), .Z(n15315) );
  ANDN U12192 ( .B(n4991), .A(n15315), .Z(n4992) );
  NAND U12193 ( .A(n15319), .B(n4992), .Z(n4993) );
  NAND U12194 ( .A(n15317), .B(n4993), .Z(n4995) );
  NANDN U12195 ( .A(x[100]), .B(n4995), .Z(n4994) );
  ANDN U12196 ( .B(y[101]), .A(x[101]), .Z(n15314) );
  ANDN U12197 ( .B(n4994), .A(n15314), .Z(n4998) );
  XNOR U12198 ( .A(n4995), .B(x[100]), .Z(n4996) );
  NAND U12199 ( .A(n4996), .B(y[100]), .Z(n4997) );
  NAND U12200 ( .A(n4998), .B(n4997), .Z(n4999) );
  NAND U12201 ( .A(n15595), .B(n4999), .Z(n5000) );
  NAND U12202 ( .A(n15313), .B(n5000), .Z(n5001) );
  AND U12203 ( .A(n15311), .B(n5001), .Z(n5003) );
  NANDN U12204 ( .A(x[104]), .B(y[104]), .Z(n15308) );
  ANDN U12205 ( .B(y[103]), .A(x[103]), .Z(n15312) );
  ANDN U12206 ( .B(n15308), .A(n15312), .Z(n5002) );
  NANDN U12207 ( .A(n5003), .B(n5002), .Z(n5004) );
  AND U12208 ( .A(n15310), .B(n5004), .Z(n5005) );
  NANDN U12209 ( .A(y[105]), .B(x[105]), .Z(n15307) );
  NAND U12210 ( .A(n5005), .B(n15307), .Z(n5006) );
  ANDN U12211 ( .B(y[106]), .A(x[106]), .Z(n15304) );
  ANDN U12212 ( .B(n5006), .A(n15304), .Z(n5007) );
  NAND U12213 ( .A(n15309), .B(n5007), .Z(n5008) );
  NANDN U12214 ( .A(y[106]), .B(x[106]), .Z(n15306) );
  AND U12215 ( .A(n5008), .B(n15306), .Z(n5009) );
  NAND U12216 ( .A(n15303), .B(n5009), .Z(n5010) );
  NAND U12217 ( .A(n15305), .B(n5010), .Z(n5011) );
  ANDN U12218 ( .B(y[108]), .A(x[108]), .Z(n15300) );
  OR U12219 ( .A(n5011), .B(n15300), .Z(n5012) );
  AND U12220 ( .A(n5013), .B(n5012), .Z(n5015) );
  NANDN U12221 ( .A(x[109]), .B(y[109]), .Z(n15301) );
  ANDN U12222 ( .B(y[110]), .A(x[110]), .Z(n15296) );
  ANDN U12223 ( .B(n15301), .A(n15296), .Z(n5014) );
  NANDN U12224 ( .A(n5015), .B(n5014), .Z(n5016) );
  AND U12225 ( .A(n15299), .B(n5016), .Z(n5017) );
  NANDN U12226 ( .A(y[111]), .B(x[111]), .Z(n15295) );
  NAND U12227 ( .A(n5017), .B(n15295), .Z(n5018) );
  NANDN U12228 ( .A(x[112]), .B(y[112]), .Z(n15293) );
  AND U12229 ( .A(n5018), .B(n15293), .Z(n5019) );
  NAND U12230 ( .A(n15297), .B(n5019), .Z(n5020) );
  NANDN U12231 ( .A(y[112]), .B(x[112]), .Z(n15294) );
  AND U12232 ( .A(n5020), .B(n15294), .Z(n5021) );
  NAND U12233 ( .A(n15288), .B(n5021), .Z(n5022) );
  NANDN U12234 ( .A(n15291), .B(n5022), .Z(n5023) );
  NANDN U12235 ( .A(x[114]), .B(y[114]), .Z(n15287) );
  NANDN U12236 ( .A(n5023), .B(n15287), .Z(n5024) );
  AND U12237 ( .A(n5025), .B(n5024), .Z(n5027) );
  NANDN U12238 ( .A(x[116]), .B(y[116]), .Z(n15283) );
  ANDN U12239 ( .B(y[115]), .A(x[115]), .Z(n15286) );
  ANDN U12240 ( .B(n15283), .A(n15286), .Z(n5026) );
  NANDN U12241 ( .A(n5027), .B(n5026), .Z(n5028) );
  AND U12242 ( .A(n15284), .B(n5028), .Z(n5029) );
  NANDN U12243 ( .A(y[117]), .B(x[117]), .Z(n15280) );
  NAND U12244 ( .A(n5029), .B(n15280), .Z(n5030) );
  ANDN U12245 ( .B(y[118]), .A(x[118]), .Z(n15278) );
  ANDN U12246 ( .B(n5030), .A(n15278), .Z(n5031) );
  NANDN U12247 ( .A(n15282), .B(n5031), .Z(n5032) );
  NANDN U12248 ( .A(y[118]), .B(x[118]), .Z(n15281) );
  AND U12249 ( .A(n5032), .B(n15281), .Z(n5033) );
  NAND U12250 ( .A(n15277), .B(n5033), .Z(n5034) );
  NAND U12251 ( .A(n15279), .B(n5034), .Z(n5035) );
  ANDN U12252 ( .B(y[120]), .A(x[120]), .Z(n15274) );
  OR U12253 ( .A(n5035), .B(n15274), .Z(n5036) );
  AND U12254 ( .A(n5037), .B(n5036), .Z(n5039) );
  NANDN U12255 ( .A(x[121]), .B(y[121]), .Z(n15275) );
  ANDN U12256 ( .B(y[122]), .A(x[122]), .Z(n15270) );
  ANDN U12257 ( .B(n15275), .A(n15270), .Z(n5038) );
  NANDN U12258 ( .A(n5039), .B(n5038), .Z(n5040) );
  AND U12259 ( .A(n15272), .B(n5040), .Z(n5041) );
  NANDN U12260 ( .A(y[123]), .B(x[123]), .Z(n15269) );
  NAND U12261 ( .A(n5041), .B(n15269), .Z(n5042) );
  NANDN U12262 ( .A(x[124]), .B(y[124]), .Z(n15267) );
  AND U12263 ( .A(n5042), .B(n15267), .Z(n5043) );
  NAND U12264 ( .A(n15271), .B(n5043), .Z(n5044) );
  NANDN U12265 ( .A(y[124]), .B(x[124]), .Z(n15268) );
  AND U12266 ( .A(n5044), .B(n15268), .Z(n5045) );
  NAND U12267 ( .A(n15265), .B(n5045), .Z(n5046) );
  NANDN U12268 ( .A(n15266), .B(n5046), .Z(n5047) );
  ANDN U12269 ( .B(y[126]), .A(x[126]), .Z(n15262) );
  OR U12270 ( .A(n5047), .B(n15262), .Z(n5048) );
  AND U12271 ( .A(n5049), .B(n5048), .Z(n5051) );
  NANDN U12272 ( .A(x[128]), .B(y[128]), .Z(n15260) );
  NANDN U12273 ( .A(x[127]), .B(y[127]), .Z(n15263) );
  AND U12274 ( .A(n15260), .B(n15263), .Z(n5050) );
  NANDN U12275 ( .A(n5051), .B(n5050), .Z(n5052) );
  AND U12276 ( .A(n5053), .B(n5052), .Z(n5054) );
  NANDN U12277 ( .A(y[129]), .B(x[129]), .Z(n15258) );
  NAND U12278 ( .A(n5054), .B(n15258), .Z(n5055) );
  NANDN U12279 ( .A(x[130]), .B(y[130]), .Z(n15256) );
  AND U12280 ( .A(n5055), .B(n15256), .Z(n5056) );
  NANDN U12281 ( .A(n15259), .B(n5056), .Z(n5057) );
  NANDN U12282 ( .A(y[130]), .B(x[130]), .Z(n15257) );
  AND U12283 ( .A(n5057), .B(n15257), .Z(n5058) );
  NAND U12284 ( .A(n15253), .B(n5058), .Z(n5059) );
  NANDN U12285 ( .A(n15255), .B(n5059), .Z(n5060) );
  NANDN U12286 ( .A(x[132]), .B(y[132]), .Z(n15252) );
  NANDN U12287 ( .A(n5060), .B(n15252), .Z(n5061) );
  AND U12288 ( .A(n5062), .B(n5061), .Z(n5064) );
  NANDN U12289 ( .A(x[134]), .B(y[134]), .Z(n15247) );
  ANDN U12290 ( .B(y[133]), .A(x[133]), .Z(n15251) );
  ANDN U12291 ( .B(n15247), .A(n15251), .Z(n5063) );
  NANDN U12292 ( .A(n5064), .B(n5063), .Z(n5065) );
  AND U12293 ( .A(n15249), .B(n5065), .Z(n5066) );
  NANDN U12294 ( .A(y[135]), .B(x[135]), .Z(n15246) );
  NAND U12295 ( .A(n5066), .B(n15246), .Z(n5067) );
  NANDN U12296 ( .A(x[136]), .B(y[136]), .Z(n15244) );
  AND U12297 ( .A(n5067), .B(n15244), .Z(n5068) );
  NAND U12298 ( .A(n15248), .B(n5068), .Z(n5069) );
  NANDN U12299 ( .A(y[136]), .B(x[136]), .Z(n15245) );
  AND U12300 ( .A(n5069), .B(n15245), .Z(n5070) );
  NAND U12301 ( .A(n15241), .B(n5070), .Z(n5071) );
  NANDN U12302 ( .A(n15243), .B(n5071), .Z(n5072) );
  NANDN U12303 ( .A(x[138]), .B(y[138]), .Z(n15240) );
  NANDN U12304 ( .A(n5072), .B(n15240), .Z(n5073) );
  AND U12305 ( .A(n5074), .B(n5073), .Z(n5076) );
  NANDN U12306 ( .A(x[140]), .B(y[140]), .Z(n15235) );
  ANDN U12307 ( .B(y[139]), .A(x[139]), .Z(n15239) );
  ANDN U12308 ( .B(n15235), .A(n15239), .Z(n5075) );
  NANDN U12309 ( .A(n5076), .B(n5075), .Z(n5077) );
  AND U12310 ( .A(n15237), .B(n5077), .Z(n5078) );
  NAND U12311 ( .A(n5079), .B(n5078), .Z(n5080) );
  NAND U12312 ( .A(n15236), .B(n5080), .Z(n5081) );
  AND U12313 ( .A(n15234), .B(n5081), .Z(n5084) );
  NANDN U12314 ( .A(x[142]), .B(y[142]), .Z(n5083) );
  NANDN U12315 ( .A(x[143]), .B(y[143]), .Z(n5082) );
  NAND U12316 ( .A(n5083), .B(n5082), .Z(n15637) );
  OR U12317 ( .A(n5084), .B(n15637), .Z(n5085) );
  NAND U12318 ( .A(n15639), .B(n5085), .Z(n5086) );
  NAND U12319 ( .A(n15232), .B(n5086), .Z(n5087) );
  NAND U12320 ( .A(n15230), .B(n5087), .Z(n5088) );
  NANDN U12321 ( .A(x[146]), .B(y[146]), .Z(n15229) );
  AND U12322 ( .A(n5088), .B(n15229), .Z(n5089) );
  NANDN U12323 ( .A(n15231), .B(n5089), .Z(n5091) );
  NANDN U12324 ( .A(y[146]), .B(x[146]), .Z(n5090) );
  AND U12325 ( .A(n5091), .B(n5090), .Z(n5092) );
  NAND U12326 ( .A(n15226), .B(n5092), .Z(n5093) );
  NANDN U12327 ( .A(n15228), .B(n5093), .Z(n5094) );
  NANDN U12328 ( .A(x[148]), .B(y[148]), .Z(n15225) );
  NANDN U12329 ( .A(n5094), .B(n15225), .Z(n5095) );
  AND U12330 ( .A(n5096), .B(n5095), .Z(n5098) );
  NANDN U12331 ( .A(x[150]), .B(y[150]), .Z(n15222) );
  ANDN U12332 ( .B(y[149]), .A(x[149]), .Z(n15224) );
  ANDN U12333 ( .B(n15222), .A(n15224), .Z(n5097) );
  NANDN U12334 ( .A(n5098), .B(n5097), .Z(n5099) );
  AND U12335 ( .A(n5100), .B(n5099), .Z(n5101) );
  NANDN U12336 ( .A(y[151]), .B(x[151]), .Z(n15220) );
  NAND U12337 ( .A(n5101), .B(n15220), .Z(n5102) );
  NANDN U12338 ( .A(x[152]), .B(y[152]), .Z(n15218) );
  AND U12339 ( .A(n5102), .B(n15218), .Z(n5103) );
  NANDN U12340 ( .A(n15221), .B(n5103), .Z(n5104) );
  NANDN U12341 ( .A(y[152]), .B(x[152]), .Z(n15219) );
  AND U12342 ( .A(n5104), .B(n15219), .Z(n5105) );
  NAND U12343 ( .A(n15215), .B(n5105), .Z(n5106) );
  NANDN U12344 ( .A(n15217), .B(n5106), .Z(n5107) );
  NANDN U12345 ( .A(x[154]), .B(y[154]), .Z(n15214) );
  NANDN U12346 ( .A(n5107), .B(n15214), .Z(n5108) );
  AND U12347 ( .A(n5109), .B(n5108), .Z(n5111) );
  NANDN U12348 ( .A(x[156]), .B(y[156]), .Z(n15209) );
  ANDN U12349 ( .B(y[155]), .A(x[155]), .Z(n15213) );
  ANDN U12350 ( .B(n15209), .A(n15213), .Z(n5110) );
  NANDN U12351 ( .A(n5111), .B(n5110), .Z(n5112) );
  AND U12352 ( .A(n15211), .B(n5112), .Z(n5113) );
  NANDN U12353 ( .A(y[157]), .B(x[157]), .Z(n15208) );
  NAND U12354 ( .A(n5113), .B(n15208), .Z(n5114) );
  ANDN U12355 ( .B(y[158]), .A(x[158]), .Z(n15205) );
  ANDN U12356 ( .B(n5114), .A(n15205), .Z(n5115) );
  NAND U12357 ( .A(n15210), .B(n5115), .Z(n5116) );
  NANDN U12358 ( .A(y[158]), .B(x[158]), .Z(n15207) );
  AND U12359 ( .A(n5116), .B(n15207), .Z(n5117) );
  NAND U12360 ( .A(n15203), .B(n5117), .Z(n5118) );
  NAND U12361 ( .A(n15206), .B(n5118), .Z(n5119) );
  NANDN U12362 ( .A(x[160]), .B(y[160]), .Z(n15202) );
  NANDN U12363 ( .A(n5119), .B(n15202), .Z(n5120) );
  AND U12364 ( .A(n5121), .B(n5120), .Z(n5123) );
  NANDN U12365 ( .A(x[162]), .B(y[162]), .Z(n15198) );
  ANDN U12366 ( .B(y[161]), .A(x[161]), .Z(n15201) );
  ANDN U12367 ( .B(n15198), .A(n15201), .Z(n5122) );
  NANDN U12368 ( .A(n5123), .B(n5122), .Z(n5124) );
  AND U12369 ( .A(n15200), .B(n5124), .Z(n5125) );
  NANDN U12370 ( .A(y[163]), .B(x[163]), .Z(n15195) );
  NAND U12371 ( .A(n5125), .B(n15195), .Z(n5126) );
  NANDN U12372 ( .A(x[164]), .B(y[164]), .Z(n15194) );
  AND U12373 ( .A(n5126), .B(n15194), .Z(n5127) );
  NANDN U12374 ( .A(n15197), .B(n5127), .Z(n5128) );
  NANDN U12375 ( .A(y[164]), .B(x[164]), .Z(n15196) );
  AND U12376 ( .A(n5128), .B(n15196), .Z(n5129) );
  NAND U12377 ( .A(n15192), .B(n5129), .Z(n5130) );
  NANDN U12378 ( .A(n15193), .B(n5130), .Z(n5131) );
  NANDN U12379 ( .A(x[166]), .B(y[166]), .Z(n15190) );
  NANDN U12380 ( .A(n5131), .B(n15190), .Z(n5132) );
  AND U12381 ( .A(n5133), .B(n5132), .Z(n5135) );
  NANDN U12382 ( .A(x[168]), .B(y[168]), .Z(n15185) );
  ANDN U12383 ( .B(y[167]), .A(x[167]), .Z(n15188) );
  ANDN U12384 ( .B(n15185), .A(n15188), .Z(n5134) );
  NANDN U12385 ( .A(n5135), .B(n5134), .Z(n5136) );
  AND U12386 ( .A(n15186), .B(n5136), .Z(n5137) );
  NANDN U12387 ( .A(y[169]), .B(x[169]), .Z(n15183) );
  NAND U12388 ( .A(n5137), .B(n15183), .Z(n5138) );
  ANDN U12389 ( .B(y[169]), .A(x[169]), .Z(n15184) );
  ANDN U12390 ( .B(n5138), .A(n15184), .Z(n5139) );
  NANDN U12391 ( .A(n15182), .B(n5139), .Z(n5141) );
  NANDN U12392 ( .A(y[170]), .B(x[170]), .Z(n5140) );
  AND U12393 ( .A(n5141), .B(n5140), .Z(n5142) );
  NAND U12394 ( .A(n15180), .B(n5142), .Z(n5143) );
  NANDN U12395 ( .A(n15181), .B(n5143), .Z(n5144) );
  ANDN U12396 ( .B(y[172]), .A(x[172]), .Z(n15176) );
  OR U12397 ( .A(n5144), .B(n15176), .Z(n5145) );
  AND U12398 ( .A(n5146), .B(n5145), .Z(n5148) );
  NANDN U12399 ( .A(x[174]), .B(y[174]), .Z(n15172) );
  NANDN U12400 ( .A(x[173]), .B(y[173]), .Z(n15178) );
  AND U12401 ( .A(n15172), .B(n15178), .Z(n5147) );
  NANDN U12402 ( .A(n5148), .B(n5147), .Z(n5149) );
  AND U12403 ( .A(n5150), .B(n5149), .Z(n5151) );
  NAND U12404 ( .A(n15167), .B(n5151), .Z(n5152) );
  NANDN U12405 ( .A(x[176]), .B(y[176]), .Z(n15166) );
  AND U12406 ( .A(n5152), .B(n15166), .Z(n5153) );
  NANDN U12407 ( .A(n15170), .B(n5153), .Z(n5155) );
  NANDN U12408 ( .A(y[176]), .B(x[176]), .Z(n5154) );
  AND U12409 ( .A(n5155), .B(n5154), .Z(n5156) );
  NAND U12410 ( .A(n15163), .B(n5156), .Z(n5157) );
  NANDN U12411 ( .A(n15165), .B(n5157), .Z(n5158) );
  NANDN U12412 ( .A(x[178]), .B(y[178]), .Z(n15162) );
  NANDN U12413 ( .A(n5158), .B(n15162), .Z(n5159) );
  AND U12414 ( .A(n5160), .B(n5159), .Z(n5162) );
  NANDN U12415 ( .A(x[180]), .B(y[180]), .Z(n15159) );
  ANDN U12416 ( .B(y[179]), .A(x[179]), .Z(n15161) );
  ANDN U12417 ( .B(n15159), .A(n15161), .Z(n5161) );
  NANDN U12418 ( .A(n5162), .B(n5161), .Z(n5163) );
  AND U12419 ( .A(n5164), .B(n5163), .Z(n5165) );
  NAND U12420 ( .A(n15157), .B(n5165), .Z(n5166) );
  NANDN U12421 ( .A(x[182]), .B(y[182]), .Z(n15156) );
  AND U12422 ( .A(n5166), .B(n15156), .Z(n5167) );
  NANDN U12423 ( .A(n15158), .B(n5167), .Z(n5169) );
  NANDN U12424 ( .A(y[182]), .B(x[182]), .Z(n5168) );
  AND U12425 ( .A(n5169), .B(n5168), .Z(n5170) );
  NAND U12426 ( .A(n15154), .B(n5170), .Z(n5171) );
  NANDN U12427 ( .A(n15155), .B(n5171), .Z(n5172) );
  ANDN U12428 ( .B(y[184]), .A(x[184]), .Z(n15151) );
  OR U12429 ( .A(n5172), .B(n15151), .Z(n5173) );
  AND U12430 ( .A(n5174), .B(n5173), .Z(n5176) );
  NANDN U12431 ( .A(x[185]), .B(y[185]), .Z(n15152) );
  ANDN U12432 ( .B(y[186]), .A(x[186]), .Z(n15146) );
  ANDN U12433 ( .B(n15152), .A(n15146), .Z(n5175) );
  NANDN U12434 ( .A(n5176), .B(n5175), .Z(n5177) );
  AND U12435 ( .A(n15149), .B(n5177), .Z(n5178) );
  NANDN U12436 ( .A(y[187]), .B(x[187]), .Z(n15145) );
  NAND U12437 ( .A(n5178), .B(n15145), .Z(n5179) );
  ANDN U12438 ( .B(y[188]), .A(x[188]), .Z(n15142) );
  ANDN U12439 ( .B(n5179), .A(n15142), .Z(n5180) );
  NAND U12440 ( .A(n15148), .B(n5180), .Z(n5181) );
  NANDN U12441 ( .A(y[188]), .B(x[188]), .Z(n15144) );
  AND U12442 ( .A(n5181), .B(n15144), .Z(n5182) );
  NAND U12443 ( .A(n15140), .B(n5182), .Z(n5183) );
  NAND U12444 ( .A(n15143), .B(n5183), .Z(n5184) );
  ANDN U12445 ( .B(y[190]), .A(x[190]), .Z(n15138) );
  OR U12446 ( .A(n5184), .B(n15138), .Z(n5185) );
  AND U12447 ( .A(n5186), .B(n5185), .Z(n5188) );
  NANDN U12448 ( .A(x[192]), .B(y[192]), .Z(n15135) );
  NANDN U12449 ( .A(x[191]), .B(y[191]), .Z(n15139) );
  AND U12450 ( .A(n15135), .B(n15139), .Z(n5187) );
  NANDN U12451 ( .A(n5188), .B(n5187), .Z(n5189) );
  AND U12452 ( .A(n15136), .B(n5189), .Z(n5190) );
  NANDN U12453 ( .A(y[193]), .B(x[193]), .Z(n15132) );
  NAND U12454 ( .A(n5190), .B(n15132), .Z(n5191) );
  NANDN U12455 ( .A(x[194]), .B(y[194]), .Z(n15131) );
  AND U12456 ( .A(n5191), .B(n15131), .Z(n5192) );
  NANDN U12457 ( .A(n15134), .B(n5192), .Z(n5193) );
  NANDN U12458 ( .A(y[194]), .B(x[194]), .Z(n15133) );
  AND U12459 ( .A(n5193), .B(n15133), .Z(n5194) );
  NAND U12460 ( .A(n15128), .B(n5194), .Z(n5195) );
  NANDN U12461 ( .A(n15130), .B(n5195), .Z(n5196) );
  ANDN U12462 ( .B(y[196]), .A(x[196]), .Z(n15126) );
  OR U12463 ( .A(n5196), .B(n15126), .Z(n5197) );
  AND U12464 ( .A(n5198), .B(n5197), .Z(n5200) );
  NANDN U12465 ( .A(x[198]), .B(y[198]), .Z(n15124) );
  NANDN U12466 ( .A(x[197]), .B(y[197]), .Z(n15127) );
  AND U12467 ( .A(n15124), .B(n15127), .Z(n5199) );
  NANDN U12468 ( .A(n5200), .B(n5199), .Z(n5201) );
  AND U12469 ( .A(n5202), .B(n5201), .Z(n5203) );
  NANDN U12470 ( .A(y[199]), .B(x[199]), .Z(n15121) );
  NAND U12471 ( .A(n5203), .B(n15121), .Z(n5204) );
  NANDN U12472 ( .A(x[200]), .B(y[200]), .Z(n15120) );
  AND U12473 ( .A(n5204), .B(n15120), .Z(n5205) );
  NANDN U12474 ( .A(n15123), .B(n5205), .Z(n5206) );
  NANDN U12475 ( .A(y[200]), .B(x[200]), .Z(n15122) );
  AND U12476 ( .A(n5206), .B(n15122), .Z(n5207) );
  NAND U12477 ( .A(n15118), .B(n5207), .Z(n5208) );
  NANDN U12478 ( .A(n15119), .B(n5208), .Z(n5209) );
  ANDN U12479 ( .B(y[202]), .A(x[202]), .Z(n15115) );
  OR U12480 ( .A(n5209), .B(n15115), .Z(n5210) );
  AND U12481 ( .A(n5211), .B(n5210), .Z(n5213) );
  NANDN U12482 ( .A(x[204]), .B(y[204]), .Z(n15112) );
  NANDN U12483 ( .A(x[203]), .B(y[203]), .Z(n15116) );
  AND U12484 ( .A(n15112), .B(n15116), .Z(n5212) );
  NANDN U12485 ( .A(n5213), .B(n5212), .Z(n5214) );
  AND U12486 ( .A(n15113), .B(n5214), .Z(n5215) );
  NANDN U12487 ( .A(y[205]), .B(x[205]), .Z(n15109) );
  NAND U12488 ( .A(n5215), .B(n15109), .Z(n5216) );
  ANDN U12489 ( .B(y[206]), .A(x[206]), .Z(n15106) );
  ANDN U12490 ( .B(n5216), .A(n15106), .Z(n5217) );
  NANDN U12491 ( .A(n15111), .B(n5217), .Z(n5218) );
  NANDN U12492 ( .A(y[206]), .B(x[206]), .Z(n15110) );
  AND U12493 ( .A(n5218), .B(n15110), .Z(n5219) );
  NAND U12494 ( .A(n15104), .B(n5219), .Z(n5220) );
  NAND U12495 ( .A(n15108), .B(n5220), .Z(n5221) );
  NANDN U12496 ( .A(x[208]), .B(y[208]), .Z(n15103) );
  NANDN U12497 ( .A(n5221), .B(n15103), .Z(n5222) );
  AND U12498 ( .A(n5223), .B(n5222), .Z(n5225) );
  NANDN U12499 ( .A(x[210]), .B(y[210]), .Z(n15100) );
  ANDN U12500 ( .B(y[209]), .A(x[209]), .Z(n15102) );
  ANDN U12501 ( .B(n15100), .A(n15102), .Z(n5224) );
  NANDN U12502 ( .A(n5225), .B(n5224), .Z(n5226) );
  AND U12503 ( .A(n5227), .B(n5226), .Z(n5228) );
  NANDN U12504 ( .A(y[211]), .B(x[211]), .Z(n15097) );
  NAND U12505 ( .A(n5228), .B(n15097), .Z(n5229) );
  NANDN U12506 ( .A(x[212]), .B(y[212]), .Z(n15096) );
  AND U12507 ( .A(n5229), .B(n15096), .Z(n5230) );
  NANDN U12508 ( .A(n15099), .B(n5230), .Z(n5231) );
  NANDN U12509 ( .A(y[212]), .B(x[212]), .Z(n15098) );
  AND U12510 ( .A(n5231), .B(n15098), .Z(n5232) );
  NAND U12511 ( .A(n15094), .B(n5232), .Z(n5233) );
  NANDN U12512 ( .A(n15095), .B(n5233), .Z(n5234) );
  ANDN U12513 ( .B(y[214]), .A(x[214]), .Z(n15091) );
  OR U12514 ( .A(n5234), .B(n15091), .Z(n5235) );
  AND U12515 ( .A(n5236), .B(n5235), .Z(n5238) );
  NANDN U12516 ( .A(x[216]), .B(y[216]), .Z(n15088) );
  NANDN U12517 ( .A(x[215]), .B(y[215]), .Z(n15092) );
  AND U12518 ( .A(n15088), .B(n15092), .Z(n5237) );
  NANDN U12519 ( .A(n5238), .B(n5237), .Z(n5239) );
  AND U12520 ( .A(n15089), .B(n5239), .Z(n5240) );
  NANDN U12521 ( .A(y[217]), .B(x[217]), .Z(n15085) );
  NAND U12522 ( .A(n5240), .B(n15085), .Z(n5241) );
  NANDN U12523 ( .A(x[218]), .B(y[218]), .Z(n15084) );
  AND U12524 ( .A(n5241), .B(n15084), .Z(n5242) );
  NANDN U12525 ( .A(n15087), .B(n5242), .Z(n5243) );
  NANDN U12526 ( .A(y[218]), .B(x[218]), .Z(n15086) );
  AND U12527 ( .A(n5243), .B(n15086), .Z(n5244) );
  NAND U12528 ( .A(n15081), .B(n5244), .Z(n5245) );
  NANDN U12529 ( .A(n15083), .B(n5245), .Z(n5246) );
  ANDN U12530 ( .B(y[220]), .A(x[220]), .Z(n15079) );
  OR U12531 ( .A(n5246), .B(n15079), .Z(n5247) );
  AND U12532 ( .A(n5248), .B(n5247), .Z(n5250) );
  NANDN U12533 ( .A(x[221]), .B(y[221]), .Z(n15080) );
  ANDN U12534 ( .B(y[222]), .A(x[222]), .Z(n15075) );
  ANDN U12535 ( .B(n15080), .A(n15075), .Z(n5249) );
  NANDN U12536 ( .A(n5250), .B(n5249), .Z(n5251) );
  AND U12537 ( .A(n15078), .B(n5251), .Z(n5252) );
  NANDN U12538 ( .A(y[223]), .B(x[223]), .Z(n15073) );
  NAND U12539 ( .A(n5252), .B(n15073), .Z(n5253) );
  ANDN U12540 ( .B(y[224]), .A(x[224]), .Z(n15071) );
  ANDN U12541 ( .B(n5253), .A(n15071), .Z(n5254) );
  NAND U12542 ( .A(n15076), .B(n5254), .Z(n5255) );
  NANDN U12543 ( .A(y[224]), .B(x[224]), .Z(n15074) );
  AND U12544 ( .A(n5255), .B(n15074), .Z(n5256) );
  NAND U12545 ( .A(n15069), .B(n5256), .Z(n5257) );
  NAND U12546 ( .A(n15072), .B(n5257), .Z(n5258) );
  NANDN U12547 ( .A(x[226]), .B(y[226]), .Z(n15068) );
  NANDN U12548 ( .A(n5258), .B(n15068), .Z(n5259) );
  AND U12549 ( .A(n5260), .B(n5259), .Z(n5262) );
  NANDN U12550 ( .A(x[228]), .B(y[228]), .Z(n15063) );
  ANDN U12551 ( .B(y[227]), .A(x[227]), .Z(n15066) );
  ANDN U12552 ( .B(n15063), .A(n15066), .Z(n5261) );
  NANDN U12553 ( .A(n5262), .B(n5261), .Z(n5263) );
  AND U12554 ( .A(n15064), .B(n5263), .Z(n5264) );
  NAND U12555 ( .A(n15061), .B(n5264), .Z(n5265) );
  NANDN U12556 ( .A(x[230]), .B(y[230]), .Z(n15060) );
  AND U12557 ( .A(n5265), .B(n15060), .Z(n5266) );
  NANDN U12558 ( .A(n15062), .B(n5266), .Z(n5268) );
  NANDN U12559 ( .A(y[230]), .B(x[230]), .Z(n5267) );
  AND U12560 ( .A(n5268), .B(n5267), .Z(n5269) );
  NAND U12561 ( .A(n15058), .B(n5269), .Z(n5270) );
  NANDN U12562 ( .A(n15059), .B(n5270), .Z(n5271) );
  ANDN U12563 ( .B(y[232]), .A(x[232]), .Z(n15055) );
  OR U12564 ( .A(n5271), .B(n15055), .Z(n5272) );
  AND U12565 ( .A(n5273), .B(n5272), .Z(n5275) );
  NANDN U12566 ( .A(x[234]), .B(y[234]), .Z(n15052) );
  NANDN U12567 ( .A(x[233]), .B(y[233]), .Z(n15056) );
  AND U12568 ( .A(n15052), .B(n15056), .Z(n5274) );
  NANDN U12569 ( .A(n5275), .B(n5274), .Z(n5276) );
  AND U12570 ( .A(n15054), .B(n5276), .Z(n5277) );
  NANDN U12571 ( .A(y[235]), .B(x[235]), .Z(n15050) );
  NAND U12572 ( .A(n5277), .B(n15050), .Z(n5278) );
  NANDN U12573 ( .A(x[236]), .B(y[236]), .Z(n15048) );
  AND U12574 ( .A(n5278), .B(n15048), .Z(n5279) );
  NANDN U12575 ( .A(n15051), .B(n5279), .Z(n5280) );
  NANDN U12576 ( .A(y[236]), .B(x[236]), .Z(n15049) );
  AND U12577 ( .A(n5280), .B(n15049), .Z(n5281) );
  NAND U12578 ( .A(n15045), .B(n5281), .Z(n5282) );
  NANDN U12579 ( .A(n15047), .B(n5282), .Z(n5283) );
  NANDN U12580 ( .A(x[238]), .B(y[238]), .Z(n15044) );
  NANDN U12581 ( .A(n5283), .B(n15044), .Z(n5284) );
  AND U12582 ( .A(n5285), .B(n5284), .Z(n5287) );
  NANDN U12583 ( .A(x[240]), .B(y[240]), .Z(n15039) );
  ANDN U12584 ( .B(y[239]), .A(x[239]), .Z(n15043) );
  ANDN U12585 ( .B(n15039), .A(n15043), .Z(n5286) );
  NANDN U12586 ( .A(n5287), .B(n5286), .Z(n5288) );
  AND U12587 ( .A(n15041), .B(n5288), .Z(n5289) );
  NAND U12588 ( .A(n15038), .B(n5289), .Z(n5290) );
  NANDN U12589 ( .A(x[242]), .B(y[242]), .Z(n15037) );
  AND U12590 ( .A(n5290), .B(n15037), .Z(n5291) );
  NAND U12591 ( .A(n15040), .B(n5291), .Z(n5293) );
  NANDN U12592 ( .A(y[242]), .B(x[242]), .Z(n5292) );
  AND U12593 ( .A(n5293), .B(n5292), .Z(n5294) );
  NAND U12594 ( .A(n15035), .B(n5294), .Z(n5295) );
  NANDN U12595 ( .A(n15036), .B(n5295), .Z(n5296) );
  NANDN U12596 ( .A(x[244]), .B(y[244]), .Z(n15033) );
  NANDN U12597 ( .A(n5296), .B(n15033), .Z(n5297) );
  AND U12598 ( .A(n5298), .B(n5297), .Z(n5300) );
  NANDN U12599 ( .A(x[246]), .B(y[246]), .Z(n15028) );
  ANDN U12600 ( .B(y[245]), .A(x[245]), .Z(n15032) );
  ANDN U12601 ( .B(n15028), .A(n15032), .Z(n5299) );
  NANDN U12602 ( .A(n5300), .B(n5299), .Z(n5301) );
  AND U12603 ( .A(n15031), .B(n5301), .Z(n5302) );
  NANDN U12604 ( .A(y[247]), .B(x[247]), .Z(n15027) );
  NAND U12605 ( .A(n5302), .B(n15027), .Z(n5303) );
  ANDN U12606 ( .B(y[248]), .A(x[248]), .Z(n15024) );
  ANDN U12607 ( .B(n5303), .A(n15024), .Z(n5304) );
  NAND U12608 ( .A(n15029), .B(n5304), .Z(n5305) );
  NANDN U12609 ( .A(y[248]), .B(x[248]), .Z(n15026) );
  AND U12610 ( .A(n5305), .B(n15026), .Z(n5306) );
  NAND U12611 ( .A(n15022), .B(n5306), .Z(n5307) );
  NAND U12612 ( .A(n15025), .B(n5307), .Z(n5308) );
  NANDN U12613 ( .A(x[250]), .B(y[250]), .Z(n15021) );
  NANDN U12614 ( .A(n5308), .B(n15021), .Z(n5309) );
  AND U12615 ( .A(n5310), .B(n5309), .Z(n5312) );
  NANDN U12616 ( .A(x[252]), .B(y[252]), .Z(n15017) );
  ANDN U12617 ( .B(y[251]), .A(x[251]), .Z(n15020) );
  ANDN U12618 ( .B(n15017), .A(n15020), .Z(n5311) );
  NANDN U12619 ( .A(n5312), .B(n5311), .Z(n5313) );
  AND U12620 ( .A(n15019), .B(n5313), .Z(n5314) );
  NAND U12621 ( .A(n15015), .B(n5314), .Z(n5315) );
  NANDN U12622 ( .A(x[254]), .B(y[254]), .Z(n15014) );
  AND U12623 ( .A(n5315), .B(n15014), .Z(n5316) );
  NANDN U12624 ( .A(n15016), .B(n5316), .Z(n5318) );
  NANDN U12625 ( .A(y[254]), .B(x[254]), .Z(n5317) );
  AND U12626 ( .A(n5318), .B(n5317), .Z(n5319) );
  NAND U12627 ( .A(n15011), .B(n5319), .Z(n5320) );
  NANDN U12628 ( .A(n15013), .B(n5320), .Z(n5321) );
  NANDN U12629 ( .A(x[256]), .B(y[256]), .Z(n15010) );
  NANDN U12630 ( .A(n5321), .B(n15010), .Z(n5322) );
  AND U12631 ( .A(n5323), .B(n5322), .Z(n5325) );
  NANDN U12632 ( .A(x[258]), .B(y[258]), .Z(n15006) );
  ANDN U12633 ( .B(y[257]), .A(x[257]), .Z(n15009) );
  ANDN U12634 ( .B(n15006), .A(n15009), .Z(n5324) );
  NANDN U12635 ( .A(n5325), .B(n5324), .Z(n5326) );
  AND U12636 ( .A(n15008), .B(n5326), .Z(n5327) );
  NAND U12637 ( .A(n15004), .B(n5327), .Z(n5328) );
  NANDN U12638 ( .A(x[260]), .B(y[260]), .Z(n15003) );
  AND U12639 ( .A(n5328), .B(n15003), .Z(n5329) );
  NANDN U12640 ( .A(n15005), .B(n5329), .Z(n5331) );
  NANDN U12641 ( .A(y[260]), .B(x[260]), .Z(n5330) );
  AND U12642 ( .A(n5331), .B(n5330), .Z(n5332) );
  NAND U12643 ( .A(n15000), .B(n5332), .Z(n5333) );
  NANDN U12644 ( .A(n15002), .B(n5333), .Z(n5335) );
  NANDN U12645 ( .A(x[262]), .B(n5335), .Z(n5334) );
  ANDN U12646 ( .B(y[263]), .A(x[263]), .Z(n14999) );
  ANDN U12647 ( .B(n5334), .A(n14999), .Z(n5338) );
  XNOR U12648 ( .A(n5335), .B(x[262]), .Z(n5336) );
  NAND U12649 ( .A(n5336), .B(y[262]), .Z(n5337) );
  NAND U12650 ( .A(n5338), .B(n5337), .Z(n5339) );
  NAND U12651 ( .A(n15760), .B(n5339), .Z(n5340) );
  NANDN U12652 ( .A(n14998), .B(n5340), .Z(n5343) );
  NANDN U12653 ( .A(y[266]), .B(x[266]), .Z(n5342) );
  NANDN U12654 ( .A(y[265]), .B(x[265]), .Z(n5341) );
  AND U12655 ( .A(n5342), .B(n5341), .Z(n14997) );
  AND U12656 ( .A(n5343), .B(n14997), .Z(n5346) );
  NANDN U12657 ( .A(x[266]), .B(y[266]), .Z(n5345) );
  NANDN U12658 ( .A(x[267]), .B(y[267]), .Z(n5344) );
  NAND U12659 ( .A(n5345), .B(n5344), .Z(n14996) );
  OR U12660 ( .A(n5346), .B(n14996), .Z(n5347) );
  NAND U12661 ( .A(n14995), .B(n5347), .Z(n5348) );
  NANDN U12662 ( .A(n15766), .B(n5348), .Z(n5349) );
  NAND U12663 ( .A(n15768), .B(n5349), .Z(n5350) );
  NANDN U12664 ( .A(n14994), .B(n5350), .Z(n5351) );
  AND U12665 ( .A(n14992), .B(n5351), .Z(n5352) );
  NANDN U12666 ( .A(x[272]), .B(y[272]), .Z(n14991) );
  NANDN U12667 ( .A(n5352), .B(n14991), .Z(n5353) );
  AND U12668 ( .A(n5354), .B(n5353), .Z(n5356) );
  NANDN U12669 ( .A(x[274]), .B(y[274]), .Z(n14987) );
  ANDN U12670 ( .B(y[273]), .A(x[273]), .Z(n14990) );
  ANDN U12671 ( .B(n14987), .A(n14990), .Z(n5355) );
  NANDN U12672 ( .A(n5356), .B(n5355), .Z(n5357) );
  AND U12673 ( .A(n14989), .B(n5357), .Z(n5358) );
  NANDN U12674 ( .A(y[275]), .B(x[275]), .Z(n14985) );
  NAND U12675 ( .A(n5358), .B(n14985), .Z(n5359) );
  ANDN U12676 ( .B(y[276]), .A(x[276]), .Z(n14982) );
  ANDN U12677 ( .B(n5359), .A(n14982), .Z(n5360) );
  NANDN U12678 ( .A(n14986), .B(n5360), .Z(n5361) );
  NANDN U12679 ( .A(y[276]), .B(x[276]), .Z(n14984) );
  AND U12680 ( .A(n5361), .B(n14984), .Z(n5362) );
  NAND U12681 ( .A(n14981), .B(n5362), .Z(n5363) );
  NAND U12682 ( .A(n14983), .B(n5363), .Z(n5364) );
  NANDN U12683 ( .A(x[278]), .B(y[278]), .Z(n14980) );
  NANDN U12684 ( .A(n5364), .B(n14980), .Z(n5365) );
  AND U12685 ( .A(n5366), .B(n5365), .Z(n5368) );
  NANDN U12686 ( .A(x[280]), .B(y[280]), .Z(n14976) );
  ANDN U12687 ( .B(y[279]), .A(x[279]), .Z(n14979) );
  ANDN U12688 ( .B(n14976), .A(n14979), .Z(n5367) );
  NANDN U12689 ( .A(n5368), .B(n5367), .Z(n5369) );
  AND U12690 ( .A(n14978), .B(n5369), .Z(n5370) );
  NANDN U12691 ( .A(y[281]), .B(x[281]), .Z(n14973) );
  NAND U12692 ( .A(n5370), .B(n14973), .Z(n5371) );
  NANDN U12693 ( .A(x[282]), .B(y[282]), .Z(n14972) );
  AND U12694 ( .A(n5371), .B(n14972), .Z(n5372) );
  NANDN U12695 ( .A(n14975), .B(n5372), .Z(n5373) );
  NANDN U12696 ( .A(y[282]), .B(x[282]), .Z(n14974) );
  AND U12697 ( .A(n5373), .B(n14974), .Z(n5374) );
  NAND U12698 ( .A(n14969), .B(n5374), .Z(n5375) );
  NANDN U12699 ( .A(n14971), .B(n5375), .Z(n5376) );
  NANDN U12700 ( .A(x[284]), .B(y[284]), .Z(n14968) );
  NANDN U12701 ( .A(n5376), .B(n14968), .Z(n5377) );
  AND U12702 ( .A(n5378), .B(n5377), .Z(n5380) );
  NANDN U12703 ( .A(x[286]), .B(y[286]), .Z(n14964) );
  ANDN U12704 ( .B(y[285]), .A(x[285]), .Z(n14967) );
  ANDN U12705 ( .B(n14964), .A(n14967), .Z(n5379) );
  NANDN U12706 ( .A(n5380), .B(n5379), .Z(n5381) );
  AND U12707 ( .A(n14966), .B(n5381), .Z(n5382) );
  NAND U12708 ( .A(n14959), .B(n5382), .Z(n5383) );
  NANDN U12709 ( .A(x[288]), .B(y[288]), .Z(n14958) );
  AND U12710 ( .A(n5383), .B(n14958), .Z(n5384) );
  NANDN U12711 ( .A(n14962), .B(n5384), .Z(n5386) );
  NANDN U12712 ( .A(y[288]), .B(x[288]), .Z(n5385) );
  AND U12713 ( .A(n5386), .B(n5385), .Z(n5387) );
  NAND U12714 ( .A(n14956), .B(n5387), .Z(n5388) );
  NANDN U12715 ( .A(n14957), .B(n5388), .Z(n5389) );
  NANDN U12716 ( .A(x[290]), .B(y[290]), .Z(n14954) );
  NANDN U12717 ( .A(n5389), .B(n14954), .Z(n5390) );
  AND U12718 ( .A(n5391), .B(n5390), .Z(n5393) );
  NANDN U12719 ( .A(x[292]), .B(y[292]), .Z(n14949) );
  ANDN U12720 ( .B(y[291]), .A(x[291]), .Z(n14953) );
  ANDN U12721 ( .B(n14949), .A(n14953), .Z(n5392) );
  NANDN U12722 ( .A(n5393), .B(n5392), .Z(n5394) );
  AND U12723 ( .A(n14952), .B(n5394), .Z(n5395) );
  NANDN U12724 ( .A(y[293]), .B(x[293]), .Z(n14948) );
  NAND U12725 ( .A(n5395), .B(n14948), .Z(n5396) );
  ANDN U12726 ( .B(y[294]), .A(x[294]), .Z(n14945) );
  ANDN U12727 ( .B(n5396), .A(n14945), .Z(n5397) );
  NAND U12728 ( .A(n14950), .B(n5397), .Z(n5398) );
  NANDN U12729 ( .A(y[294]), .B(x[294]), .Z(n14947) );
  AND U12730 ( .A(n5398), .B(n14947), .Z(n5399) );
  NAND U12731 ( .A(n14944), .B(n5399), .Z(n5400) );
  NAND U12732 ( .A(n14946), .B(n5400), .Z(n5401) );
  NANDN U12733 ( .A(x[296]), .B(y[296]), .Z(n14943) );
  NANDN U12734 ( .A(n5401), .B(n14943), .Z(n5402) );
  AND U12735 ( .A(n5403), .B(n5402), .Z(n5405) );
  NANDN U12736 ( .A(x[298]), .B(y[298]), .Z(n14938) );
  ANDN U12737 ( .B(y[297]), .A(x[297]), .Z(n14942) );
  ANDN U12738 ( .B(n14938), .A(n14942), .Z(n5404) );
  NANDN U12739 ( .A(n5405), .B(n5404), .Z(n5406) );
  AND U12740 ( .A(n14940), .B(n5406), .Z(n5407) );
  NANDN U12741 ( .A(y[299]), .B(x[299]), .Z(n14937) );
  NAND U12742 ( .A(n5407), .B(n14937), .Z(n5408) );
  ANDN U12743 ( .B(y[300]), .A(x[300]), .Z(n14934) );
  ANDN U12744 ( .B(n5408), .A(n14934), .Z(n5409) );
  NAND U12745 ( .A(n14939), .B(n5409), .Z(n5410) );
  NANDN U12746 ( .A(y[300]), .B(x[300]), .Z(n14936) );
  AND U12747 ( .A(n5410), .B(n14936), .Z(n5411) );
  NAND U12748 ( .A(n14933), .B(n5411), .Z(n5412) );
  NAND U12749 ( .A(n14935), .B(n5412), .Z(n5413) );
  NANDN U12750 ( .A(x[302]), .B(y[302]), .Z(n14932) );
  NANDN U12751 ( .A(n5413), .B(n14932), .Z(n5414) );
  AND U12752 ( .A(n5415), .B(n5414), .Z(n5417) );
  NANDN U12753 ( .A(x[304]), .B(y[304]), .Z(n14928) );
  ANDN U12754 ( .B(y[303]), .A(x[303]), .Z(n14931) );
  ANDN U12755 ( .B(n14928), .A(n14931), .Z(n5416) );
  NANDN U12756 ( .A(n5417), .B(n5416), .Z(n5418) );
  AND U12757 ( .A(n14929), .B(n5418), .Z(n5419) );
  NAND U12758 ( .A(n14926), .B(n5419), .Z(n5420) );
  NANDN U12759 ( .A(x[306]), .B(y[306]), .Z(n14925) );
  AND U12760 ( .A(n5420), .B(n14925), .Z(n5421) );
  NANDN U12761 ( .A(n14927), .B(n5421), .Z(n5423) );
  NANDN U12762 ( .A(y[306]), .B(x[306]), .Z(n5422) );
  AND U12763 ( .A(n5423), .B(n5422), .Z(n5424) );
  NAND U12764 ( .A(n14920), .B(n5424), .Z(n5425) );
  NANDN U12765 ( .A(n14923), .B(n5425), .Z(n5426) );
  NANDN U12766 ( .A(x[308]), .B(y[308]), .Z(n14919) );
  NANDN U12767 ( .A(n5426), .B(n14919), .Z(n5427) );
  AND U12768 ( .A(n5428), .B(n5427), .Z(n5430) );
  NANDN U12769 ( .A(x[310]), .B(y[310]), .Z(n14914) );
  ANDN U12770 ( .B(y[309]), .A(x[309]), .Z(n14918) );
  ANDN U12771 ( .B(n14914), .A(n14918), .Z(n5429) );
  NANDN U12772 ( .A(n5430), .B(n5429), .Z(n5431) );
  AND U12773 ( .A(n14916), .B(n5431), .Z(n5432) );
  NANDN U12774 ( .A(y[311]), .B(x[311]), .Z(n14912) );
  NAND U12775 ( .A(n5432), .B(n14912), .Z(n5433) );
  NANDN U12776 ( .A(x[312]), .B(y[312]), .Z(n14911) );
  AND U12777 ( .A(n5433), .B(n14911), .Z(n5434) );
  NAND U12778 ( .A(n14915), .B(n5434), .Z(n5435) );
  NANDN U12779 ( .A(y[312]), .B(x[312]), .Z(n14913) );
  AND U12780 ( .A(n5435), .B(n14913), .Z(n5436) );
  NAND U12781 ( .A(n14908), .B(n5436), .Z(n5437) );
  NANDN U12782 ( .A(n14909), .B(n5437), .Z(n5438) );
  ANDN U12783 ( .B(y[314]), .A(x[314]), .Z(n14905) );
  OR U12784 ( .A(n5438), .B(n14905), .Z(n5439) );
  AND U12785 ( .A(n5440), .B(n5439), .Z(n5442) );
  NANDN U12786 ( .A(x[315]), .B(y[315]), .Z(n14906) );
  ANDN U12787 ( .B(y[316]), .A(x[316]), .Z(n14901) );
  ANDN U12788 ( .B(n14906), .A(n14901), .Z(n5441) );
  NANDN U12789 ( .A(n5442), .B(n5441), .Z(n5443) );
  AND U12790 ( .A(n14903), .B(n5443), .Z(n5444) );
  NANDN U12791 ( .A(y[317]), .B(x[317]), .Z(n14900) );
  NAND U12792 ( .A(n5444), .B(n14900), .Z(n5445) );
  NANDN U12793 ( .A(x[317]), .B(y[317]), .Z(n14902) );
  AND U12794 ( .A(n5445), .B(n14902), .Z(n5446) );
  NANDN U12795 ( .A(n14899), .B(n5446), .Z(n5448) );
  NANDN U12796 ( .A(y[318]), .B(x[318]), .Z(n5447) );
  AND U12797 ( .A(n5448), .B(n5447), .Z(n5449) );
  NAND U12798 ( .A(n14897), .B(n5449), .Z(n5450) );
  NANDN U12799 ( .A(n14898), .B(n5450), .Z(n5451) );
  NANDN U12800 ( .A(x[320]), .B(y[320]), .Z(n14896) );
  NANDN U12801 ( .A(n5451), .B(n14896), .Z(n5452) );
  AND U12802 ( .A(n5453), .B(n5452), .Z(n5455) );
  NANDN U12803 ( .A(x[322]), .B(y[322]), .Z(n14891) );
  ANDN U12804 ( .B(y[321]), .A(x[321]), .Z(n14895) );
  ANDN U12805 ( .B(n14891), .A(n14895), .Z(n5454) );
  NANDN U12806 ( .A(n5455), .B(n5454), .Z(n5456) );
  AND U12807 ( .A(n14893), .B(n5456), .Z(n5457) );
  NANDN U12808 ( .A(y[323]), .B(x[323]), .Z(n14890) );
  NAND U12809 ( .A(n5457), .B(n14890), .Z(n5458) );
  NANDN U12810 ( .A(x[323]), .B(y[323]), .Z(n14892) );
  AND U12811 ( .A(n5458), .B(n14892), .Z(n5459) );
  NANDN U12812 ( .A(n14889), .B(n5459), .Z(n5461) );
  NANDN U12813 ( .A(y[324]), .B(x[324]), .Z(n5460) );
  AND U12814 ( .A(n5461), .B(n5460), .Z(n5462) );
  NAND U12815 ( .A(n14886), .B(n5462), .Z(n5463) );
  NANDN U12816 ( .A(n14888), .B(n5463), .Z(n5464) );
  NANDN U12817 ( .A(x[326]), .B(y[326]), .Z(n14885) );
  NANDN U12818 ( .A(n5464), .B(n14885), .Z(n5465) );
  AND U12819 ( .A(n5466), .B(n5465), .Z(n5468) );
  NANDN U12820 ( .A(x[328]), .B(y[328]), .Z(n14881) );
  ANDN U12821 ( .B(y[327]), .A(x[327]), .Z(n14884) );
  ANDN U12822 ( .B(n14881), .A(n14884), .Z(n5467) );
  NANDN U12823 ( .A(n5468), .B(n5467), .Z(n5469) );
  AND U12824 ( .A(n14882), .B(n5469), .Z(n5470) );
  NANDN U12825 ( .A(y[329]), .B(x[329]), .Z(n14878) );
  NAND U12826 ( .A(n5470), .B(n14878), .Z(n5471) );
  NANDN U12827 ( .A(x[330]), .B(y[330]), .Z(n14877) );
  AND U12828 ( .A(n5471), .B(n14877), .Z(n5472) );
  NANDN U12829 ( .A(n14880), .B(n5472), .Z(n5473) );
  NANDN U12830 ( .A(y[330]), .B(x[330]), .Z(n14879) );
  AND U12831 ( .A(n5473), .B(n14879), .Z(n5474) );
  NAND U12832 ( .A(n14875), .B(n5474), .Z(n5475) );
  NANDN U12833 ( .A(n14876), .B(n5475), .Z(n5476) );
  ANDN U12834 ( .B(y[332]), .A(x[332]), .Z(n14872) );
  OR U12835 ( .A(n5476), .B(n14872), .Z(n5477) );
  AND U12836 ( .A(n5478), .B(n5477), .Z(n5480) );
  NANDN U12837 ( .A(x[334]), .B(y[334]), .Z(n14869) );
  NANDN U12838 ( .A(x[333]), .B(y[333]), .Z(n14873) );
  AND U12839 ( .A(n14869), .B(n14873), .Z(n5479) );
  NANDN U12840 ( .A(n5480), .B(n5479), .Z(n5481) );
  AND U12841 ( .A(n14870), .B(n5481), .Z(n5482) );
  NANDN U12842 ( .A(y[335]), .B(x[335]), .Z(n14866) );
  NAND U12843 ( .A(n5482), .B(n14866), .Z(n5483) );
  ANDN U12844 ( .B(y[336]), .A(x[336]), .Z(n14865) );
  ANDN U12845 ( .B(n5483), .A(n14865), .Z(n5484) );
  NANDN U12846 ( .A(n14868), .B(n5484), .Z(n5485) );
  NAND U12847 ( .A(n14867), .B(n5485), .Z(n5487) );
  NANDN U12848 ( .A(y[337]), .B(n5487), .Z(n5486) );
  ANDN U12849 ( .B(x[338]), .A(y[338]), .Z(n14864) );
  ANDN U12850 ( .B(n5486), .A(n14864), .Z(n5490) );
  XNOR U12851 ( .A(n5487), .B(y[337]), .Z(n5488) );
  NAND U12852 ( .A(n5488), .B(x[337]), .Z(n5489) );
  NAND U12853 ( .A(n5490), .B(n5489), .Z(n5491) );
  NAND U12854 ( .A(n25211), .B(n5491), .Z(n5492) );
  NANDN U12855 ( .A(n25213), .B(n5492), .Z(n5493) );
  AND U12856 ( .A(n25215), .B(n5493), .Z(n5494) );
  ANDN U12857 ( .B(x[341]), .A(y[341]), .Z(n14862) );
  OR U12858 ( .A(n5494), .B(n14862), .Z(n5495) );
  NAND U12859 ( .A(n14861), .B(n5495), .Z(n5496) );
  NAND U12860 ( .A(n14863), .B(n5496), .Z(n5497) );
  ANDN U12861 ( .B(x[343]), .A(y[343]), .Z(n14858) );
  OR U12862 ( .A(n5497), .B(n14858), .Z(n5498) );
  AND U12863 ( .A(n5499), .B(n5498), .Z(n5501) );
  NANDN U12864 ( .A(y[344]), .B(x[344]), .Z(n14859) );
  ANDN U12865 ( .B(x[345]), .A(y[345]), .Z(n14854) );
  ANDN U12866 ( .B(n14859), .A(n14854), .Z(n5500) );
  NANDN U12867 ( .A(n5501), .B(n5500), .Z(n5502) );
  AND U12868 ( .A(n14857), .B(n5502), .Z(n5503) );
  NANDN U12869 ( .A(x[346]), .B(y[346]), .Z(n14852) );
  NAND U12870 ( .A(n5503), .B(n14852), .Z(n5504) );
  ANDN U12871 ( .B(x[347]), .A(y[347]), .Z(n14850) );
  ANDN U12872 ( .B(n5504), .A(n14850), .Z(n5505) );
  NAND U12873 ( .A(n14855), .B(n5505), .Z(n5506) );
  NANDN U12874 ( .A(x[347]), .B(y[347]), .Z(n14853) );
  AND U12875 ( .A(n5506), .B(n14853), .Z(n5507) );
  NAND U12876 ( .A(n14849), .B(n5507), .Z(n5508) );
  NAND U12877 ( .A(n14851), .B(n5508), .Z(n5509) );
  ANDN U12878 ( .B(x[349]), .A(y[349]), .Z(n14846) );
  OR U12879 ( .A(n5509), .B(n14846), .Z(n5510) );
  AND U12880 ( .A(n5511), .B(n5510), .Z(n5513) );
  NANDN U12881 ( .A(y[350]), .B(x[350]), .Z(n14847) );
  NANDN U12882 ( .A(y[351]), .B(x[351]), .Z(n25236) );
  AND U12883 ( .A(n14847), .B(n25236), .Z(n5512) );
  NANDN U12884 ( .A(n5513), .B(n5512), .Z(n5514) );
  XNOR U12885 ( .A(x[352]), .B(y[352]), .Z(n25235) );
  AND U12886 ( .A(n5514), .B(n25235), .Z(n5515) );
  NANDN U12887 ( .A(x[351]), .B(y[351]), .Z(n15850) );
  NAND U12888 ( .A(n5515), .B(n15850), .Z(n5516) );
  ANDN U12889 ( .B(x[353]), .A(y[353]), .Z(n14843) );
  ANDN U12890 ( .B(n5516), .A(n14843), .Z(n5517) );
  NAND U12891 ( .A(n15854), .B(n5517), .Z(n5518) );
  NANDN U12892 ( .A(x[353]), .B(y[353]), .Z(n14844) );
  AND U12893 ( .A(n5518), .B(n14844), .Z(n5519) );
  NAND U12894 ( .A(n14841), .B(n5519), .Z(n5520) );
  NANDN U12895 ( .A(n5521), .B(n5520), .Z(n5522) );
  ANDN U12896 ( .B(x[355]), .A(y[355]), .Z(n14838) );
  OR U12897 ( .A(n5522), .B(n14838), .Z(n5523) );
  AND U12898 ( .A(n5524), .B(n5523), .Z(n5526) );
  NANDN U12899 ( .A(y[357]), .B(x[357]), .Z(n14835) );
  NANDN U12900 ( .A(y[356]), .B(x[356]), .Z(n14839) );
  AND U12901 ( .A(n14835), .B(n14839), .Z(n5525) );
  NANDN U12902 ( .A(n5526), .B(n5525), .Z(n5527) );
  AND U12903 ( .A(n14837), .B(n5527), .Z(n5528) );
  NANDN U12904 ( .A(x[358]), .B(y[358]), .Z(n14832) );
  NAND U12905 ( .A(n5528), .B(n14832), .Z(n5529) );
  ANDN U12906 ( .B(x[359]), .A(y[359]), .Z(n14831) );
  ANDN U12907 ( .B(n5529), .A(n14831), .Z(n5530) );
  NANDN U12908 ( .A(n14834), .B(n5530), .Z(n5531) );
  NANDN U12909 ( .A(x[359]), .B(y[359]), .Z(n14833) );
  AND U12910 ( .A(n5531), .B(n14833), .Z(n5532) );
  NAND U12911 ( .A(n14829), .B(n5532), .Z(n5533) );
  NANDN U12912 ( .A(n5534), .B(n5533), .Z(n5535) );
  ANDN U12913 ( .B(x[361]), .A(y[361]), .Z(n14827) );
  OR U12914 ( .A(n5535), .B(n14827), .Z(n5536) );
  AND U12915 ( .A(n5537), .B(n5536), .Z(n5540) );
  NANDN U12916 ( .A(y[363]), .B(x[363]), .Z(n14823) );
  ANDN U12917 ( .B(x[362]), .A(y[362]), .Z(n5538) );
  ANDN U12918 ( .B(n14823), .A(n5538), .Z(n5539) );
  NANDN U12919 ( .A(n5540), .B(n5539), .Z(n5541) );
  AND U12920 ( .A(n14824), .B(n5541), .Z(n5542) );
  NANDN U12921 ( .A(x[364]), .B(y[364]), .Z(n14821) );
  NAND U12922 ( .A(n5542), .B(n14821), .Z(n5543) );
  NANDN U12923 ( .A(y[365]), .B(x[365]), .Z(n14819) );
  AND U12924 ( .A(n5543), .B(n14819), .Z(n5544) );
  NANDN U12925 ( .A(n14822), .B(n5544), .Z(n5545) );
  NANDN U12926 ( .A(x[365]), .B(y[365]), .Z(n14820) );
  AND U12927 ( .A(n5545), .B(n14820), .Z(n5546) );
  NAND U12928 ( .A(n14817), .B(n5546), .Z(n5547) );
  NANDN U12929 ( .A(n14818), .B(n5547), .Z(n5548) );
  ANDN U12930 ( .B(x[367]), .A(y[367]), .Z(n14815) );
  OR U12931 ( .A(n5548), .B(n14815), .Z(n5549) );
  AND U12932 ( .A(n5550), .B(n5549), .Z(n5553) );
  NANDN U12933 ( .A(y[369]), .B(x[369]), .Z(n14811) );
  ANDN U12934 ( .B(x[368]), .A(y[368]), .Z(n5551) );
  ANDN U12935 ( .B(n14811), .A(n5551), .Z(n5552) );
  NANDN U12936 ( .A(n5553), .B(n5552), .Z(n5554) );
  AND U12937 ( .A(n14812), .B(n5554), .Z(n5555) );
  NANDN U12938 ( .A(x[370]), .B(y[370]), .Z(n14809) );
  NAND U12939 ( .A(n5555), .B(n14809), .Z(n5556) );
  NANDN U12940 ( .A(y[371]), .B(x[371]), .Z(n14807) );
  AND U12941 ( .A(n5556), .B(n14807), .Z(n5557) );
  NANDN U12942 ( .A(n14810), .B(n5557), .Z(n5558) );
  NANDN U12943 ( .A(x[371]), .B(y[371]), .Z(n14808) );
  AND U12944 ( .A(n5558), .B(n14808), .Z(n5559) );
  NAND U12945 ( .A(n14805), .B(n5559), .Z(n5560) );
  NANDN U12946 ( .A(n14806), .B(n5560), .Z(n5561) );
  NANDN U12947 ( .A(y[373]), .B(x[373]), .Z(n14803) );
  NANDN U12948 ( .A(n5561), .B(n14803), .Z(n5562) );
  AND U12949 ( .A(n5563), .B(n5562), .Z(n5565) );
  NANDN U12950 ( .A(y[375]), .B(x[375]), .Z(n14799) );
  ANDN U12951 ( .B(x[374]), .A(y[374]), .Z(n14802) );
  ANDN U12952 ( .B(n14799), .A(n14802), .Z(n5564) );
  NANDN U12953 ( .A(n5565), .B(n5564), .Z(n5566) );
  AND U12954 ( .A(n14801), .B(n5566), .Z(n5567) );
  NANDN U12955 ( .A(x[376]), .B(y[376]), .Z(n14796) );
  NAND U12956 ( .A(n5567), .B(n14796), .Z(n5568) );
  ANDN U12957 ( .B(x[377]), .A(y[377]), .Z(n14794) );
  ANDN U12958 ( .B(n5568), .A(n14794), .Z(n5569) );
  NAND U12959 ( .A(n14798), .B(n5569), .Z(n5570) );
  NANDN U12960 ( .A(x[377]), .B(y[377]), .Z(n14797) );
  AND U12961 ( .A(n5570), .B(n14797), .Z(n5571) );
  NAND U12962 ( .A(n14792), .B(n5571), .Z(n5572) );
  NAND U12963 ( .A(n14795), .B(n5572), .Z(n5573) );
  ANDN U12964 ( .B(x[379]), .A(y[379]), .Z(n14790) );
  OR U12965 ( .A(n5573), .B(n14790), .Z(n5574) );
  AND U12966 ( .A(n5575), .B(n5574), .Z(n5577) );
  NANDN U12967 ( .A(y[381]), .B(x[381]), .Z(n14787) );
  NANDN U12968 ( .A(y[380]), .B(x[380]), .Z(n14791) );
  AND U12969 ( .A(n14787), .B(n14791), .Z(n5576) );
  NANDN U12970 ( .A(n5577), .B(n5576), .Z(n5578) );
  AND U12971 ( .A(n14789), .B(n5578), .Z(n5579) );
  NANDN U12972 ( .A(x[382]), .B(y[382]), .Z(n14785) );
  NAND U12973 ( .A(n5579), .B(n14785), .Z(n5580) );
  ANDN U12974 ( .B(x[383]), .A(y[383]), .Z(n14782) );
  ANDN U12975 ( .B(n5580), .A(n14782), .Z(n5581) );
  NANDN U12976 ( .A(n14786), .B(n5581), .Z(n5582) );
  NANDN U12977 ( .A(x[383]), .B(y[383]), .Z(n14784) );
  AND U12978 ( .A(n5582), .B(n14784), .Z(n5583) );
  NAND U12979 ( .A(n14780), .B(n5583), .Z(n5584) );
  NAND U12980 ( .A(n14783), .B(n5584), .Z(n5585) );
  ANDN U12981 ( .B(x[385]), .A(y[385]), .Z(n14778) );
  OR U12982 ( .A(n5585), .B(n14778), .Z(n5586) );
  AND U12983 ( .A(n5587), .B(n5586), .Z(n5589) );
  NANDN U12984 ( .A(y[386]), .B(x[386]), .Z(n14779) );
  ANDN U12985 ( .B(x[387]), .A(y[387]), .Z(n14774) );
  ANDN U12986 ( .B(n14779), .A(n14774), .Z(n5588) );
  NANDN U12987 ( .A(n5589), .B(n5588), .Z(n5590) );
  AND U12988 ( .A(n14776), .B(n5590), .Z(n5591) );
  NANDN U12989 ( .A(x[388]), .B(y[388]), .Z(n14772) );
  NAND U12990 ( .A(n5591), .B(n14772), .Z(n5592) );
  ANDN U12991 ( .B(x[389]), .A(y[389]), .Z(n14770) );
  ANDN U12992 ( .B(n5592), .A(n14770), .Z(n5593) );
  NAND U12993 ( .A(n14775), .B(n5593), .Z(n5594) );
  AND U12994 ( .A(n14773), .B(n5594), .Z(n5595) );
  NAND U12995 ( .A(n5596), .B(n5595), .Z(n5597) );
  NAND U12996 ( .A(n14771), .B(n5597), .Z(n5598) );
  AND U12997 ( .A(n14769), .B(n5598), .Z(n5601) );
  NANDN U12998 ( .A(y[391]), .B(x[391]), .Z(n5600) );
  NANDN U12999 ( .A(y[392]), .B(x[392]), .Z(n5599) );
  NAND U13000 ( .A(n5600), .B(n5599), .Z(n25301) );
  OR U13001 ( .A(n5601), .B(n25301), .Z(n5602) );
  NAND U13002 ( .A(n25303), .B(n5602), .Z(n5603) );
  NANDN U13003 ( .A(n25305), .B(n5603), .Z(n5604) );
  NAND U13004 ( .A(n25307), .B(n5604), .Z(n5605) );
  NANDN U13005 ( .A(n25309), .B(n5605), .Z(n5606) );
  AND U13006 ( .A(n25311), .B(n5606), .Z(n5607) );
  OR U13007 ( .A(n25313), .B(n5607), .Z(n5608) );
  NAND U13008 ( .A(n25315), .B(n5608), .Z(n5609) );
  NANDN U13009 ( .A(n25317), .B(n5609), .Z(n5610) );
  NAND U13010 ( .A(n25319), .B(n5610), .Z(n5611) );
  NANDN U13011 ( .A(n14767), .B(n5611), .Z(n5612) );
  AND U13012 ( .A(n14765), .B(n5612), .Z(n5615) );
  NANDN U13013 ( .A(y[403]), .B(x[403]), .Z(n14763) );
  ANDN U13014 ( .B(x[402]), .A(y[402]), .Z(n5613) );
  ANDN U13015 ( .B(n14763), .A(n5613), .Z(n5614) );
  NANDN U13016 ( .A(n5615), .B(n5614), .Z(n5616) );
  AND U13017 ( .A(n14764), .B(n5616), .Z(n5617) );
  NANDN U13018 ( .A(x[404]), .B(y[404]), .Z(n14761) );
  NAND U13019 ( .A(n5617), .B(n14761), .Z(n5618) );
  NANDN U13020 ( .A(y[405]), .B(x[405]), .Z(n14759) );
  AND U13021 ( .A(n5618), .B(n14759), .Z(n5619) );
  NANDN U13022 ( .A(n14762), .B(n5619), .Z(n5620) );
  NANDN U13023 ( .A(x[405]), .B(y[405]), .Z(n14760) );
  AND U13024 ( .A(n5620), .B(n14760), .Z(n5621) );
  NAND U13025 ( .A(n14757), .B(n5621), .Z(n5622) );
  NANDN U13026 ( .A(n14758), .B(n5622), .Z(n5623) );
  ANDN U13027 ( .B(x[407]), .A(y[407]), .Z(n14754) );
  OR U13028 ( .A(n5623), .B(n14754), .Z(n5624) );
  AND U13029 ( .A(n5625), .B(n5624), .Z(n5627) );
  NANDN U13030 ( .A(y[408]), .B(x[408]), .Z(n14755) );
  ANDN U13031 ( .B(x[409]), .A(y[409]), .Z(n14751) );
  ANDN U13032 ( .B(n14755), .A(n14751), .Z(n5626) );
  NANDN U13033 ( .A(n5627), .B(n5626), .Z(n5628) );
  AND U13034 ( .A(n14753), .B(n5628), .Z(n5629) );
  NANDN U13035 ( .A(x[410]), .B(y[410]), .Z(n14749) );
  NAND U13036 ( .A(n5629), .B(n14749), .Z(n5630) );
  NANDN U13037 ( .A(y[411]), .B(x[411]), .Z(n14747) );
  AND U13038 ( .A(n5630), .B(n14747), .Z(n5631) );
  NANDN U13039 ( .A(n5632), .B(n5631), .Z(n5633) );
  NANDN U13040 ( .A(x[411]), .B(y[411]), .Z(n14748) );
  AND U13041 ( .A(n5633), .B(n14748), .Z(n5634) );
  NAND U13042 ( .A(n14745), .B(n5634), .Z(n5635) );
  NANDN U13043 ( .A(n14746), .B(n5635), .Z(n5636) );
  NANDN U13044 ( .A(y[413]), .B(x[413]), .Z(n14743) );
  NANDN U13045 ( .A(n5636), .B(n14743), .Z(n5637) );
  AND U13046 ( .A(n5638), .B(n5637), .Z(n5640) );
  ANDN U13047 ( .B(x[414]), .A(y[414]), .Z(n14742) );
  ANDN U13048 ( .B(x[415]), .A(y[415]), .Z(n14739) );
  NOR U13049 ( .A(n14742), .B(n14739), .Z(n5639) );
  NANDN U13050 ( .A(n5640), .B(n5639), .Z(n5641) );
  AND U13051 ( .A(n14740), .B(n5641), .Z(n5642) );
  NANDN U13052 ( .A(x[416]), .B(y[416]), .Z(n14737) );
  NAND U13053 ( .A(n5642), .B(n14737), .Z(n5643) );
  ANDN U13054 ( .B(x[417]), .A(y[417]), .Z(n14734) );
  ANDN U13055 ( .B(n5643), .A(n14734), .Z(n5644) );
  NANDN U13056 ( .A(n5645), .B(n5644), .Z(n5646) );
  AND U13057 ( .A(n14736), .B(n5646), .Z(n5647) );
  NAND U13058 ( .A(n5648), .B(n5647), .Z(n5649) );
  NAND U13059 ( .A(n14735), .B(n5649), .Z(n5650) );
  AND U13060 ( .A(n14733), .B(n5650), .Z(n5653) );
  NANDN U13061 ( .A(y[419]), .B(x[419]), .Z(n5652) );
  NANDN U13062 ( .A(y[420]), .B(x[420]), .Z(n5651) );
  NAND U13063 ( .A(n5652), .B(n5651), .Z(n25357) );
  OR U13064 ( .A(n5653), .B(n25357), .Z(n5654) );
  NAND U13065 ( .A(n25359), .B(n5654), .Z(n5655) );
  NANDN U13066 ( .A(n14730), .B(n5655), .Z(n5656) );
  NANDN U13067 ( .A(x[422]), .B(y[422]), .Z(n14728) );
  NAND U13068 ( .A(n5656), .B(n14728), .Z(n5657) );
  ANDN U13069 ( .B(x[423]), .A(y[423]), .Z(n14726) );
  ANDN U13070 ( .B(n5657), .A(n14726), .Z(n5658) );
  NAND U13071 ( .A(n14731), .B(n5658), .Z(n5659) );
  NANDN U13072 ( .A(x[423]), .B(y[423]), .Z(n14729) );
  AND U13073 ( .A(n5659), .B(n14729), .Z(n5660) );
  NAND U13074 ( .A(n14725), .B(n5660), .Z(n5661) );
  NAND U13075 ( .A(n14727), .B(n5661), .Z(n5662) );
  ANDN U13076 ( .B(x[425]), .A(y[425]), .Z(n14723) );
  OR U13077 ( .A(n5662), .B(n14723), .Z(n5663) );
  AND U13078 ( .A(n5664), .B(n5663), .Z(n5667) );
  ANDN U13079 ( .B(x[427]), .A(y[427]), .Z(n14719) );
  ANDN U13080 ( .B(x[426]), .A(y[426]), .Z(n5665) );
  NOR U13081 ( .A(n14719), .B(n5665), .Z(n5666) );
  NANDN U13082 ( .A(n5667), .B(n5666), .Z(n5668) );
  AND U13083 ( .A(n14720), .B(n5668), .Z(n5669) );
  NANDN U13084 ( .A(x[428]), .B(y[428]), .Z(n14717) );
  NAND U13085 ( .A(n5669), .B(n14717), .Z(n5670) );
  NANDN U13086 ( .A(n5671), .B(n5670), .Z(n5672) );
  AND U13087 ( .A(n14716), .B(n5672), .Z(n5675) );
  NANDN U13088 ( .A(y[429]), .B(x[429]), .Z(n5674) );
  NANDN U13089 ( .A(y[430]), .B(x[430]), .Z(n5673) );
  NAND U13090 ( .A(n5674), .B(n5673), .Z(n25377) );
  OR U13091 ( .A(n5675), .B(n25377), .Z(n5676) );
  NAND U13092 ( .A(n25379), .B(n5676), .Z(n5677) );
  NANDN U13093 ( .A(n25381), .B(n5677), .Z(n5678) );
  NANDN U13094 ( .A(x[432]), .B(y[432]), .Z(n14715) );
  NAND U13095 ( .A(n5678), .B(n14715), .Z(n5679) );
  NANDN U13096 ( .A(n14713), .B(n5679), .Z(n5680) );
  AND U13097 ( .A(n14714), .B(n5680), .Z(n5681) );
  NANDN U13098 ( .A(x[434]), .B(y[434]), .Z(n14711) );
  NAND U13099 ( .A(n5681), .B(n14711), .Z(n5682) );
  NANDN U13100 ( .A(y[435]), .B(x[435]), .Z(n14709) );
  AND U13101 ( .A(n5682), .B(n14709), .Z(n5683) );
  NANDN U13102 ( .A(n5684), .B(n5683), .Z(n5685) );
  NANDN U13103 ( .A(x[435]), .B(y[435]), .Z(n14710) );
  AND U13104 ( .A(n5685), .B(n14710), .Z(n5686) );
  NAND U13105 ( .A(n14707), .B(n5686), .Z(n5687) );
  NANDN U13106 ( .A(n14708), .B(n5687), .Z(n5688) );
  ANDN U13107 ( .B(x[437]), .A(y[437]), .Z(n14705) );
  OR U13108 ( .A(n5688), .B(n14705), .Z(n5689) );
  AND U13109 ( .A(n5690), .B(n5689), .Z(n5693) );
  NANDN U13110 ( .A(y[439]), .B(x[439]), .Z(n14701) );
  ANDN U13111 ( .B(x[438]), .A(y[438]), .Z(n5691) );
  ANDN U13112 ( .B(n14701), .A(n5691), .Z(n5692) );
  NANDN U13113 ( .A(n5693), .B(n5692), .Z(n5694) );
  AND U13114 ( .A(n14702), .B(n5694), .Z(n5695) );
  NANDN U13115 ( .A(x[440]), .B(y[440]), .Z(n14698) );
  NAND U13116 ( .A(n5695), .B(n14698), .Z(n5696) );
  NANDN U13117 ( .A(y[441]), .B(x[441]), .Z(n14697) );
  AND U13118 ( .A(n5696), .B(n14697), .Z(n5697) );
  NANDN U13119 ( .A(n14700), .B(n5697), .Z(n5698) );
  NANDN U13120 ( .A(x[441]), .B(y[441]), .Z(n14699) );
  NAND U13121 ( .A(n5698), .B(n14699), .Z(n5699) );
  NANDN U13122 ( .A(n14696), .B(n5699), .Z(n5700) );
  AND U13123 ( .A(n14695), .B(n5700), .Z(n5701) );
  NANDN U13124 ( .A(y[443]), .B(x[443]), .Z(n14693) );
  NANDN U13125 ( .A(n5701), .B(n14693), .Z(n5702) );
  AND U13126 ( .A(n5703), .B(n5702), .Z(n5705) );
  NANDN U13127 ( .A(y[445]), .B(x[445]), .Z(n14689) );
  ANDN U13128 ( .B(x[444]), .A(y[444]), .Z(n14692) );
  ANDN U13129 ( .B(n14689), .A(n14692), .Z(n5704) );
  NANDN U13130 ( .A(n5705), .B(n5704), .Z(n5706) );
  AND U13131 ( .A(n14690), .B(n5706), .Z(n5707) );
  NANDN U13132 ( .A(x[446]), .B(y[446]), .Z(n14686) );
  NAND U13133 ( .A(n5707), .B(n14686), .Z(n5708) );
  ANDN U13134 ( .B(x[447]), .A(y[447]), .Z(n14684) );
  ANDN U13135 ( .B(n5708), .A(n14684), .Z(n5709) );
  NANDN U13136 ( .A(n14688), .B(n5709), .Z(n5710) );
  NANDN U13137 ( .A(x[447]), .B(y[447]), .Z(n14687) );
  AND U13138 ( .A(n5710), .B(n14687), .Z(n5711) );
  NAND U13139 ( .A(n14682), .B(n5711), .Z(n5712) );
  NAND U13140 ( .A(n14685), .B(n5712), .Z(n5713) );
  ANDN U13141 ( .B(x[449]), .A(y[449]), .Z(n14681) );
  OR U13142 ( .A(n5713), .B(n14681), .Z(n5714) );
  AND U13143 ( .A(n5715), .B(n5714), .Z(n5718) );
  ANDN U13144 ( .B(x[451]), .A(y[451]), .Z(n14676) );
  ANDN U13145 ( .B(x[450]), .A(y[450]), .Z(n5716) );
  NOR U13146 ( .A(n14676), .B(n5716), .Z(n5717) );
  NANDN U13147 ( .A(n5718), .B(n5717), .Z(n5719) );
  AND U13148 ( .A(n14678), .B(n5719), .Z(n5720) );
  NANDN U13149 ( .A(x[452]), .B(y[452]), .Z(n14674) );
  NAND U13150 ( .A(n5720), .B(n14674), .Z(n5721) );
  ANDN U13151 ( .B(x[453]), .A(y[453]), .Z(n14672) );
  ANDN U13152 ( .B(n5721), .A(n14672), .Z(n5722) );
  NAND U13153 ( .A(n14677), .B(n5722), .Z(n5723) );
  NANDN U13154 ( .A(x[453]), .B(y[453]), .Z(n14675) );
  AND U13155 ( .A(n5723), .B(n14675), .Z(n5724) );
  NAND U13156 ( .A(n14670), .B(n5724), .Z(n5725) );
  NAND U13157 ( .A(n14673), .B(n5725), .Z(n5726) );
  ANDN U13158 ( .B(x[455]), .A(y[455]), .Z(n14669) );
  OR U13159 ( .A(n5726), .B(n14669), .Z(n5727) );
  AND U13160 ( .A(n5728), .B(n5727), .Z(n5731) );
  ANDN U13161 ( .B(x[457]), .A(y[457]), .Z(n14664) );
  ANDN U13162 ( .B(x[456]), .A(y[456]), .Z(n5729) );
  NOR U13163 ( .A(n14664), .B(n5729), .Z(n5730) );
  NANDN U13164 ( .A(n5731), .B(n5730), .Z(n5732) );
  AND U13165 ( .A(n14666), .B(n5732), .Z(n5733) );
  NANDN U13166 ( .A(x[458]), .B(y[458]), .Z(n14662) );
  NAND U13167 ( .A(n5733), .B(n14662), .Z(n5734) );
  NANDN U13168 ( .A(y[459]), .B(x[459]), .Z(n14661) );
  AND U13169 ( .A(n5734), .B(n14661), .Z(n5735) );
  NAND U13170 ( .A(n14665), .B(n5735), .Z(n5736) );
  NANDN U13171 ( .A(x[459]), .B(y[459]), .Z(n14663) );
  AND U13172 ( .A(n5736), .B(n14663), .Z(n5737) );
  NAND U13173 ( .A(n14659), .B(n5737), .Z(n5738) );
  NANDN U13174 ( .A(n14660), .B(n5738), .Z(n5739) );
  ANDN U13175 ( .B(x[461]), .A(y[461]), .Z(n14656) );
  OR U13176 ( .A(n5739), .B(n14656), .Z(n5740) );
  AND U13177 ( .A(n5741), .B(n5740), .Z(n5743) );
  NANDN U13178 ( .A(y[462]), .B(x[462]), .Z(n14657) );
  ANDN U13179 ( .B(x[463]), .A(y[463]), .Z(n14653) );
  ANDN U13180 ( .B(n14657), .A(n14653), .Z(n5742) );
  NANDN U13181 ( .A(n5743), .B(n5742), .Z(n5744) );
  AND U13182 ( .A(n14654), .B(n5744), .Z(n5745) );
  NANDN U13183 ( .A(x[464]), .B(y[464]), .Z(n14651) );
  NAND U13184 ( .A(n5745), .B(n14651), .Z(n5746) );
  ANDN U13185 ( .B(x[465]), .A(y[465]), .Z(n14648) );
  ANDN U13186 ( .B(n5746), .A(n14648), .Z(n5747) );
  NANDN U13187 ( .A(n5748), .B(n5747), .Z(n5749) );
  NANDN U13188 ( .A(x[465]), .B(y[465]), .Z(n14650) );
  AND U13189 ( .A(n5749), .B(n14650), .Z(n5750) );
  NAND U13190 ( .A(n14646), .B(n5750), .Z(n5751) );
  NAND U13191 ( .A(n14649), .B(n5751), .Z(n5752) );
  ANDN U13192 ( .B(x[467]), .A(y[467]), .Z(n14644) );
  OR U13193 ( .A(n5752), .B(n14644), .Z(n5753) );
  AND U13194 ( .A(n5754), .B(n5753), .Z(n5756) );
  NANDN U13195 ( .A(y[469]), .B(x[469]), .Z(n14641) );
  NANDN U13196 ( .A(y[468]), .B(x[468]), .Z(n14645) );
  AND U13197 ( .A(n14641), .B(n14645), .Z(n5755) );
  NANDN U13198 ( .A(n5756), .B(n5755), .Z(n5757) );
  AND U13199 ( .A(n14642), .B(n5757), .Z(n5758) );
  NANDN U13200 ( .A(x[470]), .B(y[470]), .Z(n14639) );
  NAND U13201 ( .A(n5758), .B(n14639), .Z(n5759) );
  NANDN U13202 ( .A(y[471]), .B(x[471]), .Z(n14637) );
  AND U13203 ( .A(n5759), .B(n14637), .Z(n5760) );
  NANDN U13204 ( .A(n14640), .B(n5760), .Z(n5761) );
  NANDN U13205 ( .A(x[471]), .B(y[471]), .Z(n14638) );
  AND U13206 ( .A(n5761), .B(n14638), .Z(n5762) );
  NAND U13207 ( .A(n14635), .B(n5762), .Z(n5763) );
  NANDN U13208 ( .A(n14636), .B(n5763), .Z(n5764) );
  ANDN U13209 ( .B(x[473]), .A(y[473]), .Z(n14632) );
  OR U13210 ( .A(n5764), .B(n14632), .Z(n5765) );
  AND U13211 ( .A(n5766), .B(n5765), .Z(n5768) );
  NANDN U13212 ( .A(y[474]), .B(x[474]), .Z(n14633) );
  ANDN U13213 ( .B(x[475]), .A(y[475]), .Z(n14628) );
  ANDN U13214 ( .B(n14633), .A(n14628), .Z(n5767) );
  NANDN U13215 ( .A(n5768), .B(n5767), .Z(n5769) );
  AND U13216 ( .A(n14631), .B(n5769), .Z(n5770) );
  NANDN U13217 ( .A(x[476]), .B(y[476]), .Z(n14626) );
  NAND U13218 ( .A(n5770), .B(n14626), .Z(n5771) );
  NANDN U13219 ( .A(y[477]), .B(x[477]), .Z(n14625) );
  AND U13220 ( .A(n5771), .B(n14625), .Z(n5772) );
  NAND U13221 ( .A(n14629), .B(n5772), .Z(n5773) );
  NANDN U13222 ( .A(x[477]), .B(y[477]), .Z(n14627) );
  AND U13223 ( .A(n5773), .B(n14627), .Z(n5774) );
  NAND U13224 ( .A(n14622), .B(n5774), .Z(n5775) );
  NANDN U13225 ( .A(n14624), .B(n5775), .Z(n5776) );
  ANDN U13226 ( .B(x[479]), .A(y[479]), .Z(n14620) );
  OR U13227 ( .A(n5776), .B(n14620), .Z(n5777) );
  AND U13228 ( .A(n5778), .B(n5777), .Z(n5780) );
  NANDN U13229 ( .A(y[481]), .B(x[481]), .Z(n14617) );
  NANDN U13230 ( .A(y[480]), .B(x[480]), .Z(n14621) );
  AND U13231 ( .A(n14617), .B(n14621), .Z(n5779) );
  NANDN U13232 ( .A(n5780), .B(n5779), .Z(n5781) );
  AND U13233 ( .A(n14619), .B(n5781), .Z(n5782) );
  NANDN U13234 ( .A(x[482]), .B(y[482]), .Z(n14615) );
  NAND U13235 ( .A(n5782), .B(n14615), .Z(n5783) );
  NANDN U13236 ( .A(y[483]), .B(x[483]), .Z(n14613) );
  AND U13237 ( .A(n5783), .B(n14613), .Z(n5784) );
  NANDN U13238 ( .A(n14616), .B(n5784), .Z(n5785) );
  NANDN U13239 ( .A(x[483]), .B(y[483]), .Z(n14614) );
  AND U13240 ( .A(n5785), .B(n14614), .Z(n5786) );
  NAND U13241 ( .A(n14611), .B(n5786), .Z(n5787) );
  NANDN U13242 ( .A(n14612), .B(n5787), .Z(n5788) );
  ANDN U13243 ( .B(x[485]), .A(y[485]), .Z(n14609) );
  OR U13244 ( .A(n5788), .B(n14609), .Z(n5789) );
  AND U13245 ( .A(n5790), .B(n5789), .Z(n5793) );
  ANDN U13246 ( .B(x[487]), .A(y[487]), .Z(n14604) );
  ANDN U13247 ( .B(x[486]), .A(y[486]), .Z(n5791) );
  NOR U13248 ( .A(n14604), .B(n5791), .Z(n5792) );
  NANDN U13249 ( .A(n5793), .B(n5792), .Z(n5794) );
  AND U13250 ( .A(n14606), .B(n5794), .Z(n5795) );
  NANDN U13251 ( .A(x[488]), .B(y[488]), .Z(n14603) );
  NAND U13252 ( .A(n5795), .B(n14603), .Z(n5796) );
  ANDN U13253 ( .B(x[489]), .A(y[489]), .Z(n14599) );
  ANDN U13254 ( .B(n5796), .A(n14599), .Z(n5797) );
  NAND U13255 ( .A(n14605), .B(n5797), .Z(n5798) );
  NANDN U13256 ( .A(x[489]), .B(y[489]), .Z(n14602) );
  AND U13257 ( .A(n5798), .B(n14602), .Z(n5799) );
  NAND U13258 ( .A(n14598), .B(n5799), .Z(n5800) );
  NAND U13259 ( .A(n14600), .B(n5800), .Z(n5801) );
  ANDN U13260 ( .B(x[491]), .A(y[491]), .Z(n14595) );
  OR U13261 ( .A(n5801), .B(n14595), .Z(n5802) );
  AND U13262 ( .A(n5803), .B(n5802), .Z(n5805) );
  NANDN U13263 ( .A(y[492]), .B(x[492]), .Z(n14596) );
  ANDN U13264 ( .B(x[493]), .A(y[493]), .Z(n14591) );
  ANDN U13265 ( .B(n14596), .A(n14591), .Z(n5804) );
  NANDN U13266 ( .A(n5805), .B(n5804), .Z(n5806) );
  AND U13267 ( .A(n14594), .B(n5806), .Z(n5807) );
  NANDN U13268 ( .A(x[494]), .B(y[494]), .Z(n14590) );
  NAND U13269 ( .A(n5807), .B(n14590), .Z(n5808) );
  NANDN U13270 ( .A(y[495]), .B(x[495]), .Z(n14588) );
  AND U13271 ( .A(n5808), .B(n14588), .Z(n5809) );
  NAND U13272 ( .A(n14592), .B(n5809), .Z(n5810) );
  NANDN U13273 ( .A(x[495]), .B(y[495]), .Z(n14589) );
  AND U13274 ( .A(n5810), .B(n14589), .Z(n5811) );
  NAND U13275 ( .A(n14586), .B(n5811), .Z(n5812) );
  NANDN U13276 ( .A(n14587), .B(n5812), .Z(n5813) );
  ANDN U13277 ( .B(x[497]), .A(y[497]), .Z(n14583) );
  OR U13278 ( .A(n5813), .B(n14583), .Z(n5814) );
  AND U13279 ( .A(n5815), .B(n5814), .Z(n5817) );
  NANDN U13280 ( .A(y[499]), .B(x[499]), .Z(n14580) );
  NANDN U13281 ( .A(y[498]), .B(x[498]), .Z(n14584) );
  AND U13282 ( .A(n14580), .B(n14584), .Z(n5816) );
  NANDN U13283 ( .A(n5817), .B(n5816), .Z(n5818) );
  AND U13284 ( .A(n14581), .B(n5818), .Z(n5819) );
  NANDN U13285 ( .A(x[500]), .B(y[500]), .Z(n14578) );
  NAND U13286 ( .A(n5819), .B(n14578), .Z(n5820) );
  ANDN U13287 ( .B(x[501]), .A(y[501]), .Z(n14575) );
  ANDN U13288 ( .B(n5820), .A(n14575), .Z(n5821) );
  NANDN U13289 ( .A(n14579), .B(n5821), .Z(n5822) );
  NANDN U13290 ( .A(x[501]), .B(y[501]), .Z(n14577) );
  AND U13291 ( .A(n5822), .B(n14577), .Z(n5823) );
  NAND U13292 ( .A(n14573), .B(n5823), .Z(n5824) );
  NAND U13293 ( .A(n14576), .B(n5824), .Z(n5825) );
  ANDN U13294 ( .B(x[503]), .A(y[503]), .Z(n14571) );
  OR U13295 ( .A(n5825), .B(n14571), .Z(n5826) );
  AND U13296 ( .A(n5827), .B(n5826), .Z(n5829) );
  NANDN U13297 ( .A(y[505]), .B(x[505]), .Z(n14568) );
  NANDN U13298 ( .A(y[504]), .B(x[504]), .Z(n14572) );
  AND U13299 ( .A(n14568), .B(n14572), .Z(n5828) );
  NANDN U13300 ( .A(n5829), .B(n5828), .Z(n5830) );
  AND U13301 ( .A(n14569), .B(n5830), .Z(n5831) );
  NANDN U13302 ( .A(x[506]), .B(y[506]), .Z(n14566) );
  NAND U13303 ( .A(n5831), .B(n14566), .Z(n5832) );
  ANDN U13304 ( .B(x[507]), .A(y[507]), .Z(n25532) );
  ANDN U13305 ( .B(n5832), .A(n25532), .Z(n5833) );
  NANDN U13306 ( .A(n14567), .B(n5833), .Z(n5834) );
  XNOR U13307 ( .A(x[508]), .B(y[508]), .Z(n24539) );
  AND U13308 ( .A(n5834), .B(n24539), .Z(n5835) );
  NAND U13309 ( .A(n14565), .B(n5835), .Z(n5836) );
  NANDN U13310 ( .A(n16012), .B(n5836), .Z(n5837) );
  ANDN U13311 ( .B(x[509]), .A(y[509]), .Z(n14562) );
  OR U13312 ( .A(n5837), .B(n14562), .Z(n5838) );
  AND U13313 ( .A(n5839), .B(n5838), .Z(n5842) );
  ANDN U13314 ( .B(x[511]), .A(y[511]), .Z(n14557) );
  ANDN U13315 ( .B(x[510]), .A(y[510]), .Z(n5840) );
  NOR U13316 ( .A(n14557), .B(n5840), .Z(n5841) );
  NANDN U13317 ( .A(n5842), .B(n5841), .Z(n5843) );
  AND U13318 ( .A(n14559), .B(n5843), .Z(n5844) );
  NANDN U13319 ( .A(x[512]), .B(y[512]), .Z(n14556) );
  NAND U13320 ( .A(n5844), .B(n14556), .Z(n5845) );
  ANDN U13321 ( .B(x[513]), .A(y[513]), .Z(n14553) );
  ANDN U13322 ( .B(n5845), .A(n14553), .Z(n5846) );
  NAND U13323 ( .A(n14558), .B(n5846), .Z(n5847) );
  NANDN U13324 ( .A(x[513]), .B(y[513]), .Z(n14555) );
  AND U13325 ( .A(n5847), .B(n14555), .Z(n5848) );
  NAND U13326 ( .A(n14551), .B(n5848), .Z(n5849) );
  NAND U13327 ( .A(n14554), .B(n5849), .Z(n5850) );
  ANDN U13328 ( .B(x[515]), .A(y[515]), .Z(n14549) );
  OR U13329 ( .A(n5850), .B(n14549), .Z(n5851) );
  AND U13330 ( .A(n5852), .B(n5851), .Z(n5854) );
  NANDN U13331 ( .A(y[516]), .B(x[516]), .Z(n14550) );
  ANDN U13332 ( .B(x[517]), .A(y[517]), .Z(n14546) );
  ANDN U13333 ( .B(n14550), .A(n14546), .Z(n5853) );
  NANDN U13334 ( .A(n5854), .B(n5853), .Z(n5855) );
  AND U13335 ( .A(n14547), .B(n5855), .Z(n5856) );
  NANDN U13336 ( .A(x[518]), .B(y[518]), .Z(n14544) );
  NAND U13337 ( .A(n5856), .B(n14544), .Z(n5857) );
  ANDN U13338 ( .B(x[519]), .A(y[519]), .Z(n14541) );
  ANDN U13339 ( .B(n5857), .A(n14541), .Z(n5858) );
  NANDN U13340 ( .A(n5859), .B(n5858), .Z(n5860) );
  NANDN U13341 ( .A(x[519]), .B(y[519]), .Z(n14543) );
  AND U13342 ( .A(n5860), .B(n14543), .Z(n5861) );
  NAND U13343 ( .A(n14539), .B(n5861), .Z(n5862) );
  NAND U13344 ( .A(n14542), .B(n5862), .Z(n5863) );
  ANDN U13345 ( .B(x[521]), .A(y[521]), .Z(n14538) );
  OR U13346 ( .A(n5863), .B(n14538), .Z(n5864) );
  AND U13347 ( .A(n5865), .B(n5864), .Z(n5868) );
  NANDN U13348 ( .A(y[523]), .B(x[523]), .Z(n14534) );
  ANDN U13349 ( .B(x[522]), .A(y[522]), .Z(n5866) );
  ANDN U13350 ( .B(n14534), .A(n5866), .Z(n5867) );
  NANDN U13351 ( .A(n5868), .B(n5867), .Z(n5869) );
  AND U13352 ( .A(n14535), .B(n5869), .Z(n5870) );
  NANDN U13353 ( .A(x[524]), .B(y[524]), .Z(n14531) );
  NAND U13354 ( .A(n5870), .B(n14531), .Z(n5871) );
  ANDN U13355 ( .B(x[525]), .A(y[525]), .Z(n14529) );
  ANDN U13356 ( .B(n5871), .A(n14529), .Z(n5872) );
  NANDN U13357 ( .A(n14533), .B(n5872), .Z(n5873) );
  NANDN U13358 ( .A(x[525]), .B(y[525]), .Z(n14532) );
  AND U13359 ( .A(n5873), .B(n14532), .Z(n5874) );
  NAND U13360 ( .A(n14528), .B(n5874), .Z(n5875) );
  NAND U13361 ( .A(n14530), .B(n5875), .Z(n5876) );
  ANDN U13362 ( .B(x[527]), .A(y[527]), .Z(n14526) );
  OR U13363 ( .A(n5876), .B(n14526), .Z(n5877) );
  AND U13364 ( .A(n5878), .B(n5877), .Z(n5881) );
  NANDN U13365 ( .A(y[529]), .B(x[529]), .Z(n14522) );
  ANDN U13366 ( .B(x[528]), .A(y[528]), .Z(n5879) );
  ANDN U13367 ( .B(n14522), .A(n5879), .Z(n5880) );
  NANDN U13368 ( .A(n5881), .B(n5880), .Z(n5882) );
  AND U13369 ( .A(n14523), .B(n5882), .Z(n5883) );
  NANDN U13370 ( .A(x[530]), .B(y[530]), .Z(n14520) );
  NAND U13371 ( .A(n5883), .B(n14520), .Z(n5884) );
  ANDN U13372 ( .B(x[531]), .A(y[531]), .Z(n14517) );
  ANDN U13373 ( .B(n5884), .A(n14517), .Z(n5885) );
  NANDN U13374 ( .A(n14521), .B(n5885), .Z(n5886) );
  NANDN U13375 ( .A(x[531]), .B(y[531]), .Z(n14519) );
  AND U13376 ( .A(n5886), .B(n14519), .Z(n5887) );
  NAND U13377 ( .A(n14516), .B(n5887), .Z(n5888) );
  NAND U13378 ( .A(n14518), .B(n5888), .Z(n5889) );
  ANDN U13379 ( .B(x[533]), .A(y[533]), .Z(n14513) );
  OR U13380 ( .A(n5889), .B(n14513), .Z(n5890) );
  AND U13381 ( .A(n5891), .B(n5890), .Z(n5894) );
  ANDN U13382 ( .B(x[535]), .A(y[535]), .Z(n14509) );
  ANDN U13383 ( .B(x[534]), .A(y[534]), .Z(n5892) );
  NOR U13384 ( .A(n14509), .B(n5892), .Z(n5893) );
  NANDN U13385 ( .A(n5894), .B(n5893), .Z(n5895) );
  AND U13386 ( .A(n14511), .B(n5895), .Z(n5896) );
  NANDN U13387 ( .A(x[536]), .B(y[536]), .Z(n14507) );
  NAND U13388 ( .A(n5896), .B(n14507), .Z(n5897) );
  NANDN U13389 ( .A(y[537]), .B(x[537]), .Z(n14506) );
  AND U13390 ( .A(n5897), .B(n14506), .Z(n5898) );
  NAND U13391 ( .A(n14510), .B(n5898), .Z(n5899) );
  NANDN U13392 ( .A(x[537]), .B(y[537]), .Z(n14508) );
  AND U13393 ( .A(n5899), .B(n14508), .Z(n5900) );
  NAND U13394 ( .A(n14504), .B(n5900), .Z(n5901) );
  NANDN U13395 ( .A(n14505), .B(n5901), .Z(n5902) );
  ANDN U13396 ( .B(x[539]), .A(y[539]), .Z(n14501) );
  OR U13397 ( .A(n5902), .B(n14501), .Z(n5903) );
  AND U13398 ( .A(n5904), .B(n5903), .Z(n5906) );
  NANDN U13399 ( .A(y[540]), .B(x[540]), .Z(n14502) );
  ANDN U13400 ( .B(x[541]), .A(y[541]), .Z(n14498) );
  ANDN U13401 ( .B(n14502), .A(n14498), .Z(n5905) );
  NANDN U13402 ( .A(n5906), .B(n5905), .Z(n5907) );
  AND U13403 ( .A(n14499), .B(n5907), .Z(n5908) );
  NANDN U13404 ( .A(x[542]), .B(y[542]), .Z(n14496) );
  NAND U13405 ( .A(n5908), .B(n14496), .Z(n5909) );
  NANDN U13406 ( .A(y[543]), .B(x[543]), .Z(n14494) );
  AND U13407 ( .A(n5909), .B(n14494), .Z(n5910) );
  NANDN U13408 ( .A(n5911), .B(n5910), .Z(n5912) );
  NANDN U13409 ( .A(x[543]), .B(y[543]), .Z(n14495) );
  AND U13410 ( .A(n5912), .B(n14495), .Z(n5913) );
  NAND U13411 ( .A(n14492), .B(n5913), .Z(n5914) );
  NANDN U13412 ( .A(n14493), .B(n5914), .Z(n5915) );
  NANDN U13413 ( .A(y[545]), .B(x[545]), .Z(n14490) );
  NANDN U13414 ( .A(n5915), .B(n14490), .Z(n5916) );
  AND U13415 ( .A(n5917), .B(n5916), .Z(n5919) );
  NANDN U13416 ( .A(y[547]), .B(x[547]), .Z(n14486) );
  ANDN U13417 ( .B(x[546]), .A(y[546]), .Z(n14489) );
  ANDN U13418 ( .B(n14486), .A(n14489), .Z(n5918) );
  NANDN U13419 ( .A(n5919), .B(n5918), .Z(n5920) );
  AND U13420 ( .A(n14487), .B(n5920), .Z(n5921) );
  NANDN U13421 ( .A(x[548]), .B(y[548]), .Z(n14484) );
  NAND U13422 ( .A(n5921), .B(n14484), .Z(n5922) );
  ANDN U13423 ( .B(x[549]), .A(y[549]), .Z(n14481) );
  ANDN U13424 ( .B(n5922), .A(n14481), .Z(n5923) );
  NANDN U13425 ( .A(n14485), .B(n5923), .Z(n5924) );
  NANDN U13426 ( .A(x[549]), .B(y[549]), .Z(n14483) );
  AND U13427 ( .A(n5924), .B(n14483), .Z(n5925) );
  NAND U13428 ( .A(n14479), .B(n5925), .Z(n5926) );
  NAND U13429 ( .A(n14482), .B(n5926), .Z(n5927) );
  ANDN U13430 ( .B(x[551]), .A(y[551]), .Z(n14478) );
  OR U13431 ( .A(n5927), .B(n14478), .Z(n5928) );
  AND U13432 ( .A(n5929), .B(n5928), .Z(n5932) );
  ANDN U13433 ( .B(x[553]), .A(y[553]), .Z(n14474) );
  ANDN U13434 ( .B(x[552]), .A(y[552]), .Z(n5930) );
  NOR U13435 ( .A(n14474), .B(n5930), .Z(n5931) );
  NANDN U13436 ( .A(n5932), .B(n5931), .Z(n5933) );
  AND U13437 ( .A(n14475), .B(n5933), .Z(n5934) );
  NANDN U13438 ( .A(x[554]), .B(y[554]), .Z(n14472) );
  NAND U13439 ( .A(n5934), .B(n14472), .Z(n5935) );
  NANDN U13440 ( .A(n5936), .B(n5935), .Z(n5937) );
  AND U13441 ( .A(n14471), .B(n5937), .Z(n5938) );
  NANDN U13442 ( .A(x[556]), .B(y[556]), .Z(n14467) );
  NAND U13443 ( .A(n5938), .B(n14467), .Z(n5939) );
  ANDN U13444 ( .B(x[557]), .A(y[557]), .Z(n14465) );
  ANDN U13445 ( .B(n5939), .A(n14465), .Z(n5940) );
  NANDN U13446 ( .A(n14469), .B(n5940), .Z(n5941) );
  AND U13447 ( .A(n14466), .B(n5941), .Z(n5942) );
  NAND U13448 ( .A(n14468), .B(n5942), .Z(n5943) );
  NANDN U13449 ( .A(n5944), .B(n5943), .Z(n5945) );
  NANDN U13450 ( .A(x[559]), .B(y[559]), .Z(n14463) );
  NAND U13451 ( .A(n5945), .B(n14463), .Z(n5946) );
  NANDN U13452 ( .A(n14462), .B(n5946), .Z(n5947) );
  AND U13453 ( .A(n14460), .B(n5947), .Z(n5950) );
  ANDN U13454 ( .B(x[561]), .A(y[561]), .Z(n14457) );
  ANDN U13455 ( .B(x[560]), .A(y[560]), .Z(n5948) );
  NOR U13456 ( .A(n14457), .B(n5948), .Z(n5949) );
  NANDN U13457 ( .A(n5950), .B(n5949), .Z(n5951) );
  AND U13458 ( .A(n14459), .B(n5951), .Z(n5952) );
  NANDN U13459 ( .A(x[562]), .B(y[562]), .Z(n14456) );
  NAND U13460 ( .A(n5952), .B(n14456), .Z(n5953) );
  NANDN U13461 ( .A(y[563]), .B(x[563]), .Z(n14454) );
  AND U13462 ( .A(n5953), .B(n14454), .Z(n5954) );
  NAND U13463 ( .A(n14458), .B(n5954), .Z(n5955) );
  NANDN U13464 ( .A(x[563]), .B(y[563]), .Z(n14455) );
  AND U13465 ( .A(n5955), .B(n14455), .Z(n5956) );
  NAND U13466 ( .A(n14452), .B(n5956), .Z(n5957) );
  NANDN U13467 ( .A(n14453), .B(n5957), .Z(n5958) );
  ANDN U13468 ( .B(x[565]), .A(y[565]), .Z(n14450) );
  OR U13469 ( .A(n5958), .B(n14450), .Z(n5959) );
  AND U13470 ( .A(n5960), .B(n5959), .Z(n5963) );
  ANDN U13471 ( .B(x[566]), .A(y[566]), .Z(n5961) );
  ANDN U13472 ( .B(x[567]), .A(y[567]), .Z(n25634) );
  NOR U13473 ( .A(n5961), .B(n25634), .Z(n5962) );
  NANDN U13474 ( .A(n5963), .B(n5962), .Z(n5964) );
  XNOR U13475 ( .A(x[568]), .B(y[568]), .Z(n24538) );
  AND U13476 ( .A(n5964), .B(n24538), .Z(n5965) );
  NANDN U13477 ( .A(x[567]), .B(y[567]), .Z(n14447) );
  NAND U13478 ( .A(n5965), .B(n14447), .Z(n5966) );
  ANDN U13479 ( .B(x[569]), .A(y[569]), .Z(n14443) );
  ANDN U13480 ( .B(n5966), .A(n14443), .Z(n5967) );
  NANDN U13481 ( .A(n16074), .B(n5967), .Z(n5968) );
  NANDN U13482 ( .A(x[569]), .B(y[569]), .Z(n14445) );
  AND U13483 ( .A(n5968), .B(n14445), .Z(n5969) );
  NAND U13484 ( .A(n14441), .B(n5969), .Z(n5970) );
  NAND U13485 ( .A(n14444), .B(n5970), .Z(n5971) );
  NANDN U13486 ( .A(y[571]), .B(x[571]), .Z(n14440) );
  NANDN U13487 ( .A(n5971), .B(n14440), .Z(n5972) );
  AND U13488 ( .A(n5973), .B(n5972), .Z(n5975) );
  NANDN U13489 ( .A(y[573]), .B(x[573]), .Z(n14436) );
  ANDN U13490 ( .B(x[572]), .A(y[572]), .Z(n14439) );
  ANDN U13491 ( .B(n14436), .A(n14439), .Z(n5974) );
  NANDN U13492 ( .A(n5975), .B(n5974), .Z(n5976) );
  AND U13493 ( .A(n14438), .B(n5976), .Z(n5977) );
  NAND U13494 ( .A(n5978), .B(n5977), .Z(n5979) );
  NAND U13495 ( .A(n14435), .B(n5979), .Z(n5980) );
  AND U13496 ( .A(n14434), .B(n5980), .Z(n5983) );
  NANDN U13497 ( .A(y[575]), .B(x[575]), .Z(n5982) );
  NANDN U13498 ( .A(y[576]), .B(x[576]), .Z(n5981) );
  NAND U13499 ( .A(n5982), .B(n5981), .Z(n25642) );
  OR U13500 ( .A(n5983), .B(n25642), .Z(n5984) );
  NAND U13501 ( .A(n25643), .B(n5984), .Z(n5985) );
  NANDN U13502 ( .A(n14432), .B(n5985), .Z(n5986) );
  NANDN U13503 ( .A(x[578]), .B(y[578]), .Z(n14430) );
  NAND U13504 ( .A(n5986), .B(n14430), .Z(n5987) );
  ANDN U13505 ( .B(x[579]), .A(y[579]), .Z(n25647) );
  ANDN U13506 ( .B(n5987), .A(n25647), .Z(n5988) );
  NANDN U13507 ( .A(n5989), .B(n5988), .Z(n5990) );
  XNOR U13508 ( .A(x[580]), .B(y[580]), .Z(n25646) );
  AND U13509 ( .A(n5990), .B(n25646), .Z(n5991) );
  NAND U13510 ( .A(n14429), .B(n5991), .Z(n5992) );
  NANDN U13511 ( .A(n16087), .B(n5992), .Z(n5993) );
  ANDN U13512 ( .B(x[581]), .A(y[581]), .Z(n14426) );
  OR U13513 ( .A(n5993), .B(n14426), .Z(n5994) );
  AND U13514 ( .A(n5995), .B(n5994), .Z(n5998) );
  ANDN U13515 ( .B(x[583]), .A(y[583]), .Z(n14422) );
  ANDN U13516 ( .B(x[582]), .A(y[582]), .Z(n5996) );
  NOR U13517 ( .A(n14422), .B(n5996), .Z(n5997) );
  NANDN U13518 ( .A(n5998), .B(n5997), .Z(n5999) );
  AND U13519 ( .A(n14423), .B(n5999), .Z(n6000) );
  NANDN U13520 ( .A(x[584]), .B(y[584]), .Z(n14420) );
  NAND U13521 ( .A(n6000), .B(n14420), .Z(n6001) );
  NANDN U13522 ( .A(y[585]), .B(x[585]), .Z(n14418) );
  AND U13523 ( .A(n6001), .B(n14418), .Z(n6002) );
  NANDN U13524 ( .A(n6003), .B(n6002), .Z(n6004) );
  NANDN U13525 ( .A(x[585]), .B(y[585]), .Z(n14419) );
  AND U13526 ( .A(n6004), .B(n14419), .Z(n6005) );
  NAND U13527 ( .A(n14416), .B(n6005), .Z(n6006) );
  NANDN U13528 ( .A(n14417), .B(n6006), .Z(n6007) );
  ANDN U13529 ( .B(x[587]), .A(y[587]), .Z(n14414) );
  OR U13530 ( .A(n6007), .B(n14414), .Z(n6008) );
  AND U13531 ( .A(n6009), .B(n6008), .Z(n6012) );
  ANDN U13532 ( .B(x[589]), .A(y[589]), .Z(n14409) );
  ANDN U13533 ( .B(x[588]), .A(y[588]), .Z(n6010) );
  NOR U13534 ( .A(n14409), .B(n6010), .Z(n6011) );
  NANDN U13535 ( .A(n6012), .B(n6011), .Z(n6013) );
  AND U13536 ( .A(n14411), .B(n6013), .Z(n6014) );
  NAND U13537 ( .A(n6015), .B(n6014), .Z(n6016) );
  NAND U13538 ( .A(n14410), .B(n6016), .Z(n6017) );
  AND U13539 ( .A(n14408), .B(n6017), .Z(n6020) );
  NANDN U13540 ( .A(y[591]), .B(x[591]), .Z(n6019) );
  NANDN U13541 ( .A(y[592]), .B(x[592]), .Z(n6018) );
  NAND U13542 ( .A(n6019), .B(n6018), .Z(n25670) );
  OR U13543 ( .A(n6020), .B(n25670), .Z(n6021) );
  NAND U13544 ( .A(n25672), .B(n6021), .Z(n6022) );
  NANDN U13545 ( .A(n6023), .B(n6022), .Z(n6024) );
  NAND U13546 ( .A(n25676), .B(n6024), .Z(n6025) );
  NANDN U13547 ( .A(n14403), .B(n6025), .Z(n6026) );
  AND U13548 ( .A(n14402), .B(n6026), .Z(n6028) );
  NANDN U13549 ( .A(y[596]), .B(x[596]), .Z(n14404) );
  ANDN U13550 ( .B(x[597]), .A(y[597]), .Z(n14399) );
  ANDN U13551 ( .B(n14404), .A(n14399), .Z(n6027) );
  NANDN U13552 ( .A(n6028), .B(n6027), .Z(n6029) );
  AND U13553 ( .A(n14401), .B(n6029), .Z(n6030) );
  NAND U13554 ( .A(n6031), .B(n6030), .Z(n6032) );
  NAND U13555 ( .A(n14400), .B(n6032), .Z(n6033) );
  AND U13556 ( .A(n14398), .B(n6033), .Z(n6034) );
  ANDN U13557 ( .B(x[599]), .A(y[599]), .Z(n14395) );
  OR U13558 ( .A(n6034), .B(n14395), .Z(n6035) );
  NAND U13559 ( .A(n14393), .B(n6035), .Z(n6036) );
  NAND U13560 ( .A(n14396), .B(n6036), .Z(n6037) );
  ANDN U13561 ( .B(x[601]), .A(y[601]), .Z(n14391) );
  OR U13562 ( .A(n6037), .B(n14391), .Z(n6038) );
  AND U13563 ( .A(n6039), .B(n6038), .Z(n6041) );
  NANDN U13564 ( .A(y[602]), .B(x[602]), .Z(n14392) );
  ANDN U13565 ( .B(x[603]), .A(y[603]), .Z(n14387) );
  ANDN U13566 ( .B(n14392), .A(n14387), .Z(n6040) );
  NANDN U13567 ( .A(n6041), .B(n6040), .Z(n6042) );
  AND U13568 ( .A(n14389), .B(n6042), .Z(n6043) );
  NANDN U13569 ( .A(x[604]), .B(y[604]), .Z(n14386) );
  NAND U13570 ( .A(n6043), .B(n14386), .Z(n6044) );
  ANDN U13571 ( .B(x[605]), .A(y[605]), .Z(n14383) );
  ANDN U13572 ( .B(n6044), .A(n14383), .Z(n6045) );
  NAND U13573 ( .A(n14388), .B(n6045), .Z(n6046) );
  NANDN U13574 ( .A(x[605]), .B(y[605]), .Z(n14385) );
  AND U13575 ( .A(n6046), .B(n14385), .Z(n6047) );
  NAND U13576 ( .A(n14381), .B(n6047), .Z(n6048) );
  NAND U13577 ( .A(n14384), .B(n6048), .Z(n6049) );
  ANDN U13578 ( .B(x[607]), .A(y[607]), .Z(n14379) );
  OR U13579 ( .A(n6049), .B(n14379), .Z(n6050) );
  AND U13580 ( .A(n6051), .B(n6050), .Z(n6053) );
  NANDN U13581 ( .A(y[608]), .B(x[608]), .Z(n14380) );
  ANDN U13582 ( .B(x[609]), .A(y[609]), .Z(n14375) );
  ANDN U13583 ( .B(n14380), .A(n14375), .Z(n6052) );
  NANDN U13584 ( .A(n6053), .B(n6052), .Z(n6054) );
  AND U13585 ( .A(n14378), .B(n6054), .Z(n6055) );
  NANDN U13586 ( .A(x[610]), .B(y[610]), .Z(n14374) );
  NAND U13587 ( .A(n6055), .B(n14374), .Z(n6056) );
  ANDN U13588 ( .B(x[611]), .A(y[611]), .Z(n14372) );
  ANDN U13589 ( .B(n6056), .A(n14372), .Z(n6057) );
  NAND U13590 ( .A(n14376), .B(n6057), .Z(n6058) );
  NANDN U13591 ( .A(x[611]), .B(y[611]), .Z(n14373) );
  AND U13592 ( .A(n6058), .B(n14373), .Z(n6059) );
  NAND U13593 ( .A(n14370), .B(n6059), .Z(n6060) );
  NANDN U13594 ( .A(n6061), .B(n6060), .Z(n6062) );
  ANDN U13595 ( .B(x[613]), .A(y[613]), .Z(n14368) );
  OR U13596 ( .A(n6062), .B(n14368), .Z(n6063) );
  AND U13597 ( .A(n6064), .B(n6063), .Z(n6067) );
  ANDN U13598 ( .B(x[615]), .A(y[615]), .Z(n14363) );
  ANDN U13599 ( .B(x[614]), .A(y[614]), .Z(n6065) );
  NOR U13600 ( .A(n14363), .B(n6065), .Z(n6066) );
  NANDN U13601 ( .A(n6067), .B(n6066), .Z(n6068) );
  AND U13602 ( .A(n14365), .B(n6068), .Z(n6069) );
  NANDN U13603 ( .A(x[616]), .B(y[616]), .Z(n14361) );
  NAND U13604 ( .A(n6069), .B(n14361), .Z(n6070) );
  NANDN U13605 ( .A(y[617]), .B(x[617]), .Z(n14360) );
  AND U13606 ( .A(n6070), .B(n14360), .Z(n6071) );
  NAND U13607 ( .A(n14364), .B(n6071), .Z(n6072) );
  NANDN U13608 ( .A(x[617]), .B(y[617]), .Z(n14362) );
  AND U13609 ( .A(n6072), .B(n14362), .Z(n6073) );
  NAND U13610 ( .A(n14358), .B(n6073), .Z(n6074) );
  NANDN U13611 ( .A(n14359), .B(n6074), .Z(n6075) );
  NANDN U13612 ( .A(y[619]), .B(x[619]), .Z(n14356) );
  NANDN U13613 ( .A(n6075), .B(n14356), .Z(n6076) );
  AND U13614 ( .A(n6077), .B(n6076), .Z(n6079) );
  NANDN U13615 ( .A(y[621]), .B(x[621]), .Z(n14352) );
  ANDN U13616 ( .B(x[620]), .A(y[620]), .Z(n14355) );
  ANDN U13617 ( .B(n14352), .A(n14355), .Z(n6078) );
  NANDN U13618 ( .A(n6079), .B(n6078), .Z(n6080) );
  AND U13619 ( .A(n14353), .B(n6080), .Z(n6081) );
  NANDN U13620 ( .A(x[622]), .B(y[622]), .Z(n14350) );
  NAND U13621 ( .A(n6081), .B(n14350), .Z(n6082) );
  ANDN U13622 ( .B(x[623]), .A(y[623]), .Z(n14347) );
  ANDN U13623 ( .B(n6082), .A(n14347), .Z(n6083) );
  NANDN U13624 ( .A(n14351), .B(n6083), .Z(n6084) );
  AND U13625 ( .A(n14348), .B(n6084), .Z(n6085) );
  NAND U13626 ( .A(n14349), .B(n6085), .Z(n6086) );
  NANDN U13627 ( .A(n6087), .B(n6086), .Z(n6088) );
  ANDN U13628 ( .B(x[625]), .A(y[625]), .Z(n14344) );
  OR U13629 ( .A(n6088), .B(n14344), .Z(n6089) );
  AND U13630 ( .A(n6090), .B(n6089), .Z(n6093) );
  NANDN U13631 ( .A(y[627]), .B(x[627]), .Z(n14340) );
  ANDN U13632 ( .B(x[626]), .A(y[626]), .Z(n6091) );
  ANDN U13633 ( .B(n14340), .A(n6091), .Z(n6092) );
  NANDN U13634 ( .A(n6093), .B(n6092), .Z(n6094) );
  AND U13635 ( .A(n14341), .B(n6094), .Z(n6095) );
  NANDN U13636 ( .A(x[628]), .B(y[628]), .Z(n14337) );
  NAND U13637 ( .A(n6095), .B(n14337), .Z(n6096) );
  ANDN U13638 ( .B(x[629]), .A(y[629]), .Z(n14335) );
  ANDN U13639 ( .B(n6096), .A(n14335), .Z(n6097) );
  NANDN U13640 ( .A(n14339), .B(n6097), .Z(n6098) );
  NANDN U13641 ( .A(x[629]), .B(y[629]), .Z(n14338) );
  AND U13642 ( .A(n6098), .B(n14338), .Z(n6099) );
  NAND U13643 ( .A(n14334), .B(n6099), .Z(n6100) );
  NAND U13644 ( .A(n14336), .B(n6100), .Z(n6101) );
  NANDN U13645 ( .A(y[631]), .B(x[631]), .Z(n14332) );
  NANDN U13646 ( .A(n6101), .B(n14332), .Z(n6102) );
  AND U13647 ( .A(n6103), .B(n6102), .Z(n6105) );
  NANDN U13648 ( .A(y[633]), .B(x[633]), .Z(n14328) );
  ANDN U13649 ( .B(x[632]), .A(y[632]), .Z(n14331) );
  ANDN U13650 ( .B(n14328), .A(n14331), .Z(n6104) );
  NANDN U13651 ( .A(n6105), .B(n6104), .Z(n6106) );
  AND U13652 ( .A(n14329), .B(n6106), .Z(n6107) );
  NANDN U13653 ( .A(x[634]), .B(y[634]), .Z(n14326) );
  NAND U13654 ( .A(n6107), .B(n14326), .Z(n6108) );
  NANDN U13655 ( .A(y[635]), .B(x[635]), .Z(n14324) );
  AND U13656 ( .A(n6108), .B(n14324), .Z(n6109) );
  NANDN U13657 ( .A(n14327), .B(n6109), .Z(n6110) );
  NANDN U13658 ( .A(x[635]), .B(y[635]), .Z(n14325) );
  AND U13659 ( .A(n6110), .B(n14325), .Z(n6111) );
  NAND U13660 ( .A(n14321), .B(n6111), .Z(n6112) );
  NANDN U13661 ( .A(n14323), .B(n6112), .Z(n6113) );
  ANDN U13662 ( .B(x[637]), .A(y[637]), .Z(n14320) );
  OR U13663 ( .A(n6113), .B(n14320), .Z(n6114) );
  AND U13664 ( .A(n6115), .B(n6114), .Z(n6118) );
  NANDN U13665 ( .A(y[639]), .B(x[639]), .Z(n14316) );
  ANDN U13666 ( .B(x[638]), .A(y[638]), .Z(n6116) );
  ANDN U13667 ( .B(n14316), .A(n6116), .Z(n6117) );
  NANDN U13668 ( .A(n6118), .B(n6117), .Z(n6119) );
  AND U13669 ( .A(n14317), .B(n6119), .Z(n6120) );
  NANDN U13670 ( .A(x[640]), .B(y[640]), .Z(n14314) );
  NAND U13671 ( .A(n6120), .B(n14314), .Z(n6121) );
  NANDN U13672 ( .A(y[641]), .B(x[641]), .Z(n14312) );
  AND U13673 ( .A(n6121), .B(n14312), .Z(n6122) );
  NANDN U13674 ( .A(n14315), .B(n6122), .Z(n6123) );
  NANDN U13675 ( .A(x[641]), .B(y[641]), .Z(n14313) );
  AND U13676 ( .A(n6123), .B(n14313), .Z(n6124) );
  NAND U13677 ( .A(n14310), .B(n6124), .Z(n6125) );
  NANDN U13678 ( .A(n14311), .B(n6125), .Z(n6126) );
  NANDN U13679 ( .A(y[643]), .B(x[643]), .Z(n14308) );
  NANDN U13680 ( .A(n6126), .B(n14308), .Z(n6127) );
  AND U13681 ( .A(n6128), .B(n6127), .Z(n6130) );
  NANDN U13682 ( .A(y[645]), .B(x[645]), .Z(n14304) );
  ANDN U13683 ( .B(x[644]), .A(y[644]), .Z(n14307) );
  ANDN U13684 ( .B(n14304), .A(n14307), .Z(n6129) );
  NANDN U13685 ( .A(n6130), .B(n6129), .Z(n6131) );
  AND U13686 ( .A(n14306), .B(n6131), .Z(n6132) );
  NANDN U13687 ( .A(x[646]), .B(y[646]), .Z(n14301) );
  NAND U13688 ( .A(n6132), .B(n14301), .Z(n6133) );
  NAND U13689 ( .A(n14303), .B(n6133), .Z(n6134) );
  AND U13690 ( .A(n14302), .B(n6134), .Z(n6135) );
  ANDN U13691 ( .B(x[647]), .A(y[647]), .Z(n14299) );
  OR U13692 ( .A(n6135), .B(n14299), .Z(n6136) );
  NAND U13693 ( .A(n14300), .B(n6136), .Z(n6137) );
  NANDN U13694 ( .A(n6138), .B(n6137), .Z(n6139) );
  ANDN U13695 ( .B(x[649]), .A(y[649]), .Z(n14295) );
  OR U13696 ( .A(n6139), .B(n14295), .Z(n6140) );
  AND U13697 ( .A(n6141), .B(n6140), .Z(n6144) );
  ANDN U13698 ( .B(x[651]), .A(y[651]), .Z(n14291) );
  ANDN U13699 ( .B(x[650]), .A(y[650]), .Z(n6142) );
  NOR U13700 ( .A(n14291), .B(n6142), .Z(n6143) );
  NANDN U13701 ( .A(n6144), .B(n6143), .Z(n6145) );
  AND U13702 ( .A(n14293), .B(n6145), .Z(n6146) );
  NAND U13703 ( .A(n14292), .B(n6146), .Z(n6148) );
  ANDN U13704 ( .B(x[652]), .A(y[652]), .Z(n6147) );
  ANDN U13705 ( .B(n6148), .A(n6147), .Z(n6149) );
  NANDN U13706 ( .A(n14287), .B(n6149), .Z(n6150) );
  NANDN U13707 ( .A(x[653]), .B(y[653]), .Z(n14289) );
  AND U13708 ( .A(n6150), .B(n14289), .Z(n6151) );
  NAND U13709 ( .A(n14285), .B(n6151), .Z(n6152) );
  NAND U13710 ( .A(n14288), .B(n6152), .Z(n6153) );
  ANDN U13711 ( .B(x[655]), .A(y[655]), .Z(n14283) );
  OR U13712 ( .A(n6153), .B(n14283), .Z(n6154) );
  AND U13713 ( .A(n6155), .B(n6154), .Z(n6157) );
  NANDN U13714 ( .A(y[657]), .B(x[657]), .Z(n14280) );
  NANDN U13715 ( .A(y[656]), .B(x[656]), .Z(n14284) );
  AND U13716 ( .A(n14280), .B(n14284), .Z(n6156) );
  NANDN U13717 ( .A(n6157), .B(n6156), .Z(n6158) );
  AND U13718 ( .A(n14281), .B(n6158), .Z(n6159) );
  NANDN U13719 ( .A(x[658]), .B(y[658]), .Z(n14277) );
  NAND U13720 ( .A(n6159), .B(n14277), .Z(n6160) );
  ANDN U13721 ( .B(x[659]), .A(y[659]), .Z(n14276) );
  ANDN U13722 ( .B(n6160), .A(n14276), .Z(n6161) );
  NANDN U13723 ( .A(n14279), .B(n6161), .Z(n6162) );
  NANDN U13724 ( .A(x[659]), .B(y[659]), .Z(n14278) );
  AND U13725 ( .A(n6162), .B(n14278), .Z(n6163) );
  NAND U13726 ( .A(n14274), .B(n6163), .Z(n6164) );
  NANDN U13727 ( .A(n6165), .B(n6164), .Z(n6166) );
  ANDN U13728 ( .B(x[661]), .A(y[661]), .Z(n14271) );
  OR U13729 ( .A(n6166), .B(n14271), .Z(n6167) );
  AND U13730 ( .A(n14273), .B(n6167), .Z(n6168) );
  NAND U13731 ( .A(n6169), .B(n6168), .Z(n6170) );
  NAND U13732 ( .A(n14272), .B(n6170), .Z(n6171) );
  AND U13733 ( .A(n14270), .B(n6171), .Z(n6174) );
  NANDN U13734 ( .A(y[663]), .B(x[663]), .Z(n6173) );
  NANDN U13735 ( .A(y[664]), .B(x[664]), .Z(n6172) );
  NAND U13736 ( .A(n6173), .B(n6172), .Z(n25814) );
  OR U13737 ( .A(n6174), .B(n25814), .Z(n6175) );
  NAND U13738 ( .A(n25816), .B(n6175), .Z(n6176) );
  NANDN U13739 ( .A(n14267), .B(n6176), .Z(n6177) );
  NANDN U13740 ( .A(x[666]), .B(y[666]), .Z(n14265) );
  NAND U13741 ( .A(n6177), .B(n14265), .Z(n6178) );
  ANDN U13742 ( .B(x[667]), .A(y[667]), .Z(n14263) );
  ANDN U13743 ( .B(n6178), .A(n14263), .Z(n6179) );
  NAND U13744 ( .A(n14268), .B(n6179), .Z(n6180) );
  NANDN U13745 ( .A(x[667]), .B(y[667]), .Z(n14266) );
  AND U13746 ( .A(n6180), .B(n14266), .Z(n6181) );
  NAND U13747 ( .A(n14262), .B(n6181), .Z(n6182) );
  NAND U13748 ( .A(n14264), .B(n6182), .Z(n6183) );
  NANDN U13749 ( .A(y[669]), .B(x[669]), .Z(n14260) );
  NANDN U13750 ( .A(n6183), .B(n14260), .Z(n6184) );
  AND U13751 ( .A(n6185), .B(n6184), .Z(n6187) );
  ANDN U13752 ( .B(x[670]), .A(y[670]), .Z(n14259) );
  ANDN U13753 ( .B(x[671]), .A(y[671]), .Z(n14256) );
  NOR U13754 ( .A(n14259), .B(n14256), .Z(n6186) );
  NANDN U13755 ( .A(n6187), .B(n6186), .Z(n6188) );
  AND U13756 ( .A(n14257), .B(n6188), .Z(n6189) );
  NANDN U13757 ( .A(x[672]), .B(y[672]), .Z(n14254) );
  NAND U13758 ( .A(n6189), .B(n14254), .Z(n6190) );
  ANDN U13759 ( .B(x[673]), .A(y[673]), .Z(n14251) );
  ANDN U13760 ( .B(n6190), .A(n14251), .Z(n6191) );
  NANDN U13761 ( .A(n6192), .B(n6191), .Z(n6193) );
  NANDN U13762 ( .A(x[673]), .B(y[673]), .Z(n14253) );
  AND U13763 ( .A(n6193), .B(n14253), .Z(n6194) );
  NAND U13764 ( .A(n14250), .B(n6194), .Z(n6195) );
  NAND U13765 ( .A(n14252), .B(n6195), .Z(n6196) );
  ANDN U13766 ( .B(x[675]), .A(y[675]), .Z(n14248) );
  OR U13767 ( .A(n6196), .B(n14248), .Z(n6197) );
  AND U13768 ( .A(n6198), .B(n6197), .Z(n6201) );
  ANDN U13769 ( .B(x[677]), .A(y[677]), .Z(n14244) );
  ANDN U13770 ( .B(x[676]), .A(y[676]), .Z(n6199) );
  NOR U13771 ( .A(n14244), .B(n6199), .Z(n6200) );
  NANDN U13772 ( .A(n6201), .B(n6200), .Z(n6202) );
  AND U13773 ( .A(n14245), .B(n6202), .Z(n6203) );
  NANDN U13774 ( .A(x[678]), .B(y[678]), .Z(n14242) );
  NAND U13775 ( .A(n6203), .B(n14242), .Z(n6204) );
  NANDN U13776 ( .A(y[679]), .B(x[679]), .Z(n14240) );
  AND U13777 ( .A(n6204), .B(n14240), .Z(n6205) );
  NANDN U13778 ( .A(n6206), .B(n6205), .Z(n6207) );
  NANDN U13779 ( .A(x[679]), .B(y[679]), .Z(n14241) );
  AND U13780 ( .A(n6207), .B(n14241), .Z(n6208) );
  NAND U13781 ( .A(n14238), .B(n6208), .Z(n6209) );
  NANDN U13782 ( .A(n14239), .B(n6209), .Z(n6210) );
  OR U13783 ( .A(n14236), .B(n6210), .Z(n6211) );
  AND U13784 ( .A(n14237), .B(n6211), .Z(n6212) );
  NANDN U13785 ( .A(n14233), .B(n6212), .Z(n6213) );
  NAND U13786 ( .A(n6214), .B(n6213), .Z(n6215) );
  NANDN U13787 ( .A(x[683]), .B(y[683]), .Z(n14234) );
  AND U13788 ( .A(n6215), .B(n14234), .Z(n6216) );
  NAND U13789 ( .A(n14231), .B(n6216), .Z(n6217) );
  NANDN U13790 ( .A(n6218), .B(n6217), .Z(n6219) );
  ANDN U13791 ( .B(x[685]), .A(y[685]), .Z(n16195) );
  OR U13792 ( .A(n6219), .B(n16195), .Z(n6220) );
  AND U13793 ( .A(n14230), .B(n6220), .Z(n6221) );
  NANDN U13794 ( .A(x[686]), .B(y[686]), .Z(n14229) );
  NAND U13795 ( .A(n6221), .B(n14229), .Z(n6222) );
  ANDN U13796 ( .B(x[687]), .A(y[687]), .Z(n14226) );
  ANDN U13797 ( .B(n6222), .A(n14226), .Z(n6223) );
  NANDN U13798 ( .A(n6224), .B(n6223), .Z(n6225) );
  ANDN U13799 ( .B(y[688]), .A(x[688]), .Z(n25856) );
  ANDN U13800 ( .B(n6225), .A(n25856), .Z(n6226) );
  NAND U13801 ( .A(n14228), .B(n6226), .Z(n6227) );
  NAND U13802 ( .A(n25857), .B(n6227), .Z(n6228) );
  NANDN U13803 ( .A(y[688]), .B(x[688]), .Z(n14227) );
  NANDN U13804 ( .A(n6228), .B(n14227), .Z(n6229) );
  AND U13805 ( .A(n25858), .B(n6229), .Z(n6230) );
  NANDN U13806 ( .A(y[690]), .B(x[690]), .Z(n16203) );
  NANDN U13807 ( .A(y[691]), .B(x[691]), .Z(n16209) );
  AND U13808 ( .A(n16203), .B(n16209), .Z(n24536) );
  NANDN U13809 ( .A(n6230), .B(n24536), .Z(n6231) );
  NAND U13810 ( .A(n6232), .B(n6231), .Z(n6233) );
  NANDN U13811 ( .A(y[692]), .B(x[692]), .Z(n24535) );
  AND U13812 ( .A(n6233), .B(n24535), .Z(n6234) );
  NAND U13813 ( .A(n14223), .B(n6234), .Z(n6235) );
  NANDN U13814 ( .A(n14224), .B(n6235), .Z(n6236) );
  ANDN U13815 ( .B(y[694]), .A(x[694]), .Z(n14220) );
  OR U13816 ( .A(n6236), .B(n14220), .Z(n6237) );
  AND U13817 ( .A(n14222), .B(n6237), .Z(n6238) );
  NANDN U13818 ( .A(y[695]), .B(x[695]), .Z(n16215) );
  NAND U13819 ( .A(n6238), .B(n16215), .Z(n6239) );
  NAND U13820 ( .A(n14221), .B(n6239), .Z(n6240) );
  ANDN U13821 ( .B(y[696]), .A(x[696]), .Z(n16218) );
  OR U13822 ( .A(n6240), .B(n16218), .Z(n6241) );
  NAND U13823 ( .A(n6242), .B(n6241), .Z(n6243) );
  NANDN U13824 ( .A(n6244), .B(n6243), .Z(n6245) );
  NANDN U13825 ( .A(y[698]), .B(x[698]), .Z(n14218) );
  AND U13826 ( .A(n6245), .B(n14218), .Z(n6246) );
  NAND U13827 ( .A(n14214), .B(n6246), .Z(n6247) );
  NANDN U13828 ( .A(n14215), .B(n6247), .Z(n6248) );
  ANDN U13829 ( .B(y[700]), .A(x[700]), .Z(n14211) );
  OR U13830 ( .A(n6248), .B(n14211), .Z(n6249) );
  AND U13831 ( .A(n14213), .B(n6249), .Z(n6250) );
  NANDN U13832 ( .A(y[701]), .B(x[701]), .Z(n16226) );
  NAND U13833 ( .A(n6250), .B(n16226), .Z(n6251) );
  ANDN U13834 ( .B(y[702]), .A(x[702]), .Z(n16229) );
  ANDN U13835 ( .B(n6251), .A(n16229), .Z(n6252) );
  NANDN U13836 ( .A(n14210), .B(n6252), .Z(n6254) );
  NANDN U13837 ( .A(y[702]), .B(x[702]), .Z(n6253) );
  AND U13838 ( .A(n6254), .B(n6253), .Z(n6255) );
  NAND U13839 ( .A(n14209), .B(n6255), .Z(n6256) );
  NANDN U13840 ( .A(n16228), .B(n6256), .Z(n6257) );
  ANDN U13841 ( .B(y[704]), .A(x[704]), .Z(n14205) );
  OR U13842 ( .A(n6257), .B(n14205), .Z(n6258) );
  NAND U13843 ( .A(n6259), .B(n6258), .Z(n6260) );
  NANDN U13844 ( .A(x[705]), .B(y[705]), .Z(n14207) );
  AND U13845 ( .A(n6260), .B(n14207), .Z(n6261) );
  NAND U13846 ( .A(n14201), .B(n6261), .Z(n6262) );
  NAND U13847 ( .A(n14204), .B(n6262), .Z(n6263) );
  NANDN U13848 ( .A(y[707]), .B(x[707]), .Z(n14199) );
  NANDN U13849 ( .A(n6263), .B(n14199), .Z(n6264) );
  AND U13850 ( .A(n14200), .B(n6264), .Z(n6265) );
  NANDN U13851 ( .A(x[708]), .B(y[708]), .Z(n16238) );
  NAND U13852 ( .A(n6265), .B(n16238), .Z(n6266) );
  ANDN U13853 ( .B(x[709]), .A(y[709]), .Z(n14196) );
  ANDN U13854 ( .B(n6266), .A(n14196), .Z(n6267) );
  ANDN U13855 ( .B(x[708]), .A(y[708]), .Z(n14198) );
  ANDN U13856 ( .B(n6267), .A(n14198), .Z(n6269) );
  NANDN U13857 ( .A(x[710]), .B(y[710]), .Z(n14195) );
  ANDN U13858 ( .B(y[709]), .A(x[709]), .Z(n16237) );
  ANDN U13859 ( .B(n14195), .A(n16237), .Z(n6268) );
  NANDN U13860 ( .A(n6269), .B(n6268), .Z(n6270) );
  AND U13861 ( .A(n14197), .B(n6270), .Z(n6271) );
  NANDN U13862 ( .A(y[711]), .B(x[711]), .Z(n14192) );
  NAND U13863 ( .A(n6271), .B(n14192), .Z(n6272) );
  NAND U13864 ( .A(n14193), .B(n6272), .Z(n6273) );
  ANDN U13865 ( .B(y[711]), .A(x[711]), .Z(n14194) );
  OR U13866 ( .A(n6273), .B(n14194), .Z(n6274) );
  NAND U13867 ( .A(n6275), .B(n6274), .Z(n6276) );
  NANDN U13868 ( .A(n16247), .B(n6276), .Z(n6277) );
  ANDN U13869 ( .B(y[713]), .A(x[713]), .Z(n14191) );
  OR U13870 ( .A(n6277), .B(n14191), .Z(n6278) );
  AND U13871 ( .A(n6279), .B(n6278), .Z(n6280) );
  NANDN U13872 ( .A(n14189), .B(n6280), .Z(n6281) );
  NAND U13873 ( .A(n6282), .B(n6281), .Z(n6283) );
  NANDN U13874 ( .A(y[716]), .B(x[716]), .Z(n14190) );
  AND U13875 ( .A(n6283), .B(n14190), .Z(n6284) );
  NAND U13876 ( .A(n14186), .B(n6284), .Z(n6285) );
  NANDN U13877 ( .A(n14187), .B(n6285), .Z(n6286) );
  ANDN U13878 ( .B(y[718]), .A(x[718]), .Z(n14182) );
  OR U13879 ( .A(n6286), .B(n14182), .Z(n6287) );
  AND U13880 ( .A(n14185), .B(n6287), .Z(n6288) );
  NANDN U13881 ( .A(y[719]), .B(x[719]), .Z(n16255) );
  NAND U13882 ( .A(n6288), .B(n16255), .Z(n6289) );
  ANDN U13883 ( .B(y[720]), .A(x[720]), .Z(n16257) );
  ANDN U13884 ( .B(n6289), .A(n16257), .Z(n6290) );
  NANDN U13885 ( .A(n14183), .B(n6290), .Z(n6291) );
  NANDN U13886 ( .A(y[720]), .B(x[720]), .Z(n16254) );
  AND U13887 ( .A(n6291), .B(n16254), .Z(n6292) );
  NAND U13888 ( .A(n14180), .B(n6292), .Z(n6293) );
  NANDN U13889 ( .A(n16258), .B(n6293), .Z(n6294) );
  XNOR U13890 ( .A(x[722]), .B(y[722]), .Z(n14181) );
  NANDN U13891 ( .A(n6294), .B(n14181), .Z(n6295) );
  NAND U13892 ( .A(n6296), .B(n6295), .Z(n6297) );
  NANDN U13893 ( .A(x[723]), .B(y[723]), .Z(n14178) );
  AND U13894 ( .A(n6297), .B(n14178), .Z(n6298) );
  NAND U13895 ( .A(n14175), .B(n6298), .Z(n6299) );
  NANDN U13896 ( .A(n14176), .B(n6299), .Z(n6300) );
  ANDN U13897 ( .B(x[725]), .A(y[725]), .Z(n14171) );
  OR U13898 ( .A(n6300), .B(n14171), .Z(n6301) );
  NAND U13899 ( .A(n6302), .B(n6301), .Z(n6303) );
  NANDN U13900 ( .A(y[726]), .B(x[726]), .Z(n14173) );
  AND U13901 ( .A(n6303), .B(n14173), .Z(n6304) );
  NAND U13902 ( .A(n14169), .B(n6304), .Z(n6305) );
  NANDN U13903 ( .A(n16266), .B(n6305), .Z(n6306) );
  ANDN U13904 ( .B(y[728]), .A(x[728]), .Z(n14166) );
  OR U13905 ( .A(n6306), .B(n14166), .Z(n6307) );
  AND U13906 ( .A(n14170), .B(n6307), .Z(n6308) );
  NANDN U13907 ( .A(n14164), .B(n6308), .Z(n6309) );
  NAND U13908 ( .A(n6310), .B(n6309), .Z(n6311) );
  NANDN U13909 ( .A(y[730]), .B(x[730]), .Z(n14165) );
  AND U13910 ( .A(n6311), .B(n14165), .Z(n6312) );
  NAND U13911 ( .A(n16274), .B(n6312), .Z(n6313) );
  NANDN U13912 ( .A(n14162), .B(n6313), .Z(n6314) );
  ANDN U13913 ( .B(y[732]), .A(x[732]), .Z(n16277) );
  OR U13914 ( .A(n6314), .B(n16277), .Z(n6315) );
  AND U13915 ( .A(n6316), .B(n6315), .Z(n6317) );
  NANDN U13916 ( .A(y[733]), .B(x[733]), .Z(n14161) );
  NAND U13917 ( .A(n6317), .B(n14161), .Z(n6318) );
  ANDN U13918 ( .B(y[734]), .A(x[734]), .Z(n14159) );
  ANDN U13919 ( .B(n6318), .A(n14159), .Z(n6319) );
  NANDN U13920 ( .A(n16276), .B(n6319), .Z(n6321) );
  NANDN U13921 ( .A(y[734]), .B(x[734]), .Z(n6320) );
  AND U13922 ( .A(n6321), .B(n6320), .Z(n6322) );
  NAND U13923 ( .A(n14156), .B(n6322), .Z(n6323) );
  NANDN U13924 ( .A(n14158), .B(n6323), .Z(n6324) );
  XNOR U13925 ( .A(x[736]), .B(y[736]), .Z(n14157) );
  NANDN U13926 ( .A(n6324), .B(n14157), .Z(n6325) );
  NAND U13927 ( .A(n6326), .B(n6325), .Z(n6327) );
  NANDN U13928 ( .A(x[737]), .B(y[737]), .Z(n14154) );
  AND U13929 ( .A(n6327), .B(n14154), .Z(n6328) );
  NAND U13930 ( .A(n16284), .B(n6328), .Z(n6329) );
  NANDN U13931 ( .A(n14152), .B(n6329), .Z(n6330) );
  ANDN U13932 ( .B(x[739]), .A(y[739]), .Z(n14149) );
  OR U13933 ( .A(n6330), .B(n14149), .Z(n6331) );
  AND U13934 ( .A(n16285), .B(n6331), .Z(n6332) );
  NANDN U13935 ( .A(x[740]), .B(y[740]), .Z(n14148) );
  NAND U13936 ( .A(n6332), .B(n14148), .Z(n6333) );
  ANDN U13937 ( .B(x[741]), .A(y[741]), .Z(n14144) );
  ANDN U13938 ( .B(n6333), .A(n14144), .Z(n6334) );
  NANDN U13939 ( .A(n6335), .B(n6334), .Z(n6336) );
  NANDN U13940 ( .A(x[741]), .B(y[741]), .Z(n14147) );
  AND U13941 ( .A(n6336), .B(n14147), .Z(n6337) );
  NAND U13942 ( .A(n14143), .B(n6337), .Z(n6338) );
  NANDN U13943 ( .A(n6339), .B(n6338), .Z(n6340) );
  ANDN U13944 ( .B(x[743]), .A(y[743]), .Z(n14139) );
  OR U13945 ( .A(n6340), .B(n14139), .Z(n6341) );
  NAND U13946 ( .A(n6342), .B(n6341), .Z(n6343) );
  NANDN U13947 ( .A(y[744]), .B(x[744]), .Z(n14140) );
  AND U13948 ( .A(n6343), .B(n14140), .Z(n6344) );
  NAND U13949 ( .A(n14138), .B(n6344), .Z(n6345) );
  NANDN U13950 ( .A(n16292), .B(n6345), .Z(n6346) );
  ANDN U13951 ( .B(y[746]), .A(x[746]), .Z(n14135) );
  OR U13952 ( .A(n6346), .B(n14135), .Z(n6347) );
  AND U13953 ( .A(n14137), .B(n6347), .Z(n6348) );
  NANDN U13954 ( .A(n14133), .B(n6348), .Z(n6349) );
  NAND U13955 ( .A(n6350), .B(n6349), .Z(n6352) );
  NANDN U13956 ( .A(y[748]), .B(x[748]), .Z(n6351) );
  AND U13957 ( .A(n6352), .B(n6351), .Z(n6353) );
  NAND U13958 ( .A(n16300), .B(n6353), .Z(n6354) );
  NANDN U13959 ( .A(n14132), .B(n6354), .Z(n6355) );
  ANDN U13960 ( .B(y[750]), .A(x[750]), .Z(n16303) );
  OR U13961 ( .A(n6355), .B(n16303), .Z(n6356) );
  AND U13962 ( .A(n6357), .B(n6356), .Z(n6358) );
  NANDN U13963 ( .A(y[751]), .B(x[751]), .Z(n14131) );
  NAND U13964 ( .A(n6358), .B(n14131), .Z(n6359) );
  ANDN U13965 ( .B(y[752]), .A(x[752]), .Z(n14129) );
  ANDN U13966 ( .B(n6359), .A(n14129), .Z(n6360) );
  NANDN U13967 ( .A(n16302), .B(n6360), .Z(n6362) );
  NANDN U13968 ( .A(y[752]), .B(x[752]), .Z(n6361) );
  AND U13969 ( .A(n6362), .B(n6361), .Z(n6363) );
  NAND U13970 ( .A(n14127), .B(n6363), .Z(n6364) );
  NANDN U13971 ( .A(n14128), .B(n6364), .Z(n6365) );
  ANDN U13972 ( .B(y[754]), .A(x[754]), .Z(n14124) );
  OR U13973 ( .A(n6365), .B(n14124), .Z(n6366) );
  AND U13974 ( .A(n6367), .B(n6366), .Z(n6368) );
  NANDN U13975 ( .A(n14121), .B(n6368), .Z(n6369) );
  AND U13976 ( .A(n14125), .B(n6369), .Z(n6370) );
  NANDN U13977 ( .A(x[756]), .B(y[756]), .Z(n16311) );
  NAND U13978 ( .A(n6370), .B(n16311), .Z(n6371) );
  ANDN U13979 ( .B(x[757]), .A(y[757]), .Z(n14119) );
  ANDN U13980 ( .B(n6371), .A(n14119), .Z(n6372) );
  NANDN U13981 ( .A(n6373), .B(n6372), .Z(n6374) );
  NANDN U13982 ( .A(x[757]), .B(y[757]), .Z(n16310) );
  AND U13983 ( .A(n6374), .B(n16310), .Z(n6375) );
  NAND U13984 ( .A(n14118), .B(n6375), .Z(n6376) );
  NAND U13985 ( .A(n14120), .B(n6376), .Z(n6377) );
  ANDN U13986 ( .B(x[759]), .A(y[759]), .Z(n14114) );
  OR U13987 ( .A(n6377), .B(n14114), .Z(n6378) );
  AND U13988 ( .A(n14117), .B(n6378), .Z(n6379) );
  NANDN U13989 ( .A(n14112), .B(n6379), .Z(n6380) );
  AND U13990 ( .A(n6381), .B(n6380), .Z(n6382) );
  NANDN U13991 ( .A(y[761]), .B(x[761]), .Z(n16318) );
  NAND U13992 ( .A(n6382), .B(n16318), .Z(n6383) );
  ANDN U13993 ( .B(y[762]), .A(x[762]), .Z(n16321) );
  ANDN U13994 ( .B(n6383), .A(n16321), .Z(n6384) );
  NANDN U13995 ( .A(n14111), .B(n6384), .Z(n6385) );
  NANDN U13996 ( .A(y[762]), .B(x[762]), .Z(n16317) );
  AND U13997 ( .A(n6385), .B(n16317), .Z(n6386) );
  NAND U13998 ( .A(n14110), .B(n6386), .Z(n6387) );
  NANDN U13999 ( .A(n16320), .B(n6387), .Z(n6388) );
  ANDN U14000 ( .B(y[764]), .A(x[764]), .Z(n14107) );
  OR U14001 ( .A(n6388), .B(n14107), .Z(n6389) );
  NAND U14002 ( .A(n6390), .B(n6389), .Z(n6391) );
  NANDN U14003 ( .A(x[765]), .B(y[765]), .Z(n14108) );
  AND U14004 ( .A(n6391), .B(n14108), .Z(n6392) );
  NAND U14005 ( .A(n14104), .B(n6392), .Z(n6393) );
  NANDN U14006 ( .A(n14105), .B(n6393), .Z(n6394) );
  ANDN U14007 ( .B(x[767]), .A(y[767]), .Z(n14101) );
  OR U14008 ( .A(n6394), .B(n14101), .Z(n6395) );
  AND U14009 ( .A(n14103), .B(n6395), .Z(n6396) );
  NANDN U14010 ( .A(n16329), .B(n6396), .Z(n6397) );
  AND U14011 ( .A(n14102), .B(n6397), .Z(n6398) );
  NANDN U14012 ( .A(y[769]), .B(x[769]), .Z(n14099) );
  NAND U14013 ( .A(n6398), .B(n14099), .Z(n6399) );
  ANDN U14014 ( .B(y[770]), .A(x[770]), .Z(n14098) );
  ANDN U14015 ( .B(n6399), .A(n14098), .Z(n6400) );
  NANDN U14016 ( .A(n16330), .B(n6400), .Z(n6401) );
  NANDN U14017 ( .A(y[770]), .B(x[770]), .Z(n14100) );
  AND U14018 ( .A(n6401), .B(n14100), .Z(n6402) );
  NAND U14019 ( .A(n14095), .B(n6402), .Z(n6403) );
  NANDN U14020 ( .A(n14097), .B(n6403), .Z(n6404) );
  ANDN U14021 ( .B(y[772]), .A(x[772]), .Z(n14093) );
  OR U14022 ( .A(n6404), .B(n14093), .Z(n6405) );
  AND U14023 ( .A(n14096), .B(n6405), .Z(n6406) );
  NAND U14024 ( .A(n6407), .B(n6406), .Z(n6408) );
  NAND U14025 ( .A(n14094), .B(n6408), .Z(n6409) );
  AND U14026 ( .A(n14092), .B(n6409), .Z(n6412) );
  NANDN U14027 ( .A(x[774]), .B(y[774]), .Z(n6411) );
  NANDN U14028 ( .A(x[775]), .B(y[775]), .Z(n6410) );
  NAND U14029 ( .A(n6411), .B(n6410), .Z(n24514) );
  OR U14030 ( .A(n6412), .B(n24514), .Z(n6415) );
  NANDN U14031 ( .A(y[776]), .B(x[776]), .Z(n6414) );
  NANDN U14032 ( .A(y[775]), .B(x[775]), .Z(n6413) );
  AND U14033 ( .A(n6414), .B(n6413), .Z(n24513) );
  AND U14034 ( .A(n6415), .B(n24513), .Z(n6418) );
  NANDN U14035 ( .A(x[776]), .B(y[776]), .Z(n6417) );
  NANDN U14036 ( .A(x[777]), .B(y[777]), .Z(n6416) );
  NAND U14037 ( .A(n6417), .B(n6416), .Z(n25930) );
  OR U14038 ( .A(n6418), .B(n25930), .Z(n6421) );
  NANDN U14039 ( .A(y[778]), .B(x[778]), .Z(n6420) );
  NANDN U14040 ( .A(y[777]), .B(x[777]), .Z(n6419) );
  AND U14041 ( .A(n6420), .B(n6419), .Z(n25931) );
  AND U14042 ( .A(n6421), .B(n25931), .Z(n6424) );
  NANDN U14043 ( .A(x[778]), .B(y[778]), .Z(n6423) );
  NANDN U14044 ( .A(x[779]), .B(y[779]), .Z(n6422) );
  NAND U14045 ( .A(n6423), .B(n6422), .Z(n24512) );
  OR U14046 ( .A(n6424), .B(n24512), .Z(n6425) );
  NAND U14047 ( .A(n24511), .B(n6425), .Z(n6426) );
  NANDN U14048 ( .A(n24510), .B(n6426), .Z(n6427) );
  NANDN U14049 ( .A(n14090), .B(n6427), .Z(n6429) );
  ANDN U14050 ( .B(y[783]), .A(x[783]), .Z(n6431) );
  NANDN U14051 ( .A(x[782]), .B(y[782]), .Z(n6428) );
  NANDN U14052 ( .A(n6431), .B(n6428), .Z(n16346) );
  IV U14053 ( .A(n16346), .Z(n25934) );
  AND U14054 ( .A(n6429), .B(n25934), .Z(n6436) );
  NANDN U14055 ( .A(y[782]), .B(x[782]), .Z(n6430) );
  OR U14056 ( .A(n6431), .B(n6430), .Z(n6434) );
  NANDN U14057 ( .A(y[784]), .B(x[784]), .Z(n6433) );
  NANDN U14058 ( .A(y[783]), .B(x[783]), .Z(n6432) );
  AND U14059 ( .A(n6433), .B(n6432), .Z(n25935) );
  AND U14060 ( .A(n6434), .B(n25935), .Z(n6435) );
  NANDN U14061 ( .A(n6436), .B(n6435), .Z(n6437) );
  NANDN U14062 ( .A(n14089), .B(n6437), .Z(n6438) );
  AND U14063 ( .A(n14087), .B(n6438), .Z(n6439) );
  NAND U14064 ( .A(n6440), .B(n6439), .Z(n6441) );
  NAND U14065 ( .A(n6442), .B(n6441), .Z(n6443) );
  NAND U14066 ( .A(n14084), .B(n6443), .Z(n6444) );
  NANDN U14067 ( .A(n16352), .B(n6444), .Z(n6447) );
  NANDN U14068 ( .A(y[790]), .B(x[790]), .Z(n6446) );
  NANDN U14069 ( .A(y[789]), .B(x[789]), .Z(n6445) );
  AND U14070 ( .A(n6446), .B(n6445), .Z(n16354) );
  AND U14071 ( .A(n6447), .B(n16354), .Z(n6450) );
  NANDN U14072 ( .A(x[790]), .B(y[790]), .Z(n6449) );
  NANDN U14073 ( .A(x[791]), .B(y[791]), .Z(n6448) );
  NAND U14074 ( .A(n6449), .B(n6448), .Z(n14083) );
  OR U14075 ( .A(n6450), .B(n14083), .Z(n6451) );
  NAND U14076 ( .A(n14082), .B(n6451), .Z(n6452) );
  NANDN U14077 ( .A(n14081), .B(n6452), .Z(n6453) );
  NAND U14078 ( .A(n14080), .B(n6453), .Z(n6454) );
  NAND U14079 ( .A(n25946), .B(n6454), .Z(n6455) );
  NANDN U14080 ( .A(n14078), .B(n6455), .Z(n6456) );
  NANDN U14081 ( .A(x[796]), .B(y[796]), .Z(n14076) );
  NAND U14082 ( .A(n6456), .B(n14076), .Z(n6457) );
  NANDN U14083 ( .A(y[797]), .B(x[797]), .Z(n14075) );
  AND U14084 ( .A(n6457), .B(n14075), .Z(n6458) );
  NAND U14085 ( .A(n14079), .B(n6458), .Z(n6459) );
  NANDN U14086 ( .A(x[797]), .B(y[797]), .Z(n14077) );
  AND U14087 ( .A(n6459), .B(n14077), .Z(n6460) );
  NAND U14088 ( .A(n14073), .B(n6460), .Z(n6461) );
  NANDN U14089 ( .A(n14074), .B(n6461), .Z(n6462) );
  ANDN U14090 ( .B(x[799]), .A(y[799]), .Z(n14071) );
  OR U14091 ( .A(n6462), .B(n14071), .Z(n6463) );
  NAND U14092 ( .A(n6464), .B(n6463), .Z(n6466) );
  NANDN U14093 ( .A(y[800]), .B(x[800]), .Z(n6465) );
  AND U14094 ( .A(n6466), .B(n6465), .Z(n6467) );
  NAND U14095 ( .A(n14066), .B(n6467), .Z(n6468) );
  NANDN U14096 ( .A(n14068), .B(n6468), .Z(n6469) );
  NANDN U14097 ( .A(x[802]), .B(y[802]), .Z(n14065) );
  NANDN U14098 ( .A(n6469), .B(n14065), .Z(n6470) );
  AND U14099 ( .A(n14067), .B(n6470), .Z(n6471) );
  NANDN U14100 ( .A(y[803]), .B(x[803]), .Z(n14061) );
  NAND U14101 ( .A(n6471), .B(n14061), .Z(n6472) );
  ANDN U14102 ( .B(y[804]), .A(x[804]), .Z(n14058) );
  ANDN U14103 ( .B(n6472), .A(n14058), .Z(n6473) );
  NANDN U14104 ( .A(n14063), .B(n6473), .Z(n6474) );
  NANDN U14105 ( .A(y[804]), .B(x[804]), .Z(n14062) );
  AND U14106 ( .A(n6474), .B(n14062), .Z(n6475) );
  NAND U14107 ( .A(n14056), .B(n6475), .Z(n6476) );
  NAND U14108 ( .A(n14060), .B(n6476), .Z(n6477) );
  ANDN U14109 ( .B(y[806]), .A(x[806]), .Z(n14052) );
  OR U14110 ( .A(n6477), .B(n14052), .Z(n6478) );
  NAND U14111 ( .A(n6479), .B(n6478), .Z(n6480) );
  NANDN U14112 ( .A(x[807]), .B(y[807]), .Z(n14054) );
  AND U14113 ( .A(n6480), .B(n14054), .Z(n6481) );
  NAND U14114 ( .A(n14047), .B(n6481), .Z(n6482) );
  NANDN U14115 ( .A(n14049), .B(n6482), .Z(n6483) );
  OR U14116 ( .A(n14046), .B(n6483), .Z(n6484) );
  AND U14117 ( .A(n14048), .B(n6484), .Z(n6485) );
  NAND U14118 ( .A(n14044), .B(n6485), .Z(n6486) );
  AND U14119 ( .A(n6487), .B(n6486), .Z(n6488) );
  NAND U14120 ( .A(n14042), .B(n6488), .Z(n6489) );
  NANDN U14121 ( .A(x[812]), .B(y[812]), .Z(n14041) );
  AND U14122 ( .A(n6489), .B(n14041), .Z(n6490) );
  NANDN U14123 ( .A(n14043), .B(n6490), .Z(n6492) );
  NANDN U14124 ( .A(y[812]), .B(x[812]), .Z(n6491) );
  AND U14125 ( .A(n6492), .B(n6491), .Z(n6493) );
  NAND U14126 ( .A(n14039), .B(n6493), .Z(n6494) );
  NANDN U14127 ( .A(n14040), .B(n6494), .Z(n6495) );
  ANDN U14128 ( .B(y[814]), .A(x[814]), .Z(n14036) );
  OR U14129 ( .A(n6495), .B(n14036), .Z(n6496) );
  NAND U14130 ( .A(n6497), .B(n6496), .Z(n6498) );
  NANDN U14131 ( .A(x[815]), .B(y[815]), .Z(n14037) );
  AND U14132 ( .A(n6498), .B(n14037), .Z(n6499) );
  NAND U14133 ( .A(n14033), .B(n6499), .Z(n6500) );
  NAND U14134 ( .A(n14034), .B(n6500), .Z(n6501) );
  ANDN U14135 ( .B(x[817]), .A(y[817]), .Z(n14030) );
  OR U14136 ( .A(n6501), .B(n14030), .Z(n6502) );
  AND U14137 ( .A(n14032), .B(n6502), .Z(n6503) );
  NANDN U14138 ( .A(n14028), .B(n6503), .Z(n6504) );
  NAND U14139 ( .A(n6505), .B(n6504), .Z(n6506) );
  NANDN U14140 ( .A(x[819]), .B(y[819]), .Z(n14029) );
  AND U14141 ( .A(n6506), .B(n14029), .Z(n6507) );
  NAND U14142 ( .A(n14024), .B(n6507), .Z(n6508) );
  NANDN U14143 ( .A(n14026), .B(n6508), .Z(n6509) );
  ANDN U14144 ( .B(x[821]), .A(y[821]), .Z(n14022) );
  OR U14145 ( .A(n6509), .B(n14022), .Z(n6510) );
  AND U14146 ( .A(n14025), .B(n6510), .Z(n6511) );
  NANDN U14147 ( .A(x[822]), .B(y[822]), .Z(n14021) );
  NAND U14148 ( .A(n6511), .B(n14021), .Z(n6512) );
  ANDN U14149 ( .B(x[823]), .A(y[823]), .Z(n25999) );
  ANDN U14150 ( .B(n6512), .A(n25999), .Z(n6513) );
  NAND U14151 ( .A(n14023), .B(n6513), .Z(n6514) );
  NANDN U14152 ( .A(x[824]), .B(y[824]), .Z(n26000) );
  AND U14153 ( .A(n6514), .B(n26000), .Z(n6515) );
  NAND U14154 ( .A(n14020), .B(n6515), .Z(n6516) );
  NANDN U14155 ( .A(n26003), .B(n6516), .Z(n6517) );
  NANDN U14156 ( .A(x[825]), .B(y[825]), .Z(n26005) );
  AND U14157 ( .A(n6517), .B(n26005), .Z(n6518) );
  NAND U14158 ( .A(n26009), .B(n6518), .Z(n6519) );
  NANDN U14159 ( .A(n6520), .B(n6519), .Z(n6521) );
  NAND U14160 ( .A(n26012), .B(n6521), .Z(n6522) );
  NAND U14161 ( .A(n26015), .B(n6522), .Z(n6523) );
  AND U14162 ( .A(n26017), .B(n6523), .Z(n6524) );
  OR U14163 ( .A(n26019), .B(n6524), .Z(n6525) );
  AND U14164 ( .A(n6526), .B(n6525), .Z(n6528) );
  ANDN U14165 ( .B(x[833]), .A(y[833]), .Z(n14016) );
  ANDN U14166 ( .B(x[832]), .A(y[832]), .Z(n26023) );
  NOR U14167 ( .A(n14016), .B(n26023), .Z(n6527) );
  NANDN U14168 ( .A(n6528), .B(n6527), .Z(n6529) );
  AND U14169 ( .A(n14018), .B(n6529), .Z(n6530) );
  NAND U14170 ( .A(n6531), .B(n6530), .Z(n6532) );
  NAND U14171 ( .A(n14017), .B(n6532), .Z(n6533) );
  AND U14172 ( .A(n14015), .B(n6533), .Z(n6534) );
  OR U14173 ( .A(n26031), .B(n6534), .Z(n6535) );
  AND U14174 ( .A(n26033), .B(n6535), .Z(n6538) );
  NANDN U14175 ( .A(y[838]), .B(x[838]), .Z(n6537) );
  NANDN U14176 ( .A(y[837]), .B(x[837]), .Z(n6536) );
  AND U14177 ( .A(n6537), .B(n6536), .Z(n14013) );
  NANDN U14178 ( .A(n6538), .B(n14013), .Z(n6539) );
  NANDN U14179 ( .A(n16421), .B(n6539), .Z(n6540) );
  NANDN U14180 ( .A(y[839]), .B(x[839]), .Z(n14012) );
  AND U14181 ( .A(n6540), .B(n14012), .Z(n6541) );
  ANDN U14182 ( .B(y[840]), .A(x[840]), .Z(n16426) );
  OR U14183 ( .A(n6541), .B(n16426), .Z(n6542) );
  AND U14184 ( .A(n26038), .B(n6542), .Z(n6544) );
  NANDN U14185 ( .A(x[841]), .B(y[841]), .Z(n26039) );
  ANDN U14186 ( .B(y[842]), .A(x[842]), .Z(n14010) );
  ANDN U14187 ( .B(n26039), .A(n14010), .Z(n6543) );
  NANDN U14188 ( .A(n6544), .B(n6543), .Z(n6545) );
  NANDN U14189 ( .A(n6546), .B(n6545), .Z(n6547) );
  NANDN U14190 ( .A(x[844]), .B(y[844]), .Z(n26043) );
  AND U14191 ( .A(n6547), .B(n26043), .Z(n6548) );
  NAND U14192 ( .A(n14011), .B(n6548), .Z(n6549) );
  NANDN U14193 ( .A(n24509), .B(n6549), .Z(n6551) );
  NANDN U14194 ( .A(x[846]), .B(y[846]), .Z(n14008) );
  NANDN U14195 ( .A(x[845]), .B(y[845]), .Z(n24508) );
  AND U14196 ( .A(n14008), .B(n24508), .Z(n6550) );
  NAND U14197 ( .A(n6551), .B(n6550), .Z(n6552) );
  AND U14198 ( .A(n26044), .B(n6552), .Z(n6555) );
  NANDN U14199 ( .A(x[847]), .B(y[847]), .Z(n6554) );
  NANDN U14200 ( .A(x[848]), .B(y[848]), .Z(n6553) );
  NAND U14201 ( .A(n6554), .B(n6553), .Z(n14009) );
  OR U14202 ( .A(n6555), .B(n14009), .Z(n6556) );
  NANDN U14203 ( .A(n26046), .B(n6556), .Z(n6557) );
  NANDN U14204 ( .A(n26047), .B(n6557), .Z(n6558) );
  ANDN U14205 ( .B(x[850]), .A(y[850]), .Z(n26049) );
  ANDN U14206 ( .B(n6558), .A(n26049), .Z(n6559) );
  NAND U14207 ( .A(n14005), .B(n6559), .Z(n6560) );
  NANDN U14208 ( .A(n26050), .B(n6560), .Z(n6561) );
  ANDN U14209 ( .B(y[852]), .A(x[852]), .Z(n14002) );
  OR U14210 ( .A(n6561), .B(n14002), .Z(n6562) );
  AND U14211 ( .A(n14004), .B(n6562), .Z(n6563) );
  NAND U14212 ( .A(n14001), .B(n6563), .Z(n6564) );
  AND U14213 ( .A(n6565), .B(n6564), .Z(n6567) );
  NANDN U14214 ( .A(y[854]), .B(x[854]), .Z(n14000) );
  ANDN U14215 ( .B(x[855]), .A(y[855]), .Z(n13997) );
  ANDN U14216 ( .B(n14000), .A(n13997), .Z(n6566) );
  NANDN U14217 ( .A(n6567), .B(n6566), .Z(n6568) );
  NANDN U14218 ( .A(x[856]), .B(y[856]), .Z(n13996) );
  AND U14219 ( .A(n6568), .B(n13996), .Z(n6569) );
  NANDN U14220 ( .A(x[855]), .B(y[855]), .Z(n13999) );
  NAND U14221 ( .A(n6569), .B(n13999), .Z(n6570) );
  NANDN U14222 ( .A(n6571), .B(n6570), .Z(n6572) );
  AND U14223 ( .A(n26059), .B(n6572), .Z(n6573) );
  NANDN U14224 ( .A(y[858]), .B(x[858]), .Z(n16458) );
  NANDN U14225 ( .A(y[859]), .B(x[859]), .Z(n16464) );
  NAND U14226 ( .A(n16458), .B(n16464), .Z(n24507) );
  OR U14227 ( .A(n6573), .B(n24507), .Z(n6574) );
  NAND U14228 ( .A(n26060), .B(n6574), .Z(n6575) );
  NANDN U14229 ( .A(n24506), .B(n6575), .Z(n6576) );
  NAND U14230 ( .A(n26061), .B(n6576), .Z(n6577) );
  NAND U14231 ( .A(n26062), .B(n6577), .Z(n6578) );
  NANDN U14232 ( .A(n26063), .B(n6578), .Z(n6579) );
  NAND U14233 ( .A(n26064), .B(n6579), .Z(n6580) );
  ANDN U14234 ( .B(y[866]), .A(x[866]), .Z(n13992) );
  ANDN U14235 ( .B(n6580), .A(n13992), .Z(n6581) );
  NANDN U14236 ( .A(n26066), .B(n6581), .Z(n6582) );
  NANDN U14237 ( .A(y[866]), .B(x[866]), .Z(n26067) );
  AND U14238 ( .A(n6582), .B(n26067), .Z(n6583) );
  NAND U14239 ( .A(n13990), .B(n6583), .Z(n6584) );
  NAND U14240 ( .A(n13993), .B(n6584), .Z(n6585) );
  ANDN U14241 ( .B(y[868]), .A(x[868]), .Z(n13988) );
  OR U14242 ( .A(n6585), .B(n13988), .Z(n6586) );
  AND U14243 ( .A(n13991), .B(n6586), .Z(n6587) );
  NANDN U14244 ( .A(y[869]), .B(x[869]), .Z(n13987) );
  NAND U14245 ( .A(n6587), .B(n13987), .Z(n6588) );
  NANDN U14246 ( .A(x[869]), .B(y[869]), .Z(n13989) );
  AND U14247 ( .A(n6588), .B(n13989), .Z(n6589) );
  NANDN U14248 ( .A(n13986), .B(n6589), .Z(n6590) );
  NANDN U14249 ( .A(y[871]), .B(x[871]), .Z(n26073) );
  AND U14250 ( .A(n6590), .B(n26073), .Z(n6591) );
  NAND U14251 ( .A(n6592), .B(n6591), .Z(n6593) );
  NANDN U14252 ( .A(n13985), .B(n6593), .Z(n6594) );
  ANDN U14253 ( .B(y[872]), .A(x[872]), .Z(n13983) );
  OR U14254 ( .A(n6594), .B(n13983), .Z(n6595) );
  NAND U14255 ( .A(n24505), .B(n6595), .Z(n6596) );
  NANDN U14256 ( .A(n13982), .B(n6596), .Z(n6597) );
  ANDN U14257 ( .B(y[874]), .A(x[874]), .Z(n16499) );
  OR U14258 ( .A(n6597), .B(n16499), .Z(n6598) );
  AND U14259 ( .A(n6599), .B(n6598), .Z(n6601) );
  ANDN U14260 ( .B(y[876]), .A(x[876]), .Z(n16505) );
  IV U14261 ( .A(n16505), .Z(n26078) );
  ANDN U14262 ( .B(y[875]), .A(x[875]), .Z(n16500) );
  ANDN U14263 ( .B(n26078), .A(n16500), .Z(n6600) );
  NANDN U14264 ( .A(n6601), .B(n6600), .Z(n6602) );
  NANDN U14265 ( .A(y[876]), .B(x[876]), .Z(n13980) );
  NANDN U14266 ( .A(y[877]), .B(x[877]), .Z(n16510) );
  AND U14267 ( .A(n13980), .B(n16510), .Z(n24503) );
  AND U14268 ( .A(n6602), .B(n24503), .Z(n6603) );
  ANDN U14269 ( .B(y[877]), .A(x[877]), .Z(n16507) );
  ANDN U14270 ( .B(y[878]), .A(x[878]), .Z(n16515) );
  OR U14271 ( .A(n16507), .B(n16515), .Z(n26079) );
  OR U14272 ( .A(n6603), .B(n26079), .Z(n6604) );
  NAND U14273 ( .A(n26082), .B(n6604), .Z(n6605) );
  NANDN U14274 ( .A(n24502), .B(n6605), .Z(n6606) );
  NANDN U14275 ( .A(n26083), .B(n6606), .Z(n6607) );
  AND U14276 ( .A(n26084), .B(n6607), .Z(n6609) );
  NANDN U14277 ( .A(y[882]), .B(x[882]), .Z(n26085) );
  ANDN U14278 ( .B(x[883]), .A(y[883]), .Z(n13977) );
  ANDN U14279 ( .B(n26085), .A(n13977), .Z(n6608) );
  NANDN U14280 ( .A(n6609), .B(n6608), .Z(n6610) );
  NANDN U14281 ( .A(n26086), .B(n6610), .Z(n6611) );
  ANDN U14282 ( .B(y[884]), .A(x[884]), .Z(n16530) );
  OR U14283 ( .A(n6611), .B(n16530), .Z(n6612) );
  NAND U14284 ( .A(n6613), .B(n6612), .Z(n6614) );
  NANDN U14285 ( .A(x[885]), .B(y[885]), .Z(n16531) );
  AND U14286 ( .A(n6614), .B(n16531), .Z(n6615) );
  NAND U14287 ( .A(n13974), .B(n6615), .Z(n6616) );
  NAND U14288 ( .A(n26090), .B(n6616), .Z(n6617) );
  ANDN U14289 ( .B(x[886]), .A(y[886]), .Z(n13975) );
  OR U14290 ( .A(n6617), .B(n13975), .Z(n6618) );
  AND U14291 ( .A(n13973), .B(n6618), .Z(n6619) );
  NANDN U14292 ( .A(n13972), .B(n6619), .Z(n6620) );
  NANDN U14293 ( .A(y[888]), .B(x[888]), .Z(n16535) );
  NANDN U14294 ( .A(y[889]), .B(x[889]), .Z(n16540) );
  AND U14295 ( .A(n16535), .B(n16540), .Z(n24500) );
  AND U14296 ( .A(n6620), .B(n24500), .Z(n6622) );
  NANDN U14297 ( .A(x[890]), .B(y[890]), .Z(n13969) );
  ANDN U14298 ( .B(y[889]), .A(x[889]), .Z(n13971) );
  ANDN U14299 ( .B(n13969), .A(n13971), .Z(n6621) );
  NANDN U14300 ( .A(n6622), .B(n6621), .Z(n6623) );
  NANDN U14301 ( .A(y[891]), .B(x[891]), .Z(n24499) );
  AND U14302 ( .A(n6623), .B(n24499), .Z(n6624) );
  NAND U14303 ( .A(n26093), .B(n6624), .Z(n6625) );
  NANDN U14304 ( .A(x[892]), .B(y[892]), .Z(n26097) );
  AND U14305 ( .A(n6625), .B(n26097), .Z(n6626) );
  NAND U14306 ( .A(n13970), .B(n6626), .Z(n6627) );
  NANDN U14307 ( .A(n26098), .B(n6627), .Z(n6628) );
  NANDN U14308 ( .A(x[894]), .B(y[894]), .Z(n13968) );
  AND U14309 ( .A(n6628), .B(n13968), .Z(n6629) );
  NAND U14310 ( .A(n26099), .B(n6629), .Z(n6630) );
  NANDN U14311 ( .A(n6631), .B(n6630), .Z(n6632) );
  NANDN U14312 ( .A(x[896]), .B(y[896]), .Z(n26101) );
  AND U14313 ( .A(n6632), .B(n26101), .Z(n6633) );
  NAND U14314 ( .A(n13967), .B(n6633), .Z(n6634) );
  NANDN U14315 ( .A(n26102), .B(n6634), .Z(n6635) );
  NANDN U14316 ( .A(x[898]), .B(y[898]), .Z(n13961) );
  AND U14317 ( .A(n6635), .B(n13961), .Z(n6636) );
  NAND U14318 ( .A(n13965), .B(n6636), .Z(n6637) );
  NAND U14319 ( .A(n26105), .B(n6637), .Z(n6638) );
  ANDN U14320 ( .B(x[899]), .A(y[899]), .Z(n13959) );
  OR U14321 ( .A(n6638), .B(n13959), .Z(n6639) );
  AND U14322 ( .A(n26104), .B(n6639), .Z(n6640) );
  NANDN U14323 ( .A(n13958), .B(n6640), .Z(n6641) );
  AND U14324 ( .A(n13960), .B(n6641), .Z(n6642) );
  NANDN U14325 ( .A(y[901]), .B(x[901]), .Z(n16562) );
  NAND U14326 ( .A(n6642), .B(n16562), .Z(n6643) );
  ANDN U14327 ( .B(y[902]), .A(x[902]), .Z(n16565) );
  ANDN U14328 ( .B(n6643), .A(n16565), .Z(n6644) );
  NANDN U14329 ( .A(n13957), .B(n6644), .Z(n6645) );
  NANDN U14330 ( .A(y[902]), .B(x[902]), .Z(n16561) );
  AND U14331 ( .A(n6645), .B(n16561), .Z(n6646) );
  NAND U14332 ( .A(n13956), .B(n6646), .Z(n6647) );
  NANDN U14333 ( .A(n16564), .B(n6647), .Z(n6648) );
  ANDN U14334 ( .B(y[904]), .A(x[904]), .Z(n13953) );
  OR U14335 ( .A(n6648), .B(n13953), .Z(n6649) );
  NAND U14336 ( .A(n6650), .B(n6649), .Z(n6651) );
  NANDN U14337 ( .A(x[905]), .B(y[905]), .Z(n13954) );
  AND U14338 ( .A(n6651), .B(n13954), .Z(n6652) );
  NAND U14339 ( .A(n13950), .B(n6652), .Z(n6653) );
  NANDN U14340 ( .A(n26115), .B(n6653), .Z(n6654) );
  NANDN U14341 ( .A(y[906]), .B(x[906]), .Z(n13951) );
  NANDN U14342 ( .A(n6654), .B(n13951), .Z(n6655) );
  AND U14343 ( .A(n26116), .B(n6655), .Z(n6656) );
  NANDN U14344 ( .A(x[907]), .B(y[907]), .Z(n13949) );
  NAND U14345 ( .A(n6656), .B(n13949), .Z(n6657) );
  NANDN U14346 ( .A(n26117), .B(n6657), .Z(n6658) );
  AND U14347 ( .A(n26118), .B(n6658), .Z(n6659) );
  NANDN U14348 ( .A(y[910]), .B(x[910]), .Z(n13947) );
  NANDN U14349 ( .A(y[911]), .B(x[911]), .Z(n13944) );
  NAND U14350 ( .A(n13947), .B(n13944), .Z(n24495) );
  OR U14351 ( .A(n6659), .B(n24495), .Z(n6660) );
  NAND U14352 ( .A(n24494), .B(n6660), .Z(n6661) );
  NANDN U14353 ( .A(n24493), .B(n6661), .Z(n6662) );
  NAND U14354 ( .A(n24492), .B(n6662), .Z(n6663) );
  NANDN U14355 ( .A(y[915]), .B(x[915]), .Z(n13941) );
  AND U14356 ( .A(n6663), .B(n13941), .Z(n6664) );
  NANDN U14357 ( .A(n26119), .B(n6664), .Z(n6665) );
  NANDN U14358 ( .A(x[915]), .B(y[915]), .Z(n13942) );
  AND U14359 ( .A(n6665), .B(n13942), .Z(n6666) );
  NAND U14360 ( .A(n13939), .B(n6666), .Z(n6667) );
  NANDN U14361 ( .A(n13940), .B(n6667), .Z(n6668) );
  NANDN U14362 ( .A(y[917]), .B(x[917]), .Z(n13937) );
  NANDN U14363 ( .A(n6668), .B(n13937), .Z(n6669) );
  NAND U14364 ( .A(n6670), .B(n6669), .Z(n6671) );
  NANDN U14365 ( .A(n13936), .B(n6671), .Z(n6672) );
  ANDN U14366 ( .B(x[919]), .A(y[919]), .Z(n16597) );
  OR U14367 ( .A(n6672), .B(n16597), .Z(n6673) );
  AND U14368 ( .A(n6674), .B(n6673), .Z(n6678) );
  NANDN U14369 ( .A(y[920]), .B(x[920]), .Z(n26127) );
  NANDN U14370 ( .A(y[921]), .B(x[921]), .Z(n26128) );
  NAND U14371 ( .A(n26127), .B(n26128), .Z(n6676) );
  NAND U14372 ( .A(n6676), .B(n6675), .Z(n6677) );
  NANDN U14373 ( .A(n6678), .B(n6677), .Z(n6679) );
  NANDN U14374 ( .A(x[922]), .B(y[922]), .Z(n26129) );
  AND U14375 ( .A(n6679), .B(n26129), .Z(n6680) );
  NANDN U14376 ( .A(y[922]), .B(x[922]), .Z(n16602) );
  NANDN U14377 ( .A(y[923]), .B(x[923]), .Z(n16607) );
  NAND U14378 ( .A(n16602), .B(n16607), .Z(n26130) );
  OR U14379 ( .A(n6680), .B(n26130), .Z(n6681) );
  AND U14380 ( .A(n26131), .B(n6681), .Z(n6682) );
  NANDN U14381 ( .A(x[924]), .B(y[924]), .Z(n13930) );
  NAND U14382 ( .A(n6682), .B(n13930), .Z(n6683) );
  NAND U14383 ( .A(n26132), .B(n6683), .Z(n6684) );
  AND U14384 ( .A(n13931), .B(n6684), .Z(n6686) );
  NANDN U14385 ( .A(x[927]), .B(y[927]), .Z(n6690) );
  NANDN U14386 ( .A(x[926]), .B(y[926]), .Z(n6685) );
  AND U14387 ( .A(n6690), .B(n6685), .Z(n13933) );
  NAND U14388 ( .A(n6686), .B(n13933), .Z(n6691) );
  XNOR U14389 ( .A(x[927]), .B(y[927]), .Z(n6688) );
  NANDN U14390 ( .A(y[926]), .B(x[926]), .Z(n6687) );
  NAND U14391 ( .A(n6688), .B(n6687), .Z(n6689) );
  NAND U14392 ( .A(n6690), .B(n6689), .Z(n24490) );
  AND U14393 ( .A(n6691), .B(n24490), .Z(n6692) );
  ANDN U14394 ( .B(y[928]), .A(x[928]), .Z(n24489) );
  OR U14395 ( .A(n6692), .B(n24489), .Z(n6693) );
  NANDN U14396 ( .A(y[928]), .B(x[928]), .Z(n16611) );
  NANDN U14397 ( .A(y[929]), .B(x[929]), .Z(n16616) );
  AND U14398 ( .A(n16611), .B(n16616), .Z(n24488) );
  AND U14399 ( .A(n6693), .B(n24488), .Z(n6694) );
  ANDN U14400 ( .B(y[929]), .A(x[929]), .Z(n16613) );
  NANDN U14401 ( .A(x[930]), .B(y[930]), .Z(n16621) );
  NANDN U14402 ( .A(n16613), .B(n16621), .Z(n26135) );
  OR U14403 ( .A(n6694), .B(n26135), .Z(n6695) );
  NAND U14404 ( .A(n26136), .B(n6695), .Z(n6696) );
  NANDN U14405 ( .A(n26137), .B(n6696), .Z(n6697) );
  ANDN U14406 ( .B(y[932]), .A(x[932]), .Z(n13928) );
  OR U14407 ( .A(n6697), .B(n13928), .Z(n6698) );
  AND U14408 ( .A(n13927), .B(n6698), .Z(n6699) );
  NANDN U14409 ( .A(y[932]), .B(x[932]), .Z(n26138) );
  NAND U14410 ( .A(n6699), .B(n26138), .Z(n6700) );
  NANDN U14411 ( .A(x[934]), .B(y[934]), .Z(n13925) );
  AND U14412 ( .A(n6700), .B(n13925), .Z(n6701) );
  NAND U14413 ( .A(n13929), .B(n6701), .Z(n6702) );
  NANDN U14414 ( .A(y[935]), .B(x[935]), .Z(n26141) );
  AND U14415 ( .A(n6702), .B(n26141), .Z(n6703) );
  NAND U14416 ( .A(n13926), .B(n6703), .Z(n6704) );
  NANDN U14417 ( .A(n26142), .B(n6704), .Z(n6705) );
  ANDN U14418 ( .B(y[935]), .A(x[935]), .Z(n13924) );
  OR U14419 ( .A(n6705), .B(n13924), .Z(n6706) );
  AND U14420 ( .A(n26143), .B(n6706), .Z(n6709) );
  NANDN U14421 ( .A(x[938]), .B(y[938]), .Z(n6707) );
  NAND U14422 ( .A(n6708), .B(n6707), .Z(n16638) );
  ANDN U14423 ( .B(y[937]), .A(x[937]), .Z(n16633) );
  NOR U14424 ( .A(n16638), .B(n16633), .Z(n26144) );
  NANDN U14425 ( .A(n6709), .B(n26144), .Z(n6710) );
  NANDN U14426 ( .A(n26145), .B(n6710), .Z(n6713) );
  NANDN U14427 ( .A(x[940]), .B(y[940]), .Z(n6711) );
  AND U14428 ( .A(n6712), .B(n6711), .Z(n13921) );
  AND U14429 ( .A(n6713), .B(n13921), .Z(n6714) );
  OR U14430 ( .A(n6715), .B(n6714), .Z(n6716) );
  NAND U14431 ( .A(n13920), .B(n6716), .Z(n6717) );
  NANDN U14432 ( .A(n24486), .B(n6717), .Z(n6718) );
  NANDN U14433 ( .A(x[943]), .B(y[943]), .Z(n16647) );
  AND U14434 ( .A(n6718), .B(n16647), .Z(n6719) );
  NAND U14435 ( .A(n13917), .B(n6719), .Z(n6720) );
  NANDN U14436 ( .A(n13918), .B(n6720), .Z(n6721) );
  NANDN U14437 ( .A(y[945]), .B(x[945]), .Z(n13915) );
  NANDN U14438 ( .A(n6721), .B(n13915), .Z(n6722) );
  AND U14439 ( .A(n13916), .B(n6722), .Z(n6723) );
  NANDN U14440 ( .A(x[946]), .B(y[946]), .Z(n13913) );
  NAND U14441 ( .A(n6723), .B(n13913), .Z(n6724) );
  NANDN U14442 ( .A(y[947]), .B(x[947]), .Z(n13911) );
  AND U14443 ( .A(n6724), .B(n13911), .Z(n6725) );
  NANDN U14444 ( .A(n13914), .B(n6725), .Z(n6726) );
  NANDN U14445 ( .A(x[947]), .B(y[947]), .Z(n13912) );
  AND U14446 ( .A(n6726), .B(n13912), .Z(n6727) );
  NAND U14447 ( .A(n13909), .B(n6727), .Z(n6728) );
  NANDN U14448 ( .A(n13910), .B(n6728), .Z(n6729) );
  ANDN U14449 ( .B(x[949]), .A(y[949]), .Z(n13906) );
  OR U14450 ( .A(n6729), .B(n13906), .Z(n6730) );
  NAND U14451 ( .A(n6731), .B(n6730), .Z(n6732) );
  NANDN U14452 ( .A(y[950]), .B(x[950]), .Z(n13907) );
  AND U14453 ( .A(n6732), .B(n13907), .Z(n6733) );
  NAND U14454 ( .A(n13903), .B(n6733), .Z(n6734) );
  NAND U14455 ( .A(n13904), .B(n6734), .Z(n6735) );
  ANDN U14456 ( .B(y[952]), .A(x[952]), .Z(n13900) );
  OR U14457 ( .A(n6735), .B(n13900), .Z(n6736) );
  AND U14458 ( .A(n13902), .B(n6736), .Z(n6737) );
  NAND U14459 ( .A(n13899), .B(n6737), .Z(n6738) );
  AND U14460 ( .A(n13901), .B(n6738), .Z(n6739) );
  NANDN U14461 ( .A(x[954]), .B(y[954]), .Z(n13897) );
  NAND U14462 ( .A(n6739), .B(n13897), .Z(n6740) );
  NANDN U14463 ( .A(y[955]), .B(x[955]), .Z(n13895) );
  AND U14464 ( .A(n6740), .B(n13895), .Z(n6741) );
  NANDN U14465 ( .A(n13898), .B(n6741), .Z(n6742) );
  NANDN U14466 ( .A(x[955]), .B(y[955]), .Z(n13896) );
  AND U14467 ( .A(n6742), .B(n13896), .Z(n6743) );
  NAND U14468 ( .A(n16664), .B(n6743), .Z(n6744) );
  NAND U14469 ( .A(n26167), .B(n6744), .Z(n6745) );
  ANDN U14470 ( .B(x[956]), .A(y[956]), .Z(n13894) );
  OR U14471 ( .A(n6745), .B(n13894), .Z(n6746) );
  ANDN U14472 ( .B(y[958]), .A(x[958]), .Z(n26168) );
  ANDN U14473 ( .B(n6746), .A(n26168), .Z(n6747) );
  NANDN U14474 ( .A(x[957]), .B(y[957]), .Z(n16663) );
  NAND U14475 ( .A(n6747), .B(n16663), .Z(n6748) );
  NANDN U14476 ( .A(n26169), .B(n6748), .Z(n6749) );
  AND U14477 ( .A(n26171), .B(n6749), .Z(n6750) );
  OR U14478 ( .A(n26172), .B(n6750), .Z(n6751) );
  NAND U14479 ( .A(n26173), .B(n6751), .Z(n6752) );
  NANDN U14480 ( .A(n26174), .B(n6752), .Z(n6753) );
  ANDN U14481 ( .B(x[963]), .A(y[963]), .Z(n13892) );
  OR U14482 ( .A(n6753), .B(n13892), .Z(n6754) );
  AND U14483 ( .A(n26175), .B(n6754), .Z(n6755) );
  NANDN U14484 ( .A(x[964]), .B(y[964]), .Z(n13891) );
  NAND U14485 ( .A(n6755), .B(n13891), .Z(n6756) );
  ANDN U14486 ( .B(x[965]), .A(y[965]), .Z(n13888) );
  ANDN U14487 ( .B(n6756), .A(n13888), .Z(n6757) );
  NAND U14488 ( .A(n13893), .B(n6757), .Z(n6758) );
  NANDN U14489 ( .A(x[965]), .B(y[965]), .Z(n13890) );
  AND U14490 ( .A(n6758), .B(n13890), .Z(n6759) );
  NAND U14491 ( .A(n13887), .B(n6759), .Z(n6760) );
  NAND U14492 ( .A(n13889), .B(n6760), .Z(n6761) );
  ANDN U14493 ( .B(x[967]), .A(y[967]), .Z(n13884) );
  OR U14494 ( .A(n6761), .B(n13884), .Z(n6762) );
  NAND U14495 ( .A(n6763), .B(n6762), .Z(n6764) );
  NANDN U14496 ( .A(y[968]), .B(x[968]), .Z(n13885) );
  AND U14497 ( .A(n6764), .B(n13885), .Z(n6765) );
  NAND U14498 ( .A(n16693), .B(n6765), .Z(n6766) );
  NANDN U14499 ( .A(n13882), .B(n6766), .Z(n6767) );
  ANDN U14500 ( .B(y[970]), .A(x[970]), .Z(n16696) );
  OR U14501 ( .A(n6767), .B(n16696), .Z(n6768) );
  AND U14502 ( .A(n26183), .B(n6768), .Z(n6769) );
  NANDN U14503 ( .A(y[970]), .B(x[970]), .Z(n16692) );
  NAND U14504 ( .A(n6769), .B(n16692), .Z(n6770) );
  ANDN U14505 ( .B(y[971]), .A(x[971]), .Z(n16695) );
  ANDN U14506 ( .B(n6770), .A(n16695), .Z(n6771) );
  NAND U14507 ( .A(n26184), .B(n6771), .Z(n6772) );
  NAND U14508 ( .A(n26185), .B(n6772), .Z(n6773) );
  NAND U14509 ( .A(n26186), .B(n6773), .Z(n6774) );
  AND U14510 ( .A(n13879), .B(n6774), .Z(n6775) );
  NAND U14511 ( .A(n24484), .B(n6775), .Z(n6776) );
  ANDN U14512 ( .B(y[979]), .A(x[979]), .Z(n26187) );
  ANDN U14513 ( .B(n6776), .A(n26187), .Z(n6777) );
  NANDN U14514 ( .A(n13877), .B(n6777), .Z(n6778) );
  NANDN U14515 ( .A(y[980]), .B(x[980]), .Z(n13878) );
  AND U14516 ( .A(n6778), .B(n13878), .Z(n6779) );
  NAND U14517 ( .A(n13875), .B(n6779), .Z(n6780) );
  NANDN U14518 ( .A(n13876), .B(n6780), .Z(n6781) );
  ANDN U14519 ( .B(y[982]), .A(x[982]), .Z(n13872) );
  OR U14520 ( .A(n6781), .B(n13872), .Z(n6782) );
  NANDN U14521 ( .A(y[983]), .B(x[983]), .Z(n24483) );
  AND U14522 ( .A(n6782), .B(n24483), .Z(n6783) );
  NANDN U14523 ( .A(n6784), .B(n6783), .Z(n6785) );
  AND U14524 ( .A(n6786), .B(n6785), .Z(n6787) );
  OR U14525 ( .A(n26195), .B(n6787), .Z(n6788) );
  NAND U14526 ( .A(n26196), .B(n6788), .Z(n6789) );
  NANDN U14527 ( .A(n26197), .B(n6789), .Z(n6790) );
  NANDN U14528 ( .A(n24482), .B(n6790), .Z(n6791) );
  AND U14529 ( .A(n26198), .B(n6791), .Z(n6793) );
  NANDN U14530 ( .A(x[989]), .B(y[989]), .Z(n26199) );
  ANDN U14531 ( .B(y[990]), .A(x[990]), .Z(n13870) );
  ANDN U14532 ( .B(n26199), .A(n13870), .Z(n6792) );
  NANDN U14533 ( .A(n6793), .B(n6792), .Z(n6794) );
  NAND U14534 ( .A(n26200), .B(n6794), .Z(n6795) );
  NANDN U14535 ( .A(n13871), .B(n6795), .Z(n6796) );
  AND U14536 ( .A(n26202), .B(n6796), .Z(n6799) );
  NANDN U14537 ( .A(x[996]), .B(y[996]), .Z(n16756) );
  NANDN U14538 ( .A(x[994]), .B(y[994]), .Z(n6798) );
  NANDN U14539 ( .A(x[995]), .B(y[995]), .Z(n6797) );
  AND U14540 ( .A(n6798), .B(n6797), .Z(n16749) );
  NANDN U14541 ( .A(n6799), .B(n26204), .Z(n6800) );
  NANDN U14542 ( .A(n26205), .B(n6800), .Z(n6801) );
  NANDN U14543 ( .A(x[997]), .B(y[997]), .Z(n16755) );
  NANDN U14544 ( .A(x[998]), .B(y[998]), .Z(n16762) );
  AND U14545 ( .A(n16755), .B(n16762), .Z(n24481) );
  AND U14546 ( .A(n6801), .B(n24481), .Z(n6802) );
  ANDN U14547 ( .B(x[998]), .A(y[998]), .Z(n16758) );
  ANDN U14548 ( .B(x[999]), .A(y[999]), .Z(n16766) );
  OR U14549 ( .A(n16758), .B(n16766), .Z(n26206) );
  OR U14550 ( .A(n6802), .B(n26206), .Z(n6803) );
  NANDN U14551 ( .A(x[999]), .B(y[999]), .Z(n26207) );
  AND U14552 ( .A(n6803), .B(n26207), .Z(n6804) );
  NANDN U14553 ( .A(x[1000]), .B(y[1000]), .Z(n16769) );
  NAND U14554 ( .A(n6804), .B(n16769), .Z(n6805) );
  NANDN U14555 ( .A(y[1001]), .B(x[1001]), .Z(n16772) );
  AND U14556 ( .A(n6805), .B(n16772), .Z(n6806) );
  NANDN U14557 ( .A(n24480), .B(n6806), .Z(n6807) );
  NANDN U14558 ( .A(x[1001]), .B(y[1001]), .Z(n16768) );
  AND U14559 ( .A(n6807), .B(n16768), .Z(n6808) );
  NAND U14560 ( .A(n13868), .B(n6808), .Z(n6809) );
  NANDN U14561 ( .A(n16771), .B(n6809), .Z(n6810) );
  ANDN U14562 ( .B(x[1003]), .A(y[1003]), .Z(n13865) );
  OR U14563 ( .A(n6810), .B(n13865), .Z(n6811) );
  NAND U14564 ( .A(n6812), .B(n6811), .Z(n6813) );
  NANDN U14565 ( .A(y[1004]), .B(x[1004]), .Z(n13866) );
  AND U14566 ( .A(n6813), .B(n13866), .Z(n6814) );
  NAND U14567 ( .A(n13862), .B(n6814), .Z(n6815) );
  NAND U14568 ( .A(n13863), .B(n6815), .Z(n6816) );
  ANDN U14569 ( .B(y[1006]), .A(x[1006]), .Z(n13859) );
  OR U14570 ( .A(n6816), .B(n13859), .Z(n6817) );
  AND U14571 ( .A(n26214), .B(n6817), .Z(n6818) );
  NANDN U14572 ( .A(n13861), .B(n6818), .Z(n6819) );
  AND U14573 ( .A(n6820), .B(n6819), .Z(n6821) );
  OR U14574 ( .A(n26217), .B(n6821), .Z(n6822) );
  AND U14575 ( .A(n6823), .B(n6822), .Z(n6824) );
  NANDN U14576 ( .A(y[1010]), .B(x[1010]), .Z(n13858) );
  NANDN U14577 ( .A(y[1011]), .B(x[1011]), .Z(n16789) );
  NAND U14578 ( .A(n13858), .B(n16789), .Z(n24478) );
  OR U14579 ( .A(n6824), .B(n24478), .Z(n6825) );
  NANDN U14580 ( .A(x[1011]), .B(y[1011]), .Z(n24477) );
  AND U14581 ( .A(n6825), .B(n24477), .Z(n6826) );
  NANDN U14582 ( .A(x[1012]), .B(y[1012]), .Z(n13856) );
  NAND U14583 ( .A(n6826), .B(n13856), .Z(n6827) );
  NANDN U14584 ( .A(y[1013]), .B(x[1013]), .Z(n13854) );
  AND U14585 ( .A(n6827), .B(n13854), .Z(n6828) );
  NAND U14586 ( .A(n26220), .B(n6828), .Z(n6829) );
  NANDN U14587 ( .A(x[1013]), .B(y[1013]), .Z(n13855) );
  AND U14588 ( .A(n6829), .B(n13855), .Z(n6830) );
  NAND U14589 ( .A(n16794), .B(n6830), .Z(n6831) );
  NANDN U14590 ( .A(n13853), .B(n6831), .Z(n6832) );
  ANDN U14591 ( .B(x[1015]), .A(y[1015]), .Z(n13850) );
  OR U14592 ( .A(n6832), .B(n13850), .Z(n6833) );
  AND U14593 ( .A(n16793), .B(n6833), .Z(n6834) );
  NANDN U14594 ( .A(n13848), .B(n6834), .Z(n6835) );
  NAND U14595 ( .A(n13851), .B(n6835), .Z(n6836) );
  NANDN U14596 ( .A(n13847), .B(n6836), .Z(n6837) );
  NANDN U14597 ( .A(y[1018]), .B(x[1018]), .Z(n13852) );
  AND U14598 ( .A(n6837), .B(n13852), .Z(n6838) );
  NAND U14599 ( .A(n13845), .B(n6838), .Z(n6839) );
  NANDN U14600 ( .A(n13846), .B(n6839), .Z(n6840) );
  ANDN U14601 ( .B(y[1020]), .A(x[1020]), .Z(n13842) );
  OR U14602 ( .A(n6840), .B(n13842), .Z(n6841) );
  AND U14603 ( .A(n26226), .B(n6841), .Z(n6842) );
  NANDN U14604 ( .A(n13844), .B(n6842), .Z(n6843) );
  AND U14605 ( .A(n26227), .B(n6843), .Z(n6844) );
  NAND U14606 ( .A(n13843), .B(n6844), .Z(n6845) );
  NAND U14607 ( .A(n26228), .B(n6845), .Z(n6846) );
  NANDN U14608 ( .A(n26229), .B(n6846), .Z(n6847) );
  NAND U14609 ( .A(n26232), .B(n6847), .Z(n6848) );
  NANDN U14610 ( .A(n26233), .B(n6848), .Z(n6849) );
  AND U14611 ( .A(n26234), .B(n6849), .Z(n6852) );
  NANDN U14612 ( .A(x[1030]), .B(y[1030]), .Z(n6851) );
  AND U14613 ( .A(n6851), .B(n6850), .Z(n26235) );
  NANDN U14614 ( .A(n6852), .B(n26235), .Z(n6853) );
  NAND U14615 ( .A(n26236), .B(n6853), .Z(n6854) );
  NANDN U14616 ( .A(n26237), .B(n6854), .Z(n6855) );
  NAND U14617 ( .A(n26238), .B(n6855), .Z(n6856) );
  NANDN U14618 ( .A(n26239), .B(n6856), .Z(n6857) );
  AND U14619 ( .A(n26240), .B(n6857), .Z(n6861) );
  NANDN U14620 ( .A(x[1038]), .B(y[1038]), .Z(n6859) );
  NANDN U14621 ( .A(x[1037]), .B(y[1037]), .Z(n6858) );
  AND U14622 ( .A(n6859), .B(n6858), .Z(n6860) );
  NANDN U14623 ( .A(x[1039]), .B(y[1039]), .Z(n6865) );
  NAND U14624 ( .A(n6860), .B(n6865), .Z(n24474) );
  OR U14625 ( .A(n6861), .B(n24474), .Z(n6868) );
  XNOR U14626 ( .A(x[1039]), .B(y[1039]), .Z(n6863) );
  NANDN U14627 ( .A(y[1038]), .B(x[1038]), .Z(n6862) );
  NAND U14628 ( .A(n6863), .B(n6862), .Z(n6864) );
  NAND U14629 ( .A(n6865), .B(n6864), .Z(n6867) );
  NANDN U14630 ( .A(y[1040]), .B(x[1040]), .Z(n6866) );
  AND U14631 ( .A(n6867), .B(n6866), .Z(n24473) );
  AND U14632 ( .A(n6868), .B(n24473), .Z(n6871) );
  NANDN U14633 ( .A(x[1040]), .B(y[1040]), .Z(n6870) );
  NANDN U14634 ( .A(x[1041]), .B(y[1041]), .Z(n6869) );
  NAND U14635 ( .A(n6870), .B(n6869), .Z(n13841) );
  OR U14636 ( .A(n6871), .B(n13841), .Z(n6874) );
  NANDN U14637 ( .A(y[1042]), .B(x[1042]), .Z(n6873) );
  NANDN U14638 ( .A(y[1041]), .B(x[1041]), .Z(n6872) );
  AND U14639 ( .A(n6873), .B(n6872), .Z(n13840) );
  AND U14640 ( .A(n6874), .B(n13840), .Z(n6875) );
  NANDN U14641 ( .A(x[1042]), .B(y[1042]), .Z(n13839) );
  NANDN U14642 ( .A(n6875), .B(n13839), .Z(n6876) );
  NAND U14643 ( .A(n13837), .B(n6876), .Z(n6877) );
  NANDN U14644 ( .A(n13838), .B(n6877), .Z(n6878) );
  ANDN U14645 ( .B(y[1044]), .A(x[1044]), .Z(n13835) );
  OR U14646 ( .A(n6878), .B(n13835), .Z(n6879) );
  AND U14647 ( .A(n13836), .B(n6879), .Z(n6880) );
  NANDN U14648 ( .A(y[1045]), .B(x[1045]), .Z(n13833) );
  NAND U14649 ( .A(n6880), .B(n13833), .Z(n6881) );
  ANDN U14650 ( .B(y[1046]), .A(x[1046]), .Z(n13831) );
  ANDN U14651 ( .B(n6881), .A(n13831), .Z(n6882) );
  NANDN U14652 ( .A(n13834), .B(n6882), .Z(n6883) );
  NANDN U14653 ( .A(y[1047]), .B(x[1047]), .Z(n13829) );
  AND U14654 ( .A(n6883), .B(n13829), .Z(n6884) );
  NAND U14655 ( .A(n13832), .B(n6884), .Z(n6885) );
  NANDN U14656 ( .A(n26250), .B(n6885), .Z(n6886) );
  ANDN U14657 ( .B(y[1047]), .A(x[1047]), .Z(n13830) );
  OR U14658 ( .A(n6886), .B(n13830), .Z(n6887) );
  NANDN U14659 ( .A(y[1048]), .B(x[1048]), .Z(n16843) );
  NANDN U14660 ( .A(y[1049]), .B(x[1049]), .Z(n16847) );
  AND U14661 ( .A(n16843), .B(n16847), .Z(n26251) );
  AND U14662 ( .A(n6887), .B(n26251), .Z(n6889) );
  NANDN U14663 ( .A(x[1049]), .B(y[1049]), .Z(n26252) );
  ANDN U14664 ( .B(y[1050]), .A(x[1050]), .Z(n13827) );
  ANDN U14665 ( .B(n26252), .A(n13827), .Z(n6888) );
  NANDN U14666 ( .A(n6889), .B(n6888), .Z(n6890) );
  NANDN U14667 ( .A(n6891), .B(n6890), .Z(n6892) );
  NANDN U14668 ( .A(x[1051]), .B(y[1051]), .Z(n13828) );
  AND U14669 ( .A(n6892), .B(n13828), .Z(n6893) );
  NANDN U14670 ( .A(n26255), .B(n6893), .Z(n6894) );
  NANDN U14671 ( .A(n26256), .B(n6894), .Z(n6895) );
  NANDN U14672 ( .A(n26257), .B(n6895), .Z(n6896) );
  AND U14673 ( .A(n26258), .B(n6896), .Z(n6897) );
  NANDN U14674 ( .A(x[1055]), .B(y[1055]), .Z(n13823) );
  NANDN U14675 ( .A(x[1056]), .B(y[1056]), .Z(n16866) );
  NAND U14676 ( .A(n13823), .B(n16866), .Z(n24470) );
  OR U14677 ( .A(n6897), .B(n24470), .Z(n6898) );
  NAND U14678 ( .A(n26260), .B(n6898), .Z(n6899) );
  NANDN U14679 ( .A(n13822), .B(n6899), .Z(n6900) );
  NANDN U14680 ( .A(x[1058]), .B(y[1058]), .Z(n13821) );
  NANDN U14681 ( .A(n6900), .B(n13821), .Z(n6901) );
  NAND U14682 ( .A(n6902), .B(n6901), .Z(n6903) );
  NAND U14683 ( .A(n26265), .B(n6903), .Z(n6904) );
  ANDN U14684 ( .B(y[1059]), .A(x[1059]), .Z(n13820) );
  OR U14685 ( .A(n6904), .B(n13820), .Z(n6905) );
  AND U14686 ( .A(n26266), .B(n6905), .Z(n6906) );
  OR U14687 ( .A(n26267), .B(n6906), .Z(n6907) );
  NAND U14688 ( .A(n26268), .B(n6907), .Z(n6908) );
  NANDN U14689 ( .A(n13819), .B(n6908), .Z(n6909) );
  ANDN U14690 ( .B(y[1064]), .A(x[1064]), .Z(n13817) );
  OR U14691 ( .A(n6909), .B(n13817), .Z(n6910) );
  NAND U14692 ( .A(n26270), .B(n6910), .Z(n6911) );
  NANDN U14693 ( .A(n13818), .B(n6911), .Z(n6912) );
  NAND U14694 ( .A(n24469), .B(n6912), .Z(n6913) );
  ANDN U14695 ( .B(y[1068]), .A(x[1068]), .Z(n13814) );
  ANDN U14696 ( .B(n6913), .A(n13814), .Z(n6914) );
  NANDN U14697 ( .A(n24468), .B(n6914), .Z(n6915) );
  NAND U14698 ( .A(n26272), .B(n6915), .Z(n6916) );
  NANDN U14699 ( .A(n13815), .B(n6916), .Z(n6919) );
  NANDN U14700 ( .A(y[1071]), .B(x[1071]), .Z(n6918) );
  NANDN U14701 ( .A(y[1070]), .B(x[1070]), .Z(n6917) );
  AND U14702 ( .A(n6918), .B(n6917), .Z(n26274) );
  AND U14703 ( .A(n6919), .B(n26274), .Z(n6920) );
  NANDN U14704 ( .A(x[1071]), .B(y[1071]), .Z(n16898) );
  NANDN U14705 ( .A(x[1072]), .B(y[1072]), .Z(n16901) );
  NAND U14706 ( .A(n16898), .B(n16901), .Z(n24467) );
  OR U14707 ( .A(n6920), .B(n24467), .Z(n6921) );
  NAND U14708 ( .A(n26277), .B(n6921), .Z(n6922) );
  NANDN U14709 ( .A(n24466), .B(n6922), .Z(n6923) );
  NANDN U14710 ( .A(y[1074]), .B(x[1074]), .Z(n16907) );
  AND U14711 ( .A(n6923), .B(n16907), .Z(n6924) );
  NAND U14712 ( .A(n13811), .B(n6924), .Z(n6925) );
  NANDN U14713 ( .A(n13812), .B(n6925), .Z(n6926) );
  ANDN U14714 ( .B(y[1076]), .A(x[1076]), .Z(n13808) );
  OR U14715 ( .A(n6926), .B(n13808), .Z(n6927) );
  NAND U14716 ( .A(n6928), .B(n6927), .Z(n6929) );
  NANDN U14717 ( .A(x[1077]), .B(y[1077]), .Z(n13809) );
  AND U14718 ( .A(n6929), .B(n13809), .Z(n6930) );
  NAND U14719 ( .A(n13805), .B(n6930), .Z(n6931) );
  NAND U14720 ( .A(n13806), .B(n6931), .Z(n6934) );
  NANDN U14721 ( .A(y[1079]), .B(x[1079]), .Z(n6932) );
  NAND U14722 ( .A(n6933), .B(n6932), .Z(n24465) );
  OR U14723 ( .A(n6934), .B(n24465), .Z(n6935) );
  AND U14724 ( .A(n6936), .B(n6935), .Z(n6937) );
  NAND U14725 ( .A(n13802), .B(n6937), .Z(n6938) );
  NANDN U14726 ( .A(n13800), .B(n6938), .Z(n6939) );
  AND U14727 ( .A(n24463), .B(n6939), .Z(n6940) );
  OR U14728 ( .A(n26286), .B(n6940), .Z(n6941) );
  NAND U14729 ( .A(n26287), .B(n6941), .Z(n6942) );
  NANDN U14730 ( .A(n26288), .B(n6942), .Z(n6943) );
  NANDN U14731 ( .A(x[1088]), .B(y[1088]), .Z(n24462) );
  NANDN U14732 ( .A(x[1090]), .B(y[1090]), .Z(n13794) );
  NANDN U14733 ( .A(y[1092]), .B(x[1092]), .Z(n6945) );
  NANDN U14734 ( .A(y[1093]), .B(x[1093]), .Z(n6944) );
  NAND U14735 ( .A(n6945), .B(n6944), .Z(n13788) );
  NANDN U14736 ( .A(x[1093]), .B(y[1093]), .Z(n13792) );
  ANDN U14737 ( .B(y[1094]), .A(x[1094]), .Z(n13786) );
  NANDN U14738 ( .A(y[1095]), .B(x[1095]), .Z(n16944) );
  NANDN U14739 ( .A(y[1094]), .B(x[1094]), .Z(n13790) );
  XNOR U14740 ( .A(y[1103]), .B(x[1103]), .Z(n6947) );
  NANDN U14741 ( .A(x[1102]), .B(y[1102]), .Z(n6946) );
  NAND U14742 ( .A(n6947), .B(n6946), .Z(n6948) );
  NAND U14743 ( .A(n6949), .B(n6948), .Z(n6951) );
  NANDN U14744 ( .A(x[1104]), .B(y[1104]), .Z(n6950) );
  AND U14745 ( .A(n6951), .B(n6950), .Z(n24460) );
  NANDN U14746 ( .A(y[1104]), .B(x[1104]), .Z(n6953) );
  NANDN U14747 ( .A(y[1105]), .B(x[1105]), .Z(n6952) );
  NAND U14748 ( .A(n6953), .B(n6952), .Z(n26301) );
  NAND U14749 ( .A(n26302), .B(n6954), .Z(n6955) );
  NANDN U14750 ( .A(n26303), .B(n6955), .Z(n6956) );
  NAND U14751 ( .A(n26306), .B(n6956), .Z(n6957) );
  NANDN U14752 ( .A(n13778), .B(n6957), .Z(n6958) );
  AND U14753 ( .A(n13776), .B(n6958), .Z(n6960) );
  NANDN U14754 ( .A(y[1110]), .B(x[1110]), .Z(n13779) );
  ANDN U14755 ( .B(x[1111]), .A(y[1111]), .Z(n13774) );
  ANDN U14756 ( .B(n13779), .A(n13774), .Z(n6959) );
  NANDN U14757 ( .A(n6960), .B(n6959), .Z(n6961) );
  AND U14758 ( .A(n13777), .B(n6961), .Z(n6962) );
  NANDN U14759 ( .A(x[1112]), .B(y[1112]), .Z(n26309) );
  NAND U14760 ( .A(n6962), .B(n26309), .Z(n6963) );
  NANDN U14761 ( .A(n26310), .B(n6963), .Z(n6964) );
  AND U14762 ( .A(n26311), .B(n6964), .Z(n6965) );
  NANDN U14763 ( .A(x[1114]), .B(y[1114]), .Z(n16970) );
  NAND U14764 ( .A(n6965), .B(n16970), .Z(n6966) );
  NANDN U14765 ( .A(y[1115]), .B(x[1115]), .Z(n26314) );
  AND U14766 ( .A(n6966), .B(n26314), .Z(n6967) );
  NAND U14767 ( .A(n26312), .B(n6967), .Z(n6968) );
  NANDN U14768 ( .A(x[1116]), .B(y[1116]), .Z(n13771) );
  AND U14769 ( .A(n6968), .B(n13771), .Z(n6969) );
  NAND U14770 ( .A(n16969), .B(n6969), .Z(n6970) );
  NANDN U14771 ( .A(n26317), .B(n6970), .Z(n6971) );
  NANDN U14772 ( .A(x[1118]), .B(y[1118]), .Z(n13766) );
  AND U14773 ( .A(n6971), .B(n13766), .Z(n6972) );
  NAND U14774 ( .A(n26316), .B(n6972), .Z(n6973) );
  NANDN U14775 ( .A(n13769), .B(n6973), .Z(n6974) );
  NAND U14776 ( .A(n13765), .B(n6974), .Z(n6975) );
  NANDN U14777 ( .A(n13763), .B(n6975), .Z(n6976) );
  NANDN U14778 ( .A(x[1121]), .B(y[1121]), .Z(n13762) );
  AND U14779 ( .A(n6976), .B(n13762), .Z(n6977) );
  NANDN U14780 ( .A(x[1122]), .B(y[1122]), .Z(n13761) );
  NAND U14781 ( .A(n6977), .B(n13761), .Z(n6978) );
  ANDN U14782 ( .B(x[1123]), .A(y[1123]), .Z(n16980) );
  ANDN U14783 ( .B(n6978), .A(n16980), .Z(n6979) );
  NANDN U14784 ( .A(n13764), .B(n6979), .Z(n6980) );
  NANDN U14785 ( .A(x[1123]), .B(y[1123]), .Z(n13760) );
  AND U14786 ( .A(n6980), .B(n13760), .Z(n6981) );
  NAND U14787 ( .A(n16986), .B(n6981), .Z(n6982) );
  NANDN U14788 ( .A(n26325), .B(n6982), .Z(n6983) );
  NANDN U14789 ( .A(n26326), .B(n6983), .Z(n6984) );
  AND U14790 ( .A(n16994), .B(n6984), .Z(n6985) );
  NAND U14791 ( .A(n26327), .B(n6985), .Z(n6986) );
  ANDN U14792 ( .B(y[1128]), .A(x[1128]), .Z(n16997) );
  ANDN U14793 ( .B(n6986), .A(n16997), .Z(n6987) );
  NANDN U14794 ( .A(n24458), .B(n6987), .Z(n6988) );
  NANDN U14795 ( .A(y[1129]), .B(x[1129]), .Z(n24456) );
  AND U14796 ( .A(n6988), .B(n24456), .Z(n6989) );
  NAND U14797 ( .A(n16993), .B(n6989), .Z(n6990) );
  NANDN U14798 ( .A(n26329), .B(n6990), .Z(n6991) );
  ANDN U14799 ( .B(y[1129]), .A(x[1129]), .Z(n16996) );
  OR U14800 ( .A(n6991), .B(n16996), .Z(n6992) );
  NANDN U14801 ( .A(y[1130]), .B(x[1130]), .Z(n17000) );
  NANDN U14802 ( .A(y[1131]), .B(x[1131]), .Z(n17005) );
  AND U14803 ( .A(n17000), .B(n17005), .Z(n26330) );
  AND U14804 ( .A(n6992), .B(n26330), .Z(n6993) );
  ANDN U14805 ( .B(y[1131]), .A(x[1131]), .Z(n17002) );
  ANDN U14806 ( .B(y[1132]), .A(x[1132]), .Z(n17010) );
  OR U14807 ( .A(n17002), .B(n17010), .Z(n24455) );
  OR U14808 ( .A(n6993), .B(n24455), .Z(n6994) );
  NANDN U14809 ( .A(y[1132]), .B(x[1132]), .Z(n17006) );
  NANDN U14810 ( .A(y[1133]), .B(x[1133]), .Z(n13758) );
  AND U14811 ( .A(n17006), .B(n13758), .Z(n24454) );
  AND U14812 ( .A(n6994), .B(n24454), .Z(n6996) );
  ANDN U14813 ( .B(y[1134]), .A(x[1134]), .Z(n17016) );
  IV U14814 ( .A(n17016), .Z(n26335) );
  ANDN U14815 ( .B(y[1133]), .A(x[1133]), .Z(n26333) );
  ANDN U14816 ( .B(n26335), .A(n26333), .Z(n6995) );
  NANDN U14817 ( .A(n6996), .B(n6995), .Z(n6997) );
  NANDN U14818 ( .A(n6998), .B(n6997), .Z(n6999) );
  NAND U14819 ( .A(n26336), .B(n6999), .Z(n7000) );
  ANDN U14820 ( .B(x[1137]), .A(y[1137]), .Z(n13755) );
  ANDN U14821 ( .B(n7000), .A(n13755), .Z(n7002) );
  NANDN U14822 ( .A(y[1136]), .B(x[1136]), .Z(n13757) );
  ANDN U14823 ( .B(n7001), .A(n13757), .Z(n24451) );
  ANDN U14824 ( .B(n7002), .A(n24451), .Z(n7003) );
  ANDN U14825 ( .B(y[1138]), .A(x[1138]), .Z(n13753) );
  OR U14826 ( .A(n7003), .B(n13753), .Z(n7004) );
  AND U14827 ( .A(n13756), .B(n7004), .Z(n7005) );
  NANDN U14828 ( .A(y[1139]), .B(x[1139]), .Z(n13752) );
  NAND U14829 ( .A(n7005), .B(n13752), .Z(n7006) );
  ANDN U14830 ( .B(y[1140]), .A(x[1140]), .Z(n13749) );
  ANDN U14831 ( .B(n7006), .A(n13749), .Z(n7007) );
  NAND U14832 ( .A(n13754), .B(n7007), .Z(n7008) );
  NANDN U14833 ( .A(y[1140]), .B(x[1140]), .Z(n13751) );
  AND U14834 ( .A(n7008), .B(n13751), .Z(n7009) );
  NAND U14835 ( .A(n17027), .B(n7009), .Z(n7010) );
  NAND U14836 ( .A(n13750), .B(n7010), .Z(n7011) );
  ANDN U14837 ( .B(y[1142]), .A(x[1142]), .Z(n17029) );
  OR U14838 ( .A(n7011), .B(n17029), .Z(n7012) );
  NAND U14839 ( .A(n7013), .B(n7012), .Z(n7014) );
  NANDN U14840 ( .A(x[1144]), .B(y[1144]), .Z(n13744) );
  AND U14841 ( .A(n7014), .B(n13744), .Z(n7015) );
  NAND U14842 ( .A(n17030), .B(n7015), .Z(n7016) );
  NAND U14843 ( .A(n13748), .B(n7016), .Z(n7018) );
  NANDN U14844 ( .A(x[1146]), .B(y[1146]), .Z(n13743) );
  NANDN U14845 ( .A(x[1145]), .B(y[1145]), .Z(n13745) );
  AND U14846 ( .A(n13743), .B(n13745), .Z(n7017) );
  NAND U14847 ( .A(n7018), .B(n7017), .Z(n7020) );
  NANDN U14848 ( .A(y[1147]), .B(x[1147]), .Z(n13742) );
  NANDN U14849 ( .A(y[1146]), .B(x[1146]), .Z(n7019) );
  AND U14850 ( .A(n13742), .B(n7019), .Z(n24448) );
  AND U14851 ( .A(n7020), .B(n24448), .Z(n7021) );
  ANDN U14852 ( .B(y[1147]), .A(x[1147]), .Z(n17037) );
  NANDN U14853 ( .A(x[1148]), .B(y[1148]), .Z(n17043) );
  NANDN U14854 ( .A(n17037), .B(n17043), .Z(n26343) );
  OR U14855 ( .A(n7021), .B(n26343), .Z(n7022) );
  NAND U14856 ( .A(n26345), .B(n7022), .Z(n7023) );
  NANDN U14857 ( .A(n26346), .B(n7023), .Z(n7025) );
  NANDN U14858 ( .A(y[1151]), .B(x[1151]), .Z(n13741) );
  NANDN U14859 ( .A(y[1150]), .B(x[1150]), .Z(n17046) );
  AND U14860 ( .A(n13741), .B(n17046), .Z(n7024) );
  NAND U14861 ( .A(n7025), .B(n7024), .Z(n7026) );
  ANDN U14862 ( .B(y[1151]), .A(x[1151]), .Z(n26348) );
  ANDN U14863 ( .B(n7026), .A(n26348), .Z(n7027) );
  NANDN U14864 ( .A(x[1152]), .B(y[1152]), .Z(n13739) );
  NAND U14865 ( .A(n7027), .B(n13739), .Z(n7028) );
  NANDN U14866 ( .A(y[1153]), .B(x[1153]), .Z(n26350) );
  AND U14867 ( .A(n7028), .B(n26350), .Z(n7029) );
  NANDN U14868 ( .A(n13740), .B(n7029), .Z(n7030) );
  NANDN U14869 ( .A(x[1153]), .B(y[1153]), .Z(n13738) );
  AND U14870 ( .A(n7030), .B(n13738), .Z(n7031) );
  NANDN U14871 ( .A(n26351), .B(n7031), .Z(n7032) );
  NANDN U14872 ( .A(n26352), .B(n7032), .Z(n7033) );
  NAND U14873 ( .A(n26353), .B(n7033), .Z(n7034) );
  NAND U14874 ( .A(n26354), .B(n7034), .Z(n7035) );
  NANDN U14875 ( .A(n13735), .B(n7035), .Z(n7036) );
  NANDN U14876 ( .A(y[1159]), .B(x[1159]), .Z(n17067) );
  AND U14877 ( .A(n7036), .B(n17067), .Z(n7037) );
  NAND U14878 ( .A(n26355), .B(n7037), .Z(n7038) );
  NANDN U14879 ( .A(n13733), .B(n7038), .Z(n7039) );
  ANDN U14880 ( .B(y[1159]), .A(x[1159]), .Z(n13734) );
  OR U14881 ( .A(n7039), .B(n13734), .Z(n7040) );
  AND U14882 ( .A(n26361), .B(n7040), .Z(n7041) );
  NANDN U14883 ( .A(x[1161]), .B(y[1161]), .Z(n17072) );
  NANDN U14884 ( .A(x[1162]), .B(y[1162]), .Z(n17079) );
  NAND U14885 ( .A(n17072), .B(n17079), .Z(n26362) );
  OR U14886 ( .A(n7041), .B(n26362), .Z(n7042) );
  AND U14887 ( .A(n26363), .B(n7042), .Z(n7044) );
  NANDN U14888 ( .A(x[1163]), .B(y[1163]), .Z(n26364) );
  ANDN U14889 ( .B(y[1164]), .A(x[1164]), .Z(n13730) );
  ANDN U14890 ( .B(n26364), .A(n13730), .Z(n7043) );
  NANDN U14891 ( .A(n7044), .B(n7043), .Z(n7045) );
  NANDN U14892 ( .A(n26365), .B(n7045), .Z(n7046) );
  NAND U14893 ( .A(n13732), .B(n7046), .Z(n7047) );
  NANDN U14894 ( .A(n17085), .B(n7047), .Z(n7048) );
  NANDN U14895 ( .A(x[1167]), .B(y[1167]), .Z(n17087) );
  AND U14896 ( .A(n7048), .B(n17087), .Z(n7049) );
  NANDN U14897 ( .A(x[1168]), .B(y[1168]), .Z(n13727) );
  NAND U14898 ( .A(n7049), .B(n13727), .Z(n7050) );
  NANDN U14899 ( .A(y[1169]), .B(x[1169]), .Z(n13725) );
  AND U14900 ( .A(n7050), .B(n13725), .Z(n7051) );
  NANDN U14901 ( .A(n13728), .B(n7051), .Z(n7052) );
  NANDN U14902 ( .A(x[1169]), .B(y[1169]), .Z(n13726) );
  AND U14903 ( .A(n7052), .B(n13726), .Z(n7053) );
  NAND U14904 ( .A(n13723), .B(n7053), .Z(n7054) );
  NANDN U14905 ( .A(n13724), .B(n7054), .Z(n7055) );
  ANDN U14906 ( .B(x[1171]), .A(y[1171]), .Z(n13720) );
  OR U14907 ( .A(n7055), .B(n13720), .Z(n7056) );
  NAND U14908 ( .A(n7057), .B(n7056), .Z(n7058) );
  NANDN U14909 ( .A(y[1172]), .B(x[1172]), .Z(n13721) );
  AND U14910 ( .A(n7058), .B(n13721), .Z(n7059) );
  NAND U14911 ( .A(n13717), .B(n7059), .Z(n7060) );
  NAND U14912 ( .A(n13718), .B(n7060), .Z(n7061) );
  ANDN U14913 ( .B(y[1174]), .A(x[1174]), .Z(n13715) );
  OR U14914 ( .A(n7061), .B(n13715), .Z(n7062) );
  NANDN U14915 ( .A(y[1175]), .B(x[1175]), .Z(n26377) );
  AND U14916 ( .A(n7062), .B(n26377), .Z(n7063) );
  NANDN U14917 ( .A(y[1174]), .B(x[1174]), .Z(n13716) );
  NAND U14918 ( .A(n7063), .B(n13716), .Z(n7066) );
  NANDN U14919 ( .A(x[1176]), .B(y[1176]), .Z(n7065) );
  ANDN U14920 ( .B(n7065), .A(n7064), .Z(n26378) );
  AND U14921 ( .A(n7066), .B(n26378), .Z(n7067) );
  NANDN U14922 ( .A(n13714), .B(n7067), .Z(n7068) );
  NAND U14923 ( .A(n26379), .B(n7068), .Z(n7069) );
  NANDN U14924 ( .A(n24445), .B(n7069), .Z(n7070) );
  AND U14925 ( .A(n26380), .B(n7070), .Z(n7071) );
  OR U14926 ( .A(n26381), .B(n7071), .Z(n7072) );
  NAND U14927 ( .A(n26382), .B(n7072), .Z(n7073) );
  NAND U14928 ( .A(n26383), .B(n7073), .Z(n7074) );
  ANDN U14929 ( .B(y[1184]), .A(x[1184]), .Z(n13710) );
  OR U14930 ( .A(n7074), .B(n13710), .Z(n7075) );
  NAND U14931 ( .A(n26384), .B(n7075), .Z(n7076) );
  NANDN U14932 ( .A(n13711), .B(n7076), .Z(n7077) );
  NAND U14933 ( .A(n13708), .B(n7077), .Z(n7078) );
  NAND U14934 ( .A(n26387), .B(n7078), .Z(n7079) );
  NANDN U14935 ( .A(n26388), .B(n7079), .Z(n7080) );
  NAND U14936 ( .A(n13707), .B(n7080), .Z(n7081) );
  ANDN U14937 ( .B(y[1190]), .A(x[1190]), .Z(n13704) );
  OR U14938 ( .A(n7081), .B(n13704), .Z(n7082) );
  NAND U14939 ( .A(n26390), .B(n7082), .Z(n7083) );
  NANDN U14940 ( .A(n13706), .B(n7083), .Z(n7084) );
  NAND U14941 ( .A(n24444), .B(n7084), .Z(n7085) );
  NANDN U14942 ( .A(n26394), .B(n7085), .Z(n7086) );
  NANDN U14943 ( .A(y[1195]), .B(x[1195]), .Z(n13703) );
  AND U14944 ( .A(n7086), .B(n13703), .Z(n7087) );
  ANDN U14945 ( .B(y[1196]), .A(x[1196]), .Z(n24443) );
  OR U14946 ( .A(n7087), .B(n24443), .Z(n7088) );
  NAND U14947 ( .A(n24442), .B(n7088), .Z(n7089) );
  NANDN U14948 ( .A(n13701), .B(n7089), .Z(n7090) );
  ANDN U14949 ( .B(y[1197]), .A(x[1197]), .Z(n13702) );
  OR U14950 ( .A(n7090), .B(n13702), .Z(n7091) );
  NAND U14951 ( .A(n26398), .B(n7091), .Z(n7092) );
  NANDN U14952 ( .A(n13699), .B(n7092), .Z(n7093) );
  ANDN U14953 ( .B(y[1199]), .A(x[1199]), .Z(n13700) );
  OR U14954 ( .A(n7093), .B(n13700), .Z(n7094) );
  NAND U14955 ( .A(n26399), .B(n7094), .Z(n7095) );
  NANDN U14956 ( .A(n24438), .B(n7095), .Z(n7096) );
  NANDN U14957 ( .A(y[1202]), .B(x[1202]), .Z(n13698) );
  AND U14958 ( .A(n7096), .B(n13698), .Z(n7097) );
  NAND U14959 ( .A(n13697), .B(n7097), .Z(n7098) );
  NANDN U14960 ( .A(n17157), .B(n7098), .Z(n7099) );
  ANDN U14961 ( .B(y[1204]), .A(x[1204]), .Z(n13694) );
  OR U14962 ( .A(n7099), .B(n13694), .Z(n7100) );
  NAND U14963 ( .A(n7101), .B(n7100), .Z(n7102) );
  AND U14964 ( .A(n13693), .B(n7102), .Z(n7103) );
  NAND U14965 ( .A(n13695), .B(n7103), .Z(n7104) );
  NANDN U14966 ( .A(n26408), .B(n7104), .Z(n7105) );
  OR U14967 ( .A(n7106), .B(n7105), .Z(n7107) );
  AND U14968 ( .A(n17164), .B(n7107), .Z(n7108) );
  NANDN U14969 ( .A(x[1208]), .B(y[1208]), .Z(n26409) );
  NAND U14970 ( .A(n7108), .B(n26409), .Z(n7109) );
  NANDN U14971 ( .A(n26412), .B(n7109), .Z(n7110) );
  AND U14972 ( .A(n26414), .B(n7110), .Z(n7111) );
  OR U14973 ( .A(n26416), .B(n7111), .Z(n7112) );
  NAND U14974 ( .A(n26418), .B(n7112), .Z(n7113) );
  NANDN U14975 ( .A(n26420), .B(n7113), .Z(n7114) );
  NAND U14976 ( .A(n26422), .B(n7114), .Z(n7115) );
  NAND U14977 ( .A(n17192), .B(n7115), .Z(n7116) );
  NANDN U14978 ( .A(n17194), .B(n7116), .Z(n7117) );
  NAND U14979 ( .A(n17196), .B(n7117), .Z(n7118) );
  NANDN U14980 ( .A(x[1218]), .B(y[1218]), .Z(n13690) );
  AND U14981 ( .A(n7118), .B(n13690), .Z(n7119) );
  NAND U14982 ( .A(n26430), .B(n7119), .Z(n7120) );
  NAND U14983 ( .A(n7121), .B(n7120), .Z(n7122) );
  NANDN U14984 ( .A(x[1220]), .B(y[1220]), .Z(n26437) );
  AND U14985 ( .A(n7122), .B(n26437), .Z(n7123) );
  NANDN U14986 ( .A(n13689), .B(n7123), .Z(n7124) );
  AND U14987 ( .A(n26440), .B(n7124), .Z(n7126) );
  NANDN U14988 ( .A(x[1221]), .B(y[1221]), .Z(n26442) );
  ANDN U14989 ( .B(y[1222]), .A(x[1222]), .Z(n13685) );
  ANDN U14990 ( .B(n26442), .A(n13685), .Z(n7125) );
  NANDN U14991 ( .A(n7126), .B(n7125), .Z(n7127) );
  NANDN U14992 ( .A(n7128), .B(n7127), .Z(n7131) );
  NANDN U14993 ( .A(x[1224]), .B(y[1224]), .Z(n7129) );
  NAND U14994 ( .A(n7130), .B(n7129), .Z(n26448) );
  ANDN U14995 ( .B(n7131), .A(n26448), .Z(n7132) );
  NAND U14996 ( .A(n13686), .B(n7132), .Z(n7133) );
  NANDN U14997 ( .A(n26449), .B(n7133), .Z(n7134) );
  AND U14998 ( .A(n26450), .B(n7134), .Z(n7135) );
  NANDN U14999 ( .A(y[1228]), .B(x[1228]), .Z(n17216) );
  NANDN U15000 ( .A(y[1229]), .B(x[1229]), .Z(n17223) );
  NAND U15001 ( .A(n17216), .B(n17223), .Z(n24437) );
  OR U15002 ( .A(n7135), .B(n24437), .Z(n7136) );
  NAND U15003 ( .A(n26451), .B(n7136), .Z(n7137) );
  NANDN U15004 ( .A(n26452), .B(n7137), .Z(n7138) );
  XOR U15005 ( .A(x[1232]), .B(y[1232]), .Z(n13682) );
  ANDN U15006 ( .B(n7138), .A(n13682), .Z(n7139) );
  NAND U15007 ( .A(n26454), .B(n7139), .Z(n7140) );
  NANDN U15008 ( .A(n26455), .B(n7140), .Z(n7141) );
  NAND U15009 ( .A(n26456), .B(n7141), .Z(n7142) );
  ANDN U15010 ( .B(x[1235]), .A(y[1235]), .Z(n13679) );
  ANDN U15011 ( .B(n7142), .A(n13679), .Z(n7143) );
  NANDN U15012 ( .A(n26457), .B(n7143), .Z(n7144) );
  NANDN U15013 ( .A(x[1235]), .B(y[1235]), .Z(n26458) );
  AND U15014 ( .A(n7144), .B(n26458), .Z(n7145) );
  NAND U15015 ( .A(n13678), .B(n7145), .Z(n7146) );
  NAND U15016 ( .A(n13680), .B(n7146), .Z(n7147) );
  ANDN U15017 ( .B(x[1237]), .A(y[1237]), .Z(n13676) );
  OR U15018 ( .A(n7147), .B(n13676), .Z(n7148) );
  NAND U15019 ( .A(n7149), .B(n7148), .Z(n7150) );
  NANDN U15020 ( .A(n13675), .B(n7150), .Z(n7151) );
  ANDN U15021 ( .B(x[1239]), .A(y[1239]), .Z(n24436) );
  OR U15022 ( .A(n7151), .B(n24436), .Z(n7152) );
  AND U15023 ( .A(n7153), .B(n7152), .Z(n7154) );
  NANDN U15024 ( .A(y[1240]), .B(x[1240]), .Z(n17245) );
  NANDN U15025 ( .A(y[1241]), .B(x[1241]), .Z(n17250) );
  NAND U15026 ( .A(n17245), .B(n17250), .Z(n26465) );
  OR U15027 ( .A(n7154), .B(n26465), .Z(n7155) );
  NANDN U15028 ( .A(x[1241]), .B(y[1241]), .Z(n26466) );
  AND U15029 ( .A(n7155), .B(n26466), .Z(n7156) );
  NANDN U15030 ( .A(x[1242]), .B(y[1242]), .Z(n13671) );
  NAND U15031 ( .A(n7156), .B(n13671), .Z(n7157) );
  ANDN U15032 ( .B(x[1243]), .A(y[1243]), .Z(n17254) );
  ANDN U15033 ( .B(n7157), .A(n17254), .Z(n7158) );
  NANDN U15034 ( .A(n17249), .B(n7158), .Z(n7159) );
  NANDN U15035 ( .A(x[1243]), .B(y[1243]), .Z(n13670) );
  AND U15036 ( .A(n7159), .B(n13670), .Z(n7160) );
  NANDN U15037 ( .A(n26470), .B(n7160), .Z(n7161) );
  NANDN U15038 ( .A(n26471), .B(n7161), .Z(n7163) );
  NANDN U15039 ( .A(x[1246]), .B(y[1246]), .Z(n17263) );
  ANDN U15040 ( .B(y[1245]), .A(x[1245]), .Z(n26472) );
  ANDN U15041 ( .B(n17263), .A(n26472), .Z(n7162) );
  NAND U15042 ( .A(n7163), .B(n7162), .Z(n7164) );
  AND U15043 ( .A(n7165), .B(n7164), .Z(n7169) );
  NANDN U15044 ( .A(x[1248]), .B(y[1248]), .Z(n7167) );
  ANDN U15045 ( .B(n7167), .A(n7166), .Z(n26476) );
  ANDN U15046 ( .B(y[1247]), .A(x[1247]), .Z(n17262) );
  ANDN U15047 ( .B(n26476), .A(n17262), .Z(n7168) );
  NANDN U15048 ( .A(n7169), .B(n7168), .Z(n7170) );
  AND U15049 ( .A(n26477), .B(n7170), .Z(n7179) );
  ANDN U15050 ( .B(y[1250]), .A(x[1250]), .Z(n7171) );
  NAND U15051 ( .A(n7171), .B(y[1251]), .Z(n7174) );
  XOR U15052 ( .A(n7171), .B(y[1251]), .Z(n7172) );
  NANDN U15053 ( .A(x[1251]), .B(n7172), .Z(n7173) );
  NAND U15054 ( .A(n7174), .B(n7173), .Z(n7176) );
  NOR U15055 ( .A(n7176), .B(n7175), .Z(n7178) );
  NANDN U15056 ( .A(x[1252]), .B(y[1252]), .Z(n7177) );
  NAND U15057 ( .A(n7178), .B(n7177), .Z(n24435) );
  OR U15058 ( .A(n7179), .B(n24435), .Z(n7180) );
  AND U15059 ( .A(n7181), .B(n7180), .Z(n7183) );
  NANDN U15060 ( .A(x[1256]), .B(y[1256]), .Z(n13665) );
  ANDN U15061 ( .B(y[1255]), .A(x[1255]), .Z(n24433) );
  ANDN U15062 ( .B(n13665), .A(n24433), .Z(n7182) );
  NANDN U15063 ( .A(n7183), .B(n7182), .Z(n7184) );
  NANDN U15064 ( .A(y[1257]), .B(x[1257]), .Z(n13664) );
  AND U15065 ( .A(n7184), .B(n13664), .Z(n7185) );
  NANDN U15066 ( .A(y[1256]), .B(x[1256]), .Z(n13667) );
  NAND U15067 ( .A(n7185), .B(n13667), .Z(n7186) );
  NANDN U15068 ( .A(x[1257]), .B(y[1257]), .Z(n13666) );
  AND U15069 ( .A(n7186), .B(n13666), .Z(n7187) );
  NANDN U15070 ( .A(n26482), .B(n7187), .Z(n7188) );
  NANDN U15071 ( .A(n26483), .B(n7188), .Z(n7189) );
  NANDN U15072 ( .A(x[1260]), .B(y[1260]), .Z(n13663) );
  AND U15073 ( .A(n7189), .B(n13663), .Z(n7190) );
  NAND U15074 ( .A(n26484), .B(n7190), .Z(n7191) );
  NAND U15075 ( .A(n26485), .B(n7191), .Z(n7193) );
  NANDN U15076 ( .A(x[1261]), .B(y[1261]), .Z(n13662) );
  ANDN U15077 ( .B(y[1262]), .A(x[1262]), .Z(n24431) );
  ANDN U15078 ( .B(n13662), .A(n24431), .Z(n7192) );
  NAND U15079 ( .A(n7193), .B(n7192), .Z(n7194) );
  AND U15080 ( .A(n26486), .B(n7194), .Z(n7195) );
  ANDN U15081 ( .B(y[1263]), .A(x[1263]), .Z(n17290) );
  NANDN U15082 ( .A(x[1264]), .B(y[1264]), .Z(n17294) );
  NANDN U15083 ( .A(n17290), .B(n17294), .Z(n24428) );
  OR U15084 ( .A(n7195), .B(n24428), .Z(n7196) );
  NAND U15085 ( .A(n26488), .B(n7196), .Z(n7197) );
  NANDN U15086 ( .A(n24427), .B(n7197), .Z(n7198) );
  NANDN U15087 ( .A(y[1266]), .B(x[1266]), .Z(n17300) );
  AND U15088 ( .A(n7198), .B(n17300), .Z(n7199) );
  NAND U15089 ( .A(n13658), .B(n7199), .Z(n7200) );
  NANDN U15090 ( .A(n13659), .B(n7200), .Z(n7201) );
  NANDN U15091 ( .A(x[1268]), .B(y[1268]), .Z(n13656) );
  NANDN U15092 ( .A(n7201), .B(n13656), .Z(n7202) );
  AND U15093 ( .A(n13657), .B(n7202), .Z(n7203) );
  NAND U15094 ( .A(n17307), .B(n7203), .Z(n7206) );
  ANDN U15095 ( .B(y[1269]), .A(x[1269]), .Z(n13655) );
  NAND U15096 ( .A(n13655), .B(n7204), .Z(n7205) );
  NAND U15097 ( .A(n7206), .B(n7205), .Z(n7209) );
  NANDN U15098 ( .A(x[1270]), .B(y[1270]), .Z(n7208) );
  NANDN U15099 ( .A(x[1271]), .B(y[1271]), .Z(n7207) );
  NAND U15100 ( .A(n7208), .B(n7207), .Z(n17309) );
  OR U15101 ( .A(n7209), .B(n17309), .Z(n7210) );
  NAND U15102 ( .A(n24426), .B(n7210), .Z(n7211) );
  NANDN U15103 ( .A(n17314), .B(n7211), .Z(n7215) );
  NANDN U15104 ( .A(y[1274]), .B(x[1274]), .Z(n17319) );
  NANDN U15105 ( .A(y[1273]), .B(x[1273]), .Z(n17316) );
  NANDN U15106 ( .A(y[1272]), .B(x[1272]), .Z(n17311) );
  NAND U15107 ( .A(n17316), .B(n17311), .Z(n7212) );
  NAND U15108 ( .A(n7213), .B(n7212), .Z(n7214) );
  AND U15109 ( .A(n17319), .B(n7214), .Z(n26496) );
  AND U15110 ( .A(n7215), .B(n26496), .Z(n7216) );
  NAND U15111 ( .A(n13653), .B(n7216), .Z(n7217) );
  NANDN U15112 ( .A(n13654), .B(n7217), .Z(n7218) );
  ANDN U15113 ( .B(y[1276]), .A(x[1276]), .Z(n13650) );
  OR U15114 ( .A(n7218), .B(n13650), .Z(n7219) );
  AND U15115 ( .A(n13652), .B(n7219), .Z(n7220) );
  NANDN U15116 ( .A(n26500), .B(n7220), .Z(n7221) );
  AND U15117 ( .A(n7222), .B(n7221), .Z(n7223) );
  OR U15118 ( .A(n26502), .B(n7223), .Z(n7224) );
  NAND U15119 ( .A(n26504), .B(n7224), .Z(n7225) );
  NANDN U15120 ( .A(n26505), .B(n7225), .Z(n7226) );
  NAND U15121 ( .A(n26506), .B(n7226), .Z(n7227) );
  NANDN U15122 ( .A(n24425), .B(n7227), .Z(n7228) );
  AND U15123 ( .A(n26507), .B(n7228), .Z(n7229) );
  ANDN U15124 ( .B(x[1284]), .A(y[1284]), .Z(n17348) );
  NANDN U15125 ( .A(y[1285]), .B(x[1285]), .Z(n17354) );
  NANDN U15126 ( .A(n17348), .B(n17354), .Z(n24424) );
  OR U15127 ( .A(n7229), .B(n24424), .Z(n7230) );
  AND U15128 ( .A(n13647), .B(n7230), .Z(n7231) );
  NAND U15129 ( .A(n13648), .B(n7231), .Z(n7232) );
  NANDN U15130 ( .A(n26509), .B(n7232), .Z(n7235) );
  NANDN U15131 ( .A(x[1288]), .B(y[1288]), .Z(n7234) );
  NANDN U15132 ( .A(x[1287]), .B(y[1287]), .Z(n7233) );
  AND U15133 ( .A(n7234), .B(n7233), .Z(n13644) );
  AND U15134 ( .A(n7235), .B(n13644), .Z(n7238) );
  NANDN U15135 ( .A(y[1289]), .B(x[1289]), .Z(n7237) );
  NANDN U15136 ( .A(y[1288]), .B(x[1288]), .Z(n7236) );
  NAND U15137 ( .A(n7237), .B(n7236), .Z(n13642) );
  OR U15138 ( .A(n7238), .B(n13642), .Z(n7239) );
  NANDN U15139 ( .A(x[1289]), .B(y[1289]), .Z(n13641) );
  AND U15140 ( .A(n7239), .B(n13641), .Z(n7240) );
  NANDN U15141 ( .A(x[1290]), .B(y[1290]), .Z(n13640) );
  NAND U15142 ( .A(n7240), .B(n13640), .Z(n7241) );
  NANDN U15143 ( .A(y[1291]), .B(x[1291]), .Z(n13638) );
  AND U15144 ( .A(n7241), .B(n13638), .Z(n7242) );
  NANDN U15145 ( .A(n13643), .B(n7242), .Z(n7243) );
  NANDN U15146 ( .A(x[1291]), .B(y[1291]), .Z(n13639) );
  AND U15147 ( .A(n7243), .B(n13639), .Z(n7244) );
  NAND U15148 ( .A(n13636), .B(n7244), .Z(n7245) );
  NANDN U15149 ( .A(n13637), .B(n7245), .Z(n7247) );
  NANDN U15150 ( .A(y[1294]), .B(x[1294]), .Z(n7249) );
  NANDN U15151 ( .A(y[1293]), .B(x[1293]), .Z(n7246) );
  AND U15152 ( .A(n7249), .B(n7246), .Z(n24423) );
  NANDN U15153 ( .A(n7247), .B(n24423), .Z(n7251) );
  ANDN U15154 ( .B(y[1294]), .A(x[1294]), .Z(n17364) );
  NANDN U15155 ( .A(x[1293]), .B(y[1293]), .Z(n13635) );
  NANDN U15156 ( .A(n17364), .B(n13635), .Z(n7248) );
  AND U15157 ( .A(n7249), .B(n7248), .Z(n7250) );
  ANDN U15158 ( .B(n7251), .A(n7250), .Z(n7252) );
  NANDN U15159 ( .A(y[1295]), .B(x[1295]), .Z(n26516) );
  NANDN U15160 ( .A(n7252), .B(n26516), .Z(n7253) );
  NANDN U15161 ( .A(x[1298]), .B(y[1298]), .Z(n26520) );
  NANDN U15162 ( .A(x[1297]), .B(y[1297]), .Z(n13633) );
  AND U15163 ( .A(n26520), .B(n13633), .Z(n7256) );
  AND U15164 ( .A(n7253), .B(n7256), .Z(n7254) );
  ANDN U15165 ( .B(y[1295]), .A(x[1295]), .Z(n17363) );
  ANDN U15166 ( .B(n7254), .A(n17363), .Z(n7255) );
  XNOR U15167 ( .A(x[1296]), .B(y[1296]), .Z(n13634) );
  NAND U15168 ( .A(n7255), .B(n13634), .Z(n7257) );
  NANDN U15169 ( .A(y[1298]), .B(x[1298]), .Z(n13631) );
  NANDN U15170 ( .A(y[1297]), .B(x[1297]), .Z(n13630) );
  AND U15171 ( .A(n7257), .B(n24422), .Z(n7258) );
  NAND U15172 ( .A(n13628), .B(n7258), .Z(n7259) );
  NANDN U15173 ( .A(n13629), .B(n7259), .Z(n7260) );
  ANDN U15174 ( .B(y[1300]), .A(x[1300]), .Z(n13625) );
  OR U15175 ( .A(n7260), .B(n13625), .Z(n7261) );
  AND U15176 ( .A(n13627), .B(n7261), .Z(n7262) );
  NANDN U15177 ( .A(y[1301]), .B(x[1301]), .Z(n13624) );
  NAND U15178 ( .A(n7262), .B(n13624), .Z(n7263) );
  AND U15179 ( .A(n13626), .B(n7263), .Z(n7264) );
  NANDN U15180 ( .A(x[1302]), .B(y[1302]), .Z(n13622) );
  NAND U15181 ( .A(n7264), .B(n13622), .Z(n7265) );
  ANDN U15182 ( .B(x[1303]), .A(y[1303]), .Z(n17377) );
  ANDN U15183 ( .B(n7265), .A(n17377), .Z(n7266) );
  NANDN U15184 ( .A(n13623), .B(n7266), .Z(n7269) );
  NANDN U15185 ( .A(x[1304]), .B(y[1304]), .Z(n7267) );
  AND U15186 ( .A(n7268), .B(n7267), .Z(n26527) );
  AND U15187 ( .A(n7269), .B(n26527), .Z(n7270) );
  NAND U15188 ( .A(n13621), .B(n7270), .Z(n7271) );
  NANDN U15189 ( .A(n24421), .B(n7271), .Z(n7272) );
  NAND U15190 ( .A(n24420), .B(n7272), .Z(n7273) );
  NANDN U15191 ( .A(n13620), .B(n7273), .Z(n7274) );
  NANDN U15192 ( .A(x[1308]), .B(y[1308]), .Z(n13619) );
  AND U15193 ( .A(n7274), .B(n13619), .Z(n7275) );
  NANDN U15194 ( .A(y[1308]), .B(x[1308]), .Z(n17386) );
  NANDN U15195 ( .A(y[1309]), .B(x[1309]), .Z(n13618) );
  NAND U15196 ( .A(n17386), .B(n13618), .Z(n26530) );
  OR U15197 ( .A(n7275), .B(n26530), .Z(n7276) );
  NANDN U15198 ( .A(x[1309]), .B(y[1309]), .Z(n17389) );
  AND U15199 ( .A(n7276), .B(n17389), .Z(n7277) );
  NANDN U15200 ( .A(n13616), .B(n7277), .Z(n7278) );
  AND U15201 ( .A(n7279), .B(n7278), .Z(n7281) );
  NANDN U15202 ( .A(x[1311]), .B(y[1311]), .Z(n13617) );
  ANDN U15203 ( .B(y[1312]), .A(x[1312]), .Z(n24419) );
  ANDN U15204 ( .B(n13617), .A(n24419), .Z(n7280) );
  NANDN U15205 ( .A(n7281), .B(n7280), .Z(n7282) );
  NANDN U15206 ( .A(y[1312]), .B(x[1312]), .Z(n17394) );
  NANDN U15207 ( .A(y[1313]), .B(x[1313]), .Z(n13615) );
  AND U15208 ( .A(n17394), .B(n13615), .Z(n24418) );
  AND U15209 ( .A(n7282), .B(n24418), .Z(n7283) );
  ANDN U15210 ( .B(y[1313]), .A(x[1313]), .Z(n17398) );
  ANDN U15211 ( .B(y[1314]), .A(x[1314]), .Z(n17404) );
  OR U15212 ( .A(n17398), .B(n17404), .Z(n24417) );
  OR U15213 ( .A(n7283), .B(n24417), .Z(n7284) );
  NAND U15214 ( .A(n26536), .B(n7284), .Z(n7285) );
  NANDN U15215 ( .A(n26537), .B(n7285), .Z(n7286) );
  NANDN U15216 ( .A(x[1316]), .B(y[1316]), .Z(n13612) );
  NANDN U15217 ( .A(n7286), .B(n13612), .Z(n7287) );
  NAND U15218 ( .A(n26538), .B(n7287), .Z(n7288) );
  NANDN U15219 ( .A(n13611), .B(n7288), .Z(n7289) );
  ANDN U15220 ( .B(y[1318]), .A(x[1318]), .Z(n13613) );
  OR U15221 ( .A(n7289), .B(n13613), .Z(n7290) );
  NANDN U15222 ( .A(n26540), .B(n7290), .Z(n7291) );
  AND U15223 ( .A(n26541), .B(n7291), .Z(n7292) );
  OR U15224 ( .A(n26542), .B(n7292), .Z(n7293) );
  NAND U15225 ( .A(n26543), .B(n7293), .Z(n7294) );
  NANDN U15226 ( .A(n26544), .B(n7294), .Z(n7295) );
  NANDN U15227 ( .A(x[1324]), .B(y[1324]), .Z(n13608) );
  AND U15228 ( .A(n7295), .B(n13608), .Z(n7296) );
  NANDN U15229 ( .A(n26545), .B(n7296), .Z(n7297) );
  NANDN U15230 ( .A(n7298), .B(n7297), .Z(n7299) );
  AND U15231 ( .A(n26548), .B(n7299), .Z(n7300) );
  NAND U15232 ( .A(n13607), .B(n7300), .Z(n7301) );
  NANDN U15233 ( .A(n24414), .B(n7301), .Z(n7302) );
  NAND U15234 ( .A(n26549), .B(n7302), .Z(n7303) );
  NAND U15235 ( .A(n26550), .B(n7303), .Z(n7304) );
  NANDN U15236 ( .A(n13606), .B(n7304), .Z(n7305) );
  NANDN U15237 ( .A(x[1331]), .B(n7305), .Z(n7308) );
  XNOR U15238 ( .A(x[1331]), .B(n7305), .Z(n7306) );
  NAND U15239 ( .A(n7306), .B(y[1331]), .Z(n7307) );
  NAND U15240 ( .A(n7308), .B(n7307), .Z(n7309) );
  AND U15241 ( .A(n13605), .B(n7309), .Z(n7312) );
  NANDN U15242 ( .A(x[1332]), .B(y[1332]), .Z(n7311) );
  NANDN U15243 ( .A(x[1333]), .B(y[1333]), .Z(n7310) );
  NAND U15244 ( .A(n7311), .B(n7310), .Z(n26553) );
  OR U15245 ( .A(n7312), .B(n26553), .Z(n7315) );
  NANDN U15246 ( .A(y[1334]), .B(x[1334]), .Z(n7314) );
  NANDN U15247 ( .A(y[1333]), .B(x[1333]), .Z(n7313) );
  AND U15248 ( .A(n7314), .B(n7313), .Z(n26554) );
  AND U15249 ( .A(n7315), .B(n26554), .Z(n7318) );
  NANDN U15250 ( .A(x[1334]), .B(y[1334]), .Z(n7317) );
  NANDN U15251 ( .A(x[1335]), .B(y[1335]), .Z(n7316) );
  NAND U15252 ( .A(n7317), .B(n7316), .Z(n17440) );
  OR U15253 ( .A(n7318), .B(n17440), .Z(n7319) );
  NAND U15254 ( .A(n13603), .B(n7319), .Z(n7320) );
  NANDN U15255 ( .A(n17443), .B(n7320), .Z(n7321) );
  NAND U15256 ( .A(n26559), .B(n7321), .Z(n7322) );
  NAND U15257 ( .A(n26560), .B(n7322), .Z(n7323) );
  NANDN U15258 ( .A(n26561), .B(n7323), .Z(n7324) );
  AND U15259 ( .A(n26562), .B(n7324), .Z(n7325) );
  OR U15260 ( .A(n26563), .B(n7325), .Z(n7326) );
  NAND U15261 ( .A(n26564), .B(n7326), .Z(n7327) );
  NANDN U15262 ( .A(n24413), .B(n7327), .Z(n7328) );
  NANDN U15263 ( .A(x[1346]), .B(y[1346]), .Z(n26565) );
  NAND U15264 ( .A(n7328), .B(n26565), .Z(n7329) );
  NANDN U15265 ( .A(n26566), .B(n7329), .Z(n7330) );
  AND U15266 ( .A(n26567), .B(n7330), .Z(n7331) );
  OR U15267 ( .A(n26568), .B(n7331), .Z(n7332) );
  NAND U15268 ( .A(n26569), .B(n7332), .Z(n7333) );
  NANDN U15269 ( .A(n24412), .B(n7333), .Z(n7334) );
  NAND U15270 ( .A(n26570), .B(n7334), .Z(n7335) );
  NAND U15271 ( .A(n26571), .B(n7335), .Z(n7336) );
  NANDN U15272 ( .A(x[1354]), .B(y[1354]), .Z(n13594) );
  AND U15273 ( .A(n7336), .B(n13594), .Z(n7337) );
  NAND U15274 ( .A(n13597), .B(n7337), .Z(n7338) );
  NANDN U15275 ( .A(n26573), .B(n7338), .Z(n7339) );
  NANDN U15276 ( .A(x[1356]), .B(y[1356]), .Z(n13591) );
  AND U15277 ( .A(n7339), .B(n13591), .Z(n7340) );
  NAND U15278 ( .A(n13593), .B(n7340), .Z(n7341) );
  NANDN U15279 ( .A(n26578), .B(n7341), .Z(n7342) );
  NANDN U15280 ( .A(x[1358]), .B(y[1358]), .Z(n13590) );
  AND U15281 ( .A(n7342), .B(n13590), .Z(n7343) );
  NAND U15282 ( .A(n26577), .B(n7343), .Z(n7344) );
  NANDN U15283 ( .A(n7345), .B(n7344), .Z(n7347) );
  NANDN U15284 ( .A(x[1359]), .B(y[1359]), .Z(n13589) );
  NANDN U15285 ( .A(x[1360]), .B(y[1360]), .Z(n17511) );
  AND U15286 ( .A(n13589), .B(n17511), .Z(n7346) );
  NAND U15287 ( .A(n7347), .B(n7346), .Z(n7348) );
  AND U15288 ( .A(n26583), .B(n7348), .Z(n7349) );
  ANDN U15289 ( .B(y[1361]), .A(x[1361]), .Z(n17510) );
  ANDN U15290 ( .B(y[1362]), .A(x[1362]), .Z(n17517) );
  OR U15291 ( .A(n17510), .B(n17517), .Z(n26584) );
  OR U15292 ( .A(n7349), .B(n26584), .Z(n7350) );
  NANDN U15293 ( .A(y[1362]), .B(x[1362]), .Z(n24409) );
  AND U15294 ( .A(n7350), .B(n24409), .Z(n7351) );
  NANDN U15295 ( .A(y[1363]), .B(x[1363]), .Z(n17519) );
  NAND U15296 ( .A(n7351), .B(n17519), .Z(n7352) );
  ANDN U15297 ( .B(y[1364]), .A(x[1364]), .Z(n17522) );
  ANDN U15298 ( .B(n7352), .A(n17522), .Z(n7353) );
  NANDN U15299 ( .A(n26585), .B(n7353), .Z(n7354) );
  NANDN U15300 ( .A(y[1364]), .B(x[1364]), .Z(n17518) );
  AND U15301 ( .A(n7354), .B(n17518), .Z(n7355) );
  NAND U15302 ( .A(n13587), .B(n7355), .Z(n7356) );
  NANDN U15303 ( .A(n17521), .B(n7356), .Z(n7357) );
  ANDN U15304 ( .B(y[1366]), .A(x[1366]), .Z(n13584) );
  OR U15305 ( .A(n7357), .B(n13584), .Z(n7358) );
  NAND U15306 ( .A(n7359), .B(n7358), .Z(n7360) );
  NANDN U15307 ( .A(x[1367]), .B(y[1367]), .Z(n13585) );
  AND U15308 ( .A(n7360), .B(n13585), .Z(n7361) );
  NANDN U15309 ( .A(n26592), .B(n7361), .Z(n7362) );
  NANDN U15310 ( .A(n26593), .B(n7362), .Z(n7363) );
  NANDN U15311 ( .A(n24408), .B(n7363), .Z(n7364) );
  AND U15312 ( .A(n26594), .B(n7364), .Z(n7366) );
  NANDN U15313 ( .A(x[1372]), .B(y[1372]), .Z(n13581) );
  ANDN U15314 ( .B(y[1371]), .A(x[1371]), .Z(n17534) );
  ANDN U15315 ( .B(n13581), .A(n17534), .Z(n7365) );
  NANDN U15316 ( .A(n7366), .B(n7365), .Z(n7367) );
  NANDN U15317 ( .A(y[1373]), .B(x[1373]), .Z(n26598) );
  AND U15318 ( .A(n7367), .B(n26598), .Z(n7368) );
  NAND U15319 ( .A(n17540), .B(n7368), .Z(n7369) );
  NAND U15320 ( .A(n17543), .B(n7369), .Z(n7370) );
  ANDN U15321 ( .B(y[1373]), .A(x[1373]), .Z(n13580) );
  OR U15322 ( .A(n7370), .B(n13580), .Z(n7371) );
  AND U15323 ( .A(n13577), .B(n7371), .Z(n7372) );
  NANDN U15324 ( .A(y[1374]), .B(x[1374]), .Z(n26601) );
  NAND U15325 ( .A(n7372), .B(n26601), .Z(n7373) );
  NANDN U15326 ( .A(n7374), .B(n7373), .Z(n7375) );
  AND U15327 ( .A(n13578), .B(n7375), .Z(n7378) );
  NANDN U15328 ( .A(x[1378]), .B(y[1378]), .Z(n7377) );
  NANDN U15329 ( .A(x[1377]), .B(y[1377]), .Z(n7376) );
  NAND U15330 ( .A(n7377), .B(n7376), .Z(n13574) );
  OR U15331 ( .A(n7378), .B(n13574), .Z(n7381) );
  NANDN U15332 ( .A(y[1378]), .B(x[1378]), .Z(n7380) );
  NANDN U15333 ( .A(y[1379]), .B(x[1379]), .Z(n7379) );
  AND U15334 ( .A(n7380), .B(n7379), .Z(n17551) );
  AND U15335 ( .A(n7381), .B(n17551), .Z(n7382) );
  NANDN U15336 ( .A(x[1379]), .B(y[1379]), .Z(n17552) );
  NANDN U15337 ( .A(n7382), .B(n17552), .Z(n7383) );
  ANDN U15338 ( .B(y[1380]), .A(x[1380]), .Z(n13573) );
  OR U15339 ( .A(n7383), .B(n13573), .Z(n7384) );
  AND U15340 ( .A(n26608), .B(n7384), .Z(n7387) );
  NANDN U15341 ( .A(x[1382]), .B(y[1382]), .Z(n7386) );
  NANDN U15342 ( .A(x[1381]), .B(y[1381]), .Z(n7385) );
  AND U15343 ( .A(n7386), .B(n7385), .Z(n26611) );
  NANDN U15344 ( .A(n7387), .B(n26611), .Z(n7388) );
  NANDN U15345 ( .A(n26613), .B(n7388), .Z(n7389) );
  AND U15346 ( .A(n26614), .B(n7389), .Z(n7390) );
  OR U15347 ( .A(n26617), .B(n7390), .Z(n7391) );
  AND U15348 ( .A(n26619), .B(n7391), .Z(n7392) );
  OR U15349 ( .A(n26621), .B(n7392), .Z(n7393) );
  NAND U15350 ( .A(n26623), .B(n7393), .Z(n7394) );
  NANDN U15351 ( .A(n26625), .B(n7394), .Z(n7395) );
  NANDN U15352 ( .A(n26627), .B(n7395), .Z(n7396) );
  AND U15353 ( .A(n26629), .B(n7396), .Z(n7398) );
  NANDN U15354 ( .A(x[1389]), .B(y[1389]), .Z(n26630) );
  ANDN U15355 ( .B(y[1390]), .A(x[1390]), .Z(n13566) );
  ANDN U15356 ( .B(n26630), .A(n13566), .Z(n7397) );
  NANDN U15357 ( .A(n7398), .B(n7397), .Z(n7399) );
  NANDN U15358 ( .A(n26637), .B(n7399), .Z(n7400) );
  ANDN U15359 ( .B(x[1390]), .A(y[1390]), .Z(n13568) );
  OR U15360 ( .A(n7400), .B(n13568), .Z(n7401) );
  AND U15361 ( .A(n7402), .B(n7401), .Z(n7403) );
  OR U15362 ( .A(n26641), .B(n7403), .Z(n7404) );
  NAND U15363 ( .A(n26643), .B(n7404), .Z(n7405) );
  NANDN U15364 ( .A(n26645), .B(n7405), .Z(n7406) );
  ANDN U15365 ( .B(x[1395]), .A(y[1395]), .Z(n13564) );
  OR U15366 ( .A(n7406), .B(n13564), .Z(n7407) );
  AND U15367 ( .A(n13563), .B(n7407), .Z(n7408) );
  NANDN U15368 ( .A(x[1395]), .B(y[1395]), .Z(n26646) );
  NAND U15369 ( .A(n7408), .B(n26646), .Z(n7409) );
  ANDN U15370 ( .B(x[1397]), .A(y[1397]), .Z(n13560) );
  ANDN U15371 ( .B(n7409), .A(n13560), .Z(n7410) );
  NAND U15372 ( .A(n13565), .B(n7410), .Z(n7411) );
  AND U15373 ( .A(n13561), .B(n7411), .Z(n7412) );
  NAND U15374 ( .A(n13562), .B(n7412), .Z(n7413) );
  NANDN U15375 ( .A(n7414), .B(n7413), .Z(n7415) );
  OR U15376 ( .A(n26651), .B(n7415), .Z(n7416) );
  AND U15377 ( .A(n26652), .B(n7416), .Z(n7417) );
  NANDN U15378 ( .A(x[1399]), .B(y[1399]), .Z(n13558) );
  NAND U15379 ( .A(n7417), .B(n13558), .Z(n7418) );
  NANDN U15380 ( .A(n26653), .B(n7418), .Z(n7419) );
  AND U15381 ( .A(n26654), .B(n7419), .Z(n7421) );
  NANDN U15382 ( .A(y[1402]), .B(x[1402]), .Z(n7420) );
  ANDN U15383 ( .B(x[1403]), .A(y[1403]), .Z(n13556) );
  ANDN U15384 ( .B(n7420), .A(n13556), .Z(n26655) );
  NANDN U15385 ( .A(n7421), .B(n26655), .Z(n7422) );
  NAND U15386 ( .A(n26656), .B(n7422), .Z(n7423) );
  NANDN U15387 ( .A(n26657), .B(n7423), .Z(n7424) );
  NANDN U15388 ( .A(x[1406]), .B(y[1406]), .Z(n13554) );
  AND U15389 ( .A(n7424), .B(n13554), .Z(n7425) );
  NANDN U15390 ( .A(n26658), .B(n7425), .Z(n7426) );
  NANDN U15391 ( .A(n7427), .B(n7426), .Z(n7428) );
  NANDN U15392 ( .A(x[1407]), .B(y[1407]), .Z(n13553) );
  AND U15393 ( .A(n7428), .B(n13553), .Z(n7429) );
  NAND U15394 ( .A(n13552), .B(n7429), .Z(n7430) );
  NANDN U15395 ( .A(n24407), .B(n7430), .Z(n7431) );
  NANDN U15396 ( .A(x[1410]), .B(y[1410]), .Z(n13550) );
  AND U15397 ( .A(n7431), .B(n13550), .Z(n7432) );
  NAND U15398 ( .A(n17613), .B(n7432), .Z(n7433) );
  NANDN U15399 ( .A(n7434), .B(n7433), .Z(n7435) );
  NANDN U15400 ( .A(x[1412]), .B(y[1412]), .Z(n26668) );
  AND U15401 ( .A(n7435), .B(n26668), .Z(n7436) );
  NAND U15402 ( .A(n13549), .B(n7436), .Z(n7437) );
  NANDN U15403 ( .A(n24406), .B(n7437), .Z(n7439) );
  NANDN U15404 ( .A(x[1414]), .B(y[1414]), .Z(n13548) );
  NANDN U15405 ( .A(x[1413]), .B(y[1413]), .Z(n24405) );
  AND U15406 ( .A(n13548), .B(n24405), .Z(n7438) );
  NAND U15407 ( .A(n7439), .B(n7438), .Z(n7440) );
  AND U15408 ( .A(n7441), .B(n7440), .Z(n7443) );
  ANDN U15409 ( .B(y[1415]), .A(x[1415]), .Z(n13547) );
  ANDN U15410 ( .B(y[1416]), .A(x[1416]), .Z(n26672) );
  NOR U15411 ( .A(n13547), .B(n26672), .Z(n7442) );
  NANDN U15412 ( .A(n7443), .B(n7442), .Z(n7444) );
  AND U15413 ( .A(n26673), .B(n7444), .Z(n7445) );
  OR U15414 ( .A(n26674), .B(n7445), .Z(n7446) );
  NAND U15415 ( .A(n26675), .B(n7446), .Z(n7447) );
  NANDN U15416 ( .A(n26678), .B(n7447), .Z(n7448) );
  ANDN U15417 ( .B(y[1419]), .A(x[1419]), .Z(n26676) );
  OR U15418 ( .A(n7448), .B(n26676), .Z(n7449) );
  NAND U15419 ( .A(n7450), .B(n7449), .Z(n7451) );
  NANDN U15420 ( .A(n26681), .B(n7451), .Z(n7452) );
  NAND U15421 ( .A(n26682), .B(n7452), .Z(n7453) );
  NAND U15422 ( .A(n24404), .B(n7453), .Z(n7454) );
  NANDN U15423 ( .A(n26683), .B(n7454), .Z(n7455) );
  NAND U15424 ( .A(n17662), .B(n7455), .Z(n7456) );
  NANDN U15425 ( .A(x[1427]), .B(n7456), .Z(n7459) );
  XNOR U15426 ( .A(x[1427]), .B(n7456), .Z(n7457) );
  NAND U15427 ( .A(n7457), .B(y[1427]), .Z(n7458) );
  NAND U15428 ( .A(n7459), .B(n7458), .Z(n7460) );
  AND U15429 ( .A(n17665), .B(n7460), .Z(n7463) );
  NANDN U15430 ( .A(x[1428]), .B(y[1428]), .Z(n7462) );
  NANDN U15431 ( .A(x[1429]), .B(y[1429]), .Z(n7461) );
  AND U15432 ( .A(n7462), .B(n7461), .Z(n26686) );
  NANDN U15433 ( .A(n7463), .B(n26686), .Z(n7466) );
  NANDN U15434 ( .A(y[1430]), .B(x[1430]), .Z(n7465) );
  NANDN U15435 ( .A(y[1429]), .B(x[1429]), .Z(n7464) );
  NAND U15436 ( .A(n7465), .B(n7464), .Z(n26687) );
  ANDN U15437 ( .B(n7466), .A(n26687), .Z(n7469) );
  NANDN U15438 ( .A(x[1430]), .B(y[1430]), .Z(n7468) );
  NANDN U15439 ( .A(x[1431]), .B(y[1431]), .Z(n7467) );
  AND U15440 ( .A(n7468), .B(n7467), .Z(n26688) );
  NANDN U15441 ( .A(n7469), .B(n26688), .Z(n7470) );
  NANDN U15442 ( .A(n26689), .B(n7470), .Z(n7471) );
  NAND U15443 ( .A(n26690), .B(n7471), .Z(n7472) );
  ANDN U15444 ( .B(y[1434]), .A(x[1434]), .Z(n13545) );
  OR U15445 ( .A(n7472), .B(n13545), .Z(n7474) );
  NANDN U15446 ( .A(y[1434]), .B(x[1434]), .Z(n7473) );
  NANDN U15447 ( .A(y[1435]), .B(x[1435]), .Z(n13544) );
  AND U15448 ( .A(n7473), .B(n13544), .Z(n26691) );
  AND U15449 ( .A(n7474), .B(n26691), .Z(n7478) );
  NANDN U15450 ( .A(x[1436]), .B(y[1436]), .Z(n7476) );
  NANDN U15451 ( .A(x[1435]), .B(y[1435]), .Z(n7475) );
  AND U15452 ( .A(n7476), .B(n7475), .Z(n7477) );
  NANDN U15453 ( .A(x[1437]), .B(y[1437]), .Z(n7482) );
  NAND U15454 ( .A(n7477), .B(n7482), .Z(n13546) );
  OR U15455 ( .A(n7478), .B(n13546), .Z(n7485) );
  XNOR U15456 ( .A(x[1437]), .B(y[1437]), .Z(n7480) );
  NANDN U15457 ( .A(y[1436]), .B(x[1436]), .Z(n7479) );
  NAND U15458 ( .A(n7480), .B(n7479), .Z(n7481) );
  NAND U15459 ( .A(n7482), .B(n7481), .Z(n7484) );
  NANDN U15460 ( .A(y[1438]), .B(x[1438]), .Z(n7483) );
  NAND U15461 ( .A(n7484), .B(n7483), .Z(n26693) );
  ANDN U15462 ( .B(n7485), .A(n26693), .Z(n7488) );
  NANDN U15463 ( .A(x[1438]), .B(y[1438]), .Z(n7487) );
  NANDN U15464 ( .A(x[1439]), .B(y[1439]), .Z(n7486) );
  AND U15465 ( .A(n7487), .B(n7486), .Z(n26694) );
  NANDN U15466 ( .A(n7488), .B(n26694), .Z(n7491) );
  NANDN U15467 ( .A(y[1440]), .B(x[1440]), .Z(n7490) );
  NANDN U15468 ( .A(y[1439]), .B(x[1439]), .Z(n7489) );
  NAND U15469 ( .A(n7490), .B(n7489), .Z(n26696) );
  ANDN U15470 ( .B(n7491), .A(n26696), .Z(n7492) );
  ANDN U15471 ( .B(y[1440]), .A(x[1440]), .Z(n13542) );
  OR U15472 ( .A(n7492), .B(n13542), .Z(n7495) );
  NANDN U15473 ( .A(y[1441]), .B(x[1441]), .Z(n7493) );
  NAND U15474 ( .A(n7494), .B(n7493), .Z(n26698) );
  ANDN U15475 ( .B(n7495), .A(n26698), .Z(n7496) );
  OR U15476 ( .A(n7497), .B(n7496), .Z(n7498) );
  NAND U15477 ( .A(n26700), .B(n7498), .Z(n7499) );
  NANDN U15478 ( .A(n26701), .B(n7499), .Z(n7500) );
  AND U15479 ( .A(n26702), .B(n7500), .Z(n7502) );
  NANDN U15480 ( .A(x[1447]), .B(y[1447]), .Z(n26703) );
  ANDN U15481 ( .B(y[1448]), .A(x[1448]), .Z(n13536) );
  ANDN U15482 ( .B(n26703), .A(n13536), .Z(n7501) );
  NANDN U15483 ( .A(n7502), .B(n7501), .Z(n7503) );
  NANDN U15484 ( .A(n26704), .B(n7503), .Z(n7504) );
  AND U15485 ( .A(n13538), .B(n7504), .Z(n7505) );
  OR U15486 ( .A(n26706), .B(n7505), .Z(n7506) );
  NAND U15487 ( .A(n26707), .B(n7506), .Z(n7507) );
  NANDN U15488 ( .A(n26708), .B(n7507), .Z(n7508) );
  AND U15489 ( .A(n26709), .B(n7508), .Z(n7509) );
  OR U15490 ( .A(n26710), .B(n7509), .Z(n7510) );
  NAND U15491 ( .A(n26711), .B(n7510), .Z(n7511) );
  NANDN U15492 ( .A(n26712), .B(n7511), .Z(n7512) );
  NAND U15493 ( .A(n26713), .B(n7512), .Z(n7513) );
  ANDN U15494 ( .B(x[1459]), .A(y[1459]), .Z(n13533) );
  ANDN U15495 ( .B(n7513), .A(n13533), .Z(n7514) );
  NANDN U15496 ( .A(n26714), .B(n7514), .Z(n7515) );
  NAND U15497 ( .A(n26716), .B(n7515), .Z(n7516) );
  ANDN U15498 ( .B(y[1460]), .A(x[1460]), .Z(n13531) );
  OR U15499 ( .A(n7516), .B(n13531), .Z(n7517) );
  NAND U15500 ( .A(n7518), .B(n7517), .Z(n7519) );
  NANDN U15501 ( .A(x[1461]), .B(y[1461]), .Z(n13532) );
  AND U15502 ( .A(n7519), .B(n13532), .Z(n7520) );
  NAND U15503 ( .A(n13528), .B(n7520), .Z(n7521) );
  NANDN U15504 ( .A(n13525), .B(n7521), .Z(n7522) );
  ANDN U15505 ( .B(x[1462]), .A(y[1462]), .Z(n13529) );
  OR U15506 ( .A(n7522), .B(n13529), .Z(n7523) );
  AND U15507 ( .A(n13527), .B(n7523), .Z(n7524) );
  NANDN U15508 ( .A(n17714), .B(n7524), .Z(n7525) );
  NANDN U15509 ( .A(y[1464]), .B(x[1464]), .Z(n13526) );
  NANDN U15510 ( .A(y[1465]), .B(x[1465]), .Z(n17718) );
  AND U15511 ( .A(n13526), .B(n17718), .Z(n24402) );
  AND U15512 ( .A(n7525), .B(n24402), .Z(n7527) );
  NANDN U15513 ( .A(x[1466]), .B(y[1466]), .Z(n13524) );
  ANDN U15514 ( .B(y[1465]), .A(x[1465]), .Z(n17713) );
  ANDN U15515 ( .B(n13524), .A(n17713), .Z(n7526) );
  NANDN U15516 ( .A(n7527), .B(n7526), .Z(n7528) );
  AND U15517 ( .A(n26725), .B(n7528), .Z(n7529) );
  NANDN U15518 ( .A(y[1466]), .B(x[1466]), .Z(n26723) );
  AND U15519 ( .A(n7529), .B(n26723), .Z(n7531) );
  NANDN U15520 ( .A(x[1467]), .B(y[1467]), .Z(n13523) );
  ANDN U15521 ( .B(y[1468]), .A(x[1468]), .Z(n26726) );
  ANDN U15522 ( .B(n13523), .A(n26726), .Z(n7530) );
  NANDN U15523 ( .A(n7531), .B(n7530), .Z(n7532) );
  NANDN U15524 ( .A(n24401), .B(n7532), .Z(n7533) );
  AND U15525 ( .A(n26727), .B(n7533), .Z(n7534) );
  NANDN U15526 ( .A(y[1470]), .B(x[1470]), .Z(n17728) );
  NANDN U15527 ( .A(y[1471]), .B(x[1471]), .Z(n17735) );
  AND U15528 ( .A(n17728), .B(n17735), .Z(n26728) );
  NANDN U15529 ( .A(n7534), .B(n26728), .Z(n7535) );
  NAND U15530 ( .A(n7536), .B(n7535), .Z(n7537) );
  NAND U15531 ( .A(n26731), .B(n7537), .Z(n7538) );
  NANDN U15532 ( .A(n13522), .B(n7538), .Z(n7539) );
  AND U15533 ( .A(n26733), .B(n7539), .Z(n7540) );
  ANDN U15534 ( .B(y[1476]), .A(x[1476]), .Z(n17739) );
  OR U15535 ( .A(n7540), .B(n17739), .Z(n7541) );
  NANDN U15536 ( .A(n26735), .B(n7541), .Z(n7542) );
  NANDN U15537 ( .A(n26736), .B(n7542), .Z(n7543) );
  NANDN U15538 ( .A(x[1477]), .B(y[1477]), .Z(n17740) );
  NANDN U15539 ( .A(n7543), .B(n17740), .Z(n7544) );
  AND U15540 ( .A(n26737), .B(n7544), .Z(n7546) );
  NANDN U15541 ( .A(x[1479]), .B(y[1479]), .Z(n26738) );
  ANDN U15542 ( .B(y[1480]), .A(x[1480]), .Z(n13518) );
  ANDN U15543 ( .B(n26738), .A(n13518), .Z(n7545) );
  NANDN U15544 ( .A(n7546), .B(n7545), .Z(n7547) );
  AND U15545 ( .A(n26741), .B(n7547), .Z(n7548) );
  NANDN U15546 ( .A(y[1480]), .B(x[1480]), .Z(n26739) );
  AND U15547 ( .A(n7548), .B(n26739), .Z(n7550) );
  NANDN U15548 ( .A(x[1481]), .B(y[1481]), .Z(n13519) );
  ANDN U15549 ( .B(y[1482]), .A(x[1482]), .Z(n24400) );
  ANDN U15550 ( .B(n13519), .A(n24400), .Z(n7549) );
  NANDN U15551 ( .A(n7550), .B(n7549), .Z(n7551) );
  NANDN U15552 ( .A(n26742), .B(n7551), .Z(n7552) );
  AND U15553 ( .A(n26743), .B(n7552), .Z(n7554) );
  NANDN U15554 ( .A(y[1484]), .B(x[1484]), .Z(n7553) );
  ANDN U15555 ( .B(x[1485]), .A(y[1485]), .Z(n13516) );
  ANDN U15556 ( .B(n7553), .A(n13516), .Z(n26744) );
  NANDN U15557 ( .A(n7554), .B(n26744), .Z(n7555) );
  NAND U15558 ( .A(n26745), .B(n7555), .Z(n7556) );
  NANDN U15559 ( .A(n26746), .B(n7556), .Z(n7557) );
  AND U15560 ( .A(n26747), .B(n7557), .Z(n7558) );
  NAND U15561 ( .A(n13512), .B(n7558), .Z(n7559) );
  NAND U15562 ( .A(n17764), .B(n7559), .Z(n7560) );
  NANDN U15563 ( .A(n13514), .B(n7560), .Z(n7561) );
  ANDN U15564 ( .B(n7562), .A(n7561), .Z(n7565) );
  NANDN U15565 ( .A(y[1491]), .B(x[1491]), .Z(n7564) );
  NANDN U15566 ( .A(y[1492]), .B(x[1492]), .Z(n7563) );
  NAND U15567 ( .A(n7564), .B(n7563), .Z(n26751) );
  OR U15568 ( .A(n7565), .B(n26751), .Z(n7566) );
  AND U15569 ( .A(n26752), .B(n7566), .Z(n7567) );
  ANDN U15570 ( .B(x[1493]), .A(y[1493]), .Z(n13509) );
  OR U15571 ( .A(n7567), .B(n13509), .Z(n7568) );
  AND U15572 ( .A(n26754), .B(n7568), .Z(n7572) );
  ANDN U15573 ( .B(x[1495]), .A(y[1495]), .Z(n26755) );
  NANDN U15574 ( .A(y[1494]), .B(x[1494]), .Z(n13510) );
  NANDN U15575 ( .A(n26755), .B(n13510), .Z(n7569) );
  AND U15576 ( .A(n7570), .B(n7569), .Z(n7571) );
  OR U15577 ( .A(n7572), .B(n7571), .Z(n7573) );
  NAND U15578 ( .A(n26756), .B(n7573), .Z(n7574) );
  NANDN U15579 ( .A(n26757), .B(n7574), .Z(n7575) );
  AND U15580 ( .A(n26758), .B(n7575), .Z(n7576) );
  NANDN U15581 ( .A(x[1498]), .B(y[1498]), .Z(n17779) );
  NAND U15582 ( .A(n7576), .B(n17779), .Z(n7577) );
  NANDN U15583 ( .A(n7578), .B(n7577), .Z(n7579) );
  AND U15584 ( .A(n26761), .B(n7579), .Z(n7580) );
  NANDN U15585 ( .A(x[1499]), .B(y[1499]), .Z(n17778) );
  NAND U15586 ( .A(n7580), .B(n17778), .Z(n7581) );
  NANDN U15587 ( .A(n24398), .B(n7581), .Z(n7582) );
  AND U15588 ( .A(n26762), .B(n7582), .Z(n7585) );
  NANDN U15589 ( .A(y[1504]), .B(x[1504]), .Z(n7584) );
  NANDN U15590 ( .A(y[1505]), .B(x[1505]), .Z(n7583) );
  NAND U15591 ( .A(n7584), .B(n7583), .Z(n13505) );
  OR U15592 ( .A(n7585), .B(n13505), .Z(n7586) );
  NAND U15593 ( .A(n13504), .B(n7586), .Z(n7587) );
  NAND U15594 ( .A(n26766), .B(n7587), .Z(n7588) );
  NANDN U15595 ( .A(x[1509]), .B(y[1509]), .Z(n13503) );
  AND U15596 ( .A(n7588), .B(n13503), .Z(n7589) );
  NANDN U15597 ( .A(n17799), .B(n7589), .Z(n7590) );
  NAND U15598 ( .A(n26768), .B(n7590), .Z(n7591) );
  NANDN U15599 ( .A(n17798), .B(n7591), .Z(n7592) );
  ANDN U15600 ( .B(y[1512]), .A(x[1512]), .Z(n24397) );
  OR U15601 ( .A(n7592), .B(n24397), .Z(n7593) );
  NANDN U15602 ( .A(y[1512]), .B(x[1512]), .Z(n17802) );
  NANDN U15603 ( .A(y[1513]), .B(x[1513]), .Z(n17806) );
  AND U15604 ( .A(n17802), .B(n17806), .Z(n24396) );
  AND U15605 ( .A(n7593), .B(n24396), .Z(n7595) );
  NANDN U15606 ( .A(x[1514]), .B(y[1514]), .Z(n13502) );
  ANDN U15607 ( .B(y[1513]), .A(x[1513]), .Z(n26771) );
  ANDN U15608 ( .B(n13502), .A(n26771), .Z(n7594) );
  NANDN U15609 ( .A(n7595), .B(n7594), .Z(n7596) );
  AND U15610 ( .A(n7597), .B(n7596), .Z(n7599) );
  ANDN U15611 ( .B(y[1515]), .A(x[1515]), .Z(n13501) );
  ANDN U15612 ( .B(y[1516]), .A(x[1516]), .Z(n26775) );
  NOR U15613 ( .A(n13501), .B(n26775), .Z(n7598) );
  NANDN U15614 ( .A(n7599), .B(n7598), .Z(n7600) );
  NANDN U15615 ( .A(n24395), .B(n7600), .Z(n7601) );
  NANDN U15616 ( .A(x[1517]), .B(y[1517]), .Z(n17814) );
  AND U15617 ( .A(n7601), .B(n17814), .Z(n7602) );
  NAND U15618 ( .A(n13496), .B(n7602), .Z(n7603) );
  AND U15619 ( .A(n26777), .B(n7603), .Z(n7604) );
  OR U15620 ( .A(n13499), .B(n7604), .Z(n7605) );
  NAND U15621 ( .A(n13494), .B(n7605), .Z(n7606) );
  NANDN U15622 ( .A(n13498), .B(n7606), .Z(n7607) );
  ANDN U15623 ( .B(y[1524]), .A(x[1524]), .Z(n13492) );
  OR U15624 ( .A(n7607), .B(n13492), .Z(n7608) );
  AND U15625 ( .A(n13495), .B(n7608), .Z(n7609) );
  NANDN U15626 ( .A(y[1525]), .B(x[1525]), .Z(n13491) );
  AND U15627 ( .A(n7609), .B(n13491), .Z(n7610) );
  NANDN U15628 ( .A(x[1525]), .B(y[1525]), .Z(n13493) );
  NANDN U15629 ( .A(n7610), .B(n13493), .Z(n7611) );
  ANDN U15630 ( .B(y[1526]), .A(x[1526]), .Z(n17822) );
  OR U15631 ( .A(n7611), .B(n17822), .Z(n7612) );
  AND U15632 ( .A(n26784), .B(n7612), .Z(n7613) );
  NANDN U15633 ( .A(n13490), .B(n7613), .Z(n7614) );
  AND U15634 ( .A(n7615), .B(n7614), .Z(n7616) );
  NANDN U15635 ( .A(y[1528]), .B(x[1528]), .Z(n17826) );
  NANDN U15636 ( .A(y[1529]), .B(x[1529]), .Z(n17831) );
  NAND U15637 ( .A(n17826), .B(n17831), .Z(n26786) );
  OR U15638 ( .A(n7616), .B(n26786), .Z(n7617) );
  NAND U15639 ( .A(n26787), .B(n7617), .Z(n7618) );
  NANDN U15640 ( .A(n24394), .B(n7618), .Z(n7619) );
  NANDN U15641 ( .A(x[1532]), .B(y[1532]), .Z(n13488) );
  AND U15642 ( .A(n7619), .B(n13488), .Z(n7620) );
  NAND U15643 ( .A(n17837), .B(n7620), .Z(n7621) );
  NANDN U15644 ( .A(n7622), .B(n7621), .Z(n7623) );
  AND U15645 ( .A(n26791), .B(n7623), .Z(n7624) );
  NAND U15646 ( .A(n13487), .B(n7624), .Z(n7625) );
  NANDN U15647 ( .A(n26792), .B(n7625), .Z(n7626) );
  AND U15648 ( .A(n26793), .B(n7626), .Z(n7627) );
  OR U15649 ( .A(n26794), .B(n7627), .Z(n7628) );
  NAND U15650 ( .A(n26795), .B(n7628), .Z(n7629) );
  NANDN U15651 ( .A(n26797), .B(n7629), .Z(n7630) );
  ANDN U15652 ( .B(x[1541]), .A(y[1541]), .Z(n13485) );
  OR U15653 ( .A(n7630), .B(n13485), .Z(n7631) );
  AND U15654 ( .A(n13484), .B(n7631), .Z(n7632) );
  NANDN U15655 ( .A(x[1541]), .B(y[1541]), .Z(n26798) );
  NAND U15656 ( .A(n7632), .B(n26798), .Z(n7633) );
  NANDN U15657 ( .A(y[1542]), .B(x[1542]), .Z(n13486) );
  AND U15658 ( .A(n7633), .B(n13486), .Z(n7634) );
  NANDN U15659 ( .A(n13481), .B(n7634), .Z(n7636) );
  OR U15660 ( .A(n7636), .B(n7635), .Z(n7637) );
  NAND U15661 ( .A(n7638), .B(n7637), .Z(n7639) );
  NANDN U15662 ( .A(n7640), .B(n7639), .Z(n7641) );
  NANDN U15663 ( .A(x[1548]), .B(y[1548]), .Z(n26806) );
  AND U15664 ( .A(n7641), .B(n26806), .Z(n7642) );
  NANDN U15665 ( .A(x[1547]), .B(y[1547]), .Z(n17863) );
  NAND U15666 ( .A(n7642), .B(n17863), .Z(n7643) );
  NANDN U15667 ( .A(n26807), .B(n7643), .Z(n7644) );
  NANDN U15668 ( .A(x[1549]), .B(y[1549]), .Z(n17870) );
  NANDN U15669 ( .A(x[1550]), .B(y[1550]), .Z(n17876) );
  AND U15670 ( .A(n17870), .B(n17876), .Z(n26808) );
  AND U15671 ( .A(n7644), .B(n26808), .Z(n7645) );
  ANDN U15672 ( .B(x[1550]), .A(y[1550]), .Z(n17872) );
  ANDN U15673 ( .B(x[1551]), .A(y[1551]), .Z(n17880) );
  OR U15674 ( .A(n17872), .B(n17880), .Z(n24391) );
  OR U15675 ( .A(n7645), .B(n24391), .Z(n7646) );
  NANDN U15676 ( .A(x[1551]), .B(y[1551]), .Z(n24390) );
  AND U15677 ( .A(n7646), .B(n24390), .Z(n7647) );
  NAND U15678 ( .A(n13480), .B(n7647), .Z(n7648) );
  AND U15679 ( .A(n17884), .B(n7648), .Z(n7649) );
  NANDN U15680 ( .A(n26810), .B(n7649), .Z(n7650) );
  ANDN U15681 ( .B(y[1554]), .A(x[1554]), .Z(n13477) );
  ANDN U15682 ( .B(n7650), .A(n13477), .Z(n7651) );
  NANDN U15683 ( .A(n13479), .B(n7651), .Z(n7652) );
  AND U15684 ( .A(n24389), .B(n7652), .Z(n7653) );
  NANDN U15685 ( .A(n17883), .B(n7653), .Z(n7654) );
  AND U15686 ( .A(n7655), .B(n7654), .Z(n7657) );
  NANDN U15687 ( .A(y[1557]), .B(x[1557]), .Z(n13474) );
  ANDN U15688 ( .B(x[1556]), .A(y[1556]), .Z(n24388) );
  ANDN U15689 ( .B(n13474), .A(n24388), .Z(n7656) );
  NANDN U15690 ( .A(n7657), .B(n7656), .Z(n7658) );
  AND U15691 ( .A(n13475), .B(n7658), .Z(n7659) );
  NANDN U15692 ( .A(n17892), .B(n7659), .Z(n7660) );
  NANDN U15693 ( .A(y[1559]), .B(x[1559]), .Z(n24387) );
  AND U15694 ( .A(n7660), .B(n24387), .Z(n7661) );
  NANDN U15695 ( .A(n13473), .B(n7661), .Z(n7662) );
  AND U15696 ( .A(n7663), .B(n7662), .Z(n7664) );
  NANDN U15697 ( .A(y[1560]), .B(x[1560]), .Z(n13472) );
  NANDN U15698 ( .A(y[1561]), .B(x[1561]), .Z(n17899) );
  NAND U15699 ( .A(n13472), .B(n17899), .Z(n26818) );
  OR U15700 ( .A(n7664), .B(n26818), .Z(n7665) );
  AND U15701 ( .A(n26819), .B(n7665), .Z(n7666) );
  NANDN U15702 ( .A(n13471), .B(n7666), .Z(n7667) );
  NANDN U15703 ( .A(y[1563]), .B(x[1563]), .Z(n24386) );
  AND U15704 ( .A(n7667), .B(n24386), .Z(n7668) );
  NAND U15705 ( .A(n26820), .B(n7668), .Z(n7669) );
  ANDN U15706 ( .B(y[1564]), .A(x[1564]), .Z(n13468) );
  ANDN U15707 ( .B(n7669), .A(n13468), .Z(n7670) );
  NANDN U15708 ( .A(n13470), .B(n7670), .Z(n7671) );
  NANDN U15709 ( .A(y[1564]), .B(x[1564]), .Z(n24385) );
  AND U15710 ( .A(n7671), .B(n24385), .Z(n7672) );
  NAND U15711 ( .A(n13466), .B(n7672), .Z(n7673) );
  NANDN U15712 ( .A(n13469), .B(n7673), .Z(n7674) );
  ANDN U15713 ( .B(y[1566]), .A(x[1566]), .Z(n13464) );
  OR U15714 ( .A(n7674), .B(n13464), .Z(n7675) );
  NAND U15715 ( .A(n13467), .B(n7675), .Z(n7676) );
  NANDN U15716 ( .A(n13465), .B(n7676), .Z(n7677) );
  NAND U15717 ( .A(n24384), .B(n7677), .Z(n7678) );
  NAND U15718 ( .A(n26827), .B(n7678), .Z(n7679) );
  NANDN U15719 ( .A(n26828), .B(n7679), .Z(n7680) );
  AND U15720 ( .A(n26829), .B(n7680), .Z(n7681) );
  NANDN U15721 ( .A(y[1574]), .B(x[1574]), .Z(n17919) );
  NANDN U15722 ( .A(y[1575]), .B(x[1575]), .Z(n17925) );
  NAND U15723 ( .A(n17919), .B(n17925), .Z(n26830) );
  OR U15724 ( .A(n7681), .B(n26830), .Z(n7682) );
  ANDN U15725 ( .B(y[1575]), .A(x[1575]), .Z(n26831) );
  ANDN U15726 ( .B(n7682), .A(n26831), .Z(n7683) );
  NANDN U15727 ( .A(n13460), .B(n7683), .Z(n7684) );
  NAND U15728 ( .A(n26832), .B(n7684), .Z(n7685) );
  NANDN U15729 ( .A(n13459), .B(n7685), .Z(n7688) );
  NANDN U15730 ( .A(x[1578]), .B(y[1578]), .Z(n7687) );
  AND U15731 ( .A(n7687), .B(n7686), .Z(n26834) );
  NANDN U15732 ( .A(n7688), .B(n26834), .Z(n7689) );
  NAND U15733 ( .A(n26837), .B(n7689), .Z(n7690) );
  NANDN U15734 ( .A(n13457), .B(n7690), .Z(n7691) );
  AND U15735 ( .A(n7692), .B(n7691), .Z(n7695) );
  NANDN U15736 ( .A(x[1582]), .B(y[1582]), .Z(n7693) );
  NAND U15737 ( .A(n7694), .B(n7693), .Z(n13456) );
  OR U15738 ( .A(n7695), .B(n13456), .Z(n7696) );
  NAND U15739 ( .A(n26839), .B(n7696), .Z(n7697) );
  NANDN U15740 ( .A(n26840), .B(n7697), .Z(n7698) );
  NAND U15741 ( .A(n26841), .B(n7698), .Z(n7699) );
  NAND U15742 ( .A(n26842), .B(n7699), .Z(n7700) );
  AND U15743 ( .A(n13455), .B(n7700), .Z(n7701) );
  ANDN U15744 ( .B(y[1588]), .A(x[1588]), .Z(n13452) );
  OR U15745 ( .A(n7701), .B(n13452), .Z(n7702) );
  AND U15746 ( .A(n13454), .B(n7702), .Z(n7703) );
  ANDN U15747 ( .B(x[1589]), .A(y[1589]), .Z(n26845) );
  ANDN U15748 ( .B(n7703), .A(n26845), .Z(n7704) );
  NANDN U15749 ( .A(x[1589]), .B(y[1589]), .Z(n13453) );
  NANDN U15750 ( .A(n7704), .B(n13453), .Z(n7707) );
  NANDN U15751 ( .A(x[1590]), .B(y[1590]), .Z(n7706) );
  ANDN U15752 ( .B(n7706), .A(n7705), .Z(n26846) );
  NANDN U15753 ( .A(n7707), .B(n26846), .Z(n7708) );
  NAND U15754 ( .A(n17944), .B(n7708), .Z(n7709) );
  NAND U15755 ( .A(n13451), .B(n7709), .Z(n7710) );
  NAND U15756 ( .A(n13449), .B(n7710), .Z(n7711) );
  ANDN U15757 ( .B(y[1594]), .A(x[1594]), .Z(n17950) );
  ANDN U15758 ( .B(n7711), .A(n17950), .Z(n7712) );
  NANDN U15759 ( .A(n13450), .B(n7712), .Z(n7713) );
  NANDN U15760 ( .A(n26850), .B(n7713), .Z(n7714) );
  AND U15761 ( .A(n26851), .B(n7714), .Z(n7715) );
  OR U15762 ( .A(n26852), .B(n7715), .Z(n7716) );
  AND U15763 ( .A(n7717), .B(n7716), .Z(n7719) );
  NANDN U15764 ( .A(y[1598]), .B(x[1598]), .Z(n7718) );
  NANDN U15765 ( .A(y[1599]), .B(x[1599]), .Z(n17958) );
  AND U15766 ( .A(n7718), .B(n17958), .Z(n13448) );
  NANDN U15767 ( .A(n7719), .B(n13448), .Z(n7720) );
  AND U15768 ( .A(n17960), .B(n7720), .Z(n7723) );
  NANDN U15769 ( .A(y[1601]), .B(x[1601]), .Z(n7722) );
  NANDN U15770 ( .A(y[1600]), .B(x[1600]), .Z(n7721) );
  AND U15771 ( .A(n7722), .B(n7721), .Z(n26857) );
  NANDN U15772 ( .A(n7723), .B(n26857), .Z(n7724) );
  ANDN U15773 ( .B(y[1601]), .A(x[1601]), .Z(n26858) );
  ANDN U15774 ( .B(n7724), .A(n26858), .Z(n7725) );
  NANDN U15775 ( .A(x[1602]), .B(y[1602]), .Z(n17965) );
  AND U15776 ( .A(n7725), .B(n17965), .Z(n7726) );
  ANDN U15777 ( .B(n26859), .A(n7726), .Z(n7731) );
  NANDN U15778 ( .A(x[1604]), .B(y[1604]), .Z(n7728) );
  NANDN U15779 ( .A(x[1603]), .B(y[1603]), .Z(n7727) );
  AND U15780 ( .A(n7728), .B(n7727), .Z(n7730) );
  NAND U15781 ( .A(n7730), .B(n7729), .Z(n17967) );
  OR U15782 ( .A(n7731), .B(n17967), .Z(n7732) );
  NAND U15783 ( .A(n13447), .B(n7732), .Z(n7733) );
  NANDN U15784 ( .A(n13445), .B(n7733), .Z(n7734) );
  NANDN U15785 ( .A(y[1607]), .B(x[1607]), .Z(n26863) );
  AND U15786 ( .A(n7734), .B(n26863), .Z(n7735) );
  NAND U15787 ( .A(n13446), .B(n7735), .Z(n7736) );
  NANDN U15788 ( .A(n24381), .B(n7736), .Z(n7737) );
  ANDN U15789 ( .B(y[1607]), .A(x[1607]), .Z(n13444) );
  OR U15790 ( .A(n7737), .B(n13444), .Z(n7738) );
  NAND U15791 ( .A(n26864), .B(n7738), .Z(n7739) );
  NANDN U15792 ( .A(n26865), .B(n7739), .Z(n7740) );
  NANDN U15793 ( .A(n26866), .B(n7740), .Z(n7741) );
  NAND U15794 ( .A(n26867), .B(n7741), .Z(n7742) );
  NANDN U15795 ( .A(n26868), .B(n7742), .Z(n7743) );
  AND U15796 ( .A(n26869), .B(n7743), .Z(n7744) );
  ANDN U15797 ( .B(x[1612]), .A(y[1612]), .Z(n17981) );
  ANDN U15798 ( .B(x[1613]), .A(y[1613]), .Z(n17985) );
  OR U15799 ( .A(n17981), .B(n17985), .Z(n26870) );
  OR U15800 ( .A(n7744), .B(n26870), .Z(n7745) );
  AND U15801 ( .A(n26872), .B(n7745), .Z(n7746) );
  NANDN U15802 ( .A(x[1614]), .B(y[1614]), .Z(n13442) );
  NAND U15803 ( .A(n7746), .B(n13442), .Z(n7747) );
  NANDN U15804 ( .A(y[1615]), .B(x[1615]), .Z(n26875) );
  AND U15805 ( .A(n7747), .B(n26875), .Z(n7748) );
  NANDN U15806 ( .A(n26873), .B(n7748), .Z(n7749) );
  ANDN U15807 ( .B(y[1616]), .A(x[1616]), .Z(n26876) );
  ANDN U15808 ( .B(n7749), .A(n26876), .Z(n7750) );
  NANDN U15809 ( .A(n13441), .B(n7750), .Z(n7751) );
  NAND U15810 ( .A(n24380), .B(n7751), .Z(n7752) );
  NANDN U15811 ( .A(n24379), .B(n7752), .Z(n7753) );
  NANDN U15812 ( .A(y[1618]), .B(x[1618]), .Z(n24378) );
  AND U15813 ( .A(n7753), .B(n24378), .Z(n7754) );
  NANDN U15814 ( .A(n13439), .B(n7754), .Z(n7755) );
  NAND U15815 ( .A(n7756), .B(n7755), .Z(n7757) );
  AND U15816 ( .A(n13440), .B(n7757), .Z(n7758) );
  NANDN U15817 ( .A(n13437), .B(n7758), .Z(n7759) );
  NAND U15818 ( .A(n7760), .B(n7759), .Z(n7761) );
  NANDN U15819 ( .A(y[1623]), .B(x[1623]), .Z(n24376) );
  AND U15820 ( .A(n7761), .B(n24376), .Z(n7762) );
  NAND U15821 ( .A(n13438), .B(n7762), .Z(n7763) );
  NANDN U15822 ( .A(n26881), .B(n7763), .Z(n7764) );
  ANDN U15823 ( .B(y[1623]), .A(x[1623]), .Z(n13435) );
  OR U15824 ( .A(n7764), .B(n13435), .Z(n7765) );
  NANDN U15825 ( .A(y[1624]), .B(x[1624]), .Z(n18006) );
  NANDN U15826 ( .A(y[1625]), .B(x[1625]), .Z(n13434) );
  AND U15827 ( .A(n18006), .B(n13434), .Z(n26884) );
  AND U15828 ( .A(n7765), .B(n26884), .Z(n7766) );
  ANDN U15829 ( .B(y[1625]), .A(x[1625]), .Z(n18010) );
  NANDN U15830 ( .A(x[1626]), .B(y[1626]), .Z(n13432) );
  NANDN U15831 ( .A(n18010), .B(n13432), .Z(n24375) );
  OR U15832 ( .A(n7766), .B(n24375), .Z(n7767) );
  NAND U15833 ( .A(n24374), .B(n7767), .Z(n7768) );
  NANDN U15834 ( .A(n13431), .B(n7768), .Z(n7769) );
  ANDN U15835 ( .B(y[1628]), .A(x[1628]), .Z(n18019) );
  OR U15836 ( .A(n7769), .B(n18019), .Z(n7770) );
  NAND U15837 ( .A(n26887), .B(n7770), .Z(n7771) );
  NAND U15838 ( .A(n26888), .B(n7771), .Z(n7772) );
  OR U15839 ( .A(n18018), .B(n7772), .Z(n7773) );
  AND U15840 ( .A(n26890), .B(n7773), .Z(n7774) );
  NANDN U15841 ( .A(x[1631]), .B(y[1631]), .Z(n18026) );
  NANDN U15842 ( .A(x[1632]), .B(y[1632]), .Z(n18032) );
  NAND U15843 ( .A(n18026), .B(n18032), .Z(n26891) );
  OR U15844 ( .A(n7774), .B(n26891), .Z(n7775) );
  AND U15845 ( .A(n26892), .B(n7775), .Z(n7776) );
  OR U15846 ( .A(n26893), .B(n7776), .Z(n7777) );
  NAND U15847 ( .A(n26894), .B(n7777), .Z(n7778) );
  NANDN U15848 ( .A(n26895), .B(n7778), .Z(n7779) );
  ANDN U15849 ( .B(y[1636]), .A(x[1636]), .Z(n13427) );
  OR U15850 ( .A(n7779), .B(n13427), .Z(n7780) );
  NAND U15851 ( .A(n7781), .B(n7780), .Z(n7782) );
  NAND U15852 ( .A(n13428), .B(n7782), .Z(n7783) );
  OR U15853 ( .A(n26899), .B(n7783), .Z(n7784) );
  AND U15854 ( .A(n26901), .B(n7784), .Z(n7785) );
  OR U15855 ( .A(n26902), .B(n7785), .Z(n7786) );
  NAND U15856 ( .A(n26903), .B(n7786), .Z(n7787) );
  NANDN U15857 ( .A(n24373), .B(n7787), .Z(n7788) );
  NANDN U15858 ( .A(y[1642]), .B(x[1642]), .Z(n24372) );
  AND U15859 ( .A(n7788), .B(n24372), .Z(n7789) );
  NAND U15860 ( .A(n18067), .B(n7789), .Z(n7790) );
  NANDN U15861 ( .A(n24371), .B(n7790), .Z(n7791) );
  ANDN U15862 ( .B(y[1644]), .A(x[1644]), .Z(n18069) );
  OR U15863 ( .A(n7791), .B(n18069), .Z(n7792) );
  NANDN U15864 ( .A(n7793), .B(n7792), .Z(n7794) );
  AND U15865 ( .A(n7795), .B(n7794), .Z(n7796) );
  NANDN U15866 ( .A(y[1646]), .B(x[1646]), .Z(n13426) );
  NANDN U15867 ( .A(y[1647]), .B(x[1647]), .Z(n18077) );
  NAND U15868 ( .A(n13426), .B(n18077), .Z(n26907) );
  OR U15869 ( .A(n7796), .B(n26907), .Z(n7797) );
  ANDN U15870 ( .B(y[1647]), .A(x[1647]), .Z(n26908) );
  ANDN U15871 ( .B(n7797), .A(n26908), .Z(n7798) );
  NANDN U15872 ( .A(x[1648]), .B(y[1648]), .Z(n13425) );
  NAND U15873 ( .A(n7798), .B(n13425), .Z(n7799) );
  NANDN U15874 ( .A(y[1649]), .B(x[1649]), .Z(n13423) );
  AND U15875 ( .A(n7799), .B(n13423), .Z(n7800) );
  NAND U15876 ( .A(n26909), .B(n7800), .Z(n7801) );
  AND U15877 ( .A(n13424), .B(n7801), .Z(n7802) );
  NANDN U15878 ( .A(x[1650]), .B(y[1650]), .Z(n18082) );
  NAND U15879 ( .A(n7802), .B(n18082), .Z(n7803) );
  ANDN U15880 ( .B(x[1651]), .A(y[1651]), .Z(n13420) );
  ANDN U15881 ( .B(n7803), .A(n13420), .Z(n7804) );
  NANDN U15882 ( .A(n13422), .B(n7804), .Z(n7806) );
  NANDN U15883 ( .A(x[1652]), .B(y[1652]), .Z(n13419) );
  NANDN U15884 ( .A(x[1651]), .B(y[1651]), .Z(n18081) );
  AND U15885 ( .A(n13419), .B(n18081), .Z(n7805) );
  NAND U15886 ( .A(n7806), .B(n7805), .Z(n7807) );
  AND U15887 ( .A(n13421), .B(n7807), .Z(n7808) );
  NANDN U15888 ( .A(y[1653]), .B(x[1653]), .Z(n13417) );
  AND U15889 ( .A(n7808), .B(n13417), .Z(n7810) );
  NANDN U15890 ( .A(x[1654]), .B(y[1654]), .Z(n13414) );
  ANDN U15891 ( .B(y[1653]), .A(x[1653]), .Z(n13418) );
  ANDN U15892 ( .B(n13414), .A(n13418), .Z(n7809) );
  NANDN U15893 ( .A(n7810), .B(n7809), .Z(n7811) );
  NAND U15894 ( .A(n26917), .B(n7811), .Z(n7812) );
  ANDN U15895 ( .B(x[1654]), .A(y[1654]), .Z(n13416) );
  OR U15896 ( .A(n7812), .B(n13416), .Z(n7813) );
  AND U15897 ( .A(n7814), .B(n7813), .Z(n7815) );
  NANDN U15898 ( .A(y[1656]), .B(x[1656]), .Z(n18089) );
  NANDN U15899 ( .A(y[1657]), .B(x[1657]), .Z(n18093) );
  NAND U15900 ( .A(n18089), .B(n18093), .Z(n26919) );
  OR U15901 ( .A(n7815), .B(n26919), .Z(n7816) );
  ANDN U15902 ( .B(y[1657]), .A(x[1657]), .Z(n26920) );
  ANDN U15903 ( .B(n7816), .A(n26920), .Z(n7817) );
  NANDN U15904 ( .A(n13413), .B(n7817), .Z(n7818) );
  AND U15905 ( .A(n13411), .B(n7818), .Z(n7819) );
  NAND U15906 ( .A(n24368), .B(n7819), .Z(n7820) );
  NANDN U15907 ( .A(x[1660]), .B(y[1660]), .Z(n13409) );
  AND U15908 ( .A(n7820), .B(n13409), .Z(n7821) );
  NANDN U15909 ( .A(n13412), .B(n7821), .Z(n7822) );
  AND U15910 ( .A(n13410), .B(n7822), .Z(n7823) );
  NANDN U15911 ( .A(y[1661]), .B(x[1661]), .Z(n13407) );
  NAND U15912 ( .A(n7823), .B(n13407), .Z(n7824) );
  ANDN U15913 ( .B(y[1662]), .A(x[1662]), .Z(n13404) );
  ANDN U15914 ( .B(n7824), .A(n13404), .Z(n7825) );
  NANDN U15915 ( .A(n13408), .B(n7825), .Z(n7827) );
  NANDN U15916 ( .A(y[1662]), .B(x[1662]), .Z(n13406) );
  NANDN U15917 ( .A(y[1663]), .B(x[1663]), .Z(n18103) );
  AND U15918 ( .A(n13406), .B(n18103), .Z(n7826) );
  NAND U15919 ( .A(n7827), .B(n7826), .Z(n7828) );
  AND U15920 ( .A(n13405), .B(n7828), .Z(n7829) );
  AND U15921 ( .A(n26927), .B(n7829), .Z(n7832) );
  NANDN U15922 ( .A(y[1665]), .B(x[1665]), .Z(n18109) );
  ANDN U15923 ( .B(x[1664]), .A(y[1664]), .Z(n18102) );
  NAND U15924 ( .A(n18102), .B(n7830), .Z(n7831) );
  NAND U15925 ( .A(n18109), .B(n7831), .Z(n26929) );
  OR U15926 ( .A(n7832), .B(n26929), .Z(n7833) );
  ANDN U15927 ( .B(y[1666]), .A(x[1666]), .Z(n26930) );
  ANDN U15928 ( .B(n7833), .A(n26930), .Z(n7834) );
  NANDN U15929 ( .A(y[1666]), .B(x[1666]), .Z(n18107) );
  NANDN U15930 ( .A(y[1667]), .B(x[1667]), .Z(n18114) );
  NAND U15931 ( .A(n18107), .B(n18114), .Z(n26931) );
  OR U15932 ( .A(n7834), .B(n26931), .Z(n7835) );
  AND U15933 ( .A(n26932), .B(n7835), .Z(n7837) );
  ANDN U15934 ( .B(x[1669]), .A(y[1669]), .Z(n13400) );
  ANDN U15935 ( .B(x[1668]), .A(y[1668]), .Z(n26933) );
  NOR U15936 ( .A(n13400), .B(n26933), .Z(n7836) );
  NANDN U15937 ( .A(n7837), .B(n7836), .Z(n7838) );
  NANDN U15938 ( .A(n13402), .B(n7838), .Z(n7839) );
  ANDN U15939 ( .B(y[1670]), .A(x[1670]), .Z(n13398) );
  OR U15940 ( .A(n7839), .B(n13398), .Z(n7840) );
  AND U15941 ( .A(n13401), .B(n7840), .Z(n7841) );
  NANDN U15942 ( .A(y[1671]), .B(x[1671]), .Z(n13397) );
  AND U15943 ( .A(n7841), .B(n13397), .Z(n7842) );
  NANDN U15944 ( .A(x[1671]), .B(y[1671]), .Z(n13399) );
  NANDN U15945 ( .A(n7842), .B(n13399), .Z(n7844) );
  NANDN U15946 ( .A(x[1672]), .B(n7844), .Z(n7843) );
  ANDN U15947 ( .B(y[1673]), .A(x[1673]), .Z(n13395) );
  ANDN U15948 ( .B(n7843), .A(n13395), .Z(n7847) );
  XNOR U15949 ( .A(n7844), .B(x[1672]), .Z(n7845) );
  NAND U15950 ( .A(n7845), .B(y[1672]), .Z(n7846) );
  NAND U15951 ( .A(n7847), .B(n7846), .Z(n7850) );
  NANDN U15952 ( .A(y[1674]), .B(x[1674]), .Z(n7849) );
  NANDN U15953 ( .A(y[1673]), .B(x[1673]), .Z(n7848) );
  AND U15954 ( .A(n7849), .B(n7848), .Z(n24367) );
  AND U15955 ( .A(n7850), .B(n24367), .Z(n7853) );
  NANDN U15956 ( .A(x[1674]), .B(y[1674]), .Z(n7852) );
  NANDN U15957 ( .A(x[1675]), .B(y[1675]), .Z(n7851) );
  NAND U15958 ( .A(n7852), .B(n7851), .Z(n26939) );
  OR U15959 ( .A(n7853), .B(n26939), .Z(n7854) );
  NAND U15960 ( .A(n26940), .B(n7854), .Z(n7855) );
  NANDN U15961 ( .A(n26941), .B(n7855), .Z(n7856) );
  AND U15962 ( .A(n26942), .B(n7856), .Z(n7857) );
  ANDN U15963 ( .B(y[1678]), .A(x[1678]), .Z(n13393) );
  OR U15964 ( .A(n7857), .B(n13393), .Z(n7858) );
  NAND U15965 ( .A(n24366), .B(n7858), .Z(n7859) );
  NANDN U15966 ( .A(n13392), .B(n7859), .Z(n7860) );
  XNOR U15967 ( .A(y[1680]), .B(x[1680]), .Z(n13391) );
  NANDN U15968 ( .A(n7860), .B(n13391), .Z(n7861) );
  NAND U15969 ( .A(n7862), .B(n7861), .Z(n7863) );
  NANDN U15970 ( .A(n7864), .B(n7863), .Z(n7865) );
  AND U15971 ( .A(n13386), .B(n7865), .Z(n7866) );
  NANDN U15972 ( .A(y[1683]), .B(x[1683]), .Z(n13383) );
  NAND U15973 ( .A(n7866), .B(n13383), .Z(n7867) );
  NANDN U15974 ( .A(x[1683]), .B(y[1683]), .Z(n13384) );
  AND U15975 ( .A(n7867), .B(n13384), .Z(n7868) );
  NAND U15976 ( .A(n13381), .B(n7868), .Z(n7869) );
  NANDN U15977 ( .A(n18137), .B(n7869), .Z(n7870) );
  ANDN U15978 ( .B(x[1684]), .A(y[1684]), .Z(n13382) );
  OR U15979 ( .A(n7870), .B(n13382), .Z(n7871) );
  AND U15980 ( .A(n13380), .B(n7871), .Z(n7872) );
  NAND U15981 ( .A(n26953), .B(n7872), .Z(n7873) );
  NANDN U15982 ( .A(n24365), .B(n7873), .Z(n7874) );
  NANDN U15983 ( .A(x[1689]), .B(y[1689]), .Z(n13379) );
  AND U15984 ( .A(n7874), .B(n13379), .Z(n7875) );
  NANDN U15985 ( .A(x[1690]), .B(y[1690]), .Z(n13378) );
  NAND U15986 ( .A(n7875), .B(n13378), .Z(n7876) );
  NANDN U15987 ( .A(y[1691]), .B(x[1691]), .Z(n13376) );
  AND U15988 ( .A(n7876), .B(n13376), .Z(n7877) );
  NANDN U15989 ( .A(n18149), .B(n7877), .Z(n7878) );
  AND U15990 ( .A(n13377), .B(n7878), .Z(n7879) );
  NANDN U15991 ( .A(x[1692]), .B(y[1692]), .Z(n13374) );
  NAND U15992 ( .A(n7879), .B(n13374), .Z(n7880) );
  ANDN U15993 ( .B(x[1693]), .A(y[1693]), .Z(n13372) );
  ANDN U15994 ( .B(n7880), .A(n13372), .Z(n7881) );
  NANDN U15995 ( .A(n13375), .B(n7881), .Z(n7883) );
  NANDN U15996 ( .A(x[1693]), .B(y[1693]), .Z(n13373) );
  NANDN U15997 ( .A(x[1694]), .B(y[1694]), .Z(n13371) );
  AND U15998 ( .A(n13373), .B(n13371), .Z(n7882) );
  NAND U15999 ( .A(n7883), .B(n7882), .Z(n7884) );
  AND U16000 ( .A(n18157), .B(n7884), .Z(n7885) );
  NANDN U16001 ( .A(x[1695]), .B(y[1695]), .Z(n24364) );
  NANDN U16002 ( .A(x[1696]), .B(y[1696]), .Z(n26965) );
  NAND U16003 ( .A(n24364), .B(n26965), .Z(n18158) );
  OR U16004 ( .A(n7885), .B(n18158), .Z(n7886) );
  AND U16005 ( .A(n26964), .B(n7886), .Z(n7887) );
  NANDN U16006 ( .A(y[1697]), .B(x[1697]), .Z(n13370) );
  AND U16007 ( .A(n7887), .B(n13370), .Z(n7888) );
  OR U16008 ( .A(n7889), .B(n7888), .Z(n7890) );
  AND U16009 ( .A(n7891), .B(n7890), .Z(n7896) );
  NANDN U16010 ( .A(x[1701]), .B(y[1701]), .Z(n7893) );
  NANDN U16011 ( .A(x[1700]), .B(y[1700]), .Z(n7892) );
  NAND U16012 ( .A(n7893), .B(n7892), .Z(n18169) );
  ANDN U16013 ( .B(y[1699]), .A(x[1699]), .Z(n18165) );
  NAND U16014 ( .A(n18165), .B(n7894), .Z(n7895) );
  NANDN U16015 ( .A(n18169), .B(n7895), .Z(n26970) );
  OR U16016 ( .A(n7896), .B(n26970), .Z(n7897) );
  NAND U16017 ( .A(n13368), .B(n7897), .Z(n7898) );
  NANDN U16018 ( .A(n13365), .B(n7898), .Z(n7900) );
  NANDN U16019 ( .A(y[1703]), .B(x[1703]), .Z(n13364) );
  NANDN U16020 ( .A(y[1702]), .B(x[1702]), .Z(n13367) );
  AND U16021 ( .A(n13364), .B(n13367), .Z(n7899) );
  NAND U16022 ( .A(n7900), .B(n7899), .Z(n7901) );
  AND U16023 ( .A(n13366), .B(n7901), .Z(n7902) );
  NANDN U16024 ( .A(x[1704]), .B(y[1704]), .Z(n13362) );
  NAND U16025 ( .A(n7902), .B(n13362), .Z(n7903) );
  ANDN U16026 ( .B(x[1705]), .A(y[1705]), .Z(n13359) );
  ANDN U16027 ( .B(n7903), .A(n13359), .Z(n7904) );
  NANDN U16028 ( .A(n13363), .B(n7904), .Z(n7905) );
  AND U16029 ( .A(n13361), .B(n7905), .Z(n7906) );
  NANDN U16030 ( .A(x[1706]), .B(y[1706]), .Z(n13358) );
  NAND U16031 ( .A(n7906), .B(n13358), .Z(n7907) );
  ANDN U16032 ( .B(x[1707]), .A(y[1707]), .Z(n24363) );
  ANDN U16033 ( .B(n7907), .A(n24363), .Z(n7908) );
  NAND U16034 ( .A(n13360), .B(n7908), .Z(n7911) );
  NANDN U16035 ( .A(x[1708]), .B(y[1708]), .Z(n7909) );
  AND U16036 ( .A(n7910), .B(n7909), .Z(n24362) );
  AND U16037 ( .A(n7911), .B(n24362), .Z(n7912) );
  NAND U16038 ( .A(n13357), .B(n7912), .Z(n7913) );
  NANDN U16039 ( .A(n24361), .B(n7913), .Z(n7915) );
  NANDN U16040 ( .A(x[1712]), .B(y[1712]), .Z(n18187) );
  NANDN U16041 ( .A(x[1711]), .B(y[1711]), .Z(n7914) );
  AND U16042 ( .A(n18187), .B(n7914), .Z(n24360) );
  AND U16043 ( .A(n7915), .B(n24360), .Z(n7918) );
  NANDN U16044 ( .A(y[1712]), .B(x[1712]), .Z(n7917) );
  NANDN U16045 ( .A(y[1713]), .B(x[1713]), .Z(n7916) );
  NAND U16046 ( .A(n7917), .B(n7916), .Z(n18188) );
  OR U16047 ( .A(n7918), .B(n18188), .Z(n7919) );
  NAND U16048 ( .A(n13352), .B(n7919), .Z(n7920) );
  NANDN U16049 ( .A(n18191), .B(n7920), .Z(n7921) );
  NAND U16050 ( .A(n18193), .B(n7921), .Z(n7922) );
  NANDN U16051 ( .A(y[1717]), .B(x[1717]), .Z(n13351) );
  AND U16052 ( .A(n7922), .B(n13351), .Z(n7923) );
  NANDN U16053 ( .A(n18195), .B(n7923), .Z(n7924) );
  NANDN U16054 ( .A(x[1717]), .B(y[1717]), .Z(n18197) );
  AND U16055 ( .A(n7924), .B(n18197), .Z(n7925) );
  NAND U16056 ( .A(n13349), .B(n7925), .Z(n7926) );
  NANDN U16057 ( .A(n13350), .B(n7926), .Z(n7927) );
  ANDN U16058 ( .B(x[1719]), .A(y[1719]), .Z(n13346) );
  OR U16059 ( .A(n7927), .B(n13346), .Z(n7928) );
  AND U16060 ( .A(n13348), .B(n7928), .Z(n7929) );
  NANDN U16061 ( .A(n26987), .B(n7929), .Z(n7930) );
  AND U16062 ( .A(n7931), .B(n7930), .Z(n7932) );
  OR U16063 ( .A(n26990), .B(n7932), .Z(n7933) );
  NAND U16064 ( .A(n26991), .B(n7933), .Z(n7934) );
  NANDN U16065 ( .A(n26992), .B(n7934), .Z(n7935) );
  ANDN U16066 ( .B(x[1724]), .A(y[1724]), .Z(n26993) );
  ANDN U16067 ( .B(n7935), .A(n26993), .Z(n7936) );
  NAND U16068 ( .A(n18217), .B(n7936), .Z(n7937) );
  NAND U16069 ( .A(n26994), .B(n7937), .Z(n7938) );
  ANDN U16070 ( .B(y[1726]), .A(x[1726]), .Z(n13342) );
  OR U16071 ( .A(n7938), .B(n13342), .Z(n7939) );
  AND U16072 ( .A(n7940), .B(n7939), .Z(n7942) );
  NANDN U16073 ( .A(x[1728]), .B(y[1728]), .Z(n13339) );
  NANDN U16074 ( .A(x[1727]), .B(y[1727]), .Z(n13343) );
  AND U16075 ( .A(n13339), .B(n13343), .Z(n7941) );
  NANDN U16076 ( .A(n7942), .B(n7941), .Z(n7943) );
  NANDN U16077 ( .A(n13336), .B(n7943), .Z(n7944) );
  ANDN U16078 ( .B(x[1728]), .A(y[1728]), .Z(n13340) );
  OR U16079 ( .A(n7944), .B(n13340), .Z(n7945) );
  NANDN U16080 ( .A(x[1730]), .B(y[1730]), .Z(n26999) );
  AND U16081 ( .A(n7945), .B(n26999), .Z(n7946) );
  NANDN U16082 ( .A(n13338), .B(n7946), .Z(n7947) );
  AND U16083 ( .A(n27000), .B(n7947), .Z(n7948) );
  OR U16084 ( .A(n27001), .B(n7948), .Z(n7949) );
  NAND U16085 ( .A(n27002), .B(n7949), .Z(n7950) );
  NANDN U16086 ( .A(n27003), .B(n7950), .Z(n7951) );
  NANDN U16087 ( .A(y[1734]), .B(x[1734]), .Z(n27004) );
  AND U16088 ( .A(n7951), .B(n27004), .Z(n7952) );
  NAND U16089 ( .A(n13330), .B(n7952), .Z(n7953) );
  NANDN U16090 ( .A(n27005), .B(n7953), .Z(n7954) );
  ANDN U16091 ( .B(y[1736]), .A(x[1736]), .Z(n18237) );
  OR U16092 ( .A(n7954), .B(n18237), .Z(n7955) );
  NAND U16093 ( .A(n7956), .B(n7955), .Z(n7957) );
  AND U16094 ( .A(n18241), .B(n7957), .Z(n7958) );
  NAND U16095 ( .A(n18238), .B(n7958), .Z(n7959) );
  NANDN U16096 ( .A(n27009), .B(n7959), .Z(n7960) );
  ANDN U16097 ( .B(x[1739]), .A(y[1739]), .Z(n18248) );
  OR U16098 ( .A(n7960), .B(n18248), .Z(n7961) );
  AND U16099 ( .A(n18244), .B(n7961), .Z(n7962) );
  NANDN U16100 ( .A(x[1740]), .B(y[1740]), .Z(n13328) );
  NAND U16101 ( .A(n7962), .B(n13328), .Z(n7963) );
  ANDN U16102 ( .B(x[1741]), .A(y[1741]), .Z(n13326) );
  ANDN U16103 ( .B(n7963), .A(n13326), .Z(n7964) );
  NANDN U16104 ( .A(n18247), .B(n7964), .Z(n7965) );
  NANDN U16105 ( .A(x[1742]), .B(y[1742]), .Z(n24357) );
  AND U16106 ( .A(n7965), .B(n24357), .Z(n7966) );
  NANDN U16107 ( .A(x[1741]), .B(y[1741]), .Z(n13327) );
  NAND U16108 ( .A(n7966), .B(n13327), .Z(n7967) );
  ANDN U16109 ( .B(x[1742]), .A(y[1742]), .Z(n13325) );
  ANDN U16110 ( .B(n7967), .A(n13325), .Z(n7968) );
  NANDN U16111 ( .A(n24356), .B(n7968), .Z(n7969) );
  NANDN U16112 ( .A(n27014), .B(n7969), .Z(n7970) );
  AND U16113 ( .A(n27015), .B(n7970), .Z(n7972) );
  NANDN U16114 ( .A(x[1745]), .B(y[1745]), .Z(n27016) );
  ANDN U16115 ( .B(y[1746]), .A(x[1746]), .Z(n13321) );
  ANDN U16116 ( .B(n27016), .A(n13321), .Z(n7971) );
  NANDN U16117 ( .A(n7972), .B(n7971), .Z(n7973) );
  AND U16118 ( .A(n27017), .B(n7973), .Z(n7974) );
  NANDN U16119 ( .A(x[1747]), .B(y[1747]), .Z(n13322) );
  NANDN U16120 ( .A(n7974), .B(n13322), .Z(n7977) );
  NANDN U16121 ( .A(y[1748]), .B(x[1748]), .Z(n7976) );
  NANDN U16122 ( .A(y[1747]), .B(x[1747]), .Z(n7975) );
  NAND U16123 ( .A(n7976), .B(n7975), .Z(n27019) );
  ANDN U16124 ( .B(n7977), .A(n27019), .Z(n7978) );
  ANDN U16125 ( .B(n24355), .A(n7978), .Z(n7981) );
  NANDN U16126 ( .A(y[1749]), .B(x[1749]), .Z(n7980) );
  NANDN U16127 ( .A(y[1750]), .B(x[1750]), .Z(n7979) );
  NAND U16128 ( .A(n7980), .B(n7979), .Z(n27022) );
  OR U16129 ( .A(n7981), .B(n27022), .Z(n7982) );
  NAND U16130 ( .A(n27023), .B(n7982), .Z(n7983) );
  NANDN U16131 ( .A(n27024), .B(n7983), .Z(n7984) );
  NAND U16132 ( .A(n18269), .B(n7984), .Z(n7985) );
  NAND U16133 ( .A(n27026), .B(n7985), .Z(n7986) );
  AND U16134 ( .A(n27027), .B(n7986), .Z(n7987) );
  OR U16135 ( .A(n27029), .B(n7987), .Z(n7988) );
  NAND U16136 ( .A(n27030), .B(n7988), .Z(n7989) );
  NANDN U16137 ( .A(n27031), .B(n7989), .Z(n7990) );
  ANDN U16138 ( .B(x[1757]), .A(y[1757]), .Z(n13318) );
  OR U16139 ( .A(n7990), .B(n13318), .Z(n7991) );
  NAND U16140 ( .A(n7992), .B(n7991), .Z(n7993) );
  NANDN U16141 ( .A(y[1758]), .B(x[1758]), .Z(n13319) );
  AND U16142 ( .A(n7993), .B(n13319), .Z(n7994) );
  NAND U16143 ( .A(n13317), .B(n7994), .Z(n7995) );
  NANDN U16144 ( .A(n18282), .B(n7995), .Z(n7996) );
  ANDN U16145 ( .B(y[1760]), .A(x[1760]), .Z(n13314) );
  OR U16146 ( .A(n7996), .B(n13314), .Z(n7997) );
  AND U16147 ( .A(n13316), .B(n7997), .Z(n7998) );
  NANDN U16148 ( .A(y[1761]), .B(x[1761]), .Z(n18288) );
  AND U16149 ( .A(n7998), .B(n18288), .Z(n7999) );
  NANDN U16150 ( .A(x[1761]), .B(y[1761]), .Z(n13315) );
  NANDN U16151 ( .A(n7999), .B(n13315), .Z(n8000) );
  ANDN U16152 ( .B(y[1762]), .A(x[1762]), .Z(n18291) );
  OR U16153 ( .A(n8000), .B(n18291), .Z(n8001) );
  AND U16154 ( .A(n18287), .B(n8001), .Z(n8002) );
  NANDN U16155 ( .A(y[1763]), .B(x[1763]), .Z(n13313) );
  NAND U16156 ( .A(n8002), .B(n13313), .Z(n8003) );
  ANDN U16157 ( .B(y[1764]), .A(x[1764]), .Z(n27040) );
  ANDN U16158 ( .B(n8003), .A(n27040), .Z(n8004) );
  NANDN U16159 ( .A(n18290), .B(n8004), .Z(n8005) );
  AND U16160 ( .A(n27041), .B(n8005), .Z(n8006) );
  NANDN U16161 ( .A(y[1764]), .B(x[1764]), .Z(n13312) );
  AND U16162 ( .A(n8006), .B(n13312), .Z(n8007) );
  OR U16163 ( .A(n27042), .B(n8007), .Z(n8008) );
  NAND U16164 ( .A(n27043), .B(n8008), .Z(n8009) );
  NANDN U16165 ( .A(n27044), .B(n8009), .Z(n8010) );
  NANDN U16166 ( .A(x[1768]), .B(y[1768]), .Z(n13310) );
  NANDN U16167 ( .A(n8010), .B(n13310), .Z(n8011) );
  AND U16168 ( .A(n27045), .B(n8011), .Z(n8012) );
  NANDN U16169 ( .A(y[1769]), .B(x[1769]), .Z(n13308) );
  NAND U16170 ( .A(n8012), .B(n13308), .Z(n8013) );
  ANDN U16171 ( .B(y[1770]), .A(x[1770]), .Z(n13305) );
  ANDN U16172 ( .B(n8013), .A(n13305), .Z(n8014) );
  NANDN U16173 ( .A(n13309), .B(n8014), .Z(n8015) );
  NANDN U16174 ( .A(y[1770]), .B(x[1770]), .Z(n13307) );
  AND U16175 ( .A(n8015), .B(n13307), .Z(n8016) );
  NAND U16176 ( .A(n13304), .B(n8016), .Z(n8017) );
  NAND U16177 ( .A(n13306), .B(n8017), .Z(n8018) );
  ANDN U16178 ( .B(y[1772]), .A(x[1772]), .Z(n13301) );
  OR U16179 ( .A(n8018), .B(n13301), .Z(n8019) );
  AND U16180 ( .A(n8020), .B(n8019), .Z(n8021) );
  NANDN U16181 ( .A(n18310), .B(n8021), .Z(n8022) );
  AND U16182 ( .A(n8023), .B(n8022), .Z(n8025) );
  NANDN U16183 ( .A(y[1774]), .B(x[1774]), .Z(n18311) );
  NANDN U16184 ( .A(y[1775]), .B(x[1775]), .Z(n8024) );
  NAND U16185 ( .A(n18311), .B(n8024), .Z(n27053) );
  OR U16186 ( .A(n8025), .B(n27053), .Z(n8026) );
  NAND U16187 ( .A(n27054), .B(n8026), .Z(n8027) );
  NANDN U16188 ( .A(n24352), .B(n8027), .Z(n8028) );
  NAND U16189 ( .A(n24351), .B(n8028), .Z(n8029) );
  ANDN U16190 ( .B(x[1779]), .A(y[1779]), .Z(n13294) );
  ANDN U16191 ( .B(n8029), .A(n13294), .Z(n8030) );
  NANDN U16192 ( .A(n13296), .B(n8030), .Z(n8031) );
  NANDN U16193 ( .A(x[1779]), .B(y[1779]), .Z(n24350) );
  AND U16194 ( .A(n8031), .B(n24350), .Z(n8032) );
  NANDN U16195 ( .A(x[1780]), .B(y[1780]), .Z(n18330) );
  NAND U16196 ( .A(n8032), .B(n18330), .Z(n8033) );
  AND U16197 ( .A(n13295), .B(n8033), .Z(n8034) );
  NANDN U16198 ( .A(y[1781]), .B(x[1781]), .Z(n18333) );
  NAND U16199 ( .A(n8034), .B(n18333), .Z(n8035) );
  NANDN U16200 ( .A(n8036), .B(n8035), .Z(n8037) );
  AND U16201 ( .A(n18332), .B(n8037), .Z(n8038) );
  NANDN U16202 ( .A(y[1783]), .B(x[1783]), .Z(n13293) );
  NAND U16203 ( .A(n8038), .B(n13293), .Z(n8039) );
  AND U16204 ( .A(n18335), .B(n8039), .Z(n8040) );
  NANDN U16205 ( .A(n13290), .B(n8040), .Z(n8041) );
  NAND U16206 ( .A(n8042), .B(n8041), .Z(n8043) );
  NANDN U16207 ( .A(x[1785]), .B(y[1785]), .Z(n13291) );
  AND U16208 ( .A(n8043), .B(n13291), .Z(n8044) );
  NAND U16209 ( .A(n13287), .B(n8044), .Z(n8045) );
  NAND U16210 ( .A(n27064), .B(n8045), .Z(n8046) );
  ANDN U16211 ( .B(x[1786]), .A(y[1786]), .Z(n13288) );
  OR U16212 ( .A(n8046), .B(n13288), .Z(n8047) );
  NAND U16213 ( .A(n8048), .B(n8047), .Z(n8049) );
  NANDN U16214 ( .A(n27067), .B(n8049), .Z(n8050) );
  NANDN U16215 ( .A(x[1789]), .B(y[1789]), .Z(n27068) );
  AND U16216 ( .A(n8050), .B(n27068), .Z(n8051) );
  NAND U16217 ( .A(n13284), .B(n8051), .Z(n8052) );
  NAND U16218 ( .A(n27069), .B(n8052), .Z(n8053) );
  ANDN U16219 ( .B(x[1791]), .A(y[1791]), .Z(n13281) );
  OR U16220 ( .A(n8053), .B(n13281), .Z(n8054) );
  AND U16221 ( .A(n13283), .B(n8054), .Z(n8055) );
  NANDN U16222 ( .A(x[1792]), .B(y[1792]), .Z(n13280) );
  AND U16223 ( .A(n8055), .B(n13280), .Z(n8056) );
  NANDN U16224 ( .A(y[1792]), .B(x[1792]), .Z(n13282) );
  NANDN U16225 ( .A(n8056), .B(n13282), .Z(n8057) );
  ANDN U16226 ( .B(x[1793]), .A(y[1793]), .Z(n13277) );
  OR U16227 ( .A(n8057), .B(n13277), .Z(n8058) );
  AND U16228 ( .A(n13279), .B(n8058), .Z(n8059) );
  NANDN U16229 ( .A(x[1794]), .B(y[1794]), .Z(n13276) );
  AND U16230 ( .A(n8059), .B(n13276), .Z(n8060) );
  NANDN U16231 ( .A(y[1794]), .B(x[1794]), .Z(n13278) );
  NANDN U16232 ( .A(n8060), .B(n13278), .Z(n8061) );
  ANDN U16233 ( .B(x[1795]), .A(y[1795]), .Z(n13273) );
  OR U16234 ( .A(n8061), .B(n13273), .Z(n8062) );
  AND U16235 ( .A(n13275), .B(n8062), .Z(n8063) );
  NANDN U16236 ( .A(x[1796]), .B(y[1796]), .Z(n13272) );
  NAND U16237 ( .A(n8063), .B(n13272), .Z(n8064) );
  ANDN U16238 ( .B(x[1797]), .A(y[1797]), .Z(n27077) );
  ANDN U16239 ( .B(n8064), .A(n27077), .Z(n8065) );
  NAND U16240 ( .A(n13274), .B(n8065), .Z(n8066) );
  AND U16241 ( .A(n13271), .B(n8066), .Z(n8067) );
  NANDN U16242 ( .A(x[1798]), .B(y[1798]), .Z(n27078) );
  NAND U16243 ( .A(n8067), .B(n27078), .Z(n8068) );
  NANDN U16244 ( .A(n18359), .B(n8068), .Z(n8069) );
  AND U16245 ( .A(n27079), .B(n8069), .Z(n8072) );
  NANDN U16246 ( .A(y[1801]), .B(x[1801]), .Z(n8071) );
  NANDN U16247 ( .A(y[1800]), .B(x[1800]), .Z(n8070) );
  NAND U16248 ( .A(n8071), .B(n8070), .Z(n27080) );
  OR U16249 ( .A(n8072), .B(n27080), .Z(n8073) );
  AND U16250 ( .A(n13270), .B(n8073), .Z(n8074) );
  NANDN U16251 ( .A(x[1801]), .B(y[1801]), .Z(n27081) );
  NAND U16252 ( .A(n8074), .B(n27081), .Z(n8075) );
  ANDN U16253 ( .B(x[1803]), .A(y[1803]), .Z(n13267) );
  ANDN U16254 ( .B(n8075), .A(n13267), .Z(n8076) );
  NANDN U16255 ( .A(n27083), .B(n8076), .Z(n8077) );
  AND U16256 ( .A(n13269), .B(n8077), .Z(n8078) );
  NANDN U16257 ( .A(x[1804]), .B(y[1804]), .Z(n18367) );
  NAND U16258 ( .A(n8078), .B(n18367), .Z(n8079) );
  NANDN U16259 ( .A(y[1804]), .B(x[1804]), .Z(n13268) );
  AND U16260 ( .A(n8079), .B(n13268), .Z(n8080) );
  NAND U16261 ( .A(n13266), .B(n8080), .Z(n8081) );
  NANDN U16262 ( .A(n18366), .B(n8081), .Z(n8082) );
  ANDN U16263 ( .B(y[1806]), .A(x[1806]), .Z(n13263) );
  OR U16264 ( .A(n8082), .B(n13263), .Z(n8083) );
  NANDN U16265 ( .A(n8084), .B(n8083), .Z(n8085) );
  NANDN U16266 ( .A(x[1808]), .B(y[1808]), .Z(n18372) );
  AND U16267 ( .A(n8085), .B(n18372), .Z(n8086) );
  NANDN U16268 ( .A(x[1807]), .B(y[1807]), .Z(n13264) );
  NAND U16269 ( .A(n8086), .B(n13264), .Z(n8087) );
  ANDN U16270 ( .B(x[1808]), .A(y[1808]), .Z(n13261) );
  ANDN U16271 ( .B(n8087), .A(n13261), .Z(n8088) );
  NANDN U16272 ( .A(n18376), .B(n8088), .Z(n8089) );
  AND U16273 ( .A(n27092), .B(n8089), .Z(n8090) );
  NANDN U16274 ( .A(y[1810]), .B(x[1810]), .Z(n18377) );
  NANDN U16275 ( .A(y[1811]), .B(x[1811]), .Z(n18385) );
  NAND U16276 ( .A(n18377), .B(n18385), .Z(n27093) );
  OR U16277 ( .A(n8090), .B(n27093), .Z(n8091) );
  NANDN U16278 ( .A(x[1811]), .B(y[1811]), .Z(n18382) );
  AND U16279 ( .A(n8091), .B(n18382), .Z(n8092) );
  NANDN U16280 ( .A(x[1812]), .B(y[1812]), .Z(n18388) );
  NAND U16281 ( .A(n8092), .B(n18388), .Z(n8093) );
  ANDN U16282 ( .B(x[1813]), .A(y[1813]), .Z(n18390) );
  ANDN U16283 ( .B(n8093), .A(n18390), .Z(n8094) );
  NANDN U16284 ( .A(n27095), .B(n8094), .Z(n8095) );
  AND U16285 ( .A(n18387), .B(n8095), .Z(n8096) );
  NANDN U16286 ( .A(n13259), .B(n8096), .Z(n8097) );
  NAND U16287 ( .A(n8098), .B(n8097), .Z(n8099) );
  NANDN U16288 ( .A(x[1815]), .B(y[1815]), .Z(n13260) );
  AND U16289 ( .A(n8099), .B(n13260), .Z(n8100) );
  NAND U16290 ( .A(n13256), .B(n8100), .Z(n8101) );
  NANDN U16291 ( .A(n13254), .B(n8101), .Z(n8102) );
  ANDN U16292 ( .B(x[1816]), .A(y[1816]), .Z(n13257) );
  OR U16293 ( .A(n8102), .B(n13257), .Z(n8103) );
  AND U16294 ( .A(n13255), .B(n8103), .Z(n8104) );
  NANDN U16295 ( .A(n24343), .B(n8104), .Z(n8105) );
  NAND U16296 ( .A(n24342), .B(n8105), .Z(n8106) );
  NANDN U16297 ( .A(n27102), .B(n8106), .Z(n8109) );
  NANDN U16298 ( .A(y[1821]), .B(x[1821]), .Z(n8108) );
  NANDN U16299 ( .A(y[1820]), .B(x[1820]), .Z(n8107) );
  AND U16300 ( .A(n8108), .B(n8107), .Z(n27103) );
  AND U16301 ( .A(n8109), .B(n27103), .Z(n8110) );
  ANDN U16302 ( .B(y[1821]), .A(x[1821]), .Z(n18402) );
  ANDN U16303 ( .B(y[1822]), .A(x[1822]), .Z(n18404) );
  NOR U16304 ( .A(n18402), .B(n18404), .Z(n27104) );
  NANDN U16305 ( .A(n8110), .B(n27104), .Z(n8111) );
  NAND U16306 ( .A(n8112), .B(n8111), .Z(n8113) );
  ANDN U16307 ( .B(y[1823]), .A(x[1823]), .Z(n27106) );
  ANDN U16308 ( .B(n8113), .A(n27106), .Z(n8114) );
  NANDN U16309 ( .A(x[1824]), .B(y[1824]), .Z(n13251) );
  NAND U16310 ( .A(n8114), .B(n13251), .Z(n8115) );
  AND U16311 ( .A(n13253), .B(n8115), .Z(n8116) );
  NANDN U16312 ( .A(y[1825]), .B(x[1825]), .Z(n18410) );
  NAND U16313 ( .A(n8116), .B(n18410), .Z(n8117) );
  NANDN U16314 ( .A(x[1826]), .B(y[1826]), .Z(n13249) );
  AND U16315 ( .A(n8117), .B(n13249), .Z(n8118) );
  NANDN U16316 ( .A(n13250), .B(n8118), .Z(n8119) );
  NANDN U16317 ( .A(y[1826]), .B(x[1826]), .Z(n18409) );
  AND U16318 ( .A(n8119), .B(n18409), .Z(n8120) );
  NAND U16319 ( .A(n13247), .B(n8120), .Z(n8121) );
  NANDN U16320 ( .A(n13248), .B(n8121), .Z(n8122) );
  ANDN U16321 ( .B(y[1828]), .A(x[1828]), .Z(n13244) );
  OR U16322 ( .A(n8122), .B(n13244), .Z(n8123) );
  AND U16323 ( .A(n13246), .B(n8123), .Z(n8124) );
  NANDN U16324 ( .A(y[1829]), .B(x[1829]), .Z(n13243) );
  NAND U16325 ( .A(n8124), .B(n13243), .Z(n8125) );
  ANDN U16326 ( .B(y[1830]), .A(x[1830]), .Z(n13241) );
  ANDN U16327 ( .B(n8125), .A(n13241), .Z(n8126) );
  NAND U16328 ( .A(n13245), .B(n8126), .Z(n8127) );
  NANDN U16329 ( .A(y[1831]), .B(x[1831]), .Z(n13240) );
  AND U16330 ( .A(n8127), .B(n13240), .Z(n8128) );
  NANDN U16331 ( .A(n13242), .B(n8128), .Z(n8129) );
  NAND U16332 ( .A(n27117), .B(n8129), .Z(n8130) );
  NANDN U16333 ( .A(n27118), .B(n8130), .Z(n8131) );
  NANDN U16334 ( .A(x[1833]), .B(y[1833]), .Z(n13239) );
  AND U16335 ( .A(n8131), .B(n13239), .Z(n8132) );
  NANDN U16336 ( .A(x[1834]), .B(y[1834]), .Z(n13236) );
  NAND U16337 ( .A(n8132), .B(n13236), .Z(n8133) );
  ANDN U16338 ( .B(x[1835]), .A(y[1835]), .Z(n13233) );
  ANDN U16339 ( .B(n8133), .A(n13233), .Z(n8134) );
  NANDN U16340 ( .A(n13237), .B(n8134), .Z(n8136) );
  NANDN U16341 ( .A(x[1836]), .B(y[1836]), .Z(n13232) );
  NANDN U16342 ( .A(x[1835]), .B(y[1835]), .Z(n13235) );
  AND U16343 ( .A(n13232), .B(n13235), .Z(n8135) );
  NAND U16344 ( .A(n8136), .B(n8135), .Z(n8137) );
  AND U16345 ( .A(n13234), .B(n8137), .Z(n8138) );
  NANDN U16346 ( .A(y[1837]), .B(x[1837]), .Z(n13230) );
  NAND U16347 ( .A(n8138), .B(n13230), .Z(n8139) );
  NANDN U16348 ( .A(x[1838]), .B(y[1838]), .Z(n13228) );
  AND U16349 ( .A(n8139), .B(n13228), .Z(n8140) );
  NANDN U16350 ( .A(n13231), .B(n8140), .Z(n8141) );
  NANDN U16351 ( .A(y[1839]), .B(x[1839]), .Z(n27125) );
  AND U16352 ( .A(n8141), .B(n27125), .Z(n8142) );
  NANDN U16353 ( .A(y[1838]), .B(x[1838]), .Z(n13229) );
  NAND U16354 ( .A(n8142), .B(n13229), .Z(n8143) );
  ANDN U16355 ( .B(y[1839]), .A(x[1839]), .Z(n13227) );
  ANDN U16356 ( .B(n8143), .A(n13227), .Z(n8144) );
  NANDN U16357 ( .A(n18434), .B(n8144), .Z(n8145) );
  NANDN U16358 ( .A(n27127), .B(n8145), .Z(n8146) );
  AND U16359 ( .A(n27129), .B(n8146), .Z(n8147) );
  OR U16360 ( .A(n27131), .B(n8147), .Z(n8148) );
  NAND U16361 ( .A(n27133), .B(n8148), .Z(n8149) );
  NANDN U16362 ( .A(n27135), .B(n8149), .Z(n8150) );
  NANDN U16363 ( .A(y[1845]), .B(x[1845]), .Z(n13224) );
  NANDN U16364 ( .A(n8150), .B(n13224), .Z(n8151) );
  AND U16365 ( .A(n27136), .B(n8151), .Z(n8152) );
  NANDN U16366 ( .A(n13221), .B(n8152), .Z(n8153) );
  NAND U16367 ( .A(n8154), .B(n8153), .Z(n8155) );
  NAND U16368 ( .A(n13222), .B(n8155), .Z(n8156) );
  ANDN U16369 ( .B(y[1848]), .A(x[1848]), .Z(n13219) );
  OR U16370 ( .A(n8156), .B(n13219), .Z(n8157) );
  NAND U16371 ( .A(n8158), .B(n8157), .Z(n8159) );
  AND U16372 ( .A(n13220), .B(n8159), .Z(n8160) );
  NANDN U16373 ( .A(x[1850]), .B(y[1850]), .Z(n13216) );
  NAND U16374 ( .A(n8160), .B(n13216), .Z(n8161) );
  ANDN U16375 ( .B(x[1851]), .A(y[1851]), .Z(n13213) );
  ANDN U16376 ( .B(n8161), .A(n13213), .Z(n8162) );
  ANDN U16377 ( .B(x[1850]), .A(y[1850]), .Z(n13217) );
  ANDN U16378 ( .B(n8162), .A(n13217), .Z(n8164) );
  NANDN U16379 ( .A(x[1852]), .B(y[1852]), .Z(n27152) );
  ANDN U16380 ( .B(y[1851]), .A(x[1851]), .Z(n13215) );
  ANDN U16381 ( .B(n27152), .A(n13215), .Z(n8163) );
  NANDN U16382 ( .A(n8164), .B(n8163), .Z(n8165) );
  ANDN U16383 ( .B(x[1853]), .A(y[1853]), .Z(n27154) );
  ANDN U16384 ( .B(n8165), .A(n27154), .Z(n8166) );
  NANDN U16385 ( .A(y[1852]), .B(x[1852]), .Z(n13214) );
  AND U16386 ( .A(n8166), .B(n13214), .Z(n8167) );
  OR U16387 ( .A(n27156), .B(n8167), .Z(n8168) );
  NAND U16388 ( .A(n27159), .B(n8168), .Z(n8169) );
  NAND U16389 ( .A(n27160), .B(n8169), .Z(n8170) );
  ANDN U16390 ( .B(y[1856]), .A(x[1856]), .Z(n13209) );
  OR U16391 ( .A(n8170), .B(n13209), .Z(n8171) );
  AND U16392 ( .A(n27163), .B(n8171), .Z(n8172) );
  NANDN U16393 ( .A(y[1857]), .B(x[1857]), .Z(n13208) );
  NAND U16394 ( .A(n8172), .B(n13208), .Z(n8173) );
  ANDN U16395 ( .B(y[1858]), .A(x[1858]), .Z(n13205) );
  ANDN U16396 ( .B(n8173), .A(n13205), .Z(n8174) );
  NAND U16397 ( .A(n13210), .B(n8174), .Z(n8175) );
  AND U16398 ( .A(n13207), .B(n8175), .Z(n8176) );
  NANDN U16399 ( .A(y[1859]), .B(x[1859]), .Z(n13204) );
  NAND U16400 ( .A(n8176), .B(n13204), .Z(n8177) );
  NANDN U16401 ( .A(x[1860]), .B(y[1860]), .Z(n13202) );
  AND U16402 ( .A(n8177), .B(n13202), .Z(n8178) );
  NAND U16403 ( .A(n13206), .B(n8178), .Z(n8179) );
  NANDN U16404 ( .A(y[1861]), .B(x[1861]), .Z(n27171) );
  AND U16405 ( .A(n8179), .B(n27171), .Z(n8180) );
  NAND U16406 ( .A(n13203), .B(n8180), .Z(n8181) );
  NANDN U16407 ( .A(n27172), .B(n8181), .Z(n8182) );
  ANDN U16408 ( .B(y[1861]), .A(x[1861]), .Z(n13201) );
  OR U16409 ( .A(n8182), .B(n13201), .Z(n8183) );
  AND U16410 ( .A(n27173), .B(n8183), .Z(n8184) );
  OR U16411 ( .A(n27174), .B(n8184), .Z(n8185) );
  NAND U16412 ( .A(n27175), .B(n8185), .Z(n8186) );
  NANDN U16413 ( .A(n27176), .B(n8186), .Z(n8187) );
  NANDN U16414 ( .A(y[1866]), .B(x[1866]), .Z(n27177) );
  AND U16415 ( .A(n8187), .B(n27177), .Z(n8188) );
  NAND U16416 ( .A(n13200), .B(n8188), .Z(n8189) );
  NANDN U16417 ( .A(n27178), .B(n8189), .Z(n8190) );
  ANDN U16418 ( .B(y[1868]), .A(x[1868]), .Z(n13197) );
  OR U16419 ( .A(n8190), .B(n13197), .Z(n8191) );
  NAND U16420 ( .A(n8192), .B(n8191), .Z(n8193) );
  AND U16421 ( .A(n13198), .B(n8193), .Z(n8194) );
  NANDN U16422 ( .A(n13193), .B(n8194), .Z(n8195) );
  NAND U16423 ( .A(n8196), .B(n8195), .Z(n8197) );
  AND U16424 ( .A(n13194), .B(n8197), .Z(n8198) );
  NANDN U16425 ( .A(x[1872]), .B(y[1872]), .Z(n13190) );
  NAND U16426 ( .A(n8198), .B(n13190), .Z(n8199) );
  ANDN U16427 ( .B(x[1873]), .A(y[1873]), .Z(n13187) );
  ANDN U16428 ( .B(n8199), .A(n13187), .Z(n8200) );
  ANDN U16429 ( .B(x[1872]), .A(y[1872]), .Z(n13191) );
  ANDN U16430 ( .B(n8200), .A(n13191), .Z(n8202) );
  NANDN U16431 ( .A(x[1873]), .B(y[1873]), .Z(n13189) );
  ANDN U16432 ( .B(y[1874]), .A(x[1874]), .Z(n18499) );
  ANDN U16433 ( .B(n13189), .A(n18499), .Z(n8201) );
  NANDN U16434 ( .A(n8202), .B(n8201), .Z(n8203) );
  NANDN U16435 ( .A(y[1875]), .B(x[1875]), .Z(n18505) );
  AND U16436 ( .A(n8203), .B(n18505), .Z(n8204) );
  NANDN U16437 ( .A(y[1874]), .B(x[1874]), .Z(n13188) );
  AND U16438 ( .A(n8204), .B(n13188), .Z(n8205) );
  NANDN U16439 ( .A(x[1875]), .B(y[1875]), .Z(n18500) );
  NANDN U16440 ( .A(x[1876]), .B(y[1876]), .Z(n13186) );
  NAND U16441 ( .A(n18500), .B(n13186), .Z(n27189) );
  OR U16442 ( .A(n8205), .B(n27189), .Z(n8206) );
  NAND U16443 ( .A(n27190), .B(n8206), .Z(n8207) );
  NANDN U16444 ( .A(n13185), .B(n8207), .Z(n8208) );
  ANDN U16445 ( .B(y[1878]), .A(x[1878]), .Z(n18512) );
  OR U16446 ( .A(n8208), .B(n18512), .Z(n8209) );
  NANDN U16447 ( .A(y[1878]), .B(x[1878]), .Z(n27192) );
  NANDN U16448 ( .A(y[1879]), .B(x[1879]), .Z(n13183) );
  ANDN U16449 ( .B(y[1880]), .A(x[1880]), .Z(n13180) );
  NANDN U16450 ( .A(y[1881]), .B(x[1881]), .Z(n13179) );
  NANDN U16451 ( .A(x[1882]), .B(y[1882]), .Z(n13177) );
  NANDN U16452 ( .A(y[1883]), .B(x[1883]), .Z(n27198) );
  NANDN U16453 ( .A(x[1887]), .B(y[1887]), .Z(n18524) );
  NANDN U16454 ( .A(x[1888]), .B(y[1888]), .Z(n18530) );
  NAND U16455 ( .A(n18524), .B(n18530), .Z(n27203) );
  NANDN U16456 ( .A(y[1889]), .B(x[1889]), .Z(n13172) );
  ANDN U16457 ( .B(y[1890]), .A(x[1890]), .Z(n13169) );
  NAND U16458 ( .A(n27205), .B(n8210), .Z(n8211) );
  AND U16459 ( .A(n13171), .B(n8211), .Z(n8212) );
  NANDN U16460 ( .A(y[1891]), .B(x[1891]), .Z(n18535) );
  NAND U16461 ( .A(n8212), .B(n18535), .Z(n8213) );
  AND U16462 ( .A(n13170), .B(n8213), .Z(n8214) );
  NANDN U16463 ( .A(x[1892]), .B(y[1892]), .Z(n13168) );
  NAND U16464 ( .A(n8214), .B(n13168), .Z(n8215) );
  NANDN U16465 ( .A(n8216), .B(n8215), .Z(n8217) );
  AND U16466 ( .A(n13167), .B(n8217), .Z(n8218) );
  NANDN U16467 ( .A(x[1894]), .B(y[1894]), .Z(n13164) );
  NAND U16468 ( .A(n8218), .B(n13164), .Z(n8219) );
  AND U16469 ( .A(n13165), .B(n8219), .Z(n8220) );
  NANDN U16470 ( .A(y[1895]), .B(x[1895]), .Z(n13162) );
  NAND U16471 ( .A(n8220), .B(n13162), .Z(n8221) );
  ANDN U16472 ( .B(y[1896]), .A(x[1896]), .Z(n13159) );
  ANDN U16473 ( .B(n8221), .A(n13159), .Z(n8222) );
  ANDN U16474 ( .B(y[1895]), .A(x[1895]), .Z(n13163) );
  ANDN U16475 ( .B(n8222), .A(n13163), .Z(n8224) );
  ANDN U16476 ( .B(x[1896]), .A(y[1896]), .Z(n13161) );
  ANDN U16477 ( .B(x[1897]), .A(y[1897]), .Z(n27214) );
  NOR U16478 ( .A(n13161), .B(n27214), .Z(n8223) );
  NANDN U16479 ( .A(n8224), .B(n8223), .Z(n8225) );
  AND U16480 ( .A(n27215), .B(n8225), .Z(n8226) );
  NANDN U16481 ( .A(x[1897]), .B(y[1897]), .Z(n13160) );
  AND U16482 ( .A(n8226), .B(n13160), .Z(n8227) );
  OR U16483 ( .A(n27216), .B(n8227), .Z(n8228) );
  AND U16484 ( .A(n8229), .B(n8228), .Z(n8230) );
  NANDN U16485 ( .A(y[1900]), .B(x[1900]), .Z(n27218) );
  ANDN U16486 ( .B(x[1901]), .A(y[1901]), .Z(n24335) );
  ANDN U16487 ( .B(n27218), .A(n24335), .Z(n13157) );
  NANDN U16488 ( .A(n8230), .B(n13157), .Z(n8231) );
  NAND U16489 ( .A(n8232), .B(n8231), .Z(n8233) );
  NANDN U16490 ( .A(n13154), .B(n8233), .Z(n8234) );
  ANDN U16491 ( .B(y[1903]), .A(x[1903]), .Z(n18549) );
  ANDN U16492 ( .B(n8234), .A(n18549), .Z(n8235) );
  NAND U16493 ( .A(n13153), .B(n8235), .Z(n8236) );
  NANDN U16494 ( .A(n13150), .B(n8236), .Z(n8237) );
  ANDN U16495 ( .B(x[1904]), .A(y[1904]), .Z(n13155) );
  OR U16496 ( .A(n8237), .B(n13155), .Z(n8238) );
  AND U16497 ( .A(n8239), .B(n8238), .Z(n8240) );
  ANDN U16498 ( .B(x[1907]), .A(y[1907]), .Z(n13148) );
  NANDN U16499 ( .A(y[1906]), .B(x[1906]), .Z(n13151) );
  NANDN U16500 ( .A(n13148), .B(n13151), .Z(n24332) );
  OR U16501 ( .A(n8240), .B(n24332), .Z(n8241) );
  NAND U16502 ( .A(n27225), .B(n8241), .Z(n8242) );
  NANDN U16503 ( .A(n27226), .B(n8242), .Z(n8243) );
  NANDN U16504 ( .A(n27227), .B(n8243), .Z(n8244) );
  AND U16505 ( .A(n18578), .B(n8244), .Z(n8245) );
  NAND U16506 ( .A(n13147), .B(n8245), .Z(n8246) );
  ANDN U16507 ( .B(y[1912]), .A(x[1912]), .Z(n18580) );
  ANDN U16508 ( .B(n8246), .A(n18580), .Z(n8247) );
  NANDN U16509 ( .A(n27229), .B(n8247), .Z(n8248) );
  AND U16510 ( .A(n18577), .B(n8248), .Z(n8249) );
  NANDN U16511 ( .A(n13145), .B(n8249), .Z(n8250) );
  NAND U16512 ( .A(n8251), .B(n8250), .Z(n8252) );
  AND U16513 ( .A(n13146), .B(n8252), .Z(n8253) );
  ANDN U16514 ( .B(y[1915]), .A(x[1915]), .Z(n13143) );
  OR U16515 ( .A(n8253), .B(n13143), .Z(n8254) );
  NAND U16516 ( .A(n27235), .B(n8254), .Z(n8255) );
  NANDN U16517 ( .A(n18587), .B(n8255), .Z(n8256) );
  NANDN U16518 ( .A(y[1917]), .B(x[1917]), .Z(n13142) );
  NAND U16519 ( .A(n8256), .B(n13142), .Z(n8257) );
  ANDN U16520 ( .B(y[1918]), .A(x[1918]), .Z(n27238) );
  ANDN U16521 ( .B(n8257), .A(n27238), .Z(n8258) );
  NANDN U16522 ( .A(n18586), .B(n8258), .Z(n8259) );
  NANDN U16523 ( .A(y[1919]), .B(x[1919]), .Z(n13139) );
  AND U16524 ( .A(n8259), .B(n13139), .Z(n8260) );
  NANDN U16525 ( .A(y[1918]), .B(x[1918]), .Z(n13141) );
  NAND U16526 ( .A(n8260), .B(n13141), .Z(n8261) );
  NANDN U16527 ( .A(n24330), .B(n8261), .Z(n8262) );
  AND U16528 ( .A(n27240), .B(n8262), .Z(n8264) );
  NANDN U16529 ( .A(x[1922]), .B(y[1922]), .Z(n13137) );
  ANDN U16530 ( .B(y[1921]), .A(x[1921]), .Z(n18595) );
  ANDN U16531 ( .B(n13137), .A(n18595), .Z(n8263) );
  NANDN U16532 ( .A(n8264), .B(n8263), .Z(n8265) );
  NANDN U16533 ( .A(y[1922]), .B(x[1922]), .Z(n18601) );
  AND U16534 ( .A(n8265), .B(n18601), .Z(n8266) );
  NANDN U16535 ( .A(y[1923]), .B(x[1923]), .Z(n18605) );
  AND U16536 ( .A(n8266), .B(n18605), .Z(n8267) );
  NANDN U16537 ( .A(x[1923]), .B(y[1923]), .Z(n13138) );
  NANDN U16538 ( .A(n8267), .B(n13138), .Z(n8268) );
  ANDN U16539 ( .B(y[1924]), .A(x[1924]), .Z(n13135) );
  OR U16540 ( .A(n8268), .B(n13135), .Z(n8269) );
  AND U16541 ( .A(n18604), .B(n8269), .Z(n8270) );
  NANDN U16542 ( .A(y[1925]), .B(x[1925]), .Z(n13134) );
  AND U16543 ( .A(n8270), .B(n13134), .Z(n8271) );
  NANDN U16544 ( .A(x[1925]), .B(y[1925]), .Z(n13136) );
  NANDN U16545 ( .A(n8271), .B(n13136), .Z(n8272) );
  ANDN U16546 ( .B(y[1926]), .A(x[1926]), .Z(n13131) );
  OR U16547 ( .A(n8272), .B(n13131), .Z(n8273) );
  AND U16548 ( .A(n27248), .B(n8273), .Z(n8274) );
  NANDN U16549 ( .A(n13133), .B(n8274), .Z(n8275) );
  AND U16550 ( .A(n8276), .B(n8275), .Z(n8277) );
  NANDN U16551 ( .A(y[1928]), .B(x[1928]), .Z(n13130) );
  NANDN U16552 ( .A(y[1929]), .B(x[1929]), .Z(n13128) );
  NAND U16553 ( .A(n13130), .B(n13128), .Z(n27250) );
  OR U16554 ( .A(n8277), .B(n27250), .Z(n8278) );
  NAND U16555 ( .A(n27251), .B(n8278), .Z(n8279) );
  NANDN U16556 ( .A(n24328), .B(n8279), .Z(n8280) );
  NAND U16557 ( .A(n27252), .B(n8280), .Z(n8281) );
  NANDN U16558 ( .A(y[1933]), .B(x[1933]), .Z(n13124) );
  AND U16559 ( .A(n8281), .B(n13124), .Z(n8282) );
  NANDN U16560 ( .A(n18618), .B(n8282), .Z(n8283) );
  NANDN U16561 ( .A(x[1933]), .B(y[1933]), .Z(n18624) );
  AND U16562 ( .A(n8283), .B(n18624), .Z(n8284) );
  NANDN U16563 ( .A(x[1934]), .B(y[1934]), .Z(n13122) );
  NAND U16564 ( .A(n8284), .B(n13122), .Z(n8285) );
  ANDN U16565 ( .B(x[1935]), .A(y[1935]), .Z(n13119) );
  ANDN U16566 ( .B(n8285), .A(n13119), .Z(n8286) );
  NANDN U16567 ( .A(n13123), .B(n8286), .Z(n8288) );
  NANDN U16568 ( .A(x[1936]), .B(y[1936]), .Z(n13118) );
  NANDN U16569 ( .A(x[1935]), .B(y[1935]), .Z(n13121) );
  AND U16570 ( .A(n13118), .B(n13121), .Z(n8287) );
  NAND U16571 ( .A(n8288), .B(n8287), .Z(n8289) );
  AND U16572 ( .A(n13120), .B(n8289), .Z(n8290) );
  NANDN U16573 ( .A(y[1937]), .B(x[1937]), .Z(n13116) );
  AND U16574 ( .A(n8290), .B(n13116), .Z(n8292) );
  NANDN U16575 ( .A(x[1938]), .B(y[1938]), .Z(n13114) );
  ANDN U16576 ( .B(y[1937]), .A(x[1937]), .Z(n13117) );
  ANDN U16577 ( .B(n13114), .A(n13117), .Z(n8291) );
  NANDN U16578 ( .A(n8292), .B(n8291), .Z(n8293) );
  NANDN U16579 ( .A(n13115), .B(n8293), .Z(n8294) );
  ANDN U16580 ( .B(x[1939]), .A(y[1939]), .Z(n13111) );
  OR U16581 ( .A(n8294), .B(n13111), .Z(n8295) );
  NAND U16582 ( .A(n8296), .B(n8295), .Z(n8297) );
  NANDN U16583 ( .A(n8298), .B(n8297), .Z(n8299) );
  AND U16584 ( .A(n27264), .B(n8299), .Z(n8300) );
  NANDN U16585 ( .A(y[1942]), .B(x[1942]), .Z(n18638) );
  NANDN U16586 ( .A(y[1943]), .B(x[1943]), .Z(n18643) );
  AND U16587 ( .A(n18638), .B(n18643), .Z(n27266) );
  NANDN U16588 ( .A(n8300), .B(n27266), .Z(n8301) );
  NAND U16589 ( .A(n8302), .B(n8301), .Z(n8303) );
  AND U16590 ( .A(n27268), .B(n8303), .Z(n8309) );
  ANDN U16591 ( .B(y[1945]), .A(x[1945]), .Z(n13108) );
  NANDN U16592 ( .A(n8304), .B(n13108), .Z(n8307) );
  NANDN U16593 ( .A(x[1947]), .B(y[1947]), .Z(n8306) );
  NANDN U16594 ( .A(x[1946]), .B(y[1946]), .Z(n8305) );
  AND U16595 ( .A(n8306), .B(n8305), .Z(n13107) );
  AND U16596 ( .A(n8307), .B(n13107), .Z(n8308) );
  NANDN U16597 ( .A(n8309), .B(n8308), .Z(n8310) );
  NAND U16598 ( .A(n27270), .B(n8310), .Z(n8311) );
  NANDN U16599 ( .A(n27271), .B(n8311), .Z(n8312) );
  AND U16600 ( .A(n27272), .B(n8312), .Z(n8315) );
  NANDN U16601 ( .A(x[1950]), .B(y[1950]), .Z(n8314) );
  NANDN U16602 ( .A(x[1951]), .B(y[1951]), .Z(n8313) );
  NAND U16603 ( .A(n8314), .B(n8313), .Z(n27273) );
  OR U16604 ( .A(n8315), .B(n27273), .Z(n8316) );
  NAND U16605 ( .A(n24327), .B(n8316), .Z(n8317) );
  NANDN U16606 ( .A(n27274), .B(n8317), .Z(n8318) );
  NAND U16607 ( .A(n27275), .B(n8318), .Z(n8319) );
  NANDN U16608 ( .A(n27276), .B(n8319), .Z(n8322) );
  NANDN U16609 ( .A(y[1956]), .B(x[1956]), .Z(n8325) );
  NANDN U16610 ( .A(y[1955]), .B(x[1955]), .Z(n8320) );
  AND U16611 ( .A(n8325), .B(n8320), .Z(n13104) );
  NANDN U16612 ( .A(y[1954]), .B(x[1954]), .Z(n8321) );
  AND U16613 ( .A(n13104), .B(n8321), .Z(n27277) );
  AND U16614 ( .A(n8322), .B(n27277), .Z(n8327) );
  NANDN U16615 ( .A(x[1957]), .B(y[1957]), .Z(n8324) );
  NANDN U16616 ( .A(x[1956]), .B(y[1956]), .Z(n8323) );
  NAND U16617 ( .A(n8324), .B(n8323), .Z(n13106) );
  ANDN U16618 ( .B(y[1955]), .A(x[1955]), .Z(n13101) );
  NAND U16619 ( .A(n13101), .B(n8325), .Z(n8326) );
  NANDN U16620 ( .A(n13106), .B(n8326), .Z(n24326) );
  OR U16621 ( .A(n8327), .B(n24326), .Z(n8328) );
  NAND U16622 ( .A(n24325), .B(n8328), .Z(n8329) );
  NANDN U16623 ( .A(n24324), .B(n8329), .Z(n8330) );
  NAND U16624 ( .A(n24323), .B(n8330), .Z(n8331) );
  NAND U16625 ( .A(n27280), .B(n8331), .Z(n8332) );
  NANDN U16626 ( .A(n27281), .B(n8332), .Z(n8333) );
  AND U16627 ( .A(n27282), .B(n8333), .Z(n8334) );
  OR U16628 ( .A(n27283), .B(n8334), .Z(n8335) );
  NAND U16629 ( .A(n27284), .B(n8335), .Z(n8336) );
  NANDN U16630 ( .A(n27285), .B(n8336), .Z(n8337) );
  NANDN U16631 ( .A(n27286), .B(n8337), .Z(n8338) );
  ANDN U16632 ( .B(y[1966]), .A(x[1966]), .Z(n18676) );
  OR U16633 ( .A(n8338), .B(n18676), .Z(n8339) );
  NAND U16634 ( .A(n27287), .B(n8339), .Z(n8340) );
  NANDN U16635 ( .A(n18677), .B(n8340), .Z(n8341) );
  ANDN U16636 ( .B(y[1968]), .A(x[1968]), .Z(n13098) );
  OR U16637 ( .A(n8341), .B(n13098), .Z(n8342) );
  AND U16638 ( .A(n27289), .B(n8342), .Z(n8345) );
  NANDN U16639 ( .A(x[1969]), .B(y[1969]), .Z(n8344) );
  NANDN U16640 ( .A(x[1970]), .B(y[1970]), .Z(n8343) );
  NAND U16641 ( .A(n8344), .B(n8343), .Z(n13099) );
  OR U16642 ( .A(n8345), .B(n13099), .Z(n8348) );
  NANDN U16643 ( .A(y[1971]), .B(x[1971]), .Z(n8347) );
  NANDN U16644 ( .A(y[1970]), .B(x[1970]), .Z(n8346) );
  AND U16645 ( .A(n8347), .B(n8346), .Z(n27291) );
  AND U16646 ( .A(n8348), .B(n27291), .Z(n8351) );
  NANDN U16647 ( .A(x[1971]), .B(y[1971]), .Z(n8350) );
  NANDN U16648 ( .A(x[1972]), .B(y[1972]), .Z(n8349) );
  NAND U16649 ( .A(n8350), .B(n8349), .Z(n24322) );
  OR U16650 ( .A(n8351), .B(n24322), .Z(n8354) );
  NANDN U16651 ( .A(y[1973]), .B(x[1973]), .Z(n8353) );
  NANDN U16652 ( .A(y[1972]), .B(x[1972]), .Z(n8352) );
  AND U16653 ( .A(n8353), .B(n8352), .Z(n24321) );
  AND U16654 ( .A(n8354), .B(n24321), .Z(n8357) );
  NANDN U16655 ( .A(x[1973]), .B(y[1973]), .Z(n8356) );
  NANDN U16656 ( .A(x[1974]), .B(y[1974]), .Z(n8355) );
  NAND U16657 ( .A(n8356), .B(n8355), .Z(n27294) );
  OR U16658 ( .A(n8357), .B(n27294), .Z(n8360) );
  NANDN U16659 ( .A(y[1975]), .B(x[1975]), .Z(n8359) );
  NANDN U16660 ( .A(y[1974]), .B(x[1974]), .Z(n8358) );
  AND U16661 ( .A(n8359), .B(n8358), .Z(n27295) );
  AND U16662 ( .A(n8360), .B(n27295), .Z(n8361) );
  NANDN U16663 ( .A(x[1975]), .B(y[1975]), .Z(n18687) );
  NANDN U16664 ( .A(x[1976]), .B(y[1976]), .Z(n18691) );
  NAND U16665 ( .A(n18687), .B(n18691), .Z(n24320) );
  OR U16666 ( .A(n8361), .B(n24320), .Z(n8362) );
  AND U16667 ( .A(n27296), .B(n8362), .Z(n8364) );
  NANDN U16668 ( .A(x[1978]), .B(y[1978]), .Z(n13095) );
  ANDN U16669 ( .B(y[1977]), .A(x[1977]), .Z(n13096) );
  ANDN U16670 ( .B(n13095), .A(n13096), .Z(n8363) );
  NANDN U16671 ( .A(n8364), .B(n8363), .Z(n8365) );
  NAND U16672 ( .A(n27298), .B(n8365), .Z(n8366) );
  ANDN U16673 ( .B(x[1979]), .A(y[1979]), .Z(n13092) );
  OR U16674 ( .A(n8366), .B(n13092), .Z(n8367) );
  AND U16675 ( .A(n13094), .B(n8367), .Z(n8368) );
  NANDN U16676 ( .A(x[1980]), .B(y[1980]), .Z(n13091) );
  AND U16677 ( .A(n8368), .B(n13091), .Z(n8369) );
  NANDN U16678 ( .A(y[1980]), .B(x[1980]), .Z(n13093) );
  NANDN U16679 ( .A(n8369), .B(n13093), .Z(n8370) );
  NANDN U16680 ( .A(y[1981]), .B(x[1981]), .Z(n13089) );
  NANDN U16681 ( .A(n8370), .B(n13089), .Z(n8371) );
  NANDN U16682 ( .A(x[1982]), .B(y[1982]), .Z(n18700) );
  AND U16683 ( .A(n8371), .B(n18700), .Z(n8372) );
  NANDN U16684 ( .A(x[1981]), .B(y[1981]), .Z(n13090) );
  NAND U16685 ( .A(n8372), .B(n13090), .Z(n8373) );
  ANDN U16686 ( .B(x[1982]), .A(y[1982]), .Z(n13088) );
  ANDN U16687 ( .B(n8373), .A(n13088), .Z(n8374) );
  NANDN U16688 ( .A(n18704), .B(n8374), .Z(n8375) );
  AND U16689 ( .A(n27305), .B(n8375), .Z(n8376) );
  NANDN U16690 ( .A(y[1984]), .B(x[1984]), .Z(n18705) );
  NANDN U16691 ( .A(y[1985]), .B(x[1985]), .Z(n18712) );
  NAND U16692 ( .A(n18705), .B(n18712), .Z(n27306) );
  OR U16693 ( .A(n8376), .B(n27306), .Z(n8377) );
  ANDN U16694 ( .B(y[1985]), .A(x[1985]), .Z(n27307) );
  ANDN U16695 ( .B(n8377), .A(n27307), .Z(n8378) );
  NANDN U16696 ( .A(x[1986]), .B(y[1986]), .Z(n13087) );
  NAND U16697 ( .A(n8378), .B(n13087), .Z(n8379) );
  ANDN U16698 ( .B(x[1987]), .A(y[1987]), .Z(n13084) );
  ANDN U16699 ( .B(n8379), .A(n13084), .Z(n8380) );
  NANDN U16700 ( .A(n27309), .B(n8380), .Z(n8381) );
  NANDN U16701 ( .A(x[1987]), .B(y[1987]), .Z(n13086) );
  AND U16702 ( .A(n8381), .B(n13086), .Z(n8382) );
  NAND U16703 ( .A(n13083), .B(n8382), .Z(n8383) );
  NAND U16704 ( .A(n27313), .B(n8383), .Z(n8384) );
  NANDN U16705 ( .A(y[1988]), .B(x[1988]), .Z(n13085) );
  NANDN U16706 ( .A(n8384), .B(n13085), .Z(n8385) );
  AND U16707 ( .A(n13082), .B(n8385), .Z(n8386) );
  NANDN U16708 ( .A(n18719), .B(n8386), .Z(n8387) );
  AND U16709 ( .A(n27315), .B(n8387), .Z(n8388) );
  NANDN U16710 ( .A(x[1991]), .B(y[1991]), .Z(n18720) );
  NANDN U16711 ( .A(x[1992]), .B(y[1992]), .Z(n13079) );
  NAND U16712 ( .A(n18720), .B(n13079), .Z(n27316) );
  OR U16713 ( .A(n8388), .B(n27316), .Z(n8389) );
  NANDN U16714 ( .A(y[1992]), .B(x[1992]), .Z(n13080) );
  AND U16715 ( .A(n8389), .B(n13080), .Z(n8390) );
  NANDN U16716 ( .A(y[1993]), .B(x[1993]), .Z(n13077) );
  NAND U16717 ( .A(n8390), .B(n13077), .Z(n8391) );
  ANDN U16718 ( .B(y[1994]), .A(x[1994]), .Z(n13074) );
  ANDN U16719 ( .B(n8391), .A(n13074), .Z(n8392) );
  NANDN U16720 ( .A(n13078), .B(n8392), .Z(n8393) );
  NAND U16721 ( .A(n13076), .B(n8393), .Z(n8394) );
  ANDN U16722 ( .B(x[1995]), .A(y[1995]), .Z(n13072) );
  OR U16723 ( .A(n8394), .B(n13072), .Z(n8395) );
  NAND U16724 ( .A(n8396), .B(n8395), .Z(n8397) );
  AND U16725 ( .A(n13073), .B(n8397), .Z(n8398) );
  NANDN U16726 ( .A(n13070), .B(n8398), .Z(n8399) );
  NANDN U16727 ( .A(n24317), .B(n8399), .Z(n8400) );
  NANDN U16728 ( .A(n27324), .B(n8400), .Z(n8401) );
  NANDN U16729 ( .A(y[1998]), .B(x[1998]), .Z(n24318) );
  NANDN U16730 ( .A(n8401), .B(n24318), .Z(n8402) );
  AND U16731 ( .A(n24319), .B(n8402), .Z(n8403) );
  ANDN U16732 ( .B(x[2000]), .A(y[2000]), .Z(n18738) );
  NANDN U16733 ( .A(y[2001]), .B(x[2001]), .Z(n13066) );
  NANDN U16734 ( .A(n18738), .B(n13066), .Z(n27326) );
  OR U16735 ( .A(n8403), .B(n27326), .Z(n8404) );
  AND U16736 ( .A(n27329), .B(n8404), .Z(n8405) );
  NANDN U16737 ( .A(y[2002]), .B(x[2002]), .Z(n13067) );
  NANDN U16738 ( .A(y[2003]), .B(x[2003]), .Z(n18748) );
  NAND U16739 ( .A(n13067), .B(n18748), .Z(n27330) );
  OR U16740 ( .A(n8405), .B(n27330), .Z(n8406) );
  ANDN U16741 ( .B(y[2003]), .A(x[2003]), .Z(n27331) );
  ANDN U16742 ( .B(n8406), .A(n27331), .Z(n8407) );
  NANDN U16743 ( .A(n13064), .B(n8407), .Z(n8409) );
  NANDN U16744 ( .A(y[2005]), .B(x[2005]), .Z(n13063) );
  NANDN U16745 ( .A(y[2004]), .B(x[2004]), .Z(n8408) );
  AND U16746 ( .A(n13063), .B(n8408), .Z(n27332) );
  AND U16747 ( .A(n8409), .B(n27332), .Z(n8412) );
  NANDN U16748 ( .A(x[2005]), .B(y[2005]), .Z(n8411) );
  NANDN U16749 ( .A(x[2006]), .B(y[2006]), .Z(n8410) );
  NAND U16750 ( .A(n8411), .B(n8410), .Z(n13065) );
  OR U16751 ( .A(n8412), .B(n13065), .Z(n8415) );
  NANDN U16752 ( .A(y[2007]), .B(x[2007]), .Z(n8414) );
  NANDN U16753 ( .A(y[2006]), .B(x[2006]), .Z(n8413) );
  AND U16754 ( .A(n8414), .B(n8413), .Z(n24316) );
  AND U16755 ( .A(n8415), .B(n24316), .Z(n8418) );
  NANDN U16756 ( .A(x[2007]), .B(y[2007]), .Z(n8417) );
  NANDN U16757 ( .A(x[2008]), .B(y[2008]), .Z(n8416) );
  NAND U16758 ( .A(n8417), .B(n8416), .Z(n24315) );
  OR U16759 ( .A(n8418), .B(n24315), .Z(n8419) );
  AND U16760 ( .A(n27334), .B(n8419), .Z(n8421) );
  ANDN U16761 ( .B(y[2010]), .A(x[2010]), .Z(n18756) );
  ANDN U16762 ( .B(y[2009]), .A(x[2009]), .Z(n27335) );
  NOR U16763 ( .A(n18756), .B(n27335), .Z(n8420) );
  NANDN U16764 ( .A(n8421), .B(n8420), .Z(n8422) );
  AND U16765 ( .A(n27336), .B(n8422), .Z(n8425) );
  NANDN U16766 ( .A(x[2011]), .B(y[2011]), .Z(n8424) );
  NANDN U16767 ( .A(x[2012]), .B(y[2012]), .Z(n8423) );
  NAND U16768 ( .A(n8424), .B(n8423), .Z(n18758) );
  OR U16769 ( .A(n8425), .B(n18758), .Z(n8426) );
  NAND U16770 ( .A(n13062), .B(n8426), .Z(n8427) );
  NANDN U16771 ( .A(n8428), .B(n8427), .Z(n8429) );
  NANDN U16772 ( .A(y[2014]), .B(x[2014]), .Z(n18762) );
  AND U16773 ( .A(n8429), .B(n18762), .Z(n8430) );
  NAND U16774 ( .A(n13059), .B(n8430), .Z(n8431) );
  NANDN U16775 ( .A(n13060), .B(n8431), .Z(n8432) );
  NANDN U16776 ( .A(x[2016]), .B(y[2016]), .Z(n13057) );
  NANDN U16777 ( .A(n8432), .B(n13057), .Z(n8433) );
  AND U16778 ( .A(n13058), .B(n8433), .Z(n8434) );
  NANDN U16779 ( .A(y[2017]), .B(x[2017]), .Z(n13055) );
  NAND U16780 ( .A(n8434), .B(n13055), .Z(n8435) );
  ANDN U16781 ( .B(y[2018]), .A(x[2018]), .Z(n13052) );
  ANDN U16782 ( .B(n8435), .A(n13052), .Z(n8436) );
  NANDN U16783 ( .A(n13056), .B(n8436), .Z(n8437) );
  AND U16784 ( .A(n13054), .B(n8437), .Z(n8438) );
  NANDN U16785 ( .A(y[2019]), .B(x[2019]), .Z(n13051) );
  NAND U16786 ( .A(n8438), .B(n13051), .Z(n8439) );
  NANDN U16787 ( .A(n27350), .B(n8439), .Z(n8440) );
  NANDN U16788 ( .A(y[2020]), .B(x[2020]), .Z(n27349) );
  AND U16789 ( .A(n8440), .B(n27349), .Z(n8441) );
  NANDN U16790 ( .A(y[2021]), .B(x[2021]), .Z(n13048) );
  NAND U16791 ( .A(n8441), .B(n13048), .Z(n8442) );
  ANDN U16792 ( .B(y[2021]), .A(x[2021]), .Z(n13049) );
  ANDN U16793 ( .B(n8442), .A(n13049), .Z(n8443) );
  NANDN U16794 ( .A(n13047), .B(n8443), .Z(n8444) );
  NANDN U16795 ( .A(y[2023]), .B(x[2023]), .Z(n18779) );
  AND U16796 ( .A(n8444), .B(n18779), .Z(n8446) );
  NANDN U16797 ( .A(y[2022]), .B(x[2022]), .Z(n8445) );
  NAND U16798 ( .A(n8446), .B(n8445), .Z(n8447) );
  NANDN U16799 ( .A(n27354), .B(n8447), .Z(n8448) );
  AND U16800 ( .A(n27355), .B(n8448), .Z(n8449) );
  NANDN U16801 ( .A(x[2025]), .B(y[2025]), .Z(n13045) );
  NANDN U16802 ( .A(x[2026]), .B(y[2026]), .Z(n13043) );
  NAND U16803 ( .A(n13045), .B(n13043), .Z(n24314) );
  OR U16804 ( .A(n8449), .B(n24314), .Z(n8450) );
  NAND U16805 ( .A(n27356), .B(n8450), .Z(n8451) );
  NANDN U16806 ( .A(n27357), .B(n8451), .Z(n8452) );
  NANDN U16807 ( .A(n27358), .B(n8452), .Z(n8453) );
  AND U16808 ( .A(n27359), .B(n8453), .Z(n8456) );
  NANDN U16809 ( .A(y[2030]), .B(x[2030]), .Z(n8455) );
  NANDN U16810 ( .A(y[2031]), .B(x[2031]), .Z(n8454) );
  NAND U16811 ( .A(n8455), .B(n8454), .Z(n13038) );
  OR U16812 ( .A(n8456), .B(n13038), .Z(n8459) );
  NANDN U16813 ( .A(x[2032]), .B(y[2032]), .Z(n8458) );
  NANDN U16814 ( .A(x[2031]), .B(y[2031]), .Z(n8457) );
  AND U16815 ( .A(n8458), .B(n8457), .Z(n18795) );
  AND U16816 ( .A(n8459), .B(n18795), .Z(n8462) );
  NANDN U16817 ( .A(y[2032]), .B(x[2032]), .Z(n8461) );
  NANDN U16818 ( .A(y[2033]), .B(x[2033]), .Z(n8460) );
  NAND U16819 ( .A(n8461), .B(n8460), .Z(n13035) );
  OR U16820 ( .A(n8462), .B(n13035), .Z(n8465) );
  NANDN U16821 ( .A(x[2034]), .B(y[2034]), .Z(n8464) );
  NANDN U16822 ( .A(x[2033]), .B(y[2033]), .Z(n8463) );
  AND U16823 ( .A(n8464), .B(n8463), .Z(n13034) );
  AND U16824 ( .A(n8465), .B(n13034), .Z(n8466) );
  NANDN U16825 ( .A(y[2034]), .B(x[2034]), .Z(n18799) );
  NANDN U16826 ( .A(y[2035]), .B(x[2035]), .Z(n18805) );
  NAND U16827 ( .A(n18799), .B(n18805), .Z(n27365) );
  OR U16828 ( .A(n8466), .B(n27365), .Z(n8467) );
  AND U16829 ( .A(n27366), .B(n8467), .Z(n8468) );
  NANDN U16830 ( .A(y[2036]), .B(x[2036]), .Z(n18804) );
  NANDN U16831 ( .A(y[2037]), .B(x[2037]), .Z(n13033) );
  NAND U16832 ( .A(n18804), .B(n13033), .Z(n24313) );
  OR U16833 ( .A(n8468), .B(n24313), .Z(n8469) );
  NAND U16834 ( .A(n27367), .B(n8469), .Z(n8470) );
  NAND U16835 ( .A(n27368), .B(n8470), .Z(n8471) );
  ANDN U16836 ( .B(x[2039]), .A(y[2039]), .Z(n13030) );
  OR U16837 ( .A(n8471), .B(n13030), .Z(n8472) );
  NAND U16838 ( .A(n8473), .B(n8472), .Z(n8474) );
  NANDN U16839 ( .A(y[2041]), .B(x[2041]), .Z(n27372) );
  AND U16840 ( .A(n8474), .B(n27372), .Z(n8476) );
  NANDN U16841 ( .A(y[2040]), .B(x[2040]), .Z(n8475) );
  AND U16842 ( .A(n8476), .B(n8475), .Z(n8477) );
  ANDN U16843 ( .B(y[2041]), .A(x[2041]), .Z(n18817) );
  NANDN U16844 ( .A(x[2042]), .B(y[2042]), .Z(n13029) );
  NANDN U16845 ( .A(n18817), .B(n13029), .Z(n24312) );
  OR U16846 ( .A(n8477), .B(n24312), .Z(n8478) );
  NANDN U16847 ( .A(y[2042]), .B(x[2042]), .Z(n24311) );
  AND U16848 ( .A(n8478), .B(n24311), .Z(n8479) );
  NANDN U16849 ( .A(y[2043]), .B(x[2043]), .Z(n13027) );
  NAND U16850 ( .A(n8479), .B(n13027), .Z(n8480) );
  ANDN U16851 ( .B(y[2043]), .A(x[2043]), .Z(n13028) );
  ANDN U16852 ( .B(n8480), .A(n13028), .Z(n8481) );
  NANDN U16853 ( .A(n13026), .B(n8481), .Z(n8482) );
  NANDN U16854 ( .A(y[2045]), .B(x[2045]), .Z(n27378) );
  AND U16855 ( .A(n8482), .B(n27378), .Z(n8484) );
  NANDN U16856 ( .A(y[2044]), .B(x[2044]), .Z(n8483) );
  AND U16857 ( .A(n8484), .B(n8483), .Z(n8485) );
  ANDN U16858 ( .B(y[2045]), .A(x[2045]), .Z(n18825) );
  ANDN U16859 ( .B(y[2046]), .A(x[2046]), .Z(n18831) );
  OR U16860 ( .A(n18825), .B(n18831), .Z(n27379) );
  OR U16861 ( .A(n8485), .B(n27379), .Z(n8486) );
  NAND U16862 ( .A(n27380), .B(n8486), .Z(n8487) );
  NANDN U16863 ( .A(n27381), .B(n8487), .Z(n8488) );
  ANDN U16864 ( .B(y[2048]), .A(x[2048]), .Z(n13023) );
  OR U16865 ( .A(n8488), .B(n13023), .Z(n8489) );
  NAND U16866 ( .A(n8490), .B(n8489), .Z(n8491) );
  AND U16867 ( .A(n27385), .B(n8491), .Z(n8492) );
  NANDN U16868 ( .A(x[2049]), .B(y[2049]), .Z(n13024) );
  NAND U16869 ( .A(n8492), .B(n13024), .Z(n8493) );
  NANDN U16870 ( .A(n27386), .B(n8493), .Z(n8494) );
  AND U16871 ( .A(n27388), .B(n8494), .Z(n8495) );
  ANDN U16872 ( .B(x[2052]), .A(y[2052]), .Z(n18842) );
  NANDN U16873 ( .A(y[2053]), .B(x[2053]), .Z(n13021) );
  NANDN U16874 ( .A(n18842), .B(n13021), .Z(n27389) );
  OR U16875 ( .A(n8495), .B(n27389), .Z(n8496) );
  ANDN U16876 ( .B(y[2053]), .A(x[2053]), .Z(n27390) );
  ANDN U16877 ( .B(n8496), .A(n27390), .Z(n8497) );
  NANDN U16878 ( .A(x[2054]), .B(y[2054]), .Z(n18851) );
  NAND U16879 ( .A(n8497), .B(n18851), .Z(n8498) );
  NANDN U16880 ( .A(y[2055]), .B(x[2055]), .Z(n27393) );
  AND U16881 ( .A(n8498), .B(n27393), .Z(n8499) );
  NAND U16882 ( .A(n27391), .B(n8499), .Z(n8500) );
  AND U16883 ( .A(n18850), .B(n8500), .Z(n8501) );
  NANDN U16884 ( .A(x[2056]), .B(y[2056]), .Z(n13019) );
  NAND U16885 ( .A(n8501), .B(n13019), .Z(n8502) );
  NANDN U16886 ( .A(n24308), .B(n8502), .Z(n8503) );
  AND U16887 ( .A(n24309), .B(n8503), .Z(n8504) );
  NANDN U16888 ( .A(x[2058]), .B(y[2058]), .Z(n13017) );
  NAND U16889 ( .A(n8504), .B(n13017), .Z(n8505) );
  NANDN U16890 ( .A(y[2059]), .B(x[2059]), .Z(n13015) );
  AND U16891 ( .A(n8505), .B(n13015), .Z(n8506) );
  NAND U16892 ( .A(n27394), .B(n8506), .Z(n8507) );
  AND U16893 ( .A(n13016), .B(n8507), .Z(n8508) );
  NANDN U16894 ( .A(x[2060]), .B(y[2060]), .Z(n18861) );
  NAND U16895 ( .A(n8508), .B(n18861), .Z(n8509) );
  NANDN U16896 ( .A(y[2061]), .B(x[2061]), .Z(n13013) );
  AND U16897 ( .A(n8509), .B(n13013), .Z(n8510) );
  NANDN U16898 ( .A(n13014), .B(n8510), .Z(n8511) );
  NANDN U16899 ( .A(x[2062]), .B(y[2062]), .Z(n27398) );
  AND U16900 ( .A(n8511), .B(n27398), .Z(n8512) );
  NAND U16901 ( .A(n18860), .B(n8512), .Z(n8513) );
  NANDN U16902 ( .A(n13012), .B(n8513), .Z(n8514) );
  ANDN U16903 ( .B(x[2063]), .A(y[2063]), .Z(n13010) );
  OR U16904 ( .A(n8514), .B(n13010), .Z(n8515) );
  NANDN U16905 ( .A(x[2063]), .B(y[2063]), .Z(n13011) );
  NANDN U16906 ( .A(x[2064]), .B(y[2064]), .Z(n13009) );
  AND U16907 ( .A(n13011), .B(n13009), .Z(n27402) );
  AND U16908 ( .A(n8515), .B(n27402), .Z(n8517) );
  NANDN U16909 ( .A(y[2064]), .B(x[2064]), .Z(n27403) );
  ANDN U16910 ( .B(x[2065]), .A(y[2065]), .Z(n13007) );
  ANDN U16911 ( .B(n27403), .A(n13007), .Z(n8516) );
  NANDN U16912 ( .A(n8517), .B(n8516), .Z(n8518) );
  NAND U16913 ( .A(n27401), .B(n8518), .Z(n8519) );
  XNOR U16914 ( .A(x[2066]), .B(y[2066]), .Z(n13008) );
  NANDN U16915 ( .A(n8519), .B(n13008), .Z(n8520) );
  NAND U16916 ( .A(n8521), .B(n8520), .Z(n8522) );
  NANDN U16917 ( .A(n24305), .B(n8522), .Z(n8523) );
  NANDN U16918 ( .A(y[2068]), .B(x[2068]), .Z(n24306) );
  AND U16919 ( .A(n8523), .B(n24306), .Z(n8524) );
  NAND U16920 ( .A(n13005), .B(n8524), .Z(n8525) );
  NANDN U16921 ( .A(n27408), .B(n8525), .Z(n8526) );
  XOR U16922 ( .A(x[2070]), .B(y[2070]), .Z(n13004) );
  OR U16923 ( .A(n8526), .B(n13004), .Z(n8527) );
  NANDN U16924 ( .A(y[2071]), .B(x[2071]), .Z(n24304) );
  AND U16925 ( .A(n8527), .B(n24304), .Z(n8528) );
  NANDN U16926 ( .A(n8529), .B(n8528), .Z(n8530) );
  AND U16927 ( .A(n8531), .B(n8530), .Z(n8532) );
  OR U16928 ( .A(n27412), .B(n8532), .Z(n8533) );
  NAND U16929 ( .A(n27413), .B(n8533), .Z(n8534) );
  NANDN U16930 ( .A(n27414), .B(n8534), .Z(n8536) );
  NANDN U16931 ( .A(x[2076]), .B(y[2076]), .Z(n12999) );
  NANDN U16932 ( .A(x[2075]), .B(y[2075]), .Z(n27415) );
  AND U16933 ( .A(n12999), .B(n27415), .Z(n8535) );
  NAND U16934 ( .A(n8536), .B(n8535), .Z(n8538) );
  NANDN U16935 ( .A(y[2076]), .B(x[2076]), .Z(n8537) );
  NANDN U16936 ( .A(y[2077]), .B(x[2077]), .Z(n12998) );
  AND U16937 ( .A(n8537), .B(n12998), .Z(n18893) );
  AND U16938 ( .A(n8538), .B(n18893), .Z(n8541) );
  NANDN U16939 ( .A(x[2077]), .B(y[2077]), .Z(n8540) );
  NANDN U16940 ( .A(x[2078]), .B(y[2078]), .Z(n8539) );
  NAND U16941 ( .A(n8540), .B(n8539), .Z(n13000) );
  OR U16942 ( .A(n8541), .B(n13000), .Z(n8544) );
  NANDN U16943 ( .A(y[2079]), .B(x[2079]), .Z(n8543) );
  NANDN U16944 ( .A(y[2078]), .B(x[2078]), .Z(n8542) );
  AND U16945 ( .A(n8543), .B(n8542), .Z(n12997) );
  AND U16946 ( .A(n8544), .B(n12997), .Z(n8547) );
  NANDN U16947 ( .A(x[2079]), .B(y[2079]), .Z(n8546) );
  NANDN U16948 ( .A(x[2080]), .B(y[2080]), .Z(n8545) );
  NAND U16949 ( .A(n8546), .B(n8545), .Z(n12996) );
  OR U16950 ( .A(n8547), .B(n12996), .Z(n8550) );
  NANDN U16951 ( .A(y[2081]), .B(x[2081]), .Z(n8549) );
  NANDN U16952 ( .A(y[2080]), .B(x[2080]), .Z(n8548) );
  AND U16953 ( .A(n8549), .B(n8548), .Z(n27421) );
  AND U16954 ( .A(n8550), .B(n27421), .Z(n8553) );
  NANDN U16955 ( .A(x[2081]), .B(y[2081]), .Z(n8552) );
  NANDN U16956 ( .A(x[2082]), .B(y[2082]), .Z(n8551) );
  NAND U16957 ( .A(n8552), .B(n8551), .Z(n24303) );
  OR U16958 ( .A(n8553), .B(n24303), .Z(n8556) );
  NANDN U16959 ( .A(y[2083]), .B(x[2083]), .Z(n8555) );
  NANDN U16960 ( .A(y[2082]), .B(x[2082]), .Z(n8554) );
  AND U16961 ( .A(n8555), .B(n8554), .Z(n24302) );
  AND U16962 ( .A(n8556), .B(n24302), .Z(n8559) );
  NANDN U16963 ( .A(x[2083]), .B(y[2083]), .Z(n8558) );
  NANDN U16964 ( .A(x[2084]), .B(y[2084]), .Z(n8557) );
  NAND U16965 ( .A(n8558), .B(n8557), .Z(n27422) );
  OR U16966 ( .A(n8559), .B(n27422), .Z(n8560) );
  NANDN U16967 ( .A(y[2084]), .B(x[2084]), .Z(n18903) );
  NANDN U16968 ( .A(y[2085]), .B(x[2085]), .Z(n12995) );
  AND U16969 ( .A(n18903), .B(n12995), .Z(n27423) );
  AND U16970 ( .A(n8560), .B(n27423), .Z(n8561) );
  ANDN U16971 ( .B(y[2085]), .A(x[2085]), .Z(n18905) );
  NANDN U16972 ( .A(x[2086]), .B(y[2086]), .Z(n12994) );
  NANDN U16973 ( .A(n18905), .B(n12994), .Z(n24301) );
  OR U16974 ( .A(n8561), .B(n24301), .Z(n8562) );
  NANDN U16975 ( .A(y[2086]), .B(x[2086]), .Z(n24300) );
  AND U16976 ( .A(n8562), .B(n24300), .Z(n8563) );
  NANDN U16977 ( .A(y[2087]), .B(x[2087]), .Z(n12991) );
  AND U16978 ( .A(n8563), .B(n12991), .Z(n8565) );
  NANDN U16979 ( .A(x[2088]), .B(y[2088]), .Z(n12993) );
  NANDN U16980 ( .A(x[2087]), .B(y[2087]), .Z(n8564) );
  AND U16981 ( .A(n12993), .B(n8564), .Z(n27424) );
  NANDN U16982 ( .A(n8565), .B(n27424), .Z(n8566) );
  NANDN U16983 ( .A(y[2088]), .B(x[2088]), .Z(n12992) );
  AND U16984 ( .A(n8566), .B(n12992), .Z(n8567) );
  NANDN U16985 ( .A(n12990), .B(n8567), .Z(n8568) );
  NAND U16986 ( .A(n27428), .B(n8568), .Z(n8569) );
  NANDN U16987 ( .A(n12989), .B(n8569), .Z(n8570) );
  NANDN U16988 ( .A(y[2091]), .B(x[2091]), .Z(n12987) );
  NANDN U16989 ( .A(n8570), .B(n12987), .Z(n8571) );
  AND U16990 ( .A(n8572), .B(n8571), .Z(n8574) );
  NANDN U16991 ( .A(y[2093]), .B(x[2093]), .Z(n27433) );
  ANDN U16992 ( .B(x[2092]), .A(y[2092]), .Z(n12986) );
  ANDN U16993 ( .B(n27433), .A(n12986), .Z(n8573) );
  NANDN U16994 ( .A(n8574), .B(n8573), .Z(n8575) );
  NANDN U16995 ( .A(n24299), .B(n8575), .Z(n8576) );
  ANDN U16996 ( .B(y[2093]), .A(x[2093]), .Z(n12984) );
  OR U16997 ( .A(n8576), .B(n12984), .Z(n8577) );
  NAND U16998 ( .A(n24298), .B(n8577), .Z(n8578) );
  NANDN U16999 ( .A(n27434), .B(n8578), .Z(n8579) );
  NAND U17000 ( .A(n27435), .B(n8579), .Z(n8580) );
  ANDN U17001 ( .B(y[2098]), .A(x[2098]), .Z(n12981) );
  ANDN U17002 ( .B(n8580), .A(n12981), .Z(n8581) );
  NANDN U17003 ( .A(n24297), .B(n8581), .Z(n8582) );
  NANDN U17004 ( .A(y[2098]), .B(x[2098]), .Z(n24296) );
  AND U17005 ( .A(n8582), .B(n24296), .Z(n8583) );
  NANDN U17006 ( .A(y[2099]), .B(x[2099]), .Z(n18935) );
  NAND U17007 ( .A(n8583), .B(n18935), .Z(n8584) );
  AND U17008 ( .A(n12982), .B(n8584), .Z(n8585) );
  NANDN U17009 ( .A(n12978), .B(n8585), .Z(n8586) );
  NAND U17010 ( .A(n18936), .B(n8586), .Z(n8587) );
  NANDN U17011 ( .A(n12977), .B(n8587), .Z(n8588) );
  ANDN U17012 ( .B(y[2102]), .A(x[2102]), .Z(n12976) );
  OR U17013 ( .A(n8588), .B(n12976), .Z(n8589) );
  NANDN U17014 ( .A(y[2102]), .B(x[2102]), .Z(n27440) );
  AND U17015 ( .A(n8589), .B(n27440), .Z(n8590) );
  NANDN U17016 ( .A(y[2103]), .B(x[2103]), .Z(n18942) );
  NAND U17017 ( .A(n8590), .B(n18942), .Z(n8591) );
  ANDN U17018 ( .B(y[2104]), .A(x[2104]), .Z(n18945) );
  ANDN U17019 ( .B(n8591), .A(n18945), .Z(n8592) );
  NANDN U17020 ( .A(n12975), .B(n8592), .Z(n8593) );
  NANDN U17021 ( .A(y[2104]), .B(x[2104]), .Z(n18941) );
  AND U17022 ( .A(n8593), .B(n18941), .Z(n8594) );
  NAND U17023 ( .A(n12974), .B(n8594), .Z(n8595) );
  NAND U17024 ( .A(n27444), .B(n8595), .Z(n8596) );
  ANDN U17025 ( .B(y[2105]), .A(x[2105]), .Z(n18944) );
  OR U17026 ( .A(n8596), .B(n18944), .Z(n8597) );
  NAND U17027 ( .A(n8598), .B(n8597), .Z(n8599) );
  NANDN U17028 ( .A(n27446), .B(n8599), .Z(n8600) );
  AND U17029 ( .A(n27447), .B(n8600), .Z(n8601) );
  NAND U17030 ( .A(n12970), .B(n8601), .Z(n8602) );
  NAND U17031 ( .A(n27448), .B(n8602), .Z(n8603) );
  NANDN U17032 ( .A(n12969), .B(n8603), .Z(n8604) );
  ANDN U17033 ( .B(x[2111]), .A(y[2111]), .Z(n12967) );
  OR U17034 ( .A(n8604), .B(n12967), .Z(n8605) );
  AND U17035 ( .A(n27450), .B(n8605), .Z(n8606) );
  OR U17036 ( .A(n27451), .B(n8606), .Z(n8607) );
  NAND U17037 ( .A(n8608), .B(n8607), .Z(n8609) );
  NANDN U17038 ( .A(n8610), .B(n8609), .Z(n8611) );
  AND U17039 ( .A(n12964), .B(n8611), .Z(n8612) );
  NANDN U17040 ( .A(n27458), .B(n8612), .Z(n8613) );
  NAND U17041 ( .A(n27459), .B(n8613), .Z(n8614) );
  NANDN U17042 ( .A(n27460), .B(n8614), .Z(n8615) );
  NANDN U17043 ( .A(y[2118]), .B(x[2118]), .Z(n18972) );
  NANDN U17044 ( .A(y[2119]), .B(x[2119]), .Z(n12962) );
  AND U17045 ( .A(n18972), .B(n12962), .Z(n27461) );
  AND U17046 ( .A(n8615), .B(n27461), .Z(n8617) );
  NANDN U17047 ( .A(x[2120]), .B(y[2120]), .Z(n12960) );
  ANDN U17048 ( .B(y[2119]), .A(x[2119]), .Z(n24291) );
  ANDN U17049 ( .B(n12960), .A(n24291), .Z(n8616) );
  NANDN U17050 ( .A(n8617), .B(n8616), .Z(n8618) );
  NAND U17051 ( .A(n27464), .B(n8618), .Z(n8619) );
  NANDN U17052 ( .A(y[2120]), .B(x[2120]), .Z(n27462) );
  NANDN U17053 ( .A(n8619), .B(n27462), .Z(n8620) );
  AND U17054 ( .A(n8621), .B(n8620), .Z(n8622) );
  NANDN U17055 ( .A(y[2122]), .B(x[2122]), .Z(n18980) );
  NANDN U17056 ( .A(y[2123]), .B(x[2123]), .Z(n12959) );
  NAND U17057 ( .A(n18980), .B(n12959), .Z(n27466) );
  OR U17058 ( .A(n8622), .B(n27466), .Z(n8623) );
  ANDN U17059 ( .B(y[2123]), .A(x[2123]), .Z(n27467) );
  ANDN U17060 ( .B(n8623), .A(n27467), .Z(n8624) );
  NANDN U17061 ( .A(x[2124]), .B(y[2124]), .Z(n18988) );
  NAND U17062 ( .A(n8624), .B(n18988), .Z(n8625) );
  NANDN U17063 ( .A(y[2125]), .B(x[2125]), .Z(n12958) );
  AND U17064 ( .A(n8625), .B(n12958), .Z(n8626) );
  NAND U17065 ( .A(n27468), .B(n8626), .Z(n8627) );
  AND U17066 ( .A(n18987), .B(n8627), .Z(n8628) );
  NANDN U17067 ( .A(x[2126]), .B(y[2126]), .Z(n12956) );
  NAND U17068 ( .A(n8628), .B(n12956), .Z(n8629) );
  NANDN U17069 ( .A(y[2127]), .B(x[2127]), .Z(n12954) );
  AND U17070 ( .A(n8629), .B(n12954), .Z(n8630) );
  NANDN U17071 ( .A(n12957), .B(n8630), .Z(n8631) );
  ANDN U17072 ( .B(y[2128]), .A(x[2128]), .Z(n27474) );
  ANDN U17073 ( .B(n8631), .A(n27474), .Z(n8632) );
  NAND U17074 ( .A(n12955), .B(n8632), .Z(n8633) );
  NANDN U17075 ( .A(y[2129]), .B(x[2129]), .Z(n8635) );
  AND U17076 ( .A(n8635), .B(n8634), .Z(n27475) );
  NANDN U17077 ( .A(y[2134]), .B(x[2134]), .Z(n12950) );
  NANDN U17078 ( .A(y[2135]), .B(x[2135]), .Z(n19010) );
  NAND U17079 ( .A(n12950), .B(n19010), .Z(n27481) );
  ANDN U17080 ( .B(y[2136]), .A(x[2136]), .Z(n19009) );
  NANDN U17081 ( .A(x[2135]), .B(y[2135]), .Z(n8636) );
  NANDN U17082 ( .A(n19009), .B(n8636), .Z(n19006) );
  IV U17083 ( .A(n19006), .Z(n27482) );
  NANDN U17084 ( .A(y[2136]), .B(x[2136]), .Z(n12949) );
  NANDN U17085 ( .A(x[2137]), .B(y[2137]), .Z(n27485) );
  NANDN U17086 ( .A(y[2137]), .B(x[2137]), .Z(n12948) );
  ANDN U17087 ( .B(x[2138]), .A(y[2138]), .Z(n12947) );
  NANDN U17088 ( .A(y[2139]), .B(x[2139]), .Z(n27486) );
  NANDN U17089 ( .A(y[2141]), .B(x[2141]), .Z(n12944) );
  NANDN U17090 ( .A(x[2141]), .B(y[2141]), .Z(n27489) );
  ANDN U17091 ( .B(y[2142]), .A(x[2142]), .Z(n12941) );
  ANDN U17092 ( .B(n27489), .A(n12941), .Z(n8637) );
  NANDN U17093 ( .A(n8638), .B(n8637), .Z(n8639) );
  NAND U17094 ( .A(n12943), .B(n8639), .Z(n8640) );
  AND U17095 ( .A(n12940), .B(n8640), .Z(n8643) );
  NANDN U17096 ( .A(y[2144]), .B(x[2144]), .Z(n8642) );
  NANDN U17097 ( .A(y[2145]), .B(x[2145]), .Z(n8641) );
  NAND U17098 ( .A(n8642), .B(n8641), .Z(n12936) );
  OR U17099 ( .A(n8643), .B(n12936), .Z(n8644) );
  NAND U17100 ( .A(n8645), .B(n8644), .Z(n8646) );
  NANDN U17101 ( .A(y[2146]), .B(x[2146]), .Z(n12938) );
  AND U17102 ( .A(n8646), .B(n12938), .Z(n8647) );
  NAND U17103 ( .A(n19027), .B(n8647), .Z(n8648) );
  NANDN U17104 ( .A(n12934), .B(n8648), .Z(n8649) );
  ANDN U17105 ( .B(y[2148]), .A(x[2148]), .Z(n19030) );
  OR U17106 ( .A(n8649), .B(n19030), .Z(n8650) );
  AND U17107 ( .A(n19026), .B(n8650), .Z(n8651) );
  NANDN U17108 ( .A(y[2149]), .B(x[2149]), .Z(n12933) );
  NAND U17109 ( .A(n8651), .B(n12933), .Z(n8652) );
  NANDN U17110 ( .A(x[2150]), .B(y[2150]), .Z(n27497) );
  AND U17111 ( .A(n8652), .B(n27497), .Z(n8653) );
  NANDN U17112 ( .A(n19029), .B(n8653), .Z(n8654) );
  AND U17113 ( .A(n12932), .B(n8654), .Z(n8655) );
  NANDN U17114 ( .A(n12930), .B(n8655), .Z(n8656) );
  NAND U17115 ( .A(n27499), .B(n8656), .Z(n8657) );
  NANDN U17116 ( .A(n12931), .B(n8657), .Z(n8658) );
  ANDN U17117 ( .B(x[2153]), .A(y[2153]), .Z(n12928) );
  OR U17118 ( .A(n8658), .B(n12928), .Z(n8659) );
  AND U17119 ( .A(n27501), .B(n8659), .Z(n8660) );
  OR U17120 ( .A(n8661), .B(n8660), .Z(n8662) );
  NAND U17121 ( .A(n27504), .B(n8662), .Z(n8663) );
  NANDN U17122 ( .A(n27505), .B(n8663), .Z(n8664) );
  AND U17123 ( .A(n27506), .B(n8664), .Z(n8665) );
  XNOR U17124 ( .A(x[2158]), .B(y[2158]), .Z(n27507) );
  NANDN U17125 ( .A(n8665), .B(n27507), .Z(n8666) );
  NAND U17126 ( .A(n27508), .B(n8666), .Z(n8667) );
  NANDN U17127 ( .A(n27509), .B(n8667), .Z(n8668) );
  AND U17128 ( .A(n27510), .B(n8668), .Z(n8674) );
  ANDN U17129 ( .B(x[2161]), .A(y[2161]), .Z(n12925) );
  ANDN U17130 ( .B(x[2160]), .A(y[2160]), .Z(n19055) );
  OR U17131 ( .A(n12925), .B(n19055), .Z(n8669) );
  NAND U17132 ( .A(n8670), .B(n8669), .Z(n8673) );
  NANDN U17133 ( .A(y[2162]), .B(x[2162]), .Z(n8672) );
  NANDN U17134 ( .A(y[2163]), .B(x[2163]), .Z(n8671) );
  NAND U17135 ( .A(n8672), .B(n8671), .Z(n19061) );
  ANDN U17136 ( .B(n8673), .A(n19061), .Z(n27511) );
  NANDN U17137 ( .A(n8674), .B(n27511), .Z(n8675) );
  NAND U17138 ( .A(n8676), .B(n8675), .Z(n8678) );
  ANDN U17139 ( .B(x[2164]), .A(y[2164]), .Z(n27513) );
  ANDN U17140 ( .B(x[2165]), .A(y[2165]), .Z(n27515) );
  NOR U17141 ( .A(n27513), .B(n27515), .Z(n8677) );
  NAND U17142 ( .A(n8678), .B(n8677), .Z(n8679) );
  NANDN U17143 ( .A(x[2166]), .B(y[2166]), .Z(n27516) );
  AND U17144 ( .A(n8679), .B(n27516), .Z(n8680) );
  NANDN U17145 ( .A(x[2165]), .B(y[2165]), .Z(n12923) );
  NAND U17146 ( .A(n8680), .B(n12923), .Z(n8681) );
  NANDN U17147 ( .A(n27517), .B(n8681), .Z(n8682) );
  NANDN U17148 ( .A(x[2167]), .B(y[2167]), .Z(n12921) );
  NANDN U17149 ( .A(x[2168]), .B(y[2168]), .Z(n19073) );
  AND U17150 ( .A(n12921), .B(n19073), .Z(n27518) );
  AND U17151 ( .A(n8682), .B(n27518), .Z(n8683) );
  NANDN U17152 ( .A(y[2168]), .B(x[2168]), .Z(n12919) );
  NANDN U17153 ( .A(y[2169]), .B(x[2169]), .Z(n12918) );
  NAND U17154 ( .A(n12919), .B(n12918), .Z(n24286) );
  OR U17155 ( .A(n8683), .B(n24286), .Z(n8684) );
  NANDN U17156 ( .A(x[2169]), .B(y[2169]), .Z(n19072) );
  NANDN U17157 ( .A(x[2170]), .B(y[2170]), .Z(n19079) );
  AND U17158 ( .A(n19072), .B(n19079), .Z(n24285) );
  AND U17159 ( .A(n8684), .B(n24285), .Z(n8685) );
  NANDN U17160 ( .A(y[2170]), .B(x[2170]), .Z(n12917) );
  NANDN U17161 ( .A(y[2171]), .B(x[2171]), .Z(n12916) );
  NAND U17162 ( .A(n12917), .B(n12916), .Z(n27520) );
  OR U17163 ( .A(n8685), .B(n27520), .Z(n8686) );
  NAND U17164 ( .A(n27521), .B(n8686), .Z(n8687) );
  NANDN U17165 ( .A(n24284), .B(n8687), .Z(n8688) );
  NAND U17166 ( .A(n27522), .B(n8688), .Z(n8689) );
  NANDN U17167 ( .A(y[2175]), .B(x[2175]), .Z(n12914) );
  AND U17168 ( .A(n8689), .B(n12914), .Z(n8690) );
  NANDN U17169 ( .A(n19088), .B(n8690), .Z(n8691) );
  AND U17170 ( .A(n8692), .B(n8691), .Z(n8694) );
  NANDN U17171 ( .A(y[2177]), .B(x[2177]), .Z(n27527) );
  ANDN U17172 ( .B(x[2176]), .A(y[2176]), .Z(n12913) );
  ANDN U17173 ( .B(n27527), .A(n12913), .Z(n8693) );
  NANDN U17174 ( .A(n8694), .B(n8693), .Z(n8695) );
  NANDN U17175 ( .A(n24283), .B(n8695), .Z(n8696) );
  NAND U17176 ( .A(n24282), .B(n8696), .Z(n8697) );
  NAND U17177 ( .A(n12909), .B(n8697), .Z(n8698) );
  ANDN U17178 ( .B(y[2179]), .A(x[2179]), .Z(n12910) );
  OR U17179 ( .A(n8698), .B(n12910), .Z(n8700) );
  NANDN U17180 ( .A(y[2181]), .B(x[2181]), .Z(n19106) );
  NANDN U17181 ( .A(y[2180]), .B(x[2180]), .Z(n8699) );
  AND U17182 ( .A(n19106), .B(n8699), .Z(n27530) );
  AND U17183 ( .A(n8700), .B(n27530), .Z(n8703) );
  NANDN U17184 ( .A(x[2182]), .B(y[2182]), .Z(n8702) );
  NANDN U17185 ( .A(x[2181]), .B(y[2181]), .Z(n8701) );
  NAND U17186 ( .A(n8702), .B(n8701), .Z(n12906) );
  OR U17187 ( .A(n8703), .B(n12906), .Z(n8706) );
  NANDN U17188 ( .A(y[2182]), .B(x[2182]), .Z(n8705) );
  NANDN U17189 ( .A(y[2183]), .B(x[2183]), .Z(n8704) );
  NAND U17190 ( .A(n8705), .B(n8704), .Z(n19111) );
  ANDN U17191 ( .B(n8706), .A(n19111), .Z(n8707) );
  OR U17192 ( .A(n8708), .B(n8707), .Z(n8709) );
  NAND U17193 ( .A(n24281), .B(n8709), .Z(n8710) );
  NANDN U17194 ( .A(n12903), .B(n8710), .Z(n8711) );
  ANDN U17195 ( .B(y[2186]), .A(x[2186]), .Z(n19118) );
  OR U17196 ( .A(n8711), .B(n19118), .Z(n8712) );
  AND U17197 ( .A(n27536), .B(n8712), .Z(n8714) );
  NANDN U17198 ( .A(x[2187]), .B(y[2187]), .Z(n19119) );
  ANDN U17199 ( .B(y[2188]), .A(x[2188]), .Z(n24280) );
  ANDN U17200 ( .B(n19119), .A(n24280), .Z(n8713) );
  NANDN U17201 ( .A(n8714), .B(n8713), .Z(n8715) );
  NANDN U17202 ( .A(n27537), .B(n8715), .Z(n8716) );
  AND U17203 ( .A(n27538), .B(n8716), .Z(n8717) );
  OR U17204 ( .A(n27539), .B(n8717), .Z(n8718) );
  NAND U17205 ( .A(n24277), .B(n8718), .Z(n8719) );
  NANDN U17206 ( .A(n27540), .B(n8719), .Z(n8720) );
  NANDN U17207 ( .A(n27542), .B(n8720), .Z(n8721) );
  AND U17208 ( .A(n27543), .B(n8721), .Z(n8722) );
  NANDN U17209 ( .A(x[2195]), .B(y[2195]), .Z(n12894) );
  NANDN U17210 ( .A(x[2196]), .B(y[2196]), .Z(n19148) );
  NAND U17211 ( .A(n12894), .B(n19148), .Z(n27544) );
  OR U17212 ( .A(n8722), .B(n27544), .Z(n8723) );
  ANDN U17213 ( .B(x[2196]), .A(y[2196]), .Z(n27545) );
  ANDN U17214 ( .B(n8723), .A(n27545), .Z(n8724) );
  NANDN U17215 ( .A(y[2197]), .B(x[2197]), .Z(n19150) );
  AND U17216 ( .A(n8724), .B(n19150), .Z(n8726) );
  NANDN U17217 ( .A(x[2198]), .B(y[2198]), .Z(n19151) );
  NANDN U17218 ( .A(x[2197]), .B(y[2197]), .Z(n8725) );
  AND U17219 ( .A(n19151), .B(n8725), .Z(n27546) );
  NANDN U17220 ( .A(n8726), .B(n27546), .Z(n8727) );
  NANDN U17221 ( .A(n19153), .B(n8727), .Z(n8728) );
  NANDN U17222 ( .A(n12891), .B(n8728), .Z(n8729) );
  NANDN U17223 ( .A(y[2200]), .B(x[2200]), .Z(n12890) );
  AND U17224 ( .A(n8729), .B(n12890), .Z(n8730) );
  NANDN U17225 ( .A(y[2201]), .B(x[2201]), .Z(n12889) );
  NAND U17226 ( .A(n8730), .B(n12889), .Z(n8731) );
  AND U17227 ( .A(n12893), .B(n8731), .Z(n8732) );
  NANDN U17228 ( .A(n12886), .B(n8732), .Z(n8733) );
  AND U17229 ( .A(n8734), .B(n8733), .Z(n8735) );
  ANDN U17230 ( .B(n24275), .A(n8735), .Z(n8738) );
  NANDN U17231 ( .A(x[2203]), .B(y[2203]), .Z(n12887) );
  OR U17232 ( .A(n12887), .B(n8736), .Z(n8737) );
  AND U17233 ( .A(n8738), .B(n8737), .Z(n8739) );
  ANDN U17234 ( .B(x[2205]), .A(y[2205]), .Z(n27551) );
  OR U17235 ( .A(n8739), .B(n27551), .Z(n8740) );
  AND U17236 ( .A(n12885), .B(n8740), .Z(n8741) );
  ANDN U17237 ( .B(x[2206]), .A(y[2206]), .Z(n19162) );
  NANDN U17238 ( .A(y[2207]), .B(x[2207]), .Z(n12884) );
  NANDN U17239 ( .A(n19162), .B(n12884), .Z(n27556) );
  OR U17240 ( .A(n8741), .B(n27556), .Z(n8742) );
  AND U17241 ( .A(n27555), .B(n8742), .Z(n8743) );
  NANDN U17242 ( .A(x[2208]), .B(y[2208]), .Z(n12883) );
  AND U17243 ( .A(n8743), .B(n12883), .Z(n8745) );
  NANDN U17244 ( .A(y[2208]), .B(x[2208]), .Z(n8744) );
  NANDN U17245 ( .A(y[2209]), .B(x[2209]), .Z(n12882) );
  AND U17246 ( .A(n8744), .B(n12882), .Z(n27554) );
  NANDN U17247 ( .A(n8745), .B(n27554), .Z(n8746) );
  NANDN U17248 ( .A(n12880), .B(n8746), .Z(n8749) );
  NANDN U17249 ( .A(y[2210]), .B(x[2210]), .Z(n8748) );
  NANDN U17250 ( .A(y[2211]), .B(x[2211]), .Z(n8747) );
  NAND U17251 ( .A(n8748), .B(n8747), .Z(n12878) );
  ANDN U17252 ( .B(n8749), .A(n12878), .Z(n8751) );
  NANDN U17253 ( .A(x[2211]), .B(y[2211]), .Z(n12881) );
  ANDN U17254 ( .B(y[2212]), .A(x[2212]), .Z(n12876) );
  ANDN U17255 ( .B(n12881), .A(n12876), .Z(n8750) );
  NANDN U17256 ( .A(n8751), .B(n8750), .Z(n8752) );
  NANDN U17257 ( .A(n12879), .B(n8752), .Z(n8753) );
  NANDN U17258 ( .A(y[2213]), .B(x[2213]), .Z(n12875) );
  NANDN U17259 ( .A(n8753), .B(n12875), .Z(n8754) );
  AND U17260 ( .A(n12877), .B(n8754), .Z(n8755) );
  NANDN U17261 ( .A(x[2214]), .B(y[2214]), .Z(n19172) );
  AND U17262 ( .A(n8755), .B(n19172), .Z(n8756) );
  NANDN U17263 ( .A(x[2215]), .B(y[2215]), .Z(n19171) );
  ANDN U17264 ( .B(x[2219]), .A(y[2219]), .Z(n19180) );
  NANDN U17265 ( .A(x[2220]), .B(y[2220]), .Z(n27566) );
  NANDN U17266 ( .A(x[2219]), .B(y[2219]), .Z(n19177) );
  ANDN U17267 ( .B(x[2225]), .A(y[2225]), .Z(n12869) );
  AND U17268 ( .A(n8759), .B(n8758), .Z(n8760) );
  ANDN U17269 ( .B(x[2227]), .A(y[2227]), .Z(n12864) );
  ANDN U17270 ( .B(x[2226]), .A(y[2226]), .Z(n19191) );
  OR U17271 ( .A(n12864), .B(n19191), .Z(n27574) );
  OR U17272 ( .A(n8760), .B(n27574), .Z(n8761) );
  NAND U17273 ( .A(n27575), .B(n8761), .Z(n8762) );
  NANDN U17274 ( .A(n24272), .B(n8762), .Z(n8763) );
  NANDN U17275 ( .A(x[2230]), .B(y[2230]), .Z(n12861) );
  AND U17276 ( .A(n8763), .B(n12861), .Z(n8764) );
  NAND U17277 ( .A(n24271), .B(n8764), .Z(n8765) );
  NAND U17278 ( .A(n27576), .B(n8765), .Z(n8766) );
  AND U17279 ( .A(n12859), .B(n8766), .Z(n8769) );
  NANDN U17280 ( .A(y[2232]), .B(x[2232]), .Z(n8768) );
  NANDN U17281 ( .A(y[2233]), .B(x[2233]), .Z(n8767) );
  NAND U17282 ( .A(n8768), .B(n8767), .Z(n12855) );
  OR U17283 ( .A(n8769), .B(n12855), .Z(n8770) );
  NAND U17284 ( .A(n8771), .B(n8770), .Z(n8772) );
  NANDN U17285 ( .A(y[2234]), .B(x[2234]), .Z(n12857) );
  AND U17286 ( .A(n8772), .B(n12857), .Z(n8773) );
  NAND U17287 ( .A(n19203), .B(n8773), .Z(n8774) );
  NANDN U17288 ( .A(n12853), .B(n8774), .Z(n8775) );
  NANDN U17289 ( .A(x[2236]), .B(y[2236]), .Z(n12852) );
  NANDN U17290 ( .A(n8775), .B(n12852), .Z(n8776) );
  AND U17291 ( .A(n19202), .B(n8776), .Z(n8777) );
  NANDN U17292 ( .A(y[2237]), .B(x[2237]), .Z(n19207) );
  NAND U17293 ( .A(n8777), .B(n19207), .Z(n8778) );
  NANDN U17294 ( .A(x[2238]), .B(y[2238]), .Z(n27583) );
  AND U17295 ( .A(n8778), .B(n27583), .Z(n8779) );
  NANDN U17296 ( .A(n12851), .B(n8779), .Z(n8780) );
  AND U17297 ( .A(n19206), .B(n8780), .Z(n8781) );
  NAND U17298 ( .A(n27584), .B(n8781), .Z(n8788) );
  NANDN U17299 ( .A(x[2241]), .B(y[2241]), .Z(n8783) );
  NANDN U17300 ( .A(x[2240]), .B(y[2240]), .Z(n8782) );
  AND U17301 ( .A(n8783), .B(n8782), .Z(n8785) );
  NANDN U17302 ( .A(x[2242]), .B(y[2242]), .Z(n8784) );
  AND U17303 ( .A(n8785), .B(n8784), .Z(n19214) );
  NANDN U17304 ( .A(x[2239]), .B(y[2239]), .Z(n12850) );
  OR U17305 ( .A(n8786), .B(n12850), .Z(n8787) );
  AND U17306 ( .A(n19214), .B(n8787), .Z(n27586) );
  AND U17307 ( .A(n8788), .B(n27586), .Z(n8795) );
  NANDN U17308 ( .A(y[2242]), .B(x[2242]), .Z(n8790) );
  ANDN U17309 ( .B(x[2243]), .A(y[2243]), .Z(n8789) );
  ANDN U17310 ( .B(n8790), .A(n8789), .Z(n8794) );
  XNOR U17311 ( .A(x[2242]), .B(y[2242]), .Z(n8792) );
  ANDN U17312 ( .B(x[2241]), .A(y[2241]), .Z(n8791) );
  NAND U17313 ( .A(n8792), .B(n8791), .Z(n8793) );
  AND U17314 ( .A(n8794), .B(n8793), .Z(n12849) );
  NANDN U17315 ( .A(n8795), .B(n12849), .Z(n8796) );
  NANDN U17316 ( .A(n19216), .B(n8796), .Z(n8797) );
  NANDN U17317 ( .A(n19217), .B(n8797), .Z(n8798) );
  NANDN U17318 ( .A(y[2245]), .B(x[2245]), .Z(n12848) );
  NANDN U17319 ( .A(n8798), .B(n12848), .Z(n8799) );
  AND U17320 ( .A(n19219), .B(n8799), .Z(n8800) );
  NANDN U17321 ( .A(x[2246]), .B(y[2246]), .Z(n12846) );
  NAND U17322 ( .A(n8800), .B(n12846), .Z(n8801) );
  ANDN U17323 ( .B(x[2247]), .A(y[2247]), .Z(n19223) );
  ANDN U17324 ( .B(n8801), .A(n19223), .Z(n8802) );
  NANDN U17325 ( .A(n12847), .B(n8802), .Z(n8803) );
  NANDN U17326 ( .A(x[2248]), .B(y[2248]), .Z(n12844) );
  AND U17327 ( .A(n8803), .B(n12844), .Z(n8804) );
  NANDN U17328 ( .A(n12845), .B(n8804), .Z(n8805) );
  NAND U17329 ( .A(n24270), .B(n8805), .Z(n8806) );
  NANDN U17330 ( .A(n27593), .B(n8806), .Z(n8807) );
  AND U17331 ( .A(n27594), .B(n8807), .Z(n8808) );
  ANDN U17332 ( .B(y[2251]), .A(x[2251]), .Z(n27595) );
  OR U17333 ( .A(n8808), .B(n27595), .Z(n8809) );
  ANDN U17334 ( .B(y[2252]), .A(x[2252]), .Z(n19238) );
  OR U17335 ( .A(n8809), .B(n19238), .Z(n8810) );
  AND U17336 ( .A(n27596), .B(n8810), .Z(n8813) );
  NANDN U17337 ( .A(x[2253]), .B(y[2253]), .Z(n8812) );
  NANDN U17338 ( .A(x[2254]), .B(y[2254]), .Z(n8811) );
  NAND U17339 ( .A(n8812), .B(n8811), .Z(n19236) );
  OR U17340 ( .A(n8813), .B(n19236), .Z(n8814) );
  NANDN U17341 ( .A(n12839), .B(n8814), .Z(n8815) );
  NANDN U17342 ( .A(n8816), .B(n8815), .Z(n8817) );
  NANDN U17343 ( .A(y[2256]), .B(x[2256]), .Z(n12840) );
  AND U17344 ( .A(n8817), .B(n12840), .Z(n8818) );
  NAND U17345 ( .A(n12836), .B(n8818), .Z(n8819) );
  NANDN U17346 ( .A(n12837), .B(n8819), .Z(n8820) );
  ANDN U17347 ( .B(y[2258]), .A(x[2258]), .Z(n12833) );
  OR U17348 ( .A(n8820), .B(n12833), .Z(n8821) );
  AND U17349 ( .A(n12835), .B(n8821), .Z(n8822) );
  NANDN U17350 ( .A(y[2259]), .B(x[2259]), .Z(n12832) );
  NAND U17351 ( .A(n8822), .B(n12832), .Z(n8823) );
  ANDN U17352 ( .B(y[2260]), .A(x[2260]), .Z(n12829) );
  ANDN U17353 ( .B(n8823), .A(n12829), .Z(n8824) );
  NAND U17354 ( .A(n12834), .B(n8824), .Z(n8827) );
  NANDN U17355 ( .A(y[2261]), .B(x[2261]), .Z(n8825) );
  AND U17356 ( .A(n8826), .B(n8825), .Z(n27604) );
  AND U17357 ( .A(n8827), .B(n27604), .Z(n8828) );
  NAND U17358 ( .A(n12831), .B(n8828), .Z(n8829) );
  NANDN U17359 ( .A(n24268), .B(n8829), .Z(n8830) );
  NAND U17360 ( .A(n12828), .B(n8830), .Z(n8831) );
  NAND U17361 ( .A(n27606), .B(n8831), .Z(n8832) );
  NAND U17362 ( .A(n27607), .B(n8832), .Z(n8833) );
  NAND U17363 ( .A(n27608), .B(n8833), .Z(n8834) );
  NANDN U17364 ( .A(n27609), .B(n8834), .Z(n8835) );
  AND U17365 ( .A(n27610), .B(n8835), .Z(n8836) );
  NANDN U17366 ( .A(y[2269]), .B(x[2269]), .Z(n27611) );
  NANDN U17367 ( .A(n8836), .B(n27611), .Z(n8837) );
  AND U17368 ( .A(n27612), .B(n8837), .Z(n8838) );
  OR U17369 ( .A(n27613), .B(n8838), .Z(n8839) );
  NAND U17370 ( .A(n8840), .B(n8839), .Z(n8842) );
  NANDN U17371 ( .A(y[2275]), .B(x[2275]), .Z(n19266) );
  NANDN U17372 ( .A(y[2274]), .B(x[2274]), .Z(n8841) );
  AND U17373 ( .A(n19266), .B(n8841), .Z(n27615) );
  AND U17374 ( .A(n8842), .B(n27615), .Z(n8845) );
  NANDN U17375 ( .A(x[2275]), .B(y[2275]), .Z(n8844) );
  NANDN U17376 ( .A(x[2276]), .B(y[2276]), .Z(n8843) );
  NAND U17377 ( .A(n8844), .B(n8843), .Z(n19268) );
  OR U17378 ( .A(n8845), .B(n19268), .Z(n8846) );
  NAND U17379 ( .A(n24267), .B(n8846), .Z(n8847) );
  NANDN U17380 ( .A(n27618), .B(n8847), .Z(n8848) );
  AND U17381 ( .A(n27619), .B(n8848), .Z(n8849) );
  NANDN U17382 ( .A(x[2279]), .B(y[2279]), .Z(n19275) );
  NANDN U17383 ( .A(x[2280]), .B(y[2280]), .Z(n12817) );
  NAND U17384 ( .A(n19275), .B(n12817), .Z(n24266) );
  OR U17385 ( .A(n8849), .B(n24266), .Z(n8850) );
  AND U17386 ( .A(n8851), .B(n8850), .Z(n8852) );
  ANDN U17387 ( .B(y[2282]), .A(x[2282]), .Z(n24265) );
  NANDN U17388 ( .A(x[2281]), .B(y[2281]), .Z(n12818) );
  NANDN U17389 ( .A(n24265), .B(n12818), .Z(n27621) );
  OR U17390 ( .A(n8852), .B(n27621), .Z(n8853) );
  AND U17391 ( .A(n19281), .B(n8853), .Z(n8854) );
  NANDN U17392 ( .A(y[2283]), .B(x[2283]), .Z(n19286) );
  NAND U17393 ( .A(n8854), .B(n19286), .Z(n8855) );
  ANDN U17394 ( .B(y[2284]), .A(x[2284]), .Z(n19288) );
  ANDN U17395 ( .B(n8855), .A(n19288), .Z(n8856) );
  NAND U17396 ( .A(n27623), .B(n8856), .Z(n8857) );
  AND U17397 ( .A(n27622), .B(n8857), .Z(n8858) );
  NANDN U17398 ( .A(n12815), .B(n8858), .Z(n8859) );
  NAND U17399 ( .A(n8860), .B(n8859), .Z(n8861) );
  NANDN U17400 ( .A(y[2287]), .B(x[2287]), .Z(n27627) );
  NANDN U17401 ( .A(y[2286]), .B(x[2286]), .Z(n12816) );
  NANDN U17402 ( .A(y[2288]), .B(x[2288]), .Z(n27631) );
  NANDN U17403 ( .A(y[2289]), .B(x[2289]), .Z(n12813) );
  ANDN U17404 ( .B(y[2289]), .A(x[2289]), .Z(n27632) );
  NANDN U17405 ( .A(x[2295]), .B(y[2295]), .Z(n27640) );
  ANDN U17406 ( .B(y[2296]), .A(x[2296]), .Z(n19319) );
  NANDN U17407 ( .A(y[2298]), .B(x[2298]), .Z(n8863) );
  NANDN U17408 ( .A(y[2299]), .B(x[2299]), .Z(n8862) );
  NAND U17409 ( .A(n8863), .B(n8862), .Z(n12807) );
  NAND U17410 ( .A(n8865), .B(n8864), .Z(n8866) );
  AND U17411 ( .A(n12809), .B(n8866), .Z(n8867) );
  NANDN U17412 ( .A(y[2301]), .B(x[2301]), .Z(n12803) );
  NAND U17413 ( .A(n8867), .B(n12803), .Z(n8868) );
  AND U17414 ( .A(n12805), .B(n8868), .Z(n8869) );
  NAND U17415 ( .A(n12801), .B(n8869), .Z(n8870) );
  NAND U17416 ( .A(n8871), .B(n8870), .Z(n8872) );
  NANDN U17417 ( .A(n12796), .B(n8872), .Z(n8873) );
  ANDN U17418 ( .B(y[2303]), .A(x[2303]), .Z(n12800) );
  OR U17419 ( .A(n8873), .B(n12800), .Z(n8874) );
  AND U17420 ( .A(n12798), .B(n8874), .Z(n8875) );
  NAND U17421 ( .A(n24262), .B(n8875), .Z(n8876) );
  NANDN U17422 ( .A(n24261), .B(n8876), .Z(n8878) );
  NANDN U17423 ( .A(y[2308]), .B(x[2308]), .Z(n8879) );
  NANDN U17424 ( .A(y[2307]), .B(x[2307]), .Z(n8877) );
  AND U17425 ( .A(n8879), .B(n8877), .Z(n19334) );
  NANDN U17426 ( .A(y[2306]), .B(x[2306]), .Z(n12795) );
  AND U17427 ( .A(n19334), .B(n12795), .Z(n24260) );
  AND U17428 ( .A(n8878), .B(n24260), .Z(n8881) );
  NANDN U17429 ( .A(x[2307]), .B(y[2307]), .Z(n12793) );
  NANDN U17430 ( .A(n12793), .B(n8879), .Z(n8880) );
  ANDN U17431 ( .B(y[2308]), .A(x[2308]), .Z(n19338) );
  ANDN U17432 ( .B(n8880), .A(n19338), .Z(n27651) );
  NANDN U17433 ( .A(n8881), .B(n27651), .Z(n8883) );
  NANDN U17434 ( .A(y[2310]), .B(x[2310]), .Z(n8886) );
  NANDN U17435 ( .A(y[2309]), .B(x[2309]), .Z(n8882) );
  AND U17436 ( .A(n8886), .B(n8882), .Z(n27652) );
  AND U17437 ( .A(n8883), .B(n27652), .Z(n8888) );
  NANDN U17438 ( .A(x[2311]), .B(y[2311]), .Z(n8885) );
  NANDN U17439 ( .A(x[2310]), .B(y[2310]), .Z(n8884) );
  NAND U17440 ( .A(n8885), .B(n8884), .Z(n19340) );
  ANDN U17441 ( .B(y[2309]), .A(x[2309]), .Z(n19336) );
  NAND U17442 ( .A(n19336), .B(n8886), .Z(n8887) );
  NANDN U17443 ( .A(n19340), .B(n8887), .Z(n24259) );
  OR U17444 ( .A(n8888), .B(n24259), .Z(n8889) );
  NAND U17445 ( .A(n24258), .B(n8889), .Z(n8890) );
  NANDN U17446 ( .A(n19344), .B(n8890), .Z(n8891) );
  NANDN U17447 ( .A(y[2313]), .B(x[2313]), .Z(n27654) );
  NAND U17448 ( .A(n8891), .B(n27654), .Z(n8892) );
  ANDN U17449 ( .B(y[2313]), .A(x[2313]), .Z(n19343) );
  ANDN U17450 ( .B(n8892), .A(n19343), .Z(n8893) );
  NANDN U17451 ( .A(n27655), .B(n8893), .Z(n8894) );
  AND U17452 ( .A(n27656), .B(n8894), .Z(n8895) );
  OR U17453 ( .A(n27657), .B(n8895), .Z(n8896) );
  NAND U17454 ( .A(n27659), .B(n8896), .Z(n8897) );
  NANDN U17455 ( .A(n27660), .B(n8897), .Z(n8898) );
  ANDN U17456 ( .B(y[2318]), .A(x[2318]), .Z(n12791) );
  OR U17457 ( .A(n8898), .B(n12791), .Z(n8900) );
  NANDN U17458 ( .A(y[2318]), .B(x[2318]), .Z(n8899) );
  NANDN U17459 ( .A(y[2319]), .B(x[2319]), .Z(n12790) );
  AND U17460 ( .A(n8899), .B(n12790), .Z(n27661) );
  AND U17461 ( .A(n8900), .B(n27661), .Z(n8903) );
  NANDN U17462 ( .A(x[2319]), .B(y[2319]), .Z(n8902) );
  NANDN U17463 ( .A(x[2320]), .B(y[2320]), .Z(n8901) );
  NAND U17464 ( .A(n8902), .B(n8901), .Z(n12792) );
  OR U17465 ( .A(n8903), .B(n12792), .Z(n8904) );
  AND U17466 ( .A(n27663), .B(n8904), .Z(n8905) );
  OR U17467 ( .A(n27664), .B(n8905), .Z(n8906) );
  NAND U17468 ( .A(n27665), .B(n8906), .Z(n8907) );
  NANDN U17469 ( .A(n27666), .B(n8907), .Z(n8908) );
  NANDN U17470 ( .A(y[2325]), .B(x[2325]), .Z(n19374) );
  AND U17471 ( .A(n8908), .B(n19374), .Z(n8909) );
  NAND U17472 ( .A(n27667), .B(n8909), .Z(n8910) );
  NANDN U17473 ( .A(n12783), .B(n8910), .Z(n8911) );
  AND U17474 ( .A(n19376), .B(n8911), .Z(n8912) );
  NANDN U17475 ( .A(x[2327]), .B(y[2327]), .Z(n19379) );
  NANDN U17476 ( .A(x[2328]), .B(y[2328]), .Z(n19381) );
  AND U17477 ( .A(n19379), .B(n19381), .Z(n24256) );
  NANDN U17478 ( .A(n8912), .B(n24256), .Z(n8913) );
  NAND U17479 ( .A(n8914), .B(n8913), .Z(n8915) );
  NANDN U17480 ( .A(x[2329]), .B(y[2329]), .Z(n27670) );
  AND U17481 ( .A(n8915), .B(n27670), .Z(n8916) );
  NAND U17482 ( .A(n12782), .B(n8916), .Z(n8918) );
  ANDN U17483 ( .B(x[2330]), .A(y[2330]), .Z(n8917) );
  ANDN U17484 ( .B(n8918), .A(n8917), .Z(n8919) );
  NANDN U17485 ( .A(n12780), .B(n8919), .Z(n8920) );
  NAND U17486 ( .A(n27676), .B(n8920), .Z(n8921) );
  NANDN U17487 ( .A(y[2333]), .B(x[2333]), .Z(n12779) );
  AND U17488 ( .A(n8921), .B(n12779), .Z(n8922) );
  NAND U17489 ( .A(n27675), .B(n8922), .Z(n8923) );
  ANDN U17490 ( .B(y[2333]), .A(x[2333]), .Z(n27677) );
  ANDN U17491 ( .B(n8923), .A(n27677), .Z(n8924) );
  NANDN U17492 ( .A(x[2334]), .B(y[2334]), .Z(n12777) );
  NAND U17493 ( .A(n8924), .B(n12777), .Z(n8925) );
  ANDN U17494 ( .B(x[2335]), .A(y[2335]), .Z(n12774) );
  ANDN U17495 ( .B(n8925), .A(n12774), .Z(n8926) );
  NANDN U17496 ( .A(n12778), .B(n8926), .Z(n8927) );
  NANDN U17497 ( .A(x[2335]), .B(y[2335]), .Z(n12776) );
  AND U17498 ( .A(n8927), .B(n12776), .Z(n8928) );
  NAND U17499 ( .A(n19398), .B(n8928), .Z(n8929) );
  NANDN U17500 ( .A(n27690), .B(n8929), .Z(n8930) );
  NAND U17501 ( .A(n27692), .B(n8930), .Z(n8931) );
  NAND U17502 ( .A(n27693), .B(n8931), .Z(n8932) );
  NANDN U17503 ( .A(x[2340]), .B(y[2340]), .Z(n12771) );
  AND U17504 ( .A(n8932), .B(n12771), .Z(n8933) );
  NANDN U17505 ( .A(n19402), .B(n8933), .Z(n8934) );
  NANDN U17506 ( .A(y[2340]), .B(x[2340]), .Z(n19408) );
  AND U17507 ( .A(n8934), .B(n19408), .Z(n8935) );
  NANDN U17508 ( .A(y[2341]), .B(x[2341]), .Z(n12769) );
  NAND U17509 ( .A(n8935), .B(n12769), .Z(n8936) );
  ANDN U17510 ( .B(y[2342]), .A(x[2342]), .Z(n12766) );
  ANDN U17511 ( .B(n8936), .A(n12766), .Z(n8937) );
  NANDN U17512 ( .A(n12770), .B(n8937), .Z(n8939) );
  NANDN U17513 ( .A(y[2343]), .B(x[2343]), .Z(n12765) );
  NANDN U17514 ( .A(y[2342]), .B(x[2342]), .Z(n12768) );
  AND U17515 ( .A(n12765), .B(n12768), .Z(n8938) );
  NAND U17516 ( .A(n8939), .B(n8938), .Z(n8940) );
  AND U17517 ( .A(n12767), .B(n8940), .Z(n8941) );
  NANDN U17518 ( .A(x[2344]), .B(y[2344]), .Z(n12763) );
  AND U17519 ( .A(n8941), .B(n12763), .Z(n8942) );
  NANDN U17520 ( .A(y[2344]), .B(x[2344]), .Z(n12764) );
  NANDN U17521 ( .A(n8942), .B(n12764), .Z(n8943) );
  NANDN U17522 ( .A(y[2345]), .B(x[2345]), .Z(n12761) );
  NANDN U17523 ( .A(n8943), .B(n12761), .Z(n8944) );
  AND U17524 ( .A(n12762), .B(n8944), .Z(n8945) );
  NANDN U17525 ( .A(x[2346]), .B(y[2346]), .Z(n12759) );
  AND U17526 ( .A(n8945), .B(n12759), .Z(n8947) );
  NANDN U17527 ( .A(y[2347]), .B(x[2347]), .Z(n12757) );
  ANDN U17528 ( .B(x[2346]), .A(y[2346]), .Z(n12760) );
  ANDN U17529 ( .B(n12757), .A(n12760), .Z(n8946) );
  NANDN U17530 ( .A(n8947), .B(n8946), .Z(n8948) );
  NANDN U17531 ( .A(n12758), .B(n8948), .Z(n8949) );
  ANDN U17532 ( .B(y[2348]), .A(x[2348]), .Z(n12754) );
  OR U17533 ( .A(n8949), .B(n12754), .Z(n8950) );
  NAND U17534 ( .A(n8951), .B(n8950), .Z(n8952) );
  NANDN U17535 ( .A(x[2349]), .B(y[2349]), .Z(n12755) );
  AND U17536 ( .A(n8952), .B(n12755), .Z(n8953) );
  NAND U17537 ( .A(n19421), .B(n8953), .Z(n8954) );
  NANDN U17538 ( .A(n12752), .B(n8954), .Z(n8955) );
  NANDN U17539 ( .A(y[2351]), .B(x[2351]), .Z(n12751) );
  NANDN U17540 ( .A(n8955), .B(n12751), .Z(n8956) );
  ANDN U17541 ( .B(y[2352]), .A(x[2352]), .Z(n27722) );
  ANDN U17542 ( .B(n8956), .A(n27722), .Z(n8957) );
  NANDN U17543 ( .A(x[2351]), .B(y[2351]), .Z(n19420) );
  NAND U17544 ( .A(n8957), .B(n19420), .Z(n8958) );
  ANDN U17545 ( .B(x[2352]), .A(y[2352]), .Z(n12750) );
  ANDN U17546 ( .B(n8958), .A(n12750), .Z(n8959) );
  NAND U17547 ( .A(n27723), .B(n8959), .Z(n8960) );
  AND U17548 ( .A(n27724), .B(n8960), .Z(n8962) );
  NANDN U17549 ( .A(y[2354]), .B(x[2354]), .Z(n27725) );
  ANDN U17550 ( .B(x[2355]), .A(y[2355]), .Z(n12748) );
  ANDN U17551 ( .B(n27725), .A(n12748), .Z(n8961) );
  NANDN U17552 ( .A(n8962), .B(n8961), .Z(n8963) );
  NAND U17553 ( .A(n12749), .B(n8963), .Z(n8964) );
  ANDN U17554 ( .B(y[2355]), .A(x[2355]), .Z(n27726) );
  OR U17555 ( .A(n8964), .B(n27726), .Z(n8965) );
  AND U17556 ( .A(n8966), .B(n8965), .Z(n8968) );
  NANDN U17557 ( .A(x[2357]), .B(y[2357]), .Z(n19433) );
  ANDN U17558 ( .B(y[2358]), .A(x[2358]), .Z(n27730) );
  ANDN U17559 ( .B(n19433), .A(n27730), .Z(n8967) );
  NANDN U17560 ( .A(n8968), .B(n8967), .Z(n8971) );
  NANDN U17561 ( .A(y[2359]), .B(x[2359]), .Z(n8970) );
  NANDN U17562 ( .A(y[2358]), .B(x[2358]), .Z(n8969) );
  AND U17563 ( .A(n8970), .B(n8969), .Z(n27731) );
  AND U17564 ( .A(n8971), .B(n27731), .Z(n8974) );
  NANDN U17565 ( .A(x[2359]), .B(y[2359]), .Z(n8973) );
  NANDN U17566 ( .A(x[2360]), .B(y[2360]), .Z(n8972) );
  NAND U17567 ( .A(n8973), .B(n8972), .Z(n19439) );
  OR U17568 ( .A(n8974), .B(n19439), .Z(n8977) );
  NANDN U17569 ( .A(y[2361]), .B(x[2361]), .Z(n8976) );
  NANDN U17570 ( .A(y[2360]), .B(x[2360]), .Z(n8975) );
  AND U17571 ( .A(n8976), .B(n8975), .Z(n12747) );
  AND U17572 ( .A(n8977), .B(n12747), .Z(n8979) );
  NANDN U17573 ( .A(x[2361]), .B(y[2361]), .Z(n27734) );
  NANDN U17574 ( .A(x[2362]), .B(y[2362]), .Z(n8978) );
  AND U17575 ( .A(n27734), .B(n8978), .Z(n19443) );
  NANDN U17576 ( .A(n8979), .B(n19443), .Z(n8980) );
  NAND U17577 ( .A(n8981), .B(n8980), .Z(n8982) );
  NANDN U17578 ( .A(n27736), .B(n8982), .Z(n8983) );
  NAND U17579 ( .A(n27737), .B(n8983), .Z(n8984) );
  ANDN U17580 ( .B(y[2366]), .A(x[2366]), .Z(n19456) );
  ANDN U17581 ( .B(n8984), .A(n19456), .Z(n8985) );
  NANDN U17582 ( .A(n27738), .B(n8985), .Z(n8986) );
  NANDN U17583 ( .A(y[2366]), .B(x[2366]), .Z(n27739) );
  AND U17584 ( .A(n8986), .B(n27739), .Z(n8987) );
  NANDN U17585 ( .A(n12744), .B(n8987), .Z(n8988) );
  NAND U17586 ( .A(n8989), .B(n8988), .Z(n8990) );
  NANDN U17587 ( .A(y[2368]), .B(x[2368]), .Z(n12745) );
  AND U17588 ( .A(n8990), .B(n12745), .Z(n8991) );
  NAND U17589 ( .A(n12741), .B(n8991), .Z(n8992) );
  NANDN U17590 ( .A(n24253), .B(n8992), .Z(n8993) );
  ANDN U17591 ( .B(y[2369]), .A(x[2369]), .Z(n12742) );
  OR U17592 ( .A(n8993), .B(n12742), .Z(n8994) );
  NAND U17593 ( .A(n8995), .B(n8994), .Z(n8996) );
  NANDN U17594 ( .A(n27745), .B(n8996), .Z(n8997) );
  NANDN U17595 ( .A(y[2372]), .B(x[2372]), .Z(n27746) );
  AND U17596 ( .A(n8997), .B(n27746), .Z(n8998) );
  NAND U17597 ( .A(n12739), .B(n8998), .Z(n8999) );
  NAND U17598 ( .A(n27749), .B(n8999), .Z(n9000) );
  ANDN U17599 ( .B(y[2373]), .A(x[2373]), .Z(n27747) );
  OR U17600 ( .A(n9000), .B(n27747), .Z(n9001) );
  AND U17601 ( .A(n9002), .B(n9001), .Z(n9003) );
  ANDN U17602 ( .B(y[2376]), .A(x[2376]), .Z(n19476) );
  NANDN U17603 ( .A(x[2375]), .B(y[2375]), .Z(n12737) );
  NANDN U17604 ( .A(n19476), .B(n12737), .Z(n27751) );
  OR U17605 ( .A(n9003), .B(n27751), .Z(n9004) );
  AND U17606 ( .A(n27752), .B(n9004), .Z(n9005) );
  NAND U17607 ( .A(n12736), .B(n9005), .Z(n9006) );
  NANDN U17608 ( .A(x[2377]), .B(y[2377]), .Z(n19477) );
  AND U17609 ( .A(n9006), .B(n19477), .Z(n9007) );
  NANDN U17610 ( .A(x[2378]), .B(y[2378]), .Z(n19481) );
  NAND U17611 ( .A(n9007), .B(n19481), .Z(n9008) );
  ANDN U17612 ( .B(x[2379]), .A(y[2379]), .Z(n27756) );
  ANDN U17613 ( .B(n9008), .A(n27756), .Z(n9009) );
  NANDN U17614 ( .A(n12735), .B(n9009), .Z(n9010) );
  AND U17615 ( .A(n19480), .B(n9010), .Z(n9011) );
  AND U17616 ( .A(n27757), .B(n9011), .Z(n9013) );
  NANDN U17617 ( .A(y[2381]), .B(x[2381]), .Z(n12734) );
  NANDN U17618 ( .A(y[2380]), .B(x[2380]), .Z(n19484) );
  NANDN U17619 ( .A(n9013), .B(n27758), .Z(n9014) );
  AND U17620 ( .A(n27759), .B(n9014), .Z(n9018) );
  NANDN U17621 ( .A(y[2384]), .B(x[2384]), .Z(n9016) );
  NANDN U17622 ( .A(y[2383]), .B(x[2383]), .Z(n9015) );
  NAND U17623 ( .A(n9016), .B(n9015), .Z(n19491) );
  NANDN U17624 ( .A(y[2382]), .B(x[2382]), .Z(n12733) );
  NANDN U17625 ( .A(n9018), .B(n27760), .Z(n9019) );
  NAND U17626 ( .A(n27761), .B(n9019), .Z(n9020) );
  AND U17627 ( .A(n27762), .B(n9020), .Z(n9021) );
  OR U17628 ( .A(n27763), .B(n9021), .Z(n9022) );
  NAND U17629 ( .A(n27765), .B(n9022), .Z(n9023) );
  NANDN U17630 ( .A(n27766), .B(n9023), .Z(n9024) );
  NANDN U17631 ( .A(y[2390]), .B(x[2390]), .Z(n24252) );
  AND U17632 ( .A(n9024), .B(n24252), .Z(n9025) );
  ANDN U17633 ( .B(y[2391]), .A(x[2391]), .Z(n24251) );
  OR U17634 ( .A(n9025), .B(n24251), .Z(n9028) );
  NANDN U17635 ( .A(y[2392]), .B(x[2392]), .Z(n9027) );
  NANDN U17636 ( .A(y[2391]), .B(x[2391]), .Z(n9026) );
  AND U17637 ( .A(n9027), .B(n9026), .Z(n24250) );
  AND U17638 ( .A(n9028), .B(n24250), .Z(n9029) );
  ANDN U17639 ( .B(y[2392]), .A(x[2392]), .Z(n12724) );
  OR U17640 ( .A(n9029), .B(n12724), .Z(n9030) );
  NANDN U17641 ( .A(n27768), .B(n9030), .Z(n9031) );
  AND U17642 ( .A(n27769), .B(n9031), .Z(n9032) );
  OR U17643 ( .A(n27770), .B(n9032), .Z(n9033) );
  NAND U17644 ( .A(n27771), .B(n9033), .Z(n9034) );
  NANDN U17645 ( .A(n19523), .B(n9034), .Z(n9037) );
  NANDN U17646 ( .A(x[2398]), .B(y[2398]), .Z(n9036) );
  NANDN U17647 ( .A(x[2397]), .B(y[2397]), .Z(n9035) );
  AND U17648 ( .A(n9036), .B(n9035), .Z(n24249) );
  AND U17649 ( .A(n9037), .B(n24249), .Z(n9042) );
  NANDN U17650 ( .A(y[2399]), .B(x[2399]), .Z(n9039) );
  NANDN U17651 ( .A(y[2398]), .B(x[2398]), .Z(n9038) );
  AND U17652 ( .A(n9039), .B(n9038), .Z(n9041) );
  NAND U17653 ( .A(n9041), .B(n9040), .Z(n27773) );
  OR U17654 ( .A(n9042), .B(n27773), .Z(n9043) );
  NAND U17655 ( .A(n12723), .B(n9043), .Z(n9044) );
  NANDN U17656 ( .A(n27775), .B(n9044), .Z(n9047) );
  NANDN U17657 ( .A(x[2402]), .B(y[2402]), .Z(n9045) );
  AND U17658 ( .A(n9046), .B(n9045), .Z(n27778) );
  AND U17659 ( .A(n9047), .B(n27778), .Z(n9048) );
  NAND U17660 ( .A(n12722), .B(n9048), .Z(n9049) );
  NANDN U17661 ( .A(n27780), .B(n9049), .Z(n9051) );
  NANDN U17662 ( .A(x[2406]), .B(y[2406]), .Z(n12717) );
  NANDN U17663 ( .A(x[2405]), .B(y[2405]), .Z(n27781) );
  AND U17664 ( .A(n12717), .B(n27781), .Z(n9050) );
  NAND U17665 ( .A(n9051), .B(n9050), .Z(n9052) );
  AND U17666 ( .A(n27782), .B(n9052), .Z(n9053) );
  ANDN U17667 ( .B(y[2407]), .A(x[2407]), .Z(n12719) );
  OR U17668 ( .A(n9053), .B(n12719), .Z(n9054) );
  AND U17669 ( .A(n27785), .B(n9054), .Z(n9055) );
  OR U17670 ( .A(n19541), .B(n9055), .Z(n9056) );
  NAND U17671 ( .A(n27789), .B(n9056), .Z(n9057) );
  NANDN U17672 ( .A(n27790), .B(n9057), .Z(n9058) );
  AND U17673 ( .A(n27791), .B(n9058), .Z(n9059) );
  OR U17674 ( .A(n27792), .B(n9059), .Z(n9060) );
  NAND U17675 ( .A(n27793), .B(n9060), .Z(n9061) );
  NANDN U17676 ( .A(n27794), .B(n9061), .Z(n9062) );
  AND U17677 ( .A(n27797), .B(n9062), .Z(n9063) );
  OR U17678 ( .A(n19549), .B(n9063), .Z(n9064) );
  AND U17679 ( .A(n9065), .B(n9064), .Z(n9069) );
  NANDN U17680 ( .A(x[2422]), .B(y[2422]), .Z(n9067) );
  ANDN U17681 ( .B(n9067), .A(n9066), .Z(n19558) );
  NANDN U17682 ( .A(x[2421]), .B(y[2421]), .Z(n9068) );
  NAND U17683 ( .A(n19558), .B(n9068), .Z(n27800) );
  OR U17684 ( .A(n9069), .B(n27800), .Z(n9070) );
  NAND U17685 ( .A(n9071), .B(n9070), .Z(n9072) );
  NANDN U17686 ( .A(n24245), .B(n9072), .Z(n9073) );
  NANDN U17687 ( .A(n27802), .B(n9073), .Z(n9074) );
  AND U17688 ( .A(n12711), .B(n9074), .Z(n9075) );
  NAND U17689 ( .A(n12714), .B(n9075), .Z(n9076) );
  ANDN U17690 ( .B(x[2429]), .A(y[2429]), .Z(n12708) );
  ANDN U17691 ( .B(n9076), .A(n12708), .Z(n9077) );
  NANDN U17692 ( .A(n12712), .B(n9077), .Z(n9078) );
  NANDN U17693 ( .A(x[2430]), .B(y[2430]), .Z(n12707) );
  AND U17694 ( .A(n9078), .B(n12707), .Z(n9079) );
  NANDN U17695 ( .A(n12710), .B(n9079), .Z(n9080) );
  NAND U17696 ( .A(n27809), .B(n9080), .Z(n9081) );
  NANDN U17697 ( .A(n27810), .B(n9081), .Z(n9082) );
  OR U17698 ( .A(n12704), .B(n9082), .Z(n9083) );
  AND U17699 ( .A(n27811), .B(n9083), .Z(n9089) );
  NANDN U17700 ( .A(x[2433]), .B(y[2433]), .Z(n12703) );
  OR U17701 ( .A(n9084), .B(n12703), .Z(n9087) );
  NANDN U17702 ( .A(x[2435]), .B(y[2435]), .Z(n9086) );
  NANDN U17703 ( .A(x[2434]), .B(y[2434]), .Z(n9085) );
  AND U17704 ( .A(n9086), .B(n9085), .Z(n12702) );
  AND U17705 ( .A(n9087), .B(n12702), .Z(n9088) );
  NANDN U17706 ( .A(n9089), .B(n9088), .Z(n9090) );
  NANDN U17707 ( .A(n12701), .B(n9090), .Z(n9091) );
  AND U17708 ( .A(n12699), .B(n9091), .Z(n9092) );
  ANDN U17709 ( .B(x[2437]), .A(y[2437]), .Z(n12697) );
  OR U17710 ( .A(n9092), .B(n12697), .Z(n9093) );
  AND U17711 ( .A(n12700), .B(n9093), .Z(n9094) );
  NANDN U17712 ( .A(x[2438]), .B(y[2438]), .Z(n12695) );
  AND U17713 ( .A(n9094), .B(n12695), .Z(n9096) );
  NANDN U17714 ( .A(y[2438]), .B(x[2438]), .Z(n12698) );
  ANDN U17715 ( .B(x[2439]), .A(y[2439]), .Z(n12693) );
  ANDN U17716 ( .B(n12698), .A(n12693), .Z(n9095) );
  NANDN U17717 ( .A(n9096), .B(n9095), .Z(n9097) );
  AND U17718 ( .A(n12696), .B(n9097), .Z(n9098) );
  OR U17719 ( .A(n9099), .B(n9098), .Z(n9100) );
  NAND U17720 ( .A(n27817), .B(n9100), .Z(n9101) );
  NANDN U17721 ( .A(n24242), .B(n9101), .Z(n9102) );
  NAND U17722 ( .A(n9103), .B(n9102), .Z(n9104) );
  NAND U17723 ( .A(n27819), .B(n9104), .Z(n9105) );
  AND U17724 ( .A(n19599), .B(n9105), .Z(n9109) );
  NANDN U17725 ( .A(x[2445]), .B(y[2445]), .Z(n19593) );
  NANDN U17726 ( .A(x[2446]), .B(y[2446]), .Z(n19597) );
  AND U17727 ( .A(n19593), .B(n19597), .Z(n9107) );
  NANDN U17728 ( .A(n9107), .B(n9106), .Z(n9108) );
  NAND U17729 ( .A(n9109), .B(n9108), .Z(n9110) );
  NANDN U17730 ( .A(n19601), .B(n9110), .Z(n9111) );
  AND U17731 ( .A(n12690), .B(n9111), .Z(n9112) );
  NAND U17732 ( .A(n19603), .B(n9112), .Z(n9113) );
  NANDN U17733 ( .A(n9114), .B(n9113), .Z(n9115) );
  AND U17734 ( .A(n27826), .B(n9115), .Z(n9116) );
  NANDN U17735 ( .A(y[2452]), .B(x[2452]), .Z(n19609) );
  NANDN U17736 ( .A(y[2453]), .B(x[2453]), .Z(n12689) );
  NAND U17737 ( .A(n19609), .B(n12689), .Z(n27827) );
  OR U17738 ( .A(n9116), .B(n27827), .Z(n9117) );
  NAND U17739 ( .A(n27828), .B(n9117), .Z(n9118) );
  NANDN U17740 ( .A(n27829), .B(n9118), .Z(n9119) );
  NAND U17741 ( .A(n27830), .B(n9119), .Z(n9120) );
  ANDN U17742 ( .B(x[2457]), .A(y[2457]), .Z(n12683) );
  ANDN U17743 ( .B(n9120), .A(n12683), .Z(n9121) );
  NANDN U17744 ( .A(n12686), .B(n9121), .Z(n9122) );
  NANDN U17745 ( .A(x[2458]), .B(y[2458]), .Z(n19629) );
  AND U17746 ( .A(n9122), .B(n19629), .Z(n9123) );
  NAND U17747 ( .A(n27832), .B(n9123), .Z(n9124) );
  NAND U17748 ( .A(n9125), .B(n9124), .Z(n9126) );
  AND U17749 ( .A(n24240), .B(n9126), .Z(n9128) );
  NANDN U17750 ( .A(y[2460]), .B(x[2460]), .Z(n24239) );
  ANDN U17751 ( .B(x[2461]), .A(y[2461]), .Z(n12680) );
  ANDN U17752 ( .B(n24239), .A(n12680), .Z(n9127) );
  NANDN U17753 ( .A(n9128), .B(n9127), .Z(n9129) );
  NANDN U17754 ( .A(n9130), .B(n9129), .Z(n9131) );
  NANDN U17755 ( .A(y[2463]), .B(x[2463]), .Z(n12678) );
  AND U17756 ( .A(n9131), .B(n12678), .Z(n9132) );
  NANDN U17757 ( .A(y[2462]), .B(x[2462]), .Z(n12681) );
  NAND U17758 ( .A(n9132), .B(n12681), .Z(n9133) );
  NANDN U17759 ( .A(n24238), .B(n9133), .Z(n9134) );
  AND U17760 ( .A(n27841), .B(n9134), .Z(n9136) );
  NANDN U17761 ( .A(x[2466]), .B(y[2466]), .Z(n12674) );
  ANDN U17762 ( .B(y[2465]), .A(x[2465]), .Z(n12677) );
  ANDN U17763 ( .B(n12674), .A(n12677), .Z(n9135) );
  NANDN U17764 ( .A(n9136), .B(n9135), .Z(n9137) );
  NANDN U17765 ( .A(y[2466]), .B(x[2466]), .Z(n12676) );
  AND U17766 ( .A(n9137), .B(n12676), .Z(n9138) );
  NANDN U17767 ( .A(x[2467]), .B(y[2467]), .Z(n12675) );
  NANDN U17768 ( .A(n9138), .B(n12675), .Z(n9141) );
  NANDN U17769 ( .A(y[2468]), .B(x[2468]), .Z(n9140) );
  NANDN U17770 ( .A(y[2467]), .B(x[2467]), .Z(n9139) );
  AND U17771 ( .A(n9140), .B(n9139), .Z(n19648) );
  AND U17772 ( .A(n9141), .B(n19648), .Z(n9144) );
  NANDN U17773 ( .A(x[2469]), .B(y[2469]), .Z(n9143) );
  NANDN U17774 ( .A(x[2468]), .B(y[2468]), .Z(n9142) );
  NAND U17775 ( .A(n9143), .B(n9142), .Z(n12673) );
  OR U17776 ( .A(n9144), .B(n12673), .Z(n9145) );
  NANDN U17777 ( .A(y[2469]), .B(x[2469]), .Z(n19653) );
  AND U17778 ( .A(n9145), .B(n19653), .Z(n9146) );
  NANDN U17779 ( .A(x[2470]), .B(y[2470]), .Z(n12672) );
  NANDN U17780 ( .A(n9146), .B(n12672), .Z(n9147) );
  AND U17781 ( .A(n27850), .B(n9147), .Z(n9149) );
  ANDN U17782 ( .B(y[2471]), .A(x[2471]), .Z(n27849) );
  IV U17783 ( .A(n27849), .Z(n12671) );
  ANDN U17784 ( .B(y[2472]), .A(x[2472]), .Z(n12668) );
  ANDN U17785 ( .B(n12671), .A(n12668), .Z(n9148) );
  NANDN U17786 ( .A(n9149), .B(n9148), .Z(n9150) );
  AND U17787 ( .A(n27851), .B(n9150), .Z(n9155) );
  NANDN U17788 ( .A(x[2474]), .B(y[2474]), .Z(n9152) );
  NANDN U17789 ( .A(x[2473]), .B(y[2473]), .Z(n9151) );
  AND U17790 ( .A(n9152), .B(n9151), .Z(n9154) );
  NANDN U17791 ( .A(x[2475]), .B(y[2475]), .Z(n9153) );
  AND U17792 ( .A(n9154), .B(n9153), .Z(n12669) );
  NANDN U17793 ( .A(n9155), .B(n12669), .Z(n9156) );
  NANDN U17794 ( .A(n27853), .B(n9156), .Z(n9157) );
  AND U17795 ( .A(n27854), .B(n9157), .Z(n9160) );
  NANDN U17796 ( .A(y[2477]), .B(x[2477]), .Z(n9159) );
  NANDN U17797 ( .A(y[2478]), .B(x[2478]), .Z(n9158) );
  NAND U17798 ( .A(n9159), .B(n9158), .Z(n27855) );
  OR U17799 ( .A(n9160), .B(n27855), .Z(n9161) );
  AND U17800 ( .A(n27856), .B(n9161), .Z(n9162) );
  OR U17801 ( .A(n27858), .B(n9162), .Z(n9163) );
  NAND U17802 ( .A(n27859), .B(n9163), .Z(n9164) );
  NANDN U17803 ( .A(n12666), .B(n9164), .Z(n9165) );
  NANDN U17804 ( .A(x[2481]), .B(y[2481]), .Z(n27861) );
  AND U17805 ( .A(n9165), .B(n27861), .Z(n9166) );
  NAND U17806 ( .A(n12665), .B(n9166), .Z(n9167) );
  NAND U17807 ( .A(n27862), .B(n9167), .Z(n9168) );
  ANDN U17808 ( .B(x[2483]), .A(y[2483]), .Z(n12662) );
  OR U17809 ( .A(n9168), .B(n12662), .Z(n9169) );
  AND U17810 ( .A(n27866), .B(n9169), .Z(n9170) );
  NANDN U17811 ( .A(x[2483]), .B(y[2483]), .Z(n12664) );
  NAND U17812 ( .A(n9170), .B(n12664), .Z(n9171) );
  NANDN U17813 ( .A(y[2484]), .B(x[2484]), .Z(n12663) );
  AND U17814 ( .A(n9171), .B(n12663), .Z(n9172) );
  NANDN U17815 ( .A(n27867), .B(n9172), .Z(n9173) );
  AND U17816 ( .A(n27868), .B(n9173), .Z(n9174) );
  NANDN U17817 ( .A(y[2487]), .B(x[2487]), .Z(n12659) );
  ANDN U17818 ( .B(x[2486]), .A(y[2486]), .Z(n19673) );
  ANDN U17819 ( .B(n12659), .A(n19673), .Z(n27869) );
  NANDN U17820 ( .A(n9174), .B(n27869), .Z(n9175) );
  NAND U17821 ( .A(n9176), .B(n9175), .Z(n9178) );
  NANDN U17822 ( .A(y[2488]), .B(x[2488]), .Z(n27871) );
  NANDN U17823 ( .A(y[2489]), .B(x[2489]), .Z(n19682) );
  AND U17824 ( .A(n27871), .B(n19682), .Z(n9177) );
  NAND U17825 ( .A(n9178), .B(n9177), .Z(n9179) );
  AND U17826 ( .A(n27874), .B(n9179), .Z(n9180) );
  NANDN U17827 ( .A(n12657), .B(n9180), .Z(n9181) );
  NAND U17828 ( .A(n27875), .B(n9181), .Z(n9182) );
  NANDN U17829 ( .A(n9183), .B(n9182), .Z(n9184) );
  NANDN U17830 ( .A(y[2492]), .B(x[2492]), .Z(n12655) );
  NANDN U17831 ( .A(y[2493]), .B(x[2493]), .Z(n12653) );
  AND U17832 ( .A(n12655), .B(n12653), .Z(n24237) );
  AND U17833 ( .A(n9184), .B(n24237), .Z(n9186) );
  ANDN U17834 ( .B(y[2493]), .A(x[2493]), .Z(n12654) );
  ANDN U17835 ( .B(y[2494]), .A(x[2494]), .Z(n12651) );
  NOR U17836 ( .A(n12654), .B(n12651), .Z(n9185) );
  NANDN U17837 ( .A(n9186), .B(n9185), .Z(n9187) );
  NANDN U17838 ( .A(n12652), .B(n9187), .Z(n9188) );
  NAND U17839 ( .A(n27881), .B(n9188), .Z(n9189) );
  NAND U17840 ( .A(n27883), .B(n9189), .Z(n9190) );
  NANDN U17841 ( .A(n27884), .B(n9190), .Z(n9191) );
  AND U17842 ( .A(n27885), .B(n9191), .Z(n9193) );
  ANDN U17843 ( .B(y[2501]), .A(x[2501]), .Z(n19704) );
  NANDN U17844 ( .A(x[2502]), .B(y[2502]), .Z(n9192) );
  NANDN U17845 ( .A(n19704), .B(n9192), .Z(n27886) );
  OR U17846 ( .A(n9193), .B(n27886), .Z(n9194) );
  AND U17847 ( .A(n27887), .B(n9194), .Z(n9197) );
  NANDN U17848 ( .A(x[2504]), .B(y[2504]), .Z(n9196) );
  NANDN U17849 ( .A(x[2503]), .B(y[2503]), .Z(n9195) );
  AND U17850 ( .A(n9196), .B(n9195), .Z(n27888) );
  NANDN U17851 ( .A(n9197), .B(n27888), .Z(n9198) );
  NAND U17852 ( .A(n9199), .B(n9198), .Z(n9200) );
  NANDN U17853 ( .A(n9201), .B(n9200), .Z(n9202) );
  NANDN U17854 ( .A(y[2507]), .B(x[2507]), .Z(n19722) );
  AND U17855 ( .A(n9202), .B(n19722), .Z(n9203) );
  NANDN U17856 ( .A(n12648), .B(n9203), .Z(n9204) );
  NAND U17857 ( .A(n27894), .B(n9204), .Z(n9205) );
  NANDN U17858 ( .A(n27895), .B(n9205), .Z(n9206) );
  ANDN U17859 ( .B(y[2509]), .A(x[2509]), .Z(n27896) );
  ANDN U17860 ( .B(n9206), .A(n27896), .Z(n9207) );
  NAND U17861 ( .A(n19730), .B(n9207), .Z(n9208) );
  NAND U17862 ( .A(n27900), .B(n9208), .Z(n9209) );
  NANDN U17863 ( .A(y[2510]), .B(x[2510]), .Z(n27898) );
  NANDN U17864 ( .A(n9209), .B(n27898), .Z(n9210) );
  AND U17865 ( .A(n9211), .B(n9210), .Z(n9212) );
  OR U17866 ( .A(n27902), .B(n9212), .Z(n9213) );
  NAND U17867 ( .A(n27903), .B(n9213), .Z(n9214) );
  NANDN U17868 ( .A(n27904), .B(n9214), .Z(n9216) );
  NANDN U17869 ( .A(x[2516]), .B(y[2516]), .Z(n12642) );
  ANDN U17870 ( .B(y[2515]), .A(x[2515]), .Z(n27905) );
  ANDN U17871 ( .B(n12642), .A(n27905), .Z(n9215) );
  NAND U17872 ( .A(n9216), .B(n9215), .Z(n9217) );
  AND U17873 ( .A(n27906), .B(n9217), .Z(n9220) );
  NANDN U17874 ( .A(x[2517]), .B(y[2517]), .Z(n9219) );
  NANDN U17875 ( .A(x[2518]), .B(y[2518]), .Z(n9218) );
  NAND U17876 ( .A(n9219), .B(n9218), .Z(n12643) );
  OR U17877 ( .A(n9220), .B(n12643), .Z(n9223) );
  NANDN U17878 ( .A(y[2519]), .B(x[2519]), .Z(n9222) );
  NANDN U17879 ( .A(y[2518]), .B(x[2518]), .Z(n9221) );
  AND U17880 ( .A(n9222), .B(n9221), .Z(n12640) );
  AND U17881 ( .A(n9223), .B(n12640), .Z(n9226) );
  NANDN U17882 ( .A(x[2519]), .B(y[2519]), .Z(n9225) );
  NANDN U17883 ( .A(x[2520]), .B(y[2520]), .Z(n9224) );
  NAND U17884 ( .A(n9225), .B(n9224), .Z(n12639) );
  OR U17885 ( .A(n9226), .B(n12639), .Z(n9227) );
  NANDN U17886 ( .A(y[2520]), .B(x[2520]), .Z(n19749) );
  NANDN U17887 ( .A(y[2521]), .B(x[2521]), .Z(n19752) );
  AND U17888 ( .A(n19749), .B(n19752), .Z(n27910) );
  AND U17889 ( .A(n9227), .B(n27910), .Z(n9228) );
  ANDN U17890 ( .B(y[2521]), .A(x[2521]), .Z(n19751) );
  ANDN U17891 ( .B(y[2522]), .A(x[2522]), .Z(n19756) );
  OR U17892 ( .A(n19751), .B(n19756), .Z(n24236) );
  OR U17893 ( .A(n9228), .B(n24236), .Z(n9229) );
  NAND U17894 ( .A(n9230), .B(n9229), .Z(n9231) );
  NANDN U17895 ( .A(n24234), .B(n9231), .Z(n9232) );
  XOR U17896 ( .A(x[2524]), .B(y[2524]), .Z(n12637) );
  OR U17897 ( .A(n9232), .B(n12637), .Z(n9233) );
  AND U17898 ( .A(n9234), .B(n9233), .Z(n9235) );
  ANDN U17899 ( .B(y[2526]), .A(x[2526]), .Z(n19763) );
  NANDN U17900 ( .A(x[2525]), .B(y[2525]), .Z(n12636) );
  NANDN U17901 ( .A(n19763), .B(n12636), .Z(n24231) );
  OR U17902 ( .A(n9235), .B(n24231), .Z(n9236) );
  NANDN U17903 ( .A(y[2527]), .B(x[2527]), .Z(n24230) );
  AND U17904 ( .A(n9236), .B(n24230), .Z(n9237) );
  NANDN U17905 ( .A(n12634), .B(n9237), .Z(n9238) );
  AND U17906 ( .A(n9239), .B(n9238), .Z(n9240) );
  OR U17907 ( .A(n27916), .B(n9240), .Z(n9241) );
  NAND U17908 ( .A(n27917), .B(n9241), .Z(n9242) );
  NANDN U17909 ( .A(n27918), .B(n9242), .Z(n9244) );
  NANDN U17910 ( .A(x[2532]), .B(y[2532]), .Z(n9243) );
  NANDN U17911 ( .A(x[2533]), .B(y[2533]), .Z(n9245) );
  AND U17912 ( .A(n9243), .B(n9245), .Z(n19777) );
  NANDN U17913 ( .A(x[2531]), .B(y[2531]), .Z(n12629) );
  AND U17914 ( .A(n19777), .B(n12629), .Z(n27919) );
  AND U17915 ( .A(n9244), .B(n27919), .Z(n9246) );
  NANDN U17916 ( .A(y[2532]), .B(x[2532]), .Z(n12627) );
  ANDN U17917 ( .B(x[2533]), .A(y[2533]), .Z(n19781) );
  NANDN U17918 ( .A(n9246), .B(n27920), .Z(n9247) );
  NAND U17919 ( .A(n24229), .B(n9247), .Z(n9248) );
  NANDN U17920 ( .A(n27922), .B(n9248), .Z(n9249) );
  AND U17921 ( .A(n27923), .B(n9249), .Z(n9250) );
  ANDN U17922 ( .B(x[2536]), .A(y[2536]), .Z(n19785) );
  ANDN U17923 ( .B(x[2537]), .A(y[2537]), .Z(n19793) );
  OR U17924 ( .A(n19785), .B(n19793), .Z(n27924) );
  OR U17925 ( .A(n9250), .B(n27924), .Z(n9251) );
  AND U17926 ( .A(n27925), .B(n9251), .Z(n9252) );
  NANDN U17927 ( .A(x[2538]), .B(y[2538]), .Z(n12624) );
  AND U17928 ( .A(n9252), .B(n12624), .Z(n9253) );
  OR U17929 ( .A(n27926), .B(n9253), .Z(n9254) );
  AND U17930 ( .A(n9255), .B(n9254), .Z(n9258) );
  NANDN U17931 ( .A(y[2541]), .B(x[2541]), .Z(n12622) );
  ANDN U17932 ( .B(x[2540]), .A(y[2540]), .Z(n19797) );
  NAND U17933 ( .A(n9256), .B(n19797), .Z(n9257) );
  AND U17934 ( .A(n12622), .B(n9257), .Z(n24227) );
  NANDN U17935 ( .A(n9258), .B(n24227), .Z(n9259) );
  AND U17936 ( .A(n27928), .B(n9259), .Z(n9260) );
  OR U17937 ( .A(n27929), .B(n9260), .Z(n9261) );
  NAND U17938 ( .A(n27930), .B(n9261), .Z(n9262) );
  NANDN U17939 ( .A(n27931), .B(n9262), .Z(n9263) );
  NANDN U17940 ( .A(n27932), .B(n9263), .Z(n9264) );
  NANDN U17941 ( .A(y[2546]), .B(x[2546]), .Z(n19808) );
  NANDN U17942 ( .A(y[2547]), .B(x[2547]), .Z(n19816) );
  AND U17943 ( .A(n19808), .B(n19816), .Z(n27933) );
  AND U17944 ( .A(n9264), .B(n27933), .Z(n9265) );
  ANDN U17945 ( .B(y[2547]), .A(x[2547]), .Z(n19812) );
  NANDN U17946 ( .A(x[2548]), .B(y[2548]), .Z(n12614) );
  NANDN U17947 ( .A(n19812), .B(n12614), .Z(n24226) );
  OR U17948 ( .A(n9265), .B(n24226), .Z(n9266) );
  NAND U17949 ( .A(n9267), .B(n9266), .Z(n9268) );
  NANDN U17950 ( .A(n12612), .B(n9268), .Z(n9269) );
  ANDN U17951 ( .B(y[2549]), .A(x[2549]), .Z(n12613) );
  OR U17952 ( .A(n9269), .B(n12613), .Z(n9270) );
  AND U17953 ( .A(n9271), .B(n9270), .Z(n9272) );
  NANDN U17954 ( .A(x[2551]), .B(y[2551]), .Z(n19824) );
  NANDN U17955 ( .A(x[2552]), .B(y[2552]), .Z(n12610) );
  NAND U17956 ( .A(n19824), .B(n12610), .Z(n27942) );
  OR U17957 ( .A(n9272), .B(n27942), .Z(n9273) );
  NANDN U17958 ( .A(y[2552]), .B(x[2552]), .Z(n27941) );
  AND U17959 ( .A(n9273), .B(n27941), .Z(n9274) );
  NANDN U17960 ( .A(y[2553]), .B(x[2553]), .Z(n12609) );
  AND U17961 ( .A(n9274), .B(n12609), .Z(n9275) );
  NANDN U17962 ( .A(x[2553]), .B(y[2553]), .Z(n27940) );
  NANDN U17963 ( .A(n9275), .B(n27940), .Z(n9276) );
  XOR U17964 ( .A(x[2554]), .B(y[2554]), .Z(n12608) );
  OR U17965 ( .A(n9276), .B(n12608), .Z(n9277) );
  NANDN U17966 ( .A(y[2555]), .B(x[2555]), .Z(n27945) );
  AND U17967 ( .A(n9277), .B(n27945), .Z(n9278) );
  NANDN U17968 ( .A(n9279), .B(n9278), .Z(n9280) );
  AND U17969 ( .A(n9281), .B(n9280), .Z(n9282) );
  OR U17970 ( .A(n27947), .B(n9282), .Z(n9283) );
  NAND U17971 ( .A(n27948), .B(n9283), .Z(n9284) );
  NANDN U17972 ( .A(n27949), .B(n9284), .Z(n9285) );
  NANDN U17973 ( .A(x[2560]), .B(y[2560]), .Z(n12602) );
  AND U17974 ( .A(n9285), .B(n12602), .Z(n9286) );
  NAND U17975 ( .A(n27950), .B(n9286), .Z(n9287) );
  NANDN U17976 ( .A(n9288), .B(n9287), .Z(n9289) );
  AND U17977 ( .A(n12601), .B(n9289), .Z(n9290) );
  NANDN U17978 ( .A(x[2562]), .B(y[2562]), .Z(n12600) );
  NAND U17979 ( .A(n9290), .B(n12600), .Z(n9291) );
  ANDN U17980 ( .B(x[2563]), .A(y[2563]), .Z(n12598) );
  ANDN U17981 ( .B(n9291), .A(n12598), .Z(n9292) );
  NANDN U17982 ( .A(n27957), .B(n9292), .Z(n9294) );
  NANDN U17983 ( .A(x[2564]), .B(y[2564]), .Z(n12597) );
  NANDN U17984 ( .A(x[2563]), .B(y[2563]), .Z(n27956) );
  AND U17985 ( .A(n12597), .B(n27956), .Z(n9293) );
  NAND U17986 ( .A(n9294), .B(n9293), .Z(n9295) );
  AND U17987 ( .A(n12599), .B(n9295), .Z(n9296) );
  NANDN U17988 ( .A(y[2565]), .B(x[2565]), .Z(n12595) );
  NAND U17989 ( .A(n9296), .B(n12595), .Z(n9297) );
  ANDN U17990 ( .B(y[2566]), .A(x[2566]), .Z(n12593) );
  ANDN U17991 ( .B(n9297), .A(n12593), .Z(n9298) );
  NANDN U17992 ( .A(n12596), .B(n9298), .Z(n9299) );
  AND U17993 ( .A(n12594), .B(n9299), .Z(n9300) );
  NANDN U17994 ( .A(y[2567]), .B(x[2567]), .Z(n19854) );
  NAND U17995 ( .A(n9300), .B(n19854), .Z(n9301) );
  ANDN U17996 ( .B(y[2568]), .A(x[2568]), .Z(n19856) );
  ANDN U17997 ( .B(n9301), .A(n19856), .Z(n9302) );
  NANDN U17998 ( .A(n12592), .B(n9302), .Z(n9304) );
  NANDN U17999 ( .A(y[2569]), .B(x[2569]), .Z(n12591) );
  NANDN U18000 ( .A(y[2568]), .B(x[2568]), .Z(n19853) );
  AND U18001 ( .A(n12591), .B(n19853), .Z(n9303) );
  NAND U18002 ( .A(n9304), .B(n9303), .Z(n9305) );
  AND U18003 ( .A(n24223), .B(n9305), .Z(n9306) );
  NANDN U18004 ( .A(x[2570]), .B(y[2570]), .Z(n12590) );
  NAND U18005 ( .A(n9306), .B(n12590), .Z(n9307) );
  ANDN U18006 ( .B(x[2571]), .A(y[2571]), .Z(n19861) );
  ANDN U18007 ( .B(n9307), .A(n19861), .Z(n9308) );
  NANDN U18008 ( .A(n24222), .B(n9308), .Z(n9309) );
  ANDN U18009 ( .B(y[2572]), .A(x[2572]), .Z(n27966) );
  ANDN U18010 ( .B(n9309), .A(n27966), .Z(n9310) );
  NANDN U18011 ( .A(n12589), .B(n9310), .Z(n9311) );
  NAND U18012 ( .A(n9312), .B(n9311), .Z(n9313) );
  NANDN U18013 ( .A(x[2573]), .B(y[2573]), .Z(n24221) );
  AND U18014 ( .A(n9313), .B(n24221), .Z(n9314) );
  NAND U18015 ( .A(n12587), .B(n9314), .Z(n9315) );
  NANDN U18016 ( .A(n12588), .B(n9315), .Z(n9316) );
  ANDN U18017 ( .B(x[2575]), .A(y[2575]), .Z(n12584) );
  OR U18018 ( .A(n9316), .B(n12584), .Z(n9317) );
  AND U18019 ( .A(n12586), .B(n9317), .Z(n9318) );
  NAND U18020 ( .A(n12585), .B(n9318), .Z(n9320) );
  ANDN U18021 ( .B(x[2576]), .A(y[2576]), .Z(n9319) );
  ANDN U18022 ( .B(n9320), .A(n9319), .Z(n9321) );
  NANDN U18023 ( .A(n12580), .B(n9321), .Z(n9322) );
  AND U18024 ( .A(n12582), .B(n9322), .Z(n9323) );
  NAND U18025 ( .A(n12577), .B(n9323), .Z(n9324) );
  NAND U18026 ( .A(n12581), .B(n9324), .Z(n9327) );
  NANDN U18027 ( .A(x[2580]), .B(y[2580]), .Z(n9326) );
  NANDN U18028 ( .A(x[2579]), .B(y[2579]), .Z(n9325) );
  NAND U18029 ( .A(n9326), .B(n9325), .Z(n12579) );
  ANDN U18030 ( .B(n9327), .A(n12579), .Z(n9330) );
  NANDN U18031 ( .A(y[2581]), .B(x[2581]), .Z(n9329) );
  NANDN U18032 ( .A(y[2580]), .B(x[2580]), .Z(n9328) );
  NAND U18033 ( .A(n9329), .B(n9328), .Z(n19874) );
  OR U18034 ( .A(n9330), .B(n19874), .Z(n9331) );
  NANDN U18035 ( .A(x[2581]), .B(y[2581]), .Z(n19873) );
  AND U18036 ( .A(n9331), .B(n19873), .Z(n9332) );
  NANDN U18037 ( .A(n19877), .B(n9332), .Z(n9333) );
  AND U18038 ( .A(n9334), .B(n9333), .Z(n9335) );
  OR U18039 ( .A(n27977), .B(n9335), .Z(n9336) );
  NAND U18040 ( .A(n27978), .B(n9336), .Z(n9337) );
  NANDN U18041 ( .A(n27979), .B(n9337), .Z(n9338) );
  NANDN U18042 ( .A(n24219), .B(n9338), .Z(n9339) );
  NANDN U18043 ( .A(x[2587]), .B(y[2587]), .Z(n12575) );
  NANDN U18044 ( .A(x[2588]), .B(y[2588]), .Z(n12574) );
  AND U18045 ( .A(n12575), .B(n12574), .Z(n24218) );
  AND U18046 ( .A(n9339), .B(n24218), .Z(n9340) );
  OR U18047 ( .A(n27981), .B(n9340), .Z(n9341) );
  NAND U18048 ( .A(n27982), .B(n9341), .Z(n9342) );
  NANDN U18049 ( .A(n27983), .B(n9342), .Z(n9343) );
  NAND U18050 ( .A(n27984), .B(n9343), .Z(n9344) );
  AND U18051 ( .A(n9345), .B(n9344), .Z(n9347) );
  ANDN U18052 ( .B(y[2593]), .A(x[2593]), .Z(n19910) );
  IV U18053 ( .A(n19910), .Z(n27985) );
  ANDN U18054 ( .B(y[2594]), .A(x[2594]), .Z(n12565) );
  ANDN U18055 ( .B(n27985), .A(n12565), .Z(n9346) );
  NANDN U18056 ( .A(n9347), .B(n9346), .Z(n9348) );
  NANDN U18057 ( .A(y[2595]), .B(x[2595]), .Z(n27988) );
  AND U18058 ( .A(n9348), .B(n27988), .Z(n9349) );
  NANDN U18059 ( .A(y[2594]), .B(x[2594]), .Z(n12567) );
  NAND U18060 ( .A(n9349), .B(n12567), .Z(n9350) );
  NANDN U18061 ( .A(n27989), .B(n9350), .Z(n9351) );
  NANDN U18062 ( .A(y[2596]), .B(x[2596]), .Z(n19915) );
  NANDN U18063 ( .A(y[2597]), .B(x[2597]), .Z(n12564) );
  AND U18064 ( .A(n19915), .B(n12564), .Z(n27990) );
  AND U18065 ( .A(n9351), .B(n27990), .Z(n9353) );
  ANDN U18066 ( .B(y[2597]), .A(x[2597]), .Z(n19920) );
  IV U18067 ( .A(n19920), .Z(n27991) );
  ANDN U18068 ( .B(y[2598]), .A(x[2598]), .Z(n12561) );
  ANDN U18069 ( .B(n27991), .A(n12561), .Z(n9352) );
  NANDN U18070 ( .A(n9353), .B(n9352), .Z(n9354) );
  NANDN U18071 ( .A(n27992), .B(n9354), .Z(n9355) );
  AND U18072 ( .A(n24216), .B(n9355), .Z(n9356) );
  NAND U18073 ( .A(n12562), .B(n9356), .Z(n9357) );
  NANDN U18074 ( .A(n27994), .B(n9357), .Z(n9358) );
  ANDN U18075 ( .B(y[2603]), .A(x[2603]), .Z(n27995) );
  ANDN U18076 ( .B(n9358), .A(n27995), .Z(n9359) );
  NANDN U18077 ( .A(x[2604]), .B(y[2604]), .Z(n19944) );
  NAND U18078 ( .A(n9359), .B(n19944), .Z(n9360) );
  ANDN U18079 ( .B(x[2605]), .A(y[2605]), .Z(n24211) );
  ANDN U18080 ( .B(n9360), .A(n24211), .Z(n9361) );
  NANDN U18081 ( .A(n19941), .B(n9361), .Z(n9363) );
  NANDN U18082 ( .A(x[2605]), .B(y[2605]), .Z(n19943) );
  NANDN U18083 ( .A(x[2606]), .B(y[2606]), .Z(n24210) );
  AND U18084 ( .A(n19943), .B(n24210), .Z(n9362) );
  NAND U18085 ( .A(n9363), .B(n9362), .Z(n9364) );
  AND U18086 ( .A(n27997), .B(n9364), .Z(n9365) );
  OR U18087 ( .A(n27998), .B(n9365), .Z(n9366) );
  NAND U18088 ( .A(n27999), .B(n9366), .Z(n9367) );
  NANDN U18089 ( .A(n28000), .B(n9367), .Z(n9368) );
  NANDN U18090 ( .A(y[2611]), .B(x[2611]), .Z(n12556) );
  AND U18091 ( .A(n9368), .B(n12556), .Z(n9369) );
  NAND U18092 ( .A(n28001), .B(n9369), .Z(n9370) );
  NAND U18093 ( .A(n28002), .B(n9370), .Z(n9371) );
  AND U18094 ( .A(n12555), .B(n9371), .Z(n9372) );
  NANDN U18095 ( .A(y[2613]), .B(x[2613]), .Z(n12554) );
  NAND U18096 ( .A(n9372), .B(n12554), .Z(n9373) );
  NANDN U18097 ( .A(n28006), .B(n9373), .Z(n9374) );
  AND U18098 ( .A(n12551), .B(n9374), .Z(n9375) );
  NAND U18099 ( .A(n28005), .B(n9375), .Z(n9376) );
  ANDN U18100 ( .B(y[2615]), .A(x[2615]), .Z(n12552) );
  ANDN U18101 ( .B(n9376), .A(n12552), .Z(n9377) );
  NANDN U18102 ( .A(n12550), .B(n9377), .Z(n9378) );
  NANDN U18103 ( .A(y[2617]), .B(x[2617]), .Z(n12548) );
  AND U18104 ( .A(n9378), .B(n12548), .Z(n9379) );
  NANDN U18105 ( .A(n9380), .B(n9379), .Z(n9381) );
  NAND U18106 ( .A(n28011), .B(n9381), .Z(n9382) );
  NANDN U18107 ( .A(n28012), .B(n9382), .Z(n9383) );
  NANDN U18108 ( .A(x[2619]), .B(y[2619]), .Z(n28013) );
  AND U18109 ( .A(n9383), .B(n28013), .Z(n9384) );
  NAND U18110 ( .A(n12547), .B(n9384), .Z(n9385) );
  NAND U18111 ( .A(n28016), .B(n9385), .Z(n9386) );
  OR U18112 ( .A(n28014), .B(n9386), .Z(n9387) );
  AND U18113 ( .A(n12546), .B(n9387), .Z(n9388) );
  NANDN U18114 ( .A(n28017), .B(n9388), .Z(n9389) );
  AND U18115 ( .A(n28018), .B(n9389), .Z(n9390) );
  ANDN U18116 ( .B(y[2623]), .A(x[2623]), .Z(n19989) );
  NANDN U18117 ( .A(x[2624]), .B(y[2624]), .Z(n19995) );
  NANDN U18118 ( .A(n19989), .B(n19995), .Z(n28019) );
  OR U18119 ( .A(n9390), .B(n28019), .Z(n9391) );
  AND U18120 ( .A(n28020), .B(n9391), .Z(n9392) );
  NANDN U18121 ( .A(x[2631]), .B(y[2631]), .Z(n9393) );
  NANDN U18122 ( .A(x[2632]), .B(y[2632]), .Z(n12545) );
  NAND U18123 ( .A(n9393), .B(n12545), .Z(n28032) );
  NANDN U18124 ( .A(y[2632]), .B(x[2632]), .Z(n24206) );
  NANDN U18125 ( .A(y[2633]), .B(x[2633]), .Z(n12543) );
  ANDN U18126 ( .B(y[2634]), .A(x[2634]), .Z(n28035) );
  NANDN U18127 ( .A(y[2635]), .B(x[2635]), .Z(n12541) );
  ANDN U18128 ( .B(x[2637]), .A(y[2637]), .Z(n28039) );
  ANDN U18129 ( .B(x[2636]), .A(y[2636]), .Z(n24203) );
  NANDN U18130 ( .A(x[2639]), .B(y[2639]), .Z(n12540) );
  NANDN U18131 ( .A(x[2640]), .B(y[2640]), .Z(n20031) );
  AND U18132 ( .A(n12540), .B(n20031), .Z(n24202) );
  NAND U18133 ( .A(n9395), .B(n9394), .Z(n9396) );
  NANDN U18134 ( .A(x[2641]), .B(y[2641]), .Z(n28043) );
  AND U18135 ( .A(n9396), .B(n28043), .Z(n9397) );
  NANDN U18136 ( .A(n12538), .B(n9397), .Z(n9398) );
  NAND U18137 ( .A(n9399), .B(n9398), .Z(n9400) );
  AND U18138 ( .A(n12539), .B(n9400), .Z(n9401) );
  NANDN U18139 ( .A(n12534), .B(n9401), .Z(n9402) );
  NAND U18140 ( .A(n12537), .B(n9402), .Z(n9403) );
  NANDN U18141 ( .A(n12535), .B(n9403), .Z(n9406) );
  NANDN U18142 ( .A(y[2646]), .B(x[2646]), .Z(n9405) );
  NANDN U18143 ( .A(y[2647]), .B(x[2647]), .Z(n9404) );
  AND U18144 ( .A(n9405), .B(n9404), .Z(n12532) );
  AND U18145 ( .A(n9406), .B(n12532), .Z(n9407) );
  NANDN U18146 ( .A(x[2647]), .B(y[2647]), .Z(n28048) );
  NANDN U18147 ( .A(n9407), .B(n28048), .Z(n9408) );
  ANDN U18148 ( .B(y[2648]), .A(x[2648]), .Z(n12529) );
  OR U18149 ( .A(n9408), .B(n12529), .Z(n9410) );
  NANDN U18150 ( .A(y[2648]), .B(x[2648]), .Z(n9409) );
  ANDN U18151 ( .B(x[2649]), .A(y[2649]), .Z(n12530) );
  ANDN U18152 ( .B(n9409), .A(n12530), .Z(n28049) );
  AND U18153 ( .A(n9410), .B(n28049), .Z(n9413) );
  NANDN U18154 ( .A(x[2649]), .B(y[2649]), .Z(n9412) );
  NANDN U18155 ( .A(x[2650]), .B(y[2650]), .Z(n9411) );
  NAND U18156 ( .A(n9412), .B(n9411), .Z(n12531) );
  OR U18157 ( .A(n9413), .B(n12531), .Z(n9416) );
  NANDN U18158 ( .A(y[2650]), .B(x[2650]), .Z(n9415) );
  NANDN U18159 ( .A(y[2651]), .B(x[2651]), .Z(n9414) );
  NAND U18160 ( .A(n9415), .B(n9414), .Z(n28051) );
  ANDN U18161 ( .B(n9416), .A(n28051), .Z(n9418) );
  NANDN U18162 ( .A(x[2651]), .B(y[2651]), .Z(n28052) );
  ANDN U18163 ( .B(y[2652]), .A(x[2652]), .Z(n12527) );
  ANDN U18164 ( .B(n28052), .A(n12527), .Z(n9417) );
  NANDN U18165 ( .A(n9418), .B(n9417), .Z(n9419) );
  NANDN U18166 ( .A(n28053), .B(n9419), .Z(n9420) );
  ANDN U18167 ( .B(x[2653]), .A(y[2653]), .Z(n12525) );
  OR U18168 ( .A(n9420), .B(n12525), .Z(n9421) );
  AND U18169 ( .A(n12528), .B(n9421), .Z(n9422) );
  NANDN U18170 ( .A(x[2654]), .B(y[2654]), .Z(n12524) );
  AND U18171 ( .A(n9422), .B(n12524), .Z(n9423) );
  NANDN U18172 ( .A(y[2654]), .B(x[2654]), .Z(n12526) );
  NANDN U18173 ( .A(n9423), .B(n12526), .Z(n9424) );
  NANDN U18174 ( .A(y[2655]), .B(x[2655]), .Z(n12522) );
  NANDN U18175 ( .A(n9424), .B(n12522), .Z(n9425) );
  NANDN U18176 ( .A(x[2656]), .B(y[2656]), .Z(n28059) );
  AND U18177 ( .A(n9425), .B(n28059), .Z(n9426) );
  NANDN U18178 ( .A(x[2655]), .B(y[2655]), .Z(n12523) );
  NAND U18179 ( .A(n9426), .B(n12523), .Z(n9427) );
  ANDN U18180 ( .B(x[2656]), .A(y[2656]), .Z(n12521) );
  ANDN U18181 ( .B(n9427), .A(n12521), .Z(n9428) );
  NANDN U18182 ( .A(n20052), .B(n9428), .Z(n9429) );
  AND U18183 ( .A(n28061), .B(n9429), .Z(n9431) );
  NANDN U18184 ( .A(y[2658]), .B(x[2658]), .Z(n28062) );
  ANDN U18185 ( .B(x[2659]), .A(y[2659]), .Z(n12518) );
  ANDN U18186 ( .B(n28062), .A(n12518), .Z(n9430) );
  NANDN U18187 ( .A(n9431), .B(n9430), .Z(n9432) );
  NAND U18188 ( .A(n12519), .B(n9432), .Z(n9433) );
  ANDN U18189 ( .B(y[2659]), .A(x[2659]), .Z(n28063) );
  OR U18190 ( .A(n9433), .B(n28063), .Z(n9434) );
  AND U18191 ( .A(n9435), .B(n9434), .Z(n9436) );
  ANDN U18192 ( .B(y[2662]), .A(x[2662]), .Z(n20065) );
  NANDN U18193 ( .A(x[2661]), .B(y[2661]), .Z(n12517) );
  NANDN U18194 ( .A(n20065), .B(n12517), .Z(n28066) );
  OR U18195 ( .A(n9436), .B(n28066), .Z(n9437) );
  AND U18196 ( .A(n28067), .B(n9437), .Z(n9438) );
  NANDN U18197 ( .A(y[2663]), .B(x[2663]), .Z(n12515) );
  AND U18198 ( .A(n9438), .B(n12515), .Z(n9439) );
  NANDN U18199 ( .A(x[2663]), .B(y[2663]), .Z(n12516) );
  NANDN U18200 ( .A(n9439), .B(n12516), .Z(n9440) );
  XOR U18201 ( .A(x[2664]), .B(y[2664]), .Z(n12514) );
  OR U18202 ( .A(n9440), .B(n12514), .Z(n9441) );
  AND U18203 ( .A(n28071), .B(n9441), .Z(n9442) );
  NANDN U18204 ( .A(n9443), .B(n9442), .Z(n9444) );
  AND U18205 ( .A(n9445), .B(n9444), .Z(n9446) );
  NANDN U18206 ( .A(y[2666]), .B(x[2666]), .Z(n12511) );
  NANDN U18207 ( .A(y[2667]), .B(x[2667]), .Z(n12509) );
  NAND U18208 ( .A(n12511), .B(n12509), .Z(n28074) );
  OR U18209 ( .A(n9446), .B(n28074), .Z(n9447) );
  NAND U18210 ( .A(n28075), .B(n9447), .Z(n9448) );
  NANDN U18211 ( .A(n28076), .B(n9448), .Z(n9450) );
  NANDN U18212 ( .A(x[2669]), .B(y[2669]), .Z(n28077) );
  NANDN U18213 ( .A(x[2670]), .B(y[2670]), .Z(n12507) );
  AND U18214 ( .A(n28077), .B(n12507), .Z(n9449) );
  NAND U18215 ( .A(n9450), .B(n9449), .Z(n9451) );
  AND U18216 ( .A(n28078), .B(n9451), .Z(n9452) );
  OR U18217 ( .A(n28080), .B(n9452), .Z(n9453) );
  NAND U18218 ( .A(n28081), .B(n9453), .Z(n9454) );
  NANDN U18219 ( .A(n28082), .B(n9454), .Z(n9455) );
  NANDN U18220 ( .A(n24199), .B(n9455), .Z(n9456) );
  AND U18221 ( .A(n28083), .B(n9456), .Z(n9457) );
  OR U18222 ( .A(n28084), .B(n9457), .Z(n9458) );
  NAND U18223 ( .A(n28085), .B(n9458), .Z(n9459) );
  NANDN U18224 ( .A(n28086), .B(n9459), .Z(n9460) );
  NAND U18225 ( .A(n28087), .B(n9460), .Z(n9461) );
  ANDN U18226 ( .B(x[2681]), .A(y[2681]), .Z(n12501) );
  ANDN U18227 ( .B(n9461), .A(n12501), .Z(n9462) );
  NAND U18228 ( .A(n28088), .B(n9462), .Z(n9463) );
  ANDN U18229 ( .B(y[2681]), .A(x[2681]), .Z(n28090) );
  ANDN U18230 ( .B(n9463), .A(n28090), .Z(n9464) );
  NAND U18231 ( .A(n12502), .B(n9464), .Z(n9465) );
  NAND U18232 ( .A(n9466), .B(n9465), .Z(n9467) );
  AND U18233 ( .A(n20118), .B(n9467), .Z(n9468) );
  NANDN U18234 ( .A(n12497), .B(n9468), .Z(n9469) );
  NAND U18235 ( .A(n9470), .B(n9469), .Z(n9471) );
  NANDN U18236 ( .A(x[2685]), .B(y[2685]), .Z(n12498) );
  AND U18237 ( .A(n9471), .B(n12498), .Z(n9472) );
  NAND U18238 ( .A(n12494), .B(n9472), .Z(n9473) );
  NAND U18239 ( .A(n28095), .B(n9473), .Z(n9474) );
  OR U18240 ( .A(n9475), .B(n9474), .Z(n9476) );
  AND U18241 ( .A(n12493), .B(n9476), .Z(n9477) );
  AND U18242 ( .A(n28096), .B(n9477), .Z(n9478) );
  OR U18243 ( .A(n28097), .B(n9478), .Z(n9479) );
  NANDN U18244 ( .A(n28098), .B(n9479), .Z(n9480) );
  NANDN U18245 ( .A(n28099), .B(n9480), .Z(n9481) );
  ANDN U18246 ( .B(y[2691]), .A(x[2691]), .Z(n28100) );
  ANDN U18247 ( .B(n9481), .A(n28100), .Z(n9482) );
  NAND U18248 ( .A(n12489), .B(n9482), .Z(n9483) );
  NAND U18249 ( .A(n28103), .B(n9483), .Z(n9484) );
  OR U18250 ( .A(n28101), .B(n9484), .Z(n9485) );
  AND U18251 ( .A(n12488), .B(n9485), .Z(n9486) );
  NANDN U18252 ( .A(n12485), .B(n9486), .Z(n9487) );
  NANDN U18253 ( .A(y[2694]), .B(x[2694]), .Z(n12487) );
  NANDN U18254 ( .A(y[2695]), .B(x[2695]), .Z(n12483) );
  AND U18255 ( .A(n12487), .B(n12483), .Z(n28106) );
  AND U18256 ( .A(n9487), .B(n28106), .Z(n9488) );
  NANDN U18257 ( .A(x[2695]), .B(y[2695]), .Z(n12486) );
  NANDN U18258 ( .A(x[2696]), .B(y[2696]), .Z(n20142) );
  NAND U18259 ( .A(n12486), .B(n20142), .Z(n28107) );
  OR U18260 ( .A(n9488), .B(n28107), .Z(n9489) );
  NAND U18261 ( .A(n28108), .B(n9489), .Z(n9490) );
  NANDN U18262 ( .A(n24196), .B(n9490), .Z(n9491) );
  NANDN U18263 ( .A(y[2698]), .B(x[2698]), .Z(n12482) );
  AND U18264 ( .A(n9491), .B(n12482), .Z(n9492) );
  NAND U18265 ( .A(n12479), .B(n9492), .Z(n9493) );
  NANDN U18266 ( .A(n12480), .B(n9493), .Z(n9494) );
  XOR U18267 ( .A(x[2700]), .B(y[2700]), .Z(n12478) );
  OR U18268 ( .A(n9494), .B(n12478), .Z(n9495) );
  AND U18269 ( .A(n9496), .B(n9495), .Z(n9497) );
  NANDN U18270 ( .A(x[2701]), .B(y[2701]), .Z(n20152) );
  NANDN U18271 ( .A(x[2702]), .B(y[2702]), .Z(n12476) );
  NAND U18272 ( .A(n20152), .B(n12476), .Z(n24194) );
  OR U18273 ( .A(n9497), .B(n24194), .Z(n9498) );
  NANDN U18274 ( .A(y[2702]), .B(x[2702]), .Z(n24193) );
  AND U18275 ( .A(n9498), .B(n24193), .Z(n9499) );
  NANDN U18276 ( .A(y[2703]), .B(x[2703]), .Z(n12474) );
  NAND U18277 ( .A(n9499), .B(n12474), .Z(n9500) );
  ANDN U18278 ( .B(y[2703]), .A(x[2703]), .Z(n12475) );
  ANDN U18279 ( .B(n9500), .A(n12475), .Z(n9501) );
  NANDN U18280 ( .A(n12473), .B(n9501), .Z(n9502) );
  AND U18281 ( .A(n9503), .B(n9502), .Z(n9504) );
  NANDN U18282 ( .A(y[2705]), .B(x[2705]), .Z(n12472) );
  NAND U18283 ( .A(n9504), .B(n12472), .Z(n9505) );
  NANDN U18284 ( .A(n24189), .B(n9505), .Z(n9506) );
  NANDN U18285 ( .A(y[2706]), .B(x[2706]), .Z(n24188) );
  AND U18286 ( .A(n9506), .B(n24188), .Z(n9507) );
  NANDN U18287 ( .A(y[2707]), .B(x[2707]), .Z(n12471) );
  NAND U18288 ( .A(n9507), .B(n12471), .Z(n9508) );
  ANDN U18289 ( .B(y[2707]), .A(x[2707]), .Z(n24191) );
  ANDN U18290 ( .B(n9508), .A(n24191), .Z(n9509) );
  NANDN U18291 ( .A(n12470), .B(n9509), .Z(n9510) );
  AND U18292 ( .A(n9511), .B(n9510), .Z(n9512) );
  NANDN U18293 ( .A(y[2709]), .B(x[2709]), .Z(n12468) );
  NAND U18294 ( .A(n9512), .B(n12468), .Z(n9513) );
  ANDN U18295 ( .B(y[2710]), .A(x[2710]), .Z(n12464) );
  ANDN U18296 ( .B(n9513), .A(n12464), .Z(n9514) );
  NANDN U18297 ( .A(n20167), .B(n9514), .Z(n9515) );
  AND U18298 ( .A(n12469), .B(n9515), .Z(n9516) );
  OR U18299 ( .A(n12467), .B(n9516), .Z(n9517) );
  NANDN U18300 ( .A(n20172), .B(n9517), .Z(n9518) );
  NANDN U18301 ( .A(n20171), .B(n9518), .Z(n9519) );
  ANDN U18302 ( .B(y[2714]), .A(x[2714]), .Z(n12461) );
  OR U18303 ( .A(n9519), .B(n12461), .Z(n9520) );
  AND U18304 ( .A(n9521), .B(n9520), .Z(n9522) );
  OR U18305 ( .A(n9523), .B(n9522), .Z(n9524) );
  NANDN U18306 ( .A(n28125), .B(n9524), .Z(n9525) );
  NANDN U18307 ( .A(n28126), .B(n9525), .Z(n9526) );
  NANDN U18308 ( .A(y[2718]), .B(x[2718]), .Z(n20181) );
  NANDN U18309 ( .A(y[2719]), .B(x[2719]), .Z(n12459) );
  AND U18310 ( .A(n20181), .B(n12459), .Z(n24185) );
  AND U18311 ( .A(n9526), .B(n24185), .Z(n9527) );
  ANDN U18312 ( .B(y[2719]), .A(x[2719]), .Z(n20185) );
  ANDN U18313 ( .B(y[2720]), .A(x[2720]), .Z(n20191) );
  OR U18314 ( .A(n20185), .B(n20191), .Z(n28127) );
  OR U18315 ( .A(n9527), .B(n28127), .Z(n9528) );
  AND U18316 ( .A(n9529), .B(n9528), .Z(n9530) );
  NANDN U18317 ( .A(x[2722]), .B(y[2722]), .Z(n28132) );
  ANDN U18318 ( .B(y[2721]), .A(x[2721]), .Z(n20190) );
  ANDN U18319 ( .B(n28132), .A(n20190), .Z(n28131) );
  NANDN U18320 ( .A(n9530), .B(n28131), .Z(n9531) );
  NAND U18321 ( .A(n28134), .B(n9531), .Z(n9532) );
  NANDN U18322 ( .A(n28135), .B(n9532), .Z(n9533) );
  NANDN U18323 ( .A(y[2724]), .B(x[2724]), .Z(n20200) );
  AND U18324 ( .A(n9533), .B(n20200), .Z(n9534) );
  NAND U18325 ( .A(n20206), .B(n9534), .Z(n9535) );
  NANDN U18326 ( .A(n28137), .B(n9535), .Z(n9536) );
  AND U18327 ( .A(n28138), .B(n9536), .Z(n9537) );
  NANDN U18328 ( .A(x[2727]), .B(y[2727]), .Z(n20210) );
  NANDN U18329 ( .A(x[2728]), .B(y[2728]), .Z(n20217) );
  AND U18330 ( .A(n20210), .B(n20217), .Z(n24182) );
  NANDN U18331 ( .A(n9537), .B(n24182), .Z(n9538) );
  NAND U18332 ( .A(n9539), .B(n9538), .Z(n9540) );
  NANDN U18333 ( .A(x[2729]), .B(y[2729]), .Z(n12456) );
  AND U18334 ( .A(n9540), .B(n12456), .Z(n9541) );
  NAND U18335 ( .A(n20221), .B(n9541), .Z(n9542) );
  NANDN U18336 ( .A(n28144), .B(n9542), .Z(n9543) );
  ANDN U18337 ( .B(x[2730]), .A(y[2730]), .Z(n12454) );
  OR U18338 ( .A(n9543), .B(n12454), .Z(n9544) );
  NAND U18339 ( .A(n9545), .B(n9544), .Z(n9546) );
  NANDN U18340 ( .A(n24181), .B(n9546), .Z(n9547) );
  NANDN U18341 ( .A(x[2733]), .B(y[2733]), .Z(n24180) );
  AND U18342 ( .A(n9547), .B(n24180), .Z(n9548) );
  NAND U18343 ( .A(n28146), .B(n9548), .Z(n9549) );
  AND U18344 ( .A(n28147), .B(n9549), .Z(n9551) );
  NANDN U18345 ( .A(x[2735]), .B(y[2735]), .Z(n28148) );
  ANDN U18346 ( .B(y[2736]), .A(x[2736]), .Z(n12450) );
  ANDN U18347 ( .B(n28148), .A(n12450), .Z(n9550) );
  NANDN U18348 ( .A(n9551), .B(n9550), .Z(n9552) );
  NANDN U18349 ( .A(n28149), .B(n9552), .Z(n9553) );
  AND U18350 ( .A(n12451), .B(n9553), .Z(n9554) );
  NANDN U18351 ( .A(n12448), .B(n9554), .Z(n9555) );
  NAND U18352 ( .A(n24177), .B(n9555), .Z(n9556) );
  NAND U18353 ( .A(n24176), .B(n9556), .Z(n9557) );
  NANDN U18354 ( .A(x[2740]), .B(y[2740]), .Z(n12447) );
  NANDN U18355 ( .A(n9557), .B(n12447), .Z(n9558) );
  AND U18356 ( .A(n9559), .B(n9558), .Z(n9561) );
  ANDN U18357 ( .B(y[2741]), .A(x[2741]), .Z(n12446) );
  XOR U18358 ( .A(y[2742]), .B(x[2742]), .Z(n20245) );
  NOR U18359 ( .A(n12446), .B(n20245), .Z(n9560) );
  NANDN U18360 ( .A(n9561), .B(n9560), .Z(n9562) );
  AND U18361 ( .A(n28155), .B(n9562), .Z(n9563) );
  NANDN U18362 ( .A(y[2743]), .B(x[2743]), .Z(n20248) );
  NAND U18363 ( .A(n9563), .B(n20248), .Z(n9564) );
  NAND U18364 ( .A(n20249), .B(n9564), .Z(n9565) );
  ANDN U18365 ( .B(y[2743]), .A(x[2743]), .Z(n12445) );
  OR U18366 ( .A(n9565), .B(n12445), .Z(n9566) );
  NAND U18367 ( .A(n9567), .B(n9566), .Z(n9568) );
  AND U18368 ( .A(n24172), .B(n9568), .Z(n9570) );
  NANDN U18369 ( .A(y[2746]), .B(x[2746]), .Z(n24173) );
  ANDN U18370 ( .B(x[2747]), .A(y[2747]), .Z(n12441) );
  ANDN U18371 ( .B(n24173), .A(n12441), .Z(n9569) );
  NANDN U18372 ( .A(n9570), .B(n9569), .Z(n9571) );
  NAND U18373 ( .A(n28159), .B(n9571), .Z(n9572) );
  XNOR U18374 ( .A(x[2748]), .B(y[2748]), .Z(n12442) );
  NANDN U18375 ( .A(n9572), .B(n12442), .Z(n9573) );
  AND U18376 ( .A(n9574), .B(n9573), .Z(n9575) );
  ANDN U18377 ( .B(y[2749]), .A(x[2749]), .Z(n20259) );
  NANDN U18378 ( .A(x[2750]), .B(y[2750]), .Z(n12440) );
  NANDN U18379 ( .A(n20259), .B(n12440), .Z(n28163) );
  OR U18380 ( .A(n9575), .B(n28163), .Z(n9576) );
  AND U18381 ( .A(n28164), .B(n9576), .Z(n9577) );
  NANDN U18382 ( .A(y[2751]), .B(x[2751]), .Z(n12439) );
  AND U18383 ( .A(n9577), .B(n12439), .Z(n9578) );
  NANDN U18384 ( .A(x[2751]), .B(y[2751]), .Z(n28165) );
  NANDN U18385 ( .A(n9578), .B(n28165), .Z(n9579) );
  XOR U18386 ( .A(x[2752]), .B(y[2752]), .Z(n12438) );
  OR U18387 ( .A(n9579), .B(n12438), .Z(n9580) );
  AND U18388 ( .A(n9581), .B(n9580), .Z(n9582) );
  NANDN U18389 ( .A(y[2753]), .B(x[2753]), .Z(n12435) );
  AND U18390 ( .A(n9582), .B(n12435), .Z(n9584) );
  NANDN U18391 ( .A(x[2754]), .B(y[2754]), .Z(n20271) );
  ANDN U18392 ( .B(y[2753]), .A(x[2753]), .Z(n12437) );
  ANDN U18393 ( .B(n20271), .A(n12437), .Z(n9583) );
  NANDN U18394 ( .A(n9584), .B(n9583), .Z(n9585) );
  AND U18395 ( .A(n12436), .B(n9585), .Z(n9588) );
  NANDN U18396 ( .A(x[2755]), .B(y[2755]), .Z(n9587) );
  NANDN U18397 ( .A(x[2756]), .B(y[2756]), .Z(n9586) );
  NAND U18398 ( .A(n9587), .B(n9586), .Z(n20268) );
  OR U18399 ( .A(n9588), .B(n20268), .Z(n9591) );
  NANDN U18400 ( .A(y[2756]), .B(x[2756]), .Z(n9590) );
  NANDN U18401 ( .A(y[2757]), .B(x[2757]), .Z(n9589) );
  NAND U18402 ( .A(n9590), .B(n9589), .Z(n12433) );
  ANDN U18403 ( .B(n9591), .A(n12433), .Z(n9593) );
  NANDN U18404 ( .A(x[2758]), .B(y[2758]), .Z(n12430) );
  NANDN U18405 ( .A(x[2757]), .B(y[2757]), .Z(n20269) );
  AND U18406 ( .A(n12430), .B(n20269), .Z(n9592) );
  NANDN U18407 ( .A(n9593), .B(n9592), .Z(n9594) );
  NAND U18408 ( .A(n12434), .B(n9594), .Z(n9595) );
  AND U18409 ( .A(n12432), .B(n9595), .Z(n9598) );
  NANDN U18410 ( .A(y[2760]), .B(x[2760]), .Z(n9597) );
  NANDN U18411 ( .A(y[2761]), .B(x[2761]), .Z(n9596) );
  NAND U18412 ( .A(n9597), .B(n9596), .Z(n20275) );
  OR U18413 ( .A(n9598), .B(n20275), .Z(n9601) );
  NANDN U18414 ( .A(x[2762]), .B(y[2762]), .Z(n9600) );
  NANDN U18415 ( .A(x[2761]), .B(y[2761]), .Z(n9599) );
  AND U18416 ( .A(n9600), .B(n9599), .Z(n20277) );
  AND U18417 ( .A(n9601), .B(n20277), .Z(n9604) );
  NANDN U18418 ( .A(y[2762]), .B(x[2762]), .Z(n9603) );
  NANDN U18419 ( .A(y[2763]), .B(x[2763]), .Z(n9602) );
  AND U18420 ( .A(n9603), .B(n9602), .Z(n28175) );
  NANDN U18421 ( .A(n9604), .B(n28175), .Z(n9605) );
  AND U18422 ( .A(n28176), .B(n9605), .Z(n9606) );
  OR U18423 ( .A(n28177), .B(n9606), .Z(n9607) );
  NAND U18424 ( .A(n28178), .B(n9607), .Z(n9608) );
  NANDN U18425 ( .A(n28179), .B(n9608), .Z(n9609) );
  NANDN U18426 ( .A(n24171), .B(n9609), .Z(n9610) );
  AND U18427 ( .A(n12425), .B(n9610), .Z(n9611) );
  NAND U18428 ( .A(n24170), .B(n9611), .Z(n9612) );
  ANDN U18429 ( .B(y[2769]), .A(x[2769]), .Z(n12426) );
  ANDN U18430 ( .B(n9612), .A(n12426), .Z(n9613) );
  NANDN U18431 ( .A(n12424), .B(n9613), .Z(n9614) );
  NANDN U18432 ( .A(y[2771]), .B(x[2771]), .Z(n28185) );
  AND U18433 ( .A(n9614), .B(n28185), .Z(n9615) );
  NANDN U18434 ( .A(n9616), .B(n9615), .Z(n9617) );
  NAND U18435 ( .A(n28187), .B(n9617), .Z(n9618) );
  NANDN U18436 ( .A(n28188), .B(n9618), .Z(n9619) );
  ANDN U18437 ( .B(y[2773]), .A(x[2773]), .Z(n28189) );
  ANDN U18438 ( .B(n9619), .A(n28189), .Z(n9620) );
  NANDN U18439 ( .A(n12421), .B(n9620), .Z(n9621) );
  NAND U18440 ( .A(n28190), .B(n9621), .Z(n9622) );
  NANDN U18441 ( .A(n12422), .B(n9622), .Z(n9623) );
  NANDN U18442 ( .A(y[2776]), .B(x[2776]), .Z(n20314) );
  NANDN U18443 ( .A(y[2777]), .B(x[2777]), .Z(n12417) );
  AND U18444 ( .A(n20314), .B(n12417), .Z(n24169) );
  AND U18445 ( .A(n9623), .B(n24169), .Z(n9625) );
  NANDN U18446 ( .A(x[2778]), .B(y[2778]), .Z(n12419) );
  NANDN U18447 ( .A(x[2777]), .B(y[2777]), .Z(n9624) );
  AND U18448 ( .A(n12419), .B(n9624), .Z(n28192) );
  NANDN U18449 ( .A(n9625), .B(n28192), .Z(n9626) );
  NAND U18450 ( .A(n28193), .B(n9626), .Z(n9627) );
  NANDN U18451 ( .A(n28197), .B(n9627), .Z(n9628) );
  OR U18452 ( .A(n28194), .B(n9628), .Z(n9629) );
  AND U18453 ( .A(n28195), .B(n9629), .Z(n9630) );
  OR U18454 ( .A(n28198), .B(n9630), .Z(n9631) );
  NAND U18455 ( .A(n28199), .B(n9631), .Z(n9632) );
  NANDN U18456 ( .A(n28200), .B(n9632), .Z(n9633) );
  NANDN U18457 ( .A(n24168), .B(n9633), .Z(n9634) );
  AND U18458 ( .A(n28202), .B(n9634), .Z(n9636) );
  NANDN U18459 ( .A(y[2786]), .B(x[2786]), .Z(n28203) );
  ANDN U18460 ( .B(x[2787]), .A(y[2787]), .Z(n12410) );
  ANDN U18461 ( .B(n28203), .A(n12410), .Z(n9635) );
  NANDN U18462 ( .A(n9636), .B(n9635), .Z(n9637) );
  NANDN U18463 ( .A(n24167), .B(n9637), .Z(n9638) );
  XNOR U18464 ( .A(x[2788]), .B(y[2788]), .Z(n12411) );
  NANDN U18465 ( .A(n9638), .B(n12411), .Z(n9639) );
  NAND U18466 ( .A(n9640), .B(n9639), .Z(n9641) );
  NANDN U18467 ( .A(n24166), .B(n9641), .Z(n9643) );
  NANDN U18468 ( .A(y[2791]), .B(x[2791]), .Z(n12407) );
  NANDN U18469 ( .A(y[2790]), .B(x[2790]), .Z(n24165) );
  AND U18470 ( .A(n12407), .B(n24165), .Z(n9642) );
  NAND U18471 ( .A(n9643), .B(n9642), .Z(n9644) );
  ANDN U18472 ( .B(y[2791]), .A(x[2791]), .Z(n28207) );
  ANDN U18473 ( .B(n9644), .A(n28207), .Z(n9645) );
  AND U18474 ( .A(n12408), .B(n9645), .Z(n9648) );
  ANDN U18475 ( .B(x[2793]), .A(y[2793]), .Z(n20354) );
  ANDN U18476 ( .B(x[2792]), .A(y[2792]), .Z(n9646) );
  NOR U18477 ( .A(n20354), .B(n9646), .Z(n9647) );
  NANDN U18478 ( .A(n9648), .B(n9647), .Z(n9649) );
  NANDN U18479 ( .A(n24162), .B(n9649), .Z(n9650) );
  NANDN U18480 ( .A(y[2794]), .B(x[2794]), .Z(n24163) );
  AND U18481 ( .A(n9650), .B(n24163), .Z(n9651) );
  NAND U18482 ( .A(n12405), .B(n9651), .Z(n9652) );
  NAND U18483 ( .A(n28210), .B(n9652), .Z(n9653) );
  XOR U18484 ( .A(x[2796]), .B(y[2796]), .Z(n12404) );
  OR U18485 ( .A(n9653), .B(n12404), .Z(n9654) );
  AND U18486 ( .A(n9655), .B(n9654), .Z(n9656) );
  NAND U18487 ( .A(n24161), .B(n9656), .Z(n9657) );
  ANDN U18488 ( .B(y[2797]), .A(x[2797]), .Z(n20360) );
  ANDN U18489 ( .B(n9657), .A(n20360), .Z(n9658) );
  NANDN U18490 ( .A(n12403), .B(n9658), .Z(n9659) );
  AND U18491 ( .A(n28216), .B(n9659), .Z(n9661) );
  NANDN U18492 ( .A(x[2799]), .B(y[2799]), .Z(n28217) );
  ANDN U18493 ( .B(y[2800]), .A(x[2800]), .Z(n20371) );
  ANDN U18494 ( .B(n28217), .A(n20371), .Z(n9660) );
  NANDN U18495 ( .A(n9661), .B(n9660), .Z(n9662) );
  NANDN U18496 ( .A(n20367), .B(n9662), .Z(n9663) );
  NAND U18497 ( .A(n28220), .B(n9663), .Z(n9664) );
  NANDN U18498 ( .A(x[2802]), .B(y[2802]), .Z(n12402) );
  NANDN U18499 ( .A(n9664), .B(n12402), .Z(n9665) );
  NAND U18500 ( .A(n28221), .B(n9665), .Z(n9666) );
  NANDN U18501 ( .A(n20381), .B(n9666), .Z(n9667) );
  ANDN U18502 ( .B(y[2803]), .A(x[2803]), .Z(n12401) );
  OR U18503 ( .A(n9667), .B(n12401), .Z(n9668) );
  AND U18504 ( .A(n28222), .B(n9668), .Z(n9669) );
  ANDN U18505 ( .B(y[2806]), .A(x[2806]), .Z(n20392) );
  NANDN U18506 ( .A(x[2805]), .B(y[2805]), .Z(n20382) );
  NANDN U18507 ( .A(n20392), .B(n20382), .Z(n24157) );
  OR U18508 ( .A(n9669), .B(n24157), .Z(n9670) );
  NAND U18509 ( .A(n28223), .B(n9670), .Z(n9671) );
  NANDN U18510 ( .A(n28224), .B(n9671), .Z(n9672) );
  NANDN U18511 ( .A(y[2809]), .B(x[2809]), .Z(n12396) );
  AND U18512 ( .A(n9672), .B(n12396), .Z(n9673) );
  NAND U18513 ( .A(n28227), .B(n9673), .Z(n9674) );
  NAND U18514 ( .A(n28229), .B(n9674), .Z(n9675) );
  AND U18515 ( .A(n12395), .B(n9675), .Z(n9676) );
  NANDN U18516 ( .A(y[2811]), .B(x[2811]), .Z(n12394) );
  NAND U18517 ( .A(n9676), .B(n12394), .Z(n9677) );
  ANDN U18518 ( .B(y[2812]), .A(x[2812]), .Z(n20403) );
  ANDN U18519 ( .B(n9677), .A(n20403), .Z(n9678) );
  NANDN U18520 ( .A(n28231), .B(n9678), .Z(n9679) );
  NANDN U18521 ( .A(y[2812]), .B(x[2812]), .Z(n28230) );
  AND U18522 ( .A(n9679), .B(n28230), .Z(n9680) );
  NAND U18523 ( .A(n12393), .B(n9680), .Z(n9681) );
  NANDN U18524 ( .A(n12390), .B(n9681), .Z(n9682) );
  ANDN U18525 ( .B(y[2813]), .A(x[2813]), .Z(n20402) );
  OR U18526 ( .A(n9682), .B(n20402), .Z(n9683) );
  NANDN U18527 ( .A(y[2815]), .B(x[2815]), .Z(n28235) );
  AND U18528 ( .A(n9683), .B(n28235), .Z(n9684) );
  NANDN U18529 ( .A(n12392), .B(n9684), .Z(n9685) );
  NAND U18530 ( .A(n28236), .B(n9685), .Z(n9686) );
  NAND U18531 ( .A(n28237), .B(n9686), .Z(n9687) );
  ANDN U18532 ( .B(x[2817]), .A(y[2817]), .Z(n12389) );
  OR U18533 ( .A(n9687), .B(n12389), .Z(n9688) );
  AND U18534 ( .A(n9689), .B(n9688), .Z(n9692) );
  NANDN U18535 ( .A(y[2819]), .B(x[2819]), .Z(n28240) );
  ANDN U18536 ( .B(x[2818]), .A(y[2818]), .Z(n9690) );
  ANDN U18537 ( .B(n28240), .A(n9690), .Z(n9691) );
  NANDN U18538 ( .A(n9692), .B(n9691), .Z(n9693) );
  ANDN U18539 ( .B(y[2820]), .A(x[2820]), .Z(n28241) );
  ANDN U18540 ( .B(n9693), .A(n28241), .Z(n9694) );
  NANDN U18541 ( .A(x[2819]), .B(y[2819]), .Z(n20414) );
  NAND U18542 ( .A(n9694), .B(n20414), .Z(n9695) );
  NANDN U18543 ( .A(n28243), .B(n9695), .Z(n9696) );
  AND U18544 ( .A(n28244), .B(n9696), .Z(n9697) );
  NANDN U18545 ( .A(y[2822]), .B(x[2822]), .Z(n12387) );
  NANDN U18546 ( .A(y[2823]), .B(x[2823]), .Z(n12385) );
  NAND U18547 ( .A(n12387), .B(n12385), .Z(n28245) );
  OR U18548 ( .A(n9697), .B(n28245), .Z(n9698) );
  AND U18549 ( .A(n9699), .B(n9698), .Z(n9700) );
  ANDN U18550 ( .B(n9701), .A(n9700), .Z(n9704) );
  NANDN U18551 ( .A(x[2826]), .B(y[2826]), .Z(n9703) );
  AND U18552 ( .A(n9703), .B(n9702), .Z(n28250) );
  NANDN U18553 ( .A(n9704), .B(n28250), .Z(n9705) );
  NAND U18554 ( .A(n28251), .B(n9705), .Z(n9706) );
  NAND U18555 ( .A(n20436), .B(n9706), .Z(n9707) );
  NANDN U18556 ( .A(y[2829]), .B(x[2829]), .Z(n12382) );
  NAND U18557 ( .A(n9707), .B(n12382), .Z(n9708) );
  NANDN U18558 ( .A(x[2830]), .B(y[2830]), .Z(n12380) );
  AND U18559 ( .A(n9708), .B(n12380), .Z(n9709) );
  NANDN U18560 ( .A(n20435), .B(n9709), .Z(n9710) );
  NANDN U18561 ( .A(y[2830]), .B(x[2830]), .Z(n12381) );
  AND U18562 ( .A(n9710), .B(n12381), .Z(n9711) );
  NAND U18563 ( .A(n20441), .B(n9711), .Z(n9712) );
  NANDN U18564 ( .A(n28255), .B(n9712), .Z(n9713) );
  ANDN U18565 ( .B(y[2831]), .A(x[2831]), .Z(n12379) );
  OR U18566 ( .A(n9713), .B(n12379), .Z(n9714) );
  NAND U18567 ( .A(n9715), .B(n9714), .Z(n9716) );
  NANDN U18568 ( .A(n28260), .B(n9716), .Z(n9717) );
  NANDN U18569 ( .A(y[2834]), .B(x[2834]), .Z(n28261) );
  AND U18570 ( .A(n9717), .B(n28261), .Z(n9718) );
  NAND U18571 ( .A(n12376), .B(n9718), .Z(n9719) );
  NAND U18572 ( .A(n28259), .B(n9719), .Z(n9720) );
  XOR U18573 ( .A(x[2836]), .B(y[2836]), .Z(n12375) );
  OR U18574 ( .A(n9720), .B(n12375), .Z(n9721) );
  NAND U18575 ( .A(n9722), .B(n9721), .Z(n9723) );
  NANDN U18576 ( .A(n28271), .B(n9723), .Z(n9724) );
  NANDN U18577 ( .A(y[2838]), .B(x[2838]), .Z(n28273) );
  AND U18578 ( .A(n9724), .B(n28273), .Z(n9725) );
  NAND U18579 ( .A(n12373), .B(n9725), .Z(n9726) );
  NAND U18580 ( .A(n28274), .B(n9726), .Z(n9727) );
  XOR U18581 ( .A(x[2840]), .B(y[2840]), .Z(n12372) );
  OR U18582 ( .A(n9727), .B(n12372), .Z(n9728) );
  AND U18583 ( .A(n9729), .B(n9728), .Z(n9730) );
  NANDN U18584 ( .A(n20459), .B(n9730), .Z(n9731) );
  AND U18585 ( .A(n9732), .B(n9731), .Z(n9733) );
  OR U18586 ( .A(n28285), .B(n9733), .Z(n9734) );
  NAND U18587 ( .A(n28287), .B(n9734), .Z(n9735) );
  NANDN U18588 ( .A(n28288), .B(n9735), .Z(n9737) );
  NANDN U18589 ( .A(x[2846]), .B(y[2846]), .Z(n20475) );
  ANDN U18590 ( .B(y[2845]), .A(x[2845]), .Z(n28290) );
  ANDN U18591 ( .B(n20475), .A(n28290), .Z(n9736) );
  NAND U18592 ( .A(n9737), .B(n9736), .Z(n9738) );
  AND U18593 ( .A(n28292), .B(n9738), .Z(n9743) );
  NANDN U18594 ( .A(x[2848]), .B(y[2848]), .Z(n9740) );
  NANDN U18595 ( .A(x[2847]), .B(y[2847]), .Z(n9739) );
  AND U18596 ( .A(n9740), .B(n9739), .Z(n9742) );
  NAND U18597 ( .A(n9742), .B(n9741), .Z(n20476) );
  OR U18598 ( .A(n9743), .B(n20476), .Z(n9744) );
  NAND U18599 ( .A(n28297), .B(n9744), .Z(n9745) );
  NAND U18600 ( .A(n28298), .B(n9745), .Z(n9746) );
  AND U18601 ( .A(n28299), .B(n9746), .Z(n9747) );
  OR U18602 ( .A(n28300), .B(n9747), .Z(n9748) );
  NAND U18603 ( .A(n28301), .B(n9748), .Z(n9749) );
  NANDN U18604 ( .A(n28302), .B(n9749), .Z(n9750) );
  NANDN U18605 ( .A(y[2854]), .B(x[2854]), .Z(n20487) );
  NANDN U18606 ( .A(y[2855]), .B(x[2855]), .Z(n20495) );
  AND U18607 ( .A(n20487), .B(n20495), .Z(n24151) );
  AND U18608 ( .A(n9750), .B(n24151), .Z(n9751) );
  ANDN U18609 ( .B(y[2855]), .A(x[2855]), .Z(n20491) );
  NANDN U18610 ( .A(x[2856]), .B(y[2856]), .Z(n12359) );
  NANDN U18611 ( .A(n20491), .B(n12359), .Z(n28303) );
  OR U18612 ( .A(n9751), .B(n28303), .Z(n9752) );
  NANDN U18613 ( .A(y[2856]), .B(x[2856]), .Z(n12360) );
  AND U18614 ( .A(n9752), .B(n12360), .Z(n9753) );
  NANDN U18615 ( .A(y[2857]), .B(x[2857]), .Z(n12357) );
  NAND U18616 ( .A(n9753), .B(n12357), .Z(n9754) );
  ANDN U18617 ( .B(y[2857]), .A(x[2857]), .Z(n12358) );
  ANDN U18618 ( .B(n9754), .A(n12358), .Z(n9755) );
  NANDN U18619 ( .A(n12356), .B(n9755), .Z(n9757) );
  NANDN U18620 ( .A(y[2858]), .B(x[2858]), .Z(n9756) );
  AND U18621 ( .A(n9757), .B(n9756), .Z(n9758) );
  NAND U18622 ( .A(n12354), .B(n9758), .Z(n9759) );
  NANDN U18623 ( .A(n12355), .B(n9759), .Z(n9760) );
  ANDN U18624 ( .B(y[2860]), .A(x[2860]), .Z(n12351) );
  OR U18625 ( .A(n9760), .B(n12351), .Z(n9761) );
  AND U18626 ( .A(n12353), .B(n9761), .Z(n9762) );
  NANDN U18627 ( .A(y[2861]), .B(x[2861]), .Z(n12350) );
  AND U18628 ( .A(n9762), .B(n12350), .Z(n9763) );
  NANDN U18629 ( .A(x[2861]), .B(y[2861]), .Z(n12352) );
  NANDN U18630 ( .A(n9763), .B(n12352), .Z(n9764) );
  ANDN U18631 ( .B(y[2862]), .A(x[2862]), .Z(n20504) );
  OR U18632 ( .A(n9764), .B(n20504), .Z(n9765) );
  NANDN U18633 ( .A(y[2863]), .B(x[2863]), .Z(n24150) );
  AND U18634 ( .A(n9765), .B(n24150), .Z(n9766) );
  NANDN U18635 ( .A(n12349), .B(n9766), .Z(n9767) );
  AND U18636 ( .A(n9768), .B(n9767), .Z(n9769) );
  OR U18637 ( .A(n28314), .B(n9769), .Z(n9770) );
  NAND U18638 ( .A(n28315), .B(n9770), .Z(n9771) );
  NANDN U18639 ( .A(n28316), .B(n9771), .Z(n9772) );
  NANDN U18640 ( .A(x[2868]), .B(y[2868]), .Z(n12344) );
  AND U18641 ( .A(n9772), .B(n12344), .Z(n9773) );
  NAND U18642 ( .A(n28317), .B(n9773), .Z(n9774) );
  NANDN U18643 ( .A(n9775), .B(n9774), .Z(n9776) );
  NANDN U18644 ( .A(x[2870]), .B(y[2870]), .Z(n20524) );
  AND U18645 ( .A(n9776), .B(n20524), .Z(n9777) );
  NANDN U18646 ( .A(x[2869]), .B(y[2869]), .Z(n12343) );
  AND U18647 ( .A(n9777), .B(n12343), .Z(n9778) );
  NANDN U18648 ( .A(y[2870]), .B(x[2870]), .Z(n12342) );
  NANDN U18649 ( .A(y[2871]), .B(x[2871]), .Z(n12340) );
  AND U18650 ( .A(n12342), .B(n12340), .Z(n28322) );
  NANDN U18651 ( .A(n9778), .B(n28322), .Z(n9779) );
  NANDN U18652 ( .A(n28323), .B(n9779), .Z(n9780) );
  AND U18653 ( .A(n28324), .B(n9780), .Z(n9781) );
  OR U18654 ( .A(n28325), .B(n9781), .Z(n9782) );
  NAND U18655 ( .A(n24149), .B(n9782), .Z(n9783) );
  NANDN U18656 ( .A(n28326), .B(n9783), .Z(n9784) );
  NANDN U18657 ( .A(n28327), .B(n9784), .Z(n9785) );
  AND U18658 ( .A(n28328), .B(n9785), .Z(n9787) );
  ANDN U18659 ( .B(x[2879]), .A(y[2879]), .Z(n12332) );
  ANDN U18660 ( .B(x[2878]), .A(y[2878]), .Z(n28329) );
  NOR U18661 ( .A(n12332), .B(n28329), .Z(n9786) );
  NANDN U18662 ( .A(n9787), .B(n9786), .Z(n9788) );
  NANDN U18663 ( .A(n24148), .B(n9788), .Z(n9789) );
  XNOR U18664 ( .A(x[2880]), .B(y[2880]), .Z(n12333) );
  NANDN U18665 ( .A(n9789), .B(n12333), .Z(n9790) );
  AND U18666 ( .A(n9791), .B(n9790), .Z(n9794) );
  NANDN U18667 ( .A(x[2882]), .B(y[2882]), .Z(n9793) );
  NANDN U18668 ( .A(x[2881]), .B(y[2881]), .Z(n9792) );
  NAND U18669 ( .A(n9793), .B(n9792), .Z(n28334) );
  OR U18670 ( .A(n9794), .B(n28334), .Z(n9795) );
  AND U18671 ( .A(n28335), .B(n9795), .Z(n9796) );
  NANDN U18672 ( .A(n12330), .B(n9796), .Z(n9797) );
  AND U18673 ( .A(n9798), .B(n9797), .Z(n9801) );
  ANDN U18674 ( .B(x[2885]), .A(y[2885]), .Z(n20557) );
  ANDN U18675 ( .B(x[2884]), .A(y[2884]), .Z(n9799) );
  NOR U18676 ( .A(n20557), .B(n9799), .Z(n9800) );
  NANDN U18677 ( .A(n9801), .B(n9800), .Z(n9802) );
  NANDN U18678 ( .A(x[2886]), .B(y[2886]), .Z(n12327) );
  AND U18679 ( .A(n9802), .B(n12327), .Z(n9803) );
  NANDN U18680 ( .A(x[2885]), .B(y[2885]), .Z(n12328) );
  NAND U18681 ( .A(n9803), .B(n12328), .Z(n9804) );
  NANDN U18682 ( .A(n24147), .B(n9804), .Z(n9805) );
  AND U18683 ( .A(n28341), .B(n9805), .Z(n9807) );
  NANDN U18684 ( .A(y[2888]), .B(x[2888]), .Z(n9806) );
  ANDN U18685 ( .B(x[2889]), .A(y[2889]), .Z(n12325) );
  ANDN U18686 ( .B(n9806), .A(n12325), .Z(n28342) );
  NANDN U18687 ( .A(n9807), .B(n28342), .Z(n9808) );
  AND U18688 ( .A(n9809), .B(n9808), .Z(n9811) );
  NANDN U18689 ( .A(y[2890]), .B(x[2890]), .Z(n28344) );
  ANDN U18690 ( .B(x[2891]), .A(y[2891]), .Z(n12319) );
  ANDN U18691 ( .B(n28344), .A(n12319), .Z(n9810) );
  NANDN U18692 ( .A(n9811), .B(n9810), .Z(n9812) );
  NANDN U18693 ( .A(x[2892]), .B(y[2892]), .Z(n20575) );
  AND U18694 ( .A(n9812), .B(n20575), .Z(n9813) );
  NANDN U18695 ( .A(x[2891]), .B(y[2891]), .Z(n12321) );
  NAND U18696 ( .A(n9813), .B(n12321), .Z(n9814) );
  NANDN U18697 ( .A(n28349), .B(n9814), .Z(n9815) );
  AND U18698 ( .A(n28350), .B(n9815), .Z(n9816) );
  ANDN U18699 ( .B(x[2894]), .A(y[2894]), .Z(n12318) );
  ANDN U18700 ( .B(x[2895]), .A(y[2895]), .Z(n20584) );
  OR U18701 ( .A(n12318), .B(n20584), .Z(n24146) );
  OR U18702 ( .A(n9816), .B(n24146), .Z(n9817) );
  NANDN U18703 ( .A(x[2895]), .B(y[2895]), .Z(n20580) );
  NANDN U18704 ( .A(x[2896]), .B(y[2896]), .Z(n12316) );
  AND U18705 ( .A(n20580), .B(n12316), .Z(n24145) );
  AND U18706 ( .A(n9817), .B(n24145), .Z(n9819) );
  ANDN U18707 ( .B(x[2897]), .A(y[2897]), .Z(n12314) );
  ANDN U18708 ( .B(x[2896]), .A(y[2896]), .Z(n28351) );
  NOR U18709 ( .A(n12314), .B(n28351), .Z(n9818) );
  NANDN U18710 ( .A(n9819), .B(n9818), .Z(n9820) );
  AND U18711 ( .A(n28352), .B(n9820), .Z(n9821) );
  AND U18712 ( .A(n12315), .B(n9821), .Z(n9824) );
  NANDN U18713 ( .A(y[2899]), .B(x[2899]), .Z(n28355) );
  ANDN U18714 ( .B(x[2898]), .A(y[2898]), .Z(n9822) );
  ANDN U18715 ( .B(n28355), .A(n9822), .Z(n9823) );
  NANDN U18716 ( .A(n9824), .B(n9823), .Z(n9825) );
  NANDN U18717 ( .A(n24144), .B(n9825), .Z(n9826) );
  NANDN U18718 ( .A(y[2900]), .B(x[2900]), .Z(n24143) );
  AND U18719 ( .A(n9826), .B(n24143), .Z(n9827) );
  NAND U18720 ( .A(n12311), .B(n9827), .Z(n9828) );
  NANDN U18721 ( .A(n12312), .B(n9828), .Z(n9829) );
  XOR U18722 ( .A(x[2902]), .B(y[2902]), .Z(n12310) );
  OR U18723 ( .A(n9829), .B(n12310), .Z(n9830) );
  AND U18724 ( .A(n9831), .B(n9830), .Z(n9832) );
  NANDN U18725 ( .A(x[2903]), .B(y[2903]), .Z(n20598) );
  NANDN U18726 ( .A(x[2904]), .B(y[2904]), .Z(n20604) );
  NAND U18727 ( .A(n20598), .B(n20604), .Z(n28361) );
  OR U18728 ( .A(n9832), .B(n28361), .Z(n9833) );
  NANDN U18729 ( .A(y[2904]), .B(x[2904]), .Z(n20601) );
  AND U18730 ( .A(n9833), .B(n20601), .Z(n9834) );
  NANDN U18731 ( .A(n12307), .B(n9834), .Z(n9835) );
  ANDN U18732 ( .B(y[2905]), .A(x[2905]), .Z(n28364) );
  ANDN U18733 ( .B(n9835), .A(n28364), .Z(n9836) );
  NAND U18734 ( .A(n12308), .B(n9836), .Z(n9837) );
  NANDN U18735 ( .A(y[2907]), .B(x[2907]), .Z(n28367) );
  AND U18736 ( .A(n9837), .B(n28367), .Z(n9838) );
  NANDN U18737 ( .A(n9839), .B(n9838), .Z(n9840) );
  ANDN U18738 ( .B(y[2908]), .A(x[2908]), .Z(n28368) );
  ANDN U18739 ( .B(n9840), .A(n28368), .Z(n9841) );
  NANDN U18740 ( .A(n20607), .B(n9841), .Z(n9842) );
  NAND U18741 ( .A(n28369), .B(n9842), .Z(n9843) );
  NANDN U18742 ( .A(n12304), .B(n9843), .Z(n9844) );
  ANDN U18743 ( .B(y[2909]), .A(x[2909]), .Z(n28370) );
  OR U18744 ( .A(n9844), .B(n28370), .Z(n9845) );
  NANDN U18745 ( .A(y[2910]), .B(x[2910]), .Z(n12305) );
  NANDN U18746 ( .A(y[2911]), .B(x[2911]), .Z(n20618) );
  AND U18747 ( .A(n12305), .B(n20618), .Z(n28372) );
  AND U18748 ( .A(n9845), .B(n28372), .Z(n9847) );
  ANDN U18749 ( .B(y[2911]), .A(x[2911]), .Z(n12303) );
  ANDN U18750 ( .B(y[2912]), .A(x[2912]), .Z(n12300) );
  NOR U18751 ( .A(n12303), .B(n12300), .Z(n9846) );
  NANDN U18752 ( .A(n9847), .B(n9846), .Z(n9848) );
  NAND U18753 ( .A(n24142), .B(n9848), .Z(n9849) );
  NAND U18754 ( .A(n12302), .B(n9849), .Z(n9850) );
  NAND U18755 ( .A(n24140), .B(n9850), .Z(n9851) );
  NANDN U18756 ( .A(n28376), .B(n9851), .Z(n9852) );
  AND U18757 ( .A(n12298), .B(n9852), .Z(n9853) );
  ANDN U18758 ( .B(y[2918]), .A(x[2918]), .Z(n12295) );
  OR U18759 ( .A(n9853), .B(n12295), .Z(n9854) );
  AND U18760 ( .A(n9855), .B(n9854), .Z(n9857) );
  NANDN U18761 ( .A(x[2919]), .B(y[2919]), .Z(n12296) );
  ANDN U18762 ( .B(y[2920]), .A(x[2920]), .Z(n24139) );
  ANDN U18763 ( .B(n12296), .A(n24139), .Z(n9856) );
  NANDN U18764 ( .A(n9857), .B(n9856), .Z(n9858) );
  AND U18765 ( .A(n28381), .B(n9858), .Z(n9859) );
  NANDN U18766 ( .A(y[2920]), .B(x[2920]), .Z(n12294) );
  AND U18767 ( .A(n9859), .B(n12294), .Z(n9860) );
  NANDN U18768 ( .A(x[2922]), .B(y[2922]), .Z(n20633) );
  ANDN U18769 ( .B(y[2921]), .A(x[2921]), .Z(n20628) );
  ANDN U18770 ( .B(n20633), .A(n20628), .Z(n28382) );
  NANDN U18771 ( .A(n9860), .B(n28382), .Z(n9861) );
  NAND U18772 ( .A(n9862), .B(n9861), .Z(n9863) );
  AND U18773 ( .A(n12291), .B(n9863), .Z(n9864) );
  NAND U18774 ( .A(n12292), .B(n9864), .Z(n9865) );
  NANDN U18775 ( .A(n24138), .B(n9865), .Z(n9866) );
  OR U18776 ( .A(n9867), .B(n9866), .Z(n9868) );
  NANDN U18777 ( .A(x[2925]), .B(y[2925]), .Z(n20638) );
  NANDN U18778 ( .A(x[2926]), .B(y[2926]), .Z(n20642) );
  AND U18779 ( .A(n20638), .B(n20642), .Z(n24137) );
  AND U18780 ( .A(n9868), .B(n24137), .Z(n9870) );
  NANDN U18781 ( .A(y[2927]), .B(x[2927]), .Z(n12288) );
  ANDN U18782 ( .B(x[2926]), .A(y[2926]), .Z(n28387) );
  ANDN U18783 ( .B(n12288), .A(n28387), .Z(n9869) );
  NANDN U18784 ( .A(n9870), .B(n9869), .Z(n9871) );
  NANDN U18785 ( .A(n28388), .B(n9871), .Z(n9872) );
  XNOR U18786 ( .A(x[2928]), .B(y[2928]), .Z(n12289) );
  NANDN U18787 ( .A(n9872), .B(n12289), .Z(n9873) );
  ANDN U18788 ( .B(x[2929]), .A(y[2929]), .Z(n28392) );
  ANDN U18789 ( .B(n9873), .A(n28392), .Z(n9874) );
  NANDN U18790 ( .A(n9875), .B(n9874), .Z(n9876) );
  AND U18791 ( .A(n9877), .B(n9876), .Z(n9878) );
  NANDN U18792 ( .A(y[2930]), .B(x[2930]), .Z(n20649) );
  NANDN U18793 ( .A(y[2931]), .B(x[2931]), .Z(n12287) );
  AND U18794 ( .A(n20649), .B(n12287), .Z(n28394) );
  NANDN U18795 ( .A(n9878), .B(n28394), .Z(n9879) );
  AND U18796 ( .A(n28395), .B(n9879), .Z(n9880) );
  NANDN U18797 ( .A(x[2932]), .B(y[2932]), .Z(n28396) );
  AND U18798 ( .A(n9880), .B(n28396), .Z(n9881) );
  NANDN U18799 ( .A(y[2932]), .B(x[2932]), .Z(n12286) );
  ANDN U18800 ( .B(x[2933]), .A(y[2933]), .Z(n20658) );
  ANDN U18801 ( .B(n12286), .A(n20658), .Z(n28397) );
  NANDN U18802 ( .A(n9881), .B(n28397), .Z(n9882) );
  NAND U18803 ( .A(n9883), .B(n9882), .Z(n9884) );
  AND U18804 ( .A(n28399), .B(n9884), .Z(n9886) );
  NANDN U18805 ( .A(x[2935]), .B(y[2935]), .Z(n12283) );
  ANDN U18806 ( .B(y[2936]), .A(x[2936]), .Z(n24136) );
  ANDN U18807 ( .B(n12283), .A(n24136), .Z(n9885) );
  NANDN U18808 ( .A(n9886), .B(n9885), .Z(n9887) );
  NANDN U18809 ( .A(y[2936]), .B(x[2936]), .Z(n20663) );
  NANDN U18810 ( .A(y[2937]), .B(x[2937]), .Z(n12282) );
  AND U18811 ( .A(n20663), .B(n12282), .Z(n28400) );
  AND U18812 ( .A(n9887), .B(n28400), .Z(n9888) );
  ANDN U18813 ( .B(y[2937]), .A(x[2937]), .Z(n20666) );
  ANDN U18814 ( .B(y[2938]), .A(x[2938]), .Z(n20672) );
  OR U18815 ( .A(n20666), .B(n20672), .Z(n24133) );
  OR U18816 ( .A(n9888), .B(n24133), .Z(n9889) );
  NAND U18817 ( .A(n24132), .B(n9889), .Z(n9890) );
  NANDN U18818 ( .A(n28402), .B(n9890), .Z(n9891) );
  AND U18819 ( .A(n28403), .B(n9891), .Z(n9892) );
  OR U18820 ( .A(n28404), .B(n9892), .Z(n9893) );
  NAND U18821 ( .A(n28405), .B(n9893), .Z(n9894) );
  NAND U18822 ( .A(n28406), .B(n9894), .Z(n9895) );
  NANDN U18823 ( .A(n28407), .B(n9895), .Z(n9896) );
  NANDN U18824 ( .A(y[2945]), .B(x[2945]), .Z(n12271) );
  NANDN U18825 ( .A(n9896), .B(n12271), .Z(n9897) );
  NAND U18826 ( .A(n28408), .B(n9897), .Z(n9898) );
  NANDN U18827 ( .A(n24131), .B(n9898), .Z(n9899) );
  ANDN U18828 ( .B(x[2946]), .A(y[2946]), .Z(n12270) );
  OR U18829 ( .A(n9899), .B(n12270), .Z(n9900) );
  NAND U18830 ( .A(n28409), .B(n9900), .Z(n9901) );
  NANDN U18831 ( .A(n28410), .B(n9901), .Z(n9902) );
  NANDN U18832 ( .A(x[2949]), .B(y[2949]), .Z(n28411) );
  AND U18833 ( .A(n9902), .B(n28411), .Z(n9903) );
  NANDN U18834 ( .A(x[2950]), .B(y[2950]), .Z(n12268) );
  AND U18835 ( .A(n9903), .B(n12268), .Z(n9904) );
  ANDN U18836 ( .B(x[2950]), .A(y[2950]), .Z(n20698) );
  ANDN U18837 ( .B(x[2951]), .A(y[2951]), .Z(n28414) );
  OR U18838 ( .A(n20698), .B(n28414), .Z(n24128) );
  OR U18839 ( .A(n9904), .B(n24128), .Z(n9905) );
  AND U18840 ( .A(n9906), .B(n9905), .Z(n9907) );
  OR U18841 ( .A(n28416), .B(n9907), .Z(n9908) );
  NAND U18842 ( .A(n28417), .B(n9908), .Z(n9909) );
  NANDN U18843 ( .A(n28418), .B(n9909), .Z(n9910) );
  ANDN U18844 ( .B(y[2955]), .A(x[2955]), .Z(n28419) );
  ANDN U18845 ( .B(n9910), .A(n28419), .Z(n9911) );
  NANDN U18846 ( .A(x[2956]), .B(y[2956]), .Z(n12264) );
  AND U18847 ( .A(n9911), .B(n12264), .Z(n9912) );
  OR U18848 ( .A(n9913), .B(n9912), .Z(n9914) );
  AND U18849 ( .A(n9915), .B(n9914), .Z(n9916) );
  ANDN U18850 ( .B(x[2958]), .A(y[2958]), .Z(n20718) );
  ANDN U18851 ( .B(x[2959]), .A(y[2959]), .Z(n20722) );
  OR U18852 ( .A(n20718), .B(n20722), .Z(n24125) );
  OR U18853 ( .A(n9916), .B(n24125), .Z(n9917) );
  NAND U18854 ( .A(n24124), .B(n9917), .Z(n9918) );
  NANDN U18855 ( .A(n24123), .B(n9918), .Z(n9919) );
  AND U18856 ( .A(n28423), .B(n9919), .Z(n9921) );
  NANDN U18857 ( .A(y[2963]), .B(x[2963]), .Z(n20733) );
  NANDN U18858 ( .A(y[2962]), .B(x[2962]), .Z(n12258) );
  AND U18859 ( .A(n20733), .B(n12258), .Z(n9920) );
  NANDN U18860 ( .A(n9921), .B(n9920), .Z(n9922) );
  NAND U18861 ( .A(n9923), .B(n9922), .Z(n9924) );
  AND U18862 ( .A(n9925), .B(n9924), .Z(n9926) );
  NANDN U18863 ( .A(y[2965]), .B(x[2965]), .Z(n12257) );
  NAND U18864 ( .A(n9926), .B(n12257), .Z(n9927) );
  NANDN U18865 ( .A(n28432), .B(n9927), .Z(n9928) );
  NANDN U18866 ( .A(y[2966]), .B(x[2966]), .Z(n28431) );
  AND U18867 ( .A(n9928), .B(n28431), .Z(n9929) );
  NANDN U18868 ( .A(y[2967]), .B(x[2967]), .Z(n12255) );
  AND U18869 ( .A(n9929), .B(n12255), .Z(n9931) );
  NANDN U18870 ( .A(x[2967]), .B(y[2967]), .Z(n28430) );
  NANDN U18871 ( .A(x[2968]), .B(y[2968]), .Z(n28434) );
  AND U18872 ( .A(n28430), .B(n28434), .Z(n9930) );
  NANDN U18873 ( .A(n9931), .B(n9930), .Z(n9932) );
  NAND U18874 ( .A(n9933), .B(n9932), .Z(n9934) );
  AND U18875 ( .A(n28436), .B(n9934), .Z(n9935) );
  ANDN U18876 ( .B(x[2970]), .A(y[2970]), .Z(n20745) );
  NANDN U18877 ( .A(y[2971]), .B(x[2971]), .Z(n12250) );
  NANDN U18878 ( .A(n20745), .B(n12250), .Z(n28437) );
  OR U18879 ( .A(n9935), .B(n28437), .Z(n9936) );
  NANDN U18880 ( .A(x[2971]), .B(y[2971]), .Z(n12251) );
  AND U18881 ( .A(n9936), .B(n12251), .Z(n9937) );
  NANDN U18882 ( .A(x[2972]), .B(y[2972]), .Z(n12246) );
  AND U18883 ( .A(n9937), .B(n12246), .Z(n9939) );
  ANDN U18884 ( .B(x[2973]), .A(y[2973]), .Z(n12245) );
  NANDN U18885 ( .A(y[2972]), .B(x[2972]), .Z(n9938) );
  NANDN U18886 ( .A(n12245), .B(n9938), .Z(n12249) );
  OR U18887 ( .A(n9939), .B(n12249), .Z(n9940) );
  NAND U18888 ( .A(n12248), .B(n9940), .Z(n9941) );
  NANDN U18889 ( .A(n20752), .B(n9941), .Z(n9942) );
  NANDN U18890 ( .A(x[2975]), .B(y[2975]), .Z(n20754) );
  AND U18891 ( .A(n9942), .B(n20754), .Z(n9943) );
  NANDN U18892 ( .A(x[2976]), .B(y[2976]), .Z(n12243) );
  AND U18893 ( .A(n9943), .B(n12243), .Z(n9945) );
  NANDN U18894 ( .A(y[2976]), .B(x[2976]), .Z(n9944) );
  ANDN U18895 ( .B(x[2977]), .A(y[2977]), .Z(n12244) );
  ANDN U18896 ( .B(n9944), .A(n12244), .Z(n24122) );
  NANDN U18897 ( .A(n9945), .B(n24122), .Z(n9946) );
  NAND U18898 ( .A(n9947), .B(n9946), .Z(n9949) );
  ANDN U18899 ( .B(x[2979]), .A(y[2979]), .Z(n12240) );
  NANDN U18900 ( .A(y[2978]), .B(x[2978]), .Z(n9948) );
  NANDN U18901 ( .A(n12240), .B(n9948), .Z(n20759) );
  IV U18902 ( .A(n20759), .Z(n28445) );
  AND U18903 ( .A(n9949), .B(n28445), .Z(n9951) );
  NANDN U18904 ( .A(x[2979]), .B(y[2979]), .Z(n12241) );
  ANDN U18905 ( .B(y[2980]), .A(x[2980]), .Z(n20764) );
  ANDN U18906 ( .B(n12241), .A(n20764), .Z(n9950) );
  NANDN U18907 ( .A(n9951), .B(n9950), .Z(n9952) );
  AND U18908 ( .A(n28448), .B(n9952), .Z(n9953) );
  OR U18909 ( .A(n28449), .B(n9953), .Z(n9954) );
  NAND U18910 ( .A(n28450), .B(n9954), .Z(n9955) );
  NANDN U18911 ( .A(n24120), .B(n9955), .Z(n9956) );
  NANDN U18912 ( .A(y[2984]), .B(x[2984]), .Z(n20774) );
  NANDN U18913 ( .A(y[2985]), .B(x[2985]), .Z(n20781) );
  AND U18914 ( .A(n20774), .B(n20781), .Z(n24119) );
  AND U18915 ( .A(n9956), .B(n24119), .Z(n9957) );
  NANDN U18916 ( .A(x[2985]), .B(y[2985]), .Z(n12235) );
  NANDN U18917 ( .A(x[2986]), .B(y[2986]), .Z(n12234) );
  NAND U18918 ( .A(n12235), .B(n12234), .Z(n28451) );
  OR U18919 ( .A(n9957), .B(n28451), .Z(n9958) );
  NAND U18920 ( .A(n28452), .B(n9958), .Z(n9959) );
  NANDN U18921 ( .A(x[2987]), .B(y[2987]), .Z(n12233) );
  NANDN U18922 ( .A(x[2988]), .B(y[2988]), .Z(n20792) );
  AND U18923 ( .A(n12233), .B(n20792), .Z(n28453) );
  AND U18924 ( .A(n9959), .B(n28453), .Z(n9961) );
  ANDN U18925 ( .B(x[2988]), .A(y[2988]), .Z(n20787) );
  IV U18926 ( .A(n20787), .Z(n28454) );
  ANDN U18927 ( .B(x[2989]), .A(y[2989]), .Z(n12232) );
  ANDN U18928 ( .B(n28454), .A(n12232), .Z(n9960) );
  NANDN U18929 ( .A(n9961), .B(n9960), .Z(n9962) );
  NANDN U18930 ( .A(n28455), .B(n9962), .Z(n9963) );
  AND U18931 ( .A(n24118), .B(n9963), .Z(n9964) );
  NANDN U18932 ( .A(n12231), .B(n9964), .Z(n9965) );
  NAND U18933 ( .A(n28458), .B(n9965), .Z(n9966) );
  NANDN U18934 ( .A(n24114), .B(n9966), .Z(n9967) );
  NANDN U18935 ( .A(x[2993]), .B(y[2993]), .Z(n20802) );
  AND U18936 ( .A(n9967), .B(n20802), .Z(n9968) );
  NANDN U18937 ( .A(x[2994]), .B(y[2994]), .Z(n12227) );
  AND U18938 ( .A(n9968), .B(n12227), .Z(n9970) );
  NANDN U18939 ( .A(y[2995]), .B(x[2995]), .Z(n12228) );
  NANDN U18940 ( .A(y[2994]), .B(x[2994]), .Z(n9969) );
  NAND U18941 ( .A(n12228), .B(n9969), .Z(n20804) );
  OR U18942 ( .A(n9970), .B(n20804), .Z(n9971) );
  NAND U18943 ( .A(n12229), .B(n9971), .Z(n9972) );
  NANDN U18944 ( .A(n20810), .B(n9972), .Z(n9973) );
  AND U18945 ( .A(n20811), .B(n9973), .Z(n9974) );
  NANDN U18946 ( .A(x[3000]), .B(y[3000]), .Z(n12226) );
  AND U18947 ( .A(n9974), .B(n12226), .Z(n9976) );
  NANDN U18948 ( .A(y[3000]), .B(x[3000]), .Z(n28463) );
  NANDN U18949 ( .A(y[3001]), .B(x[3001]), .Z(n28465) );
  NAND U18950 ( .A(n28463), .B(n28465), .Z(n9975) );
  OR U18951 ( .A(n9976), .B(n9975), .Z(n9977) );
  AND U18952 ( .A(n12225), .B(n9977), .Z(n9978) );
  NANDN U18953 ( .A(x[3002]), .B(y[3002]), .Z(n28466) );
  AND U18954 ( .A(n9978), .B(n28466), .Z(n9979) );
  OR U18955 ( .A(n28467), .B(n9979), .Z(n9980) );
  NAND U18956 ( .A(n9981), .B(n9980), .Z(n9982) );
  NANDN U18957 ( .A(y[3004]), .B(x[3004]), .Z(n28469) );
  AND U18958 ( .A(n9982), .B(n28469), .Z(n9983) );
  NANDN U18959 ( .A(y[3005]), .B(x[3005]), .Z(n20822) );
  NAND U18960 ( .A(n9983), .B(n20822), .Z(n9984) );
  ANDN U18961 ( .B(y[3006]), .A(x[3006]), .Z(n20825) );
  ANDN U18962 ( .B(n9984), .A(n20825), .Z(n9985) );
  NANDN U18963 ( .A(n12221), .B(n9985), .Z(n9986) );
  AND U18964 ( .A(n20821), .B(n9986), .Z(n9987) );
  NANDN U18965 ( .A(y[3007]), .B(x[3007]), .Z(n12220) );
  AND U18966 ( .A(n9987), .B(n12220), .Z(n9989) );
  NANDN U18967 ( .A(x[3008]), .B(y[3008]), .Z(n12218) );
  ANDN U18968 ( .B(y[3007]), .A(x[3007]), .Z(n20824) );
  ANDN U18969 ( .B(n12218), .A(n20824), .Z(n9988) );
  NANDN U18970 ( .A(n9989), .B(n9988), .Z(n9990) );
  AND U18971 ( .A(n12219), .B(n9990), .Z(n9991) );
  NANDN U18972 ( .A(y[3009]), .B(x[3009]), .Z(n12216) );
  NAND U18973 ( .A(n9991), .B(n12216), .Z(n9992) );
  NANDN U18974 ( .A(x[3009]), .B(y[3009]), .Z(n12217) );
  AND U18975 ( .A(n9992), .B(n12217), .Z(n9993) );
  NAND U18976 ( .A(n20831), .B(n9993), .Z(n9994) );
  NANDN U18977 ( .A(n12215), .B(n9994), .Z(n9995) );
  ANDN U18978 ( .B(x[3011]), .A(y[3011]), .Z(n20833) );
  OR U18979 ( .A(n9995), .B(n20833), .Z(n9996) );
  NAND U18980 ( .A(n9997), .B(n9996), .Z(n9999) );
  ANDN U18981 ( .B(x[3012]), .A(y[3012]), .Z(n9998) );
  ANDN U18982 ( .B(n9999), .A(n9998), .Z(n10000) );
  NANDN U18983 ( .A(y[3013]), .B(x[3013]), .Z(n28478) );
  AND U18984 ( .A(n10000), .B(n28478), .Z(n10001) );
  NANDN U18985 ( .A(x[3013]), .B(y[3013]), .Z(n20837) );
  NANDN U18986 ( .A(x[3014]), .B(y[3014]), .Z(n12213) );
  AND U18987 ( .A(n20837), .B(n12213), .Z(n24111) );
  NANDN U18988 ( .A(n10001), .B(n24111), .Z(n10002) );
  NAND U18989 ( .A(n10003), .B(n10002), .Z(n10004) );
  NANDN U18990 ( .A(x[3015]), .B(y[3015]), .Z(n28480) );
  AND U18991 ( .A(n10004), .B(n28480), .Z(n10005) );
  AND U18992 ( .A(n20844), .B(n10005), .Z(n10008) );
  NANDN U18993 ( .A(y[3017]), .B(x[3017]), .Z(n28483) );
  ANDN U18994 ( .B(x[3016]), .A(y[3016]), .Z(n10006) );
  ANDN U18995 ( .B(n28483), .A(n10006), .Z(n10007) );
  NANDN U18996 ( .A(n10008), .B(n10007), .Z(n10009) );
  NANDN U18997 ( .A(n20849), .B(n10009), .Z(n10010) );
  ANDN U18998 ( .B(y[3017]), .A(x[3017]), .Z(n12212) );
  OR U18999 ( .A(n10010), .B(n12212), .Z(n10011) );
  NAND U19000 ( .A(n28485), .B(n10011), .Z(n10012) );
  NANDN U19001 ( .A(n24110), .B(n10012), .Z(n10013) );
  NAND U19002 ( .A(n28487), .B(n10013), .Z(n10014) );
  NANDN U19003 ( .A(x[3022]), .B(y[3022]), .Z(n12209) );
  AND U19004 ( .A(n10014), .B(n12209), .Z(n10015) );
  NAND U19005 ( .A(n28488), .B(n10015), .Z(n10016) );
  NANDN U19006 ( .A(n28489), .B(n10016), .Z(n10017) );
  AND U19007 ( .A(n28490), .B(n10017), .Z(n10018) );
  NANDN U19008 ( .A(x[3023]), .B(y[3023]), .Z(n12208) );
  NAND U19009 ( .A(n10018), .B(n12208), .Z(n10019) );
  NANDN U19010 ( .A(n28493), .B(n10019), .Z(n10020) );
  AND U19011 ( .A(n28494), .B(n10020), .Z(n10021) );
  OR U19012 ( .A(n28495), .B(n10021), .Z(n10022) );
  NAND U19013 ( .A(n24109), .B(n10022), .Z(n10023) );
  NANDN U19014 ( .A(n28496), .B(n10023), .Z(n10024) );
  NANDN U19015 ( .A(x[3029]), .B(y[3029]), .Z(n12202) );
  NANDN U19016 ( .A(x[3030]), .B(y[3030]), .Z(n12199) );
  AND U19017 ( .A(n12202), .B(n12199), .Z(n28497) );
  AND U19018 ( .A(n10024), .B(n28497), .Z(n10025) );
  NANDN U19019 ( .A(y[3030]), .B(x[3030]), .Z(n12200) );
  NANDN U19020 ( .A(y[3031]), .B(x[3031]), .Z(n12197) );
  AND U19021 ( .A(n12200), .B(n12197), .Z(n28498) );
  NANDN U19022 ( .A(n10025), .B(n28498), .Z(n10026) );
  NANDN U19023 ( .A(n28499), .B(n10026), .Z(n10027) );
  AND U19024 ( .A(n28500), .B(n10027), .Z(n10028) );
  NANDN U19025 ( .A(y[3033]), .B(x[3033]), .Z(n20889) );
  AND U19026 ( .A(n10028), .B(n20889), .Z(n10029) );
  NANDN U19027 ( .A(x[3033]), .B(y[3033]), .Z(n12195) );
  NANDN U19028 ( .A(x[3034]), .B(y[3034]), .Z(n24106) );
  AND U19029 ( .A(n12195), .B(n24106), .Z(n28502) );
  NANDN U19030 ( .A(n10029), .B(n28502), .Z(n10030) );
  NAND U19031 ( .A(n10031), .B(n10030), .Z(n10032) );
  AND U19032 ( .A(n28503), .B(n10032), .Z(n10033) );
  NANDN U19033 ( .A(y[3037]), .B(x[3037]), .Z(n12192) );
  ANDN U19034 ( .B(x[3036]), .A(y[3036]), .Z(n20894) );
  ANDN U19035 ( .B(n12192), .A(n20894), .Z(n28504) );
  NANDN U19036 ( .A(n10033), .B(n28504), .Z(n10034) );
  NAND U19037 ( .A(n10035), .B(n10034), .Z(n10037) );
  NANDN U19038 ( .A(y[3039]), .B(x[3039]), .Z(n12189) );
  NANDN U19039 ( .A(y[3038]), .B(x[3038]), .Z(n10036) );
  AND U19040 ( .A(n12189), .B(n10036), .Z(n24105) );
  AND U19041 ( .A(n10037), .B(n24105), .Z(n10039) );
  NANDN U19042 ( .A(x[3039]), .B(y[3039]), .Z(n12191) );
  NANDN U19043 ( .A(x[3040]), .B(y[3040]), .Z(n10038) );
  NAND U19044 ( .A(n12191), .B(n10038), .Z(n28506) );
  OR U19045 ( .A(n10039), .B(n28506), .Z(n10040) );
  NAND U19046 ( .A(n28507), .B(n10040), .Z(n10041) );
  NAND U19047 ( .A(n28508), .B(n10041), .Z(n10042) );
  NANDN U19048 ( .A(n28509), .B(n10042), .Z(n10043) );
  NANDN U19049 ( .A(x[3044]), .B(y[3044]), .Z(n12188) );
  AND U19050 ( .A(n10043), .B(n12188), .Z(n10044) );
  NAND U19051 ( .A(n28510), .B(n10044), .Z(n10045) );
  NANDN U19052 ( .A(n28511), .B(n10045), .Z(n10046) );
  AND U19053 ( .A(n28513), .B(n10046), .Z(n10047) );
  NANDN U19054 ( .A(x[3045]), .B(y[3045]), .Z(n12187) );
  AND U19055 ( .A(n10047), .B(n12187), .Z(n10048) );
  ANDN U19056 ( .B(n28517), .A(n10048), .Z(n10049) );
  NANDN U19057 ( .A(x[3047]), .B(y[3047]), .Z(n20916) );
  NANDN U19058 ( .A(x[3048]), .B(y[3048]), .Z(n20923) );
  NAND U19059 ( .A(n20916), .B(n20923), .Z(n24103) );
  OR U19060 ( .A(n10049), .B(n24103), .Z(n10050) );
  NAND U19061 ( .A(n24102), .B(n10050), .Z(n10051) );
  NANDN U19062 ( .A(n28518), .B(n10051), .Z(n10052) );
  AND U19063 ( .A(n28519), .B(n10052), .Z(n10053) );
  NANDN U19064 ( .A(x[3051]), .B(y[3051]), .Z(n12183) );
  NANDN U19065 ( .A(x[3052]), .B(y[3052]), .Z(n20932) );
  NAND U19066 ( .A(n12183), .B(n20932), .Z(n28520) );
  OR U19067 ( .A(n10053), .B(n28520), .Z(n10054) );
  NAND U19068 ( .A(n28521), .B(n10054), .Z(n10055) );
  NANDN U19069 ( .A(x[3053]), .B(y[3053]), .Z(n20933) );
  NANDN U19070 ( .A(x[3054]), .B(y[3054]), .Z(n12180) );
  AND U19071 ( .A(n20933), .B(n12180), .Z(n24101) );
  AND U19072 ( .A(n10055), .B(n24101), .Z(n10057) );
  ANDN U19073 ( .B(x[3054]), .A(y[3054]), .Z(n20937) );
  IV U19074 ( .A(n20937), .Z(n28522) );
  ANDN U19075 ( .B(x[3055]), .A(y[3055]), .Z(n12178) );
  ANDN U19076 ( .B(n28522), .A(n12178), .Z(n10056) );
  NANDN U19077 ( .A(n10057), .B(n10056), .Z(n10058) );
  NANDN U19078 ( .A(n28523), .B(n10058), .Z(n10059) );
  ANDN U19079 ( .B(x[3057]), .A(y[3057]), .Z(n28524) );
  ANDN U19080 ( .B(n10059), .A(n28524), .Z(n10060) );
  NANDN U19081 ( .A(n12177), .B(n10060), .Z(n10061) );
  NAND U19082 ( .A(n28527), .B(n10061), .Z(n10062) );
  NANDN U19083 ( .A(n24100), .B(n10062), .Z(n10064) );
  NANDN U19084 ( .A(x[3060]), .B(y[3060]), .Z(n10063) );
  NANDN U19085 ( .A(x[3061]), .B(y[3061]), .Z(n10065) );
  AND U19086 ( .A(n10063), .B(n10065), .Z(n20956) );
  NANDN U19087 ( .A(x[3059]), .B(y[3059]), .Z(n12175) );
  AND U19088 ( .A(n20956), .B(n12175), .Z(n24099) );
  AND U19089 ( .A(n10064), .B(n24099), .Z(n10069) );
  ANDN U19090 ( .B(x[3060]), .A(y[3060]), .Z(n20952) );
  NANDN U19091 ( .A(y[3062]), .B(x[3062]), .Z(n10067) );
  NANDN U19092 ( .A(y[3061]), .B(x[3061]), .Z(n10066) );
  AND U19093 ( .A(n10067), .B(n10066), .Z(n10068) );
  NANDN U19094 ( .A(y[3063]), .B(x[3063]), .Z(n10073) );
  NAND U19095 ( .A(n10068), .B(n10073), .Z(n20958) );
  NANDN U19096 ( .A(n10069), .B(n28530), .Z(n10076) );
  XNOR U19097 ( .A(y[3063]), .B(x[3063]), .Z(n10071) );
  NANDN U19098 ( .A(x[3062]), .B(y[3062]), .Z(n10070) );
  NAND U19099 ( .A(n10071), .B(n10070), .Z(n10072) );
  NAND U19100 ( .A(n10073), .B(n10072), .Z(n10075) );
  NANDN U19101 ( .A(x[3064]), .B(y[3064]), .Z(n10074) );
  AND U19102 ( .A(n10075), .B(n10074), .Z(n24098) );
  AND U19103 ( .A(n10076), .B(n24098), .Z(n10079) );
  NANDN U19104 ( .A(y[3064]), .B(x[3064]), .Z(n10078) );
  NANDN U19105 ( .A(y[3065]), .B(x[3065]), .Z(n10077) );
  NAND U19106 ( .A(n10078), .B(n10077), .Z(n28531) );
  OR U19107 ( .A(n10079), .B(n28531), .Z(n10080) );
  NAND U19108 ( .A(n10081), .B(n10080), .Z(n10082) );
  NAND U19109 ( .A(n28533), .B(n10082), .Z(n10083) );
  AND U19110 ( .A(n12174), .B(n10083), .Z(n10084) );
  AND U19111 ( .A(n28534), .B(n10084), .Z(n10085) );
  OR U19112 ( .A(n28535), .B(n10085), .Z(n10086) );
  NAND U19113 ( .A(n28536), .B(n10086), .Z(n10087) );
  NANDN U19114 ( .A(n28537), .B(n10087), .Z(n10088) );
  AND U19115 ( .A(n28538), .B(n10088), .Z(n10089) );
  NANDN U19116 ( .A(y[3072]), .B(x[3072]), .Z(n20975) );
  NANDN U19117 ( .A(y[3073]), .B(x[3073]), .Z(n12169) );
  NAND U19118 ( .A(n20975), .B(n12169), .Z(n28539) );
  OR U19119 ( .A(n10089), .B(n28539), .Z(n10090) );
  AND U19120 ( .A(n28540), .B(n10090), .Z(n10091) );
  OR U19121 ( .A(n28541), .B(n10091), .Z(n10092) );
  NAND U19122 ( .A(n28542), .B(n10092), .Z(n10093) );
  NANDN U19123 ( .A(n12164), .B(n10093), .Z(n10094) );
  NANDN U19124 ( .A(y[3076]), .B(x[3076]), .Z(n24095) );
  NANDN U19125 ( .A(n10094), .B(n24095), .Z(n10095) );
  ANDN U19126 ( .B(y[3077]), .A(x[3077]), .Z(n28544) );
  ANDN U19127 ( .B(n10095), .A(n28544), .Z(n10096) );
  AND U19128 ( .A(n12165), .B(n10096), .Z(n10097) );
  ANDN U19129 ( .B(n10098), .A(n10097), .Z(n10099) );
  ANDN U19130 ( .B(y[3080]), .A(x[3080]), .Z(n20998) );
  NANDN U19131 ( .A(x[3079]), .B(y[3079]), .Z(n12163) );
  NANDN U19132 ( .A(n20998), .B(n12163), .Z(n28548) );
  OR U19133 ( .A(n10099), .B(n28548), .Z(n10100) );
  NAND U19134 ( .A(n28549), .B(n10100), .Z(n10101) );
  NANDN U19135 ( .A(n10102), .B(n10101), .Z(n10103) );
  AND U19136 ( .A(n28551), .B(n10103), .Z(n10106) );
  NANDN U19137 ( .A(x[3084]), .B(y[3084]), .Z(n10105) );
  NANDN U19138 ( .A(x[3083]), .B(y[3083]), .Z(n10104) );
  AND U19139 ( .A(n10105), .B(n10104), .Z(n21005) );
  NANDN U19140 ( .A(n10106), .B(n21005), .Z(n10107) );
  NAND U19141 ( .A(n28553), .B(n10107), .Z(n10110) );
  NANDN U19142 ( .A(x[3086]), .B(y[3086]), .Z(n10109) );
  NANDN U19143 ( .A(x[3085]), .B(y[3085]), .Z(n10108) );
  NAND U19144 ( .A(n10109), .B(n10108), .Z(n28554) );
  ANDN U19145 ( .B(n10110), .A(n28554), .Z(n10111) );
  OR U19146 ( .A(n28555), .B(n10111), .Z(n10112) );
  NAND U19147 ( .A(n28556), .B(n10112), .Z(n10113) );
  NANDN U19148 ( .A(n28557), .B(n10113), .Z(n10114) );
  AND U19149 ( .A(n28558), .B(n10114), .Z(n10115) );
  ANDN U19150 ( .B(x[3090]), .A(y[3090]), .Z(n21019) );
  ANDN U19151 ( .B(x[3091]), .A(y[3091]), .Z(n12158) );
  NOR U19152 ( .A(n21019), .B(n12158), .Z(n28559) );
  NANDN U19153 ( .A(n10115), .B(n28559), .Z(n10116) );
  NANDN U19154 ( .A(n12161), .B(n10116), .Z(n10117) );
  AND U19155 ( .A(n28562), .B(n10117), .Z(n10118) );
  NANDN U19156 ( .A(x[3093]), .B(y[3093]), .Z(n21026) );
  NANDN U19157 ( .A(x[3094]), .B(y[3094]), .Z(n21032) );
  NAND U19158 ( .A(n21026), .B(n21032), .Z(n28563) );
  OR U19159 ( .A(n10118), .B(n28563), .Z(n10119) );
  NAND U19160 ( .A(n28564), .B(n10119), .Z(n10120) );
  NANDN U19161 ( .A(n28565), .B(n10120), .Z(n10121) );
  AND U19162 ( .A(n28566), .B(n10121), .Z(n10122) );
  NANDN U19163 ( .A(x[3097]), .B(y[3097]), .Z(n12155) );
  NANDN U19164 ( .A(x[3098]), .B(y[3098]), .Z(n21048) );
  AND U19165 ( .A(n12155), .B(n21048), .Z(n28567) );
  NANDN U19166 ( .A(n10122), .B(n28567), .Z(n10123) );
  AND U19167 ( .A(n28568), .B(n10123), .Z(n10124) );
  OR U19168 ( .A(n28569), .B(n10124), .Z(n10125) );
  NAND U19169 ( .A(n28570), .B(n10125), .Z(n10126) );
  NANDN U19170 ( .A(n28571), .B(n10126), .Z(n10127) );
  AND U19171 ( .A(n28572), .B(n10127), .Z(n10128) );
  NANDN U19172 ( .A(x[3103]), .B(y[3103]), .Z(n12153) );
  NANDN U19173 ( .A(x[3104]), .B(y[3104]), .Z(n21070) );
  NAND U19174 ( .A(n12153), .B(n21070), .Z(n28573) );
  OR U19175 ( .A(n10128), .B(n28573), .Z(n10129) );
  AND U19176 ( .A(n28574), .B(n10129), .Z(n10130) );
  NANDN U19177 ( .A(x[3105]), .B(y[3105]), .Z(n21069) );
  NANDN U19178 ( .A(x[3106]), .B(y[3106]), .Z(n21076) );
  NAND U19179 ( .A(n21069), .B(n21076), .Z(n24094) );
  OR U19180 ( .A(n10130), .B(n24094), .Z(n10131) );
  NAND U19181 ( .A(n28576), .B(n10131), .Z(n10132) );
  NANDN U19182 ( .A(n28577), .B(n10132), .Z(n10133) );
  AND U19183 ( .A(n28578), .B(n10133), .Z(n10134) );
  NANDN U19184 ( .A(x[3109]), .B(y[3109]), .Z(n12151) );
  NANDN U19185 ( .A(x[3110]), .B(y[3110]), .Z(n21092) );
  AND U19186 ( .A(n12151), .B(n21092), .Z(n28579) );
  NANDN U19187 ( .A(n10134), .B(n28579), .Z(n10135) );
  NANDN U19188 ( .A(n24093), .B(n10135), .Z(n10136) );
  NANDN U19189 ( .A(x[3111]), .B(y[3111]), .Z(n21091) );
  NANDN U19190 ( .A(x[3112]), .B(y[3112]), .Z(n21098) );
  AND U19191 ( .A(n21091), .B(n21098), .Z(n24092) );
  AND U19192 ( .A(n10136), .B(n24092), .Z(n10137) );
  OR U19193 ( .A(n28580), .B(n10137), .Z(n10138) );
  NAND U19194 ( .A(n28581), .B(n10138), .Z(n10139) );
  NANDN U19195 ( .A(n28582), .B(n10139), .Z(n10140) );
  AND U19196 ( .A(n28583), .B(n10140), .Z(n10141) );
  ANDN U19197 ( .B(x[3116]), .A(y[3116]), .Z(n21109) );
  ANDN U19198 ( .B(x[3117]), .A(y[3117]), .Z(n21119) );
  OR U19199 ( .A(n21109), .B(n21119), .Z(n28584) );
  OR U19200 ( .A(n10141), .B(n28584), .Z(n10142) );
  NANDN U19201 ( .A(x[3117]), .B(y[3117]), .Z(n21113) );
  NANDN U19202 ( .A(x[3118]), .B(y[3118]), .Z(n21120) );
  AND U19203 ( .A(n21113), .B(n21120), .Z(n24091) );
  AND U19204 ( .A(n10142), .B(n24091), .Z(n10143) );
  ANDN U19205 ( .B(x[3118]), .A(y[3118]), .Z(n21116) );
  ANDN U19206 ( .B(x[3119]), .A(y[3119]), .Z(n21126) );
  OR U19207 ( .A(n21116), .B(n21126), .Z(n28585) );
  OR U19208 ( .A(n10143), .B(n28585), .Z(n10144) );
  NAND U19209 ( .A(n28586), .B(n10144), .Z(n10145) );
  NANDN U19210 ( .A(n24090), .B(n10145), .Z(n10146) );
  NANDN U19211 ( .A(x[3121]), .B(y[3121]), .Z(n12147) );
  NANDN U19212 ( .A(x[3122]), .B(y[3122]), .Z(n21136) );
  AND U19213 ( .A(n12147), .B(n21136), .Z(n24089) );
  AND U19214 ( .A(n10146), .B(n24089), .Z(n10147) );
  ANDN U19215 ( .B(x[3122]), .A(y[3122]), .Z(n21131) );
  ANDN U19216 ( .B(x[3123]), .A(y[3123]), .Z(n21141) );
  NOR U19217 ( .A(n21131), .B(n21141), .Z(n28588) );
  NANDN U19218 ( .A(n10147), .B(n28588), .Z(n10148) );
  NANDN U19219 ( .A(n28589), .B(n10148), .Z(n10149) );
  AND U19220 ( .A(n28590), .B(n10149), .Z(n10150) );
  NANDN U19221 ( .A(x[3125]), .B(y[3125]), .Z(n21143) );
  NANDN U19222 ( .A(x[3126]), .B(y[3126]), .Z(n12146) );
  NAND U19223 ( .A(n21143), .B(n12146), .Z(n24088) );
  OR U19224 ( .A(n10150), .B(n24088), .Z(n10151) );
  NAND U19225 ( .A(n28591), .B(n10151), .Z(n10152) );
  NANDN U19226 ( .A(n28592), .B(n10152), .Z(n10153) );
  AND U19227 ( .A(n28593), .B(n10153), .Z(n10154) );
  NANDN U19228 ( .A(x[3129]), .B(y[3129]), .Z(n21157) );
  NANDN U19229 ( .A(x[3130]), .B(y[3130]), .Z(n21164) );
  AND U19230 ( .A(n21157), .B(n21164), .Z(n28594) );
  NANDN U19231 ( .A(n10154), .B(n28594), .Z(n10155) );
  AND U19232 ( .A(n28595), .B(n10155), .Z(n10156) );
  OR U19233 ( .A(n28596), .B(n10156), .Z(n10157) );
  NAND U19234 ( .A(n28597), .B(n10157), .Z(n10158) );
  NANDN U19235 ( .A(n28598), .B(n10158), .Z(n10159) );
  AND U19236 ( .A(n28599), .B(n10159), .Z(n10160) );
  NANDN U19237 ( .A(x[3135]), .B(y[3135]), .Z(n21179) );
  NANDN U19238 ( .A(x[3136]), .B(y[3136]), .Z(n21186) );
  NAND U19239 ( .A(n21179), .B(n21186), .Z(n24087) );
  OR U19240 ( .A(n10160), .B(n24087), .Z(n10161) );
  AND U19241 ( .A(n28601), .B(n10161), .Z(n10162) );
  OR U19242 ( .A(n28602), .B(n10162), .Z(n10163) );
  NAND U19243 ( .A(n28603), .B(n10163), .Z(n10164) );
  NANDN U19244 ( .A(n28604), .B(n10164), .Z(n10165) );
  AND U19245 ( .A(n28605), .B(n10165), .Z(n10166) );
  OR U19246 ( .A(n28606), .B(n10166), .Z(n10167) );
  NAND U19247 ( .A(n28607), .B(n10167), .Z(n10168) );
  NAND U19248 ( .A(n28608), .B(n10168), .Z(n10171) );
  NANDN U19249 ( .A(y[3145]), .B(x[3145]), .Z(n10170) );
  NANDN U19250 ( .A(y[3144]), .B(x[3144]), .Z(n10169) );
  NAND U19251 ( .A(n10170), .B(n10169), .Z(n28609) );
  ANDN U19252 ( .B(n10171), .A(n28609), .Z(n10174) );
  NANDN U19253 ( .A(x[3146]), .B(y[3146]), .Z(n10173) );
  NANDN U19254 ( .A(x[3145]), .B(y[3145]), .Z(n10172) );
  AND U19255 ( .A(n10173), .B(n10172), .Z(n28610) );
  NANDN U19256 ( .A(n10174), .B(n28610), .Z(n10175) );
  NANDN U19257 ( .A(n24086), .B(n10175), .Z(n10176) );
  AND U19258 ( .A(n28611), .B(n10176), .Z(n10177) );
  ANDN U19259 ( .B(x[3149]), .A(y[3149]), .Z(n21225) );
  NANDN U19260 ( .A(y[3148]), .B(x[3148]), .Z(n21218) );
  NANDN U19261 ( .A(n21225), .B(n21218), .Z(n28612) );
  OR U19262 ( .A(n10177), .B(n28612), .Z(n10178) );
  NANDN U19263 ( .A(n28613), .B(n10178), .Z(n10179) );
  NANDN U19264 ( .A(n28615), .B(n10179), .Z(n10180) );
  AND U19265 ( .A(n28616), .B(n10180), .Z(n10181) );
  ANDN U19266 ( .B(x[3152]), .A(y[3152]), .Z(n12138) );
  ANDN U19267 ( .B(x[3153]), .A(y[3153]), .Z(n21240) );
  NOR U19268 ( .A(n12138), .B(n21240), .Z(n28617) );
  NANDN U19269 ( .A(n10181), .B(n28617), .Z(n10182) );
  NANDN U19270 ( .A(n24085), .B(n10182), .Z(n10183) );
  AND U19271 ( .A(n28618), .B(n10183), .Z(n10184) );
  OR U19272 ( .A(n28619), .B(n10184), .Z(n10185) );
  NAND U19273 ( .A(n28620), .B(n10185), .Z(n10186) );
  NANDN U19274 ( .A(n28621), .B(n10186), .Z(n10187) );
  AND U19275 ( .A(n28622), .B(n10187), .Z(n10188) );
  NANDN U19276 ( .A(x[3159]), .B(y[3159]), .Z(n21257) );
  NANDN U19277 ( .A(x[3160]), .B(y[3160]), .Z(n12135) );
  NAND U19278 ( .A(n21257), .B(n12135), .Z(n28623) );
  OR U19279 ( .A(n10188), .B(n28623), .Z(n10189) );
  AND U19280 ( .A(n28624), .B(n10189), .Z(n10190) );
  ANDN U19281 ( .B(y[3162]), .A(x[3162]), .Z(n21273) );
  NANDN U19282 ( .A(x[3161]), .B(y[3161]), .Z(n12134) );
  NANDN U19283 ( .A(n21273), .B(n12134), .Z(n28625) );
  OR U19284 ( .A(n10190), .B(n28625), .Z(n10191) );
  NAND U19285 ( .A(n28626), .B(n10191), .Z(n10192) );
  NANDN U19286 ( .A(n24084), .B(n10192), .Z(n10193) );
  NANDN U19287 ( .A(y[3164]), .B(x[3164]), .Z(n12133) );
  NANDN U19288 ( .A(y[3165]), .B(x[3165]), .Z(n21282) );
  AND U19289 ( .A(n12133), .B(n21282), .Z(n24083) );
  AND U19290 ( .A(n10193), .B(n24083), .Z(n10194) );
  NANDN U19291 ( .A(x[3166]), .B(y[3166]), .Z(n21285) );
  ANDN U19292 ( .B(y[3165]), .A(x[3165]), .Z(n21279) );
  ANDN U19293 ( .B(n21285), .A(n21279), .Z(n28627) );
  NANDN U19294 ( .A(n10194), .B(n28627), .Z(n10195) );
  NANDN U19295 ( .A(n28628), .B(n10195), .Z(n10196) );
  NANDN U19296 ( .A(x[3167]), .B(y[3167]), .Z(n21284) );
  NANDN U19297 ( .A(x[3168]), .B(y[3168]), .Z(n21292) );
  AND U19298 ( .A(n21284), .B(n21292), .Z(n28631) );
  AND U19299 ( .A(n10196), .B(n28631), .Z(n10197) );
  NANDN U19300 ( .A(y[3168]), .B(x[3168]), .Z(n12130) );
  NANDN U19301 ( .A(y[3169]), .B(x[3169]), .Z(n12129) );
  NAND U19302 ( .A(n12130), .B(n12129), .Z(n24082) );
  OR U19303 ( .A(n10197), .B(n24082), .Z(n10198) );
  NAND U19304 ( .A(n24081), .B(n10198), .Z(n10199) );
  NANDN U19305 ( .A(n28632), .B(n10199), .Z(n10200) );
  AND U19306 ( .A(n28633), .B(n10200), .Z(n10201) );
  NANDN U19307 ( .A(y[3172]), .B(x[3172]), .Z(n12126) );
  NANDN U19308 ( .A(y[3173]), .B(x[3173]), .Z(n21307) );
  NAND U19309 ( .A(n12126), .B(n21307), .Z(n28634) );
  OR U19310 ( .A(n10201), .B(n28634), .Z(n10202) );
  AND U19311 ( .A(n28635), .B(n10202), .Z(n10203) );
  OR U19312 ( .A(n28636), .B(n10203), .Z(n10204) );
  NAND U19313 ( .A(n24080), .B(n10204), .Z(n10205) );
  NANDN U19314 ( .A(n28637), .B(n10205), .Z(n10206) );
  NANDN U19315 ( .A(x[3177]), .B(y[3177]), .Z(n12122) );
  NANDN U19316 ( .A(x[3178]), .B(y[3178]), .Z(n12121) );
  AND U19317 ( .A(n12122), .B(n12121), .Z(n28638) );
  AND U19318 ( .A(n10206), .B(n28638), .Z(n10207) );
  NANDN U19319 ( .A(y[3178]), .B(x[3178]), .Z(n21318) );
  NANDN U19320 ( .A(y[3179]), .B(x[3179]), .Z(n21325) );
  AND U19321 ( .A(n21318), .B(n21325), .Z(n28639) );
  NANDN U19322 ( .A(n10207), .B(n28639), .Z(n10208) );
  NANDN U19323 ( .A(n28640), .B(n10208), .Z(n10209) );
  NANDN U19324 ( .A(y[3180]), .B(x[3180]), .Z(n21324) );
  NANDN U19325 ( .A(y[3181]), .B(x[3181]), .Z(n21331) );
  AND U19326 ( .A(n21324), .B(n21331), .Z(n24079) );
  AND U19327 ( .A(n10209), .B(n24079), .Z(n10210) );
  NANDN U19328 ( .A(x[3181]), .B(y[3181]), .Z(n12118) );
  NANDN U19329 ( .A(x[3182]), .B(y[3182]), .Z(n12117) );
  NAND U19330 ( .A(n12118), .B(n12117), .Z(n28643) );
  OR U19331 ( .A(n10210), .B(n28643), .Z(n10211) );
  NAND U19332 ( .A(n28644), .B(n10211), .Z(n10212) );
  NANDN U19333 ( .A(n24078), .B(n10212), .Z(n10213) );
  NANDN U19334 ( .A(y[3184]), .B(x[3184]), .Z(n21336) );
  NANDN U19335 ( .A(y[3185]), .B(x[3185]), .Z(n21343) );
  AND U19336 ( .A(n21336), .B(n21343), .Z(n24077) );
  AND U19337 ( .A(n10213), .B(n24077), .Z(n10214) );
  NANDN U19338 ( .A(x[3185]), .B(y[3185]), .Z(n12114) );
  NANDN U19339 ( .A(x[3186]), .B(y[3186]), .Z(n12113) );
  NAND U19340 ( .A(n12114), .B(n12113), .Z(n28645) );
  OR U19341 ( .A(n10214), .B(n28645), .Z(n10215) );
  AND U19342 ( .A(n28646), .B(n10215), .Z(n10216) );
  OR U19343 ( .A(n28647), .B(n10216), .Z(n10217) );
  NAND U19344 ( .A(n28648), .B(n10217), .Z(n10218) );
  NANDN U19345 ( .A(n28649), .B(n10218), .Z(n10219) );
  NANDN U19346 ( .A(y[3190]), .B(x[3190]), .Z(n21354) );
  NANDN U19347 ( .A(y[3191]), .B(x[3191]), .Z(n21361) );
  AND U19348 ( .A(n21354), .B(n21361), .Z(n24076) );
  AND U19349 ( .A(n10219), .B(n24076), .Z(n10220) );
  NANDN U19350 ( .A(x[3191]), .B(y[3191]), .Z(n12108) );
  NANDN U19351 ( .A(x[3192]), .B(y[3192]), .Z(n12107) );
  AND U19352 ( .A(n12108), .B(n12107), .Z(n28650) );
  NANDN U19353 ( .A(n10220), .B(n28650), .Z(n10221) );
  NANDN U19354 ( .A(n28651), .B(n10221), .Z(n10222) );
  AND U19355 ( .A(n28652), .B(n10222), .Z(n10223) );
  OR U19356 ( .A(n28653), .B(n10223), .Z(n10224) );
  NAND U19357 ( .A(n24075), .B(n10224), .Z(n10225) );
  NANDN U19358 ( .A(n28655), .B(n10225), .Z(n10226) );
  NANDN U19359 ( .A(x[3197]), .B(y[3197]), .Z(n12102) );
  NANDN U19360 ( .A(x[3198]), .B(y[3198]), .Z(n12101) );
  AND U19361 ( .A(n12102), .B(n12101), .Z(n28656) );
  AND U19362 ( .A(n10226), .B(n28656), .Z(n10227) );
  NANDN U19363 ( .A(y[3198]), .B(x[3198]), .Z(n21381) );
  NANDN U19364 ( .A(y[3199]), .B(x[3199]), .Z(n12099) );
  NAND U19365 ( .A(n21381), .B(n12099), .Z(n24074) );
  OR U19366 ( .A(n10227), .B(n24074), .Z(n10228) );
  NANDN U19367 ( .A(x[3199]), .B(y[3199]), .Z(n12100) );
  NANDN U19368 ( .A(x[3200]), .B(y[3200]), .Z(n12097) );
  AND U19369 ( .A(n12100), .B(n12097), .Z(n24073) );
  AND U19370 ( .A(n10228), .B(n24073), .Z(n10229) );
  OR U19371 ( .A(n28657), .B(n10229), .Z(n10230) );
  NAND U19372 ( .A(n28658), .B(n10230), .Z(n10231) );
  NANDN U19373 ( .A(n28659), .B(n10231), .Z(n10232) );
  AND U19374 ( .A(n28660), .B(n10232), .Z(n10233) );
  NANDN U19375 ( .A(y[3204]), .B(x[3204]), .Z(n21395) );
  ANDN U19376 ( .B(x[3205]), .A(y[3205]), .Z(n21403) );
  ANDN U19377 ( .B(n21395), .A(n21403), .Z(n28661) );
  NANDN U19378 ( .A(n10233), .B(n28661), .Z(n10234) );
  NANDN U19379 ( .A(n28662), .B(n10234), .Z(n10235) );
  AND U19380 ( .A(n28663), .B(n10235), .Z(n10236) );
  OR U19381 ( .A(n28664), .B(n10236), .Z(n10237) );
  NAND U19382 ( .A(n28665), .B(n10237), .Z(n10238) );
  NANDN U19383 ( .A(n28666), .B(n10238), .Z(n10239) );
  NANDN U19384 ( .A(y[3210]), .B(x[3210]), .Z(n21412) );
  NANDN U19385 ( .A(y[3211]), .B(x[3211]), .Z(n12087) );
  AND U19386 ( .A(n21412), .B(n12087), .Z(n24072) );
  AND U19387 ( .A(n10239), .B(n24072), .Z(n10240) );
  NANDN U19388 ( .A(x[3211]), .B(y[3211]), .Z(n21416) );
  NANDN U19389 ( .A(x[3212]), .B(y[3212]), .Z(n21423) );
  NAND U19390 ( .A(n21416), .B(n21423), .Z(n28669) );
  OR U19391 ( .A(n10240), .B(n28669), .Z(n10241) );
  NANDN U19392 ( .A(y[3212]), .B(x[3212]), .Z(n12086) );
  NANDN U19393 ( .A(y[3213]), .B(x[3213]), .Z(n12085) );
  AND U19394 ( .A(n12086), .B(n12085), .Z(n28670) );
  AND U19395 ( .A(n10241), .B(n28670), .Z(n10242) );
  ANDN U19396 ( .B(y[3214]), .A(x[3214]), .Z(n21429) );
  NANDN U19397 ( .A(x[3213]), .B(y[3213]), .Z(n21422) );
  NANDN U19398 ( .A(n21429), .B(n21422), .Z(n24071) );
  OR U19399 ( .A(n10242), .B(n24071), .Z(n10243) );
  NAND U19400 ( .A(n24070), .B(n10243), .Z(n10244) );
  NANDN U19401 ( .A(n28671), .B(n10244), .Z(n10245) );
  AND U19402 ( .A(n28672), .B(n10245), .Z(n10246) );
  NANDN U19403 ( .A(x[3217]), .B(y[3217]), .Z(n12080) );
  NANDN U19404 ( .A(x[3218]), .B(y[3218]), .Z(n21440) );
  AND U19405 ( .A(n12080), .B(n21440), .Z(n28673) );
  NANDN U19406 ( .A(n10246), .B(n28673), .Z(n10247) );
  NANDN U19407 ( .A(n24069), .B(n10247), .Z(n10248) );
  NANDN U19408 ( .A(x[3219]), .B(y[3219]), .Z(n21439) );
  NANDN U19409 ( .A(x[3220]), .B(y[3220]), .Z(n21446) );
  AND U19410 ( .A(n21439), .B(n21446), .Z(n24068) );
  AND U19411 ( .A(n10248), .B(n24068), .Z(n10249) );
  OR U19412 ( .A(n28674), .B(n10249), .Z(n10250) );
  NAND U19413 ( .A(n28675), .B(n10250), .Z(n10251) );
  NANDN U19414 ( .A(n28676), .B(n10251), .Z(n10252) );
  AND U19415 ( .A(n28678), .B(n10252), .Z(n10253) );
  NANDN U19416 ( .A(y[3224]), .B(x[3224]), .Z(n21454) );
  NANDN U19417 ( .A(y[3225]), .B(x[3225]), .Z(n21461) );
  NAND U19418 ( .A(n21454), .B(n21461), .Z(n28679) );
  OR U19419 ( .A(n10253), .B(n28679), .Z(n10254) );
  NANDN U19420 ( .A(x[3225]), .B(y[3225]), .Z(n12072) );
  NANDN U19421 ( .A(x[3226]), .B(y[3226]), .Z(n12071) );
  AND U19422 ( .A(n12072), .B(n12071), .Z(n24067) );
  AND U19423 ( .A(n10254), .B(n24067), .Z(n10255) );
  NANDN U19424 ( .A(y[3226]), .B(x[3226]), .Z(n21460) );
  NANDN U19425 ( .A(y[3227]), .B(x[3227]), .Z(n21467) );
  NAND U19426 ( .A(n21460), .B(n21467), .Z(n28680) );
  OR U19427 ( .A(n10255), .B(n28680), .Z(n10256) );
  NAND U19428 ( .A(n28681), .B(n10256), .Z(n10257) );
  NANDN U19429 ( .A(n24066), .B(n10257), .Z(n10258) );
  NANDN U19430 ( .A(x[3229]), .B(y[3229]), .Z(n12068) );
  NANDN U19431 ( .A(x[3230]), .B(y[3230]), .Z(n12067) );
  AND U19432 ( .A(n12068), .B(n12067), .Z(n24065) );
  AND U19433 ( .A(n10258), .B(n24065), .Z(n10259) );
  NANDN U19434 ( .A(y[3230]), .B(x[3230]), .Z(n21472) );
  NANDN U19435 ( .A(y[3231]), .B(x[3231]), .Z(n21479) );
  AND U19436 ( .A(n21472), .B(n21479), .Z(n24064) );
  NANDN U19437 ( .A(n10259), .B(n24064), .Z(n10260) );
  NANDN U19438 ( .A(n28682), .B(n10260), .Z(n10261) );
  NANDN U19439 ( .A(y[3232]), .B(x[3232]), .Z(n21478) );
  NANDN U19440 ( .A(y[3233]), .B(x[3233]), .Z(n21485) );
  AND U19441 ( .A(n21478), .B(n21485), .Z(n28683) );
  AND U19442 ( .A(n10261), .B(n28683), .Z(n10262) );
  NANDN U19443 ( .A(x[3233]), .B(y[3233]), .Z(n12064) );
  NANDN U19444 ( .A(x[3234]), .B(y[3234]), .Z(n12063) );
  NAND U19445 ( .A(n12064), .B(n12063), .Z(n24063) );
  OR U19446 ( .A(n10262), .B(n24063), .Z(n10263) );
  NAND U19447 ( .A(n24062), .B(n10263), .Z(n10264) );
  NANDN U19448 ( .A(n28686), .B(n10264), .Z(n10265) );
  AND U19449 ( .A(n28687), .B(n10265), .Z(n10266) );
  NANDN U19450 ( .A(x[3237]), .B(y[3237]), .Z(n12060) );
  NANDN U19451 ( .A(x[3238]), .B(y[3238]), .Z(n12059) );
  NAND U19452 ( .A(n12060), .B(n12059), .Z(n28688) );
  OR U19453 ( .A(n10266), .B(n28688), .Z(n10267) );
  AND U19454 ( .A(n28689), .B(n10267), .Z(n10268) );
  OR U19455 ( .A(n28690), .B(n10268), .Z(n10269) );
  NAND U19456 ( .A(n24061), .B(n10269), .Z(n10270) );
  NANDN U19457 ( .A(n28691), .B(n10270), .Z(n10271) );
  NANDN U19458 ( .A(y[3242]), .B(x[3242]), .Z(n21508) );
  NANDN U19459 ( .A(y[3243]), .B(x[3243]), .Z(n21515) );
  AND U19460 ( .A(n21508), .B(n21515), .Z(n28692) );
  AND U19461 ( .A(n10271), .B(n28692), .Z(n10272) );
  NANDN U19462 ( .A(x[3243]), .B(y[3243]), .Z(n12054) );
  NANDN U19463 ( .A(x[3244]), .B(y[3244]), .Z(n12053) );
  AND U19464 ( .A(n12054), .B(n12053), .Z(n28693) );
  NANDN U19465 ( .A(n10272), .B(n28693), .Z(n10273) );
  NANDN U19466 ( .A(n28694), .B(n10273), .Z(n10274) );
  NANDN U19467 ( .A(x[3245]), .B(y[3245]), .Z(n12052) );
  NANDN U19468 ( .A(x[3246]), .B(y[3246]), .Z(n12051) );
  AND U19469 ( .A(n12052), .B(n12051), .Z(n24060) );
  AND U19470 ( .A(n10274), .B(n24060), .Z(n10275) );
  ANDN U19471 ( .B(x[3247]), .A(y[3247]), .Z(n21527) );
  NANDN U19472 ( .A(y[3246]), .B(x[3246]), .Z(n21520) );
  NANDN U19473 ( .A(n21527), .B(n21520), .Z(n28695) );
  OR U19474 ( .A(n10275), .B(n28695), .Z(n10276) );
  NAND U19475 ( .A(n28696), .B(n10276), .Z(n10277) );
  NANDN U19476 ( .A(n24059), .B(n10277), .Z(n10278) );
  NANDN U19477 ( .A(x[3249]), .B(y[3249]), .Z(n21530) );
  NANDN U19478 ( .A(x[3250]), .B(y[3250]), .Z(n12049) );
  AND U19479 ( .A(n21530), .B(n12049), .Z(n24058) );
  AND U19480 ( .A(n10278), .B(n24058), .Z(n10279) );
  NANDN U19481 ( .A(y[3250]), .B(x[3250]), .Z(n21534) );
  NANDN U19482 ( .A(y[3251]), .B(x[3251]), .Z(n21541) );
  NAND U19483 ( .A(n21534), .B(n21541), .Z(n28698) );
  OR U19484 ( .A(n10279), .B(n28698), .Z(n10280) );
  AND U19485 ( .A(n28699), .B(n10280), .Z(n10281) );
  OR U19486 ( .A(n28700), .B(n10281), .Z(n10282) );
  NAND U19487 ( .A(n28701), .B(n10282), .Z(n10283) );
  NANDN U19488 ( .A(n28702), .B(n10283), .Z(n10284) );
  AND U19489 ( .A(n21553), .B(n10284), .Z(n10285) );
  NANDN U19490 ( .A(x[3255]), .B(y[3255]), .Z(n28703) );
  AND U19491 ( .A(n10285), .B(n28703), .Z(n10287) );
  NANDN U19492 ( .A(y[3256]), .B(x[3256]), .Z(n10286) );
  NANDN U19493 ( .A(y[3257]), .B(x[3257]), .Z(n21559) );
  NAND U19494 ( .A(n10286), .B(n21559), .Z(n28705) );
  OR U19495 ( .A(n10287), .B(n28705), .Z(n10288) );
  NANDN U19496 ( .A(x[3257]), .B(y[3257]), .Z(n12044) );
  NANDN U19497 ( .A(x[3258]), .B(y[3258]), .Z(n12043) );
  AND U19498 ( .A(n12044), .B(n12043), .Z(n28706) );
  AND U19499 ( .A(n10288), .B(n28706), .Z(n10289) );
  NANDN U19500 ( .A(y[3258]), .B(x[3258]), .Z(n21558) );
  NANDN U19501 ( .A(y[3259]), .B(x[3259]), .Z(n21565) );
  NAND U19502 ( .A(n21558), .B(n21565), .Z(n24057) );
  OR U19503 ( .A(n10289), .B(n24057), .Z(n10290) );
  NAND U19504 ( .A(n24056), .B(n10290), .Z(n10291) );
  NANDN U19505 ( .A(n28707), .B(n10291), .Z(n10292) );
  AND U19506 ( .A(n28709), .B(n10292), .Z(n10293) );
  NANDN U19507 ( .A(y[3262]), .B(x[3262]), .Z(n21570) );
  NANDN U19508 ( .A(y[3263]), .B(x[3263]), .Z(n21577) );
  NAND U19509 ( .A(n21570), .B(n21577), .Z(n28710) );
  OR U19510 ( .A(n10293), .B(n28710), .Z(n10294) );
  AND U19511 ( .A(n28711), .B(n10294), .Z(n10295) );
  OR U19512 ( .A(n28712), .B(n10295), .Z(n10296) );
  NAND U19513 ( .A(n24055), .B(n10296), .Z(n10297) );
  NANDN U19514 ( .A(n28713), .B(n10297), .Z(n10298) );
  NANDN U19515 ( .A(x[3267]), .B(y[3267]), .Z(n12034) );
  NANDN U19516 ( .A(x[3268]), .B(y[3268]), .Z(n12033) );
  AND U19517 ( .A(n12034), .B(n12033), .Z(n28714) );
  AND U19518 ( .A(n10298), .B(n28714), .Z(n10299) );
  NANDN U19519 ( .A(y[3268]), .B(x[3268]), .Z(n21588) );
  NANDN U19520 ( .A(y[3269]), .B(x[3269]), .Z(n21595) );
  AND U19521 ( .A(n21588), .B(n21595), .Z(n28715) );
  NANDN U19522 ( .A(n10299), .B(n28715), .Z(n10300) );
  NANDN U19523 ( .A(n28716), .B(n10300), .Z(n10301) );
  NANDN U19524 ( .A(y[3270]), .B(x[3270]), .Z(n21594) );
  NANDN U19525 ( .A(y[3271]), .B(x[3271]), .Z(n21601) );
  AND U19526 ( .A(n21594), .B(n21601), .Z(n24054) );
  AND U19527 ( .A(n10301), .B(n24054), .Z(n10302) );
  NANDN U19528 ( .A(x[3271]), .B(y[3271]), .Z(n12030) );
  NANDN U19529 ( .A(x[3272]), .B(y[3272]), .Z(n12029) );
  NAND U19530 ( .A(n12030), .B(n12029), .Z(n28717) );
  OR U19531 ( .A(n10302), .B(n28717), .Z(n10303) );
  NAND U19532 ( .A(n28718), .B(n10303), .Z(n10304) );
  NANDN U19533 ( .A(n24053), .B(n10304), .Z(n10305) );
  NANDN U19534 ( .A(y[3274]), .B(x[3274]), .Z(n21606) );
  NANDN U19535 ( .A(y[3275]), .B(x[3275]), .Z(n21613) );
  AND U19536 ( .A(n21606), .B(n21613), .Z(n24052) );
  AND U19537 ( .A(n10305), .B(n24052), .Z(n10306) );
  NANDN U19538 ( .A(x[3275]), .B(y[3275]), .Z(n12026) );
  NANDN U19539 ( .A(x[3276]), .B(y[3276]), .Z(n12025) );
  NAND U19540 ( .A(n12026), .B(n12025), .Z(n28721) );
  OR U19541 ( .A(n10306), .B(n28721), .Z(n10307) );
  AND U19542 ( .A(n28722), .B(n10307), .Z(n10308) );
  OR U19543 ( .A(n28723), .B(n10308), .Z(n10309) );
  NAND U19544 ( .A(n28724), .B(n10309), .Z(n10310) );
  NANDN U19545 ( .A(n28725), .B(n10310), .Z(n10311) );
  NANDN U19546 ( .A(y[3280]), .B(x[3280]), .Z(n21626) );
  NANDN U19547 ( .A(y[3281]), .B(x[3281]), .Z(n21633) );
  AND U19548 ( .A(n21626), .B(n21633), .Z(n24051) );
  AND U19549 ( .A(n10311), .B(n24051), .Z(n10312) );
  NANDN U19550 ( .A(x[3281]), .B(y[3281]), .Z(n12022) );
  NANDN U19551 ( .A(x[3282]), .B(y[3282]), .Z(n12021) );
  AND U19552 ( .A(n12022), .B(n12021), .Z(n28726) );
  NANDN U19553 ( .A(n10312), .B(n28726), .Z(n10313) );
  NANDN U19554 ( .A(n28727), .B(n10313), .Z(n10314) );
  AND U19555 ( .A(n28728), .B(n10314), .Z(n10315) );
  OR U19556 ( .A(n28729), .B(n10315), .Z(n10316) );
  NAND U19557 ( .A(n28730), .B(n10316), .Z(n10317) );
  NANDN U19558 ( .A(n28731), .B(n10317), .Z(n10318) );
  AND U19559 ( .A(n28732), .B(n10318), .Z(n10319) );
  NANDN U19560 ( .A(y[3288]), .B(x[3288]), .Z(n21653) );
  NANDN U19561 ( .A(y[3289]), .B(x[3289]), .Z(n21660) );
  NAND U19562 ( .A(n21653), .B(n21660), .Z(n24050) );
  OR U19563 ( .A(n10319), .B(n24050), .Z(n10320) );
  AND U19564 ( .A(n10321), .B(n10320), .Z(n10322) );
  OR U19565 ( .A(n28736), .B(n10322), .Z(n10323) );
  NAND U19566 ( .A(n28737), .B(n10323), .Z(n10324) );
  NANDN U19567 ( .A(n28738), .B(n10324), .Z(n10325) );
  AND U19568 ( .A(n28739), .B(n10325), .Z(n10326) );
  NANDN U19569 ( .A(y[3294]), .B(x[3294]), .Z(n12014) );
  NANDN U19570 ( .A(y[3295]), .B(x[3295]), .Z(n12013) );
  NAND U19571 ( .A(n12014), .B(n12013), .Z(n28740) );
  OR U19572 ( .A(n10326), .B(n28740), .Z(n10327) );
  NANDN U19573 ( .A(x[3295]), .B(y[3295]), .Z(n21674) );
  NANDN U19574 ( .A(x[3296]), .B(y[3296]), .Z(n21681) );
  AND U19575 ( .A(n21674), .B(n21681), .Z(n24048) );
  AND U19576 ( .A(n10327), .B(n24048), .Z(n10328) );
  NANDN U19577 ( .A(y[3296]), .B(x[3296]), .Z(n12012) );
  NANDN U19578 ( .A(y[3297]), .B(x[3297]), .Z(n12011) );
  NAND U19579 ( .A(n12012), .B(n12011), .Z(n28741) );
  OR U19580 ( .A(n10328), .B(n28741), .Z(n10329) );
  NAND U19581 ( .A(n28742), .B(n10329), .Z(n10330) );
  NANDN U19582 ( .A(n24047), .B(n10330), .Z(n10331) );
  NANDN U19583 ( .A(x[3299]), .B(y[3299]), .Z(n12008) );
  NANDN U19584 ( .A(x[3300]), .B(y[3300]), .Z(n12005) );
  AND U19585 ( .A(n12008), .B(n12005), .Z(n24046) );
  AND U19586 ( .A(n10331), .B(n24046), .Z(n10332) );
  NANDN U19587 ( .A(y[3300]), .B(x[3300]), .Z(n12007) );
  NANDN U19588 ( .A(y[3301]), .B(x[3301]), .Z(n21692) );
  NAND U19589 ( .A(n12007), .B(n21692), .Z(n24045) );
  OR U19590 ( .A(n10332), .B(n24045), .Z(n10333) );
  AND U19591 ( .A(n10334), .B(n10333), .Z(n10335) );
  OR U19592 ( .A(n28744), .B(n10335), .Z(n10336) );
  NAND U19593 ( .A(n28745), .B(n10336), .Z(n10337) );
  NANDN U19594 ( .A(n28746), .B(n10337), .Z(n10338) );
  NANDN U19595 ( .A(x[3305]), .B(y[3305]), .Z(n12001) );
  NANDN U19596 ( .A(x[3306]), .B(y[3306]), .Z(n11998) );
  AND U19597 ( .A(n12001), .B(n11998), .Z(n24042) );
  AND U19598 ( .A(n10338), .B(n24042), .Z(n10339) );
  NANDN U19599 ( .A(y[3306]), .B(x[3306]), .Z(n11999) );
  NANDN U19600 ( .A(y[3307]), .B(x[3307]), .Z(n21708) );
  AND U19601 ( .A(n11999), .B(n21708), .Z(n28747) );
  NANDN U19602 ( .A(n10339), .B(n28747), .Z(n10340) );
  NANDN U19603 ( .A(n28748), .B(n10340), .Z(n10341) );
  AND U19604 ( .A(n28749), .B(n10341), .Z(n10342) );
  OR U19605 ( .A(n28750), .B(n10342), .Z(n10343) );
  NAND U19606 ( .A(n24041), .B(n10343), .Z(n10344) );
  NANDN U19607 ( .A(n28751), .B(n10344), .Z(n10346) );
  NANDN U19608 ( .A(y[3313]), .B(x[3313]), .Z(n21726) );
  NANDN U19609 ( .A(y[3312]), .B(x[3312]), .Z(n10345) );
  AND U19610 ( .A(n21726), .B(n10345), .Z(n28752) );
  AND U19611 ( .A(n10346), .B(n28752), .Z(n10347) );
  NANDN U19612 ( .A(x[3314]), .B(y[3314]), .Z(n11993) );
  ANDN U19613 ( .B(y[3313]), .A(x[3313]), .Z(n21723) );
  ANDN U19614 ( .B(n11993), .A(n21723), .Z(n28753) );
  NANDN U19615 ( .A(n10347), .B(n28753), .Z(n10348) );
  NANDN U19616 ( .A(n28754), .B(n10348), .Z(n10349) );
  AND U19617 ( .A(n11992), .B(n10349), .Z(n10350) );
  NANDN U19618 ( .A(x[3315]), .B(y[3315]), .Z(n28756) );
  AND U19619 ( .A(n10350), .B(n28756), .Z(n10352) );
  NANDN U19620 ( .A(y[3316]), .B(x[3316]), .Z(n10351) );
  NANDN U19621 ( .A(y[3317]), .B(x[3317]), .Z(n11990) );
  NAND U19622 ( .A(n10351), .B(n11990), .Z(n28757) );
  OR U19623 ( .A(n10352), .B(n28757), .Z(n10353) );
  AND U19624 ( .A(n28760), .B(n10353), .Z(n10354) );
  NANDN U19625 ( .A(y[3318]), .B(x[3318]), .Z(n11989) );
  NANDN U19626 ( .A(y[3319]), .B(x[3319]), .Z(n11988) );
  NAND U19627 ( .A(n11989), .B(n11988), .Z(n24040) );
  OR U19628 ( .A(n10354), .B(n24040), .Z(n10355) );
  NAND U19629 ( .A(n28761), .B(n10355), .Z(n10356) );
  NANDN U19630 ( .A(n28762), .B(n10356), .Z(n10357) );
  AND U19631 ( .A(n28763), .B(n10357), .Z(n10358) );
  NANDN U19632 ( .A(y[3322]), .B(x[3322]), .Z(n21749) );
  NANDN U19633 ( .A(y[3323]), .B(x[3323]), .Z(n21757) );
  AND U19634 ( .A(n21749), .B(n21757), .Z(n28764) );
  NANDN U19635 ( .A(n10358), .B(n28764), .Z(n10359) );
  NANDN U19636 ( .A(n24039), .B(n10359), .Z(n10360) );
  NANDN U19637 ( .A(y[3324]), .B(x[3324]), .Z(n21756) );
  NANDN U19638 ( .A(y[3325]), .B(x[3325]), .Z(n21763) );
  AND U19639 ( .A(n21756), .B(n21763), .Z(n24038) );
  AND U19640 ( .A(n10360), .B(n24038), .Z(n10361) );
  OR U19641 ( .A(n28765), .B(n10361), .Z(n10362) );
  NAND U19642 ( .A(n28766), .B(n10362), .Z(n10363) );
  NANDN U19643 ( .A(n28767), .B(n10363), .Z(n10364) );
  AND U19644 ( .A(n28768), .B(n10364), .Z(n10365) );
  NANDN U19645 ( .A(x[3329]), .B(y[3329]), .Z(n11979) );
  NANDN U19646 ( .A(x[3330]), .B(y[3330]), .Z(n11978) );
  NAND U19647 ( .A(n11979), .B(n11978), .Z(n28769) );
  OR U19648 ( .A(n10365), .B(n28769), .Z(n10366) );
  NANDN U19649 ( .A(y[3330]), .B(x[3330]), .Z(n21774) );
  NANDN U19650 ( .A(y[3331]), .B(x[3331]), .Z(n21781) );
  AND U19651 ( .A(n21774), .B(n21781), .Z(n24037) );
  AND U19652 ( .A(n10366), .B(n24037), .Z(n10367) );
  NANDN U19653 ( .A(x[3331]), .B(y[3331]), .Z(n11977) );
  NANDN U19654 ( .A(x[3332]), .B(y[3332]), .Z(n11976) );
  NAND U19655 ( .A(n11977), .B(n11976), .Z(n28770) );
  OR U19656 ( .A(n10367), .B(n28770), .Z(n10368) );
  NAND U19657 ( .A(n28773), .B(n10368), .Z(n10369) );
  NANDN U19658 ( .A(n24036), .B(n10369), .Z(n10370) );
  AND U19659 ( .A(n28774), .B(n10370), .Z(n10371) );
  NANDN U19660 ( .A(x[3335]), .B(y[3335]), .Z(n11973) );
  NANDN U19661 ( .A(x[3336]), .B(y[3336]), .Z(n21797) );
  AND U19662 ( .A(n11973), .B(n21797), .Z(n24035) );
  NANDN U19663 ( .A(n10371), .B(n24035), .Z(n10372) );
  NANDN U19664 ( .A(n28775), .B(n10372), .Z(n10373) );
  NANDN U19665 ( .A(x[3337]), .B(y[3337]), .Z(n21796) );
  NANDN U19666 ( .A(x[3338]), .B(y[3338]), .Z(n11972) );
  AND U19667 ( .A(n21796), .B(n11972), .Z(n28776) );
  AND U19668 ( .A(n10373), .B(n28776), .Z(n10374) );
  NANDN U19669 ( .A(y[3338]), .B(x[3338]), .Z(n21800) );
  NANDN U19670 ( .A(y[3339]), .B(x[3339]), .Z(n21807) );
  NAND U19671 ( .A(n21800), .B(n21807), .Z(n24034) );
  OR U19672 ( .A(n10374), .B(n24034), .Z(n10375) );
  NAND U19673 ( .A(n24033), .B(n10375), .Z(n10376) );
  NANDN U19674 ( .A(n28777), .B(n10376), .Z(n10377) );
  AND U19675 ( .A(n28778), .B(n10377), .Z(n10378) );
  NANDN U19676 ( .A(y[3342]), .B(x[3342]), .Z(n21812) );
  NANDN U19677 ( .A(y[3343]), .B(x[3343]), .Z(n21819) );
  NAND U19678 ( .A(n21812), .B(n21819), .Z(n28779) );
  OR U19679 ( .A(n10378), .B(n28779), .Z(n10379) );
  AND U19680 ( .A(n28780), .B(n10379), .Z(n10380) );
  OR U19681 ( .A(n28782), .B(n10380), .Z(n10381) );
  NAND U19682 ( .A(n24032), .B(n10381), .Z(n10382) );
  NANDN U19683 ( .A(n28783), .B(n10382), .Z(n10383) );
  NANDN U19684 ( .A(x[3347]), .B(y[3347]), .Z(n11963) );
  NANDN U19685 ( .A(x[3348]), .B(y[3348]), .Z(n11959) );
  AND U19686 ( .A(n11963), .B(n11959), .Z(n28784) );
  AND U19687 ( .A(n10383), .B(n28784), .Z(n10384) );
  NANDN U19688 ( .A(y[3348]), .B(x[3348]), .Z(n11961) );
  NANDN U19689 ( .A(y[3349]), .B(x[3349]), .Z(n11958) );
  NAND U19690 ( .A(n11961), .B(n11958), .Z(n24031) );
  OR U19691 ( .A(n10384), .B(n24031), .Z(n10385) );
  NAND U19692 ( .A(n24030), .B(n10385), .Z(n10386) );
  NANDN U19693 ( .A(n11957), .B(n10386), .Z(n10389) );
  NANDN U19694 ( .A(x[3352]), .B(y[3352]), .Z(n10388) );
  NANDN U19695 ( .A(x[3351]), .B(y[3351]), .Z(n10387) );
  AND U19696 ( .A(n10388), .B(n10387), .Z(n24029) );
  AND U19697 ( .A(n10389), .B(n24029), .Z(n10392) );
  NANDN U19698 ( .A(y[3353]), .B(x[3353]), .Z(n10391) );
  NANDN U19699 ( .A(y[3352]), .B(x[3352]), .Z(n10390) );
  NAND U19700 ( .A(n10391), .B(n10390), .Z(n28786) );
  OR U19701 ( .A(n10392), .B(n28786), .Z(n10393) );
  NANDN U19702 ( .A(n28787), .B(n10393), .Z(n10394) );
  AND U19703 ( .A(n28788), .B(n10394), .Z(n10395) );
  OR U19704 ( .A(n28789), .B(n10395), .Z(n10396) );
  NAND U19705 ( .A(n24028), .B(n10396), .Z(n10397) );
  NANDN U19706 ( .A(n28790), .B(n10397), .Z(n10398) );
  NANDN U19707 ( .A(y[3358]), .B(x[3358]), .Z(n11953) );
  NANDN U19708 ( .A(y[3359]), .B(x[3359]), .Z(n11952) );
  AND U19709 ( .A(n11953), .B(n11952), .Z(n28793) );
  AND U19710 ( .A(n10398), .B(n28793), .Z(n10399) );
  NANDN U19711 ( .A(x[3359]), .B(y[3359]), .Z(n21858) );
  NANDN U19712 ( .A(x[3360]), .B(y[3360]), .Z(n21865) );
  NAND U19713 ( .A(n21858), .B(n21865), .Z(n24027) );
  OR U19714 ( .A(n10399), .B(n24027), .Z(n10400) );
  NANDN U19715 ( .A(y[3360]), .B(x[3360]), .Z(n11951) );
  NANDN U19716 ( .A(y[3361]), .B(x[3361]), .Z(n11950) );
  AND U19717 ( .A(n11951), .B(n11950), .Z(n24026) );
  AND U19718 ( .A(n10400), .B(n24026), .Z(n10401) );
  NANDN U19719 ( .A(x[3361]), .B(y[3361]), .Z(n21864) );
  NANDN U19720 ( .A(x[3362]), .B(y[3362]), .Z(n11948) );
  NAND U19721 ( .A(n21864), .B(n11948), .Z(n28795) );
  OR U19722 ( .A(n10401), .B(n28795), .Z(n10402) );
  AND U19723 ( .A(n28796), .B(n10402), .Z(n10404) );
  XNOR U19724 ( .A(x[3364]), .B(y[3364]), .Z(n11947) );
  NANDN U19725 ( .A(x[3363]), .B(y[3363]), .Z(n24025) );
  AND U19726 ( .A(n11947), .B(n24025), .Z(n10403) );
  NANDN U19727 ( .A(n10404), .B(n10403), .Z(n10406) );
  NANDN U19728 ( .A(y[3364]), .B(x[3364]), .Z(n10405) );
  NANDN U19729 ( .A(y[3365]), .B(x[3365]), .Z(n11944) );
  AND U19730 ( .A(n10405), .B(n11944), .Z(n28797) );
  AND U19731 ( .A(n10406), .B(n28797), .Z(n10407) );
  ANDN U19732 ( .B(n10408), .A(n10407), .Z(n10410) );
  NANDN U19733 ( .A(y[3366]), .B(x[3366]), .Z(n10409) );
  NANDN U19734 ( .A(y[3367]), .B(x[3367]), .Z(n11943) );
  NAND U19735 ( .A(n10409), .B(n11943), .Z(n28800) );
  OR U19736 ( .A(n10410), .B(n28800), .Z(n10411) );
  NAND U19737 ( .A(n28801), .B(n10411), .Z(n10412) );
  NANDN U19738 ( .A(n24023), .B(n10412), .Z(n10413) );
  AND U19739 ( .A(n28803), .B(n10413), .Z(n10414) );
  NANDN U19740 ( .A(y[3370]), .B(x[3370]), .Z(n11940) );
  NANDN U19741 ( .A(y[3371]), .B(x[3371]), .Z(n21894) );
  NAND U19742 ( .A(n11940), .B(n21894), .Z(n28804) );
  OR U19743 ( .A(n10414), .B(n28804), .Z(n10415) );
  AND U19744 ( .A(n28805), .B(n10415), .Z(n10416) );
  OR U19745 ( .A(n28806), .B(n10416), .Z(n10417) );
  NAND U19746 ( .A(n28807), .B(n10417), .Z(n10418) );
  NANDN U19747 ( .A(n28808), .B(n10418), .Z(n10419) );
  NANDN U19748 ( .A(x[3375]), .B(y[3375]), .Z(n11936) );
  NANDN U19749 ( .A(x[3376]), .B(y[3376]), .Z(n11935) );
  AND U19750 ( .A(n11936), .B(n11935), .Z(n24022) );
  AND U19751 ( .A(n10419), .B(n24022), .Z(n10420) );
  NANDN U19752 ( .A(y[3376]), .B(x[3376]), .Z(n21905) );
  NANDN U19753 ( .A(y[3377]), .B(x[3377]), .Z(n21912) );
  AND U19754 ( .A(n21905), .B(n21912), .Z(n28809) );
  NANDN U19755 ( .A(n10420), .B(n28809), .Z(n10421) );
  NANDN U19756 ( .A(n28810), .B(n10421), .Z(n10422) );
  AND U19757 ( .A(n28811), .B(n10422), .Z(n10423) );
  OR U19758 ( .A(n28812), .B(n10423), .Z(n10424) );
  NAND U19759 ( .A(n24021), .B(n10424), .Z(n10425) );
  NANDN U19760 ( .A(n28813), .B(n10425), .Z(n10426) );
  NAND U19761 ( .A(n28814), .B(n10426), .Z(n10427) );
  NAND U19762 ( .A(n28815), .B(n10427), .Z(n10428) );
  NANDN U19763 ( .A(n28816), .B(n10428), .Z(n10429) );
  NANDN U19764 ( .A(x[3385]), .B(y[3385]), .Z(n11926) );
  NANDN U19765 ( .A(x[3386]), .B(y[3386]), .Z(n11925) );
  AND U19766 ( .A(n11926), .B(n11925), .Z(n24020) );
  AND U19767 ( .A(n10429), .B(n24020), .Z(n10430) );
  NANDN U19768 ( .A(y[3386]), .B(x[3386]), .Z(n21935) );
  NANDN U19769 ( .A(y[3387]), .B(x[3387]), .Z(n11923) );
  NAND U19770 ( .A(n21935), .B(n11923), .Z(n28819) );
  OR U19771 ( .A(n10430), .B(n28819), .Z(n10431) );
  NAND U19772 ( .A(n28821), .B(n10431), .Z(n10432) );
  NANDN U19773 ( .A(n24019), .B(n10432), .Z(n10435) );
  NANDN U19774 ( .A(x[3390]), .B(y[3390]), .Z(n10434) );
  NANDN U19775 ( .A(x[3389]), .B(y[3389]), .Z(n10433) );
  AND U19776 ( .A(n10434), .B(n10433), .Z(n24018) );
  AND U19777 ( .A(n10435), .B(n24018), .Z(n10438) );
  NANDN U19778 ( .A(y[3390]), .B(x[3390]), .Z(n10437) );
  NANDN U19779 ( .A(y[3391]), .B(x[3391]), .Z(n10436) );
  NAND U19780 ( .A(n10437), .B(n10436), .Z(n28822) );
  OR U19781 ( .A(n10438), .B(n28822), .Z(n10439) );
  NAND U19782 ( .A(n28823), .B(n10439), .Z(n10440) );
  NANDN U19783 ( .A(n28824), .B(n10440), .Z(n10443) );
  NANDN U19784 ( .A(x[3394]), .B(y[3394]), .Z(n10442) );
  NANDN U19785 ( .A(x[3393]), .B(y[3393]), .Z(n10441) );
  AND U19786 ( .A(n10442), .B(n10441), .Z(n28825) );
  AND U19787 ( .A(n10443), .B(n28825), .Z(n10444) );
  ANDN U19788 ( .B(x[3394]), .A(y[3394]), .Z(n21953) );
  NANDN U19789 ( .A(y[3395]), .B(x[3395]), .Z(n21958) );
  NANDN U19790 ( .A(n21953), .B(n21958), .Z(n24017) );
  OR U19791 ( .A(n10444), .B(n24017), .Z(n10445) );
  NAND U19792 ( .A(n24016), .B(n10445), .Z(n10446) );
  NANDN U19793 ( .A(n24015), .B(n10446), .Z(n10447) );
  AND U19794 ( .A(n21964), .B(n10447), .Z(n10448) );
  NANDN U19795 ( .A(x[3397]), .B(y[3397]), .Z(n24014) );
  NAND U19796 ( .A(n10448), .B(n24014), .Z(n10449) );
  NANDN U19797 ( .A(n28828), .B(n10449), .Z(n10450) );
  AND U19798 ( .A(n11920), .B(n10450), .Z(n10451) );
  NANDN U19799 ( .A(x[3399]), .B(y[3399]), .Z(n28829) );
  AND U19800 ( .A(n10451), .B(n28829), .Z(n10453) );
  NANDN U19801 ( .A(y[3400]), .B(x[3400]), .Z(n10452) );
  NANDN U19802 ( .A(y[3401]), .B(x[3401]), .Z(n11918) );
  NAND U19803 ( .A(n10452), .B(n11918), .Z(n28831) );
  OR U19804 ( .A(n10453), .B(n28831), .Z(n10454) );
  AND U19805 ( .A(n28832), .B(n10454), .Z(n10455) );
  NANDN U19806 ( .A(y[3402]), .B(x[3402]), .Z(n11917) );
  NANDN U19807 ( .A(y[3403]), .B(x[3403]), .Z(n11916) );
  NAND U19808 ( .A(n11917), .B(n11916), .Z(n24012) );
  OR U19809 ( .A(n10455), .B(n24012), .Z(n10456) );
  NAND U19810 ( .A(n28833), .B(n10456), .Z(n10457) );
  NANDN U19811 ( .A(n24011), .B(n10457), .Z(n10458) );
  AND U19812 ( .A(n21984), .B(n10458), .Z(n10459) );
  NANDN U19813 ( .A(x[3405]), .B(y[3405]), .Z(n24009) );
  AND U19814 ( .A(n10459), .B(n24009), .Z(n10461) );
  NANDN U19815 ( .A(y[3406]), .B(x[3406]), .Z(n10460) );
  NANDN U19816 ( .A(y[3407]), .B(x[3407]), .Z(n21990) );
  NAND U19817 ( .A(n10460), .B(n21990), .Z(n28834) );
  OR U19818 ( .A(n10461), .B(n28834), .Z(n10462) );
  AND U19819 ( .A(n28835), .B(n10462), .Z(n10463) );
  OR U19820 ( .A(n28836), .B(n10463), .Z(n10464) );
  NAND U19821 ( .A(n24008), .B(n10464), .Z(n10465) );
  NANDN U19822 ( .A(n28838), .B(n10465), .Z(n10466) );
  NANDN U19823 ( .A(x[3411]), .B(y[3411]), .Z(n11909) );
  NANDN U19824 ( .A(x[3412]), .B(y[3412]), .Z(n11908) );
  AND U19825 ( .A(n11909), .B(n11908), .Z(n28839) );
  AND U19826 ( .A(n10466), .B(n28839), .Z(n10467) );
  NANDN U19827 ( .A(y[3412]), .B(x[3412]), .Z(n22001) );
  NANDN U19828 ( .A(y[3413]), .B(x[3413]), .Z(n22008) );
  AND U19829 ( .A(n22001), .B(n22008), .Z(n28840) );
  NANDN U19830 ( .A(n10467), .B(n28840), .Z(n10468) );
  NANDN U19831 ( .A(n28841), .B(n10468), .Z(n10469) );
  NANDN U19832 ( .A(y[3414]), .B(x[3414]), .Z(n22007) );
  NANDN U19833 ( .A(y[3415]), .B(x[3415]), .Z(n22014) );
  AND U19834 ( .A(n22007), .B(n22014), .Z(n24007) );
  AND U19835 ( .A(n10469), .B(n24007), .Z(n10470) );
  NANDN U19836 ( .A(x[3415]), .B(y[3415]), .Z(n11905) );
  NANDN U19837 ( .A(x[3416]), .B(y[3416]), .Z(n11904) );
  NAND U19838 ( .A(n11905), .B(n11904), .Z(n28842) );
  OR U19839 ( .A(n10470), .B(n28842), .Z(n10471) );
  NAND U19840 ( .A(n28843), .B(n10471), .Z(n10472) );
  NANDN U19841 ( .A(n24006), .B(n10472), .Z(n10473) );
  NANDN U19842 ( .A(y[3418]), .B(x[3418]), .Z(n22019) );
  NANDN U19843 ( .A(y[3419]), .B(x[3419]), .Z(n22026) );
  AND U19844 ( .A(n22019), .B(n22026), .Z(n24005) );
  AND U19845 ( .A(n10473), .B(n24005), .Z(n10474) );
  NANDN U19846 ( .A(x[3419]), .B(y[3419]), .Z(n11901) );
  NANDN U19847 ( .A(x[3420]), .B(y[3420]), .Z(n11900) );
  NAND U19848 ( .A(n11901), .B(n11900), .Z(n28844) );
  OR U19849 ( .A(n10474), .B(n28844), .Z(n10475) );
  AND U19850 ( .A(n28845), .B(n10475), .Z(n10476) );
  OR U19851 ( .A(n28847), .B(n10476), .Z(n10477) );
  NAND U19852 ( .A(n28848), .B(n10477), .Z(n10478) );
  NANDN U19853 ( .A(n28849), .B(n10478), .Z(n10479) );
  NANDN U19854 ( .A(y[3424]), .B(x[3424]), .Z(n22037) );
  NANDN U19855 ( .A(y[3425]), .B(x[3425]), .Z(n22044) );
  AND U19856 ( .A(n22037), .B(n22044), .Z(n24004) );
  AND U19857 ( .A(n10479), .B(n24004), .Z(n10480) );
  NANDN U19858 ( .A(x[3425]), .B(y[3425]), .Z(n11895) );
  NANDN U19859 ( .A(x[3426]), .B(y[3426]), .Z(n11894) );
  AND U19860 ( .A(n11895), .B(n11894), .Z(n28850) );
  NANDN U19861 ( .A(n10480), .B(n28850), .Z(n10481) );
  NANDN U19862 ( .A(n28851), .B(n10481), .Z(n10482) );
  AND U19863 ( .A(n28852), .B(n10482), .Z(n10483) );
  OR U19864 ( .A(n28853), .B(n10483), .Z(n10484) );
  NAND U19865 ( .A(n24003), .B(n10484), .Z(n10485) );
  NANDN U19866 ( .A(n28854), .B(n10485), .Z(n10486) );
  NANDN U19867 ( .A(x[3431]), .B(y[3431]), .Z(n11889) );
  NANDN U19868 ( .A(x[3432]), .B(y[3432]), .Z(n11886) );
  AND U19869 ( .A(n11889), .B(n11886), .Z(n28855) );
  AND U19870 ( .A(n10486), .B(n28855), .Z(n10487) );
  NANDN U19871 ( .A(y[3432]), .B(x[3432]), .Z(n11887) );
  NANDN U19872 ( .A(y[3433]), .B(x[3433]), .Z(n11884) );
  NAND U19873 ( .A(n11887), .B(n11884), .Z(n24002) );
  OR U19874 ( .A(n10487), .B(n24002), .Z(n10488) );
  AND U19875 ( .A(n10489), .B(n10488), .Z(n10491) );
  NANDN U19876 ( .A(y[3434]), .B(x[3434]), .Z(n10490) );
  NANDN U19877 ( .A(y[3435]), .B(x[3435]), .Z(n22072) );
  NAND U19878 ( .A(n10490), .B(n22072), .Z(n24000) );
  OR U19879 ( .A(n10491), .B(n24000), .Z(n10492) );
  NAND U19880 ( .A(n28858), .B(n10492), .Z(n10493) );
  NANDN U19881 ( .A(n28859), .B(n10493), .Z(n10494) );
  NANDN U19882 ( .A(x[3437]), .B(y[3437]), .Z(n11882) );
  NANDN U19883 ( .A(x[3438]), .B(y[3438]), .Z(n11881) );
  AND U19884 ( .A(n11882), .B(n11881), .Z(n28860) );
  AND U19885 ( .A(n10494), .B(n28860), .Z(n10495) );
  NANDN U19886 ( .A(y[3438]), .B(x[3438]), .Z(n22077) );
  NANDN U19887 ( .A(y[3439]), .B(x[3439]), .Z(n22084) );
  NAND U19888 ( .A(n22077), .B(n22084), .Z(n23999) );
  OR U19889 ( .A(n10495), .B(n23999), .Z(n10496) );
  NANDN U19890 ( .A(x[3439]), .B(y[3439]), .Z(n11880) );
  NANDN U19891 ( .A(x[3440]), .B(y[3440]), .Z(n11879) );
  AND U19892 ( .A(n11880), .B(n11879), .Z(n23998) );
  AND U19893 ( .A(n10496), .B(n23998), .Z(n10497) );
  NANDN U19894 ( .A(y[3440]), .B(x[3440]), .Z(n22083) );
  NANDN U19895 ( .A(y[3441]), .B(x[3441]), .Z(n22090) );
  NAND U19896 ( .A(n22083), .B(n22090), .Z(n28861) );
  OR U19897 ( .A(n10497), .B(n28861), .Z(n10498) );
  NAND U19898 ( .A(n28862), .B(n10498), .Z(n10499) );
  NANDN U19899 ( .A(n28863), .B(n10499), .Z(n10500) );
  AND U19900 ( .A(n28864), .B(n10500), .Z(n10501) );
  OR U19901 ( .A(n28865), .B(n10501), .Z(n10502) );
  NAND U19902 ( .A(n28866), .B(n10502), .Z(n10503) );
  NANDN U19903 ( .A(n28867), .B(n10503), .Z(n10504) );
  AND U19904 ( .A(n28868), .B(n10504), .Z(n10505) );
  NANDN U19905 ( .A(y[3448]), .B(x[3448]), .Z(n11871) );
  NANDN U19906 ( .A(y[3449]), .B(x[3449]), .Z(n22110) );
  NAND U19907 ( .A(n11871), .B(n22110), .Z(n28869) );
  OR U19908 ( .A(n10505), .B(n28869), .Z(n10506) );
  AND U19909 ( .A(n22111), .B(n10506), .Z(n10507) );
  NANDN U19910 ( .A(x[3449]), .B(y[3449]), .Z(n23996) );
  AND U19911 ( .A(n10507), .B(n23996), .Z(n10509) );
  NANDN U19912 ( .A(y[3450]), .B(x[3450]), .Z(n10508) );
  NANDN U19913 ( .A(y[3451]), .B(x[3451]), .Z(n11868) );
  NAND U19914 ( .A(n10508), .B(n11868), .Z(n28871) );
  OR U19915 ( .A(n10509), .B(n28871), .Z(n10510) );
  AND U19916 ( .A(n28872), .B(n10510), .Z(n10511) );
  NANDN U19917 ( .A(y[3452]), .B(x[3452]), .Z(n11867) );
  NANDN U19918 ( .A(y[3453]), .B(x[3453]), .Z(n11864) );
  NAND U19919 ( .A(n11867), .B(n11864), .Z(n23995) );
  OR U19920 ( .A(n10511), .B(n23995), .Z(n10512) );
  NAND U19921 ( .A(n28873), .B(n10512), .Z(n10513) );
  NANDN U19922 ( .A(n23994), .B(n10513), .Z(n10514) );
  AND U19923 ( .A(n28874), .B(n10514), .Z(n10516) );
  NANDN U19924 ( .A(y[3457]), .B(x[3457]), .Z(n22130) );
  NANDN U19925 ( .A(y[3456]), .B(x[3456]), .Z(n10515) );
  NAND U19926 ( .A(n22130), .B(n10515), .Z(n11861) );
  OR U19927 ( .A(n10516), .B(n11861), .Z(n10517) );
  NAND U19928 ( .A(n11860), .B(n10517), .Z(n10518) );
  NANDN U19929 ( .A(n11859), .B(n10518), .Z(n10519) );
  AND U19930 ( .A(n28878), .B(n10519), .Z(n10520) );
  NANDN U19931 ( .A(y[3460]), .B(x[3460]), .Z(n22137) );
  NANDN U19932 ( .A(y[3461]), .B(x[3461]), .Z(n11856) );
  AND U19933 ( .A(n22137), .B(n11856), .Z(n28879) );
  NANDN U19934 ( .A(n10520), .B(n28879), .Z(n10521) );
  NANDN U19935 ( .A(n28880), .B(n10521), .Z(n10522) );
  AND U19936 ( .A(n28881), .B(n10522), .Z(n10523) );
  OR U19937 ( .A(n28882), .B(n10523), .Z(n10524) );
  NAND U19938 ( .A(n28883), .B(n10524), .Z(n10525) );
  NANDN U19939 ( .A(n28885), .B(n10525), .Z(n10526) );
  AND U19940 ( .A(n28886), .B(n10526), .Z(n10527) );
  NANDN U19941 ( .A(x[3467]), .B(y[3467]), .Z(n11849) );
  NANDN U19942 ( .A(x[3468]), .B(y[3468]), .Z(n11846) );
  AND U19943 ( .A(n11849), .B(n11846), .Z(n28887) );
  NANDN U19944 ( .A(n10527), .B(n28887), .Z(n10528) );
  NANDN U19945 ( .A(n23993), .B(n10528), .Z(n10529) );
  AND U19946 ( .A(n22163), .B(n10529), .Z(n10530) );
  NANDN U19947 ( .A(x[3469]), .B(y[3469]), .Z(n23992) );
  AND U19948 ( .A(n10530), .B(n23992), .Z(n10532) );
  NANDN U19949 ( .A(y[3470]), .B(x[3470]), .Z(n10531) );
  NANDN U19950 ( .A(y[3471]), .B(x[3471]), .Z(n11845) );
  NAND U19951 ( .A(n10531), .B(n11845), .Z(n28889) );
  OR U19952 ( .A(n10532), .B(n28889), .Z(n10533) );
  NANDN U19953 ( .A(x[3471]), .B(y[3471]), .Z(n22165) );
  NANDN U19954 ( .A(x[3472]), .B(y[3472]), .Z(n22172) );
  AND U19955 ( .A(n22165), .B(n22172), .Z(n28890) );
  AND U19956 ( .A(n10533), .B(n28890), .Z(n10534) );
  NANDN U19957 ( .A(y[3472]), .B(x[3472]), .Z(n11844) );
  NANDN U19958 ( .A(y[3473]), .B(x[3473]), .Z(n11843) );
  NAND U19959 ( .A(n11844), .B(n11843), .Z(n28891) );
  OR U19960 ( .A(n10534), .B(n28891), .Z(n10535) );
  NAND U19961 ( .A(n28892), .B(n10535), .Z(n10536) );
  NANDN U19962 ( .A(n23991), .B(n10536), .Z(n10537) );
  NANDN U19963 ( .A(x[3475]), .B(y[3475]), .Z(n22177) );
  NANDN U19964 ( .A(x[3476]), .B(y[3476]), .Z(n22184) );
  AND U19965 ( .A(n22177), .B(n22184), .Z(n23990) );
  AND U19966 ( .A(n10537), .B(n23990), .Z(n10538) );
  NANDN U19967 ( .A(y[3476]), .B(x[3476]), .Z(n11840) );
  NANDN U19968 ( .A(y[3477]), .B(x[3477]), .Z(n11839) );
  AND U19969 ( .A(n11840), .B(n11839), .Z(n28894) );
  NANDN U19970 ( .A(n10538), .B(n28894), .Z(n10539) );
  NANDN U19971 ( .A(n28895), .B(n10539), .Z(n10540) );
  AND U19972 ( .A(n28896), .B(n10540), .Z(n10541) );
  OR U19973 ( .A(n28897), .B(n10541), .Z(n10542) );
  NAND U19974 ( .A(n28898), .B(n10542), .Z(n10543) );
  NANDN U19975 ( .A(n28899), .B(n10543), .Z(n10544) );
  NAND U19976 ( .A(n28900), .B(n10544), .Z(n10545) );
  NAND U19977 ( .A(n28901), .B(n10545), .Z(n10546) );
  NANDN U19978 ( .A(n23989), .B(n10546), .Z(n10547) );
  AND U19979 ( .A(n22207), .B(n10547), .Z(n10548) );
  NAND U19980 ( .A(n28902), .B(n10548), .Z(n10550) );
  NANDN U19981 ( .A(y[3486]), .B(x[3486]), .Z(n10549) );
  NANDN U19982 ( .A(y[3487]), .B(x[3487]), .Z(n11827) );
  AND U19983 ( .A(n10549), .B(n11827), .Z(n28904) );
  AND U19984 ( .A(n10550), .B(n28904), .Z(n10551) );
  ANDN U19985 ( .B(n28905), .A(n10551), .Z(n10552) );
  OR U19986 ( .A(n28906), .B(n10552), .Z(n10553) );
  NAND U19987 ( .A(n28908), .B(n10553), .Z(n10554) );
  NANDN U19988 ( .A(n28909), .B(n10554), .Z(n10555) );
  AND U19989 ( .A(n28910), .B(n10555), .Z(n10556) );
  NANDN U19990 ( .A(y[3492]), .B(x[3492]), .Z(n11824) );
  NANDN U19991 ( .A(y[3493]), .B(x[3493]), .Z(n11823) );
  NAND U19992 ( .A(n11824), .B(n11823), .Z(n28911) );
  OR U19993 ( .A(n10556), .B(n28911), .Z(n10557) );
  NANDN U19994 ( .A(x[3493]), .B(y[3493]), .Z(n22228) );
  NANDN U19995 ( .A(x[3494]), .B(y[3494]), .Z(n22235) );
  AND U19996 ( .A(n22228), .B(n22235), .Z(n23988) );
  AND U19997 ( .A(n10557), .B(n23988), .Z(n10558) );
  NANDN U19998 ( .A(y[3494]), .B(x[3494]), .Z(n11822) );
  NANDN U19999 ( .A(y[3495]), .B(x[3495]), .Z(n11821) );
  NAND U20000 ( .A(n11822), .B(n11821), .Z(n28912) );
  OR U20001 ( .A(n10558), .B(n28912), .Z(n10559) );
  NAND U20002 ( .A(n28913), .B(n10559), .Z(n10560) );
  NANDN U20003 ( .A(n23987), .B(n10560), .Z(n10561) );
  NANDN U20004 ( .A(x[3497]), .B(y[3497]), .Z(n22240) );
  NANDN U20005 ( .A(x[3498]), .B(y[3498]), .Z(n22247) );
  AND U20006 ( .A(n22240), .B(n22247), .Z(n23986) );
  AND U20007 ( .A(n10561), .B(n23986), .Z(n10562) );
  NANDN U20008 ( .A(y[3498]), .B(x[3498]), .Z(n11818) );
  NANDN U20009 ( .A(y[3499]), .B(x[3499]), .Z(n11817) );
  AND U20010 ( .A(n11818), .B(n11817), .Z(n28914) );
  NANDN U20011 ( .A(n10562), .B(n28914), .Z(n10563) );
  NANDN U20012 ( .A(n28915), .B(n10563), .Z(n10564) );
  AND U20013 ( .A(n28916), .B(n10564), .Z(n10565) );
  OR U20014 ( .A(n28917), .B(n10565), .Z(n10566) );
  NAND U20015 ( .A(n28918), .B(n10566), .Z(n10567) );
  NANDN U20016 ( .A(n28920), .B(n10567), .Z(n10568) );
  AND U20017 ( .A(n28921), .B(n10568), .Z(n10569) );
  NANDN U20018 ( .A(x[3505]), .B(y[3505]), .Z(n22264) );
  NANDN U20019 ( .A(x[3506]), .B(y[3506]), .Z(n22271) );
  NAND U20020 ( .A(n22264), .B(n22271), .Z(n28922) );
  OR U20021 ( .A(n10569), .B(n28922), .Z(n10570) );
  NANDN U20022 ( .A(y[3506]), .B(x[3506]), .Z(n11810) );
  NANDN U20023 ( .A(y[3507]), .B(x[3507]), .Z(n11809) );
  AND U20024 ( .A(n11810), .B(n11809), .Z(n23985) );
  AND U20025 ( .A(n10570), .B(n23985), .Z(n10571) );
  NANDN U20026 ( .A(x[3507]), .B(y[3507]), .Z(n22270) );
  NANDN U20027 ( .A(x[3508]), .B(y[3508]), .Z(n22277) );
  NAND U20028 ( .A(n22270), .B(n22277), .Z(n28923) );
  OR U20029 ( .A(n10571), .B(n28923), .Z(n10572) );
  NAND U20030 ( .A(n28924), .B(n10572), .Z(n10573) );
  NANDN U20031 ( .A(n23984), .B(n10573), .Z(n10574) );
  NANDN U20032 ( .A(y[3510]), .B(x[3510]), .Z(n11806) );
  NANDN U20033 ( .A(y[3511]), .B(x[3511]), .Z(n11802) );
  AND U20034 ( .A(n11806), .B(n11802), .Z(n23983) );
  AND U20035 ( .A(n10574), .B(n23983), .Z(n10575) );
  NANDN U20036 ( .A(x[3511]), .B(y[3511]), .Z(n11804) );
  NANDN U20037 ( .A(x[3512]), .B(y[3512]), .Z(n11801) );
  AND U20038 ( .A(n11804), .B(n11801), .Z(n28925) );
  NANDN U20039 ( .A(n10575), .B(n28925), .Z(n10576) );
  NANDN U20040 ( .A(n28926), .B(n10576), .Z(n10577) );
  AND U20041 ( .A(n11800), .B(n10577), .Z(n10578) );
  NANDN U20042 ( .A(x[3513]), .B(y[3513]), .Z(n23981) );
  AND U20043 ( .A(n10578), .B(n23981), .Z(n10580) );
  NANDN U20044 ( .A(y[3514]), .B(x[3514]), .Z(n10579) );
  NANDN U20045 ( .A(y[3515]), .B(x[3515]), .Z(n11798) );
  NAND U20046 ( .A(n10579), .B(n11798), .Z(n28927) );
  OR U20047 ( .A(n10580), .B(n28927), .Z(n10581) );
  NAND U20048 ( .A(n28928), .B(n10581), .Z(n10582) );
  NANDN U20049 ( .A(y[3516]), .B(x[3516]), .Z(n11797) );
  NANDN U20050 ( .A(y[3517]), .B(x[3517]), .Z(n11795) );
  AND U20051 ( .A(n11797), .B(n11795), .Z(n23980) );
  AND U20052 ( .A(n10582), .B(n23980), .Z(n10583) );
  ANDN U20053 ( .B(n28930), .A(n10583), .Z(n10584) );
  NAND U20054 ( .A(n11796), .B(n10584), .Z(n10585) );
  NANDN U20055 ( .A(n23979), .B(n10585), .Z(n10586) );
  NANDN U20056 ( .A(x[3519]), .B(y[3519]), .Z(n22301) );
  NANDN U20057 ( .A(x[3520]), .B(y[3520]), .Z(n22306) );
  AND U20058 ( .A(n22301), .B(n22306), .Z(n23978) );
  AND U20059 ( .A(n10586), .B(n23978), .Z(n10587) );
  NANDN U20060 ( .A(y[3520]), .B(x[3520]), .Z(n11793) );
  NANDN U20061 ( .A(y[3521]), .B(x[3521]), .Z(n11791) );
  AND U20062 ( .A(n11793), .B(n11791), .Z(n28932) );
  NANDN U20063 ( .A(n10587), .B(n28932), .Z(n10588) );
  NAND U20064 ( .A(n10589), .B(n10588), .Z(n10591) );
  NANDN U20065 ( .A(y[3522]), .B(x[3522]), .Z(n10590) );
  NANDN U20066 ( .A(y[3523]), .B(x[3523]), .Z(n11788) );
  AND U20067 ( .A(n10590), .B(n11788), .Z(n23977) );
  AND U20068 ( .A(n10591), .B(n23977), .Z(n10592) );
  NOR U20069 ( .A(n11790), .B(n10592), .Z(n10593) );
  NAND U20070 ( .A(n11789), .B(n10593), .Z(n10594) );
  NANDN U20071 ( .A(n28937), .B(n10594), .Z(n10595) );
  AND U20072 ( .A(n22318), .B(n10595), .Z(n10596) );
  NANDN U20073 ( .A(n11787), .B(n10596), .Z(n10597) );
  NAND U20074 ( .A(n28940), .B(n10597), .Z(n10598) );
  NAND U20075 ( .A(n22324), .B(n10598), .Z(n10599) );
  ANDN U20076 ( .B(y[3527]), .A(x[3527]), .Z(n11786) );
  OR U20077 ( .A(n10599), .B(n11786), .Z(n10600) );
  NAND U20078 ( .A(n28942), .B(n10600), .Z(n10602) );
  NANDN U20079 ( .A(x[3529]), .B(y[3529]), .Z(n28944) );
  XNOR U20080 ( .A(x[3530]), .B(y[3530]), .Z(n11785) );
  NAND U20081 ( .A(n28944), .B(n11785), .Z(n10601) );
  ANDN U20082 ( .B(n10602), .A(n10601), .Z(n10603) );
  OR U20083 ( .A(n28945), .B(n10603), .Z(n10604) );
  NAND U20084 ( .A(n28946), .B(n10604), .Z(n10605) );
  NANDN U20085 ( .A(n28947), .B(n10605), .Z(n10606) );
  AND U20086 ( .A(n11780), .B(n10606), .Z(n10607) );
  NANDN U20087 ( .A(x[3533]), .B(y[3533]), .Z(n23974) );
  AND U20088 ( .A(n10607), .B(n23974), .Z(n10609) );
  NANDN U20089 ( .A(y[3534]), .B(x[3534]), .Z(n10608) );
  NANDN U20090 ( .A(y[3535]), .B(x[3535]), .Z(n11778) );
  NAND U20091 ( .A(n10608), .B(n11778), .Z(n28948) );
  OR U20092 ( .A(n10609), .B(n28948), .Z(n10610) );
  AND U20093 ( .A(n28949), .B(n10610), .Z(n10611) );
  OR U20094 ( .A(n28950), .B(n10611), .Z(n10612) );
  NAND U20095 ( .A(n28951), .B(n10612), .Z(n10613) );
  NANDN U20096 ( .A(n28952), .B(n10613), .Z(n10614) );
  AND U20097 ( .A(n28953), .B(n10614), .Z(n10615) );
  NANDN U20098 ( .A(y[3540]), .B(x[3540]), .Z(n22353) );
  NANDN U20099 ( .A(y[3541]), .B(x[3541]), .Z(n22360) );
  NAND U20100 ( .A(n22353), .B(n22360), .Z(n28954) );
  OR U20101 ( .A(n10615), .B(n28954), .Z(n10616) );
  AND U20102 ( .A(n28955), .B(n10616), .Z(n10617) );
  OR U20103 ( .A(n28957), .B(n10617), .Z(n10618) );
  NAND U20104 ( .A(n28958), .B(n10618), .Z(n10619) );
  NANDN U20105 ( .A(n28959), .B(n10619), .Z(n10620) );
  NAND U20106 ( .A(n23972), .B(n10620), .Z(n10621) );
  NAND U20107 ( .A(n28960), .B(n10621), .Z(n10622) );
  NANDN U20108 ( .A(n28961), .B(n10622), .Z(n10623) );
  AND U20109 ( .A(n28962), .B(n10623), .Z(n10624) );
  OR U20110 ( .A(n28963), .B(n10624), .Z(n10625) );
  NAND U20111 ( .A(n28964), .B(n10625), .Z(n10626) );
  NANDN U20112 ( .A(n28965), .B(n10626), .Z(n10627) );
  AND U20113 ( .A(n28966), .B(n10627), .Z(n10628) );
  NANDN U20114 ( .A(x[3553]), .B(y[3553]), .Z(n11757) );
  NANDN U20115 ( .A(x[3554]), .B(y[3554]), .Z(n11756) );
  NAND U20116 ( .A(n11757), .B(n11756), .Z(n28967) );
  OR U20117 ( .A(n10628), .B(n28967), .Z(n10629) );
  AND U20118 ( .A(n28968), .B(n10629), .Z(n10630) );
  OR U20119 ( .A(n28969), .B(n10630), .Z(n10631) );
  NAND U20120 ( .A(n28970), .B(n10631), .Z(n10632) );
  NAND U20121 ( .A(n28971), .B(n10632), .Z(n10633) );
  NAND U20122 ( .A(n28972), .B(n10633), .Z(n10636) );
  NANDN U20123 ( .A(x[3560]), .B(y[3560]), .Z(n10635) );
  NANDN U20124 ( .A(x[3559]), .B(y[3559]), .Z(n10634) );
  AND U20125 ( .A(n10635), .B(n10634), .Z(n11754) );
  AND U20126 ( .A(n10636), .B(n11754), .Z(n10639) );
  NANDN U20127 ( .A(y[3561]), .B(x[3561]), .Z(n10638) );
  NANDN U20128 ( .A(y[3560]), .B(x[3560]), .Z(n10637) );
  AND U20129 ( .A(n10638), .B(n10637), .Z(n28975) );
  NANDN U20130 ( .A(n10639), .B(n28975), .Z(n10640) );
  NANDN U20131 ( .A(n28976), .B(n10640), .Z(n10641) );
  NANDN U20132 ( .A(y[3562]), .B(x[3562]), .Z(n22413) );
  NANDN U20133 ( .A(y[3563]), .B(x[3563]), .Z(n11753) );
  AND U20134 ( .A(n22413), .B(n11753), .Z(n28978) );
  AND U20135 ( .A(n10641), .B(n28978), .Z(n10642) );
  ANDN U20136 ( .B(y[3563]), .A(x[3563]), .Z(n22415) );
  NANDN U20137 ( .A(x[3564]), .B(y[3564]), .Z(n11751) );
  NANDN U20138 ( .A(n22415), .B(n11751), .Z(n28979) );
  OR U20139 ( .A(n10642), .B(n28979), .Z(n10643) );
  NAND U20140 ( .A(n28980), .B(n10643), .Z(n10644) );
  NANDN U20141 ( .A(n23971), .B(n10644), .Z(n10645) );
  NANDN U20142 ( .A(y[3566]), .B(x[3566]), .Z(n11748) );
  NANDN U20143 ( .A(y[3567]), .B(x[3567]), .Z(n22427) );
  AND U20144 ( .A(n11748), .B(n22427), .Z(n23970) );
  AND U20145 ( .A(n10645), .B(n23970), .Z(n10646) );
  NANDN U20146 ( .A(x[3567]), .B(y[3567]), .Z(n22422) );
  NANDN U20147 ( .A(x[3568]), .B(y[3568]), .Z(n11747) );
  NAND U20148 ( .A(n22422), .B(n11747), .Z(n28981) );
  OR U20149 ( .A(n10646), .B(n28981), .Z(n10647) );
  AND U20150 ( .A(n28982), .B(n10647), .Z(n10648) );
  OR U20151 ( .A(n28983), .B(n10648), .Z(n10649) );
  NAND U20152 ( .A(n28984), .B(n10649), .Z(n10650) );
  NANDN U20153 ( .A(n28985), .B(n10650), .Z(n10652) );
  NANDN U20154 ( .A(y[3573]), .B(x[3573]), .Z(n11742) );
  NANDN U20155 ( .A(y[3572]), .B(x[3572]), .Z(n10651) );
  NAND U20156 ( .A(n11742), .B(n10651), .Z(n28986) );
  ANDN U20157 ( .B(n10652), .A(n28986), .Z(n10655) );
  NANDN U20158 ( .A(x[3573]), .B(y[3573]), .Z(n10654) );
  NANDN U20159 ( .A(x[3574]), .B(y[3574]), .Z(n10653) );
  AND U20160 ( .A(n10654), .B(n10653), .Z(n28987) );
  NANDN U20161 ( .A(n10655), .B(n28987), .Z(n10656) );
  NAND U20162 ( .A(n28989), .B(n10656), .Z(n10657) );
  NANDN U20163 ( .A(n28990), .B(n10657), .Z(n10658) );
  AND U20164 ( .A(n28991), .B(n10658), .Z(n10659) );
  NANDN U20165 ( .A(x[3577]), .B(y[3577]), .Z(n22450) );
  NANDN U20166 ( .A(x[3578]), .B(y[3578]), .Z(n22458) );
  AND U20167 ( .A(n22450), .B(n22458), .Z(n28992) );
  NANDN U20168 ( .A(n10659), .B(n28992), .Z(n10660) );
  NANDN U20169 ( .A(n28993), .B(n10660), .Z(n10661) );
  AND U20170 ( .A(n28994), .B(n10661), .Z(n10662) );
  OR U20171 ( .A(n28995), .B(n10662), .Z(n10663) );
  NAND U20172 ( .A(n28996), .B(n10663), .Z(n10664) );
  NANDN U20173 ( .A(n28997), .B(n10664), .Z(n10665) );
  AND U20174 ( .A(n28998), .B(n10665), .Z(n10666) );
  NANDN U20175 ( .A(y[3584]), .B(x[3584]), .Z(n11736) );
  NANDN U20176 ( .A(y[3585]), .B(x[3585]), .Z(n22480) );
  NAND U20177 ( .A(n11736), .B(n22480), .Z(n28999) );
  OR U20178 ( .A(n10666), .B(n28999), .Z(n10667) );
  AND U20179 ( .A(n29000), .B(n10667), .Z(n10668) );
  OR U20180 ( .A(n29001), .B(n10668), .Z(n10669) );
  NAND U20181 ( .A(n29002), .B(n10669), .Z(n10670) );
  NANDN U20182 ( .A(n29003), .B(n10670), .Z(n10671) );
  AND U20183 ( .A(n29004), .B(n10671), .Z(n10672) );
  NANDN U20184 ( .A(y[3590]), .B(x[3590]), .Z(n11732) );
  NANDN U20185 ( .A(y[3591]), .B(x[3591]), .Z(n11731) );
  AND U20186 ( .A(n11732), .B(n11731), .Z(n29005) );
  NANDN U20187 ( .A(n10672), .B(n29005), .Z(n10673) );
  NANDN U20188 ( .A(n23969), .B(n10673), .Z(n10674) );
  NANDN U20189 ( .A(y[3592]), .B(x[3592]), .Z(n11730) );
  NANDN U20190 ( .A(y[3593]), .B(x[3593]), .Z(n11729) );
  AND U20191 ( .A(n11730), .B(n11729), .Z(n23968) );
  AND U20192 ( .A(n10674), .B(n23968), .Z(n10675) );
  NANDN U20193 ( .A(x[3593]), .B(y[3593]), .Z(n22501) );
  NANDN U20194 ( .A(x[3594]), .B(y[3594]), .Z(n22508) );
  NAND U20195 ( .A(n22501), .B(n22508), .Z(n29008) );
  OR U20196 ( .A(n10675), .B(n29008), .Z(n10676) );
  NAND U20197 ( .A(n29009), .B(n10676), .Z(n10677) );
  NANDN U20198 ( .A(n23967), .B(n10677), .Z(n10678) );
  NANDN U20199 ( .A(y[3596]), .B(x[3596]), .Z(n11726) );
  NANDN U20200 ( .A(y[3597]), .B(x[3597]), .Z(n11725) );
  AND U20201 ( .A(n11726), .B(n11725), .Z(n23966) );
  AND U20202 ( .A(n10678), .B(n23966), .Z(n10679) );
  NANDN U20203 ( .A(x[3597]), .B(y[3597]), .Z(n22513) );
  ANDN U20204 ( .B(y[3598]), .A(x[3598]), .Z(n22520) );
  ANDN U20205 ( .B(n22513), .A(n22520), .Z(n29010) );
  NANDN U20206 ( .A(n10679), .B(n29010), .Z(n10680) );
  NANDN U20207 ( .A(n29011), .B(n10680), .Z(n10681) );
  AND U20208 ( .A(n11723), .B(n10681), .Z(n10682) );
  NANDN U20209 ( .A(x[3599]), .B(y[3599]), .Z(n23965) );
  AND U20210 ( .A(n10682), .B(n23965), .Z(n10684) );
  NANDN U20211 ( .A(y[3600]), .B(x[3600]), .Z(n10683) );
  NANDN U20212 ( .A(y[3601]), .B(x[3601]), .Z(n11721) );
  NAND U20213 ( .A(n10683), .B(n11721), .Z(n29012) );
  OR U20214 ( .A(n10684), .B(n29012), .Z(n10685) );
  AND U20215 ( .A(n29013), .B(n10685), .Z(n10686) );
  OR U20216 ( .A(n29014), .B(n10686), .Z(n10687) );
  NAND U20217 ( .A(n10688), .B(n10687), .Z(n10689) );
  NANDN U20218 ( .A(n29018), .B(n10689), .Z(n10690) );
  AND U20219 ( .A(n11717), .B(n10690), .Z(n10691) );
  NANDN U20220 ( .A(x[3605]), .B(y[3605]), .Z(n23962) );
  AND U20221 ( .A(n10691), .B(n23962), .Z(n10693) );
  NANDN U20222 ( .A(y[3606]), .B(x[3606]), .Z(n10692) );
  NANDN U20223 ( .A(y[3607]), .B(x[3607]), .Z(n11714) );
  NAND U20224 ( .A(n10692), .B(n11714), .Z(n29020) );
  OR U20225 ( .A(n10693), .B(n29020), .Z(n10694) );
  AND U20226 ( .A(n11715), .B(n10694), .Z(n10695) );
  NANDN U20227 ( .A(x[3607]), .B(y[3607]), .Z(n29022) );
  AND U20228 ( .A(n10695), .B(n29022), .Z(n10697) );
  NANDN U20229 ( .A(y[3608]), .B(x[3608]), .Z(n10696) );
  NANDN U20230 ( .A(y[3609]), .B(x[3609]), .Z(n22546) );
  NAND U20231 ( .A(n10696), .B(n22546), .Z(n29023) );
  OR U20232 ( .A(n10697), .B(n29023), .Z(n10698) );
  AND U20233 ( .A(n10699), .B(n10698), .Z(n10700) );
  OR U20234 ( .A(n29026), .B(n10700), .Z(n10701) );
  NAND U20235 ( .A(n29027), .B(n10701), .Z(n10702) );
  NANDN U20236 ( .A(n29028), .B(n10702), .Z(n10703) );
  AND U20237 ( .A(n29029), .B(n10703), .Z(n10704) );
  NANDN U20238 ( .A(y[3614]), .B(x[3614]), .Z(n11709) );
  NANDN U20239 ( .A(y[3615]), .B(x[3615]), .Z(n11706) );
  NAND U20240 ( .A(n11709), .B(n11706), .Z(n29030) );
  OR U20241 ( .A(n10704), .B(n29030), .Z(n10705) );
  AND U20242 ( .A(n29031), .B(n10705), .Z(n10706) );
  OR U20243 ( .A(n29032), .B(n10706), .Z(n10707) );
  NAND U20244 ( .A(n29034), .B(n10707), .Z(n10708) );
  NANDN U20245 ( .A(n29035), .B(n10708), .Z(n10709) );
  AND U20246 ( .A(n11699), .B(n10709), .Z(n10710) );
  NANDN U20247 ( .A(x[3619]), .B(y[3619]), .Z(n29036) );
  AND U20248 ( .A(n10710), .B(n29036), .Z(n10711) );
  OR U20249 ( .A(n29037), .B(n10711), .Z(n10712) );
  AND U20250 ( .A(n10713), .B(n10712), .Z(n10714) );
  OR U20251 ( .A(n29040), .B(n10714), .Z(n10715) );
  NAND U20252 ( .A(n29041), .B(n10715), .Z(n10716) );
  NANDN U20253 ( .A(n29042), .B(n10716), .Z(n10717) );
  AND U20254 ( .A(n29043), .B(n10717), .Z(n10718) );
  NANDN U20255 ( .A(y[3626]), .B(x[3626]), .Z(n11692) );
  NANDN U20256 ( .A(y[3627]), .B(x[3627]), .Z(n11689) );
  NAND U20257 ( .A(n11692), .B(n11689), .Z(n29044) );
  OR U20258 ( .A(n10718), .B(n29044), .Z(n10719) );
  AND U20259 ( .A(n10720), .B(n10719), .Z(n10721) );
  OR U20260 ( .A(n29047), .B(n10721), .Z(n10722) );
  NAND U20261 ( .A(n29048), .B(n10722), .Z(n10723) );
  NANDN U20262 ( .A(n29049), .B(n10723), .Z(n10724) );
  AND U20263 ( .A(n22596), .B(n10724), .Z(n10725) );
  NANDN U20264 ( .A(x[3631]), .B(y[3631]), .Z(n29051) );
  AND U20265 ( .A(n10725), .B(n29051), .Z(n10727) );
  ANDN U20266 ( .B(x[3633]), .A(y[3633]), .Z(n22604) );
  NANDN U20267 ( .A(y[3632]), .B(x[3632]), .Z(n10726) );
  NANDN U20268 ( .A(n22604), .B(n10726), .Z(n29054) );
  OR U20269 ( .A(n10727), .B(n29054), .Z(n10728) );
  AND U20270 ( .A(n22602), .B(n10728), .Z(n10729) );
  NANDN U20271 ( .A(x[3633]), .B(y[3633]), .Z(n29055) );
  AND U20272 ( .A(n10729), .B(n29055), .Z(n10731) );
  NANDN U20273 ( .A(y[3634]), .B(x[3634]), .Z(n10730) );
  NANDN U20274 ( .A(y[3635]), .B(x[3635]), .Z(n11683) );
  NAND U20275 ( .A(n10730), .B(n11683), .Z(n29057) );
  OR U20276 ( .A(n10731), .B(n29057), .Z(n10732) );
  AND U20277 ( .A(n29058), .B(n10732), .Z(n10733) );
  OR U20278 ( .A(n29059), .B(n10733), .Z(n10734) );
  NAND U20279 ( .A(n29060), .B(n10734), .Z(n10735) );
  NANDN U20280 ( .A(n29061), .B(n10735), .Z(n10736) );
  AND U20281 ( .A(n29062), .B(n10736), .Z(n10737) );
  NANDN U20282 ( .A(y[3640]), .B(x[3640]), .Z(n11680) );
  NANDN U20283 ( .A(y[3641]), .B(x[3641]), .Z(n11679) );
  AND U20284 ( .A(n11680), .B(n11679), .Z(n29063) );
  NANDN U20285 ( .A(n10737), .B(n29063), .Z(n10738) );
  NANDN U20286 ( .A(n29064), .B(n10738), .Z(n10739) );
  NANDN U20287 ( .A(y[3642]), .B(x[3642]), .Z(n11678) );
  NANDN U20288 ( .A(y[3643]), .B(x[3643]), .Z(n11677) );
  AND U20289 ( .A(n11678), .B(n11677), .Z(n29065) );
  AND U20290 ( .A(n10739), .B(n29065), .Z(n10740) );
  NANDN U20291 ( .A(x[3643]), .B(y[3643]), .Z(n22629) );
  NANDN U20292 ( .A(x[3644]), .B(y[3644]), .Z(n22636) );
  NAND U20293 ( .A(n22629), .B(n22636), .Z(n23960) );
  OR U20294 ( .A(n10740), .B(n23960), .Z(n10741) );
  NAND U20295 ( .A(n23959), .B(n10741), .Z(n10742) );
  NANDN U20296 ( .A(n29066), .B(n10742), .Z(n10743) );
  NANDN U20297 ( .A(y[3646]), .B(x[3646]), .Z(n11674) );
  NANDN U20298 ( .A(y[3647]), .B(x[3647]), .Z(n11673) );
  AND U20299 ( .A(n11674), .B(n11673), .Z(n29069) );
  AND U20300 ( .A(n10743), .B(n29069), .Z(n10744) );
  NANDN U20301 ( .A(x[3647]), .B(y[3647]), .Z(n22641) );
  NANDN U20302 ( .A(x[3648]), .B(y[3648]), .Z(n11671) );
  NAND U20303 ( .A(n22641), .B(n11671), .Z(n23958) );
  OR U20304 ( .A(n10744), .B(n23958), .Z(n10745) );
  NANDN U20305 ( .A(y[3648]), .B(x[3648]), .Z(n11672) );
  NANDN U20306 ( .A(y[3649]), .B(x[3649]), .Z(n11668) );
  AND U20307 ( .A(n11672), .B(n11668), .Z(n23957) );
  AND U20308 ( .A(n10745), .B(n23957), .Z(n10746) );
  NANDN U20309 ( .A(x[3649]), .B(y[3649]), .Z(n11670) );
  NANDN U20310 ( .A(x[3650]), .B(y[3650]), .Z(n11667) );
  AND U20311 ( .A(n11670), .B(n11667), .Z(n29070) );
  NANDN U20312 ( .A(n10746), .B(n29070), .Z(n10747) );
  NANDN U20313 ( .A(n29071), .B(n10747), .Z(n10748) );
  AND U20314 ( .A(n22655), .B(n10748), .Z(n10749) );
  NANDN U20315 ( .A(x[3651]), .B(y[3651]), .Z(n23955) );
  AND U20316 ( .A(n10749), .B(n23955), .Z(n10750) );
  OR U20317 ( .A(n29072), .B(n10750), .Z(n10751) );
  NAND U20318 ( .A(n29073), .B(n10751), .Z(n10752) );
  NANDN U20319 ( .A(n29074), .B(n10752), .Z(n10753) );
  AND U20320 ( .A(n29075), .B(n10753), .Z(n10754) );
  NANDN U20321 ( .A(y[3656]), .B(x[3656]), .Z(n11663) );
  NANDN U20322 ( .A(y[3657]), .B(x[3657]), .Z(n11662) );
  AND U20323 ( .A(n11663), .B(n11662), .Z(n29076) );
  NANDN U20324 ( .A(n10754), .B(n29076), .Z(n10755) );
  NANDN U20325 ( .A(n23954), .B(n10755), .Z(n10756) );
  NANDN U20326 ( .A(y[3658]), .B(x[3658]), .Z(n11661) );
  NANDN U20327 ( .A(y[3659]), .B(x[3659]), .Z(n11660) );
  AND U20328 ( .A(n11661), .B(n11660), .Z(n29077) );
  AND U20329 ( .A(n10756), .B(n29077), .Z(n10757) );
  NANDN U20330 ( .A(x[3659]), .B(y[3659]), .Z(n22675) );
  NANDN U20331 ( .A(x[3660]), .B(y[3660]), .Z(n22682) );
  NAND U20332 ( .A(n22675), .B(n22682), .Z(n23953) );
  OR U20333 ( .A(n10757), .B(n23953), .Z(n10758) );
  NAND U20334 ( .A(n23952), .B(n10758), .Z(n10759) );
  NANDN U20335 ( .A(n29080), .B(n10759), .Z(n10760) );
  AND U20336 ( .A(n29081), .B(n10760), .Z(n10761) );
  NANDN U20337 ( .A(x[3663]), .B(y[3663]), .Z(n11657) );
  NANDN U20338 ( .A(x[3664]), .B(y[3664]), .Z(n11653) );
  AND U20339 ( .A(n11657), .B(n11653), .Z(n29082) );
  NANDN U20340 ( .A(n10761), .B(n29082), .Z(n10762) );
  NANDN U20341 ( .A(n29083), .B(n10762), .Z(n10763) );
  XOR U20342 ( .A(x[3666]), .B(y[3666]), .Z(n22695) );
  ANDN U20343 ( .B(n10763), .A(n22695), .Z(n10764) );
  NANDN U20344 ( .A(x[3665]), .B(y[3665]), .Z(n29084) );
  AND U20345 ( .A(n10764), .B(n29084), .Z(n10766) );
  NANDN U20346 ( .A(y[3666]), .B(x[3666]), .Z(n10765) );
  NANDN U20347 ( .A(y[3667]), .B(x[3667]), .Z(n11651) );
  NAND U20348 ( .A(n10765), .B(n11651), .Z(n23951) );
  OR U20349 ( .A(n10766), .B(n23951), .Z(n10767) );
  NAND U20350 ( .A(n10768), .B(n10767), .Z(n10770) );
  NANDN U20351 ( .A(y[3668]), .B(x[3668]), .Z(n10769) );
  NANDN U20352 ( .A(y[3669]), .B(x[3669]), .Z(n11649) );
  AND U20353 ( .A(n10769), .B(n11649), .Z(n29088) );
  AND U20354 ( .A(n10770), .B(n29088), .Z(n10771) );
  NOR U20355 ( .A(n22700), .B(n10771), .Z(n10772) );
  NAND U20356 ( .A(n11650), .B(n10772), .Z(n10773) );
  NANDN U20357 ( .A(n29090), .B(n10773), .Z(n10774) );
  AND U20358 ( .A(n29091), .B(n10774), .Z(n10775) );
  OR U20359 ( .A(n29092), .B(n10775), .Z(n10776) );
  AND U20360 ( .A(n10777), .B(n10776), .Z(n10778) );
  OR U20361 ( .A(n29095), .B(n10778), .Z(n10779) );
  NAND U20362 ( .A(n29096), .B(n10779), .Z(n10780) );
  NANDN U20363 ( .A(n29097), .B(n10780), .Z(n10781) );
  AND U20364 ( .A(n29098), .B(n10781), .Z(n10782) );
  NANDN U20365 ( .A(y[3678]), .B(x[3678]), .Z(n22725) );
  NANDN U20366 ( .A(y[3679]), .B(x[3679]), .Z(n22732) );
  NAND U20367 ( .A(n22725), .B(n22732), .Z(n29099) );
  OR U20368 ( .A(n10782), .B(n29099), .Z(n10783) );
  AND U20369 ( .A(n29100), .B(n10783), .Z(n10784) );
  OR U20370 ( .A(n29101), .B(n10784), .Z(n10785) );
  NAND U20371 ( .A(n10786), .B(n10785), .Z(n10787) );
  NANDN U20372 ( .A(n29102), .B(n10787), .Z(n10788) );
  AND U20373 ( .A(n22743), .B(n10788), .Z(n10789) );
  NAND U20374 ( .A(n29103), .B(n10789), .Z(n10790) );
  NANDN U20375 ( .A(n29105), .B(n10790), .Z(n10791) );
  NANDN U20376 ( .A(x[3685]), .B(y[3685]), .Z(n22746) );
  NANDN U20377 ( .A(x[3686]), .B(y[3686]), .Z(n11637) );
  AND U20378 ( .A(n22746), .B(n11637), .Z(n29108) );
  AND U20379 ( .A(n10791), .B(n29108), .Z(n10792) );
  NANDN U20380 ( .A(y[3686]), .B(x[3686]), .Z(n11638) );
  NANDN U20381 ( .A(y[3687]), .B(x[3687]), .Z(n11635) );
  NAND U20382 ( .A(n11638), .B(n11635), .Z(n23946) );
  OR U20383 ( .A(n10792), .B(n23946), .Z(n10793) );
  NAND U20384 ( .A(n23945), .B(n10793), .Z(n10794) );
  NANDN U20385 ( .A(n29109), .B(n10794), .Z(n10795) );
  AND U20386 ( .A(n29110), .B(n10795), .Z(n10796) );
  NANDN U20387 ( .A(y[3690]), .B(x[3690]), .Z(n11632) );
  NANDN U20388 ( .A(y[3691]), .B(x[3691]), .Z(n11631) );
  NAND U20389 ( .A(n11632), .B(n11631), .Z(n29111) );
  OR U20390 ( .A(n10796), .B(n29111), .Z(n10797) );
  AND U20391 ( .A(n29112), .B(n10797), .Z(n10798) );
  NANDN U20392 ( .A(y[3692]), .B(x[3692]), .Z(n11630) );
  NANDN U20393 ( .A(y[3693]), .B(x[3693]), .Z(n11629) );
  NAND U20394 ( .A(n11630), .B(n11629), .Z(n23944) );
  OR U20395 ( .A(n10798), .B(n23944), .Z(n10799) );
  NAND U20396 ( .A(n29113), .B(n10799), .Z(n10800) );
  NAND U20397 ( .A(n29114), .B(n10800), .Z(n10801) );
  AND U20398 ( .A(n22776), .B(n10801), .Z(n10802) );
  NANDN U20399 ( .A(x[3695]), .B(y[3695]), .Z(n29116) );
  AND U20400 ( .A(n10802), .B(n29116), .Z(n10804) );
  NANDN U20401 ( .A(y[3696]), .B(x[3696]), .Z(n10803) );
  NANDN U20402 ( .A(y[3697]), .B(x[3697]), .Z(n22782) );
  NAND U20403 ( .A(n10803), .B(n22782), .Z(n29117) );
  OR U20404 ( .A(n10804), .B(n29117), .Z(n10805) );
  AND U20405 ( .A(n29119), .B(n10805), .Z(n10806) );
  OR U20406 ( .A(n29120), .B(n10806), .Z(n10807) );
  NAND U20407 ( .A(n29121), .B(n10807), .Z(n10808) );
  NANDN U20408 ( .A(n29122), .B(n10808), .Z(n10809) );
  AND U20409 ( .A(n29123), .B(n10809), .Z(n10810) );
  NANDN U20410 ( .A(y[3702]), .B(x[3702]), .Z(n22793) );
  NANDN U20411 ( .A(y[3703]), .B(x[3703]), .Z(n22799) );
  AND U20412 ( .A(n22793), .B(n22799), .Z(n23943) );
  NANDN U20413 ( .A(n10810), .B(n23943), .Z(n10811) );
  NAND U20414 ( .A(n10812), .B(n10811), .Z(n10814) );
  NANDN U20415 ( .A(y[3704]), .B(x[3704]), .Z(n10813) );
  NANDN U20416 ( .A(y[3705]), .B(x[3705]), .Z(n22806) );
  AND U20417 ( .A(n10813), .B(n22806), .Z(n29126) );
  AND U20418 ( .A(n10814), .B(n29126), .Z(n10815) );
  NANDN U20419 ( .A(x[3705]), .B(y[3705]), .Z(n11619) );
  NANDN U20420 ( .A(x[3706]), .B(y[3706]), .Z(n11618) );
  AND U20421 ( .A(n11619), .B(n11618), .Z(n29127) );
  NANDN U20422 ( .A(n10815), .B(n29127), .Z(n10816) );
  NANDN U20423 ( .A(n29128), .B(n10816), .Z(n10817) );
  AND U20424 ( .A(n29129), .B(n10817), .Z(n10818) );
  OR U20425 ( .A(n29130), .B(n10818), .Z(n10819) );
  NAND U20426 ( .A(n29131), .B(n10819), .Z(n10820) );
  NANDN U20427 ( .A(n29132), .B(n10820), .Z(n10821) );
  NANDN U20428 ( .A(x[3711]), .B(y[3711]), .Z(n11613) );
  NANDN U20429 ( .A(x[3712]), .B(y[3712]), .Z(n11612) );
  AND U20430 ( .A(n11613), .B(n11612), .Z(n23942) );
  AND U20431 ( .A(n10821), .B(n23942), .Z(n10822) );
  ANDN U20432 ( .B(x[3713]), .A(y[3713]), .Z(n22830) );
  NANDN U20433 ( .A(y[3712]), .B(x[3712]), .Z(n22823) );
  NANDN U20434 ( .A(n22830), .B(n22823), .Z(n29133) );
  OR U20435 ( .A(n10822), .B(n29133), .Z(n10823) );
  NANDN U20436 ( .A(x[3713]), .B(y[3713]), .Z(n11611) );
  NANDN U20437 ( .A(x[3714]), .B(y[3714]), .Z(n11610) );
  AND U20438 ( .A(n11611), .B(n11610), .Z(n29136) );
  AND U20439 ( .A(n10823), .B(n29136), .Z(n10824) );
  NANDN U20440 ( .A(y[3714]), .B(x[3714]), .Z(n22832) );
  NANDN U20441 ( .A(y[3715]), .B(x[3715]), .Z(n11608) );
  NAND U20442 ( .A(n22832), .B(n11608), .Z(n23941) );
  OR U20443 ( .A(n10824), .B(n23941), .Z(n10825) );
  NAND U20444 ( .A(n23940), .B(n10825), .Z(n10826) );
  NANDN U20445 ( .A(n29137), .B(n10826), .Z(n10827) );
  AND U20446 ( .A(n29138), .B(n10827), .Z(n10828) );
  NANDN U20447 ( .A(y[3718]), .B(x[3718]), .Z(n22840) );
  NANDN U20448 ( .A(y[3719]), .B(x[3719]), .Z(n22847) );
  NAND U20449 ( .A(n22840), .B(n22847), .Z(n29139) );
  OR U20450 ( .A(n10828), .B(n29139), .Z(n10829) );
  AND U20451 ( .A(n10830), .B(n10829), .Z(n10832) );
  NANDN U20452 ( .A(y[3720]), .B(x[3720]), .Z(n10831) );
  NANDN U20453 ( .A(y[3721]), .B(x[3721]), .Z(n11602) );
  NAND U20454 ( .A(n10831), .B(n11602), .Z(n29142) );
  OR U20455 ( .A(n10832), .B(n29142), .Z(n10833) );
  NAND U20456 ( .A(n29143), .B(n10833), .Z(n10834) );
  NANDN U20457 ( .A(n29144), .B(n10834), .Z(n10835) );
  AND U20458 ( .A(n29145), .B(n10835), .Z(n10836) );
  NANDN U20459 ( .A(y[3724]), .B(x[3724]), .Z(n11598) );
  NANDN U20460 ( .A(y[3725]), .B(x[3725]), .Z(n22859) );
  NAND U20461 ( .A(n11598), .B(n22859), .Z(n29146) );
  OR U20462 ( .A(n10836), .B(n29146), .Z(n10837) );
  AND U20463 ( .A(n10838), .B(n10837), .Z(n10839) );
  OR U20464 ( .A(n29150), .B(n10839), .Z(n10840) );
  NAND U20465 ( .A(n29151), .B(n10840), .Z(n10841) );
  NANDN U20466 ( .A(n29152), .B(n10841), .Z(n10842) );
  AND U20467 ( .A(n29153), .B(n10842), .Z(n10843) );
  NANDN U20468 ( .A(y[3730]), .B(x[3730]), .Z(n11590) );
  NANDN U20469 ( .A(y[3731]), .B(x[3731]), .Z(n11589) );
  NAND U20470 ( .A(n11590), .B(n11589), .Z(n29154) );
  OR U20471 ( .A(n10843), .B(n29154), .Z(n10844) );
  AND U20472 ( .A(n29155), .B(n10844), .Z(n10845) );
  OR U20473 ( .A(n29156), .B(n10845), .Z(n10846) );
  NAND U20474 ( .A(n29157), .B(n10846), .Z(n10847) );
  NANDN U20475 ( .A(n29158), .B(n10847), .Z(n10848) );
  AND U20476 ( .A(n29159), .B(n10848), .Z(n10849) );
  NANDN U20477 ( .A(y[3736]), .B(x[3736]), .Z(n11584) );
  NANDN U20478 ( .A(y[3737]), .B(x[3737]), .Z(n22895) );
  AND U20479 ( .A(n11584), .B(n22895), .Z(n23939) );
  NANDN U20480 ( .A(n10849), .B(n23939), .Z(n10850) );
  NANDN U20481 ( .A(n29160), .B(n10850), .Z(n10851) );
  AND U20482 ( .A(n29161), .B(n10851), .Z(n10852) );
  OR U20483 ( .A(n29162), .B(n10852), .Z(n10853) );
  NAND U20484 ( .A(n29163), .B(n10853), .Z(n10854) );
  NANDN U20485 ( .A(n29164), .B(n10854), .Z(n10855) );
  AND U20486 ( .A(n29165), .B(n10855), .Z(n10856) );
  NANDN U20487 ( .A(x[3743]), .B(y[3743]), .Z(n11578) );
  NANDN U20488 ( .A(x[3744]), .B(y[3744]), .Z(n11575) );
  AND U20489 ( .A(n11578), .B(n11575), .Z(n23938) );
  NANDN U20490 ( .A(n10856), .B(n23938), .Z(n10857) );
  NAND U20491 ( .A(n29167), .B(n10857), .Z(n10858) );
  AND U20492 ( .A(n11574), .B(n10858), .Z(n10859) );
  NANDN U20493 ( .A(x[3745]), .B(y[3745]), .Z(n29169) );
  AND U20494 ( .A(n10859), .B(n29169), .Z(n10861) );
  NANDN U20495 ( .A(y[3746]), .B(x[3746]), .Z(n10860) );
  NANDN U20496 ( .A(y[3747]), .B(x[3747]), .Z(n22923) );
  NAND U20497 ( .A(n10860), .B(n22923), .Z(n29170) );
  OR U20498 ( .A(n10861), .B(n29170), .Z(n10862) );
  NAND U20499 ( .A(n29171), .B(n10862), .Z(n10863) );
  NANDN U20500 ( .A(y[3748]), .B(x[3748]), .Z(n22922) );
  NANDN U20501 ( .A(y[3749]), .B(x[3749]), .Z(n22929) );
  AND U20502 ( .A(n22922), .B(n22929), .Z(n29172) );
  AND U20503 ( .A(n10863), .B(n29172), .Z(n10865) );
  XNOR U20504 ( .A(x[3750]), .B(y[3750]), .Z(n22928) );
  ANDN U20505 ( .B(y[3749]), .A(x[3749]), .Z(n11571) );
  ANDN U20506 ( .B(n22928), .A(n11571), .Z(n10864) );
  NANDN U20507 ( .A(n10865), .B(n10864), .Z(n10867) );
  NANDN U20508 ( .A(y[3750]), .B(x[3750]), .Z(n10866) );
  NANDN U20509 ( .A(y[3751]), .B(x[3751]), .Z(n22935) );
  AND U20510 ( .A(n10866), .B(n22935), .Z(n29173) );
  AND U20511 ( .A(n10867), .B(n29173), .Z(n10868) );
  NANDN U20512 ( .A(x[3751]), .B(y[3751]), .Z(n11570) );
  NANDN U20513 ( .A(x[3752]), .B(y[3752]), .Z(n22938) );
  NAND U20514 ( .A(n11570), .B(n22938), .Z(n23935) );
  OR U20515 ( .A(n10868), .B(n23935), .Z(n10869) );
  NAND U20516 ( .A(n23934), .B(n10869), .Z(n10870) );
  NANDN U20517 ( .A(n29174), .B(n10870), .Z(n10871) );
  NANDN U20518 ( .A(y[3754]), .B(x[3754]), .Z(n11568) );
  NANDN U20519 ( .A(y[3755]), .B(x[3755]), .Z(n11567) );
  AND U20520 ( .A(n11568), .B(n11567), .Z(n29175) );
  AND U20521 ( .A(n10871), .B(n29175), .Z(n10872) );
  NANDN U20522 ( .A(x[3755]), .B(y[3755]), .Z(n22943) );
  NANDN U20523 ( .A(x[3756]), .B(y[3756]), .Z(n22950) );
  NAND U20524 ( .A(n22943), .B(n22950), .Z(n29178) );
  OR U20525 ( .A(n10872), .B(n29178), .Z(n10873) );
  NANDN U20526 ( .A(y[3756]), .B(x[3756]), .Z(n11566) );
  NANDN U20527 ( .A(y[3757]), .B(x[3757]), .Z(n11565) );
  AND U20528 ( .A(n11566), .B(n11565), .Z(n29179) );
  AND U20529 ( .A(n10873), .B(n29179), .Z(n10874) );
  NANDN U20530 ( .A(x[3757]), .B(y[3757]), .Z(n22949) );
  NANDN U20531 ( .A(x[3758]), .B(y[3758]), .Z(n22956) );
  NAND U20532 ( .A(n22949), .B(n22956), .Z(n23933) );
  OR U20533 ( .A(n10874), .B(n23933), .Z(n10875) );
  NAND U20534 ( .A(n23932), .B(n10875), .Z(n10876) );
  NANDN U20535 ( .A(n29180), .B(n10876), .Z(n10877) );
  AND U20536 ( .A(n29181), .B(n10877), .Z(n10878) );
  NANDN U20537 ( .A(x[3761]), .B(y[3761]), .Z(n22961) );
  NANDN U20538 ( .A(x[3762]), .B(y[3762]), .Z(n22968) );
  AND U20539 ( .A(n22961), .B(n22968), .Z(n23931) );
  NANDN U20540 ( .A(n10878), .B(n23931), .Z(n10879) );
  NANDN U20541 ( .A(n29182), .B(n10879), .Z(n10880) );
  NANDN U20542 ( .A(x[3763]), .B(y[3763]), .Z(n22967) );
  NANDN U20543 ( .A(x[3764]), .B(y[3764]), .Z(n22974) );
  AND U20544 ( .A(n22967), .B(n22974), .Z(n29183) );
  AND U20545 ( .A(n10880), .B(n29183), .Z(n10881) );
  NANDN U20546 ( .A(y[3764]), .B(x[3764]), .Z(n11558) );
  NANDN U20547 ( .A(y[3765]), .B(x[3765]), .Z(n11557) );
  NAND U20548 ( .A(n11558), .B(n11557), .Z(n23930) );
  OR U20549 ( .A(n10881), .B(n23930), .Z(n10882) );
  NAND U20550 ( .A(n23929), .B(n10882), .Z(n10883) );
  NANDN U20551 ( .A(n29186), .B(n10883), .Z(n10884) );
  AND U20552 ( .A(n11553), .B(n10884), .Z(n10885) );
  NANDN U20553 ( .A(x[3767]), .B(y[3767]), .Z(n29188) );
  NAND U20554 ( .A(n10885), .B(n29188), .Z(n10886) );
  NANDN U20555 ( .A(n29190), .B(n10886), .Z(n10887) );
  NANDN U20556 ( .A(x[3769]), .B(y[3769]), .Z(n22983) );
  NANDN U20557 ( .A(x[3770]), .B(y[3770]), .Z(n11550) );
  AND U20558 ( .A(n22983), .B(n11550), .Z(n29191) );
  AND U20559 ( .A(n10887), .B(n29191), .Z(n10888) );
  NANDN U20560 ( .A(y[3770]), .B(x[3770]), .Z(n11551) );
  NANDN U20561 ( .A(y[3771]), .B(x[3771]), .Z(n11548) );
  NAND U20562 ( .A(n11551), .B(n11548), .Z(n23928) );
  OR U20563 ( .A(n10888), .B(n23928), .Z(n10889) );
  NAND U20564 ( .A(n23927), .B(n10889), .Z(n10890) );
  NANDN U20565 ( .A(n29192), .B(n10890), .Z(n10891) );
  NANDN U20566 ( .A(x[3773]), .B(y[3773]), .Z(n22993) );
  NANDN U20567 ( .A(x[3774]), .B(y[3774]), .Z(n23000) );
  AND U20568 ( .A(n22993), .B(n23000), .Z(n29193) );
  AND U20569 ( .A(n10891), .B(n29193), .Z(n10892) );
  NANDN U20570 ( .A(y[3774]), .B(x[3774]), .Z(n11545) );
  NANDN U20571 ( .A(y[3775]), .B(x[3775]), .Z(n11544) );
  NAND U20572 ( .A(n11545), .B(n11544), .Z(n29194) );
  OR U20573 ( .A(n10892), .B(n29194), .Z(n10893) );
  NANDN U20574 ( .A(x[3775]), .B(y[3775]), .Z(n22999) );
  NANDN U20575 ( .A(x[3776]), .B(y[3776]), .Z(n23006) );
  AND U20576 ( .A(n22999), .B(n23006), .Z(n29195) );
  AND U20577 ( .A(n10893), .B(n29195), .Z(n10894) );
  NANDN U20578 ( .A(y[3776]), .B(x[3776]), .Z(n11543) );
  NANDN U20579 ( .A(y[3777]), .B(x[3777]), .Z(n23009) );
  NAND U20580 ( .A(n11543), .B(n23009), .Z(n23926) );
  OR U20581 ( .A(n10894), .B(n23926), .Z(n10895) );
  NAND U20582 ( .A(n23925), .B(n10895), .Z(n10896) );
  NAND U20583 ( .A(n29197), .B(n10896), .Z(n10897) );
  AND U20584 ( .A(n23015), .B(n10897), .Z(n10898) );
  NANDN U20585 ( .A(x[3779]), .B(y[3779]), .Z(n29199) );
  AND U20586 ( .A(n10898), .B(n29199), .Z(n10900) );
  NANDN U20587 ( .A(y[3780]), .B(x[3780]), .Z(n10899) );
  NANDN U20588 ( .A(y[3781]), .B(x[3781]), .Z(n23021) );
  NAND U20589 ( .A(n10899), .B(n23021), .Z(n29200) );
  OR U20590 ( .A(n10900), .B(n29200), .Z(n10901) );
  AND U20591 ( .A(n29201), .B(n10901), .Z(n10902) );
  OR U20592 ( .A(n29202), .B(n10902), .Z(n10903) );
  NAND U20593 ( .A(n29203), .B(n10903), .Z(n10904) );
  NANDN U20594 ( .A(n29204), .B(n10904), .Z(n10905) );
  AND U20595 ( .A(n29205), .B(n10905), .Z(n10906) );
  NANDN U20596 ( .A(y[3786]), .B(x[3786]), .Z(n23035) );
  NANDN U20597 ( .A(y[3787]), .B(x[3787]), .Z(n23042) );
  NAND U20598 ( .A(n23035), .B(n23042), .Z(n29206) );
  OR U20599 ( .A(n10906), .B(n29206), .Z(n10907) );
  AND U20600 ( .A(n10908), .B(n10907), .Z(n10909) );
  OR U20601 ( .A(n29209), .B(n10909), .Z(n10910) );
  NAND U20602 ( .A(n29210), .B(n10910), .Z(n10911) );
  NANDN U20603 ( .A(n29211), .B(n10911), .Z(n10912) );
  AND U20604 ( .A(n11535), .B(n10912), .Z(n10913) );
  NANDN U20605 ( .A(x[3791]), .B(y[3791]), .Z(n29212) );
  AND U20606 ( .A(n10913), .B(n29212), .Z(n10914) );
  OR U20607 ( .A(n29216), .B(n10914), .Z(n10915) );
  AND U20608 ( .A(n10916), .B(n10915), .Z(n10917) );
  OR U20609 ( .A(n29218), .B(n10917), .Z(n10918) );
  NAND U20610 ( .A(n29219), .B(n10918), .Z(n10919) );
  NANDN U20611 ( .A(n29220), .B(n10919), .Z(n10920) );
  AND U20612 ( .A(n29221), .B(n10920), .Z(n10921) );
  NANDN U20613 ( .A(y[3798]), .B(x[3798]), .Z(n11528) );
  NANDN U20614 ( .A(y[3799]), .B(x[3799]), .Z(n23074) );
  NAND U20615 ( .A(n11528), .B(n23074), .Z(n29222) );
  OR U20616 ( .A(n10921), .B(n29222), .Z(n10922) );
  AND U20617 ( .A(n29223), .B(n10922), .Z(n10923) );
  OR U20618 ( .A(n29224), .B(n10923), .Z(n10924) );
  NAND U20619 ( .A(n29225), .B(n10924), .Z(n10925) );
  NANDN U20620 ( .A(n29226), .B(n10925), .Z(n10926) );
  AND U20621 ( .A(n29227), .B(n10926), .Z(n10927) );
  NANDN U20622 ( .A(y[3804]), .B(x[3804]), .Z(n23085) );
  NANDN U20623 ( .A(y[3805]), .B(x[3805]), .Z(n11521) );
  NAND U20624 ( .A(n23085), .B(n11521), .Z(n29228) );
  OR U20625 ( .A(n10927), .B(n29228), .Z(n10928) );
  NAND U20626 ( .A(n10929), .B(n10928), .Z(n10931) );
  NANDN U20627 ( .A(y[3806]), .B(x[3806]), .Z(n10930) );
  NANDN U20628 ( .A(y[3807]), .B(x[3807]), .Z(n11518) );
  AND U20629 ( .A(n10930), .B(n11518), .Z(n29231) );
  AND U20630 ( .A(n10931), .B(n29231), .Z(n10932) );
  NOR U20631 ( .A(n11520), .B(n10932), .Z(n10933) );
  NAND U20632 ( .A(n11519), .B(n10933), .Z(n10934) );
  NANDN U20633 ( .A(n23921), .B(n10934), .Z(n10935) );
  AND U20634 ( .A(n23100), .B(n10935), .Z(n10936) );
  ANDN U20635 ( .B(y[3809]), .A(x[3809]), .Z(n29235) );
  ANDN U20636 ( .B(n10936), .A(n29235), .Z(n10938) );
  ANDN U20637 ( .B(x[3811]), .A(y[3811]), .Z(n23108) );
  NANDN U20638 ( .A(y[3810]), .B(x[3810]), .Z(n10937) );
  NANDN U20639 ( .A(n23108), .B(n10937), .Z(n29236) );
  OR U20640 ( .A(n10938), .B(n29236), .Z(n10939) );
  AND U20641 ( .A(n29237), .B(n10939), .Z(n10940) );
  NAND U20642 ( .A(n23106), .B(n10940), .Z(n10941) );
  NANDN U20643 ( .A(n29239), .B(n10941), .Z(n10942) );
  AND U20644 ( .A(n10943), .B(n10942), .Z(n10944) );
  OR U20645 ( .A(n29242), .B(n10944), .Z(n10945) );
  NAND U20646 ( .A(n29243), .B(n10945), .Z(n10946) );
  NANDN U20647 ( .A(n29244), .B(n10946), .Z(n10947) );
  AND U20648 ( .A(n11513), .B(n10947), .Z(n10948) );
  NANDN U20649 ( .A(x[3817]), .B(y[3817]), .Z(n29245) );
  AND U20650 ( .A(n10948), .B(n29245), .Z(n10949) );
  OR U20651 ( .A(n29247), .B(n10949), .Z(n10950) );
  AND U20652 ( .A(n10951), .B(n10950), .Z(n10952) );
  OR U20653 ( .A(n29250), .B(n10952), .Z(n10953) );
  NAND U20654 ( .A(n29252), .B(n10953), .Z(n10954) );
  NANDN U20655 ( .A(n29253), .B(n10954), .Z(n10955) );
  AND U20656 ( .A(n29254), .B(n10955), .Z(n10956) );
  NANDN U20657 ( .A(y[3824]), .B(x[3824]), .Z(n23135) );
  NANDN U20658 ( .A(y[3825]), .B(x[3825]), .Z(n11504) );
  NAND U20659 ( .A(n23135), .B(n11504), .Z(n29255) );
  OR U20660 ( .A(n10956), .B(n29255), .Z(n10957) );
  AND U20661 ( .A(n29256), .B(n10957), .Z(n10958) );
  OR U20662 ( .A(n29257), .B(n10958), .Z(n10959) );
  NAND U20663 ( .A(n10960), .B(n10959), .Z(n10961) );
  NAND U20664 ( .A(n29258), .B(n10961), .Z(n10962) );
  AND U20665 ( .A(n23150), .B(n10962), .Z(n10963) );
  ANDN U20666 ( .B(y[3829]), .A(x[3829]), .Z(n29260) );
  ANDN U20667 ( .B(n10963), .A(n29260), .Z(n10965) );
  ANDN U20668 ( .B(x[3831]), .A(y[3831]), .Z(n23158) );
  NANDN U20669 ( .A(y[3830]), .B(x[3830]), .Z(n10964) );
  NANDN U20670 ( .A(n23158), .B(n10964), .Z(n29261) );
  OR U20671 ( .A(n10965), .B(n29261), .Z(n10966) );
  AND U20672 ( .A(n23156), .B(n10966), .Z(n10967) );
  NANDN U20673 ( .A(x[3831]), .B(y[3831]), .Z(n29262) );
  AND U20674 ( .A(n10967), .B(n29262), .Z(n10969) );
  NANDN U20675 ( .A(y[3832]), .B(x[3832]), .Z(n10968) );
  NANDN U20676 ( .A(y[3833]), .B(x[3833]), .Z(n11498) );
  NAND U20677 ( .A(n10968), .B(n11498), .Z(n23917) );
  OR U20678 ( .A(n10969), .B(n23917), .Z(n10970) );
  NANDN U20679 ( .A(x[3833]), .B(y[3833]), .Z(n11499) );
  NANDN U20680 ( .A(x[3834]), .B(y[3834]), .Z(n11496) );
  AND U20681 ( .A(n11499), .B(n11496), .Z(n23916) );
  AND U20682 ( .A(n10970), .B(n23916), .Z(n10971) );
  NANDN U20683 ( .A(y[3834]), .B(x[3834]), .Z(n11497) );
  NANDN U20684 ( .A(y[3835]), .B(x[3835]), .Z(n23165) );
  NAND U20685 ( .A(n11497), .B(n23165), .Z(n29263) );
  OR U20686 ( .A(n10971), .B(n29263), .Z(n10972) );
  NAND U20687 ( .A(n10973), .B(n10972), .Z(n10974) );
  NANDN U20688 ( .A(n29269), .B(n10974), .Z(n10975) );
  NANDN U20689 ( .A(x[3837]), .B(y[3837]), .Z(n23169) );
  NANDN U20690 ( .A(x[3838]), .B(y[3838]), .Z(n11493) );
  AND U20691 ( .A(n23169), .B(n11493), .Z(n29270) );
  AND U20692 ( .A(n10975), .B(n29270), .Z(n10976) );
  NANDN U20693 ( .A(y[3838]), .B(x[3838]), .Z(n11494) );
  NANDN U20694 ( .A(y[3839]), .B(x[3839]), .Z(n11491) );
  NAND U20695 ( .A(n11494), .B(n11491), .Z(n23915) );
  OR U20696 ( .A(n10976), .B(n23915), .Z(n10977) );
  NANDN U20697 ( .A(x[3839]), .B(y[3839]), .Z(n11492) );
  NANDN U20698 ( .A(x[3840]), .B(y[3840]), .Z(n23180) );
  AND U20699 ( .A(n11492), .B(n23180), .Z(n23914) );
  AND U20700 ( .A(n10977), .B(n23914), .Z(n10978) );
  NANDN U20701 ( .A(y[3840]), .B(x[3840]), .Z(n11490) );
  NANDN U20702 ( .A(y[3841]), .B(x[3841]), .Z(n11489) );
  NAND U20703 ( .A(n11490), .B(n11489), .Z(n23913) );
  OR U20704 ( .A(n10978), .B(n23913), .Z(n10979) );
  NAND U20705 ( .A(n29271), .B(n10979), .Z(n10980) );
  NANDN U20706 ( .A(n29272), .B(n10980), .Z(n10981) );
  AND U20707 ( .A(n11487), .B(n10981), .Z(n10982) );
  NANDN U20708 ( .A(x[3843]), .B(y[3843]), .Z(n29273) );
  AND U20709 ( .A(n10982), .B(n29273), .Z(n10983) );
  OR U20710 ( .A(n29275), .B(n10983), .Z(n10984) );
  AND U20711 ( .A(n10985), .B(n10984), .Z(n10986) );
  OR U20712 ( .A(n29276), .B(n10986), .Z(n10987) );
  NAND U20713 ( .A(n29278), .B(n10987), .Z(n10988) );
  NANDN U20714 ( .A(n29279), .B(n10988), .Z(n10989) );
  AND U20715 ( .A(n11481), .B(n10989), .Z(n10990) );
  NANDN U20716 ( .A(x[3849]), .B(y[3849]), .Z(n29280) );
  AND U20717 ( .A(n10990), .B(n29280), .Z(n10991) );
  OR U20718 ( .A(n29282), .B(n10991), .Z(n10992) );
  AND U20719 ( .A(n10993), .B(n10992), .Z(n10994) );
  OR U20720 ( .A(n29283), .B(n10994), .Z(n10995) );
  NAND U20721 ( .A(n29284), .B(n10995), .Z(n10996) );
  NANDN U20722 ( .A(n29285), .B(n10996), .Z(n10997) );
  AND U20723 ( .A(n29286), .B(n10997), .Z(n10998) );
  OR U20724 ( .A(n29287), .B(n10998), .Z(n10999) );
  AND U20725 ( .A(n11000), .B(n10999), .Z(n11001) );
  OR U20726 ( .A(n29288), .B(n11001), .Z(n11002) );
  NAND U20727 ( .A(n29289), .B(n11002), .Z(n11003) );
  NANDN U20728 ( .A(n29290), .B(n11003), .Z(n11004) );
  AND U20729 ( .A(n29291), .B(n11004), .Z(n11005) );
  NANDN U20730 ( .A(y[3862]), .B(x[3862]), .Z(n23234) );
  NANDN U20731 ( .A(y[3863]), .B(x[3863]), .Z(n11471) );
  NAND U20732 ( .A(n23234), .B(n11471), .Z(n29292) );
  OR U20733 ( .A(n11005), .B(n29292), .Z(n11006) );
  AND U20734 ( .A(n29294), .B(n11006), .Z(n11007) );
  NANDN U20735 ( .A(y[3864]), .B(x[3864]), .Z(n11470) );
  NANDN U20736 ( .A(y[3865]), .B(x[3865]), .Z(n11469) );
  NAND U20737 ( .A(n11470), .B(n11469), .Z(n29295) );
  OR U20738 ( .A(n11007), .B(n29295), .Z(n11008) );
  NAND U20739 ( .A(n29296), .B(n11008), .Z(n11009) );
  NANDN U20740 ( .A(n23906), .B(n11009), .Z(n11010) );
  NAND U20741 ( .A(n29297), .B(n11010), .Z(n11011) );
  NAND U20742 ( .A(n29298), .B(n11011), .Z(n11012) );
  NANDN U20743 ( .A(n29299), .B(n11012), .Z(n11013) );
  AND U20744 ( .A(n29300), .B(n11013), .Z(n11014) );
  OR U20745 ( .A(n29301), .B(n11014), .Z(n11015) );
  NAND U20746 ( .A(n29302), .B(n11015), .Z(n11016) );
  NANDN U20747 ( .A(n29303), .B(n11016), .Z(n11017) );
  AND U20748 ( .A(n29304), .B(n11017), .Z(n11018) );
  NANDN U20749 ( .A(x[3875]), .B(y[3875]), .Z(n11456) );
  NANDN U20750 ( .A(x[3876]), .B(y[3876]), .Z(n11453) );
  AND U20751 ( .A(n11456), .B(n11453), .Z(n23905) );
  NANDN U20752 ( .A(n11018), .B(n23905), .Z(n11019) );
  NAND U20753 ( .A(n29305), .B(n11019), .Z(n11020) );
  AND U20754 ( .A(n23280), .B(n11020), .Z(n11021) );
  NANDN U20755 ( .A(x[3877]), .B(y[3877]), .Z(n29308) );
  AND U20756 ( .A(n11021), .B(n29308), .Z(n11023) );
  NANDN U20757 ( .A(y[3878]), .B(x[3878]), .Z(n11022) );
  NANDN U20758 ( .A(y[3879]), .B(x[3879]), .Z(n11451) );
  NAND U20759 ( .A(n11022), .B(n11451), .Z(n29309) );
  OR U20760 ( .A(n11023), .B(n29309), .Z(n11024) );
  NAND U20761 ( .A(n29310), .B(n11024), .Z(n11025) );
  NANDN U20762 ( .A(y[3880]), .B(x[3880]), .Z(n11452) );
  NANDN U20763 ( .A(y[3881]), .B(x[3881]), .Z(n11447) );
  AND U20764 ( .A(n11452), .B(n11447), .Z(n29311) );
  AND U20765 ( .A(n11025), .B(n29311), .Z(n11027) );
  XNOR U20766 ( .A(x[3882]), .B(y[3882]), .Z(n11448) );
  ANDN U20767 ( .B(y[3881]), .A(x[3881]), .Z(n11449) );
  ANDN U20768 ( .B(n11448), .A(n11449), .Z(n11026) );
  NANDN U20769 ( .A(n11027), .B(n11026), .Z(n11029) );
  NANDN U20770 ( .A(y[3882]), .B(x[3882]), .Z(n11028) );
  NANDN U20771 ( .A(y[3883]), .B(x[3883]), .Z(n11446) );
  AND U20772 ( .A(n11028), .B(n11446), .Z(n29312) );
  AND U20773 ( .A(n11029), .B(n29312), .Z(n11030) );
  NANDN U20774 ( .A(x[3883]), .B(y[3883]), .Z(n23292) );
  NANDN U20775 ( .A(x[3884]), .B(y[3884]), .Z(n23298) );
  NAND U20776 ( .A(n23292), .B(n23298), .Z(n23902) );
  OR U20777 ( .A(n11030), .B(n23902), .Z(n11031) );
  NAND U20778 ( .A(n23901), .B(n11031), .Z(n11032) );
  NANDN U20779 ( .A(n29313), .B(n11032), .Z(n11033) );
  NANDN U20780 ( .A(y[3886]), .B(x[3886]), .Z(n11443) );
  NANDN U20781 ( .A(y[3887]), .B(x[3887]), .Z(n11442) );
  AND U20782 ( .A(n11443), .B(n11442), .Z(n29314) );
  AND U20783 ( .A(n11033), .B(n29314), .Z(n11034) );
  NANDN U20784 ( .A(x[3887]), .B(y[3887]), .Z(n23303) );
  NANDN U20785 ( .A(x[3888]), .B(y[3888]), .Z(n23309) );
  AND U20786 ( .A(n23303), .B(n23309), .Z(n29315) );
  NANDN U20787 ( .A(n11034), .B(n29315), .Z(n11035) );
  NANDN U20788 ( .A(n29316), .B(n11035), .Z(n11036) );
  AND U20789 ( .A(n23312), .B(n11036), .Z(n11037) );
  NANDN U20790 ( .A(x[3889]), .B(y[3889]), .Z(n29317) );
  AND U20791 ( .A(n11037), .B(n29317), .Z(n11039) );
  NANDN U20792 ( .A(y[3890]), .B(x[3890]), .Z(n11038) );
  NANDN U20793 ( .A(y[3891]), .B(x[3891]), .Z(n11439) );
  NAND U20794 ( .A(n11038), .B(n11439), .Z(n29321) );
  OR U20795 ( .A(n11039), .B(n29321), .Z(n11040) );
  NANDN U20796 ( .A(x[3891]), .B(y[3891]), .Z(n11440) );
  NANDN U20797 ( .A(x[3892]), .B(y[3892]), .Z(n11436) );
  AND U20798 ( .A(n11440), .B(n11436), .Z(n29322) );
  AND U20799 ( .A(n11040), .B(n29322), .Z(n11041) );
  NANDN U20800 ( .A(y[3892]), .B(x[3892]), .Z(n11438) );
  NANDN U20801 ( .A(y[3893]), .B(x[3893]), .Z(n11435) );
  NAND U20802 ( .A(n11438), .B(n11435), .Z(n23900) );
  OR U20803 ( .A(n11041), .B(n23900), .Z(n11042) );
  NAND U20804 ( .A(n23899), .B(n11042), .Z(n11043) );
  NAND U20805 ( .A(n29323), .B(n11043), .Z(n11044) );
  AND U20806 ( .A(n23326), .B(n11044), .Z(n11045) );
  NANDN U20807 ( .A(x[3895]), .B(y[3895]), .Z(n29325) );
  AND U20808 ( .A(n11045), .B(n29325), .Z(n11046) );
  OR U20809 ( .A(n29326), .B(n11046), .Z(n11047) );
  AND U20810 ( .A(n11048), .B(n11047), .Z(n11049) );
  OR U20811 ( .A(n29328), .B(n11049), .Z(n11050) );
  NAND U20812 ( .A(n29329), .B(n11050), .Z(n11051) );
  NANDN U20813 ( .A(n29330), .B(n11051), .Z(n11052) );
  NAND U20814 ( .A(n29331), .B(n11052), .Z(n11053) );
  NANDN U20815 ( .A(y[3902]), .B(x[3902]), .Z(n11429) );
  NANDN U20816 ( .A(y[3903]), .B(x[3903]), .Z(n11428) );
  AND U20817 ( .A(n11429), .B(n11428), .Z(n23897) );
  AND U20818 ( .A(n11053), .B(n23897), .Z(n11054) );
  ANDN U20819 ( .B(n29334), .A(n11054), .Z(n11055) );
  OR U20820 ( .A(n29335), .B(n11055), .Z(n11056) );
  NAND U20821 ( .A(n29336), .B(n11056), .Z(n11057) );
  NANDN U20822 ( .A(n29337), .B(n11057), .Z(n11058) );
  AND U20823 ( .A(n29338), .B(n11058), .Z(n11059) );
  NANDN U20824 ( .A(y[3908]), .B(x[3908]), .Z(n11423) );
  NANDN U20825 ( .A(y[3909]), .B(x[3909]), .Z(n11420) );
  NAND U20826 ( .A(n11423), .B(n11420), .Z(n29339) );
  OR U20827 ( .A(n11059), .B(n29339), .Z(n11060) );
  AND U20828 ( .A(n11061), .B(n11060), .Z(n11062) );
  OR U20829 ( .A(n29342), .B(n11062), .Z(n11063) );
  NAND U20830 ( .A(n29343), .B(n11063), .Z(n11064) );
  NANDN U20831 ( .A(n29344), .B(n11064), .Z(n11065) );
  AND U20832 ( .A(n29345), .B(n11065), .Z(n11066) );
  NANDN U20833 ( .A(y[3914]), .B(x[3914]), .Z(n11416) );
  NANDN U20834 ( .A(y[3915]), .B(x[3915]), .Z(n23382) );
  NAND U20835 ( .A(n11416), .B(n23382), .Z(n29346) );
  OR U20836 ( .A(n11066), .B(n29346), .Z(n11067) );
  AND U20837 ( .A(n29347), .B(n11067), .Z(n11068) );
  OR U20838 ( .A(n29348), .B(n11068), .Z(n11069) );
  NAND U20839 ( .A(n29349), .B(n11069), .Z(n11070) );
  NANDN U20840 ( .A(n29350), .B(n11070), .Z(n11071) );
  AND U20841 ( .A(n23394), .B(n11071), .Z(n11072) );
  NANDN U20842 ( .A(x[3919]), .B(y[3919]), .Z(n29351) );
  AND U20843 ( .A(n11072), .B(n29351), .Z(n11073) );
  OR U20844 ( .A(n29354), .B(n11073), .Z(n11074) );
  AND U20845 ( .A(n11075), .B(n11074), .Z(n11076) );
  OR U20846 ( .A(n29357), .B(n11076), .Z(n11077) );
  NAND U20847 ( .A(n29358), .B(n11077), .Z(n11078) );
  NANDN U20848 ( .A(n29359), .B(n11078), .Z(n11079) );
  AND U20849 ( .A(n29360), .B(n11079), .Z(n11080) );
  NANDN U20850 ( .A(y[3926]), .B(x[3926]), .Z(n11402) );
  NANDN U20851 ( .A(y[3927]), .B(x[3927]), .Z(n23414) );
  NAND U20852 ( .A(n11402), .B(n23414), .Z(n29361) );
  OR U20853 ( .A(n11080), .B(n29361), .Z(n11081) );
  NANDN U20854 ( .A(x[3927]), .B(y[3927]), .Z(n11401) );
  NANDN U20855 ( .A(x[3928]), .B(y[3928]), .Z(n11399) );
  AND U20856 ( .A(n11401), .B(n11399), .Z(n29362) );
  AND U20857 ( .A(n11081), .B(n29362), .Z(n11082) );
  NANDN U20858 ( .A(y[3928]), .B(x[3928]), .Z(n23412) );
  NANDN U20859 ( .A(y[3929]), .B(x[3929]), .Z(n11397) );
  NAND U20860 ( .A(n23412), .B(n11397), .Z(n23896) );
  OR U20861 ( .A(n11082), .B(n23896), .Z(n11083) );
  NAND U20862 ( .A(n23895), .B(n11083), .Z(n11084) );
  NANDN U20863 ( .A(n29363), .B(n11084), .Z(n11085) );
  NANDN U20864 ( .A(x[3931]), .B(y[3931]), .Z(n11394) );
  NANDN U20865 ( .A(x[3932]), .B(y[3932]), .Z(n23424) );
  AND U20866 ( .A(n11394), .B(n23424), .Z(n29364) );
  AND U20867 ( .A(n11085), .B(n29364), .Z(n11086) );
  NANDN U20868 ( .A(y[3932]), .B(x[3932]), .Z(n11392) );
  NANDN U20869 ( .A(y[3933]), .B(x[3933]), .Z(n23428) );
  AND U20870 ( .A(n11392), .B(n23428), .Z(n29366) );
  NANDN U20871 ( .A(n11086), .B(n29366), .Z(n11087) );
  NAND U20872 ( .A(n29367), .B(n11087), .Z(n11088) );
  NANDN U20873 ( .A(n29368), .B(n11088), .Z(n11089) );
  AND U20874 ( .A(n23434), .B(n11089), .Z(n11090) );
  NANDN U20875 ( .A(x[3935]), .B(y[3935]), .Z(n23893) );
  AND U20876 ( .A(n11090), .B(n23893), .Z(n11092) );
  NANDN U20877 ( .A(y[3936]), .B(x[3936]), .Z(n11091) );
  NANDN U20878 ( .A(y[3937]), .B(x[3937]), .Z(n11389) );
  NAND U20879 ( .A(n11091), .B(n11389), .Z(n29369) );
  OR U20880 ( .A(n11092), .B(n29369), .Z(n11093) );
  AND U20881 ( .A(n11390), .B(n11093), .Z(n11094) );
  NANDN U20882 ( .A(x[3937]), .B(y[3937]), .Z(n29370) );
  AND U20883 ( .A(n11094), .B(n29370), .Z(n11096) );
  NANDN U20884 ( .A(y[3938]), .B(x[3938]), .Z(n11095) );
  NANDN U20885 ( .A(y[3939]), .B(x[3939]), .Z(n11387) );
  NAND U20886 ( .A(n11095), .B(n11387), .Z(n29372) );
  OR U20887 ( .A(n11096), .B(n29372), .Z(n11097) );
  NANDN U20888 ( .A(x[3939]), .B(y[3939]), .Z(n11388) );
  NANDN U20889 ( .A(x[3940]), .B(y[3940]), .Z(n11385) );
  AND U20890 ( .A(n11388), .B(n11385), .Z(n29373) );
  AND U20891 ( .A(n11097), .B(n29373), .Z(n11098) );
  NANDN U20892 ( .A(y[3940]), .B(x[3940]), .Z(n11386) );
  NANDN U20893 ( .A(y[3941]), .B(x[3941]), .Z(n11383) );
  NAND U20894 ( .A(n11386), .B(n11383), .Z(n23892) );
  OR U20895 ( .A(n11098), .B(n23892), .Z(n11099) );
  NAND U20896 ( .A(n23891), .B(n11099), .Z(n11100) );
  NANDN U20897 ( .A(n29374), .B(n11100), .Z(n11101) );
  NANDN U20898 ( .A(x[3943]), .B(y[3943]), .Z(n23449) );
  NANDN U20899 ( .A(x[3944]), .B(y[3944]), .Z(n11381) );
  AND U20900 ( .A(n23449), .B(n11381), .Z(n29377) );
  AND U20901 ( .A(n11101), .B(n29377), .Z(n11102) );
  NANDN U20902 ( .A(y[3944]), .B(x[3944]), .Z(n23453) );
  NANDN U20903 ( .A(y[3945]), .B(x[3945]), .Z(n23460) );
  AND U20904 ( .A(n23453), .B(n23460), .Z(n29378) );
  NANDN U20905 ( .A(n11102), .B(n29378), .Z(n11103) );
  NAND U20906 ( .A(n29379), .B(n11103), .Z(n11104) );
  NANDN U20907 ( .A(n29380), .B(n11104), .Z(n11105) );
  AND U20908 ( .A(n23466), .B(n11105), .Z(n11106) );
  NANDN U20909 ( .A(x[3947]), .B(y[3947]), .Z(n23889) );
  NAND U20910 ( .A(n11106), .B(n23889), .Z(n11107) );
  NANDN U20911 ( .A(n29381), .B(n11107), .Z(n11108) );
  AND U20912 ( .A(n29382), .B(n11108), .Z(n11109) );
  OR U20913 ( .A(n29383), .B(n11109), .Z(n11110) );
  NAND U20914 ( .A(n29384), .B(n11110), .Z(n11111) );
  NANDN U20915 ( .A(n29385), .B(n11111), .Z(n11112) );
  AND U20916 ( .A(n29386), .B(n11112), .Z(n11113) );
  NANDN U20917 ( .A(y[3954]), .B(x[3954]), .Z(n11372) );
  NANDN U20918 ( .A(y[3955]), .B(x[3955]), .Z(n23489) );
  NAND U20919 ( .A(n11372), .B(n23489), .Z(n29387) );
  OR U20920 ( .A(n11113), .B(n29387), .Z(n11114) );
  AND U20921 ( .A(n29388), .B(n11114), .Z(n11115) );
  OR U20922 ( .A(n29389), .B(n11115), .Z(n11116) );
  NAND U20923 ( .A(n29390), .B(n11116), .Z(n11117) );
  NANDN U20924 ( .A(n29391), .B(n11117), .Z(n11118) );
  NANDN U20925 ( .A(x[3959]), .B(y[3959]), .Z(n11366) );
  NANDN U20926 ( .A(x[3960]), .B(y[3960]), .Z(n23504) );
  AND U20927 ( .A(n11366), .B(n23504), .Z(n23888) );
  AND U20928 ( .A(n11118), .B(n23888), .Z(n11119) );
  NANDN U20929 ( .A(y[3960]), .B(x[3960]), .Z(n23500) );
  NANDN U20930 ( .A(y[3961]), .B(x[3961]), .Z(n11365) );
  AND U20931 ( .A(n23500), .B(n11365), .Z(n29393) );
  NANDN U20932 ( .A(n11119), .B(n29393), .Z(n11120) );
  NANDN U20933 ( .A(n29394), .B(n11120), .Z(n11121) );
  AND U20934 ( .A(n29395), .B(n11121), .Z(n11122) );
  OR U20935 ( .A(n29396), .B(n11122), .Z(n11123) );
  NAND U20936 ( .A(n29397), .B(n11123), .Z(n11124) );
  NANDN U20937 ( .A(n29398), .B(n11124), .Z(n11125) );
  AND U20938 ( .A(n29399), .B(n11125), .Z(n11128) );
  ANDN U20939 ( .B(y[3967]), .A(x[3967]), .Z(n11356) );
  XOR U20940 ( .A(x[3968]), .B(y[3968]), .Z(n11126) );
  NOR U20941 ( .A(n11356), .B(n11126), .Z(n11127) );
  NANDN U20942 ( .A(n11128), .B(n11127), .Z(n11130) );
  NANDN U20943 ( .A(y[3968]), .B(x[3968]), .Z(n11129) );
  NANDN U20944 ( .A(y[3969]), .B(x[3969]), .Z(n11355) );
  AND U20945 ( .A(n11129), .B(n11355), .Z(n29402) );
  AND U20946 ( .A(n11130), .B(n29402), .Z(n11131) );
  NANDN U20947 ( .A(x[3969]), .B(y[3969]), .Z(n23525) );
  NANDN U20948 ( .A(x[3970]), .B(y[3970]), .Z(n11353) );
  NAND U20949 ( .A(n23525), .B(n11353), .Z(n29403) );
  OR U20950 ( .A(n11131), .B(n29403), .Z(n11132) );
  NAND U20951 ( .A(n29404), .B(n11132), .Z(n11133) );
  NANDN U20952 ( .A(n23887), .B(n11133), .Z(n11134) );
  NANDN U20953 ( .A(y[3972]), .B(x[3972]), .Z(n11350) );
  NANDN U20954 ( .A(y[3973]), .B(x[3973]), .Z(n11349) );
  AND U20955 ( .A(n11350), .B(n11349), .Z(n23886) );
  AND U20956 ( .A(n11134), .B(n23886), .Z(n11135) );
  NANDN U20957 ( .A(x[3973]), .B(y[3973]), .Z(n23535) );
  NANDN U20958 ( .A(x[3974]), .B(y[3974]), .Z(n23542) );
  NAND U20959 ( .A(n23535), .B(n23542), .Z(n29407) );
  OR U20960 ( .A(n11135), .B(n29407), .Z(n11136) );
  AND U20961 ( .A(n29409), .B(n11136), .Z(n11137) );
  OR U20962 ( .A(n29410), .B(n11137), .Z(n11138) );
  NAND U20963 ( .A(n29411), .B(n11138), .Z(n11139) );
  NANDN U20964 ( .A(n29412), .B(n11139), .Z(n11140) );
  AND U20965 ( .A(n29413), .B(n11140), .Z(n11141) );
  NANDN U20966 ( .A(x[3979]), .B(y[3979]), .Z(n11344) );
  NANDN U20967 ( .A(x[3980]), .B(y[3980]), .Z(n11343) );
  AND U20968 ( .A(n11344), .B(n11343), .Z(n23885) );
  NANDN U20969 ( .A(n11141), .B(n23885), .Z(n11142) );
  NANDN U20970 ( .A(n29414), .B(n11142), .Z(n11143) );
  AND U20971 ( .A(n29415), .B(n11143), .Z(n11144) );
  NANDN U20972 ( .A(y[3982]), .B(x[3982]), .Z(n23565) );
  NANDN U20973 ( .A(y[3983]), .B(x[3983]), .Z(n11339) );
  NAND U20974 ( .A(n23565), .B(n11339), .Z(n29416) );
  OR U20975 ( .A(n11144), .B(n29416), .Z(n11145) );
  NAND U20976 ( .A(n29417), .B(n11145), .Z(n11146) );
  NANDN U20977 ( .A(n23884), .B(n11146), .Z(n11147) );
  NANDN U20978 ( .A(x[3985]), .B(y[3985]), .Z(n11336) );
  NANDN U20979 ( .A(x[3986]), .B(y[3986]), .Z(n11335) );
  AND U20980 ( .A(n11336), .B(n11335), .Z(n23883) );
  AND U20981 ( .A(n11147), .B(n23883), .Z(n11148) );
  NANDN U20982 ( .A(y[3986]), .B(x[3986]), .Z(n23573) );
  NANDN U20983 ( .A(y[3987]), .B(x[3987]), .Z(n23580) );
  NAND U20984 ( .A(n23573), .B(n23580), .Z(n29418) );
  OR U20985 ( .A(n11148), .B(n29418), .Z(n11149) );
  NAND U20986 ( .A(n11150), .B(n11149), .Z(n11152) );
  NANDN U20987 ( .A(y[3988]), .B(x[3988]), .Z(n11151) );
  NANDN U20988 ( .A(y[3989]), .B(x[3989]), .Z(n23586) );
  AND U20989 ( .A(n11151), .B(n23586), .Z(n23882) );
  AND U20990 ( .A(n11152), .B(n23882), .Z(n11153) );
  NOR U20991 ( .A(n11334), .B(n11153), .Z(n11154) );
  NAND U20992 ( .A(n23585), .B(n11154), .Z(n11155) );
  NANDN U20993 ( .A(n29426), .B(n11155), .Z(n11156) );
  AND U20994 ( .A(n11333), .B(n11156), .Z(n11157) );
  NANDN U20995 ( .A(x[3991]), .B(y[3991]), .Z(n23880) );
  AND U20996 ( .A(n11157), .B(n23880), .Z(n11159) );
  NANDN U20997 ( .A(y[3992]), .B(x[3992]), .Z(n11158) );
  NANDN U20998 ( .A(y[3993]), .B(x[3993]), .Z(n11329) );
  NAND U20999 ( .A(n11158), .B(n11329), .Z(n29427) );
  OR U21000 ( .A(n11159), .B(n29427), .Z(n11160) );
  AND U21001 ( .A(n11330), .B(n11160), .Z(n11161) );
  NANDN U21002 ( .A(x[3993]), .B(y[3993]), .Z(n11331) );
  AND U21003 ( .A(n11161), .B(n11331), .Z(n11163) );
  NANDN U21004 ( .A(y[3994]), .B(x[3994]), .Z(n11162) );
  NANDN U21005 ( .A(y[3995]), .B(x[3995]), .Z(n11328) );
  NAND U21006 ( .A(n11162), .B(n11328), .Z(n29430) );
  OR U21007 ( .A(n11163), .B(n29430), .Z(n11164) );
  AND U21008 ( .A(n29431), .B(n11164), .Z(n11165) );
  NANDN U21009 ( .A(y[3996]), .B(x[3996]), .Z(n11327) );
  NANDN U21010 ( .A(y[3997]), .B(x[3997]), .Z(n11326) );
  NAND U21011 ( .A(n11327), .B(n11326), .Z(n23879) );
  OR U21012 ( .A(n11165), .B(n23879), .Z(n11166) );
  NAND U21013 ( .A(n29434), .B(n11166), .Z(n11167) );
  NANDN U21014 ( .A(n29435), .B(n11167), .Z(n11168) );
  NANDN U21015 ( .A(x[3999]), .B(y[3999]), .Z(n23607) );
  NANDN U21016 ( .A(x[4000]), .B(y[4000]), .Z(n11324) );
  AND U21017 ( .A(n23607), .B(n11324), .Z(n29436) );
  AND U21018 ( .A(n11168), .B(n29436), .Z(n11169) );
  NANDN U21019 ( .A(y[4000]), .B(x[4000]), .Z(n23611) );
  NANDN U21020 ( .A(y[4001]), .B(x[4001]), .Z(n23618) );
  AND U21021 ( .A(n23611), .B(n23618), .Z(n29437) );
  NANDN U21022 ( .A(n11169), .B(n29437), .Z(n11170) );
  NANDN U21023 ( .A(n29438), .B(n11170), .Z(n11171) );
  AND U21024 ( .A(n29439), .B(n11171), .Z(n11172) );
  NANDN U21025 ( .A(x[4003]), .B(y[4003]), .Z(n11321) );
  NANDN U21026 ( .A(x[4004]), .B(y[4004]), .Z(n11320) );
  NAND U21027 ( .A(n11321), .B(n11320), .Z(n29440) );
  OR U21028 ( .A(n11172), .B(n29440), .Z(n11173) );
  NAND U21029 ( .A(n29441), .B(n11173), .Z(n11174) );
  NANDN U21030 ( .A(n23878), .B(n11174), .Z(n11175) );
  NANDN U21031 ( .A(y[4006]), .B(x[4006]), .Z(n23629) );
  NANDN U21032 ( .A(y[4007]), .B(x[4007]), .Z(n23635) );
  AND U21033 ( .A(n23629), .B(n23635), .Z(n23877) );
  AND U21034 ( .A(n11175), .B(n23877), .Z(n11177) );
  XNOR U21035 ( .A(x[4008]), .B(y[4008]), .Z(n23636) );
  ANDN U21036 ( .B(y[4007]), .A(x[4007]), .Z(n11317) );
  ANDN U21037 ( .B(n23636), .A(n11317), .Z(n11176) );
  NANDN U21038 ( .A(n11177), .B(n11176), .Z(n11178) );
  AND U21039 ( .A(n29444), .B(n11178), .Z(n11179) );
  OR U21040 ( .A(n29445), .B(n11179), .Z(n11180) );
  NAND U21041 ( .A(n29446), .B(n11180), .Z(n11181) );
  NANDN U21042 ( .A(n29447), .B(n11181), .Z(n11182) );
  NAND U21043 ( .A(n29448), .B(n11182), .Z(n11183) );
  AND U21044 ( .A(n11310), .B(n11183), .Z(n11184) );
  NAND U21045 ( .A(n29449), .B(n11184), .Z(n11185) );
  NANDN U21046 ( .A(n29451), .B(n11185), .Z(n11186) );
  AND U21047 ( .A(n29452), .B(n11186), .Z(n11187) );
  NANDN U21048 ( .A(y[4016]), .B(x[4016]), .Z(n23657) );
  NANDN U21049 ( .A(y[4017]), .B(x[4017]), .Z(n23664) );
  NAND U21050 ( .A(n23657), .B(n23664), .Z(n29453) );
  OR U21051 ( .A(n11187), .B(n29453), .Z(n11188) );
  AND U21052 ( .A(n11189), .B(n11188), .Z(n11191) );
  NANDN U21053 ( .A(y[4018]), .B(x[4018]), .Z(n11190) );
  NANDN U21054 ( .A(y[4019]), .B(x[4019]), .Z(n23670) );
  NAND U21055 ( .A(n11190), .B(n23670), .Z(n29456) );
  OR U21056 ( .A(n11191), .B(n29456), .Z(n11192) );
  NAND U21057 ( .A(n29457), .B(n11192), .Z(n11193) );
  NANDN U21058 ( .A(n23875), .B(n11193), .Z(n11194) );
  NANDN U21059 ( .A(x[4021]), .B(y[4021]), .Z(n23672) );
  NANDN U21060 ( .A(x[4022]), .B(y[4022]), .Z(n11304) );
  AND U21061 ( .A(n23672), .B(n11304), .Z(n23874) );
  AND U21062 ( .A(n11194), .B(n23874), .Z(n11195) );
  NANDN U21063 ( .A(y[4022]), .B(x[4022]), .Z(n11305) );
  NANDN U21064 ( .A(y[4023]), .B(x[4023]), .Z(n11303) );
  NAND U21065 ( .A(n11305), .B(n11303), .Z(n29459) );
  OR U21066 ( .A(n11195), .B(n29459), .Z(n11196) );
  AND U21067 ( .A(n11197), .B(n11196), .Z(n11199) );
  NANDN U21068 ( .A(y[4024]), .B(x[4024]), .Z(n11198) );
  NANDN U21069 ( .A(y[4025]), .B(x[4025]), .Z(n11301) );
  NAND U21070 ( .A(n11198), .B(n11301), .Z(n29462) );
  OR U21071 ( .A(n11199), .B(n29462), .Z(n11200) );
  NAND U21072 ( .A(n29463), .B(n11200), .Z(n11201) );
  NANDN U21073 ( .A(n23873), .B(n11201), .Z(n11202) );
  NANDN U21074 ( .A(x[4027]), .B(y[4027]), .Z(n11298) );
  NANDN U21075 ( .A(x[4028]), .B(y[4028]), .Z(n23693) );
  AND U21076 ( .A(n11298), .B(n23693), .Z(n23872) );
  AND U21077 ( .A(n11202), .B(n23872), .Z(n11203) );
  NANDN U21078 ( .A(y[4028]), .B(x[4028]), .Z(n11296) );
  NANDN U21079 ( .A(y[4029]), .B(x[4029]), .Z(n11295) );
  NAND U21080 ( .A(n11296), .B(n11295), .Z(n29464) );
  OR U21081 ( .A(n11203), .B(n29464), .Z(n11204) );
  NANDN U21082 ( .A(x[4029]), .B(y[4029]), .Z(n23692) );
  NANDN U21083 ( .A(x[4030]), .B(y[4030]), .Z(n23699) );
  AND U21084 ( .A(n23692), .B(n23699), .Z(n29465) );
  AND U21085 ( .A(n11204), .B(n29465), .Z(n11205) );
  NANDN U21086 ( .A(y[4030]), .B(x[4030]), .Z(n11294) );
  NANDN U21087 ( .A(y[4031]), .B(x[4031]), .Z(n11293) );
  NAND U21088 ( .A(n11294), .B(n11293), .Z(n29466) );
  OR U21089 ( .A(n11205), .B(n29466), .Z(n11206) );
  NAND U21090 ( .A(n29469), .B(n11206), .Z(n11207) );
  NANDN U21091 ( .A(n23871), .B(n11207), .Z(n11208) );
  NANDN U21092 ( .A(x[4033]), .B(y[4033]), .Z(n23704) );
  NANDN U21093 ( .A(x[4034]), .B(y[4034]), .Z(n11291) );
  AND U21094 ( .A(n23704), .B(n11291), .Z(n23870) );
  AND U21095 ( .A(n11208), .B(n23870), .Z(n11209) );
  NANDN U21096 ( .A(y[4034]), .B(x[4034]), .Z(n23707) );
  NANDN U21097 ( .A(y[4035]), .B(x[4035]), .Z(n23714) );
  AND U21098 ( .A(n23707), .B(n23714), .Z(n29470) );
  NANDN U21099 ( .A(n11209), .B(n29470), .Z(n11210) );
  NANDN U21100 ( .A(y[4036]), .B(x[4036]), .Z(n23713) );
  NANDN U21101 ( .A(y[4037]), .B(x[4037]), .Z(n23720) );
  AND U21102 ( .A(n23713), .B(n23720), .Z(n23869) );
  NANDN U21103 ( .A(x[4037]), .B(y[4037]), .Z(n11288) );
  NANDN U21104 ( .A(x[4038]), .B(y[4038]), .Z(n11287) );
  NAND U21105 ( .A(n11288), .B(n11287), .Z(n29472) );
  NANDN U21106 ( .A(y[4040]), .B(x[4040]), .Z(n23725) );
  NANDN U21107 ( .A(y[4041]), .B(x[4041]), .Z(n23732) );
  AND U21108 ( .A(n23725), .B(n23732), .Z(n23867) );
  NANDN U21109 ( .A(x[4041]), .B(y[4041]), .Z(n11284) );
  NANDN U21110 ( .A(x[4042]), .B(y[4042]), .Z(n11283) );
  NAND U21111 ( .A(n11284), .B(n11283), .Z(n29474) );
  NANDN U21112 ( .A(y[4042]), .B(x[4042]), .Z(n23731) );
  NANDN U21113 ( .A(y[4043]), .B(x[4043]), .Z(n23740) );
  AND U21114 ( .A(n23731), .B(n23740), .Z(n29477) );
  ANDN U21115 ( .B(y[4044]), .A(x[4044]), .Z(n23744) );
  NANDN U21116 ( .A(x[4043]), .B(y[4043]), .Z(n11282) );
  NANDN U21117 ( .A(n23744), .B(n11282), .Z(n29478) );
  NANDN U21118 ( .A(y[4046]), .B(x[4046]), .Z(n23746) );
  NANDN U21119 ( .A(y[4047]), .B(x[4047]), .Z(n23753) );
  AND U21120 ( .A(n23746), .B(n23753), .Z(n23865) );
  NANDN U21121 ( .A(x[4047]), .B(y[4047]), .Z(n11280) );
  NANDN U21122 ( .A(x[4048]), .B(y[4048]), .Z(n11279) );
  NAND U21123 ( .A(n11280), .B(n11279), .Z(n29480) );
  NANDN U21124 ( .A(y[4050]), .B(x[4050]), .Z(n23758) );
  NANDN U21125 ( .A(y[4051]), .B(x[4051]), .Z(n23764) );
  AND U21126 ( .A(n23758), .B(n23764), .Z(n23863) );
  NANDN U21127 ( .A(y[4052]), .B(x[4052]), .Z(n11211) );
  NANDN U21128 ( .A(y[4053]), .B(x[4053]), .Z(n11274) );
  AND U21129 ( .A(n11211), .B(n11274), .Z(n29485) );
  NANDN U21130 ( .A(y[4056]), .B(x[4056]), .Z(n11272) );
  NANDN U21131 ( .A(y[4057]), .B(x[4057]), .Z(n11269) );
  AND U21132 ( .A(n11272), .B(n11269), .Z(n29490) );
  NANDN U21133 ( .A(y[4060]), .B(x[4060]), .Z(n11213) );
  NANDN U21134 ( .A(y[4061]), .B(x[4061]), .Z(n23789) );
  AND U21135 ( .A(n11213), .B(n23789), .Z(n29494) );
  XNOR U21136 ( .A(x[4062]), .B(y[4062]), .Z(n23788) );
  ANDN U21137 ( .B(y[4061]), .A(x[4061]), .Z(n11265) );
  NANDN U21138 ( .A(y[4062]), .B(x[4062]), .Z(n11214) );
  NANDN U21139 ( .A(y[4063]), .B(x[4063]), .Z(n23795) );
  AND U21140 ( .A(n11214), .B(n23795), .Z(n29497) );
  NANDN U21141 ( .A(x[4063]), .B(y[4063]), .Z(n11264) );
  NANDN U21142 ( .A(x[4064]), .B(y[4064]), .Z(n11263) );
  NAND U21143 ( .A(n11264), .B(n11263), .Z(n29500) );
  NANDN U21144 ( .A(y[4066]), .B(x[4066]), .Z(n23800) );
  NANDN U21145 ( .A(y[4067]), .B(x[4067]), .Z(n23805) );
  AND U21146 ( .A(n23800), .B(n23805), .Z(n23859) );
  AND U21147 ( .A(n11215), .B(n23859), .Z(n11217) );
  XNOR U21148 ( .A(x[4068]), .B(y[4068]), .Z(n23806) );
  NANDN U21149 ( .A(x[4067]), .B(y[4067]), .Z(n29502) );
  NAND U21150 ( .A(n23806), .B(n29502), .Z(n11216) );
  OR U21151 ( .A(n11217), .B(n11216), .Z(n11219) );
  NANDN U21152 ( .A(y[4068]), .B(x[4068]), .Z(n11218) );
  NANDN U21153 ( .A(y[4069]), .B(x[4069]), .Z(n11259) );
  AND U21154 ( .A(n11218), .B(n11259), .Z(n29504) );
  AND U21155 ( .A(n11219), .B(n29504), .Z(n11220) );
  ANDN U21156 ( .B(n11260), .A(n11220), .Z(n11221) );
  NANDN U21157 ( .A(x[4069]), .B(y[4069]), .Z(n23858) );
  NAND U21158 ( .A(n11221), .B(n23858), .Z(n11222) );
  NANDN U21159 ( .A(n29505), .B(n11222), .Z(n11223) );
  AND U21160 ( .A(n11257), .B(n11223), .Z(n11224) );
  NANDN U21161 ( .A(x[4071]), .B(y[4071]), .Z(n11258) );
  AND U21162 ( .A(n11224), .B(n11258), .Z(n11226) );
  NANDN U21163 ( .A(y[4072]), .B(x[4072]), .Z(n11225) );
  NANDN U21164 ( .A(y[4073]), .B(x[4073]), .Z(n11255) );
  NAND U21165 ( .A(n11225), .B(n11255), .Z(n29508) );
  OR U21166 ( .A(n11226), .B(n29508), .Z(n11227) );
  AND U21167 ( .A(n29510), .B(n11227), .Z(n11228) );
  NANDN U21168 ( .A(y[4074]), .B(x[4074]), .Z(n11254) );
  NANDN U21169 ( .A(y[4075]), .B(x[4075]), .Z(n11251) );
  NAND U21170 ( .A(n11254), .B(n11251), .Z(n29511) );
  OR U21171 ( .A(n11228), .B(n29511), .Z(n11229) );
  AND U21172 ( .A(n11252), .B(n11229), .Z(n11230) );
  NAND U21173 ( .A(n23855), .B(n11230), .Z(n11231) );
  NANDN U21174 ( .A(n29513), .B(n11231), .Z(n11232) );
  AND U21175 ( .A(n23829), .B(n11232), .Z(n11233) );
  NANDN U21176 ( .A(x[4077]), .B(y[4077]), .Z(n11250) );
  AND U21177 ( .A(n11233), .B(n11250), .Z(n11235) );
  NANDN U21178 ( .A(y[4078]), .B(x[4078]), .Z(n11234) );
  NANDN U21179 ( .A(y[4079]), .B(x[4079]), .Z(n23836) );
  NAND U21180 ( .A(n11234), .B(n23836), .Z(n29516) );
  OR U21181 ( .A(n11235), .B(n29516), .Z(n11236) );
  NANDN U21182 ( .A(x[4079]), .B(y[4079]), .Z(n11249) );
  NANDN U21183 ( .A(x[4080]), .B(y[4080]), .Z(n11248) );
  AND U21184 ( .A(n11249), .B(n11248), .Z(n29517) );
  AND U21185 ( .A(n11236), .B(n29517), .Z(n11237) );
  NANDN U21186 ( .A(y[4080]), .B(x[4080]), .Z(n23835) );
  NANDN U21187 ( .A(y[4081]), .B(x[4081]), .Z(n23842) );
  NAND U21188 ( .A(n23835), .B(n23842), .Z(n23854) );
  OR U21189 ( .A(n11237), .B(n23854), .Z(n11238) );
  NAND U21190 ( .A(n23853), .B(n11238), .Z(n11239) );
  NANDN U21191 ( .A(n29518), .B(n11239), .Z(n11240) );
  NAND U21192 ( .A(n29519), .B(n11240), .Z(n11241) );
  AND U21193 ( .A(n11242), .B(n11241), .Z(n23849) );
  AND U21194 ( .A(n11244), .B(n11243), .Z(n23847) );
  NAND U21195 ( .A(n11246), .B(n11245), .Z(n23845) );
  NAND U21196 ( .A(n11248), .B(n11247), .Z(n23839) );
  NANDN U21197 ( .A(x[4078]), .B(y[4078]), .Z(n29515) );
  NAND U21198 ( .A(n29515), .B(n11249), .Z(n23833) );
  IV U21199 ( .A(n11250), .Z(n29514) );
  ANDN U21200 ( .B(y[4076]), .A(x[4076]), .Z(n23856) );
  AND U21201 ( .A(n11252), .B(n11251), .Z(n23825) );
  NAND U21202 ( .A(n23855), .B(n11253), .Z(n23823) );
  AND U21203 ( .A(n11255), .B(n11254), .Z(n23821) );
  AND U21204 ( .A(n11257), .B(n11256), .Z(n23816) );
  IV U21205 ( .A(n11258), .Z(n29507) );
  AND U21206 ( .A(n11260), .B(n11259), .Z(n23812) );
  NANDN U21207 ( .A(x[4068]), .B(y[4068]), .Z(n29503) );
  NAND U21208 ( .A(n29503), .B(n23858), .Z(n23810) );
  AND U21209 ( .A(n11261), .B(n29502), .Z(n23804) );
  NAND U21210 ( .A(n11263), .B(n11262), .Z(n23798) );
  NANDN U21211 ( .A(x[4062]), .B(y[4062]), .Z(n29496) );
  NAND U21212 ( .A(n29496), .B(n11264), .Z(n23792) );
  IV U21213 ( .A(n11265), .Z(n29495) );
  NANDN U21214 ( .A(x[4060]), .B(y[4060]), .Z(n29493) );
  NAND U21215 ( .A(n29495), .B(n29493), .Z(n23786) );
  XNOR U21216 ( .A(x[4060]), .B(y[4060]), .Z(n11267) );
  AND U21217 ( .A(n11267), .B(n11266), .Z(n23784) );
  NANDN U21218 ( .A(x[4058]), .B(y[4058]), .Z(n23862) );
  IV U21219 ( .A(n11268), .Z(n29492) );
  AND U21220 ( .A(n23862), .B(n29492), .Z(n23782) );
  NAND U21221 ( .A(n11270), .B(n11269), .Z(n23780) );
  IV U21222 ( .A(n11271), .Z(n23861) );
  AND U21223 ( .A(n11273), .B(n11272), .Z(n23775) );
  AND U21224 ( .A(n11275), .B(n11274), .Z(n23770) );
  IV U21225 ( .A(n11276), .Z(n29482) );
  NAND U21226 ( .A(n29482), .B(n11277), .Z(n23762) );
  NAND U21227 ( .A(n11279), .B(n11278), .Z(n23756) );
  NAND U21228 ( .A(n11281), .B(n11280), .Z(n23750) );
  AND U21229 ( .A(n11283), .B(n11282), .Z(n23736) );
  AND U21230 ( .A(n11285), .B(n11284), .Z(n23730) );
  AND U21231 ( .A(n11287), .B(n11286), .Z(n23724) );
  AND U21232 ( .A(n11289), .B(n11288), .Z(n23718) );
  AND U21233 ( .A(n11291), .B(n11290), .Z(n23712) );
  NAND U21234 ( .A(n11293), .B(n11292), .Z(n23702) );
  NAND U21235 ( .A(n11295), .B(n11294), .Z(n23696) );
  NAND U21236 ( .A(n11297), .B(n11296), .Z(n23690) );
  AND U21237 ( .A(n11299), .B(n11298), .Z(n23688) );
  NAND U21238 ( .A(n11301), .B(n11300), .Z(n23686) );
  AND U21239 ( .A(n11303), .B(n11302), .Z(n23681) );
  NAND U21240 ( .A(n11304), .B(n29460), .Z(n23679) );
  AND U21241 ( .A(n11306), .B(n11305), .Z(n23677) );
  NANDN U21242 ( .A(x[4018]), .B(y[4018]), .Z(n29455) );
  NAND U21243 ( .A(n29455), .B(n11307), .Z(n23667) );
  NAND U21244 ( .A(n29454), .B(n11308), .Z(n23661) );
  ANDN U21245 ( .B(y[4014]), .A(x[4014]), .Z(n29450) );
  AND U21246 ( .A(n11310), .B(n11309), .Z(n23652) );
  AND U21247 ( .A(n29449), .B(n11311), .Z(n23650) );
  NAND U21248 ( .A(n11313), .B(n11312), .Z(n23648) );
  AND U21249 ( .A(n11315), .B(n11314), .Z(n23646) );
  NANDN U21250 ( .A(x[4008]), .B(y[4008]), .Z(n23876) );
  AND U21251 ( .A(n11316), .B(n23876), .Z(n23640) );
  IV U21252 ( .A(n11317), .Z(n29442) );
  AND U21253 ( .A(n11318), .B(n29442), .Z(n23634) );
  AND U21254 ( .A(n11320), .B(n11319), .Z(n23628) );
  AND U21255 ( .A(n11322), .B(n11321), .Z(n23622) );
  AND U21256 ( .A(n11324), .B(n11323), .Z(n23616) );
  AND U21257 ( .A(n11326), .B(n11325), .Z(n23606) );
  AND U21258 ( .A(n11328), .B(n11327), .Z(n23600) );
  AND U21259 ( .A(n11330), .B(n11329), .Z(n23595) );
  IV U21260 ( .A(n11331), .Z(n29429) );
  AND U21261 ( .A(n11333), .B(n11332), .Z(n23591) );
  ANDN U21262 ( .B(y[3990]), .A(x[3990]), .Z(n29425) );
  NANDN U21263 ( .A(x[3988]), .B(y[3988]), .Z(n29421) );
  IV U21264 ( .A(n11334), .Z(n29424) );
  NAND U21265 ( .A(n29421), .B(n29424), .Z(n23583) );
  NAND U21266 ( .A(n29423), .B(n11335), .Z(n23577) );
  NAND U21267 ( .A(n11337), .B(n11336), .Z(n23571) );
  AND U21268 ( .A(n11339), .B(n11338), .Z(n23569) );
  NAND U21269 ( .A(n11341), .B(n11340), .Z(n23567) );
  AND U21270 ( .A(n11343), .B(n11342), .Z(n23561) );
  AND U21271 ( .A(n11345), .B(n11344), .Z(n23555) );
  NAND U21272 ( .A(n11347), .B(n11346), .Z(n23545) );
  NAND U21273 ( .A(n11349), .B(n11348), .Z(n23539) );
  NAND U21274 ( .A(n11351), .B(n11350), .Z(n23533) );
  AND U21275 ( .A(n11353), .B(n11352), .Z(n23531) );
  NAND U21276 ( .A(n11355), .B(n11354), .Z(n23529) );
  IV U21277 ( .A(n11356), .Z(n29400) );
  AND U21278 ( .A(n11357), .B(n29400), .Z(n23520) );
  AND U21279 ( .A(n11359), .B(n11358), .Z(n23518) );
  NAND U21280 ( .A(n11361), .B(n11360), .Z(n23516) );
  AND U21281 ( .A(n11363), .B(n11362), .Z(n23514) );
  AND U21282 ( .A(n11365), .B(n11364), .Z(n23508) );
  NAND U21283 ( .A(n11367), .B(n11366), .Z(n23498) );
  NAND U21284 ( .A(n11369), .B(n11368), .Z(n23492) );
  NAND U21285 ( .A(n11371), .B(n11370), .Z(n23486) );
  AND U21286 ( .A(n11373), .B(n11372), .Z(n23484) );
  NAND U21287 ( .A(n11375), .B(n11374), .Z(n23482) );
  AND U21288 ( .A(n11377), .B(n11376), .Z(n23476) );
  NANDN U21289 ( .A(x[3948]), .B(y[3948]), .Z(n23890) );
  AND U21290 ( .A(n23890), .B(n11378), .Z(n23470) );
  AND U21291 ( .A(n11379), .B(n23889), .Z(n23464) );
  AND U21292 ( .A(n11381), .B(n11380), .Z(n23458) );
  AND U21293 ( .A(n11383), .B(n11382), .Z(n23448) );
  NAND U21294 ( .A(n11385), .B(n11384), .Z(n23446) );
  AND U21295 ( .A(n11387), .B(n11386), .Z(n23444) );
  NANDN U21296 ( .A(x[3938]), .B(y[3938]), .Z(n29371) );
  AND U21297 ( .A(n11388), .B(n29371), .Z(n23442) );
  NAND U21298 ( .A(n11390), .B(n11389), .Z(n23440) );
  NANDN U21299 ( .A(x[3936]), .B(y[3936]), .Z(n23894) );
  AND U21300 ( .A(n23894), .B(n29370), .Z(n23438) );
  AND U21301 ( .A(n11391), .B(n23893), .Z(n23432) );
  AND U21302 ( .A(n11393), .B(n11392), .Z(n23422) );
  NAND U21303 ( .A(n11395), .B(n11394), .Z(n23420) );
  AND U21304 ( .A(n11397), .B(n11396), .Z(n23418) );
  NAND U21305 ( .A(n11399), .B(n11398), .Z(n23416) );
  AND U21306 ( .A(n11401), .B(n11400), .Z(n23410) );
  NAND U21307 ( .A(n11403), .B(n11402), .Z(n23408) );
  AND U21308 ( .A(n11405), .B(n11404), .Z(n23406) );
  AND U21309 ( .A(n11407), .B(n11406), .Z(n23404) );
  NANDN U21310 ( .A(x[3922]), .B(y[3922]), .Z(n29356) );
  AND U21311 ( .A(n29356), .B(n11408), .Z(n23402) );
  NAND U21312 ( .A(n11410), .B(n11409), .Z(n23400) );
  NANDN U21313 ( .A(x[3920]), .B(y[3920]), .Z(n29352) );
  AND U21314 ( .A(n29352), .B(n29355), .Z(n23398) );
  AND U21315 ( .A(n11411), .B(n29351), .Z(n23392) );
  AND U21316 ( .A(n11413), .B(n11412), .Z(n23386) );
  AND U21317 ( .A(n11415), .B(n11414), .Z(n23380) );
  NAND U21318 ( .A(n11417), .B(n11416), .Z(n23378) );
  AND U21319 ( .A(n11419), .B(n11418), .Z(n23372) );
  AND U21320 ( .A(n11421), .B(n11420), .Z(n23367) );
  NAND U21321 ( .A(n11422), .B(n29340), .Z(n23365) );
  AND U21322 ( .A(n11424), .B(n11423), .Z(n23363) );
  AND U21323 ( .A(n11426), .B(n11425), .Z(n23357) );
  AND U21324 ( .A(n11428), .B(n11427), .Z(n23351) );
  AND U21325 ( .A(n11430), .B(n11429), .Z(n23345) );
  AND U21326 ( .A(n11432), .B(n11431), .Z(n23339) );
  NANDN U21327 ( .A(x[3896]), .B(y[3896]), .Z(n29324) );
  NAND U21328 ( .A(n29324), .B(n29327), .Z(n23330) );
  NAND U21329 ( .A(n11433), .B(n29325), .Z(n23324) );
  AND U21330 ( .A(n11435), .B(n11434), .Z(n23322) );
  AND U21331 ( .A(n11437), .B(n11436), .Z(n23320) );
  NAND U21332 ( .A(n11439), .B(n11438), .Z(n23318) );
  NANDN U21333 ( .A(x[3890]), .B(y[3890]), .Z(n29318) );
  AND U21334 ( .A(n11440), .B(n29318), .Z(n23316) );
  NAND U21335 ( .A(n11442), .B(n11441), .Z(n23307) );
  NAND U21336 ( .A(n11444), .B(n11443), .Z(n23301) );
  NAND U21337 ( .A(n11446), .B(n11445), .Z(n23295) );
  NANDN U21338 ( .A(x[3882]), .B(y[3882]), .Z(n23904) );
  NAND U21339 ( .A(n11448), .B(n11447), .Z(n23290) );
  IV U21340 ( .A(n11449), .Z(n23903) );
  AND U21341 ( .A(n11450), .B(n23903), .Z(n23288) );
  AND U21342 ( .A(n11452), .B(n11451), .Z(n23286) );
  AND U21343 ( .A(n11453), .B(n29308), .Z(n23277) );
  AND U21344 ( .A(n11455), .B(n11454), .Z(n23275) );
  NAND U21345 ( .A(n11457), .B(n11456), .Z(n23273) );
  AND U21346 ( .A(n11459), .B(n11458), .Z(n23271) );
  AND U21347 ( .A(n11461), .B(n11460), .Z(n23269) );
  NAND U21348 ( .A(n11463), .B(n11462), .Z(n23267) );
  AND U21349 ( .A(n11465), .B(n11464), .Z(n23261) );
  AND U21350 ( .A(n11467), .B(n11466), .Z(n23255) );
  AND U21351 ( .A(n11469), .B(n11468), .Z(n23249) );
  AND U21352 ( .A(n11471), .B(n11470), .Z(n23243) );
  AND U21353 ( .A(n11473), .B(n11472), .Z(n23233) );
  NAND U21354 ( .A(n11475), .B(n11474), .Z(n23231) );
  AND U21355 ( .A(n11476), .B(n23907), .Z(n23222) );
  NAND U21356 ( .A(n11478), .B(n11477), .Z(n23216) );
  NANDN U21357 ( .A(x[3852]), .B(y[3852]), .Z(n23910) );
  NAND U21358 ( .A(n23910), .B(n11479), .Z(n23210) );
  ANDN U21359 ( .B(y[3850]), .A(x[3850]), .Z(n29281) );
  AND U21360 ( .A(n11481), .B(n11480), .Z(n23202) );
  AND U21361 ( .A(n29280), .B(n11482), .Z(n23200) );
  NAND U21362 ( .A(n11484), .B(n11483), .Z(n23198) );
  NANDN U21363 ( .A(x[3846]), .B(y[3846]), .Z(n23912) );
  AND U21364 ( .A(n23912), .B(n11485), .Z(n23196) );
  NAND U21365 ( .A(n11487), .B(n11486), .Z(n23188) );
  NAND U21366 ( .A(n11489), .B(n11488), .Z(n23183) );
  NAND U21367 ( .A(n11491), .B(n11490), .Z(n23177) );
  AND U21368 ( .A(n11493), .B(n11492), .Z(n23175) );
  NAND U21369 ( .A(n11495), .B(n11494), .Z(n23173) );
  AND U21370 ( .A(n11496), .B(n29266), .Z(n23164) );
  NAND U21371 ( .A(n11498), .B(n11497), .Z(n23162) );
  NANDN U21372 ( .A(x[3832]), .B(y[3832]), .Z(n23918) );
  AND U21373 ( .A(n11499), .B(n23918), .Z(n23160) );
  NANDN U21374 ( .A(x[3830]), .B(y[3830]), .Z(n29259) );
  NAND U21375 ( .A(n29259), .B(n29262), .Z(n23154) );
  ANDN U21376 ( .B(y[3828]), .A(x[3828]), .Z(n23919) );
  AND U21377 ( .A(n11501), .B(n11500), .Z(n23146) );
  AND U21378 ( .A(n23920), .B(n11502), .Z(n23144) );
  NAND U21379 ( .A(n11504), .B(n11503), .Z(n23142) );
  AND U21380 ( .A(n11506), .B(n11505), .Z(n23140) );
  AND U21381 ( .A(n11508), .B(n11507), .Z(n23134) );
  NANDN U21382 ( .A(x[3820]), .B(y[3820]), .Z(n29249) );
  AND U21383 ( .A(n29249), .B(n11509), .Z(n23128) );
  NAND U21384 ( .A(n11511), .B(n11510), .Z(n23126) );
  NAND U21385 ( .A(n11513), .B(n11512), .Z(n23122) );
  NAND U21386 ( .A(n11515), .B(n11514), .Z(n23117) );
  NAND U21387 ( .A(n11517), .B(n11516), .Z(n23112) );
  NANDN U21388 ( .A(x[3812]), .B(y[3812]), .Z(n29238) );
  AND U21389 ( .A(n29238), .B(n29240), .Z(n23110) );
  NANDN U21390 ( .A(x[3810]), .B(y[3810]), .Z(n29234) );
  NAND U21391 ( .A(n29234), .B(n29237), .Z(n23104) );
  NANDN U21392 ( .A(x[3808]), .B(y[3808]), .Z(n23923) );
  AND U21393 ( .A(n11519), .B(n11518), .Z(n23096) );
  NANDN U21394 ( .A(x[3806]), .B(y[3806]), .Z(n29230) );
  IV U21395 ( .A(n11520), .Z(n23922) );
  AND U21396 ( .A(n29230), .B(n23922), .Z(n23094) );
  NAND U21397 ( .A(n11522), .B(n11521), .Z(n23092) );
  AND U21398 ( .A(n11523), .B(n29229), .Z(n23090) );
  AND U21399 ( .A(n11525), .B(n11524), .Z(n23084) );
  AND U21400 ( .A(n11527), .B(n11526), .Z(n23078) );
  AND U21401 ( .A(n11529), .B(n11528), .Z(n23068) );
  AND U21402 ( .A(n11531), .B(n11530), .Z(n23062) );
  AND U21403 ( .A(n11533), .B(n11532), .Z(n23057) );
  AND U21404 ( .A(n11535), .B(n11534), .Z(n23053) );
  NAND U21405 ( .A(n29212), .B(n11536), .Z(n23051) );
  NANDN U21406 ( .A(x[3788]), .B(y[3788]), .Z(n29208) );
  NAND U21407 ( .A(n29208), .B(n11537), .Z(n23045) );
  NAND U21408 ( .A(n11538), .B(n29207), .Z(n23039) );
  AND U21409 ( .A(n11540), .B(n11539), .Z(n23025) );
  NANDN U21410 ( .A(x[3780]), .B(y[3780]), .Z(n29198) );
  AND U21411 ( .A(n29198), .B(n11541), .Z(n23019) );
  AND U21412 ( .A(n11542), .B(n29199), .Z(n23013) );
  NAND U21413 ( .A(n11544), .B(n11543), .Z(n23003) );
  NAND U21414 ( .A(n11546), .B(n11545), .Z(n22997) );
  NAND U21415 ( .A(n11548), .B(n11547), .Z(n22991) );
  AND U21416 ( .A(n11550), .B(n11549), .Z(n22989) );
  NAND U21417 ( .A(n11552), .B(n11551), .Z(n22987) );
  AND U21418 ( .A(n11554), .B(n11553), .Z(n22982) );
  NAND U21419 ( .A(n11555), .B(n29188), .Z(n22980) );
  AND U21420 ( .A(n11557), .B(n11556), .Z(n22978) );
  AND U21421 ( .A(n11559), .B(n11558), .Z(n22972) );
  AND U21422 ( .A(n11561), .B(n11560), .Z(n22966) );
  AND U21423 ( .A(n11563), .B(n11562), .Z(n22960) );
  AND U21424 ( .A(n11565), .B(n11564), .Z(n22954) );
  AND U21425 ( .A(n11567), .B(n11566), .Z(n22948) );
  AND U21426 ( .A(n11569), .B(n11568), .Z(n22942) );
  NANDN U21427 ( .A(x[3750]), .B(y[3750]), .Z(n23937) );
  NAND U21428 ( .A(n23937), .B(n11570), .Z(n22932) );
  IV U21429 ( .A(n11571), .Z(n23936) );
  NAND U21430 ( .A(n23936), .B(n11572), .Z(n22926) );
  ANDN U21431 ( .B(y[3746]), .A(x[3746]), .Z(n29168) );
  AND U21432 ( .A(n11574), .B(n11573), .Z(n22917) );
  AND U21433 ( .A(n29169), .B(n11575), .Z(n22915) );
  NAND U21434 ( .A(n11577), .B(n11576), .Z(n22913) );
  AND U21435 ( .A(n11579), .B(n11578), .Z(n22911) );
  AND U21436 ( .A(n11581), .B(n11580), .Z(n22905) );
  AND U21437 ( .A(n11583), .B(n11582), .Z(n22899) );
  NAND U21438 ( .A(n11585), .B(n11584), .Z(n22889) );
  NAND U21439 ( .A(n11587), .B(n11586), .Z(n22883) );
  NAND U21440 ( .A(n11589), .B(n11588), .Z(n22877) );
  NAND U21441 ( .A(n11591), .B(n11590), .Z(n22871) );
  AND U21442 ( .A(n11593), .B(n11592), .Z(n22869) );
  NAND U21443 ( .A(n11595), .B(n11594), .Z(n22867) );
  AND U21444 ( .A(n11596), .B(n29147), .Z(n22858) );
  AND U21445 ( .A(n11598), .B(n11597), .Z(n22856) );
  NAND U21446 ( .A(n11600), .B(n11599), .Z(n22854) );
  AND U21447 ( .A(n11602), .B(n11601), .Z(n22852) );
  NANDN U21448 ( .A(x[3720]), .B(y[3720]), .Z(n29141) );
  NAND U21449 ( .A(n29141), .B(n11603), .Z(n22850) );
  NAND U21450 ( .A(n11604), .B(n29140), .Z(n22844) );
  NAND U21451 ( .A(n11606), .B(n11605), .Z(n22838) );
  AND U21452 ( .A(n11608), .B(n11607), .Z(n22836) );
  NAND U21453 ( .A(n11610), .B(n11609), .Z(n22834) );
  AND U21454 ( .A(n11612), .B(n11611), .Z(n22828) );
  AND U21455 ( .A(n11614), .B(n11613), .Z(n22822) );
  AND U21456 ( .A(n11616), .B(n11615), .Z(n22816) );
  AND U21457 ( .A(n11618), .B(n11617), .Z(n22810) );
  NANDN U21458 ( .A(x[3704]), .B(y[3704]), .Z(n29125) );
  AND U21459 ( .A(n29125), .B(n11619), .Z(n22804) );
  IV U21460 ( .A(n11620), .Z(n29124) );
  AND U21461 ( .A(n11621), .B(n29124), .Z(n22798) );
  AND U21462 ( .A(n11623), .B(n11622), .Z(n22792) );
  AND U21463 ( .A(n11625), .B(n11624), .Z(n22786) );
  NANDN U21464 ( .A(x[3696]), .B(y[3696]), .Z(n29115) );
  AND U21465 ( .A(n29115), .B(n11626), .Z(n22780) );
  AND U21466 ( .A(n11627), .B(n29116), .Z(n22774) );
  NAND U21467 ( .A(n11629), .B(n11628), .Z(n22772) );
  AND U21468 ( .A(n11631), .B(n11630), .Z(n22766) );
  NAND U21469 ( .A(n11633), .B(n11632), .Z(n22760) );
  NAND U21470 ( .A(n11635), .B(n11634), .Z(n22754) );
  AND U21471 ( .A(n11637), .B(n11636), .Z(n22752) );
  NAND U21472 ( .A(n11639), .B(n11638), .Z(n22750) );
  NAND U21473 ( .A(n11640), .B(n23947), .Z(n22735) );
  NAND U21474 ( .A(n11642), .B(n11641), .Z(n22729) );
  NAND U21475 ( .A(n11644), .B(n11643), .Z(n22723) );
  AND U21476 ( .A(n11646), .B(n11645), .Z(n22721) );
  AND U21477 ( .A(n11648), .B(n11647), .Z(n22709) );
  AND U21478 ( .A(n11650), .B(n11649), .Z(n22704) );
  ANDN U21479 ( .B(y[3668]), .A(x[3668]), .Z(n29087) );
  NAND U21480 ( .A(n11652), .B(n11651), .Z(n22699) );
  NANDN U21481 ( .A(x[3666]), .B(y[3666]), .Z(n29085) );
  AND U21482 ( .A(n29085), .B(n29086), .Z(n22697) );
  AND U21483 ( .A(n11653), .B(n29084), .Z(n22691) );
  OR U21484 ( .A(n11655), .B(n11654), .Z(n11656) );
  AND U21485 ( .A(n11657), .B(n11656), .Z(n22687) );
  NAND U21486 ( .A(n29081), .B(n11658), .Z(n22685) );
  NAND U21487 ( .A(n11660), .B(n11659), .Z(n22679) );
  NAND U21488 ( .A(n11662), .B(n11661), .Z(n22673) );
  NAND U21489 ( .A(n11664), .B(n11663), .Z(n22667) );
  NAND U21490 ( .A(n11666), .B(n11665), .Z(n22661) );
  AND U21491 ( .A(n11667), .B(n23955), .Z(n22652) );
  AND U21492 ( .A(n11669), .B(n11668), .Z(n22650) );
  NAND U21493 ( .A(n11671), .B(n11670), .Z(n22648) );
  AND U21494 ( .A(n11673), .B(n11672), .Z(n22646) );
  AND U21495 ( .A(n11675), .B(n11674), .Z(n22640) );
  AND U21496 ( .A(n11677), .B(n11676), .Z(n22634) );
  AND U21497 ( .A(n11679), .B(n11678), .Z(n22628) );
  AND U21498 ( .A(n11681), .B(n11680), .Z(n22622) );
  NAND U21499 ( .A(n11683), .B(n11682), .Z(n22608) );
  NANDN U21500 ( .A(x[3634]), .B(y[3634]), .Z(n29056) );
  AND U21501 ( .A(n29056), .B(n11684), .Z(n22606) );
  NANDN U21502 ( .A(x[3632]), .B(y[3632]), .Z(n29050) );
  NAND U21503 ( .A(n29050), .B(n29055), .Z(n22600) );
  NAND U21504 ( .A(n29051), .B(n11685), .Z(n22594) );
  AND U21505 ( .A(n11687), .B(n11686), .Z(n22592) );
  NANDN U21506 ( .A(x[3628]), .B(y[3628]), .Z(n29046) );
  AND U21507 ( .A(n29046), .B(n11688), .Z(n22590) );
  NAND U21508 ( .A(n11690), .B(n11689), .Z(n22588) );
  AND U21509 ( .A(n11691), .B(n29045), .Z(n22586) );
  NAND U21510 ( .A(n11693), .B(n11692), .Z(n22584) );
  AND U21511 ( .A(n11695), .B(n11694), .Z(n22578) );
  AND U21512 ( .A(n11697), .B(n11696), .Z(n22573) );
  AND U21513 ( .A(n11699), .B(n11698), .Z(n22569) );
  AND U21514 ( .A(n11700), .B(n29036), .Z(n22567) );
  NAND U21515 ( .A(n11702), .B(n11701), .Z(n22565) );
  AND U21516 ( .A(n11704), .B(n11703), .Z(n22563) );
  NAND U21517 ( .A(n11706), .B(n11705), .Z(n22561) );
  AND U21518 ( .A(n11708), .B(n11707), .Z(n22559) );
  NAND U21519 ( .A(n11710), .B(n11709), .Z(n22557) );
  AND U21520 ( .A(n11712), .B(n11711), .Z(n22555) );
  NANDN U21521 ( .A(x[3610]), .B(y[3610]), .Z(n29025) );
  NAND U21522 ( .A(n29025), .B(n11713), .Z(n22549) );
  NANDN U21523 ( .A(x[3608]), .B(y[3608]), .Z(n29021) );
  NAND U21524 ( .A(n29021), .B(n29024), .Z(n22543) );
  AND U21525 ( .A(n11715), .B(n11714), .Z(n22541) );
  AND U21526 ( .A(n11717), .B(n11716), .Z(n22537) );
  NANDN U21527 ( .A(x[3604]), .B(y[3604]), .Z(n29016) );
  NAND U21528 ( .A(n23962), .B(n29016), .Z(n22535) );
  AND U21529 ( .A(n11719), .B(n11718), .Z(n22533) );
  AND U21530 ( .A(n11721), .B(n11720), .Z(n22528) );
  ANDN U21531 ( .B(y[3600]), .A(x[3600]), .Z(n23964) );
  NAND U21532 ( .A(n11723), .B(n11722), .Z(n22523) );
  AND U21533 ( .A(n11725), .B(n11724), .Z(n22518) );
  AND U21534 ( .A(n11727), .B(n11726), .Z(n22512) );
  AND U21535 ( .A(n11729), .B(n11728), .Z(n22506) );
  AND U21536 ( .A(n11731), .B(n11730), .Z(n22500) );
  AND U21537 ( .A(n11733), .B(n11732), .Z(n22494) );
  AND U21538 ( .A(n11735), .B(n11734), .Z(n22488) );
  AND U21539 ( .A(n11737), .B(n11736), .Z(n22474) );
  AND U21540 ( .A(n11739), .B(n11738), .Z(n22468) );
  AND U21541 ( .A(n11741), .B(n11740), .Z(n22462) );
  NAND U21542 ( .A(n11743), .B(n11742), .Z(n22442) );
  AND U21543 ( .A(n11745), .B(n11744), .Z(n22437) );
  AND U21544 ( .A(n11747), .B(n11746), .Z(n22431) );
  AND U21545 ( .A(n11749), .B(n11748), .Z(n22421) );
  NAND U21546 ( .A(n11751), .B(n11750), .Z(n22419) );
  AND U21547 ( .A(n11753), .B(n11752), .Z(n22417) );
  IV U21548 ( .A(n11754), .Z(n28973) );
  NAND U21549 ( .A(n11756), .B(n11755), .Z(n22398) );
  NAND U21550 ( .A(n11758), .B(n11757), .Z(n22392) );
  NAND U21551 ( .A(n11760), .B(n11759), .Z(n22386) );
  AND U21552 ( .A(n11762), .B(n11761), .Z(n22384) );
  NAND U21553 ( .A(n11764), .B(n11763), .Z(n22382) );
  AND U21554 ( .A(n11766), .B(n11765), .Z(n22376) );
  AND U21555 ( .A(n11768), .B(n11767), .Z(n22370) );
  AND U21556 ( .A(n11770), .B(n11769), .Z(n22364) );
  AND U21557 ( .A(n11772), .B(n11771), .Z(n22358) );
  AND U21558 ( .A(n11774), .B(n11773), .Z(n22352) );
  NAND U21559 ( .A(n11776), .B(n11775), .Z(n22350) );
  AND U21560 ( .A(n11778), .B(n11777), .Z(n22344) );
  AND U21561 ( .A(n11780), .B(n11779), .Z(n22339) );
  AND U21562 ( .A(n11781), .B(n23974), .Z(n22337) );
  NAND U21563 ( .A(n11783), .B(n11782), .Z(n22335) );
  AND U21564 ( .A(n11785), .B(n11784), .Z(n22330) );
  NANDN U21565 ( .A(x[3528]), .B(y[3528]), .Z(n23976) );
  NAND U21566 ( .A(n28944), .B(n23976), .Z(n22328) );
  IV U21567 ( .A(n11786), .Z(n23975) );
  NANDN U21568 ( .A(x[3526]), .B(y[3526]), .Z(n28939) );
  NAND U21569 ( .A(n23975), .B(n28939), .Z(n22322) );
  IV U21570 ( .A(n11787), .Z(n28938) );
  NANDN U21571 ( .A(x[3524]), .B(y[3524]), .Z(n28936) );
  NAND U21572 ( .A(n28938), .B(n28936), .Z(n22316) );
  AND U21573 ( .A(n11789), .B(n11788), .Z(n22314) );
  NANDN U21574 ( .A(x[3522]), .B(y[3522]), .Z(n28933) );
  IV U21575 ( .A(n11790), .Z(n28935) );
  AND U21576 ( .A(n28933), .B(n28935), .Z(n22312) );
  NAND U21577 ( .A(n11792), .B(n11791), .Z(n22310) );
  AND U21578 ( .A(n11794), .B(n11793), .Z(n22304) );
  ANDN U21579 ( .B(y[3518]), .A(x[3518]), .Z(n28931) );
  NAND U21580 ( .A(n11796), .B(n11795), .Z(n22299) );
  NAND U21581 ( .A(n11798), .B(n11797), .Z(n22294) );
  NANDN U21582 ( .A(x[3514]), .B(y[3514]), .Z(n23982) );
  NAND U21583 ( .A(n11800), .B(n11799), .Z(n22289) );
  AND U21584 ( .A(n11801), .B(n23981), .Z(n22287) );
  AND U21585 ( .A(n11803), .B(n11802), .Z(n22285) );
  NAND U21586 ( .A(n11805), .B(n11804), .Z(n22283) );
  AND U21587 ( .A(n11807), .B(n11806), .Z(n22281) );
  AND U21588 ( .A(n11809), .B(n11808), .Z(n22275) );
  AND U21589 ( .A(n11811), .B(n11810), .Z(n22269) );
  AND U21590 ( .A(n11813), .B(n11812), .Z(n22263) );
  AND U21591 ( .A(n11815), .B(n11814), .Z(n22257) );
  AND U21592 ( .A(n11817), .B(n11816), .Z(n22251) );
  AND U21593 ( .A(n11819), .B(n11818), .Z(n22245) );
  AND U21594 ( .A(n11821), .B(n11820), .Z(n22239) );
  AND U21595 ( .A(n11823), .B(n11822), .Z(n22233) );
  AND U21596 ( .A(n11825), .B(n11824), .Z(n22227) );
  NAND U21597 ( .A(n11827), .B(n11826), .Z(n22213) );
  NANDN U21598 ( .A(x[3486]), .B(y[3486]), .Z(n28903) );
  AND U21599 ( .A(n28903), .B(n11828), .Z(n22211) );
  NAND U21600 ( .A(n28902), .B(n11829), .Z(n22205) );
  NAND U21601 ( .A(n11831), .B(n11830), .Z(n22199) );
  AND U21602 ( .A(n11833), .B(n11832), .Z(n22197) );
  NAND U21603 ( .A(n11835), .B(n11834), .Z(n22195) );
  AND U21604 ( .A(n11837), .B(n11836), .Z(n22193) );
  NAND U21605 ( .A(n11839), .B(n11838), .Z(n22187) );
  NAND U21606 ( .A(n11841), .B(n11840), .Z(n22181) );
  NAND U21607 ( .A(n11843), .B(n11842), .Z(n22175) );
  NAND U21608 ( .A(n11845), .B(n11844), .Z(n22169) );
  NANDN U21609 ( .A(x[3470]), .B(y[3470]), .Z(n28888) );
  AND U21610 ( .A(n11846), .B(n23992), .Z(n22160) );
  AND U21611 ( .A(n11848), .B(n11847), .Z(n22158) );
  NAND U21612 ( .A(n11850), .B(n11849), .Z(n22156) );
  AND U21613 ( .A(n11852), .B(n11851), .Z(n22154) );
  AND U21614 ( .A(n11854), .B(n11853), .Z(n22148) );
  AND U21615 ( .A(n11856), .B(n11855), .Z(n22142) );
  NAND U21616 ( .A(n11858), .B(n11857), .Z(n22140) );
  IV U21617 ( .A(n11859), .Z(n28877) );
  IV U21618 ( .A(n11860), .Z(n28876) );
  IV U21619 ( .A(n11861), .Z(n28875) );
  AND U21620 ( .A(n11862), .B(n28875), .Z(n22128) );
  AND U21621 ( .A(n11864), .B(n11863), .Z(n22122) );
  AND U21622 ( .A(n11866), .B(n11865), .Z(n22120) );
  NAND U21623 ( .A(n11868), .B(n11867), .Z(n22118) );
  AND U21624 ( .A(n11869), .B(n23996), .Z(n22109) );
  AND U21625 ( .A(n11871), .B(n11870), .Z(n22107) );
  NAND U21626 ( .A(n11873), .B(n11872), .Z(n22105) );
  AND U21627 ( .A(n11875), .B(n11874), .Z(n22103) );
  AND U21628 ( .A(n11877), .B(n11876), .Z(n22097) );
  NAND U21629 ( .A(n11879), .B(n11878), .Z(n22087) );
  NAND U21630 ( .A(n11881), .B(n11880), .Z(n22081) );
  NAND U21631 ( .A(n11883), .B(n11882), .Z(n22075) );
  ANDN U21632 ( .B(y[3434]), .A(x[3434]), .Z(n28856) );
  AND U21633 ( .A(n11885), .B(n11884), .Z(n22066) );
  AND U21634 ( .A(n11886), .B(n24001), .Z(n22064) );
  NAND U21635 ( .A(n11888), .B(n11887), .Z(n22062) );
  AND U21636 ( .A(n11890), .B(n11889), .Z(n22060) );
  AND U21637 ( .A(n11892), .B(n11891), .Z(n22054) );
  AND U21638 ( .A(n11894), .B(n11893), .Z(n22048) );
  AND U21639 ( .A(n11896), .B(n11895), .Z(n22042) );
  AND U21640 ( .A(n11898), .B(n11897), .Z(n22036) );
  AND U21641 ( .A(n11900), .B(n11899), .Z(n22030) );
  AND U21642 ( .A(n11902), .B(n11901), .Z(n22024) );
  AND U21643 ( .A(n11904), .B(n11903), .Z(n22018) );
  AND U21644 ( .A(n11906), .B(n11905), .Z(n22012) );
  AND U21645 ( .A(n11908), .B(n11907), .Z(n22006) );
  AND U21646 ( .A(n11910), .B(n11909), .Z(n22000) );
  AND U21647 ( .A(n11912), .B(n11911), .Z(n21994) );
  NANDN U21648 ( .A(x[3406]), .B(y[3406]), .Z(n24010) );
  AND U21649 ( .A(n24010), .B(n11913), .Z(n21988) );
  AND U21650 ( .A(n11914), .B(n24009), .Z(n21982) );
  NAND U21651 ( .A(n11916), .B(n11915), .Z(n21980) );
  AND U21652 ( .A(n11918), .B(n11917), .Z(n21974) );
  AND U21653 ( .A(n11920), .B(n11919), .Z(n21969) );
  ANDN U21654 ( .B(y[3398]), .A(x[3398]), .Z(n24013) );
  AND U21655 ( .A(n11921), .B(n24014), .Z(n21961) );
  NAND U21656 ( .A(n11923), .B(n11922), .Z(n21942) );
  AND U21657 ( .A(n11925), .B(n11924), .Z(n21940) );
  AND U21658 ( .A(n11927), .B(n11926), .Z(n21934) );
  AND U21659 ( .A(n11929), .B(n11928), .Z(n21928) );
  AND U21660 ( .A(n11931), .B(n11930), .Z(n21922) );
  AND U21661 ( .A(n11933), .B(n11932), .Z(n21916) );
  AND U21662 ( .A(n11935), .B(n11934), .Z(n21910) );
  AND U21663 ( .A(n11937), .B(n11936), .Z(n21904) );
  AND U21664 ( .A(n11939), .B(n11938), .Z(n21898) );
  AND U21665 ( .A(n11941), .B(n11940), .Z(n21888) );
  AND U21666 ( .A(n11943), .B(n11942), .Z(n21882) );
  AND U21667 ( .A(n11945), .B(n11944), .Z(n21877) );
  AND U21668 ( .A(n11947), .B(n11946), .Z(n21873) );
  NAND U21669 ( .A(n11948), .B(n24025), .Z(n21871) );
  AND U21670 ( .A(n11950), .B(n11949), .Z(n21869) );
  AND U21671 ( .A(n11952), .B(n11951), .Z(n21863) );
  AND U21672 ( .A(n11954), .B(n11953), .Z(n21857) );
  AND U21673 ( .A(n11956), .B(n11955), .Z(n21847) );
  IV U21674 ( .A(n11957), .Z(n28785) );
  AND U21675 ( .A(n11958), .B(n28785), .Z(n21835) );
  AND U21676 ( .A(n11960), .B(n11959), .Z(n21833) );
  NAND U21677 ( .A(n11962), .B(n11961), .Z(n21831) );
  AND U21678 ( .A(n11964), .B(n11963), .Z(n21829) );
  AND U21679 ( .A(n11966), .B(n11965), .Z(n21823) );
  AND U21680 ( .A(n11968), .B(n11967), .Z(n21817) );
  AND U21681 ( .A(n11970), .B(n11969), .Z(n21811) );
  AND U21682 ( .A(n11972), .B(n11971), .Z(n21805) );
  AND U21683 ( .A(n11974), .B(n11973), .Z(n21791) );
  AND U21684 ( .A(n11976), .B(n11975), .Z(n21785) );
  AND U21685 ( .A(n11978), .B(n11977), .Z(n21779) );
  AND U21686 ( .A(n11980), .B(n11979), .Z(n21773) );
  AND U21687 ( .A(n11982), .B(n11981), .Z(n21767) );
  AND U21688 ( .A(n11984), .B(n11983), .Z(n21761) );
  NAND U21689 ( .A(n11986), .B(n11985), .Z(n21747) );
  AND U21690 ( .A(n11988), .B(n11987), .Z(n21745) );
  AND U21691 ( .A(n11990), .B(n11989), .Z(n21739) );
  AND U21692 ( .A(n11992), .B(n11991), .Z(n21734) );
  NAND U21693 ( .A(n11993), .B(n28756), .Z(n21732) );
  AND U21694 ( .A(n11994), .B(n28752), .Z(n21722) );
  AND U21695 ( .A(n11996), .B(n11995), .Z(n21716) );
  AND U21696 ( .A(n11998), .B(n11997), .Z(n21706) );
  NAND U21697 ( .A(n12000), .B(n11999), .Z(n21704) );
  AND U21698 ( .A(n12002), .B(n12001), .Z(n21702) );
  NAND U21699 ( .A(n12004), .B(n12003), .Z(n21700) );
  AND U21700 ( .A(n12005), .B(n24043), .Z(n21691) );
  AND U21701 ( .A(n12007), .B(n12006), .Z(n21689) );
  NAND U21702 ( .A(n12009), .B(n12008), .Z(n21687) );
  AND U21703 ( .A(n12011), .B(n12010), .Z(n21685) );
  AND U21704 ( .A(n12013), .B(n12012), .Z(n21679) );
  AND U21705 ( .A(n12015), .B(n12014), .Z(n21673) );
  NANDN U21706 ( .A(x[3290]), .B(y[3290]), .Z(n28733) );
  NAND U21707 ( .A(n28733), .B(n12016), .Z(n21663) );
  NAND U21708 ( .A(n24049), .B(n12017), .Z(n21657) );
  AND U21709 ( .A(n12019), .B(n12018), .Z(n21643) );
  AND U21710 ( .A(n12021), .B(n12020), .Z(n21637) );
  AND U21711 ( .A(n12023), .B(n12022), .Z(n21631) );
  AND U21712 ( .A(n12025), .B(n12024), .Z(n21617) );
  AND U21713 ( .A(n12027), .B(n12026), .Z(n21611) );
  AND U21714 ( .A(n12029), .B(n12028), .Z(n21605) );
  AND U21715 ( .A(n12031), .B(n12030), .Z(n21599) );
  AND U21716 ( .A(n12033), .B(n12032), .Z(n21593) );
  AND U21717 ( .A(n12035), .B(n12034), .Z(n21587) );
  AND U21718 ( .A(n12037), .B(n12036), .Z(n21581) );
  AND U21719 ( .A(n12039), .B(n12038), .Z(n21575) );
  AND U21720 ( .A(n12041), .B(n12040), .Z(n21569) );
  AND U21721 ( .A(n12043), .B(n12042), .Z(n21563) );
  NANDN U21722 ( .A(x[3256]), .B(y[3256]), .Z(n28704) );
  AND U21723 ( .A(n28704), .B(n12044), .Z(n21557) );
  AND U21724 ( .A(n12045), .B(n28703), .Z(n21551) );
  AND U21725 ( .A(n12047), .B(n12046), .Z(n21545) );
  AND U21726 ( .A(n12049), .B(n12048), .Z(n21539) );
  AND U21727 ( .A(n12051), .B(n12050), .Z(n21525) );
  AND U21728 ( .A(n12053), .B(n12052), .Z(n21519) );
  AND U21729 ( .A(n12055), .B(n12054), .Z(n21513) );
  AND U21730 ( .A(n12057), .B(n12056), .Z(n21507) );
  AND U21731 ( .A(n12059), .B(n12058), .Z(n21501) );
  AND U21732 ( .A(n12061), .B(n12060), .Z(n21495) );
  AND U21733 ( .A(n12063), .B(n12062), .Z(n21489) );
  AND U21734 ( .A(n12065), .B(n12064), .Z(n21483) );
  AND U21735 ( .A(n12067), .B(n12066), .Z(n21477) );
  AND U21736 ( .A(n12069), .B(n12068), .Z(n21471) );
  AND U21737 ( .A(n12071), .B(n12070), .Z(n21465) );
  AND U21738 ( .A(n12073), .B(n12072), .Z(n21459) );
  NAND U21739 ( .A(n12075), .B(n12074), .Z(n21449) );
  NAND U21740 ( .A(n12077), .B(n12076), .Z(n21443) );
  NAND U21741 ( .A(n12079), .B(n12078), .Z(n21437) );
  AND U21742 ( .A(n12081), .B(n12080), .Z(n21435) );
  NAND U21743 ( .A(n12083), .B(n12082), .Z(n21433) );
  AND U21744 ( .A(n12085), .B(n12084), .Z(n21427) );
  AND U21745 ( .A(n12087), .B(n12086), .Z(n21421) );
  AND U21746 ( .A(n12089), .B(n12088), .Z(n21411) );
  AND U21747 ( .A(n12091), .B(n12090), .Z(n21405) );
  NAND U21748 ( .A(n12093), .B(n12092), .Z(n21399) );
  NAND U21749 ( .A(n12095), .B(n12094), .Z(n21393) );
  NAND U21750 ( .A(n12097), .B(n12096), .Z(n21387) );
  AND U21751 ( .A(n12099), .B(n12098), .Z(n21385) );
  NAND U21752 ( .A(n12101), .B(n12100), .Z(n21383) );
  AND U21753 ( .A(n12103), .B(n12102), .Z(n21377) );
  AND U21754 ( .A(n12105), .B(n12104), .Z(n21371) );
  AND U21755 ( .A(n12107), .B(n12106), .Z(n21365) );
  AND U21756 ( .A(n12109), .B(n12108), .Z(n21359) );
  AND U21757 ( .A(n12111), .B(n12110), .Z(n21353) );
  AND U21758 ( .A(n12113), .B(n12112), .Z(n21347) );
  AND U21759 ( .A(n12115), .B(n12114), .Z(n21341) );
  AND U21760 ( .A(n12117), .B(n12116), .Z(n21335) );
  AND U21761 ( .A(n12119), .B(n12118), .Z(n21329) );
  AND U21762 ( .A(n12121), .B(n12120), .Z(n21323) );
  AND U21763 ( .A(n12123), .B(n12122), .Z(n21317) );
  AND U21764 ( .A(n12125), .B(n12124), .Z(n21311) );
  NAND U21765 ( .A(n12127), .B(n12126), .Z(n21301) );
  NAND U21766 ( .A(n12129), .B(n12128), .Z(n21295) );
  NAND U21767 ( .A(n12131), .B(n12130), .Z(n21289) );
  AND U21768 ( .A(n12133), .B(n12132), .Z(n21275) );
  AND U21769 ( .A(n12135), .B(n12134), .Z(n21265) );
  AND U21770 ( .A(n12137), .B(n12136), .Z(n21243) );
  ANDN U21771 ( .B(n12139), .A(n12138), .Z(n21233) );
  AND U21772 ( .A(n12140), .B(n28607), .Z(n21205) );
  AND U21773 ( .A(n12142), .B(n12141), .Z(n21195) );
  AND U21774 ( .A(n12144), .B(n12143), .Z(n21173) );
  AND U21775 ( .A(n12146), .B(n12145), .Z(n21151) );
  AND U21776 ( .A(n12148), .B(n12147), .Z(n21129) );
  AND U21777 ( .A(n12150), .B(n12149), .Z(n21107) );
  AND U21778 ( .A(n12152), .B(n12151), .Z(n21085) );
  AND U21779 ( .A(n12154), .B(n12153), .Z(n21063) );
  AND U21780 ( .A(n12156), .B(n12155), .Z(n21041) );
  OR U21781 ( .A(n12158), .B(n12157), .Z(n12159) );
  AND U21782 ( .A(n12160), .B(n12159), .Z(n21025) );
  IV U21783 ( .A(n12161), .Z(n28561) );
  AND U21784 ( .A(n12162), .B(n28561), .Z(n21023) );
  XNOR U21785 ( .A(y[3087]), .B(x[3087]), .Z(n21012) );
  NANDN U21786 ( .A(x[3078]), .B(y[3078]), .Z(n28546) );
  NAND U21787 ( .A(n28546), .B(n12163), .Z(n20993) );
  AND U21788 ( .A(n12167), .B(n12166), .Z(n20984) );
  NAND U21789 ( .A(n12169), .B(n12168), .Z(n20982) );
  AND U21790 ( .A(n12171), .B(n12170), .Z(n20980) );
  AND U21791 ( .A(n12172), .B(n28536), .Z(n20974) );
  AND U21792 ( .A(n12176), .B(n12175), .Z(n20950) );
  AND U21793 ( .A(n12180), .B(n12179), .Z(n20941) );
  AND U21794 ( .A(n12182), .B(n12181), .Z(n20931) );
  NAND U21795 ( .A(n12184), .B(n12183), .Z(n20929) );
  AND U21796 ( .A(n12186), .B(n12185), .Z(n20927) );
  AND U21797 ( .A(n12188), .B(n12187), .Z(n28515) );
  XNOR U21798 ( .A(x[3040]), .B(y[3040]), .Z(n20904) );
  NAND U21799 ( .A(n12190), .B(n12189), .Z(n24104) );
  AND U21800 ( .A(n12191), .B(n24104), .Z(n20902) );
  NAND U21801 ( .A(n24105), .B(n12192), .Z(n20900) );
  IV U21802 ( .A(n12193), .Z(n28505) );
  AND U21803 ( .A(n12194), .B(n28505), .Z(n20898) );
  AND U21804 ( .A(n12196), .B(n12195), .Z(n20887) );
  NAND U21805 ( .A(n28500), .B(n12197), .Z(n20885) );
  AND U21806 ( .A(n12199), .B(n12198), .Z(n20883) );
  NAND U21807 ( .A(n12201), .B(n12200), .Z(n20881) );
  AND U21808 ( .A(n12203), .B(n12202), .Z(n20879) );
  NAND U21809 ( .A(n12205), .B(n12204), .Z(n20877) );
  AND U21810 ( .A(n12207), .B(n12206), .Z(n20875) );
  AND U21811 ( .A(n12209), .B(n12208), .Z(n28492) );
  AND U21812 ( .A(n28488), .B(n12210), .Z(n20858) );
  NAND U21813 ( .A(n28483), .B(n12211), .Z(n20848) );
  AND U21814 ( .A(n12213), .B(n28480), .Z(n20842) );
  IV U21815 ( .A(n12214), .Z(n28479) );
  NAND U21816 ( .A(n28479), .B(n28478), .Z(n20840) );
  NANDN U21817 ( .A(x[3012]), .B(y[3012]), .Z(n24112) );
  NAND U21818 ( .A(n12218), .B(n12217), .Z(n28474) );
  AND U21819 ( .A(n12220), .B(n12219), .Z(n24113) );
  AND U21820 ( .A(n12223), .B(n28469), .Z(n20819) );
  NAND U21821 ( .A(n28468), .B(n28466), .Z(n20817) );
  AND U21822 ( .A(n28465), .B(n12224), .Z(n20815) );
  NAND U21823 ( .A(n12226), .B(n12225), .Z(n28464) );
  AND U21824 ( .A(n12230), .B(n24115), .Z(n20796) );
  AND U21825 ( .A(n12234), .B(n12233), .Z(n20785) );
  AND U21826 ( .A(n12236), .B(n12235), .Z(n20779) );
  AND U21827 ( .A(n12238), .B(n12237), .Z(n20773) );
  OR U21828 ( .A(n12240), .B(n12239), .Z(n12242) );
  AND U21829 ( .A(n12242), .B(n12241), .Z(n28447) );
  OR U21830 ( .A(n28443), .B(n12244), .Z(n20758) );
  OR U21831 ( .A(n12246), .B(n12245), .Z(n12247) );
  AND U21832 ( .A(n12248), .B(n12247), .Z(n28440) );
  IV U21833 ( .A(n12249), .Z(n28439) );
  AND U21834 ( .A(n12250), .B(n28439), .Z(n20750) );
  IV U21835 ( .A(n12251), .Z(n28438) );
  NOR U21836 ( .A(n28438), .B(n12252), .Z(n20748) );
  AND U21837 ( .A(n28434), .B(n12253), .Z(n20743) );
  AND U21838 ( .A(n12256), .B(n28430), .Z(n20740) );
  NAND U21839 ( .A(n28431), .B(n12257), .Z(n28429) );
  NANDN U21840 ( .A(x[2964]), .B(y[2964]), .Z(n28428) );
  IV U21841 ( .A(n12258), .Z(n28425) );
  NANDN U21842 ( .A(n28425), .B(n12259), .Z(n12261) );
  ANDN U21843 ( .B(n12261), .A(n12260), .Z(n20730) );
  AND U21844 ( .A(n12262), .B(n24126), .Z(n20721) );
  AND U21845 ( .A(n12264), .B(n12263), .Z(n28421) );
  NAND U21846 ( .A(n28420), .B(n12265), .Z(n20715) );
  NOR U21847 ( .A(n12266), .B(n28419), .Z(n20713) );
  NAND U21848 ( .A(n12268), .B(n12267), .Z(n28415) );
  AND U21849 ( .A(n12269), .B(n28411), .Z(n20696) );
  NANDN U21850 ( .A(n28407), .B(n12272), .Z(n12274) );
  ANDN U21851 ( .B(n12274), .A(n12273), .Z(n20684) );
  AND U21852 ( .A(n12276), .B(n12275), .Z(n20679) );
  NAND U21853 ( .A(n12278), .B(n12277), .Z(n20677) );
  AND U21854 ( .A(n12280), .B(n12279), .Z(n20675) );
  AND U21855 ( .A(n12282), .B(n12281), .Z(n20669) );
  AND U21856 ( .A(n12284), .B(n12283), .Z(n24135) );
  IV U21857 ( .A(n12285), .Z(n28398) );
  AND U21858 ( .A(n28396), .B(n28398), .Z(n20656) );
  NAND U21859 ( .A(n12287), .B(n12286), .Z(n20654) );
  AND U21860 ( .A(n28395), .B(n28393), .Z(n20652) );
  AND U21861 ( .A(n12289), .B(n12288), .Z(n28390) );
  ANDN U21862 ( .B(y[2924]), .A(x[2924]), .Z(n28386) );
  AND U21863 ( .A(n12291), .B(n12290), .Z(n28385) );
  IV U21864 ( .A(n12292), .Z(n28384) );
  AND U21865 ( .A(n12294), .B(n12293), .Z(n28380) );
  ANDN U21866 ( .B(n12296), .A(n12295), .Z(n28379) );
  NAND U21867 ( .A(n12300), .B(n12299), .Z(n12301) );
  NAND U21868 ( .A(n12302), .B(n12301), .Z(n24141) );
  IV U21869 ( .A(n12303), .Z(n28373) );
  ANDN U21870 ( .B(n28373), .A(n12304), .Z(n28371) );
  AND U21871 ( .A(n12306), .B(n12305), .Z(n20615) );
  IV U21872 ( .A(n12309), .Z(n28359) );
  NANDN U21873 ( .A(x[2902]), .B(y[2902]), .Z(n28358) );
  IV U21874 ( .A(n12312), .Z(n28356) );
  AND U21875 ( .A(n12313), .B(n28356), .Z(n20595) );
  NAND U21876 ( .A(n24143), .B(n28355), .Z(n20593) );
  AND U21877 ( .A(n28352), .B(n12316), .Z(n20587) );
  NOR U21878 ( .A(n12318), .B(n12317), .Z(n20578) );
  IV U21879 ( .A(n12319), .Z(n28346) );
  AND U21880 ( .A(n12320), .B(n28346), .Z(n20572) );
  NAND U21881 ( .A(n12322), .B(n12321), .Z(n28345) );
  IV U21882 ( .A(n12323), .Z(n28343) );
  NANDN U21883 ( .A(n28343), .B(n12324), .Z(n12326) );
  ANDN U21884 ( .B(n12326), .A(n12325), .Z(n20568) );
  IV U21885 ( .A(n12327), .Z(n28340) );
  NANDN U21886 ( .A(x[2884]), .B(y[2884]), .Z(n12329) );
  NAND U21887 ( .A(n12329), .B(n12328), .Z(n28338) );
  ANDN U21888 ( .B(y[2880]), .A(x[2880]), .Z(n28332) );
  AND U21889 ( .A(n12335), .B(n12334), .Z(n20537) );
  NAND U21890 ( .A(n12337), .B(n12336), .Z(n20535) );
  AND U21891 ( .A(n12339), .B(n12338), .Z(n20533) );
  AND U21892 ( .A(n12341), .B(n12340), .Z(n20527) );
  AND U21893 ( .A(n28320), .B(n12342), .Z(n20521) );
  NAND U21894 ( .A(n12344), .B(n12343), .Z(n28319) );
  AND U21895 ( .A(n12345), .B(n28318), .Z(n20518) );
  AND U21896 ( .A(n12347), .B(n12346), .Z(n20513) );
  AND U21897 ( .A(n12348), .B(n24150), .Z(n20508) );
  NAND U21898 ( .A(n12354), .B(n12353), .Z(n28308) );
  IV U21899 ( .A(n12358), .Z(n28305) );
  AND U21900 ( .A(n12359), .B(n28305), .Z(n20498) );
  IV U21901 ( .A(n12360), .Z(n28304) );
  NAND U21902 ( .A(n12362), .B(n12361), .Z(n20485) );
  AND U21903 ( .A(n12364), .B(n12363), .Z(n20483) );
  NAND U21904 ( .A(n28298), .B(n12365), .Z(n20481) );
  AND U21905 ( .A(n28297), .B(n12366), .Z(n20479) );
  AND U21906 ( .A(n12367), .B(n28292), .Z(n20473) );
  AND U21907 ( .A(n12369), .B(n12368), .Z(n20468) );
  NANDN U21908 ( .A(x[2840]), .B(y[2840]), .Z(n12371) );
  NAND U21909 ( .A(n12371), .B(n12370), .Z(n28279) );
  NAND U21910 ( .A(n28274), .B(n12374), .Z(n20456) );
  AND U21911 ( .A(n28269), .B(n28273), .Z(n20454) );
  NAND U21912 ( .A(n12377), .B(n28259), .Z(n20448) );
  AND U21913 ( .A(n28261), .B(n12378), .Z(n28257) );
  NAND U21914 ( .A(n12382), .B(n12381), .Z(n24152) );
  AND U21915 ( .A(n28249), .B(n12383), .Z(n20431) );
  AND U21916 ( .A(n12385), .B(n12384), .Z(n20428) );
  AND U21917 ( .A(n12387), .B(n12386), .Z(n20423) );
  AND U21918 ( .A(n28240), .B(n12388), .Z(n20418) );
  IV U21919 ( .A(n12390), .Z(n28234) );
  NAND U21920 ( .A(n28234), .B(n12391), .Z(n20407) );
  AND U21921 ( .A(n12394), .B(n28230), .Z(n24156) );
  AND U21922 ( .A(n12396), .B(n12395), .Z(n24155) );
  NAND U21923 ( .A(n12398), .B(n12397), .Z(n20396) );
  AND U21924 ( .A(n12399), .B(n28227), .Z(n20394) );
  NAND U21925 ( .A(n24158), .B(n12400), .Z(n20380) );
  IV U21926 ( .A(n12403), .Z(n28215) );
  NANDN U21927 ( .A(x[2792]), .B(y[2792]), .Z(n24164) );
  AND U21928 ( .A(n12406), .B(n24164), .Z(n20353) );
  AND U21929 ( .A(n12408), .B(n12407), .Z(n28208) );
  NANDN U21930 ( .A(x[2788]), .B(y[2788]), .Z(n28205) );
  NAND U21931 ( .A(n28205), .B(n12409), .Z(n20345) );
  AND U21932 ( .A(n12413), .B(n12412), .Z(n20336) );
  AND U21933 ( .A(n12415), .B(n12414), .Z(n20330) );
  NAND U21934 ( .A(n12417), .B(n12416), .Z(n12418) );
  NAND U21935 ( .A(n12419), .B(n12418), .Z(n20317) );
  AND U21936 ( .A(n12423), .B(n28185), .Z(n20305) );
  IV U21937 ( .A(n12426), .Z(n28180) );
  NAND U21938 ( .A(n28180), .B(n12427), .Z(n20299) );
  AND U21939 ( .A(n12428), .B(n24170), .Z(n20297) );
  OR U21940 ( .A(n12430), .B(n12429), .Z(n12431) );
  AND U21941 ( .A(n12432), .B(n12431), .Z(n28172) );
  AND U21942 ( .A(n12436), .B(n12435), .Z(n28169) );
  NAND U21943 ( .A(n28165), .B(n12440), .Z(n20264) );
  AND U21944 ( .A(n28162), .B(n28164), .Z(n20262) );
  NAND U21945 ( .A(n12443), .B(n28159), .Z(n20256) );
  NAND U21946 ( .A(n24178), .B(n12449), .Z(n20238) );
  AND U21947 ( .A(n28148), .B(n28146), .Z(n20231) );
  NAND U21948 ( .A(n12453), .B(n12452), .Z(n20229) );
  AND U21949 ( .A(n24180), .B(n28145), .Z(n20227) );
  IV U21950 ( .A(n12456), .Z(n28140) );
  NOR U21951 ( .A(n28133), .B(n12457), .Z(n20194) );
  AND U21952 ( .A(n12459), .B(n12458), .Z(n20188) );
  IV U21953 ( .A(n12460), .Z(n28124) );
  NAND U21954 ( .A(n12464), .B(n12463), .Z(n12465) );
  ANDN U21955 ( .B(n12465), .A(n20171), .Z(n12466) );
  NANDN U21956 ( .A(n12467), .B(n12466), .Z(n24186) );
  AND U21957 ( .A(n12469), .B(n12468), .Z(n24187) );
  AND U21958 ( .A(n12472), .B(n24188), .Z(n28116) );
  ANDN U21959 ( .B(y[2704]), .A(x[2704]), .Z(n28115) );
  IV U21960 ( .A(n12475), .Z(n24195) );
  AND U21961 ( .A(n12476), .B(n24195), .Z(n20157) );
  NAND U21962 ( .A(n24193), .B(n12477), .Z(n28113) );
  IV U21963 ( .A(n12480), .Z(n28110) );
  AND U21964 ( .A(n12481), .B(n28110), .Z(n20150) );
  IV U21965 ( .A(n12482), .Z(n28109) );
  AND U21966 ( .A(n12484), .B(n12483), .Z(n20141) );
  IV U21967 ( .A(n12485), .Z(n28104) );
  NAND U21968 ( .A(n28104), .B(n12486), .Z(n20139) );
  AND U21969 ( .A(n28103), .B(n12487), .Z(n20137) );
  AND U21970 ( .A(n12489), .B(n12488), .Z(n28102) );
  NOR U21971 ( .A(n12490), .B(n28101), .Z(n20134) );
  ANDN U21972 ( .B(n12491), .A(n28096), .Z(n20128) );
  AND U21973 ( .A(n12492), .B(n28095), .Z(n20126) );
  NAND U21974 ( .A(n12494), .B(n12493), .Z(n24197) );
  XNOR U21975 ( .A(x[2686]), .B(y[2686]), .Z(n12495) );
  AND U21976 ( .A(n12496), .B(n12495), .Z(n24198) );
  AND U21977 ( .A(n12500), .B(n12499), .Z(n28093) );
  AND U21978 ( .A(n12504), .B(n12503), .Z(n20098) );
  NAND U21979 ( .A(n12506), .B(n12505), .Z(n20088) );
  AND U21980 ( .A(n12510), .B(n12509), .Z(n20075) );
  AND U21981 ( .A(n28071), .B(n12511), .Z(n20069) );
  NANDN U21982 ( .A(x[2664]), .B(y[2664]), .Z(n12513) );
  NAND U21983 ( .A(n12513), .B(n12512), .Z(n28070) );
  IV U21984 ( .A(n12516), .Z(n28068) );
  AND U21985 ( .A(n28067), .B(n28065), .Z(n20062) );
  NANDN U21986 ( .A(x[2660]), .B(y[2660]), .Z(n24200) );
  NAND U21987 ( .A(n24200), .B(n12517), .Z(n20060) );
  NAND U21988 ( .A(n28059), .B(n12520), .Z(n20051) );
  NAND U21989 ( .A(n12524), .B(n12523), .Z(n28057) );
  IV U21990 ( .A(n12532), .Z(n28047) );
  NAND U21991 ( .A(n12537), .B(n12536), .Z(n28045) );
  AND U21992 ( .A(n12540), .B(n28038), .Z(n20026) );
  AND U21993 ( .A(n12543), .B(n12542), .Z(n28034) );
  IV U21994 ( .A(n12544), .Z(n28033) );
  NAND U21995 ( .A(n28033), .B(n12545), .Z(n20012) );
  XNOR U21996 ( .A(y[2624]), .B(x[2624]), .Z(n19993) );
  AND U21997 ( .A(n12547), .B(n12546), .Z(n28015) );
  IV U21998 ( .A(n12548), .Z(n28010) );
  NOR U21999 ( .A(n28010), .B(n12549), .Z(n19976) );
  IV U22000 ( .A(n12552), .Z(n28003) );
  NAND U22001 ( .A(n28003), .B(n12553), .Z(n19970) );
  AND U22002 ( .A(n12554), .B(n28005), .Z(n24209) );
  AND U22003 ( .A(n12556), .B(n12555), .Z(n24208) );
  NAND U22004 ( .A(n12558), .B(n12557), .Z(n19962) );
  AND U22005 ( .A(n12559), .B(n28001), .Z(n19960) );
  NOR U22006 ( .A(n24211), .B(n12560), .Z(n19947) );
  XNOR U22007 ( .A(y[2602]), .B(x[2602]), .Z(n19935) );
  AND U22008 ( .A(n12564), .B(n12563), .Z(n19923) );
  IV U22009 ( .A(n12565), .Z(n27987) );
  NAND U22010 ( .A(n27987), .B(n12566), .Z(n19914) );
  AND U22011 ( .A(n12568), .B(n12567), .Z(n27986) );
  AND U22012 ( .A(n12570), .B(n12569), .Z(n19904) );
  NAND U22013 ( .A(n12572), .B(n12571), .Z(n19902) );
  AND U22014 ( .A(n12574), .B(n12573), .Z(n19900) );
  AND U22015 ( .A(n12576), .B(n12575), .Z(n19894) );
  NANDN U22016 ( .A(x[2576]), .B(y[2576]), .Z(n12583) );
  NAND U22017 ( .A(n12583), .B(n12582), .Z(n27973) );
  NAND U22018 ( .A(n12587), .B(n12586), .Z(n27971) );
  IV U22019 ( .A(n12588), .Z(n27970) );
  AND U22020 ( .A(n27967), .B(n27970), .Z(n19867) );
  NAND U22021 ( .A(n12595), .B(n12594), .Z(n27961) );
  AND U22022 ( .A(n12600), .B(n27956), .Z(n27955) );
  AND U22023 ( .A(n12602), .B(n12601), .Z(n27953) );
  IV U22024 ( .A(n12603), .Z(n27951) );
  AND U22025 ( .A(n27950), .B(n12604), .Z(n19841) );
  NAND U22026 ( .A(n27945), .B(n12605), .Z(n19832) );
  NANDN U22027 ( .A(x[2554]), .B(y[2554]), .Z(n12607) );
  AND U22028 ( .A(n12607), .B(n12606), .Z(n27944) );
  AND U22029 ( .A(n12610), .B(n27940), .Z(n19828) );
  NAND U22030 ( .A(n27941), .B(n12611), .Z(n27939) );
  IV U22031 ( .A(n12612), .Z(n27938) );
  IV U22032 ( .A(n12613), .Z(n27936) );
  AND U22033 ( .A(n12614), .B(n27936), .Z(n19819) );
  IV U22034 ( .A(n12615), .Z(n27935) );
  NAND U22035 ( .A(n12617), .B(n12616), .Z(n19806) );
  AND U22036 ( .A(n12619), .B(n12618), .Z(n19804) );
  NAND U22037 ( .A(n27928), .B(n12620), .Z(n19802) );
  AND U22038 ( .A(n12622), .B(n12621), .Z(n19800) );
  NAND U22039 ( .A(n12624), .B(n12623), .Z(n12625) );
  NAND U22040 ( .A(n12626), .B(n12625), .Z(n24228) );
  NAND U22041 ( .A(n12628), .B(n12627), .Z(n19775) );
  AND U22042 ( .A(n12630), .B(n12629), .Z(n19773) );
  NAND U22043 ( .A(n12632), .B(n12631), .Z(n19771) );
  AND U22044 ( .A(n27915), .B(n12633), .Z(n19769) );
  IV U22045 ( .A(n12634), .Z(n24232) );
  AND U22046 ( .A(n12635), .B(n24232), .Z(n27913) );
  NANDN U22047 ( .A(x[2524]), .B(y[2524]), .Z(n24233) );
  NAND U22048 ( .A(n24233), .B(n12636), .Z(n19760) );
  IV U22049 ( .A(n12639), .Z(n27909) );
  IV U22050 ( .A(n12640), .Z(n27908) );
  AND U22051 ( .A(n12645), .B(n12644), .Z(n19738) );
  AND U22052 ( .A(n27900), .B(n12646), .Z(n19733) );
  AND U22053 ( .A(n12647), .B(n27898), .Z(n19728) );
  XNOR U22054 ( .A(x[2502]), .B(y[2502]), .Z(n19711) );
  AND U22055 ( .A(n12651), .B(n12650), .Z(n27882) );
  IV U22056 ( .A(n12652), .Z(n27880) );
  AND U22057 ( .A(n12653), .B(n27880), .Z(n19691) );
  IV U22058 ( .A(n12654), .Z(n27879) );
  NAND U22059 ( .A(n27879), .B(n27877), .Z(n19689) );
  AND U22060 ( .A(n12656), .B(n12655), .Z(n19687) );
  NAND U22061 ( .A(n27874), .B(n27876), .Z(n19685) );
  NAND U22062 ( .A(n27871), .B(n12659), .Z(n19678) );
  IV U22063 ( .A(n12660), .Z(n27870) );
  AND U22064 ( .A(n12661), .B(n27870), .Z(n19676) );
  AND U22065 ( .A(n12665), .B(n12664), .Z(n27864) );
  AND U22066 ( .A(n27859), .B(n27861), .Z(n19665) );
  NAND U22067 ( .A(n27851), .B(n12670), .Z(n19657) );
  AND U22068 ( .A(n12672), .B(n12671), .Z(n27848) );
  IV U22069 ( .A(n12673), .Z(n27846) );
  AND U22070 ( .A(n12675), .B(n12674), .Z(n27844) );
  IV U22071 ( .A(n12676), .Z(n27843) );
  IV U22072 ( .A(n12677), .Z(n27842) );
  IV U22073 ( .A(n12678), .Z(n27840) );
  AND U22074 ( .A(n27839), .B(n12679), .Z(n19637) );
  AND U22075 ( .A(n12682), .B(n24239), .Z(n27835) );
  NAND U22076 ( .A(n27832), .B(n12685), .Z(n19625) );
  IV U22077 ( .A(n12686), .Z(n27831) );
  AND U22078 ( .A(n12687), .B(n27831), .Z(n19623) );
  AND U22079 ( .A(n12689), .B(n12688), .Z(n19617) );
  NAND U22080 ( .A(n12691), .B(n12690), .Z(n19608) );
  NAND U22081 ( .A(n12696), .B(n12695), .Z(n27816) );
  NAND U22082 ( .A(n12700), .B(n12699), .Z(n27814) );
  IV U22083 ( .A(n12701), .Z(n27813) );
  AND U22084 ( .A(n12706), .B(n27811), .Z(n19575) );
  IV U22085 ( .A(n12707), .Z(n27807) );
  IV U22086 ( .A(n12708), .Z(n27806) );
  AND U22087 ( .A(n12709), .B(n27806), .Z(n19571) );
  IV U22088 ( .A(n12712), .Z(n27804) );
  AND U22089 ( .A(n12713), .B(n27804), .Z(n19568) );
  IV U22090 ( .A(n12714), .Z(n27803) );
  AND U22091 ( .A(n12716), .B(n12715), .Z(n19563) );
  NAND U22092 ( .A(n12721), .B(n12720), .Z(n19533) );
  AND U22093 ( .A(n12723), .B(n12722), .Z(n27774) );
  IV U22094 ( .A(n12724), .Z(n27767) );
  NAND U22095 ( .A(n12726), .B(n12725), .Z(n19501) );
  AND U22096 ( .A(n12728), .B(n12727), .Z(n19499) );
  NAND U22097 ( .A(n12730), .B(n12729), .Z(n19497) );
  AND U22098 ( .A(n12732), .B(n12731), .Z(n19495) );
  NAND U22099 ( .A(n12734), .B(n12733), .Z(n19488) );
  NAND U22100 ( .A(n27749), .B(n12737), .Z(n19472) );
  AND U22101 ( .A(n12739), .B(n12738), .Z(n27748) );
  AND U22102 ( .A(n12741), .B(n12740), .Z(n24254) );
  AND U22103 ( .A(n12746), .B(n27739), .Z(n19455) );
  IV U22104 ( .A(n12747), .Z(n27733) );
  NAND U22105 ( .A(n12763), .B(n12762), .Z(n27708) );
  NAND U22106 ( .A(n12765), .B(n12764), .Z(n27706) );
  NAND U22107 ( .A(n12769), .B(n12768), .Z(n27702) );
  NOR U22108 ( .A(n12773), .B(n12772), .Z(n19401) );
  IV U22109 ( .A(n12774), .Z(n27685) );
  AND U22110 ( .A(n12775), .B(n27685), .Z(n19395) );
  NAND U22111 ( .A(n12777), .B(n12776), .Z(n27684) );
  ANDN U22112 ( .B(y[2330]), .A(x[2330]), .Z(n27672) );
  AND U22113 ( .A(n12782), .B(n12781), .Z(n27671) );
  IV U22114 ( .A(n12783), .Z(n27668) );
  AND U22115 ( .A(n12784), .B(n27668), .Z(n19373) );
  AND U22116 ( .A(n12785), .B(n27667), .Z(n19371) );
  NAND U22117 ( .A(n12787), .B(n12786), .Z(n19369) );
  AND U22118 ( .A(n12789), .B(n12788), .Z(n19367) );
  NAND U22119 ( .A(n12794), .B(n12793), .Z(n19332) );
  AND U22120 ( .A(n12795), .B(n24262), .Z(n19330) );
  IV U22121 ( .A(n12796), .Z(n27650) );
  NAND U22122 ( .A(n27650), .B(n12797), .Z(n19328) );
  AND U22123 ( .A(n12799), .B(n12798), .Z(n27647) );
  NAND U22124 ( .A(n12803), .B(n12802), .Z(n27645) );
  AND U22125 ( .A(n12805), .B(n12804), .Z(n27644) );
  IV U22126 ( .A(n12806), .Z(n19317) );
  NAND U22127 ( .A(n19317), .B(n12807), .Z(n12808) );
  NAND U22128 ( .A(n12809), .B(n12808), .Z(n27643) );
  AND U22129 ( .A(n12810), .B(n27640), .Z(n19313) );
  AND U22130 ( .A(n27636), .B(n12811), .Z(n19307) );
  NAND U22131 ( .A(n27626), .B(n12814), .Z(n19293) );
  AND U22132 ( .A(n12818), .B(n12817), .Z(n19280) );
  IV U22133 ( .A(n12819), .Z(n27620) );
  OR U22134 ( .A(n12821), .B(n12820), .Z(n12822) );
  AND U22135 ( .A(n12823), .B(n12822), .Z(n19263) );
  AND U22136 ( .A(n27611), .B(n12824), .Z(n19260) );
  NANDN U22137 ( .A(y[2268]), .B(x[2268]), .Z(n12825) );
  NAND U22138 ( .A(n12826), .B(n12825), .Z(n19257) );
  NAND U22139 ( .A(n27607), .B(n12827), .Z(n19254) );
  IV U22140 ( .A(n12828), .Z(n27605) );
  IV U22141 ( .A(n12829), .Z(n27603) );
  NAND U22142 ( .A(n27603), .B(n12830), .Z(n19247) );
  AND U22143 ( .A(n12832), .B(n12831), .Z(n27602) );
  AND U22144 ( .A(n12836), .B(n12835), .Z(n27600) );
  NANDN U22145 ( .A(n27595), .B(n12841), .Z(n12843) );
  ANDN U22146 ( .B(n12843), .A(n12842), .Z(n19234) );
  IV U22147 ( .A(n12844), .Z(n27592) );
  AND U22148 ( .A(n27583), .B(n12850), .Z(n19210) );
  NANDN U22149 ( .A(n12858), .B(n12855), .Z(n12856) );
  AND U22150 ( .A(n12857), .B(n12856), .Z(n27578) );
  AND U22151 ( .A(n12862), .B(n24271), .Z(n12866) );
  OR U22152 ( .A(n12864), .B(n12863), .Z(n12865) );
  AND U22153 ( .A(n12866), .B(n12865), .Z(n19198) );
  AND U22154 ( .A(n12867), .B(n27576), .Z(n19196) );
  AND U22155 ( .A(n27575), .B(n24271), .Z(n12868) );
  NAND U22156 ( .A(n24273), .B(n12868), .Z(n19194) );
  IV U22157 ( .A(n12869), .Z(n27573) );
  AND U22158 ( .A(n12871), .B(n12870), .Z(n27570) );
  AND U22159 ( .A(n12872), .B(n27566), .Z(n19184) );
  NAND U22160 ( .A(n27554), .B(n12884), .Z(n19166) );
  AND U22161 ( .A(n12885), .B(n27555), .Z(n27552) );
  NAND U22162 ( .A(n12889), .B(n12888), .Z(n24276) );
  IV U22163 ( .A(n12890), .Z(n19152) );
  NANDN U22164 ( .A(n19152), .B(n12891), .Z(n12892) );
  AND U22165 ( .A(n12893), .B(n12892), .Z(n27548) );
  AND U22166 ( .A(n12895), .B(n12894), .Z(n19143) );
  AND U22167 ( .A(n12897), .B(n12896), .Z(n19137) );
  AND U22168 ( .A(n12899), .B(n12898), .Z(n19131) );
  AND U22169 ( .A(n12900), .B(n24278), .Z(n19122) );
  AND U22170 ( .A(n12902), .B(n12901), .Z(n19117) );
  IV U22171 ( .A(n12903), .Z(n27535) );
  NAND U22172 ( .A(n27534), .B(n27535), .Z(n19115) );
  ANDN U22173 ( .B(y[2180]), .A(x[2180]), .Z(n12904) );
  NAND U22174 ( .A(n12904), .B(n19106), .Z(n12905) );
  AND U22175 ( .A(n12905), .B(n19112), .Z(n12907) );
  ANDN U22176 ( .B(n12907), .A(n12906), .Z(n27532) );
  AND U22177 ( .A(n12909), .B(n12908), .Z(n19105) );
  IV U22178 ( .A(n12910), .Z(n27528) );
  NAND U22179 ( .A(n27528), .B(n12911), .Z(n19103) );
  IV U22180 ( .A(n12912), .Z(n27526) );
  AND U22181 ( .A(n12916), .B(n12915), .Z(n19083) );
  AND U22182 ( .A(n12918), .B(n12917), .Z(n19077) );
  AND U22183 ( .A(n12920), .B(n12919), .Z(n19071) );
  NAND U22184 ( .A(n27516), .B(n12921), .Z(n19069) );
  NAND U22185 ( .A(n12925), .B(n12924), .Z(n19059) );
  NAND U22186 ( .A(n27507), .B(n12926), .Z(n19052) );
  AND U22187 ( .A(n12927), .B(n27506), .Z(n19050) );
  IV U22188 ( .A(n12930), .Z(n27498) );
  IV U22189 ( .A(n12931), .Z(n27500) );
  AND U22190 ( .A(n27498), .B(n27500), .Z(n19037) );
  AND U22191 ( .A(n12933), .B(n12932), .Z(n24289) );
  NAND U22192 ( .A(n12939), .B(n12936), .Z(n12937) );
  AND U22193 ( .A(n12938), .B(n12937), .Z(n27493) );
  AND U22194 ( .A(n12944), .B(n12943), .Z(n27491) );
  AND U22195 ( .A(n12945), .B(n27489), .Z(n19021) );
  AND U22196 ( .A(n27486), .B(n12946), .Z(n19019) );
  IV U22197 ( .A(n12947), .Z(n27487) );
  AND U22198 ( .A(n12949), .B(n12948), .Z(n27483) );
  AND U22199 ( .A(n12950), .B(n27479), .Z(n19004) );
  NAND U22200 ( .A(n12956), .B(n12955), .Z(n27471) );
  AND U22201 ( .A(n12959), .B(n27468), .Z(n18986) );
  AND U22202 ( .A(n12961), .B(n12960), .Z(n27463) );
  AND U22203 ( .A(n27462), .B(n12962), .Z(n18978) );
  AND U22204 ( .A(n27457), .B(n12963), .Z(n18969) );
  NAND U22205 ( .A(n12965), .B(n12964), .Z(n27456) );
  AND U22206 ( .A(n12966), .B(n27454), .Z(n18966) );
  IV U22207 ( .A(n12967), .Z(n27449) );
  AND U22208 ( .A(n12968), .B(n27449), .Z(n18961) );
  NAND U22209 ( .A(n12972), .B(n12971), .Z(n18954) );
  AND U22210 ( .A(n27445), .B(n27447), .Z(n18952) );
  AND U22211 ( .A(n12974), .B(n12973), .Z(n24294) );
  OR U22212 ( .A(n12978), .B(n12977), .Z(n12979) );
  AND U22213 ( .A(n12980), .B(n12979), .Z(n27439) );
  AND U22214 ( .A(n12983), .B(n24296), .Z(n18933) );
  NAND U22215 ( .A(n27430), .B(n12988), .Z(n18916) );
  IV U22216 ( .A(n12989), .Z(n27429) );
  IV U22217 ( .A(n12990), .Z(n27426) );
  AND U22218 ( .A(n27429), .B(n27426), .Z(n18914) );
  NAND U22219 ( .A(n27424), .B(n12994), .Z(n18909) );
  AND U22220 ( .A(n12995), .B(n24300), .Z(n18907) );
  IV U22221 ( .A(n12996), .Z(n27420) );
  IV U22222 ( .A(n12997), .Z(n27419) );
  NOR U22223 ( .A(n13002), .B(n13001), .Z(n18887) );
  AND U22224 ( .A(n13003), .B(n24304), .Z(n18882) );
  AND U22225 ( .A(n24306), .B(n13006), .Z(n27407) );
  NAND U22226 ( .A(n13009), .B(n27401), .Z(n18868) );
  NAND U22227 ( .A(n27398), .B(n13011), .Z(n18865) );
  NAND U22228 ( .A(n13017), .B(n13016), .Z(n27395) );
  AND U22229 ( .A(n13018), .B(n27394), .Z(n18857) );
  NAND U22230 ( .A(n24309), .B(n13019), .Z(n24310) );
  AND U22231 ( .A(n27393), .B(n13020), .Z(n18854) );
  AND U22232 ( .A(n13021), .B(n27391), .Z(n18849) );
  AND U22233 ( .A(n13022), .B(n27384), .Z(n18837) );
  AND U22234 ( .A(n13025), .B(n27378), .Z(n18828) );
  IV U22235 ( .A(n13028), .Z(n27375) );
  NAND U22236 ( .A(n27375), .B(n13029), .Z(n18822) );
  AND U22237 ( .A(n27372), .B(n24311), .Z(n18820) );
  NAND U22238 ( .A(n27369), .B(n13032), .Z(n18814) );
  AND U22239 ( .A(n27368), .B(n13033), .Z(n18812) );
  IV U22240 ( .A(n13034), .Z(n27364) );
  IV U22241 ( .A(n13035), .Z(n27363) );
  OR U22242 ( .A(n13037), .B(n13036), .Z(n13039) );
  IV U22243 ( .A(n13038), .Z(n27361) );
  AND U22244 ( .A(n13039), .B(n27361), .Z(n18794) );
  AND U22245 ( .A(n13040), .B(n27359), .Z(n18792) );
  NAND U22246 ( .A(n13042), .B(n13041), .Z(n18790) );
  AND U22247 ( .A(n13044), .B(n13043), .Z(n18788) );
  AND U22248 ( .A(n13046), .B(n13045), .Z(n18782) );
  NANDN U22249 ( .A(x[2022]), .B(y[2022]), .Z(n27352) );
  IV U22250 ( .A(n13049), .Z(n27348) );
  AND U22251 ( .A(n13050), .B(n27348), .Z(n18772) );
  NAND U22252 ( .A(n27349), .B(n13051), .Z(n27347) );
  IV U22253 ( .A(n13052), .Z(n27346) );
  AND U22254 ( .A(n13053), .B(n27346), .Z(n18769) );
  NAND U22255 ( .A(n13055), .B(n13054), .Z(n27345) );
  NAND U22256 ( .A(n13059), .B(n13058), .Z(n27342) );
  IV U22257 ( .A(n13062), .Z(n27338) );
  AND U22258 ( .A(n13067), .B(n13066), .Z(n18743) );
  AND U22259 ( .A(n13069), .B(n13068), .Z(n18735) );
  AND U22260 ( .A(n27322), .B(n13071), .Z(n18732) );
  NAND U22261 ( .A(n13077), .B(n13076), .Z(n27319) );
  IV U22262 ( .A(n13078), .Z(n27318) );
  AND U22263 ( .A(n13079), .B(n27318), .Z(n18727) );
  IV U22264 ( .A(n13080), .Z(n27317) );
  NAND U22265 ( .A(n27313), .B(n13081), .Z(n18718) );
  AND U22266 ( .A(n13083), .B(n13082), .Z(n27312) );
  AND U22267 ( .A(n13087), .B(n13086), .Z(n27310) );
  NAND U22268 ( .A(n13091), .B(n13090), .Z(n27301) );
  NAND U22269 ( .A(n13095), .B(n13094), .Z(n27299) );
  IV U22270 ( .A(n13096), .Z(n27297) );
  AND U22271 ( .A(n13100), .B(n27287), .Z(n18674) );
  OR U22272 ( .A(n13102), .B(n13101), .Z(n13103) );
  NAND U22273 ( .A(n13104), .B(n13103), .Z(n13105) );
  NANDN U22274 ( .A(n13106), .B(n13105), .Z(n18658) );
  AND U22275 ( .A(n27277), .B(n27275), .Z(n18656) );
  NAND U22276 ( .A(n13114), .B(n13113), .Z(n27260) );
  NAND U22277 ( .A(n13122), .B(n13121), .Z(n27256) );
  NAND U22278 ( .A(n13126), .B(n13125), .Z(n18617) );
  AND U22279 ( .A(n13128), .B(n13127), .Z(n18615) );
  NAND U22280 ( .A(n24329), .B(n13129), .Z(n18613) );
  AND U22281 ( .A(n27248), .B(n13130), .Z(n18611) );
  AND U22282 ( .A(n13138), .B(n13137), .Z(n27243) );
  IV U22283 ( .A(n13139), .Z(n27239) );
  NOR U22284 ( .A(n27239), .B(n13140), .Z(n18594) );
  AND U22285 ( .A(n13142), .B(n13141), .Z(n24331) );
  IV U22286 ( .A(n13147), .Z(n27228) );
  NOR U22287 ( .A(n13149), .B(n13148), .Z(n18566) );
  IV U22288 ( .A(n13150), .Z(n27223) );
  AND U22289 ( .A(n13151), .B(n27223), .Z(n18560) );
  NAND U22290 ( .A(n13153), .B(n13152), .Z(n27222) );
  NANDN U22291 ( .A(n18549), .B(n13154), .Z(n13156) );
  IV U22292 ( .A(n13155), .Z(n24333) );
  AND U22293 ( .A(n13156), .B(n24333), .Z(n18557) );
  AND U22294 ( .A(n13158), .B(n13157), .Z(n18548) );
  NAND U22295 ( .A(n13166), .B(n13165), .Z(n27210) );
  AND U22296 ( .A(n13168), .B(n13167), .Z(n24337) );
  NAND U22297 ( .A(n13172), .B(n13171), .Z(n27207) );
  NAND U22298 ( .A(n27204), .B(n13173), .Z(n18528) );
  AND U22299 ( .A(n13175), .B(n13174), .Z(n18523) );
  AND U22300 ( .A(n13177), .B(n13176), .Z(n27197) );
  AND U22301 ( .A(n13183), .B(n13182), .Z(n27194) );
  AND U22302 ( .A(n13184), .B(n27192), .Z(n18510) );
  IV U22303 ( .A(n13185), .Z(n27191) );
  NAND U22304 ( .A(n27191), .B(n13186), .Z(n18508) );
  AND U22305 ( .A(n13190), .B(n13189), .Z(n27184) );
  AND U22306 ( .A(n13196), .B(n13195), .Z(n27181) );
  NAND U22307 ( .A(n13204), .B(n13203), .Z(n24339) );
  AND U22308 ( .A(n13208), .B(n13207), .Z(n27167) );
  AND U22309 ( .A(n27163), .B(n13211), .Z(n18466) );
  NAND U22310 ( .A(n27160), .B(n13212), .Z(n18464) );
  NAND U22311 ( .A(n13224), .B(n13223), .Z(n27139) );
  AND U22312 ( .A(n13225), .B(n27129), .Z(n18441) );
  NAND U22313 ( .A(n27125), .B(n13226), .Z(n18433) );
  AND U22314 ( .A(n13230), .B(n13229), .Z(n24340) );
  NAND U22315 ( .A(n13236), .B(n13235), .Z(n27121) );
  IV U22316 ( .A(n13237), .Z(n27120) );
  AND U22317 ( .A(n13238), .B(n27120), .Z(n18426) );
  IV U22318 ( .A(n13239), .Z(n27119) );
  IV U22319 ( .A(n13240), .Z(n27116) );
  IV U22320 ( .A(n13241), .Z(n27115) );
  NAND U22321 ( .A(n13247), .B(n13246), .Z(n24341) );
  IV U22322 ( .A(n13254), .Z(n27101) );
  AND U22323 ( .A(n13256), .B(n13255), .Z(n24344) );
  AND U22324 ( .A(n13266), .B(n13265), .Z(n24345) );
  NAND U22325 ( .A(n13270), .B(n13269), .Z(n27084) );
  AND U22326 ( .A(n13272), .B(n13271), .Z(n24347) );
  AND U22327 ( .A(n13276), .B(n13275), .Z(n27074) );
  AND U22328 ( .A(n13280), .B(n13279), .Z(n27072) );
  AND U22329 ( .A(n13284), .B(n13283), .Z(n27070) );
  AND U22330 ( .A(n27064), .B(n13285), .Z(n18343) );
  AND U22331 ( .A(n13287), .B(n13286), .Z(n27063) );
  NAND U22332 ( .A(n13293), .B(n13292), .Z(n27060) );
  IV U22333 ( .A(n13296), .Z(n27057) );
  NAND U22334 ( .A(n27057), .B(n13297), .Z(n18324) );
  AND U22335 ( .A(n13299), .B(n13298), .Z(n18322) );
  XNOR U22336 ( .A(y[1775]), .B(x[1775]), .Z(n18316) );
  IV U22337 ( .A(n13300), .Z(n27052) );
  XNOR U22338 ( .A(y[1772]), .B(x[1772]), .Z(n13303) );
  AND U22339 ( .A(n13304), .B(n13303), .Z(n27049) );
  AND U22340 ( .A(n13308), .B(n13307), .Z(n27047) );
  AND U22341 ( .A(n27045), .B(n13311), .Z(n18304) );
  AND U22342 ( .A(n13313), .B(n13312), .Z(n24353) );
  AND U22343 ( .A(n13317), .B(n13316), .Z(n24354) );
  NAND U22344 ( .A(n27026), .B(n13320), .Z(n18271) );
  NAND U22345 ( .A(n27017), .B(n13323), .Z(n18261) );
  AND U22346 ( .A(n13324), .B(n27016), .Z(n18259) );
  AND U22347 ( .A(n13328), .B(n13327), .Z(n27012) );
  NAND U22348 ( .A(n13332), .B(n13331), .Z(n18229) );
  AND U22349 ( .A(n13334), .B(n13333), .Z(n18227) );
  NAND U22350 ( .A(n26999), .B(n13335), .Z(n18225) );
  IV U22351 ( .A(n13336), .Z(n26998) );
  AND U22352 ( .A(n13337), .B(n26998), .Z(n18223) );
  AND U22353 ( .A(n13344), .B(n26994), .Z(n18215) );
  AND U22354 ( .A(n26988), .B(n13345), .Z(n18206) );
  NAND U22355 ( .A(n13349), .B(n13348), .Z(n26985) );
  IV U22356 ( .A(n13352), .Z(n26979) );
  NAND U22357 ( .A(n13354), .B(n13353), .Z(n13356) );
  NAND U22358 ( .A(n13356), .B(n13355), .Z(n18181) );
  AND U22359 ( .A(n13358), .B(n13357), .Z(n26977) );
  AND U22360 ( .A(n13362), .B(n13361), .Z(n26974) );
  NAND U22361 ( .A(n13368), .B(n13367), .Z(n26971) );
  AND U22362 ( .A(n13370), .B(n13369), .Z(n26967) );
  IV U22363 ( .A(n13371), .Z(n26962) );
  IV U22364 ( .A(n13372), .Z(n26961) );
  NAND U22365 ( .A(n13374), .B(n13373), .Z(n26958) );
  NAND U22366 ( .A(n13378), .B(n13377), .Z(n26956) );
  IV U22367 ( .A(n13379), .Z(n26954) );
  NAND U22368 ( .A(n13381), .B(n13380), .Z(n26951) );
  NAND U22369 ( .A(n13385), .B(n13384), .Z(n26949) );
  AND U22370 ( .A(n13387), .B(n13386), .Z(n26948) );
  NANDN U22371 ( .A(x[1680]), .B(y[1680]), .Z(n13389) );
  NAND U22372 ( .A(n13389), .B(n13388), .Z(n26947) );
  AND U22373 ( .A(n13391), .B(n13390), .Z(n18131) );
  IV U22374 ( .A(n13392), .Z(n26945) );
  IV U22375 ( .A(n13393), .Z(n26943) );
  NAND U22376 ( .A(n26945), .B(n26943), .Z(n18129) );
  AND U22377 ( .A(n26942), .B(n13394), .Z(n18127) );
  NANDN U22378 ( .A(y[1672]), .B(x[1672]), .Z(n13396) );
  NAND U22379 ( .A(n13397), .B(n13396), .Z(n26937) );
  IV U22380 ( .A(n13402), .Z(n26934) );
  AND U22381 ( .A(n13403), .B(n26934), .Z(n18117) );
  NAND U22382 ( .A(n13407), .B(n13406), .Z(n26924) );
  NAND U22383 ( .A(n13411), .B(n13410), .Z(n26922) );
  AND U22384 ( .A(n13415), .B(n13414), .Z(n26916) );
  NAND U22385 ( .A(n13425), .B(n13424), .Z(n26910) );
  AND U22386 ( .A(n13426), .B(n26905), .Z(n18073) );
  AND U22387 ( .A(n13429), .B(n26896), .Z(n18044) );
  NAND U22388 ( .A(n26887), .B(n13430), .Z(n18017) );
  IV U22389 ( .A(n13431), .Z(n26886) );
  NAND U22390 ( .A(n26886), .B(n13432), .Z(n18015) );
  AND U22391 ( .A(n13434), .B(n13433), .Z(n18013) );
  NOR U22392 ( .A(n13443), .B(n26866), .Z(n17977) );
  AND U22393 ( .A(n13447), .B(n13446), .Z(n26861) );
  IV U22394 ( .A(n13448), .Z(n26855) );
  IV U22395 ( .A(n13449), .Z(n26848) );
  NAND U22396 ( .A(n13455), .B(n13454), .Z(n24383) );
  OR U22397 ( .A(n13460), .B(n13459), .Z(n13461) );
  AND U22398 ( .A(n13462), .B(n13461), .Z(n26833) );
  AND U22399 ( .A(n13467), .B(n13466), .Z(n26825) );
  IV U22400 ( .A(n13468), .Z(n26823) );
  IV U22401 ( .A(n13469), .Z(n26824) );
  NAND U22402 ( .A(n26823), .B(n26824), .Z(n17906) );
  NAND U22403 ( .A(n26819), .B(n26817), .Z(n17898) );
  AND U22404 ( .A(n13472), .B(n24387), .Z(n17896) );
  NANDN U22405 ( .A(x[1556]), .B(y[1556]), .Z(n13476) );
  NAND U22406 ( .A(n13476), .B(n13475), .Z(n26814) );
  IV U22407 ( .A(n13481), .Z(n26801) );
  AND U22408 ( .A(n13482), .B(n26801), .Z(n17857) );
  AND U22409 ( .A(n13484), .B(n13483), .Z(n26800) );
  AND U22410 ( .A(n13488), .B(n13487), .Z(n24393) );
  IV U22411 ( .A(n13489), .Z(n26785) );
  AND U22412 ( .A(n26777), .B(n13500), .Z(n17817) );
  IV U22413 ( .A(n13503), .Z(n26767) );
  IV U22414 ( .A(n13504), .Z(n26764) );
  IV U22415 ( .A(n13505), .Z(n26763) );
  NANDN U22416 ( .A(n26761), .B(n13506), .Z(n17785) );
  NAND U22417 ( .A(n13508), .B(n13507), .Z(n17777) );
  OR U22418 ( .A(n13516), .B(n13515), .Z(n13517) );
  AND U22419 ( .A(n26745), .B(n13517), .Z(n17761) );
  ANDN U22420 ( .B(n26738), .A(n26736), .Z(n17746) );
  NAND U22421 ( .A(n13524), .B(n13523), .Z(n26724) );
  IV U22422 ( .A(n13525), .Z(n26720) );
  AND U22423 ( .A(n13526), .B(n26720), .Z(n17712) );
  AND U22424 ( .A(n13528), .B(n13527), .Z(n24403) );
  AND U22425 ( .A(n13535), .B(n26716), .Z(n17706) );
  NAND U22426 ( .A(n26668), .B(n24405), .Z(n17622) );
  NAND U22427 ( .A(n13550), .B(n13549), .Z(n26666) );
  AND U22428 ( .A(n13551), .B(n26665), .Z(n17616) );
  IV U22429 ( .A(n13552), .Z(n26662) );
  NAND U22430 ( .A(n13554), .B(n13553), .Z(n26660) );
  OR U22431 ( .A(n13556), .B(n13555), .Z(n13557) );
  AND U22432 ( .A(n26656), .B(n13557), .Z(n17601) );
  NANDN U22433 ( .A(x[1398]), .B(y[1398]), .Z(n13559) );
  AND U22434 ( .A(n13559), .B(n13558), .Z(n26650) );
  AND U22435 ( .A(n13563), .B(n13562), .Z(n26648) );
  IV U22436 ( .A(n13568), .Z(n26633) );
  NAND U22437 ( .A(n26633), .B(n13569), .Z(n17573) );
  AND U22438 ( .A(n26630), .B(n13570), .Z(n17571) );
  NAND U22439 ( .A(n13572), .B(n13571), .Z(n17569) );
  IV U22440 ( .A(n13573), .Z(n26606) );
  NAND U22441 ( .A(n13578), .B(n13577), .Z(n26602) );
  NANDN U22442 ( .A(x[1374]), .B(y[1374]), .Z(n13579) );
  AND U22443 ( .A(n13579), .B(n26600), .Z(n26599) );
  NOR U22444 ( .A(n13583), .B(n13582), .Z(n17533) );
  AND U22445 ( .A(n13588), .B(n24409), .Z(n17514) );
  NAND U22446 ( .A(n13590), .B(n13589), .Z(n26580) );
  NAND U22447 ( .A(n26577), .B(n13591), .Z(n26576) );
  AND U22448 ( .A(n24411), .B(n13592), .Z(n17500) );
  NAND U22449 ( .A(n13594), .B(n13593), .Z(n24410) );
  AND U22450 ( .A(n13596), .B(n13595), .Z(n17497) );
  IV U22451 ( .A(n13597), .Z(n26572) );
  NOR U22452 ( .A(n26572), .B(n13598), .Z(n17495) );
  NAND U22453 ( .A(n13600), .B(n13599), .Z(n17470) );
  AND U22454 ( .A(n13602), .B(n13601), .Z(n17454) );
  IV U22455 ( .A(n13603), .Z(n26557) );
  NANDN U22456 ( .A(y[1331]), .B(x[1331]), .Z(n13604) );
  AND U22457 ( .A(n13605), .B(n13604), .Z(n26552) );
  NAND U22458 ( .A(n13608), .B(n13607), .Z(n24416) );
  NOR U22459 ( .A(n13609), .B(n26545), .Z(n17423) );
  AND U22460 ( .A(n13615), .B(n13614), .Z(n17401) );
  AND U22461 ( .A(n26533), .B(n13618), .Z(n17392) );
  IV U22462 ( .A(n13619), .Z(n26529) );
  IV U22463 ( .A(n13620), .Z(n26528) );
  NAND U22464 ( .A(n13622), .B(n13621), .Z(n26525) );
  AND U22465 ( .A(n13628), .B(n13627), .Z(n26522) );
  IV U22466 ( .A(n13629), .Z(n26521) );
  NAND U22467 ( .A(n26521), .B(n26520), .Z(n17372) );
  AND U22468 ( .A(n13631), .B(n13630), .Z(n17370) );
  NANDN U22469 ( .A(x[1296]), .B(y[1296]), .Z(n13632) );
  NAND U22470 ( .A(n13633), .B(n13632), .Z(n26517) );
  AND U22471 ( .A(n13634), .B(n26516), .Z(n17367) );
  AND U22472 ( .A(n13636), .B(n13635), .Z(n26514) );
  NAND U22473 ( .A(n13640), .B(n13639), .Z(n26512) );
  IV U22474 ( .A(n13641), .Z(n13645) );
  AND U22475 ( .A(n13647), .B(n13646), .Z(n17356) );
  IV U22476 ( .A(n13648), .Z(n26508) );
  NOR U22477 ( .A(n26508), .B(n13649), .Z(n17352) );
  NAND U22478 ( .A(n13653), .B(n13652), .Z(n26498) );
  IV U22479 ( .A(n13654), .Z(n26497) );
  NAND U22480 ( .A(n13658), .B(n13657), .Z(n26491) );
  IV U22481 ( .A(n13659), .Z(n26490) );
  AND U22482 ( .A(n13661), .B(n13660), .Z(n17293) );
  NAND U22483 ( .A(n13663), .B(n13662), .Z(n24429) );
  ANDN U22484 ( .B(n26484), .A(n26482), .Z(n17280) );
  IV U22485 ( .A(n13664), .Z(n26481) );
  AND U22486 ( .A(n13666), .B(n13665), .Z(n26480) );
  AND U22487 ( .A(n13668), .B(n13667), .Z(n24432) );
  AND U22488 ( .A(n26473), .B(n13669), .Z(n17261) );
  NAND U22489 ( .A(n13671), .B(n13670), .Z(n26468) );
  IV U22490 ( .A(n13672), .Z(n26464) );
  ANDN U22491 ( .B(n26466), .A(n26464), .Z(n17248) );
  NAND U22492 ( .A(n13674), .B(n13673), .Z(n26463) );
  AND U22493 ( .A(n13678), .B(n13677), .Z(n26460) );
  AND U22494 ( .A(n13681), .B(n26458), .Z(n17239) );
  NANDN U22495 ( .A(x[1232]), .B(y[1232]), .Z(n26453) );
  NOR U22496 ( .A(n13683), .B(n13682), .Z(n17231) );
  AND U22497 ( .A(n26447), .B(n13684), .Z(n17209) );
  AND U22498 ( .A(n26443), .B(n13687), .Z(n17206) );
  NAND U22499 ( .A(n26437), .B(n26442), .Z(n17204) );
  AND U22500 ( .A(n26436), .B(n13688), .Z(n17202) );
  XNOR U22501 ( .A(x[1213]), .B(y[1213]), .Z(n17187) );
  NOR U22502 ( .A(n26408), .B(n13691), .Z(n17168) );
  AND U22503 ( .A(n13693), .B(n13692), .Z(n26404) );
  IV U22504 ( .A(n13698), .Z(n26400) );
  IV U22505 ( .A(n13699), .Z(n24441) );
  IV U22506 ( .A(n13702), .Z(n26397) );
  ANDN U22507 ( .B(n26397), .A(n24443), .Z(n17142) );
  IV U22508 ( .A(n13703), .Z(n26396) );
  IV U22509 ( .A(n13707), .Z(n26389) );
  IV U22510 ( .A(n13708), .Z(n26386) );
  NANDN U22511 ( .A(n26378), .B(n13712), .Z(n17100) );
  AND U22512 ( .A(n13713), .B(n26377), .Z(n17098) );
  AND U22513 ( .A(n13717), .B(n13716), .Z(n24446) );
  NAND U22514 ( .A(n13719), .B(n13718), .Z(n26374) );
  NAND U22515 ( .A(n13727), .B(n13726), .Z(n26370) );
  IV U22516 ( .A(n13728), .Z(n26369) );
  NAND U22517 ( .A(n13730), .B(n13729), .Z(n13731) );
  NAND U22518 ( .A(n13732), .B(n13731), .Z(n26366) );
  IV U22519 ( .A(n13733), .Z(n26360) );
  AND U22520 ( .A(n13737), .B(n13736), .Z(n17060) );
  NAND U22521 ( .A(n13739), .B(n13738), .Z(n24447) );
  NANDN U22522 ( .A(n13743), .B(n13742), .Z(n26344) );
  AND U22523 ( .A(n13752), .B(n13751), .Z(n26338) );
  AND U22524 ( .A(n13757), .B(n24453), .Z(n17019) );
  AND U22525 ( .A(n13758), .B(n26334), .Z(n17013) );
  AND U22526 ( .A(n13759), .B(n26327), .Z(n16989) );
  NAND U22527 ( .A(n13761), .B(n13760), .Z(n26322) );
  IV U22528 ( .A(n13762), .Z(n13768) );
  IV U22529 ( .A(n13769), .Z(n26318) );
  AND U22530 ( .A(n13770), .B(n26318), .Z(n16976) );
  AND U22531 ( .A(n13771), .B(n26316), .Z(n26315) );
  AND U22532 ( .A(n26314), .B(n13772), .Z(n16973) );
  AND U22533 ( .A(n13773), .B(n26312), .Z(n16968) );
  NAND U22534 ( .A(n26311), .B(n26309), .Z(n16966) );
  IV U22535 ( .A(n13774), .Z(n26308) );
  AND U22536 ( .A(n13775), .B(n26308), .Z(n16964) );
  AND U22537 ( .A(n13777), .B(n13776), .Z(n24459) );
  ANDN U22538 ( .B(n13779), .A(n13778), .Z(n26307) );
  OR U22539 ( .A(n13781), .B(n13780), .Z(n13782) );
  NAND U22540 ( .A(n13783), .B(n13782), .Z(n13784) );
  NANDN U22541 ( .A(n13785), .B(n13784), .Z(n16952) );
  NAND U22542 ( .A(n13792), .B(n13788), .Z(n13789) );
  AND U22543 ( .A(n13790), .B(n13789), .Z(n26294) );
  IV U22544 ( .A(n13795), .Z(n26291) );
  NAND U22545 ( .A(n26291), .B(n13796), .Z(n16935) );
  AND U22546 ( .A(n13797), .B(n26289), .Z(n16933) );
  IV U22547 ( .A(n13800), .Z(n26285) );
  AND U22548 ( .A(n13805), .B(n13804), .Z(n26283) );
  NAND U22549 ( .A(n13807), .B(n13806), .Z(n26282) );
  IV U22550 ( .A(n13812), .Z(n26279) );
  IV U22551 ( .A(n13819), .Z(n26269) );
  IV U22552 ( .A(n13822), .Z(n26261) );
  NAND U22553 ( .A(n13824), .B(n13823), .Z(n16860) );
  AND U22554 ( .A(n13826), .B(n13825), .Z(n16858) );
  ANDN U22555 ( .B(n26252), .A(n26250), .Z(n16846) );
  IV U22556 ( .A(n13829), .Z(n26249) );
  AND U22557 ( .A(n13833), .B(n13832), .Z(n24472) );
  AND U22558 ( .A(n13837), .B(n13836), .Z(n26244) );
  IV U22559 ( .A(n13840), .Z(n26242) );
  IV U22560 ( .A(n13841), .Z(n26241) );
  NAND U22561 ( .A(n13856), .B(n13855), .Z(n24476) );
  AND U22562 ( .A(n13858), .B(n13857), .Z(n16785) );
  NAND U22563 ( .A(n13864), .B(n13863), .Z(n26211) );
  XNOR U22564 ( .A(y[982]), .B(x[982]), .Z(n13874) );
  AND U22565 ( .A(n13875), .B(n13874), .Z(n26192) );
  AND U22566 ( .A(n13879), .B(n13878), .Z(n26190) );
  ANDN U22567 ( .B(n13880), .A(n26184), .Z(n16701) );
  AND U22568 ( .A(n26183), .B(n13881), .Z(n16699) );
  AND U22569 ( .A(n13887), .B(n13886), .Z(n26179) );
  AND U22570 ( .A(n13891), .B(n13890), .Z(n26177) );
  NAND U22571 ( .A(n13897), .B(n13896), .Z(n26164) );
  AND U22572 ( .A(n13903), .B(n13902), .Z(n26161) );
  NAND U22573 ( .A(n13905), .B(n13904), .Z(n26160) );
  NAND U22574 ( .A(n13913), .B(n13912), .Z(n26156) );
  NAND U22575 ( .A(n13917), .B(n13916), .Z(n26154) );
  IV U22576 ( .A(n13918), .Z(n26153) );
  AND U22577 ( .A(n13919), .B(n26153), .Z(n16650) );
  IV U22578 ( .A(n13920), .Z(n26149) );
  IV U22579 ( .A(n13921), .Z(n26147) );
  AND U22580 ( .A(n13923), .B(n13922), .Z(n16636) );
  NAND U22581 ( .A(n13927), .B(n13926), .Z(n24487) );
  XNOR U22582 ( .A(y[930]), .B(x[930]), .Z(n16619) );
  NAND U22583 ( .A(n26129), .B(n26131), .Z(n16605) );
  NAND U22584 ( .A(n13935), .B(n13934), .Z(n26125) );
  NAND U22585 ( .A(n13939), .B(n13938), .Z(n26123) );
  IV U22586 ( .A(n13942), .Z(n26120) );
  NAND U22587 ( .A(n13944), .B(n13943), .Z(n16582) );
  AND U22588 ( .A(n13946), .B(n13945), .Z(n16580) );
  NAND U22589 ( .A(n13948), .B(n13947), .Z(n16578) );
  AND U22590 ( .A(n13950), .B(n13949), .Z(n26114) );
  NAND U22591 ( .A(n13952), .B(n13951), .Z(n26113) );
  AND U22592 ( .A(n26104), .B(n13961), .Z(n13966) );
  NAND U22593 ( .A(n13962), .B(n26105), .Z(n13963) );
  NAND U22594 ( .A(n13966), .B(n13963), .Z(n13964) );
  AND U22595 ( .A(n26106), .B(n13964), .Z(n16559) );
  AND U22596 ( .A(n13966), .B(n13965), .Z(n26103) );
  NAND U22597 ( .A(n26103), .B(n26101), .Z(n16557) );
  NAND U22598 ( .A(n13968), .B(n13967), .Z(n24498) );
  NAND U22599 ( .A(n26097), .B(n26099), .Z(n16548) );
  AND U22600 ( .A(n13970), .B(n13969), .Z(n26096) );
  IV U22601 ( .A(n13971), .Z(n26092) );
  IV U22602 ( .A(n13972), .Z(n26091) );
  NAND U22603 ( .A(n26092), .B(n26091), .Z(n16539) );
  NAND U22604 ( .A(n13974), .B(n13973), .Z(n24501) );
  AND U22605 ( .A(n13979), .B(n26085), .Z(n16525) );
  AND U22606 ( .A(n13980), .B(n24504), .Z(n16503) );
  AND U22607 ( .A(n13981), .B(n26076), .Z(n16498) );
  IV U22608 ( .A(n13982), .Z(n26075) );
  IV U22609 ( .A(n13983), .Z(n26074) );
  NAND U22610 ( .A(n26075), .B(n26074), .Z(n16496) );
  AND U22611 ( .A(n26073), .B(n13984), .Z(n16494) );
  AND U22612 ( .A(n13991), .B(n13990), .Z(n26069) );
  AND U22613 ( .A(n13995), .B(n13994), .Z(n16473) );
  IV U22614 ( .A(n13996), .Z(n26057) );
  IV U22615 ( .A(n13997), .Z(n26055) );
  AND U22616 ( .A(n26056), .B(n26055), .Z(n16453) );
  NAND U22617 ( .A(n13999), .B(n13998), .Z(n26054) );
  AND U22618 ( .A(n14001), .B(n14000), .Z(n26053) );
  AND U22619 ( .A(n14005), .B(n14004), .Z(n26051) );
  NOR U22620 ( .A(n14006), .B(n26050), .Z(n16447) );
  AND U22621 ( .A(n26043), .B(n24508), .Z(n16437) );
  IV U22622 ( .A(n14012), .Z(n26036) );
  IV U22623 ( .A(n14013), .Z(n26034) );
  NANDN U22624 ( .A(x[834]), .B(y[834]), .Z(n14014) );
  AND U22625 ( .A(n14015), .B(n14014), .Z(n26029) );
  AND U22626 ( .A(n14019), .B(n14018), .Z(n26025) );
  AND U22627 ( .A(n26000), .B(n26005), .Z(n16393) );
  AND U22628 ( .A(n14021), .B(n14020), .Z(n25997) );
  AND U22629 ( .A(n14025), .B(n14024), .Z(n25993) );
  AND U22630 ( .A(n14033), .B(n14032), .Z(n25985) );
  NAND U22631 ( .A(n14035), .B(n14034), .Z(n25983) );
  XNOR U22632 ( .A(x[810]), .B(y[810]), .Z(n14045) );
  NANDN U22633 ( .A(n14046), .B(n14045), .Z(n25971) );
  AND U22634 ( .A(n14048), .B(n14047), .Z(n25969) );
  IV U22635 ( .A(n14049), .Z(n14051) );
  NAND U22636 ( .A(n14051), .B(n14050), .Z(n25967) );
  IV U22637 ( .A(n14052), .Z(n14053) );
  AND U22638 ( .A(n14054), .B(n14053), .Z(n25965) );
  IV U22639 ( .A(n14055), .Z(n14057) );
  NAND U22640 ( .A(n14057), .B(n14056), .Z(n25963) );
  IV U22641 ( .A(n14058), .Z(n14059) );
  AND U22642 ( .A(n14060), .B(n14059), .Z(n25961) );
  NAND U22643 ( .A(n14062), .B(n14061), .Z(n25959) );
  IV U22644 ( .A(n14063), .Z(n14064) );
  AND U22645 ( .A(n14065), .B(n14064), .Z(n25957) );
  NAND U22646 ( .A(n14067), .B(n14066), .Z(n25955) );
  XNOR U22647 ( .A(x[800]), .B(y[800]), .Z(n14070) );
  NANDN U22648 ( .A(n14071), .B(n14070), .Z(n25951) );
  AND U22649 ( .A(n14077), .B(n14076), .Z(n25948) );
  IV U22650 ( .A(n14080), .Z(n25945) );
  IV U22651 ( .A(n14081), .Z(n25944) );
  IV U22652 ( .A(n14082), .Z(n25943) );
  IV U22653 ( .A(n14083), .Z(n25942) );
  IV U22654 ( .A(n14084), .Z(n25939) );
  NANDN U22655 ( .A(y[786]), .B(x[786]), .Z(n14088) );
  NAND U22656 ( .A(n14088), .B(n14087), .Z(n25937) );
  IV U22657 ( .A(n14089), .Z(n25936) );
  NANDN U22658 ( .A(y[773]), .B(x[773]), .Z(n14091) );
  AND U22659 ( .A(n14092), .B(n14091), .Z(n25929) );
  AND U22660 ( .A(n14096), .B(n14095), .Z(n25927) );
  AND U22661 ( .A(n14100), .B(n14099), .Z(n24515) );
  NAND U22662 ( .A(n14104), .B(n14103), .Z(n24516) );
  IV U22663 ( .A(n14111), .Z(n14113) );
  ANDN U22664 ( .B(n14113), .A(n14112), .Z(n25917) );
  XNOR U22665 ( .A(x[760]), .B(y[760]), .Z(n14116) );
  IV U22666 ( .A(n14114), .Z(n14115) );
  AND U22667 ( .A(n14116), .B(n14115), .Z(n25916) );
  NAND U22668 ( .A(n14118), .B(n14117), .Z(n25915) );
  XNOR U22669 ( .A(x[756]), .B(y[756]), .Z(n14123) );
  IV U22670 ( .A(n14121), .Z(n14122) );
  AND U22671 ( .A(n14123), .B(n14122), .Z(n25913) );
  XNOR U22672 ( .A(x[754]), .B(y[754]), .Z(n14126) );
  AND U22673 ( .A(n14127), .B(n14126), .Z(n25909) );
  XNOR U22674 ( .A(x[752]), .B(y[752]), .Z(n14130) );
  AND U22675 ( .A(n14131), .B(n14130), .Z(n24519) );
  AND U22676 ( .A(n14138), .B(n14137), .Z(n24521) );
  IV U22677 ( .A(n14141), .Z(n14142) );
  AND U22678 ( .A(n14143), .B(n14142), .Z(n25901) );
  XNOR U22679 ( .A(y[742]), .B(x[742]), .Z(n14146) );
  IV U22680 ( .A(n14144), .Z(n14145) );
  AND U22681 ( .A(n14146), .B(n14145), .Z(n25900) );
  NAND U22682 ( .A(n14148), .B(n14147), .Z(n25899) );
  XNOR U22683 ( .A(x[740]), .B(y[740]), .Z(n14151) );
  IV U22684 ( .A(n14149), .Z(n14150) );
  AND U22685 ( .A(n14151), .B(n14150), .Z(n25898) );
  NANDN U22686 ( .A(x[736]), .B(y[736]), .Z(n14155) );
  NAND U22687 ( .A(n14155), .B(n14154), .Z(n24523) );
  AND U22688 ( .A(n14157), .B(n14156), .Z(n25895) );
  XNOR U22689 ( .A(y[734]), .B(x[734]), .Z(n14160) );
  AND U22690 ( .A(n14161), .B(n14160), .Z(n24524) );
  IV U22691 ( .A(n14166), .Z(n14167) );
  AND U22692 ( .A(n14168), .B(n14167), .Z(n25890) );
  AND U22693 ( .A(n14170), .B(n14169), .Z(n24526) );
  IV U22694 ( .A(n14171), .Z(n14172) );
  AND U22695 ( .A(n14173), .B(n14172), .Z(n25888) );
  NANDN U22696 ( .A(x[722]), .B(y[722]), .Z(n14179) );
  NAND U22697 ( .A(n14179), .B(n14178), .Z(n25884) );
  AND U22698 ( .A(n14181), .B(n14180), .Z(n24527) );
  IV U22699 ( .A(n14182), .Z(n14184) );
  ANDN U22700 ( .B(n14184), .A(n14183), .Z(n25882) );
  AND U22701 ( .A(n14186), .B(n14185), .Z(n25881) );
  AND U22702 ( .A(n14193), .B(n14192), .Z(n25876) );
  ANDN U22703 ( .B(n14195), .A(n14194), .Z(n25875) );
  NAND U22704 ( .A(n14201), .B(n14200), .Z(n24530) );
  IV U22705 ( .A(n14202), .Z(n14203) );
  AND U22706 ( .A(n14204), .B(n14203), .Z(n25870) );
  IV U22707 ( .A(n14205), .Z(n14206) );
  AND U22708 ( .A(n14207), .B(n14206), .Z(n25869) );
  XNOR U22709 ( .A(y[704]), .B(x[704]), .Z(n14208) );
  AND U22710 ( .A(n14209), .B(n14208), .Z(n24531) );
  IV U22711 ( .A(n14210), .Z(n14212) );
  ANDN U22712 ( .B(n14212), .A(n14211), .Z(n25867) );
  AND U22713 ( .A(n14214), .B(n14213), .Z(n25866) );
  IV U22714 ( .A(n14215), .Z(n14216) );
  AND U22715 ( .A(n14217), .B(n14216), .Z(n25865) );
  AND U22716 ( .A(n14219), .B(n14218), .Z(n24533) );
  AND U22717 ( .A(n14223), .B(n14222), .Z(n25861) );
  NAND U22718 ( .A(n14229), .B(n14228), .Z(n24537) );
  AND U22719 ( .A(n14231), .B(n14230), .Z(n25853) );
  XNOR U22720 ( .A(x[682]), .B(y[682]), .Z(n14235) );
  NANDN U22721 ( .A(n14236), .B(n14235), .Z(n25850) );
  AND U22722 ( .A(n14238), .B(n14237), .Z(n25848) );
  AND U22723 ( .A(n14242), .B(n14241), .Z(n25844) );
  XNOR U22724 ( .A(y[678]), .B(x[678]), .Z(n14243) );
  NANDN U22725 ( .A(n14244), .B(n14243), .Z(n25842) );
  AND U22726 ( .A(n14246), .B(n14245), .Z(n25840) );
  XNOR U22727 ( .A(x[676]), .B(y[676]), .Z(n14247) );
  NANDN U22728 ( .A(n14248), .B(n14247), .Z(n25838) );
  AND U22729 ( .A(n14250), .B(n14249), .Z(n25836) );
  AND U22730 ( .A(n14254), .B(n14253), .Z(n25832) );
  XNOR U22731 ( .A(x[672]), .B(y[672]), .Z(n14255) );
  NANDN U22732 ( .A(n14256), .B(n14255), .Z(n25830) );
  AND U22733 ( .A(n14258), .B(n14257), .Z(n25828) );
  AND U22734 ( .A(n14262), .B(n14261), .Z(n25824) );
  AND U22735 ( .A(n14266), .B(n14265), .Z(n25820) );
  NANDN U22736 ( .A(x[662]), .B(y[662]), .Z(n14269) );
  AND U22737 ( .A(n14270), .B(n14269), .Z(n25812) );
  AND U22738 ( .A(n14274), .B(n14273), .Z(n25808) );
  XNOR U22739 ( .A(x[660]), .B(y[660]), .Z(n14275) );
  NANDN U22740 ( .A(n14276), .B(n14275), .Z(n25806) );
  AND U22741 ( .A(n14278), .B(n14277), .Z(n25804) );
  AND U22742 ( .A(n14282), .B(n14281), .Z(n25800) );
  AND U22743 ( .A(n14286), .B(n14285), .Z(n25796) );
  NANDN U22744 ( .A(x[652]), .B(y[652]), .Z(n14290) );
  AND U22745 ( .A(n14290), .B(n14289), .Z(n25792) );
  NANDN U22746 ( .A(x[650]), .B(y[650]), .Z(n14294) );
  AND U22747 ( .A(n14294), .B(n14293), .Z(n25788) );
  NANDN U22748 ( .A(x[648]), .B(y[648]), .Z(n14298) );
  AND U22749 ( .A(n14298), .B(n14297), .Z(n25784) );
  AND U22750 ( .A(n14302), .B(n14301), .Z(n25780) );
  NAND U22751 ( .A(n14304), .B(n14303), .Z(n25778) );
  AND U22752 ( .A(n14306), .B(n14305), .Z(n25776) );
  AND U22753 ( .A(n14310), .B(n14309), .Z(n25772) );
  AND U22754 ( .A(n14314), .B(n14313), .Z(n25768) );
  AND U22755 ( .A(n14318), .B(n14317), .Z(n25764) );
  XNOR U22756 ( .A(y[638]), .B(x[638]), .Z(n14319) );
  NANDN U22757 ( .A(n14320), .B(n14319), .Z(n25762) );
  AND U22758 ( .A(n14322), .B(n14321), .Z(n25760) );
  AND U22759 ( .A(n14326), .B(n14325), .Z(n25756) );
  AND U22760 ( .A(n14330), .B(n14329), .Z(n25752) );
  AND U22761 ( .A(n14334), .B(n14333), .Z(n25748) );
  AND U22762 ( .A(n14338), .B(n14337), .Z(n25744) );
  AND U22763 ( .A(n14342), .B(n14341), .Z(n25740) );
  XNOR U22764 ( .A(x[626]), .B(y[626]), .Z(n14343) );
  NANDN U22765 ( .A(n14344), .B(n14343), .Z(n25738) );
  NANDN U22766 ( .A(x[624]), .B(y[624]), .Z(n14346) );
  AND U22767 ( .A(n14346), .B(n14345), .Z(n25736) );
  AND U22768 ( .A(n14350), .B(n14349), .Z(n25732) );
  AND U22769 ( .A(n14354), .B(n14353), .Z(n25728) );
  AND U22770 ( .A(n14358), .B(n14357), .Z(n25724) );
  AND U22771 ( .A(n14362), .B(n14361), .Z(n25720) );
  AND U22772 ( .A(n14366), .B(n14365), .Z(n25716) );
  XNOR U22773 ( .A(x[614]), .B(y[614]), .Z(n14367) );
  NANDN U22774 ( .A(n14368), .B(n14367), .Z(n25714) );
  AND U22775 ( .A(n14370), .B(n14369), .Z(n25712) );
  XNOR U22776 ( .A(x[612]), .B(y[612]), .Z(n14371) );
  NANDN U22777 ( .A(n14372), .B(n14371), .Z(n25710) );
  AND U22778 ( .A(n14374), .B(n14373), .Z(n25708) );
  AND U22779 ( .A(n14378), .B(n14377), .Z(n25704) );
  AND U22780 ( .A(n14382), .B(n14381), .Z(n25700) );
  AND U22781 ( .A(n14386), .B(n14385), .Z(n25696) );
  AND U22782 ( .A(n14390), .B(n14389), .Z(n25692) );
  AND U22783 ( .A(n14394), .B(n14393), .Z(n25688) );
  NANDN U22784 ( .A(x[598]), .B(y[598]), .Z(n14397) );
  AND U22785 ( .A(n14398), .B(n14397), .Z(n25684) );
  AND U22786 ( .A(n14402), .B(n14401), .Z(n25680) );
  XNOR U22787 ( .A(y[594]), .B(x[594]), .Z(n14406) );
  NAND U22788 ( .A(n14406), .B(n14405), .Z(n25674) );
  NANDN U22789 ( .A(x[590]), .B(y[590]), .Z(n14407) );
  AND U22790 ( .A(n14408), .B(n14407), .Z(n25668) );
  AND U22791 ( .A(n14412), .B(n14411), .Z(n25664) );
  XNOR U22792 ( .A(x[588]), .B(y[588]), .Z(n14413) );
  NANDN U22793 ( .A(n14414), .B(n14413), .Z(n25662) );
  AND U22794 ( .A(n14416), .B(n14415), .Z(n25660) );
  AND U22795 ( .A(n14420), .B(n14419), .Z(n25656) );
  XNOR U22796 ( .A(y[584]), .B(x[584]), .Z(n14421) );
  NANDN U22797 ( .A(n14422), .B(n14421), .Z(n25654) );
  AND U22798 ( .A(n14424), .B(n14423), .Z(n25652) );
  XNOR U22799 ( .A(x[582]), .B(y[582]), .Z(n14425) );
  NANDN U22800 ( .A(n14426), .B(n14425), .Z(n25650) );
  NANDN U22801 ( .A(x[580]), .B(y[580]), .Z(n14428) );
  AND U22802 ( .A(n14428), .B(n14427), .Z(n25648) );
  AND U22803 ( .A(n14430), .B(n14429), .Z(n25645) );
  XNOR U22804 ( .A(y[578]), .B(x[578]), .Z(n14431) );
  NANDN U22805 ( .A(n14432), .B(n14431), .Z(n25644) );
  NANDN U22806 ( .A(x[574]), .B(y[574]), .Z(n14433) );
  AND U22807 ( .A(n14434), .B(n14433), .Z(n25641) );
  NAND U22808 ( .A(n14436), .B(n14435), .Z(n25640) );
  AND U22809 ( .A(n14438), .B(n14437), .Z(n25639) );
  AND U22810 ( .A(n14442), .B(n14441), .Z(n25637) );
  NANDN U22811 ( .A(x[568]), .B(y[568]), .Z(n14446) );
  AND U22812 ( .A(n14446), .B(n14445), .Z(n25635) );
  AND U22813 ( .A(n14448), .B(n14447), .Z(n25633) );
  XNOR U22814 ( .A(x[566]), .B(y[566]), .Z(n14449) );
  NANDN U22815 ( .A(n14450), .B(n14449), .Z(n25632) );
  AND U22816 ( .A(n14452), .B(n14451), .Z(n25630) );
  AND U22817 ( .A(n14456), .B(n14455), .Z(n25626) );
  AND U22818 ( .A(n14460), .B(n14459), .Z(n25622) );
  XNOR U22819 ( .A(x[560]), .B(y[560]), .Z(n14461) );
  NANDN U22820 ( .A(n14462), .B(n14461), .Z(n25620) );
  NANDN U22821 ( .A(x[558]), .B(y[558]), .Z(n14464) );
  AND U22822 ( .A(n14464), .B(n14463), .Z(n25618) );
  AND U22823 ( .A(n14468), .B(n14467), .Z(n25614) );
  AND U22824 ( .A(n14472), .B(n14471), .Z(n25610) );
  XNOR U22825 ( .A(x[554]), .B(y[554]), .Z(n14473) );
  NANDN U22826 ( .A(n14474), .B(n14473), .Z(n25608) );
  AND U22827 ( .A(n14476), .B(n14475), .Z(n25606) );
  XNOR U22828 ( .A(y[552]), .B(x[552]), .Z(n14477) );
  NANDN U22829 ( .A(n14478), .B(n14477), .Z(n25604) );
  AND U22830 ( .A(n14480), .B(n14479), .Z(n25602) );
  AND U22831 ( .A(n14484), .B(n14483), .Z(n25598) );
  AND U22832 ( .A(n14488), .B(n14487), .Z(n25594) );
  AND U22833 ( .A(n14492), .B(n14491), .Z(n25590) );
  AND U22834 ( .A(n14496), .B(n14495), .Z(n25586) );
  XNOR U22835 ( .A(y[542]), .B(x[542]), .Z(n14497) );
  NANDN U22836 ( .A(n14498), .B(n14497), .Z(n25584) );
  AND U22837 ( .A(n14500), .B(n14499), .Z(n25582) );
  AND U22838 ( .A(n14504), .B(n14503), .Z(n25578) );
  AND U22839 ( .A(n14508), .B(n14507), .Z(n25574) );
  NANDN U22840 ( .A(x[534]), .B(y[534]), .Z(n14512) );
  AND U22841 ( .A(n14512), .B(n14511), .Z(n25570) );
  AND U22842 ( .A(n14516), .B(n14515), .Z(n25566) );
  AND U22843 ( .A(n14520), .B(n14519), .Z(n25562) );
  AND U22844 ( .A(n14524), .B(n14523), .Z(n25558) );
  XNOR U22845 ( .A(x[528]), .B(y[528]), .Z(n14525) );
  NANDN U22846 ( .A(n14526), .B(n14525), .Z(n25556) );
  AND U22847 ( .A(n14528), .B(n14527), .Z(n25554) );
  AND U22848 ( .A(n14532), .B(n14531), .Z(n25550) );
  AND U22849 ( .A(n14536), .B(n14535), .Z(n25548) );
  XNOR U22850 ( .A(x[522]), .B(y[522]), .Z(n14537) );
  NANDN U22851 ( .A(n14538), .B(n14537), .Z(n25547) );
  AND U22852 ( .A(n14540), .B(n14539), .Z(n25546) );
  AND U22853 ( .A(n14544), .B(n14543), .Z(n25544) );
  XNOR U22854 ( .A(y[518]), .B(x[518]), .Z(n14545) );
  NANDN U22855 ( .A(n14546), .B(n14545), .Z(n25543) );
  AND U22856 ( .A(n14548), .B(n14547), .Z(n25542) );
  AND U22857 ( .A(n14552), .B(n14551), .Z(n25540) );
  AND U22858 ( .A(n14556), .B(n14555), .Z(n25538) );
  AND U22859 ( .A(n14560), .B(n14559), .Z(n25536) );
  XNOR U22860 ( .A(y[510]), .B(x[510]), .Z(n14561) );
  NANDN U22861 ( .A(n14562), .B(n14561), .Z(n25535) );
  NANDN U22862 ( .A(x[508]), .B(y[508]), .Z(n14564) );
  AND U22863 ( .A(n14564), .B(n14563), .Z(n25534) );
  AND U22864 ( .A(n14566), .B(n14565), .Z(n25531) );
  AND U22865 ( .A(n14570), .B(n14569), .Z(n25527) );
  AND U22866 ( .A(n14574), .B(n14573), .Z(n25523) );
  AND U22867 ( .A(n14578), .B(n14577), .Z(n25519) );
  AND U22868 ( .A(n14582), .B(n14581), .Z(n25515) );
  AND U22869 ( .A(n14586), .B(n14585), .Z(n25511) );
  AND U22870 ( .A(n14590), .B(n14589), .Z(n25507) );
  AND U22871 ( .A(n14594), .B(n14593), .Z(n25503) );
  AND U22872 ( .A(n14598), .B(n14597), .Z(n25499) );
  IV U22873 ( .A(n14599), .Z(n14601) );
  NAND U22874 ( .A(n14601), .B(n14600), .Z(n25497) );
  AND U22875 ( .A(n14603), .B(n14602), .Z(n25495) );
  AND U22876 ( .A(n14607), .B(n14606), .Z(n25491) );
  XNOR U22877 ( .A(y[486]), .B(x[486]), .Z(n14608) );
  NANDN U22878 ( .A(n14609), .B(n14608), .Z(n25489) );
  AND U22879 ( .A(n14611), .B(n14610), .Z(n25487) );
  AND U22880 ( .A(n14615), .B(n14614), .Z(n25483) );
  AND U22881 ( .A(n14619), .B(n14618), .Z(n25479) );
  AND U22882 ( .A(n14623), .B(n14622), .Z(n25475) );
  AND U22883 ( .A(n14627), .B(n14626), .Z(n25471) );
  AND U22884 ( .A(n14631), .B(n14630), .Z(n25467) );
  AND U22885 ( .A(n14635), .B(n14634), .Z(n25463) );
  AND U22886 ( .A(n14639), .B(n14638), .Z(n25459) );
  AND U22887 ( .A(n14643), .B(n14642), .Z(n25455) );
  AND U22888 ( .A(n14647), .B(n14646), .Z(n25451) );
  AND U22889 ( .A(n14651), .B(n14650), .Z(n25447) );
  XNOR U22890 ( .A(x[464]), .B(y[464]), .Z(n14652) );
  NANDN U22891 ( .A(n14653), .B(n14652), .Z(n25445) );
  AND U22892 ( .A(n14655), .B(n14654), .Z(n25443) );
  AND U22893 ( .A(n14659), .B(n14658), .Z(n25439) );
  AND U22894 ( .A(n14663), .B(n14662), .Z(n25435) );
  AND U22895 ( .A(n14667), .B(n14666), .Z(n25431) );
  XNOR U22896 ( .A(x[456]), .B(y[456]), .Z(n14668) );
  NANDN U22897 ( .A(n14669), .B(n14668), .Z(n25429) );
  AND U22898 ( .A(n14671), .B(n14670), .Z(n25427) );
  AND U22899 ( .A(n14675), .B(n14674), .Z(n25423) );
  AND U22900 ( .A(n14679), .B(n14678), .Z(n25419) );
  XNOR U22901 ( .A(x[450]), .B(y[450]), .Z(n14680) );
  NANDN U22902 ( .A(n14681), .B(n14680), .Z(n25417) );
  AND U22903 ( .A(n14683), .B(n14682), .Z(n25415) );
  AND U22904 ( .A(n14687), .B(n14686), .Z(n25411) );
  AND U22905 ( .A(n14691), .B(n14690), .Z(n25407) );
  AND U22906 ( .A(n14695), .B(n14694), .Z(n25403) );
  AND U22907 ( .A(n14699), .B(n14698), .Z(n25399) );
  AND U22908 ( .A(n14703), .B(n14702), .Z(n25395) );
  XNOR U22909 ( .A(x[438]), .B(y[438]), .Z(n14704) );
  NANDN U22910 ( .A(n14705), .B(n14704), .Z(n25393) );
  AND U22911 ( .A(n14707), .B(n14706), .Z(n25391) );
  AND U22912 ( .A(n14711), .B(n14710), .Z(n25387) );
  XNOR U22913 ( .A(x[434]), .B(y[434]), .Z(n14712) );
  NANDN U22914 ( .A(n14713), .B(n14712), .Z(n25385) );
  AND U22915 ( .A(n14715), .B(n14714), .Z(n25383) );
  AND U22916 ( .A(n14717), .B(n14716), .Z(n25375) );
  XNOR U22917 ( .A(y[428]), .B(x[428]), .Z(n14718) );
  NANDN U22918 ( .A(n14719), .B(n14718), .Z(n25373) );
  AND U22919 ( .A(n14721), .B(n14720), .Z(n25371) );
  XNOR U22920 ( .A(y[426]), .B(x[426]), .Z(n14722) );
  NANDN U22921 ( .A(n14723), .B(n14722), .Z(n25369) );
  AND U22922 ( .A(n14725), .B(n14724), .Z(n25367) );
  AND U22923 ( .A(n14729), .B(n14728), .Z(n25363) );
  NANDN U22924 ( .A(x[418]), .B(y[418]), .Z(n14732) );
  AND U22925 ( .A(n14733), .B(n14732), .Z(n25355) );
  AND U22926 ( .A(n14737), .B(n14736), .Z(n25351) );
  XNOR U22927 ( .A(x[416]), .B(y[416]), .Z(n14738) );
  NANDN U22928 ( .A(n14739), .B(n14738), .Z(n25349) );
  AND U22929 ( .A(n14741), .B(n14740), .Z(n25347) );
  AND U22930 ( .A(n14745), .B(n14744), .Z(n25343) );
  AND U22931 ( .A(n14749), .B(n14748), .Z(n25339) );
  XNOR U22932 ( .A(x[410]), .B(y[410]), .Z(n14750) );
  NANDN U22933 ( .A(n14751), .B(n14750), .Z(n25337) );
  AND U22934 ( .A(n14753), .B(n14752), .Z(n25335) );
  AND U22935 ( .A(n14757), .B(n14756), .Z(n25331) );
  AND U22936 ( .A(n14761), .B(n14760), .Z(n25327) );
  AND U22937 ( .A(n14765), .B(n14764), .Z(n25323) );
  XNOR U22938 ( .A(x[402]), .B(y[402]), .Z(n14766) );
  NANDN U22939 ( .A(n14767), .B(n14766), .Z(n25321) );
  NANDN U22940 ( .A(x[390]), .B(y[390]), .Z(n14768) );
  AND U22941 ( .A(n14769), .B(n14768), .Z(n25299) );
  AND U22942 ( .A(n14773), .B(n14772), .Z(n25295) );
  AND U22943 ( .A(n14777), .B(n14776), .Z(n25291) );
  AND U22944 ( .A(n14781), .B(n14780), .Z(n25287) );
  AND U22945 ( .A(n14785), .B(n14784), .Z(n25283) );
  AND U22946 ( .A(n14789), .B(n14788), .Z(n25279) );
  AND U22947 ( .A(n14793), .B(n14792), .Z(n25275) );
  AND U22948 ( .A(n14797), .B(n14796), .Z(n25271) );
  NAND U22949 ( .A(n14799), .B(n14798), .Z(n25269) );
  AND U22950 ( .A(n14801), .B(n14800), .Z(n25267) );
  AND U22951 ( .A(n14805), .B(n14804), .Z(n25263) );
  AND U22952 ( .A(n14809), .B(n14808), .Z(n25259) );
  AND U22953 ( .A(n14813), .B(n14812), .Z(n25255) );
  XNOR U22954 ( .A(x[368]), .B(y[368]), .Z(n14814) );
  NANDN U22955 ( .A(n14815), .B(n14814), .Z(n25253) );
  AND U22956 ( .A(n14817), .B(n14816), .Z(n25251) );
  AND U22957 ( .A(n14821), .B(n14820), .Z(n25249) );
  AND U22958 ( .A(n14825), .B(n14824), .Z(n25247) );
  XNOR U22959 ( .A(x[362]), .B(y[362]), .Z(n14826) );
  NANDN U22960 ( .A(n14827), .B(n14826), .Z(n25246) );
  AND U22961 ( .A(n14829), .B(n14828), .Z(n25245) );
  XNOR U22962 ( .A(x[360]), .B(y[360]), .Z(n14830) );
  NANDN U22963 ( .A(n14831), .B(n14830), .Z(n25244) );
  AND U22964 ( .A(n14833), .B(n14832), .Z(n25243) );
  AND U22965 ( .A(n14837), .B(n14836), .Z(n25241) );
  AND U22966 ( .A(n14841), .B(n14840), .Z(n25239) );
  XNOR U22967 ( .A(y[354]), .B(x[354]), .Z(n14842) );
  NANDN U22968 ( .A(n14843), .B(n14842), .Z(n25238) );
  NANDN U22969 ( .A(x[352]), .B(y[352]), .Z(n14845) );
  AND U22970 ( .A(n14845), .B(n14844), .Z(n25237) );
  AND U22971 ( .A(n14849), .B(n14848), .Z(n25231) );
  AND U22972 ( .A(n14853), .B(n14852), .Z(n25227) );
  AND U22973 ( .A(n14857), .B(n14856), .Z(n25223) );
  AND U22974 ( .A(n14861), .B(n14860), .Z(n25219) );
  NAND U22975 ( .A(n14867), .B(n14866), .Z(n25205) );
  NAND U22976 ( .A(n14871), .B(n14870), .Z(n25201) );
  NAND U22977 ( .A(n14875), .B(n14874), .Z(n25197) );
  NAND U22978 ( .A(n14879), .B(n14878), .Z(n25193) );
  NAND U22979 ( .A(n14883), .B(n14882), .Z(n25189) );
  NAND U22980 ( .A(n14887), .B(n14886), .Z(n25185) );
  AND U22981 ( .A(n14892), .B(n14891), .Z(n25179) );
  NAND U22982 ( .A(n14894), .B(n14893), .Z(n25177) );
  NAND U22983 ( .A(n14904), .B(n14903), .Z(n25165) );
  NAND U22984 ( .A(n14908), .B(n14907), .Z(n25161) );
  IV U22985 ( .A(n14909), .Z(n14910) );
  AND U22986 ( .A(n14911), .B(n14910), .Z(n25159) );
  NAND U22987 ( .A(n14913), .B(n14912), .Z(n25157) );
  AND U22988 ( .A(n14915), .B(n14914), .Z(n25155) );
  NAND U22989 ( .A(n14917), .B(n14916), .Z(n25153) );
  IV U22990 ( .A(n14920), .Z(n14922) );
  XNOR U22991 ( .A(x[308]), .B(y[308]), .Z(n14921) );
  NANDN U22992 ( .A(n14922), .B(n14921), .Z(n25149) );
  IV U22993 ( .A(n14923), .Z(n14924) );
  AND U22994 ( .A(n14925), .B(n14924), .Z(n25147) );
  NAND U22995 ( .A(n14930), .B(n14929), .Z(n25141) );
  NAND U22996 ( .A(n14937), .B(n14936), .Z(n25133) );
  AND U22997 ( .A(n14939), .B(n14938), .Z(n25131) );
  NAND U22998 ( .A(n14941), .B(n14940), .Z(n25129) );
  NAND U22999 ( .A(n14948), .B(n14947), .Z(n25121) );
  AND U23000 ( .A(n14950), .B(n14949), .Z(n25119) );
  NAND U23001 ( .A(n14952), .B(n14951), .Z(n25117) );
  NAND U23002 ( .A(n14956), .B(n14955), .Z(n25113) );
  IV U23003 ( .A(n14959), .Z(n14961) );
  XNOR U23004 ( .A(x[288]), .B(y[288]), .Z(n14960) );
  NANDN U23005 ( .A(n14961), .B(n14960), .Z(n25109) );
  IV U23006 ( .A(n14962), .Z(n14963) );
  AND U23007 ( .A(n14964), .B(n14963), .Z(n25107) );
  NAND U23008 ( .A(n14966), .B(n14965), .Z(n25105) );
  NAND U23009 ( .A(n14970), .B(n14969), .Z(n25101) );
  NAND U23010 ( .A(n14974), .B(n14973), .Z(n25097) );
  NAND U23011 ( .A(n14978), .B(n14977), .Z(n25093) );
  NAND U23012 ( .A(n14985), .B(n14984), .Z(n25085) );
  NAND U23013 ( .A(n14989), .B(n14988), .Z(n25081) );
  NAND U23014 ( .A(n14993), .B(n14992), .Z(n25077) );
  IV U23015 ( .A(n14994), .Z(n25075) );
  IV U23016 ( .A(n14995), .Z(n25068) );
  IV U23017 ( .A(n14996), .Z(n25066) );
  IV U23018 ( .A(n14997), .Z(n25065) );
  IV U23019 ( .A(n14998), .Z(n25063) );
  NANDN U23020 ( .A(y[262]), .B(x[262]), .Z(n15001) );
  NAND U23021 ( .A(n15001), .B(n15000), .Z(n25057) );
  NAND U23022 ( .A(n15008), .B(n15007), .Z(n25049) );
  NAND U23023 ( .A(n15012), .B(n15011), .Z(n25045) );
  NAND U23024 ( .A(n15019), .B(n15018), .Z(n25037) );
  NAND U23025 ( .A(n15023), .B(n15022), .Z(n25033) );
  NAND U23026 ( .A(n15027), .B(n15026), .Z(n25029) );
  AND U23027 ( .A(n15029), .B(n15028), .Z(n25027) );
  NAND U23028 ( .A(n15031), .B(n15030), .Z(n25025) );
  NAND U23029 ( .A(n15035), .B(n15034), .Z(n25021) );
  AND U23030 ( .A(n15040), .B(n15039), .Z(n25015) );
  NAND U23031 ( .A(n15042), .B(n15041), .Z(n25013) );
  NAND U23032 ( .A(n15046), .B(n15045), .Z(n25009) );
  NAND U23033 ( .A(n15050), .B(n15049), .Z(n25005) );
  NAND U23034 ( .A(n15054), .B(n15053), .Z(n25001) );
  NAND U23035 ( .A(n15058), .B(n15057), .Z(n24997) );
  NAND U23036 ( .A(n15065), .B(n15064), .Z(n24989) );
  IV U23037 ( .A(n15066), .Z(n15067) );
  AND U23038 ( .A(n15068), .B(n15067), .Z(n24987) );
  NAND U23039 ( .A(n15070), .B(n15069), .Z(n24985) );
  NAND U23040 ( .A(n15074), .B(n15073), .Z(n24981) );
  NAND U23041 ( .A(n15078), .B(n15077), .Z(n24977) );
  NAND U23042 ( .A(n15082), .B(n15081), .Z(n24973) );
  NAND U23043 ( .A(n15086), .B(n15085), .Z(n24969) );
  NAND U23044 ( .A(n15090), .B(n15089), .Z(n24965) );
  NAND U23045 ( .A(n15094), .B(n15093), .Z(n24961) );
  NAND U23046 ( .A(n15098), .B(n15097), .Z(n24957) );
  NAND U23047 ( .A(n15105), .B(n15104), .Z(n24949) );
  IV U23048 ( .A(n15106), .Z(n15107) );
  AND U23049 ( .A(n15108), .B(n15107), .Z(n24947) );
  NAND U23050 ( .A(n15110), .B(n15109), .Z(n24945) );
  NAND U23051 ( .A(n15114), .B(n15113), .Z(n24941) );
  NAND U23052 ( .A(n15118), .B(n15117), .Z(n24937) );
  NAND U23053 ( .A(n15122), .B(n15121), .Z(n24933) );
  NAND U23054 ( .A(n15129), .B(n15128), .Z(n24925) );
  NAND U23055 ( .A(n15133), .B(n15132), .Z(n24921) );
  NAND U23056 ( .A(n15137), .B(n15136), .Z(n24917) );
  NAND U23057 ( .A(n15141), .B(n15140), .Z(n24913) );
  NAND U23058 ( .A(n15145), .B(n15144), .Z(n24909) );
  IV U23059 ( .A(n15146), .Z(n15147) );
  AND U23060 ( .A(n15148), .B(n15147), .Z(n24907) );
  NAND U23061 ( .A(n15150), .B(n15149), .Z(n24905) );
  NAND U23062 ( .A(n15154), .B(n15153), .Z(n24901) );
  NAND U23063 ( .A(n15164), .B(n15163), .Z(n24889) );
  IV U23064 ( .A(n15167), .Z(n15169) );
  XNOR U23065 ( .A(y[176]), .B(x[176]), .Z(n15168) );
  NANDN U23066 ( .A(n15169), .B(n15168), .Z(n24885) );
  IV U23067 ( .A(n15170), .Z(n15171) );
  AND U23068 ( .A(n15172), .B(n15171), .Z(n24883) );
  IV U23069 ( .A(n15173), .Z(n15175) );
  XNOR U23070 ( .A(x[174]), .B(y[174]), .Z(n15174) );
  NANDN U23071 ( .A(n15175), .B(n15174), .Z(n24881) );
  IV U23072 ( .A(n15176), .Z(n15177) );
  AND U23073 ( .A(n15178), .B(n15177), .Z(n24879) );
  NAND U23074 ( .A(n15180), .B(n15179), .Z(n24877) );
  NAND U23075 ( .A(n15187), .B(n15186), .Z(n24869) );
  IV U23076 ( .A(n15188), .Z(n15189) );
  AND U23077 ( .A(n15190), .B(n15189), .Z(n24867) );
  NAND U23078 ( .A(n15192), .B(n15191), .Z(n24865) );
  NAND U23079 ( .A(n15196), .B(n15195), .Z(n24861) );
  NAND U23080 ( .A(n15200), .B(n15199), .Z(n24857) );
  NAND U23081 ( .A(n15204), .B(n15203), .Z(n24853) );
  NAND U23082 ( .A(n15208), .B(n15207), .Z(n24849) );
  AND U23083 ( .A(n15210), .B(n15209), .Z(n24847) );
  NAND U23084 ( .A(n15212), .B(n15211), .Z(n24845) );
  NAND U23085 ( .A(n15216), .B(n15215), .Z(n24841) );
  NAND U23086 ( .A(n15220), .B(n15219), .Z(n24837) );
  NAND U23087 ( .A(n15227), .B(n15226), .Z(n24829) );
  NANDN U23088 ( .A(y[141]), .B(x[141]), .Z(n15233) );
  AND U23089 ( .A(n15234), .B(n15233), .Z(n24816) );
  AND U23090 ( .A(n15236), .B(n15235), .Z(n24815) );
  NAND U23091 ( .A(n15238), .B(n15237), .Z(n24813) );
  NAND U23092 ( .A(n15242), .B(n15241), .Z(n24809) );
  NAND U23093 ( .A(n15246), .B(n15245), .Z(n24805) );
  AND U23094 ( .A(n15248), .B(n15247), .Z(n24803) );
  NAND U23095 ( .A(n15250), .B(n15249), .Z(n24801) );
  NAND U23096 ( .A(n15254), .B(n15253), .Z(n24797) );
  NAND U23097 ( .A(n15258), .B(n15257), .Z(n24793) );
  NAND U23098 ( .A(n15265), .B(n15264), .Z(n24785) );
  NAND U23099 ( .A(n15269), .B(n15268), .Z(n24781) );
  NAND U23100 ( .A(n15273), .B(n15272), .Z(n24777) );
  NAND U23101 ( .A(n15277), .B(n15276), .Z(n24773) );
  NAND U23102 ( .A(n15281), .B(n15280), .Z(n24769) );
  NAND U23103 ( .A(n15285), .B(n15284), .Z(n24765) );
  IV U23104 ( .A(n15288), .Z(n15290) );
  XNOR U23105 ( .A(x[114]), .B(y[114]), .Z(n15289) );
  NANDN U23106 ( .A(n15290), .B(n15289), .Z(n24761) );
  IV U23107 ( .A(n15291), .Z(n15292) );
  AND U23108 ( .A(n15293), .B(n15292), .Z(n24759) );
  NAND U23109 ( .A(n15295), .B(n15294), .Z(n24757) );
  NAND U23110 ( .A(n15299), .B(n15298), .Z(n24753) );
  NAND U23111 ( .A(n15303), .B(n15302), .Z(n24749) );
  NAND U23112 ( .A(n15307), .B(n15306), .Z(n24745) );
  AND U23113 ( .A(n15309), .B(n15308), .Z(n24743) );
  NAND U23114 ( .A(n15311), .B(n15310), .Z(n24741) );
  AND U23115 ( .A(n15317), .B(n15316), .Z(n24731) );
  NANDN U23116 ( .A(x[96]), .B(y[96]), .Z(n15321) );
  AND U23117 ( .A(n15321), .B(n15320), .Z(n24727) );
  AND U23118 ( .A(n15325), .B(n15324), .Z(n24723) );
  AND U23119 ( .A(n15329), .B(n15328), .Z(n24719) );
  NAND U23120 ( .A(n15331), .B(n15330), .Z(n24717) );
  AND U23121 ( .A(n15333), .B(n15332), .Z(n24715) );
  AND U23122 ( .A(n15337), .B(n15336), .Z(n24711) );
  AND U23123 ( .A(n15341), .B(n15340), .Z(n24707) );
  AND U23124 ( .A(n15345), .B(n15344), .Z(n24703) );
  XNOR U23125 ( .A(x[84]), .B(y[84]), .Z(n15346) );
  NANDN U23126 ( .A(n15347), .B(n15346), .Z(n24701) );
  AND U23127 ( .A(n15349), .B(n15348), .Z(n24699) );
  AND U23128 ( .A(n15353), .B(n15352), .Z(n24695) );
  XNOR U23129 ( .A(x[80]), .B(y[80]), .Z(n15354) );
  NANDN U23130 ( .A(n15355), .B(n15354), .Z(n24693) );
  NANDN U23131 ( .A(x[76]), .B(y[76]), .Z(n15356) );
  AND U23132 ( .A(n15357), .B(n15356), .Z(n24687) );
  AND U23133 ( .A(n15361), .B(n15360), .Z(n24683) );
  AND U23134 ( .A(n15365), .B(n15364), .Z(n24679) );
  NANDN U23135 ( .A(x[69]), .B(y[69]), .Z(n15368) );
  AND U23136 ( .A(n15368), .B(n15367), .Z(n24671) );
  AND U23137 ( .A(n15372), .B(n15371), .Z(n24667) );
  NANDN U23138 ( .A(x[60]), .B(y[60]), .Z(n15375) );
  AND U23139 ( .A(n15376), .B(n15375), .Z(n24655) );
  AND U23140 ( .A(n15380), .B(n15379), .Z(n24651) );
  AND U23141 ( .A(n15384), .B(n15383), .Z(n24647) );
  AND U23142 ( .A(n15388), .B(n15387), .Z(n24643) );
  XNOR U23143 ( .A(x[54]), .B(y[54]), .Z(n15389) );
  NANDN U23144 ( .A(n15390), .B(n15389), .Z(n24641) );
  AND U23145 ( .A(n15392), .B(n15391), .Z(n24639) );
  AND U23146 ( .A(n15396), .B(n15395), .Z(n24635) );
  AND U23147 ( .A(n15400), .B(n15399), .Z(n24631) );
  AND U23148 ( .A(n15404), .B(n15403), .Z(n24627) );
  AND U23149 ( .A(n15408), .B(n15407), .Z(n24623) );
  AND U23150 ( .A(n15412), .B(n15411), .Z(n24619) );
  AND U23151 ( .A(n15416), .B(n15415), .Z(n24615) );
  AND U23152 ( .A(n15420), .B(n15419), .Z(n24611) );
  XNOR U23153 ( .A(x[38]), .B(y[38]), .Z(n15421) );
  NANDN U23154 ( .A(n15422), .B(n15421), .Z(n24609) );
  NANDN U23155 ( .A(x[36]), .B(y[36]), .Z(n15424) );
  AND U23156 ( .A(n15424), .B(n15423), .Z(n24607) );
  AND U23157 ( .A(n15428), .B(n15427), .Z(n24603) );
  AND U23158 ( .A(n15432), .B(n15431), .Z(n24599) );
  XNOR U23159 ( .A(x[32]), .B(y[32]), .Z(n15433) );
  NANDN U23160 ( .A(n15434), .B(n15433), .Z(n24597) );
  NANDN U23161 ( .A(x[30]), .B(y[30]), .Z(n15436) );
  AND U23162 ( .A(n15436), .B(n15435), .Z(n24595) );
  AND U23163 ( .A(n15440), .B(n15439), .Z(n24591) );
  AND U23164 ( .A(n15444), .B(n15443), .Z(n24587) );
  XNOR U23165 ( .A(x[26]), .B(y[26]), .Z(n15445) );
  NANDN U23166 ( .A(n15446), .B(n15445), .Z(n24585) );
  AND U23167 ( .A(n15448), .B(n15447), .Z(n24583) );
  AND U23168 ( .A(n15452), .B(n15451), .Z(n24579) );
  AND U23169 ( .A(n15456), .B(n15455), .Z(n24575) );
  AND U23170 ( .A(n15460), .B(n15459), .Z(n24571) );
  AND U23171 ( .A(n15464), .B(n15463), .Z(n24567) );
  AND U23172 ( .A(n15468), .B(n15467), .Z(n24563) );
  AND U23173 ( .A(n15472), .B(n15471), .Z(n24559) );
  AND U23174 ( .A(n15476), .B(n15475), .Z(n24555) );
  AND U23175 ( .A(n15480), .B(n15479), .Z(n24551) );
  NAND U23176 ( .A(n15482), .B(n15481), .Z(n24549) );
  AND U23177 ( .A(n15484), .B(n15483), .Z(n24547) );
  AND U23178 ( .A(n15488), .B(n15487), .Z(n24543) );
  NANDN U23179 ( .A(x[0]), .B(y[0]), .Z(n15491) );
  NAND U23180 ( .A(n15492), .B(n15491), .Z(n15493) );
  NANDN U23181 ( .A(n15494), .B(n15493), .Z(n15495) );
  NAND U23182 ( .A(n15496), .B(n15495), .Z(n15497) );
  NANDN U23183 ( .A(n24541), .B(n15497), .Z(n15498) );
  AND U23184 ( .A(n24543), .B(n15498), .Z(n15499) );
  OR U23185 ( .A(n24545), .B(n15499), .Z(n15500) );
  NAND U23186 ( .A(n24547), .B(n15500), .Z(n15501) );
  NANDN U23187 ( .A(n24549), .B(n15501), .Z(n15502) );
  NAND U23188 ( .A(n24551), .B(n15502), .Z(n15503) );
  NANDN U23189 ( .A(n24553), .B(n15503), .Z(n15504) );
  AND U23190 ( .A(n24555), .B(n15504), .Z(n15505) );
  OR U23191 ( .A(n24557), .B(n15505), .Z(n15506) );
  NAND U23192 ( .A(n24559), .B(n15506), .Z(n15507) );
  NANDN U23193 ( .A(n24561), .B(n15507), .Z(n15508) );
  NAND U23194 ( .A(n24563), .B(n15508), .Z(n15509) );
  NANDN U23195 ( .A(n24565), .B(n15509), .Z(n15510) );
  AND U23196 ( .A(n24567), .B(n15510), .Z(n15511) );
  OR U23197 ( .A(n24569), .B(n15511), .Z(n15512) );
  NAND U23198 ( .A(n24571), .B(n15512), .Z(n15513) );
  NANDN U23199 ( .A(n24573), .B(n15513), .Z(n15514) );
  NAND U23200 ( .A(n24575), .B(n15514), .Z(n15515) );
  NANDN U23201 ( .A(n24577), .B(n15515), .Z(n15516) );
  AND U23202 ( .A(n24579), .B(n15516), .Z(n15517) );
  OR U23203 ( .A(n24581), .B(n15517), .Z(n15518) );
  NAND U23204 ( .A(n24583), .B(n15518), .Z(n15519) );
  NANDN U23205 ( .A(n24585), .B(n15519), .Z(n15520) );
  NAND U23206 ( .A(n24587), .B(n15520), .Z(n15521) );
  NANDN U23207 ( .A(n24589), .B(n15521), .Z(n15522) );
  AND U23208 ( .A(n24591), .B(n15522), .Z(n15523) );
  OR U23209 ( .A(n24593), .B(n15523), .Z(n15524) );
  NAND U23210 ( .A(n24595), .B(n15524), .Z(n15525) );
  NANDN U23211 ( .A(n24597), .B(n15525), .Z(n15526) );
  NAND U23212 ( .A(n24599), .B(n15526), .Z(n15527) );
  NANDN U23213 ( .A(n24601), .B(n15527), .Z(n15528) );
  AND U23214 ( .A(n24603), .B(n15528), .Z(n15529) );
  OR U23215 ( .A(n24605), .B(n15529), .Z(n15530) );
  NAND U23216 ( .A(n24607), .B(n15530), .Z(n15531) );
  NANDN U23217 ( .A(n24609), .B(n15531), .Z(n15532) );
  NAND U23218 ( .A(n24611), .B(n15532), .Z(n15533) );
  NANDN U23219 ( .A(n24613), .B(n15533), .Z(n15534) );
  AND U23220 ( .A(n24615), .B(n15534), .Z(n15535) );
  OR U23221 ( .A(n24617), .B(n15535), .Z(n15536) );
  NAND U23222 ( .A(n24619), .B(n15536), .Z(n15537) );
  NANDN U23223 ( .A(n24621), .B(n15537), .Z(n15538) );
  NAND U23224 ( .A(n24623), .B(n15538), .Z(n15539) );
  NANDN U23225 ( .A(n24625), .B(n15539), .Z(n15540) );
  AND U23226 ( .A(n24627), .B(n15540), .Z(n15541) );
  OR U23227 ( .A(n24629), .B(n15541), .Z(n15542) );
  NAND U23228 ( .A(n24631), .B(n15542), .Z(n15543) );
  NANDN U23229 ( .A(n24633), .B(n15543), .Z(n15544) );
  NAND U23230 ( .A(n24635), .B(n15544), .Z(n15545) );
  NANDN U23231 ( .A(n24637), .B(n15545), .Z(n15546) );
  AND U23232 ( .A(n24639), .B(n15546), .Z(n15547) );
  OR U23233 ( .A(n24641), .B(n15547), .Z(n15548) );
  NAND U23234 ( .A(n24643), .B(n15548), .Z(n15549) );
  NANDN U23235 ( .A(n24645), .B(n15549), .Z(n15550) );
  NAND U23236 ( .A(n24647), .B(n15550), .Z(n15551) );
  NANDN U23237 ( .A(n24649), .B(n15551), .Z(n15552) );
  AND U23238 ( .A(n24651), .B(n15552), .Z(n15553) );
  OR U23239 ( .A(n24653), .B(n15553), .Z(n15554) );
  NAND U23240 ( .A(n24655), .B(n15554), .Z(n15555) );
  NANDN U23241 ( .A(n24657), .B(n15555), .Z(n15556) );
  NAND U23242 ( .A(n24659), .B(n15556), .Z(n15557) );
  NANDN U23243 ( .A(n24661), .B(n15557), .Z(n15558) );
  AND U23244 ( .A(n24663), .B(n15558), .Z(n15559) );
  OR U23245 ( .A(n24665), .B(n15559), .Z(n15560) );
  NAND U23246 ( .A(n24667), .B(n15560), .Z(n15561) );
  NANDN U23247 ( .A(n24669), .B(n15561), .Z(n15562) );
  NAND U23248 ( .A(n24671), .B(n15562), .Z(n15563) );
  NAND U23249 ( .A(n24672), .B(n15563), .Z(n15564) );
  AND U23250 ( .A(n24675), .B(n15564), .Z(n15565) );
  OR U23251 ( .A(n24677), .B(n15565), .Z(n15566) );
  NAND U23252 ( .A(n24679), .B(n15566), .Z(n15567) );
  NANDN U23253 ( .A(n24681), .B(n15567), .Z(n15568) );
  NAND U23254 ( .A(n24683), .B(n15568), .Z(n15569) );
  NANDN U23255 ( .A(n24685), .B(n15569), .Z(n15570) );
  AND U23256 ( .A(n24687), .B(n15570), .Z(n15571) );
  OR U23257 ( .A(n24689), .B(n15571), .Z(n15572) );
  NAND U23258 ( .A(n24691), .B(n15572), .Z(n15573) );
  NANDN U23259 ( .A(n24693), .B(n15573), .Z(n15574) );
  NAND U23260 ( .A(n24695), .B(n15574), .Z(n15575) );
  NANDN U23261 ( .A(n24697), .B(n15575), .Z(n15576) );
  AND U23262 ( .A(n24699), .B(n15576), .Z(n15577) );
  OR U23263 ( .A(n24701), .B(n15577), .Z(n15578) );
  NAND U23264 ( .A(n24703), .B(n15578), .Z(n15579) );
  NANDN U23265 ( .A(n24705), .B(n15579), .Z(n15580) );
  NAND U23266 ( .A(n24707), .B(n15580), .Z(n15581) );
  NANDN U23267 ( .A(n24709), .B(n15581), .Z(n15582) );
  AND U23268 ( .A(n24711), .B(n15582), .Z(n15583) );
  OR U23269 ( .A(n24713), .B(n15583), .Z(n15584) );
  NAND U23270 ( .A(n24715), .B(n15584), .Z(n15585) );
  NANDN U23271 ( .A(n24717), .B(n15585), .Z(n15586) );
  NAND U23272 ( .A(n24719), .B(n15586), .Z(n15587) );
  NANDN U23273 ( .A(n24721), .B(n15587), .Z(n15588) );
  AND U23274 ( .A(n24723), .B(n15588), .Z(n15589) );
  OR U23275 ( .A(n24725), .B(n15589), .Z(n15590) );
  NAND U23276 ( .A(n24727), .B(n15590), .Z(n15591) );
  NANDN U23277 ( .A(n24729), .B(n15591), .Z(n15592) );
  NAND U23278 ( .A(n24731), .B(n15592), .Z(n15593) );
  NANDN U23279 ( .A(n24733), .B(n15593), .Z(n15594) );
  AND U23280 ( .A(n24735), .B(n15594), .Z(n15596) );
  IV U23281 ( .A(n15595), .Z(n24737) );
  OR U23282 ( .A(n15596), .B(n24737), .Z(n15597) );
  NAND U23283 ( .A(n24739), .B(n15597), .Z(n15598) );
  NANDN U23284 ( .A(n24741), .B(n15598), .Z(n15599) );
  NAND U23285 ( .A(n24743), .B(n15599), .Z(n15600) );
  NANDN U23286 ( .A(n24745), .B(n15600), .Z(n15601) );
  AND U23287 ( .A(n24747), .B(n15601), .Z(n15602) );
  OR U23288 ( .A(n24749), .B(n15602), .Z(n15603) );
  NAND U23289 ( .A(n24751), .B(n15603), .Z(n15604) );
  NANDN U23290 ( .A(n24753), .B(n15604), .Z(n15605) );
  NAND U23291 ( .A(n24755), .B(n15605), .Z(n15606) );
  NANDN U23292 ( .A(n24757), .B(n15606), .Z(n15607) );
  AND U23293 ( .A(n24759), .B(n15607), .Z(n15608) );
  OR U23294 ( .A(n24761), .B(n15608), .Z(n15609) );
  NAND U23295 ( .A(n24763), .B(n15609), .Z(n15610) );
  NANDN U23296 ( .A(n24765), .B(n15610), .Z(n15611) );
  NAND U23297 ( .A(n24767), .B(n15611), .Z(n15612) );
  NANDN U23298 ( .A(n24769), .B(n15612), .Z(n15613) );
  AND U23299 ( .A(n24771), .B(n15613), .Z(n15614) );
  OR U23300 ( .A(n24773), .B(n15614), .Z(n15615) );
  NAND U23301 ( .A(n24775), .B(n15615), .Z(n15616) );
  NANDN U23302 ( .A(n24777), .B(n15616), .Z(n15617) );
  NAND U23303 ( .A(n24779), .B(n15617), .Z(n15618) );
  NANDN U23304 ( .A(n24781), .B(n15618), .Z(n15619) );
  AND U23305 ( .A(n24783), .B(n15619), .Z(n15620) );
  OR U23306 ( .A(n24785), .B(n15620), .Z(n15621) );
  NAND U23307 ( .A(n24787), .B(n15621), .Z(n15622) );
  NANDN U23308 ( .A(n24789), .B(n15622), .Z(n15623) );
  NAND U23309 ( .A(n24791), .B(n15623), .Z(n15624) );
  NANDN U23310 ( .A(n24793), .B(n15624), .Z(n15625) );
  AND U23311 ( .A(n24795), .B(n15625), .Z(n15626) );
  OR U23312 ( .A(n24797), .B(n15626), .Z(n15627) );
  NAND U23313 ( .A(n24799), .B(n15627), .Z(n15628) );
  NANDN U23314 ( .A(n24801), .B(n15628), .Z(n15629) );
  NAND U23315 ( .A(n24803), .B(n15629), .Z(n15630) );
  NANDN U23316 ( .A(n24805), .B(n15630), .Z(n15631) );
  AND U23317 ( .A(n24807), .B(n15631), .Z(n15632) );
  OR U23318 ( .A(n24809), .B(n15632), .Z(n15633) );
  NAND U23319 ( .A(n24811), .B(n15633), .Z(n15634) );
  NANDN U23320 ( .A(n24813), .B(n15634), .Z(n15635) );
  NAND U23321 ( .A(n24815), .B(n15635), .Z(n15636) );
  NAND U23322 ( .A(n24816), .B(n15636), .Z(n15638) );
  IV U23323 ( .A(n15637), .Z(n24819) );
  AND U23324 ( .A(n15638), .B(n24819), .Z(n15640) );
  IV U23325 ( .A(n15639), .Z(n24821) );
  OR U23326 ( .A(n15640), .B(n24821), .Z(n15641) );
  NAND U23327 ( .A(n24823), .B(n15641), .Z(n15642) );
  NANDN U23328 ( .A(n24825), .B(n15642), .Z(n15643) );
  NAND U23329 ( .A(n24827), .B(n15643), .Z(n15644) );
  NANDN U23330 ( .A(n24829), .B(n15644), .Z(n15645) );
  AND U23331 ( .A(n24831), .B(n15645), .Z(n15646) );
  OR U23332 ( .A(n24833), .B(n15646), .Z(n15647) );
  NAND U23333 ( .A(n24835), .B(n15647), .Z(n15648) );
  NANDN U23334 ( .A(n24837), .B(n15648), .Z(n15649) );
  NAND U23335 ( .A(n24839), .B(n15649), .Z(n15650) );
  NANDN U23336 ( .A(n24841), .B(n15650), .Z(n15651) );
  AND U23337 ( .A(n24843), .B(n15651), .Z(n15652) );
  OR U23338 ( .A(n24845), .B(n15652), .Z(n15653) );
  NAND U23339 ( .A(n24847), .B(n15653), .Z(n15654) );
  NANDN U23340 ( .A(n24849), .B(n15654), .Z(n15655) );
  NAND U23341 ( .A(n24851), .B(n15655), .Z(n15656) );
  NANDN U23342 ( .A(n24853), .B(n15656), .Z(n15657) );
  AND U23343 ( .A(n24855), .B(n15657), .Z(n15658) );
  OR U23344 ( .A(n24857), .B(n15658), .Z(n15659) );
  NAND U23345 ( .A(n24859), .B(n15659), .Z(n15660) );
  NANDN U23346 ( .A(n24861), .B(n15660), .Z(n15661) );
  NAND U23347 ( .A(n24863), .B(n15661), .Z(n15662) );
  NANDN U23348 ( .A(n24865), .B(n15662), .Z(n15663) );
  AND U23349 ( .A(n24867), .B(n15663), .Z(n15664) );
  OR U23350 ( .A(n24869), .B(n15664), .Z(n15665) );
  NAND U23351 ( .A(n24871), .B(n15665), .Z(n15666) );
  NANDN U23352 ( .A(n24873), .B(n15666), .Z(n15667) );
  NAND U23353 ( .A(n24875), .B(n15667), .Z(n15668) );
  NANDN U23354 ( .A(n24877), .B(n15668), .Z(n15669) );
  AND U23355 ( .A(n24879), .B(n15669), .Z(n15670) );
  OR U23356 ( .A(n24881), .B(n15670), .Z(n15671) );
  NAND U23357 ( .A(n24883), .B(n15671), .Z(n15672) );
  NANDN U23358 ( .A(n24885), .B(n15672), .Z(n15673) );
  NAND U23359 ( .A(n24887), .B(n15673), .Z(n15674) );
  NANDN U23360 ( .A(n24889), .B(n15674), .Z(n15675) );
  AND U23361 ( .A(n24891), .B(n15675), .Z(n15676) );
  OR U23362 ( .A(n24893), .B(n15676), .Z(n15677) );
  NAND U23363 ( .A(n24895), .B(n15677), .Z(n15678) );
  NANDN U23364 ( .A(n24897), .B(n15678), .Z(n15679) );
  NAND U23365 ( .A(n24899), .B(n15679), .Z(n15680) );
  NANDN U23366 ( .A(n24901), .B(n15680), .Z(n15681) );
  AND U23367 ( .A(n24903), .B(n15681), .Z(n15682) );
  OR U23368 ( .A(n24905), .B(n15682), .Z(n15683) );
  NAND U23369 ( .A(n24907), .B(n15683), .Z(n15684) );
  NANDN U23370 ( .A(n24909), .B(n15684), .Z(n15685) );
  NAND U23371 ( .A(n24911), .B(n15685), .Z(n15686) );
  NANDN U23372 ( .A(n24913), .B(n15686), .Z(n15687) );
  AND U23373 ( .A(n24915), .B(n15687), .Z(n15688) );
  OR U23374 ( .A(n24917), .B(n15688), .Z(n15689) );
  NAND U23375 ( .A(n24919), .B(n15689), .Z(n15690) );
  NANDN U23376 ( .A(n24921), .B(n15690), .Z(n15691) );
  NAND U23377 ( .A(n24923), .B(n15691), .Z(n15692) );
  NANDN U23378 ( .A(n24925), .B(n15692), .Z(n15693) );
  AND U23379 ( .A(n24927), .B(n15693), .Z(n15694) );
  OR U23380 ( .A(n24929), .B(n15694), .Z(n15695) );
  NAND U23381 ( .A(n24931), .B(n15695), .Z(n15696) );
  NANDN U23382 ( .A(n24933), .B(n15696), .Z(n15697) );
  NAND U23383 ( .A(n24935), .B(n15697), .Z(n15698) );
  NANDN U23384 ( .A(n24937), .B(n15698), .Z(n15699) );
  AND U23385 ( .A(n24939), .B(n15699), .Z(n15700) );
  OR U23386 ( .A(n24941), .B(n15700), .Z(n15701) );
  NAND U23387 ( .A(n24943), .B(n15701), .Z(n15702) );
  NANDN U23388 ( .A(n24945), .B(n15702), .Z(n15703) );
  NAND U23389 ( .A(n24947), .B(n15703), .Z(n15704) );
  NANDN U23390 ( .A(n24949), .B(n15704), .Z(n15705) );
  AND U23391 ( .A(n24951), .B(n15705), .Z(n15706) );
  OR U23392 ( .A(n24953), .B(n15706), .Z(n15707) );
  NAND U23393 ( .A(n24955), .B(n15707), .Z(n15708) );
  NANDN U23394 ( .A(n24957), .B(n15708), .Z(n15709) );
  NAND U23395 ( .A(n24959), .B(n15709), .Z(n15710) );
  NANDN U23396 ( .A(n24961), .B(n15710), .Z(n15711) );
  AND U23397 ( .A(n24963), .B(n15711), .Z(n15712) );
  OR U23398 ( .A(n24965), .B(n15712), .Z(n15713) );
  NAND U23399 ( .A(n24967), .B(n15713), .Z(n15714) );
  NANDN U23400 ( .A(n24969), .B(n15714), .Z(n15715) );
  NAND U23401 ( .A(n24971), .B(n15715), .Z(n15716) );
  NANDN U23402 ( .A(n24973), .B(n15716), .Z(n15717) );
  AND U23403 ( .A(n24975), .B(n15717), .Z(n15718) );
  OR U23404 ( .A(n24977), .B(n15718), .Z(n15719) );
  NAND U23405 ( .A(n24979), .B(n15719), .Z(n15720) );
  NANDN U23406 ( .A(n24981), .B(n15720), .Z(n15721) );
  NAND U23407 ( .A(n24983), .B(n15721), .Z(n15722) );
  NANDN U23408 ( .A(n24985), .B(n15722), .Z(n15723) );
  AND U23409 ( .A(n24987), .B(n15723), .Z(n15724) );
  OR U23410 ( .A(n24989), .B(n15724), .Z(n15725) );
  NAND U23411 ( .A(n24991), .B(n15725), .Z(n15726) );
  NANDN U23412 ( .A(n24993), .B(n15726), .Z(n15727) );
  NAND U23413 ( .A(n24995), .B(n15727), .Z(n15728) );
  NANDN U23414 ( .A(n24997), .B(n15728), .Z(n15729) );
  AND U23415 ( .A(n24999), .B(n15729), .Z(n15730) );
  OR U23416 ( .A(n25001), .B(n15730), .Z(n15731) );
  NAND U23417 ( .A(n25003), .B(n15731), .Z(n15732) );
  NANDN U23418 ( .A(n25005), .B(n15732), .Z(n15733) );
  NAND U23419 ( .A(n25007), .B(n15733), .Z(n15734) );
  NANDN U23420 ( .A(n25009), .B(n15734), .Z(n15735) );
  AND U23421 ( .A(n25011), .B(n15735), .Z(n15736) );
  OR U23422 ( .A(n25013), .B(n15736), .Z(n15737) );
  NAND U23423 ( .A(n25015), .B(n15737), .Z(n15738) );
  NANDN U23424 ( .A(n25017), .B(n15738), .Z(n15739) );
  NAND U23425 ( .A(n25019), .B(n15739), .Z(n15740) );
  NANDN U23426 ( .A(n25021), .B(n15740), .Z(n15741) );
  AND U23427 ( .A(n25023), .B(n15741), .Z(n15742) );
  OR U23428 ( .A(n25025), .B(n15742), .Z(n15743) );
  NAND U23429 ( .A(n25027), .B(n15743), .Z(n15744) );
  NANDN U23430 ( .A(n25029), .B(n15744), .Z(n15745) );
  NAND U23431 ( .A(n25031), .B(n15745), .Z(n15746) );
  NANDN U23432 ( .A(n25033), .B(n15746), .Z(n15747) );
  AND U23433 ( .A(n25035), .B(n15747), .Z(n15748) );
  OR U23434 ( .A(n25037), .B(n15748), .Z(n15749) );
  NAND U23435 ( .A(n25039), .B(n15749), .Z(n15750) );
  NANDN U23436 ( .A(n25041), .B(n15750), .Z(n15751) );
  NAND U23437 ( .A(n25043), .B(n15751), .Z(n15752) );
  NANDN U23438 ( .A(n25045), .B(n15752), .Z(n15753) );
  AND U23439 ( .A(n25047), .B(n15753), .Z(n15754) );
  OR U23440 ( .A(n25049), .B(n15754), .Z(n15755) );
  NAND U23441 ( .A(n25051), .B(n15755), .Z(n15756) );
  NANDN U23442 ( .A(n25053), .B(n15756), .Z(n15757) );
  NAND U23443 ( .A(n25055), .B(n15757), .Z(n15758) );
  NANDN U23444 ( .A(n25057), .B(n15758), .Z(n15759) );
  AND U23445 ( .A(n25059), .B(n15759), .Z(n15761) );
  IV U23446 ( .A(n15760), .Z(n25061) );
  OR U23447 ( .A(n15761), .B(n25061), .Z(n15762) );
  NAND U23448 ( .A(n25063), .B(n15762), .Z(n15763) );
  NANDN U23449 ( .A(n25065), .B(n15763), .Z(n15764) );
  NAND U23450 ( .A(n25066), .B(n15764), .Z(n15765) );
  NANDN U23451 ( .A(n25068), .B(n15765), .Z(n15767) );
  IV U23452 ( .A(n15766), .Z(n25071) );
  AND U23453 ( .A(n15767), .B(n25071), .Z(n15769) );
  IV U23454 ( .A(n15768), .Z(n25073) );
  OR U23455 ( .A(n15769), .B(n25073), .Z(n15770) );
  NAND U23456 ( .A(n25075), .B(n15770), .Z(n15771) );
  NANDN U23457 ( .A(n25077), .B(n15771), .Z(n15772) );
  NAND U23458 ( .A(n25079), .B(n15772), .Z(n15773) );
  NANDN U23459 ( .A(n25081), .B(n15773), .Z(n15774) );
  AND U23460 ( .A(n25083), .B(n15774), .Z(n15775) );
  OR U23461 ( .A(n25085), .B(n15775), .Z(n15776) );
  NAND U23462 ( .A(n25087), .B(n15776), .Z(n15777) );
  NANDN U23463 ( .A(n25089), .B(n15777), .Z(n15778) );
  NAND U23464 ( .A(n25091), .B(n15778), .Z(n15779) );
  NANDN U23465 ( .A(n25093), .B(n15779), .Z(n15780) );
  AND U23466 ( .A(n25095), .B(n15780), .Z(n15781) );
  OR U23467 ( .A(n25097), .B(n15781), .Z(n15782) );
  NAND U23468 ( .A(n25099), .B(n15782), .Z(n15783) );
  NANDN U23469 ( .A(n25101), .B(n15783), .Z(n15784) );
  NAND U23470 ( .A(n25103), .B(n15784), .Z(n15785) );
  NANDN U23471 ( .A(n25105), .B(n15785), .Z(n15786) );
  AND U23472 ( .A(n25107), .B(n15786), .Z(n15787) );
  OR U23473 ( .A(n25109), .B(n15787), .Z(n15788) );
  NAND U23474 ( .A(n25111), .B(n15788), .Z(n15789) );
  NANDN U23475 ( .A(n25113), .B(n15789), .Z(n15790) );
  NAND U23476 ( .A(n25115), .B(n15790), .Z(n15791) );
  NANDN U23477 ( .A(n25117), .B(n15791), .Z(n15792) );
  AND U23478 ( .A(n25119), .B(n15792), .Z(n15793) );
  OR U23479 ( .A(n25121), .B(n15793), .Z(n15794) );
  NAND U23480 ( .A(n25123), .B(n15794), .Z(n15795) );
  NANDN U23481 ( .A(n25125), .B(n15795), .Z(n15796) );
  NAND U23482 ( .A(n25127), .B(n15796), .Z(n15797) );
  NANDN U23483 ( .A(n25129), .B(n15797), .Z(n15798) );
  AND U23484 ( .A(n25131), .B(n15798), .Z(n15799) );
  OR U23485 ( .A(n25133), .B(n15799), .Z(n15800) );
  NAND U23486 ( .A(n25135), .B(n15800), .Z(n15801) );
  NANDN U23487 ( .A(n25137), .B(n15801), .Z(n15802) );
  NAND U23488 ( .A(n25139), .B(n15802), .Z(n15803) );
  NANDN U23489 ( .A(n25141), .B(n15803), .Z(n15804) );
  AND U23490 ( .A(n25143), .B(n15804), .Z(n15805) );
  OR U23491 ( .A(n25145), .B(n15805), .Z(n15806) );
  NAND U23492 ( .A(n25147), .B(n15806), .Z(n15807) );
  NANDN U23493 ( .A(n25149), .B(n15807), .Z(n15808) );
  NAND U23494 ( .A(n25151), .B(n15808), .Z(n15809) );
  NANDN U23495 ( .A(n25153), .B(n15809), .Z(n15810) );
  AND U23496 ( .A(n25155), .B(n15810), .Z(n15811) );
  OR U23497 ( .A(n25157), .B(n15811), .Z(n15812) );
  NAND U23498 ( .A(n25159), .B(n15812), .Z(n15813) );
  NANDN U23499 ( .A(n25161), .B(n15813), .Z(n15814) );
  NAND U23500 ( .A(n25163), .B(n15814), .Z(n15815) );
  NANDN U23501 ( .A(n25165), .B(n15815), .Z(n15816) );
  AND U23502 ( .A(n25167), .B(n15816), .Z(n15817) );
  OR U23503 ( .A(n25169), .B(n15817), .Z(n15818) );
  NAND U23504 ( .A(n25171), .B(n15818), .Z(n15819) );
  NANDN U23505 ( .A(n25173), .B(n15819), .Z(n15820) );
  NAND U23506 ( .A(n25175), .B(n15820), .Z(n15821) );
  NANDN U23507 ( .A(n25177), .B(n15821), .Z(n15822) );
  AND U23508 ( .A(n25179), .B(n15822), .Z(n15823) );
  OR U23509 ( .A(n25181), .B(n15823), .Z(n15824) );
  NAND U23510 ( .A(n25183), .B(n15824), .Z(n15825) );
  NANDN U23511 ( .A(n25185), .B(n15825), .Z(n15826) );
  NAND U23512 ( .A(n25187), .B(n15826), .Z(n15827) );
  NANDN U23513 ( .A(n25189), .B(n15827), .Z(n15828) );
  AND U23514 ( .A(n25191), .B(n15828), .Z(n15829) );
  OR U23515 ( .A(n25193), .B(n15829), .Z(n15830) );
  NAND U23516 ( .A(n25195), .B(n15830), .Z(n15831) );
  NANDN U23517 ( .A(n25197), .B(n15831), .Z(n15832) );
  NAND U23518 ( .A(n25199), .B(n15832), .Z(n15833) );
  NANDN U23519 ( .A(n25201), .B(n15833), .Z(n15834) );
  AND U23520 ( .A(n25203), .B(n15834), .Z(n15835) );
  OR U23521 ( .A(n25205), .B(n15835), .Z(n15836) );
  NAND U23522 ( .A(n25207), .B(n15836), .Z(n15837) );
  NAND U23523 ( .A(n25209), .B(n15837), .Z(n15838) );
  NAND U23524 ( .A(n25211), .B(n15838), .Z(n15839) );
  NANDN U23525 ( .A(n25213), .B(n15839), .Z(n15840) );
  AND U23526 ( .A(n25215), .B(n15840), .Z(n15841) );
  OR U23527 ( .A(n25217), .B(n15841), .Z(n15842) );
  NAND U23528 ( .A(n25219), .B(n15842), .Z(n15843) );
  NANDN U23529 ( .A(n25221), .B(n15843), .Z(n15844) );
  NAND U23530 ( .A(n25223), .B(n15844), .Z(n15845) );
  NANDN U23531 ( .A(n25225), .B(n15845), .Z(n15846) );
  AND U23532 ( .A(n25227), .B(n15846), .Z(n15847) );
  OR U23533 ( .A(n25229), .B(n15847), .Z(n15848) );
  NAND U23534 ( .A(n25231), .B(n15848), .Z(n15849) );
  NANDN U23535 ( .A(n25233), .B(n15849), .Z(n15852) );
  AND U23536 ( .A(n15851), .B(n15850), .Z(n25234) );
  NAND U23537 ( .A(n15852), .B(n25234), .Z(n15853) );
  AND U23538 ( .A(n15854), .B(n15853), .Z(n15855) );
  NAND U23539 ( .A(n15855), .B(n25236), .Z(n15856) );
  NAND U23540 ( .A(n25237), .B(n15856), .Z(n15857) );
  NANDN U23541 ( .A(n25238), .B(n15857), .Z(n15858) );
  AND U23542 ( .A(n25239), .B(n15858), .Z(n15859) );
  OR U23543 ( .A(n25240), .B(n15859), .Z(n15860) );
  NAND U23544 ( .A(n25241), .B(n15860), .Z(n15861) );
  NANDN U23545 ( .A(n25242), .B(n15861), .Z(n15862) );
  NAND U23546 ( .A(n25243), .B(n15862), .Z(n15863) );
  NANDN U23547 ( .A(n25244), .B(n15863), .Z(n15864) );
  AND U23548 ( .A(n25245), .B(n15864), .Z(n15865) );
  OR U23549 ( .A(n25246), .B(n15865), .Z(n15866) );
  NAND U23550 ( .A(n25247), .B(n15866), .Z(n15867) );
  NANDN U23551 ( .A(n25248), .B(n15867), .Z(n15868) );
  NAND U23552 ( .A(n25249), .B(n15868), .Z(n15869) );
  NANDN U23553 ( .A(n25250), .B(n15869), .Z(n15870) );
  AND U23554 ( .A(n25251), .B(n15870), .Z(n15871) );
  OR U23555 ( .A(n25253), .B(n15871), .Z(n15872) );
  NAND U23556 ( .A(n25255), .B(n15872), .Z(n15873) );
  NANDN U23557 ( .A(n25257), .B(n15873), .Z(n15874) );
  NAND U23558 ( .A(n25259), .B(n15874), .Z(n15875) );
  NANDN U23559 ( .A(n25261), .B(n15875), .Z(n15876) );
  AND U23560 ( .A(n25263), .B(n15876), .Z(n15877) );
  OR U23561 ( .A(n25265), .B(n15877), .Z(n15878) );
  NAND U23562 ( .A(n25267), .B(n15878), .Z(n15879) );
  NANDN U23563 ( .A(n25269), .B(n15879), .Z(n15880) );
  NAND U23564 ( .A(n25271), .B(n15880), .Z(n15881) );
  NANDN U23565 ( .A(n25273), .B(n15881), .Z(n15882) );
  AND U23566 ( .A(n25275), .B(n15882), .Z(n15883) );
  OR U23567 ( .A(n25277), .B(n15883), .Z(n15884) );
  NAND U23568 ( .A(n25279), .B(n15884), .Z(n15885) );
  NANDN U23569 ( .A(n25281), .B(n15885), .Z(n15886) );
  NAND U23570 ( .A(n25283), .B(n15886), .Z(n15887) );
  NANDN U23571 ( .A(n25285), .B(n15887), .Z(n15888) );
  AND U23572 ( .A(n25287), .B(n15888), .Z(n15889) );
  OR U23573 ( .A(n25289), .B(n15889), .Z(n15890) );
  NAND U23574 ( .A(n25291), .B(n15890), .Z(n15891) );
  NANDN U23575 ( .A(n25293), .B(n15891), .Z(n15892) );
  NAND U23576 ( .A(n25295), .B(n15892), .Z(n15893) );
  NANDN U23577 ( .A(n25297), .B(n15893), .Z(n15894) );
  AND U23578 ( .A(n25299), .B(n15894), .Z(n15895) );
  OR U23579 ( .A(n25301), .B(n15895), .Z(n15896) );
  NAND U23580 ( .A(n25303), .B(n15896), .Z(n15897) );
  NANDN U23581 ( .A(n25305), .B(n15897), .Z(n15898) );
  NAND U23582 ( .A(n25307), .B(n15898), .Z(n15899) );
  NANDN U23583 ( .A(n25309), .B(n15899), .Z(n15900) );
  AND U23584 ( .A(n25311), .B(n15900), .Z(n15901) );
  OR U23585 ( .A(n25313), .B(n15901), .Z(n15902) );
  NAND U23586 ( .A(n25315), .B(n15902), .Z(n15903) );
  NANDN U23587 ( .A(n25317), .B(n15903), .Z(n15904) );
  NAND U23588 ( .A(n25319), .B(n15904), .Z(n15905) );
  NANDN U23589 ( .A(n25321), .B(n15905), .Z(n15906) );
  AND U23590 ( .A(n25323), .B(n15906), .Z(n15907) );
  OR U23591 ( .A(n25325), .B(n15907), .Z(n15908) );
  NAND U23592 ( .A(n25327), .B(n15908), .Z(n15909) );
  NANDN U23593 ( .A(n25329), .B(n15909), .Z(n15910) );
  NAND U23594 ( .A(n25331), .B(n15910), .Z(n15911) );
  NANDN U23595 ( .A(n25333), .B(n15911), .Z(n15912) );
  AND U23596 ( .A(n25335), .B(n15912), .Z(n15913) );
  OR U23597 ( .A(n25337), .B(n15913), .Z(n15914) );
  NAND U23598 ( .A(n25339), .B(n15914), .Z(n15915) );
  NANDN U23599 ( .A(n25341), .B(n15915), .Z(n15916) );
  NAND U23600 ( .A(n25343), .B(n15916), .Z(n15917) );
  NANDN U23601 ( .A(n25345), .B(n15917), .Z(n15918) );
  AND U23602 ( .A(n25347), .B(n15918), .Z(n15919) );
  OR U23603 ( .A(n25349), .B(n15919), .Z(n15920) );
  NAND U23604 ( .A(n25351), .B(n15920), .Z(n15921) );
  NANDN U23605 ( .A(n25353), .B(n15921), .Z(n15922) );
  NAND U23606 ( .A(n25355), .B(n15922), .Z(n15923) );
  NANDN U23607 ( .A(n25357), .B(n15923), .Z(n15924) );
  AND U23608 ( .A(n25359), .B(n15924), .Z(n15925) );
  OR U23609 ( .A(n25361), .B(n15925), .Z(n15926) );
  NAND U23610 ( .A(n25363), .B(n15926), .Z(n15927) );
  NANDN U23611 ( .A(n25365), .B(n15927), .Z(n15928) );
  NAND U23612 ( .A(n25367), .B(n15928), .Z(n15929) );
  NANDN U23613 ( .A(n25369), .B(n15929), .Z(n15930) );
  AND U23614 ( .A(n25371), .B(n15930), .Z(n15931) );
  OR U23615 ( .A(n25373), .B(n15931), .Z(n15932) );
  NAND U23616 ( .A(n25375), .B(n15932), .Z(n15933) );
  NANDN U23617 ( .A(n25377), .B(n15933), .Z(n15934) );
  NAND U23618 ( .A(n25379), .B(n15934), .Z(n15935) );
  NANDN U23619 ( .A(n25381), .B(n15935), .Z(n15936) );
  AND U23620 ( .A(n25383), .B(n15936), .Z(n15937) );
  OR U23621 ( .A(n25385), .B(n15937), .Z(n15938) );
  NAND U23622 ( .A(n25387), .B(n15938), .Z(n15939) );
  NANDN U23623 ( .A(n25389), .B(n15939), .Z(n15940) );
  NAND U23624 ( .A(n25391), .B(n15940), .Z(n15941) );
  NANDN U23625 ( .A(n25393), .B(n15941), .Z(n15942) );
  AND U23626 ( .A(n25395), .B(n15942), .Z(n15943) );
  OR U23627 ( .A(n25397), .B(n15943), .Z(n15944) );
  NAND U23628 ( .A(n25399), .B(n15944), .Z(n15945) );
  NANDN U23629 ( .A(n25401), .B(n15945), .Z(n15946) );
  NAND U23630 ( .A(n25403), .B(n15946), .Z(n15947) );
  NANDN U23631 ( .A(n25405), .B(n15947), .Z(n15948) );
  AND U23632 ( .A(n25407), .B(n15948), .Z(n15949) );
  OR U23633 ( .A(n25409), .B(n15949), .Z(n15950) );
  NAND U23634 ( .A(n25411), .B(n15950), .Z(n15951) );
  NANDN U23635 ( .A(n25413), .B(n15951), .Z(n15952) );
  NAND U23636 ( .A(n25415), .B(n15952), .Z(n15953) );
  NANDN U23637 ( .A(n25417), .B(n15953), .Z(n15954) );
  AND U23638 ( .A(n25419), .B(n15954), .Z(n15955) );
  OR U23639 ( .A(n25421), .B(n15955), .Z(n15956) );
  NAND U23640 ( .A(n25423), .B(n15956), .Z(n15957) );
  NANDN U23641 ( .A(n25425), .B(n15957), .Z(n15958) );
  NAND U23642 ( .A(n25427), .B(n15958), .Z(n15959) );
  NANDN U23643 ( .A(n25429), .B(n15959), .Z(n15960) );
  AND U23644 ( .A(n25431), .B(n15960), .Z(n15961) );
  OR U23645 ( .A(n25433), .B(n15961), .Z(n15962) );
  NAND U23646 ( .A(n25435), .B(n15962), .Z(n15963) );
  NANDN U23647 ( .A(n25437), .B(n15963), .Z(n15964) );
  NAND U23648 ( .A(n25439), .B(n15964), .Z(n15965) );
  NANDN U23649 ( .A(n25441), .B(n15965), .Z(n15966) );
  AND U23650 ( .A(n25443), .B(n15966), .Z(n15967) );
  OR U23651 ( .A(n25445), .B(n15967), .Z(n15968) );
  NAND U23652 ( .A(n25447), .B(n15968), .Z(n15969) );
  NANDN U23653 ( .A(n25449), .B(n15969), .Z(n15970) );
  NAND U23654 ( .A(n25451), .B(n15970), .Z(n15971) );
  NANDN U23655 ( .A(n25453), .B(n15971), .Z(n15972) );
  AND U23656 ( .A(n25455), .B(n15972), .Z(n15973) );
  OR U23657 ( .A(n25457), .B(n15973), .Z(n15974) );
  NAND U23658 ( .A(n25459), .B(n15974), .Z(n15975) );
  NANDN U23659 ( .A(n25461), .B(n15975), .Z(n15976) );
  NAND U23660 ( .A(n25463), .B(n15976), .Z(n15977) );
  NANDN U23661 ( .A(n25465), .B(n15977), .Z(n15978) );
  AND U23662 ( .A(n25467), .B(n15978), .Z(n15979) );
  OR U23663 ( .A(n25469), .B(n15979), .Z(n15980) );
  NAND U23664 ( .A(n25471), .B(n15980), .Z(n15981) );
  NANDN U23665 ( .A(n25473), .B(n15981), .Z(n15982) );
  NAND U23666 ( .A(n25475), .B(n15982), .Z(n15983) );
  NANDN U23667 ( .A(n25477), .B(n15983), .Z(n15984) );
  AND U23668 ( .A(n25479), .B(n15984), .Z(n15985) );
  OR U23669 ( .A(n25481), .B(n15985), .Z(n15986) );
  NAND U23670 ( .A(n25483), .B(n15986), .Z(n15987) );
  NANDN U23671 ( .A(n25485), .B(n15987), .Z(n15988) );
  NAND U23672 ( .A(n25487), .B(n15988), .Z(n15989) );
  NANDN U23673 ( .A(n25489), .B(n15989), .Z(n15990) );
  AND U23674 ( .A(n25491), .B(n15990), .Z(n15991) );
  OR U23675 ( .A(n25493), .B(n15991), .Z(n15992) );
  NAND U23676 ( .A(n25495), .B(n15992), .Z(n15993) );
  NANDN U23677 ( .A(n25497), .B(n15993), .Z(n15994) );
  NAND U23678 ( .A(n25499), .B(n15994), .Z(n15995) );
  NANDN U23679 ( .A(n25501), .B(n15995), .Z(n15996) );
  AND U23680 ( .A(n25503), .B(n15996), .Z(n15997) );
  OR U23681 ( .A(n25505), .B(n15997), .Z(n15998) );
  NAND U23682 ( .A(n25507), .B(n15998), .Z(n15999) );
  NANDN U23683 ( .A(n25509), .B(n15999), .Z(n16000) );
  NAND U23684 ( .A(n25511), .B(n16000), .Z(n16001) );
  NANDN U23685 ( .A(n25513), .B(n16001), .Z(n16002) );
  AND U23686 ( .A(n25515), .B(n16002), .Z(n16003) );
  OR U23687 ( .A(n25517), .B(n16003), .Z(n16004) );
  NAND U23688 ( .A(n25519), .B(n16004), .Z(n16005) );
  NANDN U23689 ( .A(n25521), .B(n16005), .Z(n16006) );
  NAND U23690 ( .A(n25523), .B(n16006), .Z(n16007) );
  NANDN U23691 ( .A(n25525), .B(n16007), .Z(n16008) );
  AND U23692 ( .A(n25527), .B(n16008), .Z(n16009) );
  OR U23693 ( .A(n25529), .B(n16009), .Z(n16010) );
  NAND U23694 ( .A(n25531), .B(n16010), .Z(n16011) );
  NANDN U23695 ( .A(n25532), .B(n16011), .Z(n16013) );
  OR U23696 ( .A(n16013), .B(n16012), .Z(n16014) );
  NAND U23697 ( .A(n25534), .B(n16014), .Z(n16015) );
  NANDN U23698 ( .A(n25535), .B(n16015), .Z(n16016) );
  NAND U23699 ( .A(n25536), .B(n16016), .Z(n16017) );
  NANDN U23700 ( .A(n25537), .B(n16017), .Z(n16018) );
  AND U23701 ( .A(n25538), .B(n16018), .Z(n16019) );
  OR U23702 ( .A(n25539), .B(n16019), .Z(n16020) );
  NAND U23703 ( .A(n25540), .B(n16020), .Z(n16021) );
  NANDN U23704 ( .A(n25541), .B(n16021), .Z(n16022) );
  NAND U23705 ( .A(n25542), .B(n16022), .Z(n16023) );
  NANDN U23706 ( .A(n25543), .B(n16023), .Z(n16024) );
  AND U23707 ( .A(n25544), .B(n16024), .Z(n16025) );
  OR U23708 ( .A(n25545), .B(n16025), .Z(n16026) );
  NAND U23709 ( .A(n25546), .B(n16026), .Z(n16027) );
  NANDN U23710 ( .A(n25547), .B(n16027), .Z(n16028) );
  NAND U23711 ( .A(n25548), .B(n16028), .Z(n16029) );
  NANDN U23712 ( .A(n25549), .B(n16029), .Z(n16030) );
  AND U23713 ( .A(n25550), .B(n16030), .Z(n16031) );
  OR U23714 ( .A(n25552), .B(n16031), .Z(n16032) );
  NAND U23715 ( .A(n25554), .B(n16032), .Z(n16033) );
  NANDN U23716 ( .A(n25556), .B(n16033), .Z(n16034) );
  NAND U23717 ( .A(n25558), .B(n16034), .Z(n16035) );
  NANDN U23718 ( .A(n25560), .B(n16035), .Z(n16036) );
  AND U23719 ( .A(n25562), .B(n16036), .Z(n16037) );
  OR U23720 ( .A(n25564), .B(n16037), .Z(n16038) );
  NAND U23721 ( .A(n25566), .B(n16038), .Z(n16039) );
  NANDN U23722 ( .A(n25568), .B(n16039), .Z(n16040) );
  NAND U23723 ( .A(n25570), .B(n16040), .Z(n16041) );
  NANDN U23724 ( .A(n25572), .B(n16041), .Z(n16042) );
  AND U23725 ( .A(n25574), .B(n16042), .Z(n16043) );
  OR U23726 ( .A(n25576), .B(n16043), .Z(n16044) );
  NAND U23727 ( .A(n25578), .B(n16044), .Z(n16045) );
  NANDN U23728 ( .A(n25580), .B(n16045), .Z(n16046) );
  NAND U23729 ( .A(n25582), .B(n16046), .Z(n16047) );
  NANDN U23730 ( .A(n25584), .B(n16047), .Z(n16048) );
  AND U23731 ( .A(n25586), .B(n16048), .Z(n16049) );
  OR U23732 ( .A(n25588), .B(n16049), .Z(n16050) );
  NAND U23733 ( .A(n25590), .B(n16050), .Z(n16051) );
  NANDN U23734 ( .A(n25592), .B(n16051), .Z(n16052) );
  NAND U23735 ( .A(n25594), .B(n16052), .Z(n16053) );
  NANDN U23736 ( .A(n25596), .B(n16053), .Z(n16054) );
  AND U23737 ( .A(n25598), .B(n16054), .Z(n16055) );
  OR U23738 ( .A(n25600), .B(n16055), .Z(n16056) );
  NAND U23739 ( .A(n25602), .B(n16056), .Z(n16057) );
  NANDN U23740 ( .A(n25604), .B(n16057), .Z(n16058) );
  NAND U23741 ( .A(n25606), .B(n16058), .Z(n16059) );
  NANDN U23742 ( .A(n25608), .B(n16059), .Z(n16060) );
  AND U23743 ( .A(n25610), .B(n16060), .Z(n16061) );
  OR U23744 ( .A(n25612), .B(n16061), .Z(n16062) );
  NAND U23745 ( .A(n25614), .B(n16062), .Z(n16063) );
  NANDN U23746 ( .A(n25616), .B(n16063), .Z(n16064) );
  NAND U23747 ( .A(n25618), .B(n16064), .Z(n16065) );
  NANDN U23748 ( .A(n25620), .B(n16065), .Z(n16066) );
  AND U23749 ( .A(n25622), .B(n16066), .Z(n16067) );
  OR U23750 ( .A(n25624), .B(n16067), .Z(n16068) );
  NAND U23751 ( .A(n25626), .B(n16068), .Z(n16069) );
  NANDN U23752 ( .A(n25628), .B(n16069), .Z(n16070) );
  NAND U23753 ( .A(n25630), .B(n16070), .Z(n16071) );
  NANDN U23754 ( .A(n25632), .B(n16071), .Z(n16072) );
  AND U23755 ( .A(n25633), .B(n16072), .Z(n16073) );
  NOR U23756 ( .A(n16074), .B(n16073), .Z(n16075) );
  NANDN U23757 ( .A(n25634), .B(n16075), .Z(n16076) );
  AND U23758 ( .A(n25635), .B(n16076), .Z(n16077) );
  OR U23759 ( .A(n25636), .B(n16077), .Z(n16078) );
  NAND U23760 ( .A(n25637), .B(n16078), .Z(n16079) );
  NANDN U23761 ( .A(n25638), .B(n16079), .Z(n16080) );
  NAND U23762 ( .A(n25639), .B(n16080), .Z(n16081) );
  NANDN U23763 ( .A(n25640), .B(n16081), .Z(n16082) );
  AND U23764 ( .A(n25641), .B(n16082), .Z(n16083) );
  OR U23765 ( .A(n25642), .B(n16083), .Z(n16084) );
  NAND U23766 ( .A(n25643), .B(n16084), .Z(n16085) );
  NANDN U23767 ( .A(n25644), .B(n16085), .Z(n16086) );
  NAND U23768 ( .A(n25645), .B(n16086), .Z(n16088) );
  ANDN U23769 ( .B(n16088), .A(n16087), .Z(n16089) );
  NANDN U23770 ( .A(n25647), .B(n16089), .Z(n16090) );
  NAND U23771 ( .A(n25648), .B(n16090), .Z(n16091) );
  NANDN U23772 ( .A(n25650), .B(n16091), .Z(n16092) );
  AND U23773 ( .A(n25652), .B(n16092), .Z(n16093) );
  OR U23774 ( .A(n25654), .B(n16093), .Z(n16094) );
  NAND U23775 ( .A(n25656), .B(n16094), .Z(n16095) );
  NANDN U23776 ( .A(n25658), .B(n16095), .Z(n16096) );
  NAND U23777 ( .A(n25660), .B(n16096), .Z(n16097) );
  NANDN U23778 ( .A(n25662), .B(n16097), .Z(n16098) );
  AND U23779 ( .A(n25664), .B(n16098), .Z(n16099) );
  OR U23780 ( .A(n25666), .B(n16099), .Z(n16100) );
  NAND U23781 ( .A(n25668), .B(n16100), .Z(n16101) );
  NANDN U23782 ( .A(n25670), .B(n16101), .Z(n16102) );
  NAND U23783 ( .A(n25672), .B(n16102), .Z(n16103) );
  NANDN U23784 ( .A(n25674), .B(n16103), .Z(n16104) );
  AND U23785 ( .A(n25676), .B(n16104), .Z(n16105) );
  OR U23786 ( .A(n25678), .B(n16105), .Z(n16106) );
  NAND U23787 ( .A(n25680), .B(n16106), .Z(n16107) );
  NANDN U23788 ( .A(n25682), .B(n16107), .Z(n16108) );
  NAND U23789 ( .A(n25684), .B(n16108), .Z(n16109) );
  NANDN U23790 ( .A(n25686), .B(n16109), .Z(n16110) );
  AND U23791 ( .A(n25688), .B(n16110), .Z(n16111) );
  OR U23792 ( .A(n25690), .B(n16111), .Z(n16112) );
  NAND U23793 ( .A(n25692), .B(n16112), .Z(n16113) );
  NANDN U23794 ( .A(n25694), .B(n16113), .Z(n16114) );
  NAND U23795 ( .A(n25696), .B(n16114), .Z(n16115) );
  NANDN U23796 ( .A(n25698), .B(n16115), .Z(n16116) );
  AND U23797 ( .A(n25700), .B(n16116), .Z(n16117) );
  OR U23798 ( .A(n25702), .B(n16117), .Z(n16118) );
  NAND U23799 ( .A(n25704), .B(n16118), .Z(n16119) );
  NANDN U23800 ( .A(n25706), .B(n16119), .Z(n16120) );
  NAND U23801 ( .A(n25708), .B(n16120), .Z(n16121) );
  NANDN U23802 ( .A(n25710), .B(n16121), .Z(n16122) );
  AND U23803 ( .A(n25712), .B(n16122), .Z(n16123) );
  OR U23804 ( .A(n25714), .B(n16123), .Z(n16124) );
  NAND U23805 ( .A(n25716), .B(n16124), .Z(n16125) );
  NANDN U23806 ( .A(n25718), .B(n16125), .Z(n16126) );
  NAND U23807 ( .A(n25720), .B(n16126), .Z(n16127) );
  NANDN U23808 ( .A(n25722), .B(n16127), .Z(n16128) );
  AND U23809 ( .A(n25724), .B(n16128), .Z(n16129) );
  OR U23810 ( .A(n25726), .B(n16129), .Z(n16130) );
  NAND U23811 ( .A(n25728), .B(n16130), .Z(n16131) );
  NANDN U23812 ( .A(n25730), .B(n16131), .Z(n16132) );
  NAND U23813 ( .A(n25732), .B(n16132), .Z(n16133) );
  NANDN U23814 ( .A(n25734), .B(n16133), .Z(n16134) );
  AND U23815 ( .A(n25736), .B(n16134), .Z(n16135) );
  OR U23816 ( .A(n25738), .B(n16135), .Z(n16136) );
  NAND U23817 ( .A(n25740), .B(n16136), .Z(n16137) );
  NANDN U23818 ( .A(n25742), .B(n16137), .Z(n16138) );
  NAND U23819 ( .A(n25744), .B(n16138), .Z(n16139) );
  NANDN U23820 ( .A(n25746), .B(n16139), .Z(n16140) );
  AND U23821 ( .A(n25748), .B(n16140), .Z(n16141) );
  OR U23822 ( .A(n25750), .B(n16141), .Z(n16142) );
  NAND U23823 ( .A(n25752), .B(n16142), .Z(n16143) );
  NANDN U23824 ( .A(n25754), .B(n16143), .Z(n16144) );
  NAND U23825 ( .A(n25756), .B(n16144), .Z(n16145) );
  NANDN U23826 ( .A(n25758), .B(n16145), .Z(n16146) );
  AND U23827 ( .A(n25760), .B(n16146), .Z(n16147) );
  OR U23828 ( .A(n25762), .B(n16147), .Z(n16148) );
  NAND U23829 ( .A(n25764), .B(n16148), .Z(n16149) );
  NANDN U23830 ( .A(n25766), .B(n16149), .Z(n16150) );
  NAND U23831 ( .A(n25768), .B(n16150), .Z(n16151) );
  NANDN U23832 ( .A(n25770), .B(n16151), .Z(n16152) );
  AND U23833 ( .A(n25772), .B(n16152), .Z(n16153) );
  OR U23834 ( .A(n25774), .B(n16153), .Z(n16154) );
  NAND U23835 ( .A(n25776), .B(n16154), .Z(n16155) );
  NANDN U23836 ( .A(n25778), .B(n16155), .Z(n16156) );
  NAND U23837 ( .A(n25780), .B(n16156), .Z(n16157) );
  NANDN U23838 ( .A(n25782), .B(n16157), .Z(n16158) );
  AND U23839 ( .A(n25784), .B(n16158), .Z(n16159) );
  OR U23840 ( .A(n25786), .B(n16159), .Z(n16160) );
  NAND U23841 ( .A(n25788), .B(n16160), .Z(n16161) );
  NANDN U23842 ( .A(n25790), .B(n16161), .Z(n16162) );
  NAND U23843 ( .A(n25792), .B(n16162), .Z(n16163) );
  NANDN U23844 ( .A(n25794), .B(n16163), .Z(n16164) );
  AND U23845 ( .A(n25796), .B(n16164), .Z(n16165) );
  OR U23846 ( .A(n25798), .B(n16165), .Z(n16166) );
  NAND U23847 ( .A(n25800), .B(n16166), .Z(n16167) );
  NANDN U23848 ( .A(n25802), .B(n16167), .Z(n16168) );
  NAND U23849 ( .A(n25804), .B(n16168), .Z(n16169) );
  NANDN U23850 ( .A(n25806), .B(n16169), .Z(n16170) );
  AND U23851 ( .A(n25808), .B(n16170), .Z(n16171) );
  OR U23852 ( .A(n25810), .B(n16171), .Z(n16172) );
  NAND U23853 ( .A(n25812), .B(n16172), .Z(n16173) );
  NANDN U23854 ( .A(n25814), .B(n16173), .Z(n16174) );
  NAND U23855 ( .A(n25816), .B(n16174), .Z(n16175) );
  NANDN U23856 ( .A(n25818), .B(n16175), .Z(n16176) );
  AND U23857 ( .A(n25820), .B(n16176), .Z(n16177) );
  OR U23858 ( .A(n25822), .B(n16177), .Z(n16178) );
  NAND U23859 ( .A(n25824), .B(n16178), .Z(n16179) );
  NANDN U23860 ( .A(n25826), .B(n16179), .Z(n16180) );
  NAND U23861 ( .A(n25828), .B(n16180), .Z(n16181) );
  NANDN U23862 ( .A(n25830), .B(n16181), .Z(n16182) );
  AND U23863 ( .A(n25832), .B(n16182), .Z(n16183) );
  OR U23864 ( .A(n25834), .B(n16183), .Z(n16184) );
  NAND U23865 ( .A(n25836), .B(n16184), .Z(n16185) );
  NANDN U23866 ( .A(n25838), .B(n16185), .Z(n16186) );
  NAND U23867 ( .A(n25840), .B(n16186), .Z(n16187) );
  NANDN U23868 ( .A(n25842), .B(n16187), .Z(n16188) );
  AND U23869 ( .A(n25844), .B(n16188), .Z(n16189) );
  OR U23870 ( .A(n25846), .B(n16189), .Z(n16190) );
  NAND U23871 ( .A(n25848), .B(n16190), .Z(n16191) );
  NANDN U23872 ( .A(n25850), .B(n16191), .Z(n16192) );
  NAND U23873 ( .A(n25851), .B(n16192), .Z(n16193) );
  NANDN U23874 ( .A(n25852), .B(n16193), .Z(n16194) );
  AND U23875 ( .A(n25853), .B(n16194), .Z(n16196) );
  NANDN U23876 ( .A(n16196), .B(n25854), .Z(n16197) );
  NANDN U23877 ( .A(n24537), .B(n16197), .Z(n16198) );
  AND U23878 ( .A(n25855), .B(n16198), .Z(n16199) );
  NOR U23879 ( .A(n16199), .B(n25856), .Z(n16200) );
  NANDN U23880 ( .A(n16201), .B(n16200), .Z(n16202) );
  AND U23881 ( .A(n16203), .B(n16202), .Z(n16204) );
  NAND U23882 ( .A(n16204), .B(n25857), .Z(n16206) );
  ANDN U23883 ( .B(n16206), .A(n16205), .Z(n16207) );
  NANDN U23884 ( .A(n16208), .B(n16207), .Z(n16211) );
  AND U23885 ( .A(n16209), .B(n24535), .Z(n16210) );
  NAND U23886 ( .A(n16211), .B(n16210), .Z(n16212) );
  NAND U23887 ( .A(n25860), .B(n16212), .Z(n16213) );
  NAND U23888 ( .A(n25861), .B(n16213), .Z(n16214) );
  NAND U23889 ( .A(n25862), .B(n16214), .Z(n16217) );
  AND U23890 ( .A(n16216), .B(n16215), .Z(n24534) );
  AND U23891 ( .A(n16217), .B(n24534), .Z(n16220) );
  NANDN U23892 ( .A(n16220), .B(n25864), .Z(n16221) );
  NAND U23893 ( .A(n24533), .B(n16221), .Z(n16222) );
  NAND U23894 ( .A(n25865), .B(n16222), .Z(n16223) );
  NAND U23895 ( .A(n25866), .B(n16223), .Z(n16224) );
  NAND U23896 ( .A(n25867), .B(n16224), .Z(n16227) );
  XNOR U23897 ( .A(y[702]), .B(x[702]), .Z(n16225) );
  AND U23898 ( .A(n16226), .B(n16225), .Z(n24532) );
  AND U23899 ( .A(n16227), .B(n24532), .Z(n16231) );
  IV U23900 ( .A(n16228), .Z(n16230) );
  ANDN U23901 ( .B(n16230), .A(n16229), .Z(n25868) );
  NANDN U23902 ( .A(n16231), .B(n25868), .Z(n16232) );
  NAND U23903 ( .A(n24531), .B(n16232), .Z(n16233) );
  NAND U23904 ( .A(n25869), .B(n16233), .Z(n16234) );
  NAND U23905 ( .A(n25870), .B(n16234), .Z(n16235) );
  NANDN U23906 ( .A(n24530), .B(n16235), .Z(n16236) );
  AND U23907 ( .A(n25871), .B(n16236), .Z(n16239) );
  NANDN U23908 ( .A(n16239), .B(n25872), .Z(n16240) );
  NAND U23909 ( .A(n25874), .B(n16240), .Z(n16241) );
  NAND U23910 ( .A(n25875), .B(n16241), .Z(n16242) );
  NAND U23911 ( .A(n25876), .B(n16242), .Z(n16243) );
  NAND U23912 ( .A(n25877), .B(n16243), .Z(n16246) );
  XNOR U23913 ( .A(y[714]), .B(x[714]), .Z(n16244) );
  AND U23914 ( .A(n16245), .B(n16244), .Z(n24529) );
  AND U23915 ( .A(n16246), .B(n24529), .Z(n16249) );
  NANDN U23916 ( .A(n16249), .B(n25878), .Z(n16250) );
  NAND U23917 ( .A(n25879), .B(n16250), .Z(n16251) );
  NAND U23918 ( .A(n25880), .B(n16251), .Z(n16252) );
  NAND U23919 ( .A(n25881), .B(n16252), .Z(n16253) );
  NAND U23920 ( .A(n25882), .B(n16253), .Z(n16256) );
  AND U23921 ( .A(n16255), .B(n16254), .Z(n24528) );
  AND U23922 ( .A(n16256), .B(n24528), .Z(n16260) );
  IV U23923 ( .A(n16257), .Z(n16259) );
  ANDN U23924 ( .B(n16259), .A(n16258), .Z(n25883) );
  NANDN U23925 ( .A(n16260), .B(n25883), .Z(n16261) );
  NAND U23926 ( .A(n24527), .B(n16261), .Z(n16262) );
  NANDN U23927 ( .A(n25884), .B(n16262), .Z(n16263) );
  NAND U23928 ( .A(n25885), .B(n16263), .Z(n16264) );
  NAND U23929 ( .A(n25887), .B(n16264), .Z(n16265) );
  AND U23930 ( .A(n25888), .B(n16265), .Z(n16268) );
  ANDN U23931 ( .B(n16267), .A(n16266), .Z(n25889) );
  NANDN U23932 ( .A(n16268), .B(n25889), .Z(n16269) );
  NAND U23933 ( .A(n24526), .B(n16269), .Z(n16270) );
  NAND U23934 ( .A(n25890), .B(n16270), .Z(n16271) );
  NAND U23935 ( .A(n25891), .B(n16271), .Z(n16272) );
  NAND U23936 ( .A(n25892), .B(n16272), .Z(n16275) );
  XNOR U23937 ( .A(x[732]), .B(y[732]), .Z(n16273) );
  AND U23938 ( .A(n16274), .B(n16273), .Z(n24525) );
  AND U23939 ( .A(n16275), .B(n24525), .Z(n16278) );
  NANDN U23940 ( .A(n16278), .B(n25893), .Z(n16279) );
  NAND U23941 ( .A(n24524), .B(n16279), .Z(n16280) );
  NAND U23942 ( .A(n25894), .B(n16280), .Z(n16281) );
  NAND U23943 ( .A(n25895), .B(n16281), .Z(n16282) );
  NANDN U23944 ( .A(n24523), .B(n16282), .Z(n16283) );
  AND U23945 ( .A(n25896), .B(n16283), .Z(n16286) );
  NAND U23946 ( .A(n16285), .B(n16284), .Z(n24522) );
  OR U23947 ( .A(n16286), .B(n24522), .Z(n16287) );
  NAND U23948 ( .A(n25898), .B(n16287), .Z(n16288) );
  NANDN U23949 ( .A(n25899), .B(n16288), .Z(n16289) );
  NAND U23950 ( .A(n25900), .B(n16289), .Z(n16290) );
  NAND U23951 ( .A(n25901), .B(n16290), .Z(n16291) );
  AND U23952 ( .A(n25902), .B(n16291), .Z(n16294) );
  ANDN U23953 ( .B(n16293), .A(n16292), .Z(n25903) );
  NANDN U23954 ( .A(n16294), .B(n25903), .Z(n16295) );
  NAND U23955 ( .A(n24521), .B(n16295), .Z(n16296) );
  NAND U23956 ( .A(n25904), .B(n16296), .Z(n16297) );
  NAND U23957 ( .A(n25905), .B(n16297), .Z(n16298) );
  NAND U23958 ( .A(n25906), .B(n16298), .Z(n16301) );
  XNOR U23959 ( .A(y[750]), .B(x[750]), .Z(n16299) );
  AND U23960 ( .A(n16300), .B(n16299), .Z(n24520) );
  AND U23961 ( .A(n16301), .B(n24520), .Z(n16304) );
  NANDN U23962 ( .A(n16304), .B(n25907), .Z(n16305) );
  NAND U23963 ( .A(n24519), .B(n16305), .Z(n16306) );
  NAND U23964 ( .A(n25908), .B(n16306), .Z(n16307) );
  NAND U23965 ( .A(n25909), .B(n16307), .Z(n16308) );
  NAND U23966 ( .A(n25912), .B(n16308), .Z(n16309) );
  AND U23967 ( .A(n25913), .B(n16309), .Z(n16312) );
  NAND U23968 ( .A(n16311), .B(n16310), .Z(n24518) );
  OR U23969 ( .A(n16312), .B(n24518), .Z(n16313) );
  NAND U23970 ( .A(n25914), .B(n16313), .Z(n16314) );
  NANDN U23971 ( .A(n25915), .B(n16314), .Z(n16315) );
  NAND U23972 ( .A(n25916), .B(n16315), .Z(n16316) );
  NAND U23973 ( .A(n25917), .B(n16316), .Z(n16319) );
  AND U23974 ( .A(n16318), .B(n16317), .Z(n24517) );
  AND U23975 ( .A(n16319), .B(n24517), .Z(n16323) );
  IV U23976 ( .A(n16320), .Z(n16322) );
  ANDN U23977 ( .B(n16322), .A(n16321), .Z(n25918) );
  NANDN U23978 ( .A(n16323), .B(n25918), .Z(n16324) );
  NAND U23979 ( .A(n25919), .B(n16324), .Z(n16325) );
  NAND U23980 ( .A(n25920), .B(n16325), .Z(n16326) );
  NAND U23981 ( .A(n25921), .B(n16326), .Z(n16327) );
  NANDN U23982 ( .A(n24516), .B(n16327), .Z(n16328) );
  AND U23983 ( .A(n25922), .B(n16328), .Z(n16331) );
  NANDN U23984 ( .A(n16331), .B(n25923), .Z(n16332) );
  NAND U23985 ( .A(n24515), .B(n16332), .Z(n16333) );
  NAND U23986 ( .A(n25926), .B(n16333), .Z(n16334) );
  NAND U23987 ( .A(n25927), .B(n16334), .Z(n16335) );
  NAND U23988 ( .A(n25928), .B(n16335), .Z(n16336) );
  AND U23989 ( .A(n25929), .B(n16336), .Z(n16337) );
  OR U23990 ( .A(n16337), .B(n24514), .Z(n16338) );
  NAND U23991 ( .A(n24513), .B(n16338), .Z(n16339) );
  NANDN U23992 ( .A(n25930), .B(n16339), .Z(n16340) );
  NAND U23993 ( .A(n25931), .B(n16340), .Z(n16341) );
  NANDN U23994 ( .A(n24512), .B(n16341), .Z(n16342) );
  AND U23995 ( .A(n16342), .B(n24511), .Z(n16343) );
  OR U23996 ( .A(n16343), .B(n24510), .Z(n16344) );
  NAND U23997 ( .A(n25933), .B(n16344), .Z(n16345) );
  NANDN U23998 ( .A(n16346), .B(n16345), .Z(n16347) );
  NAND U23999 ( .A(n25935), .B(n16347), .Z(n16348) );
  NAND U24000 ( .A(n25936), .B(n16348), .Z(n16349) );
  NANDN U24001 ( .A(n25937), .B(n16349), .Z(n16350) );
  NAND U24002 ( .A(n25938), .B(n16350), .Z(n16351) );
  NANDN U24003 ( .A(n25939), .B(n16351), .Z(n16353) );
  IV U24004 ( .A(n16352), .Z(n25940) );
  AND U24005 ( .A(n16353), .B(n25940), .Z(n16355) );
  IV U24006 ( .A(n16354), .Z(n25941) );
  OR U24007 ( .A(n16355), .B(n25941), .Z(n16356) );
  NAND U24008 ( .A(n25942), .B(n16356), .Z(n16357) );
  NANDN U24009 ( .A(n25943), .B(n16357), .Z(n16358) );
  NAND U24010 ( .A(n25944), .B(n16358), .Z(n16359) );
  NANDN U24011 ( .A(n25945), .B(n16359), .Z(n16360) );
  AND U24012 ( .A(n25946), .B(n16360), .Z(n16361) );
  OR U24013 ( .A(n25947), .B(n16361), .Z(n16362) );
  NAND U24014 ( .A(n25948), .B(n16362), .Z(n16363) );
  NANDN U24015 ( .A(n25949), .B(n16363), .Z(n16364) );
  NAND U24016 ( .A(n25950), .B(n16364), .Z(n16365) );
  NANDN U24017 ( .A(n25951), .B(n16365), .Z(n16366) );
  AND U24018 ( .A(n25953), .B(n16366), .Z(n16367) );
  OR U24019 ( .A(n25955), .B(n16367), .Z(n16368) );
  NAND U24020 ( .A(n25957), .B(n16368), .Z(n16369) );
  NANDN U24021 ( .A(n25959), .B(n16369), .Z(n16370) );
  NAND U24022 ( .A(n25961), .B(n16370), .Z(n16371) );
  NANDN U24023 ( .A(n25963), .B(n16371), .Z(n16372) );
  AND U24024 ( .A(n25965), .B(n16372), .Z(n16373) );
  OR U24025 ( .A(n25967), .B(n16373), .Z(n16374) );
  NAND U24026 ( .A(n25969), .B(n16374), .Z(n16375) );
  NANDN U24027 ( .A(n25971), .B(n16375), .Z(n16376) );
  NAND U24028 ( .A(n25973), .B(n16376), .Z(n16377) );
  NANDN U24029 ( .A(n25975), .B(n16377), .Z(n16378) );
  AND U24030 ( .A(n25977), .B(n16378), .Z(n16379) );
  OR U24031 ( .A(n25979), .B(n16379), .Z(n16380) );
  NAND U24032 ( .A(n25981), .B(n16380), .Z(n16381) );
  NANDN U24033 ( .A(n25983), .B(n16381), .Z(n16382) );
  NAND U24034 ( .A(n25985), .B(n16382), .Z(n16383) );
  NANDN U24035 ( .A(n25987), .B(n16383), .Z(n16384) );
  AND U24036 ( .A(n25989), .B(n16384), .Z(n16385) );
  OR U24037 ( .A(n25990), .B(n16385), .Z(n16386) );
  NAND U24038 ( .A(n25993), .B(n16386), .Z(n16387) );
  NANDN U24039 ( .A(n25995), .B(n16387), .Z(n16388) );
  NAND U24040 ( .A(n25997), .B(n16388), .Z(n16389) );
  ANDN U24041 ( .B(n16389), .A(n25999), .Z(n16390) );
  NANDN U24042 ( .A(n16391), .B(n16390), .Z(n16392) );
  NAND U24043 ( .A(n16393), .B(n16392), .Z(n16395) );
  IV U24044 ( .A(n16394), .Z(n26006) );
  ANDN U24045 ( .B(n16395), .A(n26006), .Z(n16396) );
  NANDN U24046 ( .A(n16397), .B(n16396), .Z(n16400) );
  AND U24047 ( .A(n26009), .B(n16398), .Z(n16399) );
  NAND U24048 ( .A(n16400), .B(n16399), .Z(n16401) );
  NAND U24049 ( .A(n26011), .B(n16401), .Z(n16404) );
  NANDN U24050 ( .A(y[828]), .B(n16404), .Z(n16403) );
  ANDN U24051 ( .B(n16403), .A(n16402), .Z(n16407) );
  XNOR U24052 ( .A(n16404), .B(y[828]), .Z(n16405) );
  NAND U24053 ( .A(n16405), .B(x[828]), .Z(n16406) );
  NAND U24054 ( .A(n16407), .B(n16406), .Z(n16408) );
  NAND U24055 ( .A(n26017), .B(n16408), .Z(n16409) );
  NANDN U24056 ( .A(n16410), .B(n16409), .Z(n16411) );
  AND U24057 ( .A(n26021), .B(n16411), .Z(n16412) );
  NOR U24058 ( .A(n26023), .B(n16412), .Z(n16413) );
  NANDN U24059 ( .A(n16414), .B(n16413), .Z(n16415) );
  AND U24060 ( .A(n26025), .B(n16415), .Z(n16416) );
  OR U24061 ( .A(n26027), .B(n16416), .Z(n16417) );
  NAND U24062 ( .A(n26029), .B(n16417), .Z(n16418) );
  NANDN U24063 ( .A(n26031), .B(n16418), .Z(n16419) );
  NAND U24064 ( .A(n26033), .B(n16419), .Z(n16420) );
  NANDN U24065 ( .A(n26034), .B(n16420), .Z(n16422) );
  IV U24066 ( .A(n16421), .Z(n26035) );
  AND U24067 ( .A(n16422), .B(n26035), .Z(n16423) );
  NOR U24068 ( .A(n26036), .B(n16423), .Z(n16424) );
  NANDN U24069 ( .A(n16425), .B(n16424), .Z(n16427) );
  IV U24070 ( .A(n16426), .Z(n26037) );
  AND U24071 ( .A(n16427), .B(n26037), .Z(n16428) );
  NAND U24072 ( .A(n26039), .B(n16428), .Z(n16429) );
  AND U24073 ( .A(n16429), .B(n26040), .Z(n16430) );
  NANDN U24074 ( .A(n16431), .B(n16430), .Z(n16432) );
  NAND U24075 ( .A(n26041), .B(n16432), .Z(n16433) );
  ANDN U24076 ( .B(n16433), .A(n26042), .Z(n16434) );
  NANDN U24077 ( .A(n16435), .B(n16434), .Z(n16436) );
  NAND U24078 ( .A(n16437), .B(n16436), .Z(n16438) );
  AND U24079 ( .A(n26044), .B(n16438), .Z(n16439) );
  NANDN U24080 ( .A(n16440), .B(n16439), .Z(n16441) );
  NAND U24081 ( .A(n26045), .B(n16441), .Z(n16442) );
  NANDN U24082 ( .A(n26046), .B(n16442), .Z(n16443) );
  AND U24083 ( .A(n16444), .B(n16443), .Z(n16445) );
  OR U24084 ( .A(n26049), .B(n16445), .Z(n16446) );
  NAND U24085 ( .A(n16447), .B(n16446), .Z(n16448) );
  NAND U24086 ( .A(n26051), .B(n16448), .Z(n16449) );
  NANDN U24087 ( .A(n26052), .B(n16449), .Z(n16450) );
  AND U24088 ( .A(n26053), .B(n16450), .Z(n16451) );
  OR U24089 ( .A(n26054), .B(n16451), .Z(n16452) );
  AND U24090 ( .A(n16453), .B(n16452), .Z(n16455) );
  NOR U24091 ( .A(n16455), .B(n16454), .Z(n16456) );
  NANDN U24092 ( .A(n26057), .B(n16456), .Z(n16457) );
  AND U24093 ( .A(n16458), .B(n16457), .Z(n16459) );
  NAND U24094 ( .A(n16459), .B(n26058), .Z(n16461) );
  ANDN U24095 ( .B(n16461), .A(n16460), .Z(n16462) );
  NANDN U24096 ( .A(n16463), .B(n16462), .Z(n16467) );
  AND U24097 ( .A(n16465), .B(n16464), .Z(n16466) );
  NAND U24098 ( .A(n16467), .B(n16466), .Z(n16468) );
  NANDN U24099 ( .A(n16469), .B(n16468), .Z(n16471) );
  OR U24100 ( .A(n16471), .B(n16470), .Z(n16472) );
  AND U24101 ( .A(n16473), .B(n16472), .Z(n16475) );
  NOR U24102 ( .A(n16475), .B(n16474), .Z(n16476) );
  NANDN U24103 ( .A(n16477), .B(n16476), .Z(n16478) );
  AND U24104 ( .A(n16479), .B(n16478), .Z(n16481) );
  NAND U24105 ( .A(n16481), .B(n16480), .Z(n16483) );
  ANDN U24106 ( .B(n16483), .A(n16482), .Z(n16484) );
  NANDN U24107 ( .A(n26066), .B(n16484), .Z(n16487) );
  AND U24108 ( .A(n16485), .B(n26067), .Z(n16486) );
  NAND U24109 ( .A(n16487), .B(n16486), .Z(n16488) );
  NANDN U24110 ( .A(n26068), .B(n16488), .Z(n16489) );
  NAND U24111 ( .A(n26069), .B(n16489), .Z(n16490) );
  NANDN U24112 ( .A(n26070), .B(n16490), .Z(n16491) );
  AND U24113 ( .A(n26071), .B(n16491), .Z(n16492) );
  OR U24114 ( .A(n26072), .B(n16492), .Z(n16493) );
  AND U24115 ( .A(n16494), .B(n16493), .Z(n16495) );
  OR U24116 ( .A(n16496), .B(n16495), .Z(n16497) );
  AND U24117 ( .A(n16498), .B(n16497), .Z(n16501) );
  NANDN U24118 ( .A(n16501), .B(n26077), .Z(n16502) );
  AND U24119 ( .A(n16503), .B(n16502), .Z(n16504) );
  NOR U24120 ( .A(n16505), .B(n16504), .Z(n16506) );
  NANDN U24121 ( .A(n16507), .B(n16506), .Z(n16508) );
  AND U24122 ( .A(n16509), .B(n16508), .Z(n16511) );
  NAND U24123 ( .A(n16511), .B(n16510), .Z(n16513) );
  ANDN U24124 ( .B(n16513), .A(n16512), .Z(n16514) );
  NANDN U24125 ( .A(n16515), .B(n16514), .Z(n16519) );
  AND U24126 ( .A(n16517), .B(n16516), .Z(n16518) );
  NAND U24127 ( .A(n16519), .B(n16518), .Z(n16520) );
  NANDN U24128 ( .A(n16521), .B(n16520), .Z(n16523) );
  OR U24129 ( .A(n16523), .B(n16522), .Z(n16524) );
  AND U24130 ( .A(n16525), .B(n16524), .Z(n16526) );
  NOR U24131 ( .A(n26086), .B(n16526), .Z(n16527) );
  NANDN U24132 ( .A(n16528), .B(n16527), .Z(n16529) );
  AND U24133 ( .A(n26087), .B(n16529), .Z(n16532) );
  NANDN U24134 ( .A(n16532), .B(n26088), .Z(n16533) );
  NAND U24135 ( .A(n26089), .B(n16533), .Z(n16534) );
  NANDN U24136 ( .A(n24501), .B(n16534), .Z(n16537) );
  AND U24137 ( .A(n16535), .B(n26090), .Z(n16536) );
  NAND U24138 ( .A(n16537), .B(n16536), .Z(n16538) );
  NANDN U24139 ( .A(n16539), .B(n16538), .Z(n16542) );
  AND U24140 ( .A(n16540), .B(n26093), .Z(n16541) );
  NAND U24141 ( .A(n16542), .B(n16541), .Z(n16543) );
  NAND U24142 ( .A(n26096), .B(n16543), .Z(n16546) );
  AND U24143 ( .A(n16544), .B(n24499), .Z(n16545) );
  NAND U24144 ( .A(n16546), .B(n16545), .Z(n16547) );
  NANDN U24145 ( .A(n16548), .B(n16547), .Z(n16551) );
  AND U24146 ( .A(n16549), .B(n26100), .Z(n16550) );
  NAND U24147 ( .A(n16551), .B(n16550), .Z(n16552) );
  NANDN U24148 ( .A(n24498), .B(n16552), .Z(n16555) );
  AND U24149 ( .A(n16553), .B(n24497), .Z(n16554) );
  NAND U24150 ( .A(n16555), .B(n16554), .Z(n16556) );
  NANDN U24151 ( .A(n16557), .B(n16556), .Z(n16558) );
  NAND U24152 ( .A(n16559), .B(n16558), .Z(n16560) );
  NAND U24153 ( .A(n26107), .B(n16560), .Z(n16563) );
  AND U24154 ( .A(n16562), .B(n16561), .Z(n24496) );
  AND U24155 ( .A(n16563), .B(n24496), .Z(n16566) );
  NANDN U24156 ( .A(n16566), .B(n26110), .Z(n16567) );
  NAND U24157 ( .A(n26111), .B(n16567), .Z(n16568) );
  NAND U24158 ( .A(n26112), .B(n16568), .Z(n16569) );
  NANDN U24159 ( .A(n26113), .B(n16569), .Z(n16570) );
  AND U24160 ( .A(n26114), .B(n16570), .Z(n16571) );
  NOR U24161 ( .A(n16571), .B(n26115), .Z(n16572) );
  NANDN U24162 ( .A(n16573), .B(n16572), .Z(n16574) );
  AND U24163 ( .A(n16575), .B(n16574), .Z(n16576) );
  AND U24164 ( .A(n16576), .B(n26116), .Z(n16577) );
  OR U24165 ( .A(n16578), .B(n16577), .Z(n16579) );
  NAND U24166 ( .A(n16580), .B(n16579), .Z(n16581) );
  NANDN U24167 ( .A(n16582), .B(n16581), .Z(n16586) );
  AND U24168 ( .A(n16584), .B(n16583), .Z(n16585) );
  NAND U24169 ( .A(n16586), .B(n16585), .Z(n16587) );
  NANDN U24170 ( .A(n16588), .B(n16587), .Z(n16589) );
  OR U24171 ( .A(n16589), .B(n26119), .Z(n16590) );
  AND U24172 ( .A(n16591), .B(n16590), .Z(n16592) );
  NANDN U24173 ( .A(n26120), .B(n16592), .Z(n16593) );
  NAND U24174 ( .A(n26122), .B(n16593), .Z(n16594) );
  NANDN U24175 ( .A(n26123), .B(n16594), .Z(n16595) );
  NAND U24176 ( .A(n26124), .B(n16595), .Z(n16596) );
  NANDN U24177 ( .A(n26125), .B(n16596), .Z(n16598) );
  IV U24178 ( .A(n16597), .Z(n26126) );
  AND U24179 ( .A(n16598), .B(n26126), .Z(n16599) );
  NAND U24180 ( .A(n16599), .B(n26127), .Z(n16600) );
  NAND U24181 ( .A(n24491), .B(n16600), .Z(n16601) );
  AND U24182 ( .A(n16602), .B(n16601), .Z(n16603) );
  NAND U24183 ( .A(n16603), .B(n26128), .Z(n16604) );
  NANDN U24184 ( .A(n16605), .B(n16604), .Z(n16606) );
  AND U24185 ( .A(n16607), .B(n16606), .Z(n16608) );
  NAND U24186 ( .A(n16608), .B(n26132), .Z(n16609) );
  NAND U24187 ( .A(n26133), .B(n16609), .Z(n16610) );
  AND U24188 ( .A(n16611), .B(n16610), .Z(n16612) );
  NAND U24189 ( .A(n24490), .B(n16612), .Z(n16614) );
  ANDN U24190 ( .B(n16614), .A(n16613), .Z(n16615) );
  NANDN U24191 ( .A(n24489), .B(n16615), .Z(n16617) );
  AND U24192 ( .A(n16617), .B(n16616), .Z(n16618) );
  NAND U24193 ( .A(n16619), .B(n16618), .Z(n16620) );
  NAND U24194 ( .A(n16621), .B(n16620), .Z(n16622) );
  AND U24195 ( .A(n16623), .B(n16622), .Z(n16624) );
  OR U24196 ( .A(n16624), .B(n26137), .Z(n16625) );
  NAND U24197 ( .A(n26138), .B(n16625), .Z(n16626) );
  NANDN U24198 ( .A(n26139), .B(n16626), .Z(n16627) );
  NANDN U24199 ( .A(n24487), .B(n16627), .Z(n16628) );
  AND U24200 ( .A(n26140), .B(n16628), .Z(n16629) );
  ANDN U24201 ( .B(n16630), .A(n16629), .Z(n16631) );
  NAND U24202 ( .A(n26141), .B(n16631), .Z(n16632) );
  NANDN U24203 ( .A(n16633), .B(n16632), .Z(n16634) );
  OR U24204 ( .A(n16634), .B(n26142), .Z(n16635) );
  NAND U24205 ( .A(n16636), .B(n16635), .Z(n16637) );
  NANDN U24206 ( .A(n16638), .B(n16637), .Z(n16641) );
  AND U24207 ( .A(n16639), .B(n26146), .Z(n16640) );
  NAND U24208 ( .A(n16641), .B(n16640), .Z(n16642) );
  NANDN U24209 ( .A(n26147), .B(n16642), .Z(n16645) );
  AND U24210 ( .A(n16643), .B(n26148), .Z(n16644) );
  NAND U24211 ( .A(n16645), .B(n16644), .Z(n16646) );
  NANDN U24212 ( .A(n26149), .B(n16646), .Z(n16648) );
  IV U24213 ( .A(n16647), .Z(n26152) );
  OR U24214 ( .A(n16648), .B(n26152), .Z(n16649) );
  AND U24215 ( .A(n16650), .B(n16649), .Z(n16651) );
  OR U24216 ( .A(n26154), .B(n16651), .Z(n16652) );
  NAND U24217 ( .A(n26155), .B(n16652), .Z(n16653) );
  NANDN U24218 ( .A(n26156), .B(n16653), .Z(n16654) );
  NAND U24219 ( .A(n26157), .B(n16654), .Z(n16655) );
  NANDN U24220 ( .A(n26158), .B(n16655), .Z(n16656) );
  AND U24221 ( .A(n26159), .B(n16656), .Z(n16657) );
  OR U24222 ( .A(n26160), .B(n16657), .Z(n16658) );
  NAND U24223 ( .A(n26161), .B(n16658), .Z(n16659) );
  NANDN U24224 ( .A(n26162), .B(n16659), .Z(n16660) );
  NAND U24225 ( .A(n26163), .B(n16660), .Z(n16661) );
  NANDN U24226 ( .A(n26164), .B(n16661), .Z(n16662) );
  AND U24227 ( .A(n26165), .B(n16662), .Z(n16665) );
  NAND U24228 ( .A(n16664), .B(n16663), .Z(n26166) );
  OR U24229 ( .A(n16665), .B(n26166), .Z(n16666) );
  AND U24230 ( .A(n16667), .B(n16666), .Z(n16668) );
  NAND U24231 ( .A(n16668), .B(n26167), .Z(n16670) );
  ANDN U24232 ( .B(n16670), .A(n16669), .Z(n16671) );
  NANDN U24233 ( .A(n26168), .B(n16671), .Z(n16675) );
  AND U24234 ( .A(n16673), .B(n16672), .Z(n16674) );
  NAND U24235 ( .A(n16675), .B(n16674), .Z(n16676) );
  NANDN U24236 ( .A(n16677), .B(n16676), .Z(n16678) );
  OR U24237 ( .A(n16679), .B(n16678), .Z(n16680) );
  AND U24238 ( .A(n16681), .B(n16680), .Z(n16682) );
  NANDN U24239 ( .A(n26174), .B(n16682), .Z(n16683) );
  AND U24240 ( .A(n16684), .B(n16683), .Z(n16685) );
  NAND U24241 ( .A(n16685), .B(n26175), .Z(n16686) );
  NANDN U24242 ( .A(n26176), .B(n16686), .Z(n16687) );
  AND U24243 ( .A(n26177), .B(n16687), .Z(n16688) );
  OR U24244 ( .A(n26178), .B(n16688), .Z(n16689) );
  NAND U24245 ( .A(n26179), .B(n16689), .Z(n16690) );
  NANDN U24246 ( .A(n26180), .B(n16690), .Z(n16691) );
  NAND U24247 ( .A(n26181), .B(n16691), .Z(n16694) );
  AND U24248 ( .A(n16693), .B(n16692), .Z(n24485) );
  AND U24249 ( .A(n16694), .B(n24485), .Z(n16697) );
  NANDN U24250 ( .A(n16697), .B(n26182), .Z(n16698) );
  AND U24251 ( .A(n16699), .B(n16698), .Z(n16700) );
  OR U24252 ( .A(n16701), .B(n16700), .Z(n16702) );
  AND U24253 ( .A(n16703), .B(n16702), .Z(n16704) );
  OR U24254 ( .A(n16705), .B(n16704), .Z(n16706) );
  NAND U24255 ( .A(n16707), .B(n16706), .Z(n16708) );
  NAND U24256 ( .A(n16709), .B(n16708), .Z(n16713) );
  AND U24257 ( .A(n16711), .B(n16710), .Z(n16712) );
  NAND U24258 ( .A(n16713), .B(n16712), .Z(n16714) );
  NAND U24259 ( .A(n16715), .B(n16714), .Z(n16716) );
  OR U24260 ( .A(n16716), .B(n26187), .Z(n16717) );
  NAND U24261 ( .A(n26190), .B(n16717), .Z(n16718) );
  NAND U24262 ( .A(n26191), .B(n16718), .Z(n16719) );
  NAND U24263 ( .A(n26192), .B(n16719), .Z(n16720) );
  NAND U24264 ( .A(n26193), .B(n16720), .Z(n16721) );
  AND U24265 ( .A(n16722), .B(n16721), .Z(n16723) );
  NAND U24266 ( .A(n24483), .B(n16723), .Z(n16725) );
  ANDN U24267 ( .B(n16725), .A(n16724), .Z(n16726) );
  NANDN U24268 ( .A(n26194), .B(n16726), .Z(n16730) );
  AND U24269 ( .A(n16728), .B(n16727), .Z(n16729) );
  NAND U24270 ( .A(n16730), .B(n16729), .Z(n16731) );
  NANDN U24271 ( .A(n16732), .B(n16731), .Z(n16733) );
  OR U24272 ( .A(n16734), .B(n16733), .Z(n16735) );
  AND U24273 ( .A(n16736), .B(n16735), .Z(n16737) );
  NANDN U24274 ( .A(n16738), .B(n16737), .Z(n16739) );
  AND U24275 ( .A(n16740), .B(n16739), .Z(n16741) );
  NAND U24276 ( .A(n26199), .B(n16741), .Z(n16742) );
  AND U24277 ( .A(n26200), .B(n16742), .Z(n16743) );
  NANDN U24278 ( .A(n16744), .B(n16743), .Z(n16745) );
  NAND U24279 ( .A(n26201), .B(n16745), .Z(n16746) );
  NANDN U24280 ( .A(n16747), .B(n16746), .Z(n16748) );
  AND U24281 ( .A(n16749), .B(n16748), .Z(n16753) );
  NAND U24282 ( .A(n16751), .B(n16750), .Z(n16752) );
  OR U24283 ( .A(n16753), .B(n16752), .Z(n16754) );
  AND U24284 ( .A(n16755), .B(n16754), .Z(n16757) );
  NAND U24285 ( .A(n16757), .B(n16756), .Z(n16759) );
  ANDN U24286 ( .B(n16759), .A(n16758), .Z(n16760) );
  NANDN U24287 ( .A(n16761), .B(n16760), .Z(n16764) );
  AND U24288 ( .A(n16762), .B(n26207), .Z(n16763) );
  NAND U24289 ( .A(n16764), .B(n16763), .Z(n16765) );
  NANDN U24290 ( .A(n16766), .B(n16765), .Z(n16767) );
  OR U24291 ( .A(n16767), .B(n24480), .Z(n16770) );
  AND U24292 ( .A(n16769), .B(n16768), .Z(n24479) );
  AND U24293 ( .A(n16770), .B(n24479), .Z(n16773) );
  NANDN U24294 ( .A(n16773), .B(n26208), .Z(n16774) );
  NANDN U24295 ( .A(n26209), .B(n16774), .Z(n16775) );
  AND U24296 ( .A(n26210), .B(n16775), .Z(n16776) );
  OR U24297 ( .A(n26211), .B(n16776), .Z(n16777) );
  NAND U24298 ( .A(n26212), .B(n16777), .Z(n16778) );
  NANDN U24299 ( .A(n26213), .B(n16778), .Z(n16781) );
  AND U24300 ( .A(n16779), .B(n26214), .Z(n16780) );
  NAND U24301 ( .A(n16781), .B(n16780), .Z(n16782) );
  NANDN U24302 ( .A(n26218), .B(n16782), .Z(n16783) );
  OR U24303 ( .A(n16783), .B(n26215), .Z(n16784) );
  AND U24304 ( .A(n16785), .B(n16784), .Z(n16787) );
  NAND U24305 ( .A(n24477), .B(n26219), .Z(n16786) );
  OR U24306 ( .A(n16787), .B(n16786), .Z(n16788) );
  AND U24307 ( .A(n16789), .B(n16788), .Z(n16790) );
  NAND U24308 ( .A(n16790), .B(n26220), .Z(n16791) );
  NANDN U24309 ( .A(n24476), .B(n16791), .Z(n16792) );
  AND U24310 ( .A(n26221), .B(n16792), .Z(n16795) );
  NAND U24311 ( .A(n16794), .B(n16793), .Z(n24475) );
  OR U24312 ( .A(n16795), .B(n24475), .Z(n16796) );
  AND U24313 ( .A(n26222), .B(n16796), .Z(n16797) );
  OR U24314 ( .A(n26223), .B(n16797), .Z(n16798) );
  NAND U24315 ( .A(n26224), .B(n16798), .Z(n16799) );
  NANDN U24316 ( .A(n26225), .B(n16799), .Z(n16802) );
  AND U24317 ( .A(n16800), .B(n26226), .Z(n16801) );
  NAND U24318 ( .A(n16802), .B(n16801), .Z(n16803) );
  NAND U24319 ( .A(n26227), .B(n16803), .Z(n16804) );
  NAND U24320 ( .A(n16805), .B(n16804), .Z(n16806) );
  NANDN U24321 ( .A(n16807), .B(n16806), .Z(n16808) );
  AND U24322 ( .A(n16809), .B(n16808), .Z(n16811) );
  NAND U24323 ( .A(n16811), .B(n16810), .Z(n16813) );
  ANDN U24324 ( .B(n16813), .A(n16812), .Z(n16814) );
  NANDN U24325 ( .A(n16815), .B(n16814), .Z(n16819) );
  AND U24326 ( .A(n16817), .B(n16816), .Z(n16818) );
  NAND U24327 ( .A(n16819), .B(n16818), .Z(n16820) );
  NAND U24328 ( .A(n16821), .B(n16820), .Z(n16825) );
  AND U24329 ( .A(n16823), .B(n16822), .Z(n16824) );
  NAND U24330 ( .A(n16825), .B(n16824), .Z(n16826) );
  NAND U24331 ( .A(n26235), .B(n16826), .Z(n16827) );
  NAND U24332 ( .A(n16828), .B(n16827), .Z(n16829) );
  NANDN U24333 ( .A(n26237), .B(n16829), .Z(n16830) );
  AND U24334 ( .A(n26238), .B(n16830), .Z(n16831) );
  OR U24335 ( .A(n26239), .B(n16831), .Z(n16832) );
  NAND U24336 ( .A(n26240), .B(n16832), .Z(n16833) );
  NANDN U24337 ( .A(n24474), .B(n16833), .Z(n16834) );
  NAND U24338 ( .A(n24473), .B(n16834), .Z(n16835) );
  NAND U24339 ( .A(n26241), .B(n16835), .Z(n16836) );
  NANDN U24340 ( .A(n26242), .B(n16836), .Z(n16837) );
  NAND U24341 ( .A(n26243), .B(n16837), .Z(n16838) );
  NAND U24342 ( .A(n26244), .B(n16838), .Z(n16839) );
  NAND U24343 ( .A(n26245), .B(n16839), .Z(n16840) );
  NAND U24344 ( .A(n24472), .B(n16840), .Z(n16841) );
  NAND U24345 ( .A(n26248), .B(n16841), .Z(n16842) );
  AND U24346 ( .A(n16843), .B(n16842), .Z(n16844) );
  NANDN U24347 ( .A(n26249), .B(n16844), .Z(n16845) );
  NAND U24348 ( .A(n16846), .B(n16845), .Z(n16849) );
  AND U24349 ( .A(n16847), .B(n26253), .Z(n16848) );
  NAND U24350 ( .A(n16849), .B(n16848), .Z(n16850) );
  NAND U24351 ( .A(n26254), .B(n16850), .Z(n16853) );
  AND U24352 ( .A(n16851), .B(n24471), .Z(n16852) );
  NAND U24353 ( .A(n16853), .B(n16852), .Z(n16854) );
  NANDN U24354 ( .A(n16855), .B(n16854), .Z(n16856) );
  OR U24355 ( .A(n16856), .B(n26255), .Z(n16857) );
  NAND U24356 ( .A(n16858), .B(n16857), .Z(n16859) );
  NANDN U24357 ( .A(n16860), .B(n16859), .Z(n16864) );
  NOR U24358 ( .A(n16862), .B(n16861), .Z(n16863) );
  NAND U24359 ( .A(n16864), .B(n16863), .Z(n16865) );
  AND U24360 ( .A(n16866), .B(n16865), .Z(n16867) );
  NAND U24361 ( .A(n26261), .B(n16867), .Z(n16868) );
  ANDN U24362 ( .B(n16868), .A(n26262), .Z(n16869) );
  NANDN U24363 ( .A(n16870), .B(n16869), .Z(n16871) );
  NAND U24364 ( .A(n26263), .B(n16871), .Z(n16872) );
  ANDN U24365 ( .B(n16872), .A(n26264), .Z(n16873) );
  NANDN U24366 ( .A(n16874), .B(n16873), .Z(n16877) );
  AND U24367 ( .A(n16875), .B(n26265), .Z(n16876) );
  NAND U24368 ( .A(n16877), .B(n16876), .Z(n16878) );
  NANDN U24369 ( .A(n16879), .B(n16878), .Z(n16880) );
  OR U24370 ( .A(n16881), .B(n16880), .Z(n16882) );
  AND U24371 ( .A(n16883), .B(n16882), .Z(n16884) );
  NAND U24372 ( .A(n26269), .B(n16884), .Z(n16885) );
  AND U24373 ( .A(n26270), .B(n16885), .Z(n16886) );
  NANDN U24374 ( .A(n16887), .B(n16886), .Z(n16888) );
  NAND U24375 ( .A(n26271), .B(n16888), .Z(n16889) );
  NAND U24376 ( .A(n16890), .B(n16889), .Z(n16891) );
  NANDN U24377 ( .A(n24468), .B(n16891), .Z(n16894) );
  AND U24378 ( .A(n26272), .B(n16892), .Z(n16893) );
  NAND U24379 ( .A(n16894), .B(n16893), .Z(n16895) );
  NAND U24380 ( .A(n26273), .B(n16895), .Z(n16896) );
  NAND U24381 ( .A(n26274), .B(n16896), .Z(n16897) );
  NAND U24382 ( .A(n16898), .B(n16897), .Z(n16899) );
  NANDN U24383 ( .A(n16900), .B(n16899), .Z(n16904) );
  AND U24384 ( .A(n16902), .B(n16901), .Z(n16903) );
  NAND U24385 ( .A(n16904), .B(n16903), .Z(n16905) );
  NANDN U24386 ( .A(n16906), .B(n16905), .Z(n16908) );
  IV U24387 ( .A(n16907), .Z(n26278) );
  OR U24388 ( .A(n16908), .B(n26278), .Z(n16909) );
  AND U24389 ( .A(n16910), .B(n16909), .Z(n16911) );
  NAND U24390 ( .A(n26279), .B(n16911), .Z(n16912) );
  NANDN U24391 ( .A(n26280), .B(n16912), .Z(n16913) );
  AND U24392 ( .A(n26281), .B(n16913), .Z(n16914) );
  OR U24393 ( .A(n26282), .B(n16914), .Z(n16915) );
  NAND U24394 ( .A(n26283), .B(n16915), .Z(n16916) );
  NANDN U24395 ( .A(n24465), .B(n16916), .Z(n16917) );
  NANDN U24396 ( .A(n26284), .B(n16917), .Z(n16918) );
  NAND U24397 ( .A(n26285), .B(n16918), .Z(n16919) );
  AND U24398 ( .A(n24464), .B(n16919), .Z(n16920) );
  NANDN U24399 ( .A(n16921), .B(n16920), .Z(n16922) );
  AND U24400 ( .A(n16923), .B(n16922), .Z(n16924) );
  ANDN U24401 ( .B(n16925), .A(n16924), .Z(n16926) );
  NAND U24402 ( .A(n16927), .B(n16926), .Z(n16928) );
  NANDN U24403 ( .A(n16929), .B(n16928), .Z(n16931) );
  OR U24404 ( .A(n16931), .B(n16930), .Z(n16932) );
  NAND U24405 ( .A(n16933), .B(n16932), .Z(n16934) );
  NANDN U24406 ( .A(n16935), .B(n16934), .Z(n16939) );
  AND U24407 ( .A(n24462), .B(n24461), .Z(n16937) );
  OR U24408 ( .A(n16937), .B(n16936), .Z(n16938) );
  AND U24409 ( .A(n16939), .B(n16938), .Z(n16940) );
  NANDN U24410 ( .A(n16940), .B(n26292), .Z(n16941) );
  NAND U24411 ( .A(n26293), .B(n16941), .Z(n16942) );
  NAND U24412 ( .A(n26294), .B(n16942), .Z(n16943) );
  NAND U24413 ( .A(n26295), .B(n16943), .Z(n16945) );
  IV U24414 ( .A(n16944), .Z(n26296) );
  ANDN U24415 ( .B(n16945), .A(n26296), .Z(n16946) );
  NANDN U24416 ( .A(n16947), .B(n16946), .Z(n16948) );
  NAND U24417 ( .A(n26297), .B(n16948), .Z(n16950) );
  ANDN U24418 ( .B(n16950), .A(n16949), .Z(n16951) );
  NANDN U24419 ( .A(n16952), .B(n16951), .Z(n16953) );
  NAND U24420 ( .A(n26299), .B(n16953), .Z(n16954) );
  NANDN U24421 ( .A(n16955), .B(n16954), .Z(n16956) );
  AND U24422 ( .A(n16956), .B(n24460), .Z(n16957) );
  OR U24423 ( .A(n16957), .B(n26301), .Z(n16958) );
  AND U24424 ( .A(n16958), .B(n26302), .Z(n16959) );
  OR U24425 ( .A(n16959), .B(n26303), .Z(n16960) );
  NAND U24426 ( .A(n26306), .B(n16960), .Z(n16961) );
  NAND U24427 ( .A(n26307), .B(n16961), .Z(n16962) );
  NAND U24428 ( .A(n24459), .B(n16962), .Z(n16963) );
  AND U24429 ( .A(n16964), .B(n16963), .Z(n16965) );
  OR U24430 ( .A(n16966), .B(n16965), .Z(n16967) );
  AND U24431 ( .A(n16968), .B(n16967), .Z(n16971) );
  NAND U24432 ( .A(n16970), .B(n16969), .Z(n26313) );
  OR U24433 ( .A(n16971), .B(n26313), .Z(n16972) );
  NAND U24434 ( .A(n16973), .B(n16972), .Z(n16974) );
  NAND U24435 ( .A(n26315), .B(n16974), .Z(n16975) );
  AND U24436 ( .A(n16976), .B(n16975), .Z(n16977) );
  OR U24437 ( .A(n26319), .B(n16977), .Z(n16978) );
  NAND U24438 ( .A(n26321), .B(n16978), .Z(n16979) );
  NANDN U24439 ( .A(n26322), .B(n16979), .Z(n16983) );
  IV U24440 ( .A(n16980), .Z(n26323) );
  AND U24441 ( .A(n16981), .B(n26323), .Z(n16982) );
  NAND U24442 ( .A(n16983), .B(n16982), .Z(n16984) );
  NANDN U24443 ( .A(n16985), .B(n16984), .Z(n16987) );
  IV U24444 ( .A(n16986), .Z(n26324) );
  OR U24445 ( .A(n16987), .B(n26324), .Z(n16988) );
  AND U24446 ( .A(n16989), .B(n16988), .Z(n16990) );
  NOR U24447 ( .A(n24458), .B(n16990), .Z(n16991) );
  NANDN U24448 ( .A(n16992), .B(n16991), .Z(n16995) );
  AND U24449 ( .A(n16994), .B(n16993), .Z(n24457) );
  AND U24450 ( .A(n16995), .B(n24457), .Z(n16998) );
  NANDN U24451 ( .A(n16998), .B(n26328), .Z(n16999) );
  AND U24452 ( .A(n17000), .B(n16999), .Z(n17001) );
  NAND U24453 ( .A(n24456), .B(n17001), .Z(n17003) );
  ANDN U24454 ( .B(n17003), .A(n17002), .Z(n17004) );
  NANDN U24455 ( .A(n26329), .B(n17004), .Z(n17008) );
  AND U24456 ( .A(n17006), .B(n17005), .Z(n17007) );
  NAND U24457 ( .A(n17008), .B(n17007), .Z(n17009) );
  NANDN U24458 ( .A(n17010), .B(n17009), .Z(n17011) );
  OR U24459 ( .A(n17011), .B(n26333), .Z(n17012) );
  NAND U24460 ( .A(n17013), .B(n17012), .Z(n17014) );
  NANDN U24461 ( .A(n17015), .B(n17014), .Z(n17017) );
  OR U24462 ( .A(n17017), .B(n17016), .Z(n17018) );
  AND U24463 ( .A(n17019), .B(n17018), .Z(n17020) );
  OR U24464 ( .A(n17021), .B(n17020), .Z(n17022) );
  NAND U24465 ( .A(n24452), .B(n17022), .Z(n17023) );
  NANDN U24466 ( .A(n26337), .B(n17023), .Z(n17024) );
  NAND U24467 ( .A(n26338), .B(n17024), .Z(n17025) );
  NANDN U24468 ( .A(n26339), .B(n17025), .Z(n17028) );
  XNOR U24469 ( .A(x[1142]), .B(y[1142]), .Z(n17026) );
  AND U24470 ( .A(n17027), .B(n17026), .Z(n24450) );
  AND U24471 ( .A(n17028), .B(n24450), .Z(n17031) );
  NANDN U24472 ( .A(n17031), .B(n26340), .Z(n17032) );
  NAND U24473 ( .A(n26341), .B(n17032), .Z(n17033) );
  NANDN U24474 ( .A(n24449), .B(n17033), .Z(n17034) );
  NAND U24475 ( .A(n24448), .B(n17034), .Z(n17035) );
  AND U24476 ( .A(n26344), .B(n17035), .Z(n17036) );
  NANDN U24477 ( .A(n17037), .B(n17036), .Z(n17038) );
  AND U24478 ( .A(n17039), .B(n17038), .Z(n17040) );
  ANDN U24479 ( .B(n17041), .A(n17040), .Z(n17042) );
  NAND U24480 ( .A(n17043), .B(n17042), .Z(n17044) );
  NANDN U24481 ( .A(n17045), .B(n17044), .Z(n17047) );
  IV U24482 ( .A(n17046), .Z(n26347) );
  OR U24483 ( .A(n17047), .B(n26347), .Z(n17048) );
  AND U24484 ( .A(n17049), .B(n17048), .Z(n17050) );
  NANDN U24485 ( .A(n26348), .B(n17050), .Z(n17051) );
  NAND U24486 ( .A(n26349), .B(n17051), .Z(n17052) );
  NANDN U24487 ( .A(n24447), .B(n17052), .Z(n17055) );
  AND U24488 ( .A(n17053), .B(n26350), .Z(n17054) );
  NAND U24489 ( .A(n17055), .B(n17054), .Z(n17056) );
  NANDN U24490 ( .A(n17057), .B(n17056), .Z(n17058) );
  OR U24491 ( .A(n17058), .B(n26351), .Z(n17059) );
  NAND U24492 ( .A(n17060), .B(n17059), .Z(n17061) );
  NAND U24493 ( .A(n17062), .B(n17061), .Z(n17065) );
  AND U24494 ( .A(n17063), .B(n26355), .Z(n17064) );
  NAND U24495 ( .A(n17065), .B(n17064), .Z(n17066) );
  NAND U24496 ( .A(n26358), .B(n17066), .Z(n17070) );
  IV U24497 ( .A(n17067), .Z(n26359) );
  NOR U24498 ( .A(n26359), .B(n17068), .Z(n17069) );
  NAND U24499 ( .A(n17070), .B(n17069), .Z(n17071) );
  AND U24500 ( .A(n17072), .B(n17071), .Z(n17073) );
  NAND U24501 ( .A(n26360), .B(n17073), .Z(n17075) );
  ANDN U24502 ( .B(n17075), .A(n17074), .Z(n17076) );
  NANDN U24503 ( .A(n17077), .B(n17076), .Z(n17078) );
  AND U24504 ( .A(n17079), .B(n17078), .Z(n17080) );
  NAND U24505 ( .A(n26364), .B(n17080), .Z(n17081) );
  NANDN U24506 ( .A(n26365), .B(n17081), .Z(n17083) );
  OR U24507 ( .A(n17083), .B(n17082), .Z(n17084) );
  NANDN U24508 ( .A(n26366), .B(n17084), .Z(n17086) );
  IV U24509 ( .A(n17085), .Z(n26367) );
  AND U24510 ( .A(n17086), .B(n26367), .Z(n17088) );
  IV U24511 ( .A(n17087), .Z(n26368) );
  OR U24512 ( .A(n17088), .B(n26368), .Z(n17089) );
  NAND U24513 ( .A(n26369), .B(n17089), .Z(n17090) );
  NANDN U24514 ( .A(n26370), .B(n17090), .Z(n17091) );
  NAND U24515 ( .A(n26371), .B(n17091), .Z(n17092) );
  NANDN U24516 ( .A(n26372), .B(n17092), .Z(n17093) );
  AND U24517 ( .A(n26373), .B(n17093), .Z(n17094) );
  OR U24518 ( .A(n26374), .B(n17094), .Z(n17095) );
  NAND U24519 ( .A(n24446), .B(n17095), .Z(n17096) );
  NAND U24520 ( .A(n26375), .B(n17096), .Z(n17097) );
  NAND U24521 ( .A(n17098), .B(n17097), .Z(n17099) );
  NAND U24522 ( .A(n17100), .B(n17099), .Z(n17101) );
  NAND U24523 ( .A(n17102), .B(n17101), .Z(n17103) );
  NAND U24524 ( .A(n17104), .B(n17103), .Z(n17105) );
  NANDN U24525 ( .A(n17106), .B(n17105), .Z(n17108) );
  OR U24526 ( .A(n17108), .B(n17107), .Z(n17109) );
  AND U24527 ( .A(n17110), .B(n17109), .Z(n17112) );
  NAND U24528 ( .A(n17112), .B(n17111), .Z(n17114) );
  ANDN U24529 ( .B(n17114), .A(n17113), .Z(n17115) );
  NANDN U24530 ( .A(n17116), .B(n17115), .Z(n17117) );
  AND U24531 ( .A(n17118), .B(n17117), .Z(n17119) );
  NAND U24532 ( .A(n26383), .B(n17119), .Z(n17120) );
  NAND U24533 ( .A(n26384), .B(n17120), .Z(n17122) );
  OR U24534 ( .A(n17122), .B(n17121), .Z(n17123) );
  NAND U24535 ( .A(n26385), .B(n17123), .Z(n17124) );
  NANDN U24536 ( .A(n26386), .B(n17124), .Z(n17125) );
  NAND U24537 ( .A(n17126), .B(n17125), .Z(n17127) );
  NAND U24538 ( .A(n17128), .B(n17127), .Z(n17129) );
  NANDN U24539 ( .A(n26389), .B(n17129), .Z(n17130) );
  OR U24540 ( .A(n17131), .B(n17130), .Z(n17132) );
  AND U24541 ( .A(n26390), .B(n17132), .Z(n17134) );
  NAND U24542 ( .A(n17134), .B(n17133), .Z(n17135) );
  NAND U24543 ( .A(n26391), .B(n17135), .Z(n17136) );
  AND U24544 ( .A(n17136), .B(n24444), .Z(n17137) );
  OR U24545 ( .A(n17137), .B(n26394), .Z(n17138) );
  AND U24546 ( .A(n17139), .B(n17138), .Z(n17140) );
  NANDN U24547 ( .A(n26396), .B(n17140), .Z(n17141) );
  NAND U24548 ( .A(n17142), .B(n17141), .Z(n17146) );
  AND U24549 ( .A(n17144), .B(n17143), .Z(n17145) );
  NAND U24550 ( .A(n17146), .B(n17145), .Z(n17147) );
  NAND U24551 ( .A(n24440), .B(n17147), .Z(n17150) );
  ANDN U24552 ( .B(n24439), .A(n17148), .Z(n17149) );
  NAND U24553 ( .A(n17150), .B(n17149), .Z(n17151) );
  AND U24554 ( .A(n17152), .B(n17151), .Z(n17153) );
  NAND U24555 ( .A(n24441), .B(n17153), .Z(n17155) );
  ANDN U24556 ( .B(n17155), .A(n17154), .Z(n17156) );
  NANDN U24557 ( .A(n26400), .B(n17156), .Z(n17160) );
  IV U24558 ( .A(n17157), .Z(n26401) );
  AND U24559 ( .A(n17158), .B(n26401), .Z(n17159) );
  NAND U24560 ( .A(n17160), .B(n17159), .Z(n17161) );
  NANDN U24561 ( .A(n26402), .B(n17161), .Z(n17162) );
  NAND U24562 ( .A(n26403), .B(n17162), .Z(n17163) );
  AND U24563 ( .A(n26404), .B(n17163), .Z(n17166) );
  NANDN U24564 ( .A(x[1206]), .B(y[1206]), .Z(n17165) );
  AND U24565 ( .A(n17165), .B(n17164), .Z(n26406) );
  NANDN U24566 ( .A(n17166), .B(n26406), .Z(n17167) );
  NAND U24567 ( .A(n17168), .B(n17167), .Z(n17171) );
  AND U24568 ( .A(n17169), .B(n26409), .Z(n17170) );
  NAND U24569 ( .A(n17171), .B(n17170), .Z(n17172) );
  NANDN U24570 ( .A(n17173), .B(n17172), .Z(n17174) );
  OR U24571 ( .A(n17175), .B(n17174), .Z(n17176) );
  AND U24572 ( .A(n17177), .B(n17176), .Z(n17179) );
  NAND U24573 ( .A(n17179), .B(n17178), .Z(n17181) );
  ANDN U24574 ( .B(n17181), .A(n17180), .Z(n17182) );
  NANDN U24575 ( .A(n17183), .B(n17182), .Z(n17185) );
  AND U24576 ( .A(n17185), .B(n17184), .Z(n17186) );
  NAND U24577 ( .A(n17187), .B(n17186), .Z(n17188) );
  NAND U24578 ( .A(n17189), .B(n17188), .Z(n17190) );
  AND U24579 ( .A(n17191), .B(n17190), .Z(n17193) );
  IV U24580 ( .A(n17192), .Z(n26424) );
  OR U24581 ( .A(n17193), .B(n26424), .Z(n17195) );
  IV U24582 ( .A(n17194), .Z(n26425) );
  AND U24583 ( .A(n17195), .B(n26425), .Z(n17197) );
  IV U24584 ( .A(n17196), .Z(n26427) );
  OR U24585 ( .A(n17197), .B(n26427), .Z(n17198) );
  NAND U24586 ( .A(n26430), .B(n17198), .Z(n17199) );
  NANDN U24587 ( .A(n26432), .B(n17199), .Z(n17200) );
  NAND U24588 ( .A(n26434), .B(n17200), .Z(n17201) );
  AND U24589 ( .A(n17202), .B(n17201), .Z(n17203) );
  OR U24590 ( .A(n17204), .B(n17203), .Z(n17205) );
  NAND U24591 ( .A(n17206), .B(n17205), .Z(n17207) );
  NANDN U24592 ( .A(n26446), .B(n17207), .Z(n17208) );
  NAND U24593 ( .A(n17209), .B(n17208), .Z(n17210) );
  NANDN U24594 ( .A(n26448), .B(n17210), .Z(n17211) );
  AND U24595 ( .A(n17212), .B(n17211), .Z(n17214) );
  OR U24596 ( .A(n17214), .B(n17213), .Z(n17215) );
  AND U24597 ( .A(n17216), .B(n17215), .Z(n17218) );
  NAND U24598 ( .A(n17218), .B(n17217), .Z(n17220) );
  ANDN U24599 ( .B(n17220), .A(n17219), .Z(n17221) );
  NANDN U24600 ( .A(n17222), .B(n17221), .Z(n17226) );
  AND U24601 ( .A(n17224), .B(n17223), .Z(n17225) );
  NAND U24602 ( .A(n17226), .B(n17225), .Z(n17227) );
  NAND U24603 ( .A(n26454), .B(n17227), .Z(n17229) );
  OR U24604 ( .A(n17229), .B(n17228), .Z(n17230) );
  NAND U24605 ( .A(n17231), .B(n17230), .Z(n17232) );
  AND U24606 ( .A(n17233), .B(n17232), .Z(n17234) );
  NAND U24607 ( .A(n26453), .B(n17234), .Z(n17235) );
  NANDN U24608 ( .A(n17236), .B(n17235), .Z(n17237) );
  OR U24609 ( .A(n17237), .B(n26457), .Z(n17238) );
  AND U24610 ( .A(n17239), .B(n17238), .Z(n17240) );
  OR U24611 ( .A(n26459), .B(n17240), .Z(n17241) );
  NAND U24612 ( .A(n26460), .B(n17241), .Z(n17242) );
  NAND U24613 ( .A(n26462), .B(n17242), .Z(n17243) );
  NANDN U24614 ( .A(n26463), .B(n17243), .Z(n17244) );
  AND U24615 ( .A(n17245), .B(n17244), .Z(n17246) );
  NANDN U24616 ( .A(n24436), .B(n17246), .Z(n17247) );
  NAND U24617 ( .A(n17248), .B(n17247), .Z(n17252) );
  IV U24618 ( .A(n17249), .Z(n26467) );
  AND U24619 ( .A(n17250), .B(n26467), .Z(n17251) );
  NAND U24620 ( .A(n17252), .B(n17251), .Z(n17253) );
  NANDN U24621 ( .A(n26468), .B(n17253), .Z(n17257) );
  IV U24622 ( .A(n17254), .Z(n26469) );
  AND U24623 ( .A(n17255), .B(n26469), .Z(n17256) );
  NAND U24624 ( .A(n17257), .B(n17256), .Z(n17258) );
  NANDN U24625 ( .A(n26470), .B(n17258), .Z(n17259) );
  OR U24626 ( .A(n17259), .B(n26472), .Z(n17260) );
  AND U24627 ( .A(n17261), .B(n17260), .Z(n17264) );
  OR U24628 ( .A(n17264), .B(n26474), .Z(n17265) );
  AND U24629 ( .A(n17266), .B(n17265), .Z(n17267) );
  NAND U24630 ( .A(n17267), .B(n26475), .Z(n17268) );
  NAND U24631 ( .A(n26476), .B(n17268), .Z(n17269) );
  AND U24632 ( .A(n17270), .B(n17269), .Z(n17271) );
  OR U24633 ( .A(n17271), .B(n24435), .Z(n17272) );
  NAND U24634 ( .A(n24434), .B(n17272), .Z(n17273) );
  NANDN U24635 ( .A(n24433), .B(n17273), .Z(n17274) );
  NAND U24636 ( .A(n24432), .B(n17274), .Z(n17275) );
  NAND U24637 ( .A(n26480), .B(n17275), .Z(n17276) );
  AND U24638 ( .A(n17277), .B(n17276), .Z(n17278) );
  NANDN U24639 ( .A(n26481), .B(n17278), .Z(n17279) );
  NAND U24640 ( .A(n17280), .B(n17279), .Z(n17284) );
  AND U24641 ( .A(n17282), .B(n17281), .Z(n17283) );
  NAND U24642 ( .A(n17284), .B(n17283), .Z(n17285) );
  NANDN U24643 ( .A(n24429), .B(n17285), .Z(n17288) );
  AND U24644 ( .A(n17286), .B(n24430), .Z(n17287) );
  NAND U24645 ( .A(n17288), .B(n17287), .Z(n17289) );
  NANDN U24646 ( .A(n17290), .B(n17289), .Z(n17291) );
  OR U24647 ( .A(n17291), .B(n24431), .Z(n17292) );
  NAND U24648 ( .A(n17293), .B(n17292), .Z(n17297) );
  AND U24649 ( .A(n17295), .B(n17294), .Z(n17296) );
  NAND U24650 ( .A(n17297), .B(n17296), .Z(n17298) );
  NANDN U24651 ( .A(n17299), .B(n17298), .Z(n17301) );
  IV U24652 ( .A(n17300), .Z(n26489) );
  OR U24653 ( .A(n17301), .B(n26489), .Z(n17302) );
  AND U24654 ( .A(n17303), .B(n17302), .Z(n17304) );
  NAND U24655 ( .A(n26490), .B(n17304), .Z(n17305) );
  NANDN U24656 ( .A(n26491), .B(n17305), .Z(n17306) );
  AND U24657 ( .A(n26492), .B(n17306), .Z(n17308) );
  IV U24658 ( .A(n17307), .Z(n26493) );
  OR U24659 ( .A(n17308), .B(n26493), .Z(n17310) );
  IV U24660 ( .A(n17309), .Z(n26494) );
  AND U24661 ( .A(n17310), .B(n26494), .Z(n17313) );
  NAND U24662 ( .A(n24426), .B(n17311), .Z(n17312) );
  OR U24663 ( .A(n17313), .B(n17312), .Z(n17315) );
  IV U24664 ( .A(n17314), .Z(n26495) );
  AND U24665 ( .A(n17315), .B(n26495), .Z(n17321) );
  OR U24666 ( .A(n17317), .B(n17316), .Z(n17318) );
  AND U24667 ( .A(n17319), .B(n17318), .Z(n17320) );
  NANDN U24668 ( .A(n17321), .B(n17320), .Z(n17322) );
  NAND U24669 ( .A(n26497), .B(n17322), .Z(n17323) );
  NANDN U24670 ( .A(n26498), .B(n17323), .Z(n17324) );
  NAND U24671 ( .A(n26499), .B(n17324), .Z(n17325) );
  ANDN U24672 ( .B(n17325), .A(n26500), .Z(n17326) );
  NANDN U24673 ( .A(n17327), .B(n17326), .Z(n17330) );
  AND U24674 ( .A(n17328), .B(n26501), .Z(n17329) );
  NAND U24675 ( .A(n17330), .B(n17329), .Z(n17331) );
  NANDN U24676 ( .A(n17332), .B(n17331), .Z(n17333) );
  OR U24677 ( .A(n17334), .B(n17333), .Z(n17335) );
  AND U24678 ( .A(n17336), .B(n17335), .Z(n17338) );
  NAND U24679 ( .A(n17338), .B(n17337), .Z(n17340) );
  ANDN U24680 ( .B(n17340), .A(n17339), .Z(n17341) );
  NANDN U24681 ( .A(n17342), .B(n17341), .Z(n17346) );
  AND U24682 ( .A(n17344), .B(n17343), .Z(n17345) );
  NAND U24683 ( .A(n17346), .B(n17345), .Z(n17347) );
  NANDN U24684 ( .A(n17348), .B(n17347), .Z(n17350) );
  OR U24685 ( .A(n17350), .B(n17349), .Z(n17351) );
  NAND U24686 ( .A(n17352), .B(n17351), .Z(n17353) );
  AND U24687 ( .A(n17354), .B(n17353), .Z(n17355) );
  AND U24688 ( .A(n17356), .B(n17355), .Z(n17357) );
  OR U24689 ( .A(n26510), .B(n17357), .Z(n17358) );
  NAND U24690 ( .A(n26511), .B(n17358), .Z(n17359) );
  NANDN U24691 ( .A(n26512), .B(n17359), .Z(n17360) );
  NAND U24692 ( .A(n26513), .B(n17360), .Z(n17361) );
  NAND U24693 ( .A(n26514), .B(n17361), .Z(n17362) );
  AND U24694 ( .A(n17362), .B(n24423), .Z(n17365) );
  NANDN U24695 ( .A(n17365), .B(n26515), .Z(n17366) );
  NAND U24696 ( .A(n17367), .B(n17366), .Z(n17368) );
  NANDN U24697 ( .A(n26517), .B(n17368), .Z(n17369) );
  NAND U24698 ( .A(n17370), .B(n17369), .Z(n17371) );
  NANDN U24699 ( .A(n17372), .B(n17371), .Z(n17373) );
  AND U24700 ( .A(n26522), .B(n17373), .Z(n17374) );
  OR U24701 ( .A(n26523), .B(n17374), .Z(n17375) );
  NAND U24702 ( .A(n26524), .B(n17375), .Z(n17376) );
  NANDN U24703 ( .A(n26525), .B(n17376), .Z(n17380) );
  IV U24704 ( .A(n17377), .Z(n26526) );
  ANDN U24705 ( .B(n26526), .A(n17378), .Z(n17379) );
  NAND U24706 ( .A(n17380), .B(n17379), .Z(n17381) );
  AND U24707 ( .A(n17381), .B(n26527), .Z(n17383) );
  OR U24708 ( .A(n17383), .B(n17382), .Z(n17384) );
  AND U24709 ( .A(n17384), .B(n24420), .Z(n17385) );
  ANDN U24710 ( .B(n17386), .A(n17385), .Z(n17387) );
  NAND U24711 ( .A(n26528), .B(n17387), .Z(n17388) );
  NANDN U24712 ( .A(n26529), .B(n17388), .Z(n17390) );
  IV U24713 ( .A(n17389), .Z(n26531) );
  OR U24714 ( .A(n17390), .B(n26531), .Z(n17391) );
  NAND U24715 ( .A(n17392), .B(n17391), .Z(n17393) );
  NANDN U24716 ( .A(n26534), .B(n17393), .Z(n17396) );
  AND U24717 ( .A(n17394), .B(n26535), .Z(n17395) );
  NAND U24718 ( .A(n17396), .B(n17395), .Z(n17397) );
  NANDN U24719 ( .A(n17398), .B(n17397), .Z(n17399) );
  OR U24720 ( .A(n17399), .B(n24419), .Z(n17400) );
  NAND U24721 ( .A(n17401), .B(n17400), .Z(n17402) );
  NANDN U24722 ( .A(n26537), .B(n17402), .Z(n17403) );
  OR U24723 ( .A(n17404), .B(n17403), .Z(n17405) );
  AND U24724 ( .A(n26538), .B(n17405), .Z(n17406) );
  NANDN U24725 ( .A(n17407), .B(n17406), .Z(n17408) );
  AND U24726 ( .A(n26539), .B(n17408), .Z(n17409) );
  OR U24727 ( .A(n26540), .B(n17409), .Z(n17410) );
  NAND U24728 ( .A(n17411), .B(n17410), .Z(n17412) );
  NANDN U24729 ( .A(n17413), .B(n17412), .Z(n17417) );
  AND U24730 ( .A(n17415), .B(n17414), .Z(n17416) );
  NAND U24731 ( .A(n17417), .B(n17416), .Z(n17418) );
  NANDN U24732 ( .A(n17419), .B(n17418), .Z(n17421) );
  OR U24733 ( .A(n17421), .B(n17420), .Z(n17422) );
  NAND U24734 ( .A(n17423), .B(n17422), .Z(n17426) );
  AND U24735 ( .A(n17424), .B(n26547), .Z(n17425) );
  NAND U24736 ( .A(n17426), .B(n17425), .Z(n17427) );
  NANDN U24737 ( .A(n24416), .B(n17427), .Z(n17430) );
  ANDN U24738 ( .B(n24415), .A(n17428), .Z(n17429) );
  NAND U24739 ( .A(n17430), .B(n17429), .Z(n17431) );
  AND U24740 ( .A(n26548), .B(n17431), .Z(n17433) );
  OR U24741 ( .A(n17433), .B(n17432), .Z(n17434) );
  AND U24742 ( .A(n26549), .B(n17434), .Z(n17435) );
  NANDN U24743 ( .A(n17435), .B(n26550), .Z(n17436) );
  NAND U24744 ( .A(n26551), .B(n17436), .Z(n17437) );
  AND U24745 ( .A(n26552), .B(n17437), .Z(n17438) );
  OR U24746 ( .A(n17438), .B(n26553), .Z(n17439) );
  AND U24747 ( .A(n17439), .B(n26554), .Z(n17441) );
  IV U24748 ( .A(n17440), .Z(n26555) );
  NANDN U24749 ( .A(n17441), .B(n26555), .Z(n17442) );
  NANDN U24750 ( .A(n26557), .B(n17442), .Z(n17444) );
  IV U24751 ( .A(n17443), .Z(n26558) );
  AND U24752 ( .A(n17444), .B(n26558), .Z(n17445) );
  OR U24753 ( .A(n17446), .B(n17445), .Z(n17447) );
  NAND U24754 ( .A(n17448), .B(n17447), .Z(n17449) );
  NANDN U24755 ( .A(n17450), .B(n17449), .Z(n17452) );
  OR U24756 ( .A(n17452), .B(n17451), .Z(n17453) );
  NAND U24757 ( .A(n17454), .B(n17453), .Z(n17458) );
  AND U24758 ( .A(n17456), .B(n17455), .Z(n17457) );
  NAND U24759 ( .A(n17458), .B(n17457), .Z(n17459) );
  NANDN U24760 ( .A(n17460), .B(n17459), .Z(n17461) );
  OR U24761 ( .A(n17462), .B(n17461), .Z(n17463) );
  AND U24762 ( .A(n17464), .B(n17463), .Z(n17465) );
  NANDN U24763 ( .A(n17466), .B(n17465), .Z(n17467) );
  NAND U24764 ( .A(n17468), .B(n17467), .Z(n17469) );
  NANDN U24765 ( .A(n17470), .B(n17469), .Z(n17473) );
  AND U24766 ( .A(n17471), .B(n26565), .Z(n17472) );
  NAND U24767 ( .A(n17473), .B(n17472), .Z(n17474) );
  NANDN U24768 ( .A(n17475), .B(n17474), .Z(n17476) );
  OR U24769 ( .A(n17477), .B(n17476), .Z(n17478) );
  AND U24770 ( .A(n17479), .B(n17478), .Z(n17481) );
  NAND U24771 ( .A(n17481), .B(n17480), .Z(n17483) );
  ANDN U24772 ( .B(n17483), .A(n17482), .Z(n17484) );
  NANDN U24773 ( .A(n17485), .B(n17484), .Z(n17489) );
  AND U24774 ( .A(n17487), .B(n17486), .Z(n17488) );
  NAND U24775 ( .A(n17489), .B(n17488), .Z(n17490) );
  NANDN U24776 ( .A(n17491), .B(n17490), .Z(n17493) );
  OR U24777 ( .A(n17493), .B(n17492), .Z(n17494) );
  NAND U24778 ( .A(n17495), .B(n17494), .Z(n17496) );
  AND U24779 ( .A(n17497), .B(n17496), .Z(n17498) );
  OR U24780 ( .A(n24410), .B(n17498), .Z(n17499) );
  NAND U24781 ( .A(n17500), .B(n17499), .Z(n17501) );
  NANDN U24782 ( .A(n26576), .B(n17501), .Z(n17504) );
  AND U24783 ( .A(n17502), .B(n26579), .Z(n17503) );
  NAND U24784 ( .A(n17504), .B(n17503), .Z(n17505) );
  NANDN U24785 ( .A(n26580), .B(n17505), .Z(n17508) );
  AND U24786 ( .A(n17506), .B(n26581), .Z(n17507) );
  NAND U24787 ( .A(n17508), .B(n17507), .Z(n17509) );
  NANDN U24788 ( .A(n17510), .B(n17509), .Z(n17512) );
  IV U24789 ( .A(n17511), .Z(n26582) );
  OR U24790 ( .A(n17512), .B(n26582), .Z(n17513) );
  AND U24791 ( .A(n17514), .B(n17513), .Z(n17515) );
  NOR U24792 ( .A(n26585), .B(n17515), .Z(n17516) );
  NANDN U24793 ( .A(n17517), .B(n17516), .Z(n17520) );
  AND U24794 ( .A(n17519), .B(n17518), .Z(n26586) );
  AND U24795 ( .A(n17520), .B(n26586), .Z(n17523) );
  NANDN U24796 ( .A(n17523), .B(n26588), .Z(n17524) );
  NAND U24797 ( .A(n26589), .B(n17524), .Z(n17525) );
  NAND U24798 ( .A(n26590), .B(n17525), .Z(n17528) );
  AND U24799 ( .A(n17526), .B(n26591), .Z(n17527) );
  NAND U24800 ( .A(n17528), .B(n17527), .Z(n17529) );
  NANDN U24801 ( .A(n17530), .B(n17529), .Z(n17531) );
  OR U24802 ( .A(n17531), .B(n26592), .Z(n17532) );
  NAND U24803 ( .A(n17533), .B(n17532), .Z(n17537) );
  IV U24804 ( .A(n17534), .Z(n26595) );
  AND U24805 ( .A(n17535), .B(n26595), .Z(n17536) );
  NAND U24806 ( .A(n17537), .B(n17536), .Z(n17538) );
  NANDN U24807 ( .A(n17539), .B(n17538), .Z(n17541) );
  IV U24808 ( .A(n17540), .Z(n26596) );
  OR U24809 ( .A(n17541), .B(n26596), .Z(n17542) );
  AND U24810 ( .A(n26597), .B(n17542), .Z(n17545) );
  NAND U24811 ( .A(n26598), .B(n17543), .Z(n17544) );
  OR U24812 ( .A(n17545), .B(n17544), .Z(n17546) );
  AND U24813 ( .A(n26599), .B(n17546), .Z(n17547) );
  OR U24814 ( .A(n26602), .B(n17547), .Z(n17548) );
  NAND U24815 ( .A(n26603), .B(n17548), .Z(n17549) );
  NANDN U24816 ( .A(n17550), .B(n17549), .Z(n17553) );
  OR U24817 ( .A(n17553), .B(n26605), .Z(n17554) );
  NAND U24818 ( .A(n26606), .B(n17554), .Z(n17555) );
  NANDN U24819 ( .A(n17556), .B(n17555), .Z(n17557) );
  NAND U24820 ( .A(n26611), .B(n17557), .Z(n17558) );
  NANDN U24821 ( .A(n26613), .B(n17558), .Z(n17559) );
  AND U24822 ( .A(n26614), .B(n17559), .Z(n17560) );
  OR U24823 ( .A(n26617), .B(n17560), .Z(n17561) );
  AND U24824 ( .A(n26619), .B(n17561), .Z(n17562) );
  NOR U24825 ( .A(n17562), .B(n26621), .Z(n17563) );
  NANDN U24826 ( .A(n17564), .B(n17563), .Z(n17565) );
  AND U24827 ( .A(n17566), .B(n17565), .Z(n17567) );
  AND U24828 ( .A(n17567), .B(n26623), .Z(n17568) );
  OR U24829 ( .A(n17569), .B(n17568), .Z(n17570) );
  NAND U24830 ( .A(n17571), .B(n17570), .Z(n17572) );
  NANDN U24831 ( .A(n17573), .B(n17572), .Z(n17574) );
  NAND U24832 ( .A(n26635), .B(n17574), .Z(n17575) );
  ANDN U24833 ( .B(n17575), .A(n26637), .Z(n17576) );
  NANDN U24834 ( .A(n17577), .B(n17576), .Z(n17580) );
  AND U24835 ( .A(n17578), .B(n26639), .Z(n17579) );
  NAND U24836 ( .A(n17580), .B(n17579), .Z(n17581) );
  NANDN U24837 ( .A(n17582), .B(n17581), .Z(n17583) );
  OR U24838 ( .A(n26645), .B(n17583), .Z(n17584) );
  AND U24839 ( .A(n17585), .B(n17584), .Z(n17586) );
  NAND U24840 ( .A(n17586), .B(n26646), .Z(n17587) );
  NANDN U24841 ( .A(n26647), .B(n17587), .Z(n17588) );
  AND U24842 ( .A(n26648), .B(n17588), .Z(n17589) );
  OR U24843 ( .A(n26649), .B(n17589), .Z(n17590) );
  NAND U24844 ( .A(n26650), .B(n17590), .Z(n17591) );
  NANDN U24845 ( .A(n17592), .B(n17591), .Z(n17593) );
  OR U24846 ( .A(n26651), .B(n17593), .Z(n17594) );
  AND U24847 ( .A(n17595), .B(n17594), .Z(n17596) );
  NAND U24848 ( .A(n17596), .B(n26652), .Z(n17597) );
  AND U24849 ( .A(n26655), .B(n17597), .Z(n17598) );
  NANDN U24850 ( .A(n17599), .B(n17598), .Z(n17600) );
  NAND U24851 ( .A(n17601), .B(n17600), .Z(n17602) );
  NAND U24852 ( .A(n17603), .B(n17602), .Z(n17604) );
  NANDN U24853 ( .A(n26658), .B(n17604), .Z(n17607) );
  AND U24854 ( .A(n26659), .B(n17605), .Z(n17606) );
  NAND U24855 ( .A(n17607), .B(n17606), .Z(n17608) );
  NANDN U24856 ( .A(n26660), .B(n17608), .Z(n17611) );
  AND U24857 ( .A(n17609), .B(n26661), .Z(n17610) );
  NAND U24858 ( .A(n17611), .B(n17610), .Z(n17612) );
  NANDN U24859 ( .A(n26662), .B(n17612), .Z(n17614) );
  IV U24860 ( .A(n17613), .Z(n26664) );
  OR U24861 ( .A(n17614), .B(n26664), .Z(n17615) );
  NAND U24862 ( .A(n17616), .B(n17615), .Z(n17617) );
  NANDN U24863 ( .A(n26666), .B(n17617), .Z(n17620) );
  AND U24864 ( .A(n17618), .B(n26667), .Z(n17619) );
  NAND U24865 ( .A(n17620), .B(n17619), .Z(n17621) );
  NANDN U24866 ( .A(n17622), .B(n17621), .Z(n17625) );
  AND U24867 ( .A(n17623), .B(n26669), .Z(n17624) );
  NAND U24868 ( .A(n17625), .B(n17624), .Z(n17626) );
  NANDN U24869 ( .A(n26670), .B(n17626), .Z(n17629) );
  AND U24870 ( .A(n17627), .B(n26671), .Z(n17628) );
  NAND U24871 ( .A(n17629), .B(n17628), .Z(n17630) );
  NANDN U24872 ( .A(n17631), .B(n17630), .Z(n17632) );
  OR U24873 ( .A(n26672), .B(n17632), .Z(n17633) );
  AND U24874 ( .A(n17634), .B(n17633), .Z(n17636) );
  NAND U24875 ( .A(n17636), .B(n17635), .Z(n17638) );
  ANDN U24876 ( .B(n17638), .A(n17637), .Z(n17639) );
  NANDN U24877 ( .A(n26676), .B(n17639), .Z(n17642) );
  AND U24878 ( .A(n26677), .B(n17640), .Z(n17641) );
  NAND U24879 ( .A(n17642), .B(n17641), .Z(n17643) );
  NANDN U24880 ( .A(n26678), .B(n17643), .Z(n17644) );
  OR U24881 ( .A(n17645), .B(n17644), .Z(n17646) );
  AND U24882 ( .A(n17647), .B(n17646), .Z(n17648) );
  NANDN U24883 ( .A(n26679), .B(n17648), .Z(n17649) );
  AND U24884 ( .A(n17650), .B(n17649), .Z(n17652) );
  NAND U24885 ( .A(n17652), .B(n17651), .Z(n17654) );
  ANDN U24886 ( .B(n17654), .A(n17653), .Z(n17655) );
  NANDN U24887 ( .A(n17656), .B(n17655), .Z(n17657) );
  AND U24888 ( .A(n17658), .B(n17657), .Z(n17660) );
  OR U24889 ( .A(n17660), .B(n17659), .Z(n17663) );
  NANDN U24890 ( .A(x[1427]), .B(y[1427]), .Z(n17661) );
  AND U24891 ( .A(n17662), .B(n17661), .Z(n26684) );
  AND U24892 ( .A(n17663), .B(n26684), .Z(n17666) );
  NANDN U24893 ( .A(y[1427]), .B(x[1427]), .Z(n17664) );
  NAND U24894 ( .A(n17665), .B(n17664), .Z(n26685) );
  OR U24895 ( .A(n17666), .B(n26685), .Z(n17667) );
  NAND U24896 ( .A(n26686), .B(n17667), .Z(n17668) );
  NANDN U24897 ( .A(n26687), .B(n17668), .Z(n17669) );
  NAND U24898 ( .A(n26688), .B(n17669), .Z(n17670) );
  NANDN U24899 ( .A(n26689), .B(n17670), .Z(n17671) );
  AND U24900 ( .A(n26690), .B(n17671), .Z(n17672) );
  NANDN U24901 ( .A(n17672), .B(n26691), .Z(n17673) );
  NAND U24902 ( .A(n26692), .B(n17673), .Z(n17674) );
  NANDN U24903 ( .A(n26693), .B(n17674), .Z(n17675) );
  NAND U24904 ( .A(n26694), .B(n17675), .Z(n17676) );
  NANDN U24905 ( .A(n26696), .B(n17676), .Z(n17677) );
  AND U24906 ( .A(n26697), .B(n17677), .Z(n17678) );
  OR U24907 ( .A(n26698), .B(n17678), .Z(n17679) );
  NAND U24908 ( .A(n26699), .B(n17679), .Z(n17680) );
  NANDN U24909 ( .A(n17681), .B(n17680), .Z(n17683) );
  NAND U24910 ( .A(n17683), .B(n17682), .Z(n17685) );
  ANDN U24911 ( .B(n17685), .A(n17684), .Z(n17686) );
  NANDN U24912 ( .A(n17687), .B(n17686), .Z(n17688) );
  AND U24913 ( .A(n17689), .B(n17688), .Z(n17690) );
  NAND U24914 ( .A(n26703), .B(n17690), .Z(n17691) );
  NANDN U24915 ( .A(n26704), .B(n17691), .Z(n17692) );
  OR U24916 ( .A(n17693), .B(n17692), .Z(n17694) );
  AND U24917 ( .A(n26705), .B(n17694), .Z(n17695) );
  OR U24918 ( .A(n17695), .B(n26706), .Z(n17696) );
  AND U24919 ( .A(n26707), .B(n17696), .Z(n17697) );
  OR U24920 ( .A(n26708), .B(n17697), .Z(n17698) );
  NAND U24921 ( .A(n26709), .B(n17698), .Z(n17699) );
  NANDN U24922 ( .A(n26710), .B(n17699), .Z(n17700) );
  NAND U24923 ( .A(n26711), .B(n17700), .Z(n17701) );
  NANDN U24924 ( .A(n26712), .B(n17701), .Z(n17702) );
  AND U24925 ( .A(n17703), .B(n17702), .Z(n17704) );
  OR U24926 ( .A(n26714), .B(n17704), .Z(n17705) );
  AND U24927 ( .A(n17706), .B(n17705), .Z(n17707) );
  OR U24928 ( .A(n26717), .B(n17707), .Z(n17708) );
  NAND U24929 ( .A(n26718), .B(n17708), .Z(n17709) );
  NAND U24930 ( .A(n26719), .B(n17709), .Z(n17710) );
  NAND U24931 ( .A(n24403), .B(n17710), .Z(n17711) );
  AND U24932 ( .A(n17712), .B(n17711), .Z(n17716) );
  IV U24933 ( .A(n17713), .Z(n26722) );
  IV U24934 ( .A(n17714), .Z(n26721) );
  NAND U24935 ( .A(n26722), .B(n26721), .Z(n17715) );
  OR U24936 ( .A(n17716), .B(n17715), .Z(n17717) );
  AND U24937 ( .A(n17717), .B(n26723), .Z(n17719) );
  NAND U24938 ( .A(n17719), .B(n17718), .Z(n17720) );
  NANDN U24939 ( .A(n26724), .B(n17720), .Z(n17721) );
  AND U24940 ( .A(n17722), .B(n17721), .Z(n17723) );
  NAND U24941 ( .A(n17723), .B(n26725), .Z(n17725) );
  ANDN U24942 ( .B(n17725), .A(n17724), .Z(n17726) );
  NANDN U24943 ( .A(n26726), .B(n17726), .Z(n17730) );
  AND U24944 ( .A(n17728), .B(n17727), .Z(n17729) );
  NAND U24945 ( .A(n17730), .B(n17729), .Z(n17731) );
  NANDN U24946 ( .A(n17732), .B(n17731), .Z(n17733) );
  OR U24947 ( .A(n26730), .B(n17733), .Z(n17734) );
  AND U24948 ( .A(n26731), .B(n17734), .Z(n17736) );
  NAND U24949 ( .A(n17736), .B(n17735), .Z(n17737) );
  NAND U24950 ( .A(n26732), .B(n17737), .Z(n17738) );
  AND U24951 ( .A(n26733), .B(n17738), .Z(n17741) );
  OR U24952 ( .A(n17741), .B(n26734), .Z(n17742) );
  AND U24953 ( .A(n17743), .B(n17742), .Z(n17744) );
  NANDN U24954 ( .A(n26735), .B(n17744), .Z(n17745) );
  NAND U24955 ( .A(n17746), .B(n17745), .Z(n17749) );
  AND U24956 ( .A(n17747), .B(n26739), .Z(n17748) );
  NAND U24957 ( .A(n17749), .B(n17748), .Z(n17750) );
  NANDN U24958 ( .A(n26740), .B(n17750), .Z(n17753) );
  AND U24959 ( .A(n17751), .B(n26741), .Z(n17752) );
  NAND U24960 ( .A(n17753), .B(n17752), .Z(n17754) );
  NANDN U24961 ( .A(n17755), .B(n17754), .Z(n17756) );
  OR U24962 ( .A(n17756), .B(n24400), .Z(n17757) );
  AND U24963 ( .A(n26744), .B(n17757), .Z(n17758) );
  NANDN U24964 ( .A(n17759), .B(n17758), .Z(n17760) );
  NAND U24965 ( .A(n17761), .B(n17760), .Z(n17762) );
  NANDN U24966 ( .A(n26746), .B(n17762), .Z(n17763) );
  AND U24967 ( .A(n26747), .B(n17763), .Z(n17765) );
  IV U24968 ( .A(n17764), .Z(n26749) );
  OR U24969 ( .A(n17765), .B(n26749), .Z(n17766) );
  NAND U24970 ( .A(n26750), .B(n17766), .Z(n17767) );
  NANDN U24971 ( .A(n26751), .B(n17767), .Z(n17768) );
  NAND U24972 ( .A(n26752), .B(n17768), .Z(n17769) );
  NANDN U24973 ( .A(n26753), .B(n17769), .Z(n17770) );
  AND U24974 ( .A(n26754), .B(n17770), .Z(n17771) );
  NOR U24975 ( .A(n17771), .B(n26755), .Z(n17772) );
  NANDN U24976 ( .A(n17773), .B(n17772), .Z(n17774) );
  AND U24977 ( .A(n26756), .B(n17774), .Z(n17775) );
  NAND U24978 ( .A(n17775), .B(n26758), .Z(n17776) );
  NANDN U24979 ( .A(n17777), .B(n17776), .Z(n17780) );
  AND U24980 ( .A(n17779), .B(n17778), .Z(n24399) );
  AND U24981 ( .A(n17780), .B(n24399), .Z(n17781) );
  NOR U24982 ( .A(n26760), .B(n17781), .Z(n17782) );
  NAND U24983 ( .A(n17783), .B(n17782), .Z(n17784) );
  NAND U24984 ( .A(n17785), .B(n17784), .Z(n17786) );
  OR U24985 ( .A(n17787), .B(n17786), .Z(n17788) );
  AND U24986 ( .A(n17789), .B(n17788), .Z(n17790) );
  OR U24987 ( .A(n17791), .B(n17790), .Z(n17792) );
  NAND U24988 ( .A(n26763), .B(n17792), .Z(n17793) );
  NANDN U24989 ( .A(n26764), .B(n17793), .Z(n17794) );
  NAND U24990 ( .A(n26766), .B(n17794), .Z(n17795) );
  NANDN U24991 ( .A(n26767), .B(n17795), .Z(n17796) );
  AND U24992 ( .A(n17797), .B(n17796), .Z(n17800) );
  NANDN U24993 ( .A(n17800), .B(n26770), .Z(n17801) );
  AND U24994 ( .A(n17802), .B(n17801), .Z(n17803) );
  NAND U24995 ( .A(n26769), .B(n17803), .Z(n17804) );
  ANDN U24996 ( .B(n17804), .A(n24397), .Z(n17805) );
  NANDN U24997 ( .A(n26771), .B(n17805), .Z(n17808) );
  AND U24998 ( .A(n26772), .B(n17806), .Z(n17807) );
  NAND U24999 ( .A(n17808), .B(n17807), .Z(n17809) );
  NANDN U25000 ( .A(n26773), .B(n17809), .Z(n17812) );
  AND U25001 ( .A(n17810), .B(n26774), .Z(n17811) );
  NAND U25002 ( .A(n17812), .B(n17811), .Z(n17813) );
  NANDN U25003 ( .A(n26775), .B(n17813), .Z(n17815) );
  IV U25004 ( .A(n17814), .Z(n26776) );
  OR U25005 ( .A(n17815), .B(n26776), .Z(n17816) );
  NAND U25006 ( .A(n17817), .B(n17816), .Z(n17818) );
  NANDN U25007 ( .A(n26778), .B(n17818), .Z(n17819) );
  NAND U25008 ( .A(n26779), .B(n17819), .Z(n17820) );
  NANDN U25009 ( .A(n26781), .B(n17820), .Z(n17821) );
  AND U25010 ( .A(n26782), .B(n17821), .Z(n17824) );
  OR U25011 ( .A(n17824), .B(n26783), .Z(n17825) );
  AND U25012 ( .A(n17826), .B(n17825), .Z(n17827) );
  NAND U25013 ( .A(n17827), .B(n26784), .Z(n17829) );
  ANDN U25014 ( .B(n17829), .A(n17828), .Z(n17830) );
  NANDN U25015 ( .A(n26785), .B(n17830), .Z(n17834) );
  AND U25016 ( .A(n17832), .B(n17831), .Z(n17833) );
  NAND U25017 ( .A(n17834), .B(n17833), .Z(n17835) );
  NANDN U25018 ( .A(n17836), .B(n17835), .Z(n17838) );
  IV U25019 ( .A(n17837), .Z(n26788) );
  OR U25020 ( .A(n17838), .B(n26788), .Z(n17839) );
  AND U25021 ( .A(n26789), .B(n17839), .Z(n17840) );
  NANDN U25022 ( .A(n17841), .B(n17840), .Z(n17842) );
  NAND U25023 ( .A(n24393), .B(n17842), .Z(n17843) );
  NANDN U25024 ( .A(n17844), .B(n17843), .Z(n17845) );
  OR U25025 ( .A(n17845), .B(n26790), .Z(n17846) );
  NAND U25026 ( .A(n26791), .B(n17846), .Z(n17847) );
  NANDN U25027 ( .A(n17848), .B(n17847), .Z(n17849) );
  NAND U25028 ( .A(n26793), .B(n17849), .Z(n17850) );
  NANDN U25029 ( .A(n26794), .B(n17850), .Z(n17851) );
  AND U25030 ( .A(n26795), .B(n17851), .Z(n17852) );
  OR U25031 ( .A(n26797), .B(n17852), .Z(n17853) );
  NAND U25032 ( .A(n26798), .B(n17853), .Z(n17854) );
  NANDN U25033 ( .A(n26799), .B(n17854), .Z(n17855) );
  NAND U25034 ( .A(n26800), .B(n17855), .Z(n17856) );
  AND U25035 ( .A(n17857), .B(n17856), .Z(n17859) );
  IV U25036 ( .A(n17858), .Z(n26802) );
  OR U25037 ( .A(n17859), .B(n26802), .Z(n17860) );
  AND U25038 ( .A(n17861), .B(n17860), .Z(n17862) );
  NANDN U25039 ( .A(n26804), .B(n17862), .Z(n17865) );
  AND U25040 ( .A(n17864), .B(n17863), .Z(n24392) );
  AND U25041 ( .A(n17865), .B(n24392), .Z(n17868) );
  NAND U25042 ( .A(n26805), .B(n17866), .Z(n17867) );
  OR U25043 ( .A(n17868), .B(n17867), .Z(n17869) );
  AND U25044 ( .A(n17870), .B(n17869), .Z(n17871) );
  NAND U25045 ( .A(n26806), .B(n17871), .Z(n17873) );
  ANDN U25046 ( .B(n17873), .A(n17872), .Z(n17874) );
  NANDN U25047 ( .A(n17875), .B(n17874), .Z(n17878) );
  AND U25048 ( .A(n17876), .B(n24390), .Z(n17877) );
  NAND U25049 ( .A(n17878), .B(n17877), .Z(n17879) );
  NANDN U25050 ( .A(n17880), .B(n17879), .Z(n17881) );
  OR U25051 ( .A(n26810), .B(n17881), .Z(n17882) );
  AND U25052 ( .A(n26811), .B(n17882), .Z(n17885) );
  NANDN U25053 ( .A(n17885), .B(n26812), .Z(n17886) );
  AND U25054 ( .A(n26813), .B(n17886), .Z(n17889) );
  AND U25055 ( .A(n17887), .B(n24389), .Z(n17888) );
  NANDN U25056 ( .A(n17889), .B(n17888), .Z(n17890) );
  NANDN U25057 ( .A(n26814), .B(n17890), .Z(n17891) );
  AND U25058 ( .A(n26815), .B(n17891), .Z(n17894) );
  NANDN U25059 ( .A(n17894), .B(n26816), .Z(n17895) );
  NAND U25060 ( .A(n17896), .B(n17895), .Z(n17897) );
  NANDN U25061 ( .A(n17898), .B(n17897), .Z(n17901) );
  AND U25062 ( .A(n17899), .B(n26820), .Z(n17900) );
  NAND U25063 ( .A(n17901), .B(n17900), .Z(n17902) );
  NAND U25064 ( .A(n26821), .B(n17902), .Z(n17904) );
  AND U25065 ( .A(n24385), .B(n24386), .Z(n17903) );
  NAND U25066 ( .A(n17904), .B(n17903), .Z(n17905) );
  NANDN U25067 ( .A(n17906), .B(n17905), .Z(n17907) );
  NAND U25068 ( .A(n26825), .B(n17907), .Z(n17908) );
  NAND U25069 ( .A(n26826), .B(n17908), .Z(n17909) );
  AND U25070 ( .A(n17909), .B(n24384), .Z(n17910) );
  OR U25071 ( .A(n17911), .B(n17910), .Z(n17912) );
  NAND U25072 ( .A(n17913), .B(n17912), .Z(n17914) );
  NANDN U25073 ( .A(n17915), .B(n17914), .Z(n17916) );
  OR U25074 ( .A(n17917), .B(n17916), .Z(n17918) );
  AND U25075 ( .A(n17919), .B(n17918), .Z(n17921) );
  NAND U25076 ( .A(n17921), .B(n17920), .Z(n17923) );
  ANDN U25077 ( .B(n17923), .A(n17922), .Z(n17924) );
  NANDN U25078 ( .A(n26831), .B(n17924), .Z(n17927) );
  AND U25079 ( .A(n26832), .B(n17925), .Z(n17926) );
  NAND U25080 ( .A(n17927), .B(n17926), .Z(n17928) );
  NANDN U25081 ( .A(n26833), .B(n17928), .Z(n17930) );
  NAND U25082 ( .A(n17930), .B(n17929), .Z(n17931) );
  NAND U25083 ( .A(n26834), .B(n17931), .Z(n17932) );
  AND U25084 ( .A(n26835), .B(n17932), .Z(n17934) );
  NAND U25085 ( .A(n17934), .B(n17933), .Z(n17935) );
  NANDN U25086 ( .A(n26838), .B(n17935), .Z(n17936) );
  AND U25087 ( .A(n26839), .B(n17936), .Z(n17937) );
  OR U25088 ( .A(n17937), .B(n26840), .Z(n17938) );
  AND U25089 ( .A(n26841), .B(n17938), .Z(n17939) );
  NANDN U25090 ( .A(n17939), .B(n26842), .Z(n17940) );
  NANDN U25091 ( .A(n24383), .B(n17940), .Z(n17941) );
  AND U25092 ( .A(n26843), .B(n17941), .Z(n17942) );
  OR U25093 ( .A(n26845), .B(n17942), .Z(n17943) );
  AND U25094 ( .A(n26846), .B(n17943), .Z(n17945) );
  NANDN U25095 ( .A(n17945), .B(n17944), .Z(n17946) );
  AND U25096 ( .A(n26847), .B(n17946), .Z(n17947) );
  NOR U25097 ( .A(n26848), .B(n17947), .Z(n17948) );
  NANDN U25098 ( .A(n17949), .B(n17948), .Z(n17951) );
  IV U25099 ( .A(n17950), .Z(n26849) );
  AND U25100 ( .A(n17951), .B(n26849), .Z(n17952) );
  OR U25101 ( .A(n17953), .B(n17952), .Z(n17954) );
  AND U25102 ( .A(n26851), .B(n17954), .Z(n17955) );
  OR U25103 ( .A(n26852), .B(n17955), .Z(n17956) );
  NAND U25104 ( .A(n26854), .B(n17956), .Z(n17957) );
  NANDN U25105 ( .A(n26855), .B(n17957), .Z(n17961) );
  NAND U25106 ( .A(n17961), .B(n26856), .Z(n17962) );
  AND U25107 ( .A(n26857), .B(n17962), .Z(n17963) );
  OR U25108 ( .A(n26858), .B(n17963), .Z(n17964) );
  AND U25109 ( .A(n26859), .B(n17964), .Z(n17968) );
  NANDN U25110 ( .A(n17968), .B(n26860), .Z(n17969) );
  NAND U25111 ( .A(n26861), .B(n17969), .Z(n17970) );
  NAND U25112 ( .A(n26862), .B(n17970), .Z(n17973) );
  AND U25113 ( .A(n17971), .B(n26863), .Z(n17972) );
  NAND U25114 ( .A(n17973), .B(n17972), .Z(n17974) );
  NANDN U25115 ( .A(n24381), .B(n17974), .Z(n17975) );
  OR U25116 ( .A(n17975), .B(n26865), .Z(n17976) );
  NAND U25117 ( .A(n17977), .B(n17976), .Z(n17978) );
  NAND U25118 ( .A(n26867), .B(n17978), .Z(n17979) );
  ANDN U25119 ( .B(n17979), .A(n26868), .Z(n17980) );
  NANDN U25120 ( .A(n17981), .B(n17980), .Z(n17983) );
  AND U25121 ( .A(n26869), .B(n26872), .Z(n17982) );
  NAND U25122 ( .A(n17983), .B(n17982), .Z(n17984) );
  NANDN U25123 ( .A(n17985), .B(n17984), .Z(n17986) );
  OR U25124 ( .A(n17986), .B(n26873), .Z(n17987) );
  NAND U25125 ( .A(n26874), .B(n17987), .Z(n17988) );
  AND U25126 ( .A(n17989), .B(n17988), .Z(n17990) );
  NAND U25127 ( .A(n17990), .B(n26875), .Z(n17992) );
  ANDN U25128 ( .B(n17992), .A(n17991), .Z(n17993) );
  NANDN U25129 ( .A(n26876), .B(n17993), .Z(n17996) );
  AND U25130 ( .A(n17994), .B(n24378), .Z(n17995) );
  NAND U25131 ( .A(n17996), .B(n17995), .Z(n17997) );
  NANDN U25132 ( .A(n17998), .B(n17997), .Z(n17999) );
  OR U25133 ( .A(n26877), .B(n17999), .Z(n18000) );
  AND U25134 ( .A(n26878), .B(n18000), .Z(n18003) );
  NAND U25135 ( .A(n18002), .B(n18001), .Z(n24377) );
  OR U25136 ( .A(n18003), .B(n24377), .Z(n18004) );
  NAND U25137 ( .A(n26879), .B(n18004), .Z(n18005) );
  NAND U25138 ( .A(n26880), .B(n18005), .Z(n18008) );
  AND U25139 ( .A(n18006), .B(n24376), .Z(n18007) );
  NAND U25140 ( .A(n18008), .B(n18007), .Z(n18009) );
  NANDN U25141 ( .A(n18010), .B(n18009), .Z(n18011) );
  OR U25142 ( .A(n18011), .B(n26881), .Z(n18012) );
  NAND U25143 ( .A(n18013), .B(n18012), .Z(n18014) );
  NANDN U25144 ( .A(n18015), .B(n18014), .Z(n18016) );
  NANDN U25145 ( .A(n18017), .B(n18016), .Z(n18022) );
  OR U25146 ( .A(n18019), .B(n18018), .Z(n18020) );
  AND U25147 ( .A(n18021), .B(n18020), .Z(n26889) );
  ANDN U25148 ( .B(n18022), .A(n26889), .Z(n18023) );
  OR U25149 ( .A(n18024), .B(n18023), .Z(n18025) );
  AND U25150 ( .A(n18026), .B(n18025), .Z(n18027) );
  NAND U25151 ( .A(n18027), .B(n26888), .Z(n18029) );
  ANDN U25152 ( .B(n18029), .A(n18028), .Z(n18030) );
  NANDN U25153 ( .A(n18031), .B(n18030), .Z(n18035) );
  AND U25154 ( .A(n18033), .B(n18032), .Z(n18034) );
  NAND U25155 ( .A(n18035), .B(n18034), .Z(n18036) );
  NANDN U25156 ( .A(n18037), .B(n18036), .Z(n18038) );
  OR U25157 ( .A(n18039), .B(n18038), .Z(n18040) );
  AND U25158 ( .A(n18041), .B(n18040), .Z(n18042) );
  NANDN U25159 ( .A(n26895), .B(n18042), .Z(n18043) );
  NAND U25160 ( .A(n18044), .B(n18043), .Z(n18045) );
  NANDN U25161 ( .A(n26897), .B(n18045), .Z(n18048) );
  AND U25162 ( .A(n18046), .B(n26898), .Z(n18047) );
  NAND U25163 ( .A(n18048), .B(n18047), .Z(n18049) );
  NANDN U25164 ( .A(n18050), .B(n18049), .Z(n18051) );
  OR U25165 ( .A(n26899), .B(n18051), .Z(n18052) );
  AND U25166 ( .A(n18053), .B(n18052), .Z(n18054) );
  OR U25167 ( .A(n18055), .B(n18054), .Z(n18056) );
  NAND U25168 ( .A(n18057), .B(n18056), .Z(n18058) );
  NANDN U25169 ( .A(n18059), .B(n18058), .Z(n18062) );
  AND U25170 ( .A(n18060), .B(n24372), .Z(n18061) );
  NAND U25171 ( .A(n18062), .B(n18061), .Z(n18063) );
  NANDN U25172 ( .A(n18064), .B(n18063), .Z(n18065) );
  OR U25173 ( .A(n18065), .B(n24371), .Z(n18068) );
  AND U25174 ( .A(n18067), .B(n18066), .Z(n24370) );
  AND U25175 ( .A(n18068), .B(n24370), .Z(n18071) );
  NANDN U25176 ( .A(n18071), .B(n26904), .Z(n18072) );
  AND U25177 ( .A(n18073), .B(n18072), .Z(n18074) );
  NOR U25178 ( .A(n18074), .B(n26908), .Z(n18075) );
  NANDN U25179 ( .A(n26906), .B(n18075), .Z(n18076) );
  AND U25180 ( .A(n18077), .B(n18076), .Z(n18078) );
  NAND U25181 ( .A(n18078), .B(n26909), .Z(n18079) );
  NANDN U25182 ( .A(n26910), .B(n18079), .Z(n18080) );
  AND U25183 ( .A(n26911), .B(n18080), .Z(n18083) );
  NAND U25184 ( .A(n18082), .B(n18081), .Z(n24369) );
  OR U25185 ( .A(n18083), .B(n24369), .Z(n18084) );
  NAND U25186 ( .A(n26913), .B(n18084), .Z(n18085) );
  NAND U25187 ( .A(n26914), .B(n18085), .Z(n18086) );
  NAND U25188 ( .A(n26915), .B(n18086), .Z(n18087) );
  NAND U25189 ( .A(n26916), .B(n18087), .Z(n18088) );
  AND U25190 ( .A(n18089), .B(n18088), .Z(n18090) );
  NAND U25191 ( .A(n18090), .B(n26917), .Z(n18091) );
  ANDN U25192 ( .B(n18091), .A(n26918), .Z(n18092) );
  NANDN U25193 ( .A(n26920), .B(n18092), .Z(n18095) );
  AND U25194 ( .A(n18093), .B(n24368), .Z(n18094) );
  NAND U25195 ( .A(n18095), .B(n18094), .Z(n18096) );
  NAND U25196 ( .A(n26921), .B(n18096), .Z(n18097) );
  NANDN U25197 ( .A(n26922), .B(n18097), .Z(n18098) );
  AND U25198 ( .A(n26923), .B(n18098), .Z(n18099) );
  OR U25199 ( .A(n26924), .B(n18099), .Z(n18100) );
  NAND U25200 ( .A(n26925), .B(n18100), .Z(n18101) );
  NANDN U25201 ( .A(n18102), .B(n18101), .Z(n18104) );
  IV U25202 ( .A(n18103), .Z(n26926) );
  OR U25203 ( .A(n18104), .B(n26926), .Z(n18105) );
  AND U25204 ( .A(n26927), .B(n18105), .Z(n18106) );
  ANDN U25205 ( .B(n18107), .A(n18106), .Z(n18108) );
  NAND U25206 ( .A(n18109), .B(n18108), .Z(n18110) );
  NANDN U25207 ( .A(n18111), .B(n18110), .Z(n18112) );
  OR U25208 ( .A(n26930), .B(n18112), .Z(n18113) );
  AND U25209 ( .A(n18114), .B(n18113), .Z(n18115) );
  NANDN U25210 ( .A(n26933), .B(n18115), .Z(n18116) );
  AND U25211 ( .A(n18117), .B(n18116), .Z(n18118) );
  OR U25212 ( .A(n26935), .B(n18118), .Z(n18119) );
  NAND U25213 ( .A(n26936), .B(n18119), .Z(n18120) );
  NANDN U25214 ( .A(n26937), .B(n18120), .Z(n18121) );
  NAND U25215 ( .A(n26938), .B(n18121), .Z(n18122) );
  NAND U25216 ( .A(n24367), .B(n18122), .Z(n18123) );
  NANDN U25217 ( .A(n26939), .B(n18123), .Z(n18124) );
  AND U25218 ( .A(n18124), .B(n26940), .Z(n18125) );
  OR U25219 ( .A(n18125), .B(n26941), .Z(n18126) );
  NAND U25220 ( .A(n18127), .B(n18126), .Z(n18128) );
  NANDN U25221 ( .A(n18129), .B(n18128), .Z(n18130) );
  NAND U25222 ( .A(n18131), .B(n18130), .Z(n18132) );
  NANDN U25223 ( .A(n26947), .B(n18132), .Z(n18133) );
  AND U25224 ( .A(n26948), .B(n18133), .Z(n18134) );
  OR U25225 ( .A(n26949), .B(n18134), .Z(n18135) );
  NAND U25226 ( .A(n26950), .B(n18135), .Z(n18136) );
  NANDN U25227 ( .A(n26951), .B(n18136), .Z(n18140) );
  IV U25228 ( .A(n18137), .Z(n26952) );
  ANDN U25229 ( .B(n26952), .A(n18138), .Z(n18139) );
  NAND U25230 ( .A(n18140), .B(n18139), .Z(n18141) );
  AND U25231 ( .A(n18141), .B(n26953), .Z(n18147) );
  OR U25232 ( .A(n18143), .B(n18142), .Z(n18144) );
  AND U25233 ( .A(n18145), .B(n18144), .Z(n18146) );
  NANDN U25234 ( .A(n18147), .B(n18146), .Z(n18148) );
  NANDN U25235 ( .A(n26954), .B(n18148), .Z(n18150) );
  IV U25236 ( .A(n18149), .Z(n26955) );
  AND U25237 ( .A(n18150), .B(n26955), .Z(n18151) );
  OR U25238 ( .A(n26956), .B(n18151), .Z(n18152) );
  NAND U25239 ( .A(n26957), .B(n18152), .Z(n18153) );
  NANDN U25240 ( .A(n26958), .B(n18153), .Z(n18154) );
  NAND U25241 ( .A(n26961), .B(n18154), .Z(n18155) );
  NANDN U25242 ( .A(n26962), .B(n18155), .Z(n18156) );
  AND U25243 ( .A(n18157), .B(n18156), .Z(n18159) );
  OR U25244 ( .A(n18159), .B(n18158), .Z(n18160) );
  AND U25245 ( .A(n26964), .B(n18160), .Z(n18162) );
  IV U25246 ( .A(n18161), .Z(n26966) );
  OR U25247 ( .A(n18162), .B(n26966), .Z(n18163) );
  NAND U25248 ( .A(n26967), .B(n18163), .Z(n18164) );
  NANDN U25249 ( .A(n18165), .B(n18164), .Z(n18166) );
  NANDN U25250 ( .A(n18166), .B(n26968), .Z(n18167) );
  NAND U25251 ( .A(n26969), .B(n18167), .Z(n18168) );
  NANDN U25252 ( .A(n18169), .B(n18168), .Z(n18170) );
  NANDN U25253 ( .A(n26971), .B(n18170), .Z(n18171) );
  AND U25254 ( .A(n26972), .B(n18171), .Z(n18172) );
  OR U25255 ( .A(n26973), .B(n18172), .Z(n18173) );
  NAND U25256 ( .A(n26974), .B(n18173), .Z(n18174) );
  NANDN U25257 ( .A(n26975), .B(n18174), .Z(n18175) );
  NAND U25258 ( .A(n26977), .B(n18175), .Z(n18176) );
  ANDN U25259 ( .B(n18176), .A(n24363), .Z(n18177) );
  NANDN U25260 ( .A(n18178), .B(n18177), .Z(n18179) );
  NAND U25261 ( .A(n24362), .B(n18179), .Z(n18180) );
  NAND U25262 ( .A(n18181), .B(n18180), .Z(n18182) );
  NANDN U25263 ( .A(y[1711]), .B(n18182), .Z(n18185) );
  XNOR U25264 ( .A(y[1711]), .B(n18182), .Z(n18183) );
  NAND U25265 ( .A(n18183), .B(x[1711]), .Z(n18184) );
  NAND U25266 ( .A(n18185), .B(n18184), .Z(n18186) );
  AND U25267 ( .A(n18187), .B(n18186), .Z(n18189) );
  IV U25268 ( .A(n18188), .Z(n26978) );
  NANDN U25269 ( .A(n18189), .B(n26978), .Z(n18190) );
  NANDN U25270 ( .A(n26979), .B(n18190), .Z(n18192) );
  IV U25271 ( .A(n18191), .Z(n26980) );
  AND U25272 ( .A(n18192), .B(n26980), .Z(n18194) );
  IV U25273 ( .A(n18193), .Z(n26981) );
  OR U25274 ( .A(n18194), .B(n26981), .Z(n18196) );
  IV U25275 ( .A(n18195), .Z(n26982) );
  AND U25276 ( .A(n18196), .B(n26982), .Z(n18198) );
  IV U25277 ( .A(n18197), .Z(n26983) );
  OR U25278 ( .A(n18198), .B(n26983), .Z(n18199) );
  AND U25279 ( .A(n26984), .B(n18199), .Z(n18200) );
  OR U25280 ( .A(n26985), .B(n18200), .Z(n18201) );
  NAND U25281 ( .A(n26986), .B(n18201), .Z(n18202) );
  NANDN U25282 ( .A(n18203), .B(n18202), .Z(n18204) );
  OR U25283 ( .A(n18204), .B(n26987), .Z(n18205) );
  NAND U25284 ( .A(n18206), .B(n18205), .Z(n18207) );
  NANDN U25285 ( .A(n18208), .B(n18207), .Z(n18209) );
  OR U25286 ( .A(n18210), .B(n18209), .Z(n18211) );
  AND U25287 ( .A(n18212), .B(n18211), .Z(n18213) );
  NANDN U25288 ( .A(n26993), .B(n18213), .Z(n18214) );
  AND U25289 ( .A(n18215), .B(n18214), .Z(n18218) );
  NAND U25290 ( .A(n18217), .B(n18216), .Z(n24359) );
  OR U25291 ( .A(n18218), .B(n24359), .Z(n18219) );
  NAND U25292 ( .A(n26995), .B(n18219), .Z(n18220) );
  NAND U25293 ( .A(n26996), .B(n18220), .Z(n18221) );
  NAND U25294 ( .A(n26997), .B(n18221), .Z(n18222) );
  AND U25295 ( .A(n18223), .B(n18222), .Z(n18224) );
  OR U25296 ( .A(n18225), .B(n18224), .Z(n18226) );
  NAND U25297 ( .A(n18227), .B(n18226), .Z(n18228) );
  NANDN U25298 ( .A(n18229), .B(n18228), .Z(n18232) );
  AND U25299 ( .A(n18230), .B(n27004), .Z(n18231) );
  NAND U25300 ( .A(n18232), .B(n18231), .Z(n18233) );
  NANDN U25301 ( .A(n18234), .B(n18233), .Z(n18235) );
  OR U25302 ( .A(n27005), .B(n18235), .Z(n18236) );
  AND U25303 ( .A(n27006), .B(n18236), .Z(n18239) );
  NANDN U25304 ( .A(n18239), .B(n27008), .Z(n18240) );
  NAND U25305 ( .A(n18241), .B(n18240), .Z(n18243) );
  OR U25306 ( .A(n18243), .B(n18242), .Z(n18246) );
  NANDN U25307 ( .A(x[1738]), .B(y[1738]), .Z(n18245) );
  AND U25308 ( .A(n18245), .B(n18244), .Z(n24358) );
  AND U25309 ( .A(n18246), .B(n24358), .Z(n18249) );
  NANDN U25310 ( .A(n18249), .B(n27011), .Z(n18250) );
  NAND U25311 ( .A(n27012), .B(n18250), .Z(n18251) );
  NAND U25312 ( .A(n27013), .B(n18251), .Z(n18254) );
  AND U25313 ( .A(n18252), .B(n24357), .Z(n18253) );
  NAND U25314 ( .A(n18254), .B(n18253), .Z(n18255) );
  NANDN U25315 ( .A(n18256), .B(n18255), .Z(n18257) );
  OR U25316 ( .A(n18257), .B(n24356), .Z(n18258) );
  AND U25317 ( .A(n18259), .B(n18258), .Z(n18260) );
  OR U25318 ( .A(n18261), .B(n18260), .Z(n18262) );
  NAND U25319 ( .A(n27018), .B(n18262), .Z(n18263) );
  NANDN U25320 ( .A(n27019), .B(n18263), .Z(n18264) );
  NAND U25321 ( .A(n24355), .B(n18264), .Z(n18265) );
  NANDN U25322 ( .A(n27022), .B(n18265), .Z(n18266) );
  AND U25323 ( .A(n18266), .B(n27023), .Z(n18267) );
  OR U25324 ( .A(n18267), .B(n27024), .Z(n18268) );
  NAND U25325 ( .A(n18269), .B(n18268), .Z(n18270) );
  NANDN U25326 ( .A(n18271), .B(n18270), .Z(n18274) );
  AND U25327 ( .A(n18272), .B(n27027), .Z(n18273) );
  NAND U25328 ( .A(n18274), .B(n18273), .Z(n18275) );
  NANDN U25329 ( .A(n27031), .B(n18275), .Z(n18276) );
  OR U25330 ( .A(n18277), .B(n18276), .Z(n18278) );
  AND U25331 ( .A(n18279), .B(n18278), .Z(n18280) );
  NANDN U25332 ( .A(n27032), .B(n18280), .Z(n18281) );
  AND U25333 ( .A(n27033), .B(n18281), .Z(n18284) );
  NANDN U25334 ( .A(n18284), .B(n27034), .Z(n18285) );
  NAND U25335 ( .A(n24354), .B(n18285), .Z(n18286) );
  NAND U25336 ( .A(n27035), .B(n18286), .Z(n18289) );
  AND U25337 ( .A(n18288), .B(n18287), .Z(n27037) );
  AND U25338 ( .A(n18289), .B(n27037), .Z(n18292) );
  NANDN U25339 ( .A(n18292), .B(n27039), .Z(n18293) );
  NAND U25340 ( .A(n24353), .B(n18293), .Z(n18294) );
  NANDN U25341 ( .A(n18295), .B(n18294), .Z(n18296) );
  OR U25342 ( .A(n27040), .B(n18296), .Z(n18297) );
  AND U25343 ( .A(n18298), .B(n18297), .Z(n18299) );
  NAND U25344 ( .A(n18299), .B(n27041), .Z(n18301) );
  ANDN U25345 ( .B(n18301), .A(n18300), .Z(n18302) );
  NANDN U25346 ( .A(n27044), .B(n18302), .Z(n18303) );
  NAND U25347 ( .A(n18304), .B(n18303), .Z(n18305) );
  NANDN U25348 ( .A(n27046), .B(n18305), .Z(n18306) );
  AND U25349 ( .A(n27047), .B(n18306), .Z(n18307) );
  OR U25350 ( .A(n27048), .B(n18307), .Z(n18308) );
  NAND U25351 ( .A(n27049), .B(n18308), .Z(n18309) );
  NANDN U25352 ( .A(n27050), .B(n18309), .Z(n18313) );
  IV U25353 ( .A(n18310), .Z(n27051) );
  AND U25354 ( .A(n18311), .B(n27051), .Z(n18312) );
  NAND U25355 ( .A(n18313), .B(n18312), .Z(n18314) );
  NANDN U25356 ( .A(n27052), .B(n18314), .Z(n18315) );
  NAND U25357 ( .A(n18316), .B(n18315), .Z(n18318) );
  AND U25358 ( .A(n18318), .B(n18317), .Z(n18320) );
  NANDN U25359 ( .A(n18320), .B(n18319), .Z(n18321) );
  NAND U25360 ( .A(n18322), .B(n18321), .Z(n18323) );
  NANDN U25361 ( .A(n18324), .B(n18323), .Z(n18325) );
  AND U25362 ( .A(n18325), .B(n24350), .Z(n18327) );
  NAND U25363 ( .A(n18327), .B(n18326), .Z(n18328) );
  NAND U25364 ( .A(n27058), .B(n18328), .Z(n18331) );
  AND U25365 ( .A(n18330), .B(n18329), .Z(n27059) );
  AND U25366 ( .A(n18331), .B(n27059), .Z(n18334) );
  NAND U25367 ( .A(n18333), .B(n18332), .Z(n24349) );
  OR U25368 ( .A(n18334), .B(n24349), .Z(n18337) );
  AND U25369 ( .A(n18336), .B(n18335), .Z(n24348) );
  AND U25370 ( .A(n18337), .B(n24348), .Z(n18338) );
  OR U25371 ( .A(n27060), .B(n18338), .Z(n18339) );
  NAND U25372 ( .A(n27061), .B(n18339), .Z(n18340) );
  NANDN U25373 ( .A(n27062), .B(n18340), .Z(n18341) );
  NAND U25374 ( .A(n27063), .B(n18341), .Z(n18342) );
  AND U25375 ( .A(n18343), .B(n18342), .Z(n18345) );
  NAND U25376 ( .A(n27068), .B(n27066), .Z(n18344) );
  OR U25377 ( .A(n18345), .B(n18344), .Z(n18346) );
  AND U25378 ( .A(n27069), .B(n18346), .Z(n18347) );
  NANDN U25379 ( .A(n18348), .B(n18347), .Z(n18349) );
  AND U25380 ( .A(n27070), .B(n18349), .Z(n18350) );
  OR U25381 ( .A(n27071), .B(n18350), .Z(n18351) );
  NAND U25382 ( .A(n27072), .B(n18351), .Z(n18352) );
  NANDN U25383 ( .A(n27073), .B(n18352), .Z(n18353) );
  AND U25384 ( .A(n27074), .B(n18353), .Z(n18354) );
  OR U25385 ( .A(n27075), .B(n18354), .Z(n18355) );
  NAND U25386 ( .A(n24347), .B(n18355), .Z(n18356) );
  NANDN U25387 ( .A(n27077), .B(n18356), .Z(n18357) );
  AND U25388 ( .A(n27078), .B(n18357), .Z(n18358) );
  OR U25389 ( .A(n18359), .B(n18358), .Z(n18360) );
  NAND U25390 ( .A(n27079), .B(n18360), .Z(n18361) );
  NANDN U25391 ( .A(n27080), .B(n18361), .Z(n18362) );
  AND U25392 ( .A(n27081), .B(n18362), .Z(n18363) );
  OR U25393 ( .A(n27083), .B(n18363), .Z(n18364) );
  NANDN U25394 ( .A(n27084), .B(n18364), .Z(n18365) );
  AND U25395 ( .A(n27086), .B(n18365), .Z(n18368) );
  NANDN U25396 ( .A(n18368), .B(n27087), .Z(n18369) );
  NAND U25397 ( .A(n24345), .B(n18369), .Z(n18370) );
  NANDN U25398 ( .A(n27088), .B(n18370), .Z(n18371) );
  NAND U25399 ( .A(n27089), .B(n18371), .Z(n18373) );
  IV U25400 ( .A(n18372), .Z(n27090) );
  ANDN U25401 ( .B(n18373), .A(n27090), .Z(n18374) );
  NANDN U25402 ( .A(n18375), .B(n18374), .Z(n18379) );
  IV U25403 ( .A(n18376), .Z(n27091) );
  AND U25404 ( .A(n18377), .B(n27091), .Z(n18378) );
  NAND U25405 ( .A(n18379), .B(n18378), .Z(n18380) );
  NANDN U25406 ( .A(n18381), .B(n18380), .Z(n18383) );
  IV U25407 ( .A(n18382), .Z(n27094) );
  OR U25408 ( .A(n18383), .B(n27094), .Z(n18384) );
  AND U25409 ( .A(n18385), .B(n18384), .Z(n18386) );
  NANDN U25410 ( .A(n27095), .B(n18386), .Z(n18389) );
  AND U25411 ( .A(n18388), .B(n18387), .Z(n27096) );
  AND U25412 ( .A(n18389), .B(n27096), .Z(n18392) );
  NANDN U25413 ( .A(n18392), .B(n27097), .Z(n18393) );
  NAND U25414 ( .A(n27098), .B(n18393), .Z(n18394) );
  NAND U25415 ( .A(n27100), .B(n18394), .Z(n18395) );
  NAND U25416 ( .A(n24344), .B(n18395), .Z(n18396) );
  NAND U25417 ( .A(n27101), .B(n18396), .Z(n18397) );
  NANDN U25418 ( .A(n24343), .B(n18397), .Z(n18398) );
  AND U25419 ( .A(n18398), .B(n24342), .Z(n18399) );
  OR U25420 ( .A(n18399), .B(n27102), .Z(n18400) );
  NAND U25421 ( .A(n27103), .B(n18400), .Z(n18401) );
  NANDN U25422 ( .A(n18402), .B(n18401), .Z(n18403) );
  NAND U25423 ( .A(n18403), .B(n27105), .Z(n18405) );
  ANDN U25424 ( .B(n18405), .A(n18404), .Z(n18406) );
  NANDN U25425 ( .A(n27106), .B(n18406), .Z(n18407) );
  NAND U25426 ( .A(n27107), .B(n18407), .Z(n18408) );
  AND U25427 ( .A(n27108), .B(n18408), .Z(n18411) );
  NAND U25428 ( .A(n18410), .B(n18409), .Z(n27109) );
  OR U25429 ( .A(n18411), .B(n27109), .Z(n18412) );
  NAND U25430 ( .A(n27110), .B(n18412), .Z(n18413) );
  NANDN U25431 ( .A(n24341), .B(n18413), .Z(n18414) );
  NANDN U25432 ( .A(n27113), .B(n18414), .Z(n18415) );
  AND U25433 ( .A(n27114), .B(n18415), .Z(n18416) );
  ANDN U25434 ( .B(n18417), .A(n18416), .Z(n18418) );
  NAND U25435 ( .A(n27115), .B(n18418), .Z(n18419) );
  NANDN U25436 ( .A(n27116), .B(n18419), .Z(n18420) );
  OR U25437 ( .A(n18421), .B(n18420), .Z(n18422) );
  AND U25438 ( .A(n18423), .B(n18422), .Z(n18424) );
  NANDN U25439 ( .A(n27119), .B(n18424), .Z(n18425) );
  AND U25440 ( .A(n18426), .B(n18425), .Z(n18427) );
  OR U25441 ( .A(n27121), .B(n18427), .Z(n18428) );
  NAND U25442 ( .A(n27122), .B(n18428), .Z(n18429) );
  NANDN U25443 ( .A(n27123), .B(n18429), .Z(n18430) );
  NAND U25444 ( .A(n24340), .B(n18430), .Z(n18431) );
  NAND U25445 ( .A(n27124), .B(n18431), .Z(n18432) );
  NANDN U25446 ( .A(n18433), .B(n18432), .Z(n18437) );
  IV U25447 ( .A(n18434), .Z(n27126) );
  OR U25448 ( .A(n18435), .B(n27126), .Z(n18436) );
  AND U25449 ( .A(n18437), .B(n18436), .Z(n18438) );
  OR U25450 ( .A(n18439), .B(n18438), .Z(n18440) );
  AND U25451 ( .A(n18441), .B(n18440), .Z(n18442) );
  NOR U25452 ( .A(n18442), .B(n27135), .Z(n18443) );
  NANDN U25453 ( .A(n18444), .B(n18443), .Z(n18445) );
  AND U25454 ( .A(n27136), .B(n18445), .Z(n18447) );
  NAND U25455 ( .A(n18447), .B(n18446), .Z(n18448) );
  NANDN U25456 ( .A(n27139), .B(n18448), .Z(n18449) );
  AND U25457 ( .A(n27141), .B(n18449), .Z(n18452) );
  NAND U25458 ( .A(n18451), .B(n18450), .Z(n27143) );
  OR U25459 ( .A(n18452), .B(n27143), .Z(n18453) );
  AND U25460 ( .A(n27145), .B(n18453), .Z(n18454) );
  OR U25461 ( .A(n27147), .B(n18454), .Z(n18455) );
  NAND U25462 ( .A(n27149), .B(n18455), .Z(n18456) );
  NAND U25463 ( .A(n27150), .B(n18456), .Z(n18459) );
  AND U25464 ( .A(n18457), .B(n27152), .Z(n18458) );
  NAND U25465 ( .A(n18459), .B(n18458), .Z(n18460) );
  NANDN U25466 ( .A(n18461), .B(n18460), .Z(n18462) );
  OR U25467 ( .A(n18462), .B(n27154), .Z(n18463) );
  NANDN U25468 ( .A(n18464), .B(n18463), .Z(n18465) );
  AND U25469 ( .A(n18466), .B(n18465), .Z(n18467) );
  OR U25470 ( .A(n27164), .B(n18467), .Z(n18468) );
  NAND U25471 ( .A(n27167), .B(n18468), .Z(n18469) );
  NANDN U25472 ( .A(n27169), .B(n18469), .Z(n18470) );
  NANDN U25473 ( .A(n24339), .B(n18470), .Z(n18471) );
  AND U25474 ( .A(n27170), .B(n18471), .Z(n18472) );
  ANDN U25475 ( .B(n18473), .A(n18472), .Z(n18474) );
  NAND U25476 ( .A(n27171), .B(n18474), .Z(n18475) );
  NANDN U25477 ( .A(n18476), .B(n18475), .Z(n18477) );
  OR U25478 ( .A(n27172), .B(n18477), .Z(n18478) );
  AND U25479 ( .A(n18479), .B(n18478), .Z(n18481) );
  NAND U25480 ( .A(n18481), .B(n18480), .Z(n18483) );
  ANDN U25481 ( .B(n18483), .A(n18482), .Z(n18484) );
  NANDN U25482 ( .A(n18485), .B(n18484), .Z(n18488) );
  AND U25483 ( .A(n18486), .B(n27177), .Z(n18487) );
  NAND U25484 ( .A(n18488), .B(n18487), .Z(n18489) );
  NANDN U25485 ( .A(n27178), .B(n18489), .Z(n18491) );
  OR U25486 ( .A(n18491), .B(n18490), .Z(n18492) );
  NAND U25487 ( .A(n27179), .B(n18492), .Z(n18493) );
  NANDN U25488 ( .A(n27180), .B(n18493), .Z(n18494) );
  NAND U25489 ( .A(n27181), .B(n18494), .Z(n18495) );
  AND U25490 ( .A(n27182), .B(n18495), .Z(n18496) );
  OR U25491 ( .A(n27183), .B(n18496), .Z(n18497) );
  NAND U25492 ( .A(n27184), .B(n18497), .Z(n18498) );
  NANDN U25493 ( .A(n27185), .B(n18498), .Z(n18502) );
  IV U25494 ( .A(n18499), .Z(n27186) );
  AND U25495 ( .A(n18500), .B(n27186), .Z(n18501) );
  NAND U25496 ( .A(n18502), .B(n18501), .Z(n18503) );
  NANDN U25497 ( .A(n18504), .B(n18503), .Z(n18506) );
  IV U25498 ( .A(n18505), .Z(n27187) );
  OR U25499 ( .A(n18506), .B(n27187), .Z(n18507) );
  NANDN U25500 ( .A(n18508), .B(n18507), .Z(n18509) );
  AND U25501 ( .A(n18510), .B(n18509), .Z(n18513) );
  NANDN U25502 ( .A(n18513), .B(n27193), .Z(n18514) );
  NAND U25503 ( .A(n27194), .B(n18514), .Z(n18515) );
  NAND U25504 ( .A(n27195), .B(n18515), .Z(n18516) );
  NANDN U25505 ( .A(n27196), .B(n18516), .Z(n18517) );
  AND U25506 ( .A(n27197), .B(n18517), .Z(n18518) );
  ANDN U25507 ( .B(n18519), .A(n18518), .Z(n18520) );
  NAND U25508 ( .A(n27198), .B(n18520), .Z(n18521) );
  NAND U25509 ( .A(n27199), .B(n18521), .Z(n18522) );
  AND U25510 ( .A(n18523), .B(n18522), .Z(n18526) );
  AND U25511 ( .A(n27201), .B(n18524), .Z(n18525) );
  NANDN U25512 ( .A(n18526), .B(n18525), .Z(n18527) );
  NANDN U25513 ( .A(n18528), .B(n18527), .Z(n18529) );
  AND U25514 ( .A(n27205), .B(n18529), .Z(n18531) );
  NAND U25515 ( .A(n18531), .B(n18530), .Z(n18532) );
  NANDN U25516 ( .A(n27207), .B(n18532), .Z(n18533) );
  AND U25517 ( .A(n27209), .B(n18533), .Z(n18536) );
  NAND U25518 ( .A(n18535), .B(n18534), .Z(n24338) );
  OR U25519 ( .A(n18536), .B(n24338), .Z(n18537) );
  NAND U25520 ( .A(n24337), .B(n18537), .Z(n18538) );
  NANDN U25521 ( .A(n27210), .B(n18538), .Z(n18539) );
  AND U25522 ( .A(n27211), .B(n18539), .Z(n18540) );
  OR U25523 ( .A(n27212), .B(n18540), .Z(n18541) );
  NAND U25524 ( .A(n27213), .B(n18541), .Z(n18542) );
  NANDN U25525 ( .A(n18543), .B(n18542), .Z(n18544) );
  OR U25526 ( .A(n27214), .B(n18544), .Z(n18545) );
  AND U25527 ( .A(n27215), .B(n18545), .Z(n18546) );
  NANDN U25528 ( .A(n27217), .B(n18546), .Z(n18547) );
  AND U25529 ( .A(n18548), .B(n18547), .Z(n18555) );
  ANDN U25530 ( .B(n18550), .A(n18549), .Z(n27220) );
  NAND U25531 ( .A(n18552), .B(n18551), .Z(n27219) );
  NANDN U25532 ( .A(n24335), .B(n27219), .Z(n18553) );
  AND U25533 ( .A(n27220), .B(n18553), .Z(n18554) );
  NANDN U25534 ( .A(n18555), .B(n18554), .Z(n18556) );
  AND U25535 ( .A(n18557), .B(n18556), .Z(n18558) );
  OR U25536 ( .A(n27222), .B(n18558), .Z(n18559) );
  NAND U25537 ( .A(n18560), .B(n18559), .Z(n18561) );
  NANDN U25538 ( .A(n18562), .B(n18561), .Z(n18564) );
  IV U25539 ( .A(n18563), .Z(n27224) );
  OR U25540 ( .A(n18564), .B(n27224), .Z(n18565) );
  NAND U25541 ( .A(n18566), .B(n18565), .Z(n18570) );
  AND U25542 ( .A(n18568), .B(n18567), .Z(n18569) );
  NAND U25543 ( .A(n18570), .B(n18569), .Z(n18571) );
  NANDN U25544 ( .A(n27228), .B(n18571), .Z(n18572) );
  OR U25545 ( .A(n18573), .B(n18572), .Z(n18574) );
  AND U25546 ( .A(n18575), .B(n18574), .Z(n18576) );
  NANDN U25547 ( .A(n27229), .B(n18576), .Z(n18579) );
  AND U25548 ( .A(n18578), .B(n18577), .Z(n27230) );
  AND U25549 ( .A(n18579), .B(n27230), .Z(n18582) );
  NANDN U25550 ( .A(n18582), .B(n27231), .Z(n18583) );
  NAND U25551 ( .A(n27232), .B(n18583), .Z(n18584) );
  NAND U25552 ( .A(n27233), .B(n18584), .Z(n18585) );
  AND U25553 ( .A(n18585), .B(n27235), .Z(n18588) );
  NANDN U25554 ( .A(n18588), .B(n27237), .Z(n18589) );
  NAND U25555 ( .A(n24331), .B(n18589), .Z(n18590) );
  NANDN U25556 ( .A(n18591), .B(n18590), .Z(n18592) );
  OR U25557 ( .A(n18592), .B(n27238), .Z(n18593) );
  NAND U25558 ( .A(n18594), .B(n18593), .Z(n18598) );
  IV U25559 ( .A(n18595), .Z(n27241) );
  AND U25560 ( .A(n18596), .B(n27241), .Z(n18597) );
  NAND U25561 ( .A(n18598), .B(n18597), .Z(n18599) );
  NANDN U25562 ( .A(n18600), .B(n18599), .Z(n18602) );
  IV U25563 ( .A(n18601), .Z(n27242) );
  OR U25564 ( .A(n18602), .B(n27242), .Z(n18603) );
  AND U25565 ( .A(n27243), .B(n18603), .Z(n18606) );
  NAND U25566 ( .A(n18605), .B(n18604), .Z(n27244) );
  OR U25567 ( .A(n18606), .B(n27244), .Z(n18607) );
  NAND U25568 ( .A(n27245), .B(n18607), .Z(n18608) );
  NAND U25569 ( .A(n27246), .B(n18608), .Z(n18609) );
  NAND U25570 ( .A(n27247), .B(n18609), .Z(n18610) );
  AND U25571 ( .A(n18611), .B(n18610), .Z(n18612) );
  OR U25572 ( .A(n18613), .B(n18612), .Z(n18614) );
  NAND U25573 ( .A(n18615), .B(n18614), .Z(n18616) );
  NANDN U25574 ( .A(n18617), .B(n18616), .Z(n18621) );
  IV U25575 ( .A(n18618), .Z(n27253) );
  AND U25576 ( .A(n18619), .B(n27253), .Z(n18620) );
  NAND U25577 ( .A(n18621), .B(n18620), .Z(n18622) );
  NANDN U25578 ( .A(n18623), .B(n18622), .Z(n18625) );
  IV U25579 ( .A(n18624), .Z(n27254) );
  OR U25580 ( .A(n18625), .B(n27254), .Z(n18626) );
  AND U25581 ( .A(n27255), .B(n18626), .Z(n18627) );
  OR U25582 ( .A(n27256), .B(n18627), .Z(n18628) );
  NAND U25583 ( .A(n27257), .B(n18628), .Z(n18629) );
  NANDN U25584 ( .A(n27258), .B(n18629), .Z(n18630) );
  AND U25585 ( .A(n27259), .B(n18630), .Z(n18631) );
  OR U25586 ( .A(n27260), .B(n18631), .Z(n18632) );
  NAND U25587 ( .A(n27261), .B(n18632), .Z(n18633) );
  NANDN U25588 ( .A(n18634), .B(n18633), .Z(n18636) );
  IV U25589 ( .A(n18635), .Z(n27262) );
  OR U25590 ( .A(n18636), .B(n27262), .Z(n18637) );
  AND U25591 ( .A(n18638), .B(n18637), .Z(n18639) );
  NAND U25592 ( .A(n18639), .B(n27263), .Z(n18641) );
  ANDN U25593 ( .B(n18641), .A(n18640), .Z(n18642) );
  NANDN U25594 ( .A(n27267), .B(n18642), .Z(n18645) );
  AND U25595 ( .A(n27268), .B(n18643), .Z(n18644) );
  NAND U25596 ( .A(n18645), .B(n18644), .Z(n18646) );
  NANDN U25597 ( .A(n27269), .B(n18646), .Z(n18647) );
  AND U25598 ( .A(n27270), .B(n18647), .Z(n18648) );
  OR U25599 ( .A(n27271), .B(n18648), .Z(n18649) );
  NAND U25600 ( .A(n27272), .B(n18649), .Z(n18650) );
  NANDN U25601 ( .A(n27273), .B(n18650), .Z(n18651) );
  NAND U25602 ( .A(n24327), .B(n18651), .Z(n18652) );
  ANDN U25603 ( .B(n18652), .A(n27274), .Z(n18653) );
  NANDN U25604 ( .A(n18654), .B(n18653), .Z(n18655) );
  AND U25605 ( .A(n18656), .B(n18655), .Z(n18657) );
  OR U25606 ( .A(n18658), .B(n18657), .Z(n18659) );
  NAND U25607 ( .A(n24325), .B(n18659), .Z(n18660) );
  NANDN U25608 ( .A(n24324), .B(n18660), .Z(n18661) );
  NAND U25609 ( .A(n24323), .B(n18661), .Z(n18662) );
  NAND U25610 ( .A(n27280), .B(n18662), .Z(n18663) );
  NANDN U25611 ( .A(n27281), .B(n18663), .Z(n18666) );
  AND U25612 ( .A(n18664), .B(n27282), .Z(n18665) );
  NAND U25613 ( .A(n18666), .B(n18665), .Z(n18667) );
  NANDN U25614 ( .A(n18668), .B(n18667), .Z(n18669) );
  OR U25615 ( .A(n27283), .B(n18669), .Z(n18670) );
  AND U25616 ( .A(n18671), .B(n18670), .Z(n18672) );
  NANDN U25617 ( .A(n27286), .B(n18672), .Z(n18673) );
  AND U25618 ( .A(n18674), .B(n18673), .Z(n18678) );
  NANDN U25619 ( .A(n18678), .B(n27288), .Z(n18679) );
  NAND U25620 ( .A(n27289), .B(n18679), .Z(n18680) );
  NAND U25621 ( .A(n27290), .B(n18680), .Z(n18681) );
  AND U25622 ( .A(n18681), .B(n27291), .Z(n18682) );
  OR U25623 ( .A(n18682), .B(n24322), .Z(n18683) );
  NAND U25624 ( .A(n24321), .B(n18683), .Z(n18684) );
  NANDN U25625 ( .A(n27294), .B(n18684), .Z(n18685) );
  NAND U25626 ( .A(n27295), .B(n18685), .Z(n18686) );
  NAND U25627 ( .A(n18687), .B(n18686), .Z(n18688) );
  NANDN U25628 ( .A(n18689), .B(n18688), .Z(n18690) );
  AND U25629 ( .A(n18691), .B(n18690), .Z(n18692) );
  NAND U25630 ( .A(n27297), .B(n18692), .Z(n18695) );
  NAND U25631 ( .A(n27298), .B(n18693), .Z(n18694) );
  ANDN U25632 ( .B(n18695), .A(n18694), .Z(n18696) );
  OR U25633 ( .A(n27299), .B(n18696), .Z(n18697) );
  NAND U25634 ( .A(n27300), .B(n18697), .Z(n18698) );
  NANDN U25635 ( .A(n27301), .B(n18698), .Z(n18699) );
  NAND U25636 ( .A(n27302), .B(n18699), .Z(n18701) );
  IV U25637 ( .A(n18700), .Z(n27303) );
  ANDN U25638 ( .B(n18701), .A(n27303), .Z(n18702) );
  NANDN U25639 ( .A(n18703), .B(n18702), .Z(n18707) );
  IV U25640 ( .A(n18704), .Z(n27304) );
  AND U25641 ( .A(n18705), .B(n27304), .Z(n18706) );
  NAND U25642 ( .A(n18707), .B(n18706), .Z(n18708) );
  NANDN U25643 ( .A(n27307), .B(n18708), .Z(n18709) );
  OR U25644 ( .A(n18710), .B(n18709), .Z(n18711) );
  AND U25645 ( .A(n18712), .B(n18711), .Z(n18713) );
  NANDN U25646 ( .A(n27309), .B(n18713), .Z(n18714) );
  AND U25647 ( .A(n27310), .B(n18714), .Z(n18715) );
  OR U25648 ( .A(n27311), .B(n18715), .Z(n18716) );
  NAND U25649 ( .A(n27312), .B(n18716), .Z(n18717) );
  NANDN U25650 ( .A(n18718), .B(n18717), .Z(n18722) );
  IV U25651 ( .A(n18719), .Z(n27314) );
  AND U25652 ( .A(n18720), .B(n27314), .Z(n18721) );
  NAND U25653 ( .A(n18722), .B(n18721), .Z(n18723) );
  NANDN U25654 ( .A(n27317), .B(n18723), .Z(n18725) );
  OR U25655 ( .A(n18725), .B(n18724), .Z(n18726) );
  NAND U25656 ( .A(n18727), .B(n18726), .Z(n18728) );
  NANDN U25657 ( .A(n27319), .B(n18728), .Z(n18729) );
  NAND U25658 ( .A(n27320), .B(n18729), .Z(n18730) );
  NANDN U25659 ( .A(n27321), .B(n18730), .Z(n18731) );
  AND U25660 ( .A(n18732), .B(n18731), .Z(n18733) );
  OR U25661 ( .A(n27323), .B(n18733), .Z(n18734) );
  NAND U25662 ( .A(n18735), .B(n18734), .Z(n18736) );
  NANDN U25663 ( .A(n27324), .B(n18736), .Z(n18737) );
  OR U25664 ( .A(n18738), .B(n18737), .Z(n18739) );
  AND U25665 ( .A(n18740), .B(n18739), .Z(n18741) );
  NANDN U25666 ( .A(n27325), .B(n18741), .Z(n18742) );
  AND U25667 ( .A(n18743), .B(n18742), .Z(n18744) );
  NOR U25668 ( .A(n18744), .B(n27331), .Z(n18745) );
  NANDN U25669 ( .A(n18746), .B(n18745), .Z(n18747) );
  AND U25670 ( .A(n18747), .B(n27332), .Z(n18749) );
  NAND U25671 ( .A(n18749), .B(n18748), .Z(n18750) );
  NAND U25672 ( .A(n27333), .B(n18750), .Z(n18751) );
  AND U25673 ( .A(n18751), .B(n24316), .Z(n18752) );
  OR U25674 ( .A(n18752), .B(n24315), .Z(n18753) );
  NAND U25675 ( .A(n27334), .B(n18753), .Z(n18754) );
  NANDN U25676 ( .A(n27335), .B(n18754), .Z(n18755) );
  AND U25677 ( .A(n27336), .B(n18755), .Z(n18759) );
  NANDN U25678 ( .A(n18759), .B(n27337), .Z(n18760) );
  NANDN U25679 ( .A(n27338), .B(n18760), .Z(n18761) );
  AND U25680 ( .A(n27339), .B(n18761), .Z(n18763) );
  IV U25681 ( .A(n18762), .Z(n27340) );
  OR U25682 ( .A(n18763), .B(n27340), .Z(n18764) );
  AND U25683 ( .A(n27341), .B(n18764), .Z(n18765) );
  OR U25684 ( .A(n27342), .B(n18765), .Z(n18766) );
  NAND U25685 ( .A(n27344), .B(n18766), .Z(n18767) );
  NANDN U25686 ( .A(n27345), .B(n18767), .Z(n18768) );
  AND U25687 ( .A(n18769), .B(n18768), .Z(n18770) );
  OR U25688 ( .A(n27347), .B(n18770), .Z(n18771) );
  NAND U25689 ( .A(n18772), .B(n18771), .Z(n18773) );
  NANDN U25690 ( .A(n27351), .B(n18773), .Z(n18774) );
  AND U25691 ( .A(n18775), .B(n18774), .Z(n18776) );
  NAND U25692 ( .A(n27352), .B(n18776), .Z(n18777) );
  NANDN U25693 ( .A(n18778), .B(n18777), .Z(n18780) );
  IV U25694 ( .A(n18779), .Z(n27353) );
  OR U25695 ( .A(n18780), .B(n27353), .Z(n18781) );
  NAND U25696 ( .A(n18782), .B(n18781), .Z(n18783) );
  NANDN U25697 ( .A(n18784), .B(n18783), .Z(n18786) );
  OR U25698 ( .A(n18786), .B(n18785), .Z(n18787) );
  AND U25699 ( .A(n18788), .B(n18787), .Z(n18789) );
  OR U25700 ( .A(n18790), .B(n18789), .Z(n18791) );
  NAND U25701 ( .A(n18792), .B(n18791), .Z(n18793) );
  AND U25702 ( .A(n18794), .B(n18793), .Z(n18796) );
  IV U25703 ( .A(n18795), .Z(n27362) );
  OR U25704 ( .A(n18796), .B(n27362), .Z(n18797) );
  NAND U25705 ( .A(n27363), .B(n18797), .Z(n18798) );
  NANDN U25706 ( .A(n27364), .B(n18798), .Z(n18800) );
  NAND U25707 ( .A(n18800), .B(n18799), .Z(n18801) );
  NANDN U25708 ( .A(n18802), .B(n18801), .Z(n18803) );
  AND U25709 ( .A(n18804), .B(n18803), .Z(n18806) );
  NAND U25710 ( .A(n18806), .B(n18805), .Z(n18808) );
  ANDN U25711 ( .B(n18808), .A(n18807), .Z(n18809) );
  NANDN U25712 ( .A(n18810), .B(n18809), .Z(n18811) );
  AND U25713 ( .A(n18812), .B(n18811), .Z(n18813) );
  OR U25714 ( .A(n18814), .B(n18813), .Z(n18815) );
  NAND U25715 ( .A(n27370), .B(n18815), .Z(n18816) );
  NANDN U25716 ( .A(n18817), .B(n18816), .Z(n18818) );
  ANDN U25717 ( .B(y[2040]), .A(x[2040]), .Z(n27371) );
  OR U25718 ( .A(n18818), .B(n27371), .Z(n18819) );
  AND U25719 ( .A(n18820), .B(n18819), .Z(n18821) );
  OR U25720 ( .A(n18822), .B(n18821), .Z(n18823) );
  NAND U25721 ( .A(n27376), .B(n18823), .Z(n18824) );
  NANDN U25722 ( .A(n18825), .B(n18824), .Z(n18826) );
  ANDN U25723 ( .B(y[2044]), .A(x[2044]), .Z(n27377) );
  OR U25724 ( .A(n18826), .B(n27377), .Z(n18827) );
  AND U25725 ( .A(n18828), .B(n18827), .Z(n18829) );
  NOR U25726 ( .A(n27381), .B(n18829), .Z(n18830) );
  NANDN U25727 ( .A(n18831), .B(n18830), .Z(n18832) );
  AND U25728 ( .A(n18833), .B(n18832), .Z(n18834) );
  NAND U25729 ( .A(n27382), .B(n18834), .Z(n18835) );
  NAND U25730 ( .A(n27383), .B(n18835), .Z(n18836) );
  AND U25731 ( .A(n18837), .B(n18836), .Z(n18838) );
  ANDN U25732 ( .B(n18839), .A(n18838), .Z(n18840) );
  NAND U25733 ( .A(n27385), .B(n18840), .Z(n18841) );
  NANDN U25734 ( .A(n18842), .B(n18841), .Z(n18843) );
  OR U25735 ( .A(n18844), .B(n18843), .Z(n18845) );
  AND U25736 ( .A(n18846), .B(n18845), .Z(n18847) );
  NANDN U25737 ( .A(n27390), .B(n18847), .Z(n18848) );
  AND U25738 ( .A(n18849), .B(n18848), .Z(n18852) );
  NAND U25739 ( .A(n18851), .B(n18850), .Z(n27392) );
  OR U25740 ( .A(n18852), .B(n27392), .Z(n18853) );
  NAND U25741 ( .A(n18854), .B(n18853), .Z(n18855) );
  NANDN U25742 ( .A(n24310), .B(n18855), .Z(n18856) );
  NAND U25743 ( .A(n18857), .B(n18856), .Z(n18858) );
  NANDN U25744 ( .A(n27395), .B(n18858), .Z(n18859) );
  AND U25745 ( .A(n27396), .B(n18859), .Z(n18862) );
  NAND U25746 ( .A(n18861), .B(n18860), .Z(n24307) );
  OR U25747 ( .A(n18862), .B(n24307), .Z(n18863) );
  NAND U25748 ( .A(n27397), .B(n18863), .Z(n18864) );
  NANDN U25749 ( .A(n18865), .B(n18864), .Z(n18866) );
  AND U25750 ( .A(n27399), .B(n18866), .Z(n18867) );
  OR U25751 ( .A(n18868), .B(n18867), .Z(n18869) );
  NAND U25752 ( .A(n27405), .B(n18869), .Z(n18870) );
  NANDN U25753 ( .A(n18871), .B(n18870), .Z(n18872) );
  ANDN U25754 ( .B(y[2066]), .A(x[2066]), .Z(n27406) );
  OR U25755 ( .A(n18872), .B(n27406), .Z(n18873) );
  NAND U25756 ( .A(n27407), .B(n18873), .Z(n18874) );
  NANDN U25757 ( .A(n27408), .B(n18874), .Z(n18875) );
  OR U25758 ( .A(n18876), .B(n18875), .Z(n18877) );
  AND U25759 ( .A(n27409), .B(n18877), .Z(n18880) );
  NANDN U25760 ( .A(x[2070]), .B(y[2070]), .Z(n18879) );
  NAND U25761 ( .A(n18879), .B(n18878), .Z(n27410) );
  OR U25762 ( .A(n18880), .B(n27410), .Z(n18881) );
  NAND U25763 ( .A(n18882), .B(n18881), .Z(n18883) );
  NANDN U25764 ( .A(n18884), .B(n18883), .Z(n18885) );
  OR U25765 ( .A(n18885), .B(n27411), .Z(n18886) );
  NAND U25766 ( .A(n18887), .B(n18886), .Z(n18890) );
  AND U25767 ( .A(n18888), .B(n27415), .Z(n18889) );
  NAND U25768 ( .A(n18890), .B(n18889), .Z(n18891) );
  NANDN U25769 ( .A(n18892), .B(n18891), .Z(n18894) );
  IV U25770 ( .A(n18893), .Z(n27416) );
  OR U25771 ( .A(n18894), .B(n27416), .Z(n18895) );
  NAND U25772 ( .A(n27417), .B(n18895), .Z(n18896) );
  NANDN U25773 ( .A(n27419), .B(n18896), .Z(n18897) );
  NAND U25774 ( .A(n27420), .B(n18897), .Z(n18898) );
  NAND U25775 ( .A(n27421), .B(n18898), .Z(n18899) );
  NANDN U25776 ( .A(n24303), .B(n18899), .Z(n18900) );
  AND U25777 ( .A(n18900), .B(n24302), .Z(n18901) );
  OR U25778 ( .A(n18901), .B(n27422), .Z(n18902) );
  NAND U25779 ( .A(n18903), .B(n18902), .Z(n18904) );
  NANDN U25780 ( .A(n18905), .B(n18904), .Z(n18906) );
  AND U25781 ( .A(n18907), .B(n18906), .Z(n18908) );
  OR U25782 ( .A(n18909), .B(n18908), .Z(n18910) );
  NANDN U25783 ( .A(n27425), .B(n18910), .Z(n18911) );
  NANDN U25784 ( .A(n18912), .B(n18911), .Z(n18913) );
  AND U25785 ( .A(n18914), .B(n18913), .Z(n18915) );
  OR U25786 ( .A(n18916), .B(n18915), .Z(n18917) );
  NAND U25787 ( .A(n27431), .B(n18917), .Z(n18918) );
  NAND U25788 ( .A(n27432), .B(n18918), .Z(n18921) );
  AND U25789 ( .A(n18919), .B(n27433), .Z(n18920) );
  NAND U25790 ( .A(n18921), .B(n18920), .Z(n18922) );
  NANDN U25791 ( .A(n18923), .B(n18922), .Z(n18924) );
  OR U25792 ( .A(n18924), .B(n24299), .Z(n18925) );
  AND U25793 ( .A(n18926), .B(n18925), .Z(n18928) );
  NAND U25794 ( .A(n18928), .B(n18927), .Z(n18930) );
  ANDN U25795 ( .B(n18930), .A(n18929), .Z(n18931) );
  NANDN U25796 ( .A(n24297), .B(n18931), .Z(n18932) );
  NAND U25797 ( .A(n18933), .B(n18932), .Z(n18934) );
  NAND U25798 ( .A(n27436), .B(n18934), .Z(n18937) );
  AND U25799 ( .A(n18936), .B(n18935), .Z(n24295) );
  AND U25800 ( .A(n18937), .B(n24295), .Z(n18938) );
  OR U25801 ( .A(n27439), .B(n18938), .Z(n18939) );
  NAND U25802 ( .A(n27440), .B(n18939), .Z(n18940) );
  NAND U25803 ( .A(n27441), .B(n18940), .Z(n18943) );
  AND U25804 ( .A(n18942), .B(n18941), .Z(n27442) );
  AND U25805 ( .A(n18943), .B(n27442), .Z(n18946) );
  NANDN U25806 ( .A(n18946), .B(n27443), .Z(n18947) );
  NAND U25807 ( .A(n24294), .B(n18947), .Z(n18948) );
  NANDN U25808 ( .A(n18949), .B(n18948), .Z(n18950) );
  NANDN U25809 ( .A(n18950), .B(n27444), .Z(n18951) );
  AND U25810 ( .A(n18952), .B(n18951), .Z(n18953) );
  OR U25811 ( .A(n18954), .B(n18953), .Z(n18955) );
  NAND U25812 ( .A(n24292), .B(n18955), .Z(n18956) );
  NANDN U25813 ( .A(n18957), .B(n18956), .Z(n18959) );
  IV U25814 ( .A(n18958), .Z(n24293) );
  OR U25815 ( .A(n18959), .B(n24293), .Z(n18960) );
  AND U25816 ( .A(n18961), .B(n18960), .Z(n18964) );
  NAND U25817 ( .A(n27453), .B(n18962), .Z(n18963) );
  OR U25818 ( .A(n18964), .B(n18963), .Z(n18965) );
  AND U25819 ( .A(n18966), .B(n18965), .Z(n18967) );
  OR U25820 ( .A(n27456), .B(n18967), .Z(n18968) );
  NAND U25821 ( .A(n18969), .B(n18968), .Z(n18970) );
  NANDN U25822 ( .A(n27458), .B(n18970), .Z(n18974) );
  AND U25823 ( .A(n18972), .B(n18971), .Z(n18973) );
  NAND U25824 ( .A(n18974), .B(n18973), .Z(n18975) );
  NANDN U25825 ( .A(n27460), .B(n18975), .Z(n18976) );
  OR U25826 ( .A(n18976), .B(n24291), .Z(n18977) );
  NAND U25827 ( .A(n18978), .B(n18977), .Z(n18979) );
  NAND U25828 ( .A(n27463), .B(n18979), .Z(n18982) );
  AND U25829 ( .A(n18980), .B(n27464), .Z(n18981) );
  NAND U25830 ( .A(n18982), .B(n18981), .Z(n18983) );
  NANDN U25831 ( .A(n27465), .B(n18983), .Z(n18984) );
  OR U25832 ( .A(n18984), .B(n27467), .Z(n18985) );
  AND U25833 ( .A(n18986), .B(n18985), .Z(n18989) );
  NAND U25834 ( .A(n18988), .B(n18987), .Z(n24290) );
  OR U25835 ( .A(n18989), .B(n24290), .Z(n18990) );
  NAND U25836 ( .A(n27470), .B(n18990), .Z(n18991) );
  NANDN U25837 ( .A(n27471), .B(n18991), .Z(n18992) );
  NAND U25838 ( .A(n27473), .B(n18992), .Z(n18993) );
  ANDN U25839 ( .B(n18993), .A(n27474), .Z(n18994) );
  NANDN U25840 ( .A(n18995), .B(n18994), .Z(n18996) );
  AND U25841 ( .A(n18996), .B(n27475), .Z(n18997) );
  OR U25842 ( .A(n18998), .B(n18997), .Z(n18999) );
  NAND U25843 ( .A(n27477), .B(n18999), .Z(n19000) );
  NANDN U25844 ( .A(n27478), .B(n19000), .Z(n19002) );
  OR U25845 ( .A(n19002), .B(n19001), .Z(n19003) );
  NAND U25846 ( .A(n19004), .B(n19003), .Z(n19005) );
  NANDN U25847 ( .A(n19006), .B(n19005), .Z(n19008) );
  OR U25848 ( .A(n19008), .B(n19007), .Z(n19012) );
  OR U25849 ( .A(n19010), .B(n19009), .Z(n19011) );
  AND U25850 ( .A(n19012), .B(n19011), .Z(n19013) );
  AND U25851 ( .A(n27483), .B(n19013), .Z(n19014) );
  NANDN U25852 ( .A(n19014), .B(n27485), .Z(n19015) );
  NAND U25853 ( .A(n27487), .B(n19015), .Z(n19016) );
  NANDN U25854 ( .A(n19017), .B(n19016), .Z(n19018) );
  NAND U25855 ( .A(n19019), .B(n19018), .Z(n19020) );
  NAND U25856 ( .A(n19021), .B(n19020), .Z(n19022) );
  NAND U25857 ( .A(n27491), .B(n19022), .Z(n19023) );
  NAND U25858 ( .A(n27492), .B(n19023), .Z(n19024) );
  NAND U25859 ( .A(n27493), .B(n19024), .Z(n19025) );
  NAND U25860 ( .A(n27494), .B(n19025), .Z(n19028) );
  AND U25861 ( .A(n19027), .B(n19026), .Z(n27495) );
  AND U25862 ( .A(n19028), .B(n27495), .Z(n19031) );
  NANDN U25863 ( .A(n19031), .B(n27496), .Z(n19032) );
  NAND U25864 ( .A(n24289), .B(n19032), .Z(n19033) );
  NANDN U25865 ( .A(n19034), .B(n19033), .Z(n19035) );
  NANDN U25866 ( .A(n19035), .B(n27497), .Z(n19036) );
  NAND U25867 ( .A(n19037), .B(n19036), .Z(n19038) );
  NANDN U25868 ( .A(n19039), .B(n19038), .Z(n19040) );
  OR U25869 ( .A(n19041), .B(n19040), .Z(n19042) );
  AND U25870 ( .A(n24287), .B(n19042), .Z(n19043) );
  ANDN U25871 ( .B(n19044), .A(n19043), .Z(n19045) );
  NAND U25872 ( .A(n24288), .B(n19045), .Z(n19046) );
  NANDN U25873 ( .A(n19047), .B(n19046), .Z(n19048) );
  OR U25874 ( .A(n19048), .B(n27502), .Z(n19049) );
  AND U25875 ( .A(n19050), .B(n19049), .Z(n19051) );
  OR U25876 ( .A(n19052), .B(n19051), .Z(n19053) );
  NAND U25877 ( .A(n27508), .B(n19053), .Z(n19054) );
  NANDN U25878 ( .A(n19055), .B(n19054), .Z(n19056) );
  OR U25879 ( .A(n27509), .B(n19056), .Z(n19057) );
  AND U25880 ( .A(n27510), .B(n19057), .Z(n19058) );
  ANDN U25881 ( .B(n19059), .A(n19058), .Z(n19060) );
  NANDN U25882 ( .A(n19061), .B(n19060), .Z(n19062) );
  AND U25883 ( .A(n27512), .B(n19062), .Z(n19063) );
  OR U25884 ( .A(n27513), .B(n19063), .Z(n19064) );
  NAND U25885 ( .A(n27514), .B(n19064), .Z(n19065) );
  NANDN U25886 ( .A(n19066), .B(n19065), .Z(n19067) );
  OR U25887 ( .A(n19067), .B(n27515), .Z(n19068) );
  NANDN U25888 ( .A(n19069), .B(n19068), .Z(n19070) );
  AND U25889 ( .A(n19071), .B(n19070), .Z(n19075) );
  NAND U25890 ( .A(n19073), .B(n19072), .Z(n19074) );
  OR U25891 ( .A(n19075), .B(n19074), .Z(n19076) );
  AND U25892 ( .A(n19077), .B(n19076), .Z(n19081) );
  NAND U25893 ( .A(n19079), .B(n19078), .Z(n19080) );
  OR U25894 ( .A(n19081), .B(n19080), .Z(n19082) );
  AND U25895 ( .A(n19083), .B(n19082), .Z(n19085) );
  NOR U25896 ( .A(n19085), .B(n19084), .Z(n19086) );
  NANDN U25897 ( .A(n19087), .B(n19086), .Z(n19089) );
  IV U25898 ( .A(n19088), .Z(n27523) );
  AND U25899 ( .A(n19089), .B(n27523), .Z(n19090) );
  NANDN U25900 ( .A(n19091), .B(n19090), .Z(n19092) );
  AND U25901 ( .A(n19092), .B(n27524), .Z(n19093) );
  NANDN U25902 ( .A(n19094), .B(n19093), .Z(n19095) );
  AND U25903 ( .A(n27525), .B(n19095), .Z(n19096) );
  NOR U25904 ( .A(n27526), .B(n19096), .Z(n19097) );
  NANDN U25905 ( .A(n19098), .B(n19097), .Z(n19099) );
  AND U25906 ( .A(n27527), .B(n19099), .Z(n19101) );
  NAND U25907 ( .A(n19101), .B(n19100), .Z(n19102) );
  NANDN U25908 ( .A(n19103), .B(n19102), .Z(n19104) );
  AND U25909 ( .A(n19105), .B(n19104), .Z(n19107) );
  NAND U25910 ( .A(n19107), .B(n19106), .Z(n19108) );
  NAND U25911 ( .A(n27532), .B(n19108), .Z(n19109) );
  AND U25912 ( .A(n19110), .B(n19109), .Z(n19113) );
  NAND U25913 ( .A(n19112), .B(n19111), .Z(n27533) );
  NAND U25914 ( .A(n19113), .B(n27533), .Z(n19114) );
  NANDN U25915 ( .A(n19115), .B(n19114), .Z(n19116) );
  AND U25916 ( .A(n19117), .B(n19116), .Z(n19120) );
  NANDN U25917 ( .A(n19120), .B(n24279), .Z(n19121) );
  NAND U25918 ( .A(n19122), .B(n19121), .Z(n19123) );
  NANDN U25919 ( .A(n19124), .B(n19123), .Z(n19125) );
  OR U25920 ( .A(n24280), .B(n19125), .Z(n19126) );
  AND U25921 ( .A(n19127), .B(n19126), .Z(n19128) );
  NANDN U25922 ( .A(n19129), .B(n19128), .Z(n19130) );
  AND U25923 ( .A(n19131), .B(n19130), .Z(n19135) );
  NAND U25924 ( .A(n19133), .B(n19132), .Z(n19134) );
  OR U25925 ( .A(n19135), .B(n19134), .Z(n19136) );
  AND U25926 ( .A(n19137), .B(n19136), .Z(n19141) );
  NAND U25927 ( .A(n19139), .B(n19138), .Z(n19140) );
  OR U25928 ( .A(n19141), .B(n19140), .Z(n19142) );
  AND U25929 ( .A(n19143), .B(n19142), .Z(n19144) );
  NOR U25930 ( .A(n19144), .B(n27545), .Z(n19145) );
  NANDN U25931 ( .A(n19146), .B(n19145), .Z(n19147) );
  AND U25932 ( .A(n19148), .B(n19147), .Z(n19149) );
  AND U25933 ( .A(n19149), .B(n27546), .Z(n19154) );
  OR U25934 ( .A(n19154), .B(n27547), .Z(n19155) );
  NAND U25935 ( .A(n27548), .B(n19155), .Z(n19156) );
  NANDN U25936 ( .A(n24276), .B(n19156), .Z(n19157) );
  AND U25937 ( .A(n27549), .B(n19157), .Z(n19159) );
  OR U25938 ( .A(n19159), .B(n19158), .Z(n19160) );
  NAND U25939 ( .A(n24275), .B(n19160), .Z(n19161) );
  NANDN U25940 ( .A(n19162), .B(n19161), .Z(n19163) );
  OR U25941 ( .A(n19163), .B(n27551), .Z(n19164) );
  NAND U25942 ( .A(n27552), .B(n19164), .Z(n19165) );
  NANDN U25943 ( .A(n19166), .B(n19165), .Z(n19167) );
  NAND U25944 ( .A(n27557), .B(n19167), .Z(n19168) );
  NAND U25945 ( .A(n27558), .B(n19168), .Z(n19169) );
  NAND U25946 ( .A(n27559), .B(n19169), .Z(n19170) );
  AND U25947 ( .A(n27560), .B(n19170), .Z(n19173) );
  NAND U25948 ( .A(n19172), .B(n19171), .Z(n27561) );
  OR U25949 ( .A(n19173), .B(n27561), .Z(n19174) );
  AND U25950 ( .A(n27562), .B(n19174), .Z(n19175) );
  NANDN U25951 ( .A(n19175), .B(n27563), .Z(n19176) );
  NAND U25952 ( .A(n27564), .B(n19176), .Z(n19179) );
  NANDN U25953 ( .A(x[2218]), .B(y[2218]), .Z(n19178) );
  AND U25954 ( .A(n19178), .B(n19177), .Z(n24274) );
  AND U25955 ( .A(n19179), .B(n24274), .Z(n19182) );
  NANDN U25956 ( .A(n19182), .B(n27565), .Z(n19183) );
  AND U25957 ( .A(n19184), .B(n19183), .Z(n19185) );
  NANDN U25958 ( .A(n19185), .B(n27567), .Z(n19186) );
  AND U25959 ( .A(n19187), .B(n19186), .Z(n19188) );
  OR U25960 ( .A(n19188), .B(n27569), .Z(n19189) );
  NAND U25961 ( .A(n27570), .B(n19189), .Z(n19190) );
  NANDN U25962 ( .A(n19191), .B(n19190), .Z(n19192) );
  ANDN U25963 ( .B(n27573), .A(n19192), .Z(n19193) );
  OR U25964 ( .A(n19194), .B(n19193), .Z(n19195) );
  AND U25965 ( .A(n19196), .B(n19195), .Z(n19197) );
  NANDN U25966 ( .A(n19198), .B(n19197), .Z(n19199) );
  NAND U25967 ( .A(n27577), .B(n19199), .Z(n19200) );
  NAND U25968 ( .A(n27578), .B(n19200), .Z(n19201) );
  AND U25969 ( .A(n27579), .B(n19201), .Z(n19204) );
  NAND U25970 ( .A(n19203), .B(n19202), .Z(n27580) );
  OR U25971 ( .A(n19204), .B(n27580), .Z(n19205) );
  AND U25972 ( .A(n27581), .B(n19205), .Z(n19208) );
  NAND U25973 ( .A(n19207), .B(n19206), .Z(n27582) );
  OR U25974 ( .A(n19208), .B(n27582), .Z(n19209) );
  NAND U25975 ( .A(n19210), .B(n19209), .Z(n19211) );
  NANDN U25976 ( .A(n19212), .B(n19211), .Z(n19213) );
  NAND U25977 ( .A(n19214), .B(n19213), .Z(n19215) );
  AND U25978 ( .A(n27587), .B(n19215), .Z(n19220) );
  NANDN U25979 ( .A(n19217), .B(n19216), .Z(n19218) );
  AND U25980 ( .A(n19219), .B(n19218), .Z(n27588) );
  NANDN U25981 ( .A(n19220), .B(n27588), .Z(n19221) );
  NAND U25982 ( .A(n27589), .B(n19221), .Z(n19222) );
  NANDN U25983 ( .A(n27590), .B(n19222), .Z(n19226) );
  IV U25984 ( .A(n19223), .Z(n27591) );
  AND U25985 ( .A(n19224), .B(n27591), .Z(n19225) );
  NAND U25986 ( .A(n19226), .B(n19225), .Z(n19227) );
  NANDN U25987 ( .A(n27592), .B(n19227), .Z(n19228) );
  OR U25988 ( .A(n19229), .B(n19228), .Z(n19230) );
  AND U25989 ( .A(n27594), .B(n19230), .Z(n19232) );
  NAND U25990 ( .A(n19232), .B(n19231), .Z(n19233) );
  NANDN U25991 ( .A(n19234), .B(n19233), .Z(n19235) );
  AND U25992 ( .A(n27596), .B(n19235), .Z(n19240) );
  NANDN U25993 ( .A(n19240), .B(n24269), .Z(n19241) );
  NAND U25994 ( .A(n27597), .B(n19241), .Z(n19242) );
  NANDN U25995 ( .A(n27598), .B(n19242), .Z(n19243) );
  AND U25996 ( .A(n27600), .B(n19243), .Z(n19244) );
  OR U25997 ( .A(n27601), .B(n19244), .Z(n19245) );
  NAND U25998 ( .A(n27602), .B(n19245), .Z(n19246) );
  NANDN U25999 ( .A(n19247), .B(n19246), .Z(n19248) );
  AND U26000 ( .A(n19248), .B(n27604), .Z(n19250) );
  NANDN U26001 ( .A(n19250), .B(n19249), .Z(n19251) );
  NANDN U26002 ( .A(n27605), .B(n19251), .Z(n19252) );
  AND U26003 ( .A(n27606), .B(n19252), .Z(n19253) );
  OR U26004 ( .A(n19254), .B(n19253), .Z(n19255) );
  NAND U26005 ( .A(n27608), .B(n19255), .Z(n19256) );
  NANDN U26006 ( .A(n19257), .B(n19256), .Z(n19258) );
  NAND U26007 ( .A(n27610), .B(n19258), .Z(n19259) );
  AND U26008 ( .A(n19260), .B(n19259), .Z(n19261) );
  NANDN U26009 ( .A(n19261), .B(n27612), .Z(n19262) );
  AND U26010 ( .A(n19263), .B(n19262), .Z(n19264) );
  OR U26011 ( .A(n27614), .B(n19264), .Z(n19265) );
  AND U26012 ( .A(n19265), .B(n27615), .Z(n19269) );
  NANDN U26013 ( .A(n19269), .B(n27617), .Z(n19270) );
  NAND U26014 ( .A(n24267), .B(n19270), .Z(n19271) );
  NANDN U26015 ( .A(n27618), .B(n19271), .Z(n19272) );
  NAND U26016 ( .A(n19273), .B(n19272), .Z(n19274) );
  NAND U26017 ( .A(n19275), .B(n19274), .Z(n19276) );
  NANDN U26018 ( .A(n27620), .B(n19276), .Z(n19278) );
  OR U26019 ( .A(n19278), .B(n19277), .Z(n19279) );
  AND U26020 ( .A(n19280), .B(n19279), .Z(n19283) );
  NAND U26021 ( .A(n19282), .B(n19281), .Z(n24264) );
  OR U26022 ( .A(n19283), .B(n24264), .Z(n19284) );
  AND U26023 ( .A(n27623), .B(n19284), .Z(n19285) );
  NANDN U26024 ( .A(n24265), .B(n19285), .Z(n19287) );
  AND U26025 ( .A(n19286), .B(n27622), .Z(n24263) );
  AND U26026 ( .A(n19287), .B(n24263), .Z(n19290) );
  NANDN U26027 ( .A(n19290), .B(n27624), .Z(n19291) );
  NAND U26028 ( .A(n27625), .B(n19291), .Z(n19292) );
  NANDN U26029 ( .A(n19293), .B(n19292), .Z(n19295) );
  AND U26030 ( .A(n27631), .B(n27627), .Z(n19294) );
  NAND U26031 ( .A(n19295), .B(n19294), .Z(n19296) );
  NANDN U26032 ( .A(n19297), .B(n19296), .Z(n19298) );
  OR U26033 ( .A(n19298), .B(n27632), .Z(n19299) );
  AND U26034 ( .A(n27633), .B(n19299), .Z(n19302) );
  NANDN U26035 ( .A(n19302), .B(n27634), .Z(n19303) );
  AND U26036 ( .A(n19304), .B(n19303), .Z(n19305) );
  NANDN U26037 ( .A(n27635), .B(n19305), .Z(n19306) );
  NAND U26038 ( .A(n19307), .B(n19306), .Z(n19308) );
  NANDN U26039 ( .A(n19309), .B(n19308), .Z(n19311) );
  OR U26040 ( .A(n19311), .B(n19310), .Z(n19312) );
  AND U26041 ( .A(n19313), .B(n19312), .Z(n19316) );
  NAND U26042 ( .A(n27641), .B(n19314), .Z(n19315) );
  OR U26043 ( .A(n19316), .B(n19315), .Z(n19321) );
  AND U26044 ( .A(n19321), .B(n27642), .Z(n19322) );
  OR U26045 ( .A(n27643), .B(n19322), .Z(n19323) );
  NAND U26046 ( .A(n27644), .B(n19323), .Z(n19324) );
  NANDN U26047 ( .A(n27645), .B(n19324), .Z(n19325) );
  NAND U26048 ( .A(n27646), .B(n19325), .Z(n19326) );
  NAND U26049 ( .A(n27647), .B(n19326), .Z(n19327) );
  NANDN U26050 ( .A(n19328), .B(n19327), .Z(n19329) );
  AND U26051 ( .A(n19330), .B(n19329), .Z(n19331) );
  OR U26052 ( .A(n19332), .B(n19331), .Z(n19333) );
  NAND U26053 ( .A(n19334), .B(n19333), .Z(n19335) );
  NANDN U26054 ( .A(n19336), .B(n19335), .Z(n19337) );
  OR U26055 ( .A(n19338), .B(n19337), .Z(n19339) );
  AND U26056 ( .A(n19339), .B(n27652), .Z(n19341) );
  OR U26057 ( .A(n19341), .B(n19340), .Z(n19342) );
  AND U26058 ( .A(n19342), .B(n24258), .Z(n19345) );
  NANDN U26059 ( .A(n19345), .B(n27653), .Z(n19346) );
  AND U26060 ( .A(n19347), .B(n19346), .Z(n19348) );
  NAND U26061 ( .A(n19348), .B(n27654), .Z(n19350) );
  ANDN U26062 ( .B(n19350), .A(n19349), .Z(n19351) );
  NANDN U26063 ( .A(n27655), .B(n19351), .Z(n19354) );
  ANDN U26064 ( .B(n27659), .A(n19352), .Z(n19353) );
  NAND U26065 ( .A(n19354), .B(n19353), .Z(n19359) );
  NANDN U26066 ( .A(n27660), .B(n19355), .Z(n19357) );
  ANDN U26067 ( .B(n19357), .A(n19356), .Z(n19358) );
  ANDN U26068 ( .B(n19359), .A(n19358), .Z(n19360) );
  NANDN U26069 ( .A(n19360), .B(n27661), .Z(n19361) );
  NAND U26070 ( .A(n27662), .B(n19361), .Z(n19362) );
  NANDN U26071 ( .A(n19363), .B(n19362), .Z(n19364) );
  NAND U26072 ( .A(n19365), .B(n19364), .Z(n19366) );
  AND U26073 ( .A(n19367), .B(n19366), .Z(n19368) );
  OR U26074 ( .A(n19369), .B(n19368), .Z(n19370) );
  NAND U26075 ( .A(n19371), .B(n19370), .Z(n19372) );
  AND U26076 ( .A(n19373), .B(n19372), .Z(n19377) );
  OR U26077 ( .A(n19377), .B(n24257), .Z(n19378) );
  NAND U26078 ( .A(n19379), .B(n19378), .Z(n19380) );
  NANDN U26079 ( .A(n27669), .B(n19380), .Z(n19383) );
  AND U26080 ( .A(n19381), .B(n27670), .Z(n19382) );
  NAND U26081 ( .A(n19383), .B(n19382), .Z(n19384) );
  NAND U26082 ( .A(n27671), .B(n19384), .Z(n19386) );
  AND U26083 ( .A(n19386), .B(n19385), .Z(n19387) );
  NANDN U26084 ( .A(n27672), .B(n19387), .Z(n19388) );
  NAND U26085 ( .A(n27674), .B(n19388), .Z(n19389) );
  NANDN U26086 ( .A(n19390), .B(n19389), .Z(n19391) );
  OR U26087 ( .A(n27677), .B(n19391), .Z(n19392) );
  AND U26088 ( .A(n27682), .B(n19392), .Z(n19393) );
  OR U26089 ( .A(n27684), .B(n19393), .Z(n19394) );
  NAND U26090 ( .A(n19395), .B(n19394), .Z(n19396) );
  NANDN U26091 ( .A(n19397), .B(n19396), .Z(n19399) );
  IV U26092 ( .A(n19398), .Z(n27687) );
  OR U26093 ( .A(n19399), .B(n27687), .Z(n19400) );
  NAND U26094 ( .A(n19401), .B(n19400), .Z(n19405) );
  IV U26095 ( .A(n19402), .Z(n27695) );
  AND U26096 ( .A(n19403), .B(n27695), .Z(n19404) );
  NAND U26097 ( .A(n19405), .B(n19404), .Z(n19406) );
  NANDN U26098 ( .A(n19407), .B(n19406), .Z(n19409) );
  IV U26099 ( .A(n19408), .Z(n27697) );
  OR U26100 ( .A(n19409), .B(n27697), .Z(n19410) );
  AND U26101 ( .A(n27700), .B(n19410), .Z(n19411) );
  OR U26102 ( .A(n27702), .B(n19411), .Z(n19412) );
  NAND U26103 ( .A(n27704), .B(n19412), .Z(n19413) );
  NANDN U26104 ( .A(n27706), .B(n19413), .Z(n19414) );
  NANDN U26105 ( .A(n27708), .B(n19414), .Z(n19415) );
  AND U26106 ( .A(n27710), .B(n19415), .Z(n19416) );
  OR U26107 ( .A(n27712), .B(n19416), .Z(n19417) );
  NAND U26108 ( .A(n27714), .B(n19417), .Z(n19418) );
  NANDN U26109 ( .A(n27716), .B(n19418), .Z(n19419) );
  AND U26110 ( .A(n27718), .B(n19419), .Z(n19422) );
  NAND U26111 ( .A(n19421), .B(n19420), .Z(n27719) );
  OR U26112 ( .A(n19422), .B(n27719), .Z(n19423) );
  NAND U26113 ( .A(n27721), .B(n19423), .Z(n19424) );
  NANDN U26114 ( .A(n19425), .B(n19424), .Z(n19426) );
  OR U26115 ( .A(n27722), .B(n19426), .Z(n19427) );
  AND U26116 ( .A(n27723), .B(n19427), .Z(n19428) );
  NAND U26117 ( .A(n19428), .B(n27725), .Z(n19430) );
  ANDN U26118 ( .B(n19430), .A(n19429), .Z(n19431) );
  NANDN U26119 ( .A(n27726), .B(n19431), .Z(n19432) );
  AND U26120 ( .A(n27727), .B(n19432), .Z(n19435) );
  NANDN U26121 ( .A(x[2356]), .B(y[2356]), .Z(n19434) );
  AND U26122 ( .A(n19434), .B(n19433), .Z(n27728) );
  NANDN U26123 ( .A(n19435), .B(n27728), .Z(n19436) );
  NAND U26124 ( .A(n27729), .B(n19436), .Z(n19437) );
  NANDN U26125 ( .A(n27730), .B(n19437), .Z(n19438) );
  AND U26126 ( .A(n19438), .B(n27731), .Z(n19440) );
  IV U26127 ( .A(n19439), .Z(n27732) );
  NANDN U26128 ( .A(n19440), .B(n27732), .Z(n19441) );
  NANDN U26129 ( .A(n27733), .B(n19441), .Z(n19442) );
  AND U26130 ( .A(n19443), .B(n19442), .Z(n19444) );
  OR U26131 ( .A(n19445), .B(n19444), .Z(n19446) );
  NAND U26132 ( .A(n19447), .B(n19446), .Z(n19448) );
  NANDN U26133 ( .A(n19449), .B(n19448), .Z(n19450) );
  OR U26134 ( .A(n24255), .B(n19450), .Z(n19451) );
  AND U26135 ( .A(n19452), .B(n19451), .Z(n19453) );
  NANDN U26136 ( .A(n27738), .B(n19453), .Z(n19454) );
  AND U26137 ( .A(n19455), .B(n19454), .Z(n19458) );
  NANDN U26138 ( .A(n19458), .B(n27740), .Z(n19459) );
  NAND U26139 ( .A(n27741), .B(n19459), .Z(n19460) );
  NAND U26140 ( .A(n27742), .B(n19460), .Z(n19461) );
  NAND U26141 ( .A(n24254), .B(n19461), .Z(n19462) );
  ANDN U26142 ( .B(n19462), .A(n24253), .Z(n19463) );
  NANDN U26143 ( .A(n19464), .B(n19463), .Z(n19466) );
  AND U26144 ( .A(n27743), .B(n27746), .Z(n19465) );
  NAND U26145 ( .A(n19466), .B(n19465), .Z(n19467) );
  NANDN U26146 ( .A(n19468), .B(n19467), .Z(n19469) );
  OR U26147 ( .A(n19469), .B(n27747), .Z(n19470) );
  NAND U26148 ( .A(n27748), .B(n19470), .Z(n19471) );
  NANDN U26149 ( .A(n19472), .B(n19471), .Z(n19474) );
  AND U26150 ( .A(n27750), .B(n27752), .Z(n19473) );
  NAND U26151 ( .A(n19474), .B(n19473), .Z(n19475) );
  NANDN U26152 ( .A(n19476), .B(n19475), .Z(n19478) );
  IV U26153 ( .A(n19477), .Z(n27753) );
  OR U26154 ( .A(n19478), .B(n27753), .Z(n19479) );
  AND U26155 ( .A(n27754), .B(n19479), .Z(n19482) );
  NAND U26156 ( .A(n19481), .B(n19480), .Z(n27755) );
  OR U26157 ( .A(n19482), .B(n27755), .Z(n19483) );
  AND U26158 ( .A(n19484), .B(n19483), .Z(n19485) );
  NANDN U26159 ( .A(n27756), .B(n19485), .Z(n19486) );
  AND U26160 ( .A(n27757), .B(n19486), .Z(n19487) );
  OR U26161 ( .A(n19488), .B(n19487), .Z(n19489) );
  NAND U26162 ( .A(n27759), .B(n19489), .Z(n19490) );
  NANDN U26163 ( .A(n19491), .B(n19490), .Z(n19492) );
  NAND U26164 ( .A(n19493), .B(n19492), .Z(n19494) );
  AND U26165 ( .A(n19495), .B(n19494), .Z(n19496) );
  OR U26166 ( .A(n19497), .B(n19496), .Z(n19498) );
  NAND U26167 ( .A(n19499), .B(n19498), .Z(n19500) );
  NANDN U26168 ( .A(n19501), .B(n19500), .Z(n19504) );
  AND U26169 ( .A(n19502), .B(n24252), .Z(n19503) );
  NAND U26170 ( .A(n19504), .B(n19503), .Z(n19505) );
  NANDN U26171 ( .A(n19506), .B(n19505), .Z(n19507) );
  OR U26172 ( .A(n19507), .B(n24251), .Z(n19508) );
  AND U26173 ( .A(n19508), .B(n24250), .Z(n19509) );
  ANDN U26174 ( .B(n19510), .A(n19509), .Z(n19511) );
  NAND U26175 ( .A(n27767), .B(n19511), .Z(n19512) );
  NANDN U26176 ( .A(n19513), .B(n19512), .Z(n19514) );
  OR U26177 ( .A(n27768), .B(n19514), .Z(n19515) );
  AND U26178 ( .A(n19516), .B(n19515), .Z(n19519) );
  NANDN U26179 ( .A(n19519), .B(y[2395]), .Z(n19518) );
  ANDN U26180 ( .B(n19518), .A(n19517), .Z(n19522) );
  XNOR U26181 ( .A(y[2395]), .B(n19519), .Z(n19520) );
  NANDN U26182 ( .A(x[2395]), .B(n19520), .Z(n19521) );
  NAND U26183 ( .A(n19522), .B(n19521), .Z(n19524) );
  IV U26184 ( .A(n19523), .Z(n27772) );
  AND U26185 ( .A(n19524), .B(n27772), .Z(n19525) );
  ANDN U26186 ( .B(n24249), .A(n19525), .Z(n19526) );
  OR U26187 ( .A(n19526), .B(n27773), .Z(n19527) );
  NAND U26188 ( .A(n27774), .B(n19527), .Z(n19528) );
  NANDN U26189 ( .A(n19529), .B(n19528), .Z(n19530) );
  OR U26190 ( .A(n19530), .B(n27775), .Z(n19531) );
  AND U26191 ( .A(n19531), .B(n27778), .Z(n19532) );
  ANDN U26192 ( .B(n19533), .A(n19532), .Z(n19534) );
  NANDN U26193 ( .A(n19535), .B(n19534), .Z(n19536) );
  AND U26194 ( .A(n19536), .B(n27781), .Z(n19537) );
  NANDN U26195 ( .A(n19537), .B(n27782), .Z(n19538) );
  NAND U26196 ( .A(n27784), .B(n19538), .Z(n19539) );
  AND U26197 ( .A(n27785), .B(n19539), .Z(n19540) );
  OR U26198 ( .A(n19541), .B(n19540), .Z(n19542) );
  NAND U26199 ( .A(n27789), .B(n19542), .Z(n19543) );
  NANDN U26200 ( .A(n27790), .B(n19543), .Z(n19544) );
  AND U26201 ( .A(n27791), .B(n19544), .Z(n19545) );
  OR U26202 ( .A(n27792), .B(n19545), .Z(n19546) );
  NAND U26203 ( .A(n27793), .B(n19546), .Z(n19547) );
  NANDN U26204 ( .A(n27794), .B(n19547), .Z(n19548) );
  AND U26205 ( .A(n27797), .B(n19548), .Z(n19550) );
  OR U26206 ( .A(n19550), .B(n19549), .Z(n19551) );
  AND U26207 ( .A(n27799), .B(n19551), .Z(n19552) );
  OR U26208 ( .A(n19552), .B(n27800), .Z(n19553) );
  AND U26209 ( .A(n19554), .B(n19553), .Z(n19559) );
  NAND U26210 ( .A(n19556), .B(n19555), .Z(n19557) );
  NAND U26211 ( .A(n19558), .B(n19557), .Z(n24246) );
  AND U26212 ( .A(n19559), .B(n24246), .Z(n19560) );
  OR U26213 ( .A(n19561), .B(n19560), .Z(n19562) );
  NAND U26214 ( .A(n19563), .B(n19562), .Z(n19564) );
  NANDN U26215 ( .A(n27803), .B(n19564), .Z(n19566) );
  OR U26216 ( .A(n19566), .B(n19565), .Z(n19567) );
  AND U26217 ( .A(n19568), .B(n19567), .Z(n19569) );
  OR U26218 ( .A(n27805), .B(n19569), .Z(n19570) );
  NAND U26219 ( .A(n19571), .B(n19570), .Z(n19572) );
  NANDN U26220 ( .A(n27807), .B(n19572), .Z(n19573) );
  OR U26221 ( .A(n19573), .B(n27810), .Z(n19574) );
  AND U26222 ( .A(n19575), .B(n19574), .Z(n19576) );
  OR U26223 ( .A(n27812), .B(n19576), .Z(n19577) );
  NAND U26224 ( .A(n27813), .B(n19577), .Z(n19578) );
  NANDN U26225 ( .A(n27814), .B(n19578), .Z(n19579) );
  NAND U26226 ( .A(n27815), .B(n19579), .Z(n19580) );
  NANDN U26227 ( .A(n27816), .B(n19580), .Z(n19581) );
  AND U26228 ( .A(n24243), .B(n19581), .Z(n19582) );
  OR U26229 ( .A(n19583), .B(n19582), .Z(n19584) );
  AND U26230 ( .A(n19585), .B(n19584), .Z(n19586) );
  NAND U26231 ( .A(n19586), .B(n24244), .Z(n19588) );
  ANDN U26232 ( .B(n19588), .A(n19587), .Z(n19589) );
  NANDN U26233 ( .A(n19590), .B(n19589), .Z(n19591) );
  AND U26234 ( .A(n19592), .B(n19591), .Z(n19595) );
  NAND U26235 ( .A(n19594), .B(n19593), .Z(n27818) );
  OR U26236 ( .A(n19595), .B(n27818), .Z(n19596) );
  AND U26237 ( .A(n27819), .B(n19596), .Z(n19600) );
  OR U26238 ( .A(n19600), .B(n27820), .Z(n19602) );
  IV U26239 ( .A(n19601), .Z(n27821) );
  AND U26240 ( .A(n19602), .B(n27821), .Z(n19604) );
  IV U26241 ( .A(n19603), .Z(n27822) );
  OR U26242 ( .A(n19604), .B(n27822), .Z(n19605) );
  NAND U26243 ( .A(n19606), .B(n19605), .Z(n19607) );
  NANDN U26244 ( .A(n19608), .B(n19607), .Z(n19611) );
  AND U26245 ( .A(n19609), .B(n27825), .Z(n19610) );
  NAND U26246 ( .A(n19611), .B(n19610), .Z(n19612) );
  NANDN U26247 ( .A(n19613), .B(n19612), .Z(n19615) );
  OR U26248 ( .A(n19615), .B(n19614), .Z(n19616) );
  NAND U26249 ( .A(n19617), .B(n19616), .Z(n19618) );
  NANDN U26250 ( .A(n19619), .B(n19618), .Z(n19621) );
  OR U26251 ( .A(n19621), .B(n19620), .Z(n19622) );
  AND U26252 ( .A(n19623), .B(n19622), .Z(n19624) );
  OR U26253 ( .A(n19625), .B(n19624), .Z(n19626) );
  NAND U26254 ( .A(n27833), .B(n19626), .Z(n19627) );
  NANDN U26255 ( .A(n19628), .B(n19627), .Z(n19630) );
  IV U26256 ( .A(n19629), .Z(n27834) );
  OR U26257 ( .A(n19630), .B(n27834), .Z(n19631) );
  NAND U26258 ( .A(n27835), .B(n19631), .Z(n19632) );
  AND U26259 ( .A(n19633), .B(n19632), .Z(n19634) );
  NAND U26260 ( .A(n19634), .B(n27836), .Z(n19635) );
  NANDN U26261 ( .A(n27837), .B(n19635), .Z(n19636) );
  AND U26262 ( .A(n19637), .B(n19636), .Z(n19638) );
  NOR U26263 ( .A(n27840), .B(n19638), .Z(n19639) );
  NANDN U26264 ( .A(n19640), .B(n19639), .Z(n19641) );
  AND U26265 ( .A(n19642), .B(n19641), .Z(n19643) );
  NAND U26266 ( .A(n27842), .B(n19643), .Z(n19645) );
  ANDN U26267 ( .B(n19645), .A(n19644), .Z(n19646) );
  NANDN U26268 ( .A(n27843), .B(n19646), .Z(n19647) );
  AND U26269 ( .A(n27844), .B(n19647), .Z(n19649) );
  IV U26270 ( .A(n19648), .Z(n27845) );
  OR U26271 ( .A(n19649), .B(n27845), .Z(n19650) );
  NAND U26272 ( .A(n27846), .B(n19650), .Z(n19651) );
  NANDN U26273 ( .A(n19652), .B(n19651), .Z(n19654) );
  IV U26274 ( .A(n19653), .Z(n27847) );
  OR U26275 ( .A(n19654), .B(n27847), .Z(n19655) );
  NAND U26276 ( .A(n27848), .B(n19655), .Z(n19656) );
  NANDN U26277 ( .A(n19657), .B(n19656), .Z(n19658) );
  NAND U26278 ( .A(n27852), .B(n19658), .Z(n19659) );
  NANDN U26279 ( .A(n27853), .B(n19659), .Z(n19660) );
  AND U26280 ( .A(n27854), .B(n19660), .Z(n19661) );
  OR U26281 ( .A(n19661), .B(n27855), .Z(n19662) );
  AND U26282 ( .A(n27856), .B(n19662), .Z(n19663) );
  OR U26283 ( .A(n27858), .B(n19663), .Z(n19664) );
  AND U26284 ( .A(n19665), .B(n19664), .Z(n19666) );
  OR U26285 ( .A(n27860), .B(n19666), .Z(n19667) );
  NAND U26286 ( .A(n27864), .B(n19667), .Z(n19668) );
  NANDN U26287 ( .A(n27865), .B(n19668), .Z(n19671) );
  AND U26288 ( .A(n19669), .B(n27866), .Z(n19670) );
  NAND U26289 ( .A(n19671), .B(n19670), .Z(n19672) );
  NANDN U26290 ( .A(n19673), .B(n19672), .Z(n19674) );
  OR U26291 ( .A(n19674), .B(n27867), .Z(n19675) );
  AND U26292 ( .A(n19676), .B(n19675), .Z(n19677) );
  OR U26293 ( .A(n19678), .B(n19677), .Z(n19679) );
  NAND U26294 ( .A(n27872), .B(n19679), .Z(n19680) );
  NANDN U26295 ( .A(n19681), .B(n19680), .Z(n19683) );
  IV U26296 ( .A(n19682), .Z(n27873) );
  OR U26297 ( .A(n19683), .B(n27873), .Z(n19684) );
  NANDN U26298 ( .A(n19685), .B(n19684), .Z(n19686) );
  AND U26299 ( .A(n19687), .B(n19686), .Z(n19688) );
  OR U26300 ( .A(n19689), .B(n19688), .Z(n19690) );
  NAND U26301 ( .A(n19691), .B(n19690), .Z(n19692) );
  NANDN U26302 ( .A(n27882), .B(n19692), .Z(n19693) );
  OR U26303 ( .A(n19694), .B(n19693), .Z(n19695) );
  AND U26304 ( .A(n19696), .B(n19695), .Z(n19697) );
  ANDN U26305 ( .B(n19698), .A(n19697), .Z(n19699) );
  NANDN U26306 ( .A(n19700), .B(n19699), .Z(n19701) );
  AND U26307 ( .A(n27885), .B(n19701), .Z(n19703) );
  AND U26308 ( .A(n19703), .B(n19702), .Z(n19709) );
  OR U26309 ( .A(n19705), .B(n19704), .Z(n19706) );
  AND U26310 ( .A(n19707), .B(n19706), .Z(n19708) );
  NOR U26311 ( .A(n19709), .B(n19708), .Z(n19710) );
  NAND U26312 ( .A(n19711), .B(n19710), .Z(n19712) );
  NAND U26313 ( .A(n27887), .B(n19712), .Z(n19713) );
  AND U26314 ( .A(n27888), .B(n19713), .Z(n19714) );
  OR U26315 ( .A(n27889), .B(n19714), .Z(n19715) );
  NAND U26316 ( .A(n27890), .B(n19715), .Z(n19716) );
  NANDN U26317 ( .A(n27891), .B(n19716), .Z(n19719) );
  AND U26318 ( .A(n19717), .B(n27892), .Z(n19718) );
  NAND U26319 ( .A(n19719), .B(n19718), .Z(n19720) );
  NANDN U26320 ( .A(n19721), .B(n19720), .Z(n19723) );
  IV U26321 ( .A(n19722), .Z(n27893) );
  OR U26322 ( .A(n19723), .B(n27893), .Z(n19724) );
  AND U26323 ( .A(n19725), .B(n19724), .Z(n19726) );
  NANDN U26324 ( .A(n27896), .B(n19726), .Z(n19727) );
  AND U26325 ( .A(n19728), .B(n19727), .Z(n19731) );
  NAND U26326 ( .A(n19730), .B(n19729), .Z(n27899) );
  OR U26327 ( .A(n19731), .B(n27899), .Z(n19732) );
  NAND U26328 ( .A(n19733), .B(n19732), .Z(n19734) );
  NANDN U26329 ( .A(n19735), .B(n19734), .Z(n19736) );
  OR U26330 ( .A(n19736), .B(n27901), .Z(n19737) );
  AND U26331 ( .A(n19738), .B(n19737), .Z(n19739) );
  NOR U26332 ( .A(n19739), .B(n27905), .Z(n19740) );
  NANDN U26333 ( .A(n19741), .B(n19740), .Z(n19742) );
  AND U26334 ( .A(n27906), .B(n19742), .Z(n19743) );
  NANDN U26335 ( .A(n19744), .B(n19743), .Z(n19745) );
  NAND U26336 ( .A(n27907), .B(n19745), .Z(n19746) );
  NANDN U26337 ( .A(n27908), .B(n19746), .Z(n19747) );
  NAND U26338 ( .A(n27909), .B(n19747), .Z(n19748) );
  NAND U26339 ( .A(n19749), .B(n19748), .Z(n19750) );
  NANDN U26340 ( .A(n19751), .B(n19750), .Z(n19754) );
  AND U26341 ( .A(n19752), .B(n24235), .Z(n19753) );
  NAND U26342 ( .A(n19754), .B(n19753), .Z(n19755) );
  NANDN U26343 ( .A(n19756), .B(n19755), .Z(n19757) );
  OR U26344 ( .A(n19757), .B(n24234), .Z(n19758) );
  AND U26345 ( .A(n27912), .B(n19758), .Z(n19759) );
  OR U26346 ( .A(n19760), .B(n19759), .Z(n19761) );
  NAND U26347 ( .A(n27913), .B(n19761), .Z(n19762) );
  NANDN U26348 ( .A(n19763), .B(n19762), .Z(n19764) );
  OR U26349 ( .A(n27914), .B(n19764), .Z(n19765) );
  AND U26350 ( .A(n19765), .B(n24230), .Z(n19766) );
  NANDN U26351 ( .A(n19767), .B(n19766), .Z(n19768) );
  NAND U26352 ( .A(n19769), .B(n19768), .Z(n19770) );
  NANDN U26353 ( .A(n19771), .B(n19770), .Z(n19772) );
  AND U26354 ( .A(n19773), .B(n19772), .Z(n19774) );
  OR U26355 ( .A(n19775), .B(n19774), .Z(n19776) );
  NAND U26356 ( .A(n19777), .B(n19776), .Z(n19778) );
  NANDN U26357 ( .A(n19779), .B(n19778), .Z(n19780) );
  OR U26358 ( .A(n19781), .B(n19780), .Z(n19782) );
  AND U26359 ( .A(n19783), .B(n19782), .Z(n19784) );
  NAND U26360 ( .A(n24229), .B(n19784), .Z(n19786) );
  ANDN U26361 ( .B(n19786), .A(n19785), .Z(n19787) );
  NANDN U26362 ( .A(n19788), .B(n19787), .Z(n19791) );
  AND U26363 ( .A(n19789), .B(n27925), .Z(n19790) );
  NAND U26364 ( .A(n19791), .B(n19790), .Z(n19792) );
  NANDN U26365 ( .A(n19793), .B(n19792), .Z(n19794) );
  OR U26366 ( .A(n19794), .B(n27926), .Z(n19795) );
  NAND U26367 ( .A(n24228), .B(n19795), .Z(n19796) );
  NANDN U26368 ( .A(n19797), .B(n19796), .Z(n19798) );
  NAND U26369 ( .A(n27927), .B(n19798), .Z(n19799) );
  AND U26370 ( .A(n19800), .B(n19799), .Z(n19801) );
  OR U26371 ( .A(n19802), .B(n19801), .Z(n19803) );
  NAND U26372 ( .A(n19804), .B(n19803), .Z(n19805) );
  NANDN U26373 ( .A(n19806), .B(n19805), .Z(n19810) );
  AND U26374 ( .A(n19808), .B(n19807), .Z(n19809) );
  NAND U26375 ( .A(n19810), .B(n19809), .Z(n19811) );
  NANDN U26376 ( .A(n19812), .B(n19811), .Z(n19813) );
  OR U26377 ( .A(n19814), .B(n19813), .Z(n19815) );
  AND U26378 ( .A(n19816), .B(n19815), .Z(n19817) );
  NANDN U26379 ( .A(n27935), .B(n19817), .Z(n19818) );
  AND U26380 ( .A(n19819), .B(n19818), .Z(n19822) );
  NAND U26381 ( .A(n19821), .B(n19820), .Z(n27937) );
  OR U26382 ( .A(n19822), .B(n27937), .Z(n19823) );
  AND U26383 ( .A(n19824), .B(n19823), .Z(n19825) );
  NAND U26384 ( .A(n27938), .B(n19825), .Z(n19826) );
  NANDN U26385 ( .A(n27939), .B(n19826), .Z(n19827) );
  AND U26386 ( .A(n19828), .B(n19827), .Z(n19829) );
  OR U26387 ( .A(n27943), .B(n19829), .Z(n19830) );
  NAND U26388 ( .A(n27944), .B(n19830), .Z(n19831) );
  NANDN U26389 ( .A(n19832), .B(n19831), .Z(n19835) );
  AND U26390 ( .A(n19833), .B(n27946), .Z(n19834) );
  NAND U26391 ( .A(n19835), .B(n19834), .Z(n19836) );
  NANDN U26392 ( .A(n19837), .B(n19836), .Z(n19839) );
  OR U26393 ( .A(n19839), .B(n19838), .Z(n19840) );
  NAND U26394 ( .A(n19841), .B(n19840), .Z(n19842) );
  NANDN U26395 ( .A(n27951), .B(n19842), .Z(n19844) );
  OR U26396 ( .A(n19844), .B(n19843), .Z(n19845) );
  NAND U26397 ( .A(n27953), .B(n19845), .Z(n19846) );
  NANDN U26398 ( .A(n27957), .B(n19846), .Z(n19847) );
  NANDN U26399 ( .A(n19847), .B(n27954), .Z(n19848) );
  AND U26400 ( .A(n27955), .B(n19848), .Z(n19849) );
  OR U26401 ( .A(n27959), .B(n19849), .Z(n19850) );
  NAND U26402 ( .A(n27960), .B(n19850), .Z(n19851) );
  NANDN U26403 ( .A(n27961), .B(n19851), .Z(n19852) );
  NAND U26404 ( .A(n27962), .B(n19852), .Z(n19855) );
  AND U26405 ( .A(n19854), .B(n19853), .Z(n24225) );
  AND U26406 ( .A(n19855), .B(n24225), .Z(n19858) );
  IV U26407 ( .A(n19856), .Z(n27963) );
  AND U26408 ( .A(n24223), .B(n27963), .Z(n19857) );
  NANDN U26409 ( .A(n19858), .B(n19857), .Z(n19859) );
  NANDN U26410 ( .A(n27964), .B(n19859), .Z(n19860) );
  AND U26411 ( .A(n24224), .B(n19860), .Z(n19863) );
  OR U26412 ( .A(n19863), .B(n27965), .Z(n19864) );
  AND U26413 ( .A(n19864), .B(n24221), .Z(n19865) );
  NANDN U26414 ( .A(n27966), .B(n19865), .Z(n19866) );
  AND U26415 ( .A(n19867), .B(n19866), .Z(n19868) );
  OR U26416 ( .A(n27971), .B(n19868), .Z(n19869) );
  NAND U26417 ( .A(n27972), .B(n19869), .Z(n19870) );
  NANDN U26418 ( .A(n27973), .B(n19870), .Z(n19871) );
  NAND U26419 ( .A(n27974), .B(n19871), .Z(n19872) );
  NANDN U26420 ( .A(n24220), .B(n19872), .Z(n19875) );
  AND U26421 ( .A(n19874), .B(n19873), .Z(n27975) );
  ANDN U26422 ( .B(n19875), .A(n27975), .Z(n19876) );
  OR U26423 ( .A(n19877), .B(n19876), .Z(n19878) );
  NAND U26424 ( .A(n19879), .B(n19878), .Z(n19880) );
  NANDN U26425 ( .A(n19881), .B(n19880), .Z(n19882) );
  AND U26426 ( .A(n19883), .B(n19882), .Z(n19884) );
  NAND U26427 ( .A(n27976), .B(n19884), .Z(n19888) );
  NAND U26428 ( .A(n19886), .B(n19885), .Z(n19887) );
  ANDN U26429 ( .B(n19888), .A(n19887), .Z(n19892) );
  NAND U26430 ( .A(n19890), .B(n19889), .Z(n19891) );
  OR U26431 ( .A(n19892), .B(n19891), .Z(n19893) );
  AND U26432 ( .A(n19894), .B(n19893), .Z(n19898) );
  NAND U26433 ( .A(n19896), .B(n19895), .Z(n19897) );
  OR U26434 ( .A(n19898), .B(n19897), .Z(n19899) );
  AND U26435 ( .A(n19900), .B(n19899), .Z(n19901) );
  OR U26436 ( .A(n19902), .B(n19901), .Z(n19903) );
  NAND U26437 ( .A(n19904), .B(n19903), .Z(n19907) );
  AND U26438 ( .A(n19905), .B(n24217), .Z(n19906) );
  NAND U26439 ( .A(n19907), .B(n19906), .Z(n19908) );
  NANDN U26440 ( .A(n19909), .B(n19908), .Z(n19911) );
  OR U26441 ( .A(n19911), .B(n19910), .Z(n19912) );
  NAND U26442 ( .A(n27986), .B(n19912), .Z(n19913) );
  NANDN U26443 ( .A(n19914), .B(n19913), .Z(n19917) );
  AND U26444 ( .A(n19915), .B(n27988), .Z(n19916) );
  NAND U26445 ( .A(n19917), .B(n19916), .Z(n19918) );
  NANDN U26446 ( .A(n19919), .B(n19918), .Z(n19921) );
  OR U26447 ( .A(n19921), .B(n19920), .Z(n19922) );
  NAND U26448 ( .A(n19923), .B(n19922), .Z(n19924) );
  NAND U26449 ( .A(n24214), .B(n19924), .Z(n19927) );
  AND U26450 ( .A(n19925), .B(n24213), .Z(n19926) );
  NAND U26451 ( .A(n19927), .B(n19926), .Z(n19928) );
  NANDN U26452 ( .A(n19929), .B(n19928), .Z(n19930) );
  OR U26453 ( .A(n19931), .B(n19930), .Z(n19932) );
  AND U26454 ( .A(n19933), .B(n19932), .Z(n19934) );
  NAND U26455 ( .A(n19935), .B(n19934), .Z(n19936) );
  NAND U26456 ( .A(n19937), .B(n19936), .Z(n19938) );
  AND U26457 ( .A(n19939), .B(n19938), .Z(n19940) );
  OR U26458 ( .A(n27995), .B(n19940), .Z(n19942) );
  IV U26459 ( .A(n19941), .Z(n27996) );
  AND U26460 ( .A(n19942), .B(n27996), .Z(n19945) );
  AND U26461 ( .A(n19944), .B(n19943), .Z(n24212) );
  NANDN U26462 ( .A(n19945), .B(n24212), .Z(n19946) );
  NAND U26463 ( .A(n19947), .B(n19946), .Z(n19950) );
  AND U26464 ( .A(n19948), .B(n24210), .Z(n19949) );
  NAND U26465 ( .A(n19950), .B(n19949), .Z(n19951) );
  NANDN U26466 ( .A(n19952), .B(n19951), .Z(n19953) );
  OR U26467 ( .A(n19954), .B(n19953), .Z(n19955) );
  AND U26468 ( .A(n19956), .B(n19955), .Z(n19957) );
  NANDN U26469 ( .A(n19958), .B(n19957), .Z(n19959) );
  AND U26470 ( .A(n19960), .B(n19959), .Z(n19961) );
  OR U26471 ( .A(n19962), .B(n19961), .Z(n19963) );
  NAND U26472 ( .A(n24208), .B(n19963), .Z(n19964) );
  NANDN U26473 ( .A(n19965), .B(n19964), .Z(n19967) );
  IV U26474 ( .A(n19966), .Z(n24207) );
  OR U26475 ( .A(n19967), .B(n24207), .Z(n19968) );
  AND U26476 ( .A(n24209), .B(n19968), .Z(n19969) );
  OR U26477 ( .A(n19970), .B(n19969), .Z(n19971) );
  NAND U26478 ( .A(n28008), .B(n19971), .Z(n19972) );
  NANDN U26479 ( .A(n19973), .B(n19972), .Z(n19974) );
  ANDN U26480 ( .B(y[2616]), .A(x[2616]), .Z(n28009) );
  OR U26481 ( .A(n19974), .B(n28009), .Z(n19975) );
  NAND U26482 ( .A(n19976), .B(n19975), .Z(n19979) );
  AND U26483 ( .A(n19977), .B(n28013), .Z(n19978) );
  NAND U26484 ( .A(n19979), .B(n19978), .Z(n19980) );
  NANDN U26485 ( .A(n19981), .B(n19980), .Z(n19982) );
  OR U26486 ( .A(n28014), .B(n19982), .Z(n19983) );
  AND U26487 ( .A(n28015), .B(n19983), .Z(n19984) );
  ANDN U26488 ( .B(n19985), .A(n19984), .Z(n19986) );
  NAND U26489 ( .A(n28016), .B(n19986), .Z(n19987) );
  NANDN U26490 ( .A(n28017), .B(n19987), .Z(n19988) );
  OR U26491 ( .A(n19989), .B(n19988), .Z(n19990) );
  AND U26492 ( .A(n19991), .B(n19990), .Z(n19992) );
  NAND U26493 ( .A(n19993), .B(n19992), .Z(n19994) );
  NAND U26494 ( .A(n19995), .B(n19994), .Z(n19996) );
  AND U26495 ( .A(n19997), .B(n19996), .Z(n19998) );
  OR U26496 ( .A(n19999), .B(n19998), .Z(n20000) );
  AND U26497 ( .A(n28023), .B(n20000), .Z(n20001) );
  OR U26498 ( .A(n20001), .B(n28026), .Z(n20002) );
  AND U26499 ( .A(n28029), .B(n20002), .Z(n20003) );
  OR U26500 ( .A(n20003), .B(n28030), .Z(n20004) );
  AND U26501 ( .A(n20005), .B(n20004), .Z(n20006) );
  NAND U26502 ( .A(n20006), .B(y[2631]), .Z(n20009) );
  XOR U26503 ( .A(n20006), .B(y[2631]), .Z(n20007) );
  NANDN U26504 ( .A(x[2631]), .B(n20007), .Z(n20008) );
  NAND U26505 ( .A(n20009), .B(n20008), .Z(n20010) );
  AND U26506 ( .A(n20010), .B(n24206), .Z(n20011) );
  OR U26507 ( .A(n20012), .B(n20011), .Z(n20013) );
  NAND U26508 ( .A(n28034), .B(n20013), .Z(n20014) );
  NANDN U26509 ( .A(n20015), .B(n20014), .Z(n20016) );
  OR U26510 ( .A(n20016), .B(n28035), .Z(n20017) );
  AND U26511 ( .A(n28036), .B(n20017), .Z(n20018) );
  ANDN U26512 ( .B(n20019), .A(n20018), .Z(n20020) );
  NAND U26513 ( .A(n20021), .B(n20020), .Z(n20022) );
  NANDN U26514 ( .A(n28039), .B(n20022), .Z(n20024) );
  OR U26515 ( .A(n20024), .B(n20023), .Z(n20025) );
  AND U26516 ( .A(n20026), .B(n20025), .Z(n20027) );
  NOR U26517 ( .A(n28042), .B(n20027), .Z(n20028) );
  NANDN U26518 ( .A(n20029), .B(n20028), .Z(n20030) );
  AND U26519 ( .A(n20030), .B(n28043), .Z(n20032) );
  AND U26520 ( .A(n20032), .B(n20031), .Z(n20035) );
  XNOR U26521 ( .A(y[2642]), .B(x[2642]), .Z(n20033) );
  NANDN U26522 ( .A(n20034), .B(n20033), .Z(n24201) );
  OR U26523 ( .A(n20035), .B(n24201), .Z(n20036) );
  AND U26524 ( .A(n28044), .B(n20036), .Z(n20037) );
  OR U26525 ( .A(n28045), .B(n20037), .Z(n20038) );
  NAND U26526 ( .A(n28046), .B(n20038), .Z(n20039) );
  NANDN U26527 ( .A(n28047), .B(n20039), .Z(n20040) );
  AND U26528 ( .A(n28048), .B(n20040), .Z(n20041) );
  NANDN U26529 ( .A(n20041), .B(n28049), .Z(n20042) );
  NAND U26530 ( .A(n28050), .B(n20042), .Z(n20043) );
  NANDN U26531 ( .A(n28051), .B(n20043), .Z(n20044) );
  AND U26532 ( .A(n28052), .B(n20044), .Z(n20045) );
  OR U26533 ( .A(n20045), .B(n28053), .Z(n20046) );
  NANDN U26534 ( .A(n28055), .B(n20046), .Z(n20047) );
  AND U26535 ( .A(n28056), .B(n20047), .Z(n20048) );
  OR U26536 ( .A(n28057), .B(n20048), .Z(n20049) );
  NAND U26537 ( .A(n28058), .B(n20049), .Z(n20050) );
  NANDN U26538 ( .A(n20051), .B(n20050), .Z(n20054) );
  IV U26539 ( .A(n20052), .Z(n28060) );
  AND U26540 ( .A(n28062), .B(n28060), .Z(n20053) );
  NAND U26541 ( .A(n20054), .B(n20053), .Z(n20055) );
  NANDN U26542 ( .A(n20056), .B(n20055), .Z(n20057) );
  OR U26543 ( .A(n28063), .B(n20057), .Z(n20058) );
  AND U26544 ( .A(n28064), .B(n20058), .Z(n20059) );
  OR U26545 ( .A(n20060), .B(n20059), .Z(n20061) );
  NAND U26546 ( .A(n20062), .B(n20061), .Z(n20063) );
  NANDN U26547 ( .A(n28068), .B(n20063), .Z(n20064) );
  OR U26548 ( .A(n20065), .B(n20064), .Z(n20066) );
  AND U26549 ( .A(n28069), .B(n20066), .Z(n20067) );
  OR U26550 ( .A(n28070), .B(n20067), .Z(n20068) );
  NAND U26551 ( .A(n20069), .B(n20068), .Z(n20070) );
  NANDN U26552 ( .A(n20071), .B(n20070), .Z(n20073) );
  IV U26553 ( .A(n20072), .Z(n28072) );
  OR U26554 ( .A(n20073), .B(n28072), .Z(n20074) );
  AND U26555 ( .A(n20075), .B(n20074), .Z(n20076) );
  ANDN U26556 ( .B(n28077), .A(n20076), .Z(n20077) );
  NANDN U26557 ( .A(n20078), .B(n20077), .Z(n20079) );
  AND U26558 ( .A(n28078), .B(n20079), .Z(n20080) );
  NANDN U26559 ( .A(n20081), .B(n20080), .Z(n20082) );
  AND U26560 ( .A(n20083), .B(n20082), .Z(n20084) );
  NANDN U26561 ( .A(n28079), .B(n20084), .Z(n20085) );
  NAND U26562 ( .A(n20086), .B(n20085), .Z(n20087) );
  NANDN U26563 ( .A(n20088), .B(n20087), .Z(n20092) );
  AND U26564 ( .A(n20090), .B(n20089), .Z(n20091) );
  NAND U26565 ( .A(n20092), .B(n20091), .Z(n20093) );
  NANDN U26566 ( .A(n20094), .B(n20093), .Z(n20096) );
  OR U26567 ( .A(n20096), .B(n20095), .Z(n20097) );
  NAND U26568 ( .A(n20098), .B(n20097), .Z(n20099) );
  NANDN U26569 ( .A(n20100), .B(n20099), .Z(n20101) );
  OR U26570 ( .A(n20102), .B(n20101), .Z(n20103) );
  AND U26571 ( .A(n20104), .B(n20103), .Z(n20106) );
  NAND U26572 ( .A(n20106), .B(n20105), .Z(n20108) );
  ANDN U26573 ( .B(n20108), .A(n20107), .Z(n20109) );
  NANDN U26574 ( .A(n20110), .B(n20109), .Z(n20113) );
  AND U26575 ( .A(n20111), .B(n28088), .Z(n20112) );
  NAND U26576 ( .A(n20113), .B(n20112), .Z(n20114) );
  NANDN U26577 ( .A(n20115), .B(n20114), .Z(n20116) );
  OR U26578 ( .A(n28090), .B(n20116), .Z(n20117) );
  AND U26579 ( .A(n28091), .B(n20117), .Z(n20120) );
  NANDN U26580 ( .A(x[2682]), .B(y[2682]), .Z(n20119) );
  NAND U26581 ( .A(n20119), .B(n20118), .Z(n28092) );
  OR U26582 ( .A(n20120), .B(n28092), .Z(n20121) );
  NAND U26583 ( .A(n28093), .B(n20121), .Z(n20122) );
  NAND U26584 ( .A(n28094), .B(n20122), .Z(n20123) );
  NAND U26585 ( .A(n24198), .B(n20123), .Z(n20124) );
  NANDN U26586 ( .A(n24197), .B(n20124), .Z(n20125) );
  AND U26587 ( .A(n20126), .B(n20125), .Z(n20127) );
  OR U26588 ( .A(n20128), .B(n20127), .Z(n20129) );
  NAND U26589 ( .A(n20130), .B(n20129), .Z(n20131) );
  NANDN U26590 ( .A(n28098), .B(n20131), .Z(n20132) );
  OR U26591 ( .A(n20132), .B(n28100), .Z(n20133) );
  NAND U26592 ( .A(n20134), .B(n20133), .Z(n20135) );
  NAND U26593 ( .A(n28102), .B(n20135), .Z(n20136) );
  AND U26594 ( .A(n20137), .B(n20136), .Z(n20138) );
  OR U26595 ( .A(n20139), .B(n20138), .Z(n20140) );
  NAND U26596 ( .A(n20141), .B(n20140), .Z(n20145) );
  AND U26597 ( .A(n20143), .B(n20142), .Z(n20144) );
  NAND U26598 ( .A(n20145), .B(n20144), .Z(n20146) );
  NANDN U26599 ( .A(n28109), .B(n20146), .Z(n20148) );
  OR U26600 ( .A(n20148), .B(n20147), .Z(n20149) );
  NAND U26601 ( .A(n20150), .B(n20149), .Z(n20151) );
  NANDN U26602 ( .A(n28111), .B(n20151), .Z(n20153) );
  AND U26603 ( .A(n20153), .B(n20152), .Z(n20154) );
  NANDN U26604 ( .A(x[2700]), .B(y[2700]), .Z(n28112) );
  AND U26605 ( .A(n20154), .B(n28112), .Z(n20155) );
  OR U26606 ( .A(n28113), .B(n20155), .Z(n20156) );
  NAND U26607 ( .A(n20157), .B(n20156), .Z(n20158) );
  NANDN U26608 ( .A(n28114), .B(n20158), .Z(n20160) );
  AND U26609 ( .A(n20160), .B(n20159), .Z(n20161) );
  NANDN U26610 ( .A(n28115), .B(n20161), .Z(n20162) );
  NAND U26611 ( .A(n28116), .B(n20162), .Z(n20163) );
  NANDN U26612 ( .A(n20164), .B(n20163), .Z(n20165) );
  OR U26613 ( .A(n20165), .B(n24191), .Z(n20166) );
  AND U26614 ( .A(n28118), .B(n20166), .Z(n20168) );
  NANDN U26615 ( .A(n20168), .B(n28119), .Z(n20169) );
  NAND U26616 ( .A(n24187), .B(n20169), .Z(n20170) );
  NANDN U26617 ( .A(n24186), .B(n20170), .Z(n20174) );
  AND U26618 ( .A(n28120), .B(n28121), .Z(n20173) );
  NAND U26619 ( .A(n20174), .B(n20173), .Z(n20175) );
  NANDN U26620 ( .A(n28122), .B(n20175), .Z(n20178) );
  AND U26621 ( .A(n28123), .B(n20176), .Z(n20177) );
  NAND U26622 ( .A(n20178), .B(n20177), .Z(n20179) );
  NANDN U26623 ( .A(n28124), .B(n20179), .Z(n20183) );
  AND U26624 ( .A(n20181), .B(n20180), .Z(n20182) );
  NAND U26625 ( .A(n20183), .B(n20182), .Z(n20184) );
  NANDN U26626 ( .A(n28126), .B(n20184), .Z(n20186) );
  OR U26627 ( .A(n20186), .B(n20185), .Z(n20187) );
  NAND U26628 ( .A(n20188), .B(n20187), .Z(n20189) );
  NANDN U26629 ( .A(n20190), .B(n20189), .Z(n20192) );
  OR U26630 ( .A(n20192), .B(n20191), .Z(n20193) );
  NAND U26631 ( .A(n20194), .B(n20193), .Z(n20197) );
  AND U26632 ( .A(n20195), .B(n28132), .Z(n20196) );
  NAND U26633 ( .A(n20197), .B(n20196), .Z(n20198) );
  NANDN U26634 ( .A(n20199), .B(n20198), .Z(n20201) );
  IV U26635 ( .A(n20200), .Z(n28136) );
  OR U26636 ( .A(n20201), .B(n28136), .Z(n20202) );
  AND U26637 ( .A(n20203), .B(n20202), .Z(n20205) );
  NAND U26638 ( .A(n20205), .B(n20204), .Z(n20207) );
  IV U26639 ( .A(n20206), .Z(n24184) );
  ANDN U26640 ( .B(n20207), .A(n24184), .Z(n20208) );
  NANDN U26641 ( .A(n20209), .B(n20208), .Z(n20212) );
  AND U26642 ( .A(n20210), .B(n24183), .Z(n20211) );
  NAND U26643 ( .A(n20212), .B(n20211), .Z(n20213) );
  NANDN U26644 ( .A(n20214), .B(n20213), .Z(n20215) );
  OR U26645 ( .A(n20215), .B(n28139), .Z(n20216) );
  AND U26646 ( .A(n20217), .B(n20216), .Z(n20218) );
  NANDN U26647 ( .A(n28140), .B(n20218), .Z(n20219) );
  AND U26648 ( .A(n28142), .B(n20219), .Z(n20222) );
  NAND U26649 ( .A(n20221), .B(n20220), .Z(n28143) );
  OR U26650 ( .A(n20222), .B(n28143), .Z(n20223) );
  AND U26651 ( .A(n20224), .B(n20223), .Z(n20225) );
  NANDN U26652 ( .A(n28144), .B(n20225), .Z(n20226) );
  AND U26653 ( .A(n20227), .B(n20226), .Z(n20228) );
  OR U26654 ( .A(n20229), .B(n20228), .Z(n20230) );
  NAND U26655 ( .A(n20231), .B(n20230), .Z(n20232) );
  NANDN U26656 ( .A(n20233), .B(n20232), .Z(n20234) );
  OR U26657 ( .A(n20235), .B(n20234), .Z(n20236) );
  AND U26658 ( .A(n24179), .B(n20236), .Z(n20237) );
  OR U26659 ( .A(n20238), .B(n20237), .Z(n20239) );
  NAND U26660 ( .A(n28150), .B(n20239), .Z(n20240) );
  NAND U26661 ( .A(n28151), .B(n20240), .Z(n20242) );
  OR U26662 ( .A(n20242), .B(n20241), .Z(n20243) );
  NAND U26663 ( .A(n28154), .B(n20243), .Z(n20244) );
  NANDN U26664 ( .A(n20245), .B(n20244), .Z(n20246) );
  OR U26665 ( .A(n28156), .B(n20246), .Z(n20247) );
  AND U26666 ( .A(n28157), .B(n20247), .Z(n20250) );
  NAND U26667 ( .A(n20249), .B(n20248), .Z(n24175) );
  OR U26668 ( .A(n20250), .B(n24175), .Z(n20251) );
  NANDN U26669 ( .A(x[2744]), .B(y[2744]), .Z(n24174) );
  AND U26670 ( .A(n20251), .B(n24174), .Z(n20252) );
  NANDN U26671 ( .A(n20253), .B(n20252), .Z(n20254) );
  AND U26672 ( .A(n28158), .B(n20254), .Z(n20255) );
  OR U26673 ( .A(n20256), .B(n20255), .Z(n20257) );
  NAND U26674 ( .A(n28160), .B(n20257), .Z(n20258) );
  NANDN U26675 ( .A(n20259), .B(n20258), .Z(n20260) );
  ANDN U26676 ( .B(y[2748]), .A(x[2748]), .Z(n28161) );
  OR U26677 ( .A(n20260), .B(n28161), .Z(n20261) );
  AND U26678 ( .A(n20262), .B(n20261), .Z(n20263) );
  OR U26679 ( .A(n20264), .B(n20263), .Z(n20265) );
  NAND U26680 ( .A(n28167), .B(n20265), .Z(n20266) );
  NANDN U26681 ( .A(n28168), .B(n20266), .Z(n20267) );
  AND U26682 ( .A(n28169), .B(n20267), .Z(n20272) );
  NANDN U26683 ( .A(n20272), .B(n28170), .Z(n20273) );
  NAND U26684 ( .A(n28171), .B(n20273), .Z(n20274) );
  NAND U26685 ( .A(n28172), .B(n20274), .Z(n20276) );
  IV U26686 ( .A(n20275), .Z(n28173) );
  AND U26687 ( .A(n20276), .B(n28173), .Z(n20278) );
  IV U26688 ( .A(n20277), .Z(n28174) );
  OR U26689 ( .A(n20278), .B(n28174), .Z(n20279) );
  AND U26690 ( .A(n28175), .B(n20279), .Z(n20280) );
  OR U26691 ( .A(n20281), .B(n20280), .Z(n20282) );
  AND U26692 ( .A(n20283), .B(n20282), .Z(n20284) );
  ANDN U26693 ( .B(n20285), .A(n20284), .Z(n20286) );
  NAND U26694 ( .A(n20287), .B(n20286), .Z(n20288) );
  NANDN U26695 ( .A(n20289), .B(n20288), .Z(n20290) );
  OR U26696 ( .A(n20291), .B(n20290), .Z(n20292) );
  AND U26697 ( .A(n20293), .B(n20292), .Z(n20294) );
  NANDN U26698 ( .A(n20295), .B(n20294), .Z(n20296) );
  AND U26699 ( .A(n20297), .B(n20296), .Z(n20298) );
  OR U26700 ( .A(n20299), .B(n20298), .Z(n20300) );
  NAND U26701 ( .A(n28181), .B(n20300), .Z(n20301) );
  NANDN U26702 ( .A(n20302), .B(n20301), .Z(n20303) );
  ANDN U26703 ( .B(y[2770]), .A(x[2770]), .Z(n28182) );
  OR U26704 ( .A(n20303), .B(n28182), .Z(n20304) );
  AND U26705 ( .A(n20305), .B(n20304), .Z(n20306) );
  NOR U26706 ( .A(n20306), .B(n28189), .Z(n20307) );
  NANDN U26707 ( .A(n20308), .B(n20307), .Z(n20309) );
  AND U26708 ( .A(n20309), .B(n28190), .Z(n20311) );
  NAND U26709 ( .A(n20311), .B(n20310), .Z(n20312) );
  NAND U26710 ( .A(n28191), .B(n20312), .Z(n20313) );
  AND U26711 ( .A(n20314), .B(n20313), .Z(n20315) );
  NANDN U26712 ( .A(n20315), .B(n28192), .Z(n20316) );
  NAND U26713 ( .A(n20317), .B(n20316), .Z(n20318) );
  NANDN U26714 ( .A(n28194), .B(n20318), .Z(n20319) );
  AND U26715 ( .A(n20320), .B(n20319), .Z(n20321) );
  NAND U26716 ( .A(n20322), .B(n20321), .Z(n20325) );
  NANDN U26717 ( .A(n28197), .B(n20323), .Z(n20324) );
  ANDN U26718 ( .B(n20325), .A(n20324), .Z(n20328) );
  NAND U26719 ( .A(n28196), .B(n20326), .Z(n20327) );
  OR U26720 ( .A(n20328), .B(n20327), .Z(n20329) );
  AND U26721 ( .A(n20330), .B(n20329), .Z(n20334) );
  NAND U26722 ( .A(n20332), .B(n20331), .Z(n20333) );
  OR U26723 ( .A(n20334), .B(n20333), .Z(n20335) );
  AND U26724 ( .A(n20336), .B(n20335), .Z(n20337) );
  ANDN U26725 ( .B(n20338), .A(n20337), .Z(n20339) );
  NAND U26726 ( .A(n28203), .B(n20339), .Z(n20340) );
  NANDN U26727 ( .A(n20341), .B(n20340), .Z(n20342) );
  OR U26728 ( .A(n20342), .B(n24167), .Z(n20343) );
  NAND U26729 ( .A(n28204), .B(n20343), .Z(n20344) );
  NANDN U26730 ( .A(n20345), .B(n20344), .Z(n20347) );
  AND U26731 ( .A(n28206), .B(n24165), .Z(n20346) );
  NAND U26732 ( .A(n20347), .B(n20346), .Z(n20348) );
  NANDN U26733 ( .A(n20349), .B(n20348), .Z(n20350) );
  OR U26734 ( .A(n28207), .B(n20350), .Z(n20351) );
  AND U26735 ( .A(n28208), .B(n20351), .Z(n20352) );
  ANDN U26736 ( .B(n20353), .A(n20352), .Z(n20355) );
  NANDN U26737 ( .A(n20355), .B(n28209), .Z(n20356) );
  AND U26738 ( .A(n28210), .B(n20356), .Z(n20357) );
  NANDN U26739 ( .A(n20358), .B(n20357), .Z(n20359) );
  AND U26740 ( .A(n28213), .B(n20359), .Z(n20361) );
  NANDN U26741 ( .A(n20361), .B(n28214), .Z(n20362) );
  AND U26742 ( .A(n20362), .B(n24161), .Z(n20363) );
  NANDN U26743 ( .A(n20364), .B(n20363), .Z(n20365) );
  AND U26744 ( .A(n20365), .B(n28217), .Z(n20366) );
  NAND U26745 ( .A(n28215), .B(n20366), .Z(n20368) );
  IV U26746 ( .A(n20367), .Z(n28219) );
  AND U26747 ( .A(n20368), .B(n28219), .Z(n20369) );
  NANDN U26748 ( .A(n20370), .B(n20369), .Z(n20375) );
  IV U26749 ( .A(n20371), .Z(n28218) );
  AND U26750 ( .A(n28220), .B(n28218), .Z(n20373) );
  OR U26751 ( .A(n20373), .B(n20372), .Z(n20374) );
  AND U26752 ( .A(n20375), .B(n20374), .Z(n20376) );
  OR U26753 ( .A(n20377), .B(n20376), .Z(n20378) );
  NAND U26754 ( .A(n24159), .B(n20378), .Z(n20379) );
  NANDN U26755 ( .A(n20380), .B(n20379), .Z(n20384) );
  IV U26756 ( .A(n20381), .Z(n24160) );
  AND U26757 ( .A(n20382), .B(n24160), .Z(n20383) );
  NAND U26758 ( .A(n20384), .B(n20383), .Z(n20385) );
  NANDN U26759 ( .A(n20386), .B(n20385), .Z(n20387) );
  OR U26760 ( .A(n20388), .B(n20387), .Z(n20389) );
  AND U26761 ( .A(n20390), .B(n20389), .Z(n20391) );
  NANDN U26762 ( .A(n20392), .B(n20391), .Z(n20393) );
  AND U26763 ( .A(n20394), .B(n20393), .Z(n20395) );
  OR U26764 ( .A(n20396), .B(n20395), .Z(n20397) );
  NAND U26765 ( .A(n24155), .B(n20397), .Z(n20398) );
  NANDN U26766 ( .A(n28231), .B(n20398), .Z(n20400) );
  IV U26767 ( .A(n20399), .Z(n24154) );
  OR U26768 ( .A(n20400), .B(n24154), .Z(n20401) );
  AND U26769 ( .A(n24156), .B(n20401), .Z(n20404) );
  NANDN U26770 ( .A(n20404), .B(n28232), .Z(n20405) );
  NAND U26771 ( .A(n28233), .B(n20405), .Z(n20406) );
  NANDN U26772 ( .A(n20407), .B(n20406), .Z(n20409) );
  AND U26773 ( .A(n28237), .B(n28235), .Z(n20408) );
  NAND U26774 ( .A(n20409), .B(n20408), .Z(n20410) );
  NANDN U26775 ( .A(n20411), .B(n20410), .Z(n20412) );
  OR U26776 ( .A(n28238), .B(n20412), .Z(n20413) );
  AND U26777 ( .A(n28239), .B(n20413), .Z(n20416) );
  NAND U26778 ( .A(n20415), .B(n20414), .Z(n24153) );
  OR U26779 ( .A(n20416), .B(n24153), .Z(n20417) );
  NAND U26780 ( .A(n20418), .B(n20417), .Z(n20419) );
  NANDN U26781 ( .A(n20420), .B(n20419), .Z(n20421) );
  OR U26782 ( .A(n20421), .B(n28241), .Z(n20422) );
  AND U26783 ( .A(n20423), .B(n20422), .Z(n20426) );
  NAND U26784 ( .A(n28246), .B(n20424), .Z(n20425) );
  OR U26785 ( .A(n20426), .B(n20425), .Z(n20427) );
  AND U26786 ( .A(n20428), .B(n20427), .Z(n20429) );
  NANDN U26787 ( .A(n20429), .B(n28248), .Z(n20430) );
  AND U26788 ( .A(n20431), .B(n20430), .Z(n20432) );
  NANDN U26789 ( .A(n20432), .B(n28250), .Z(n20433) );
  AND U26790 ( .A(n20434), .B(n20433), .Z(n20437) );
  NANDN U26791 ( .A(n20437), .B(n28252), .Z(n20438) );
  NANDN U26792 ( .A(n24152), .B(n20438), .Z(n20439) );
  AND U26793 ( .A(n28253), .B(n20439), .Z(n20442) );
  NAND U26794 ( .A(n20441), .B(n20440), .Z(n28254) );
  OR U26795 ( .A(n20442), .B(n28254), .Z(n20443) );
  AND U26796 ( .A(n20444), .B(n20443), .Z(n20445) );
  NANDN U26797 ( .A(n28255), .B(n20445), .Z(n20446) );
  AND U26798 ( .A(n28257), .B(n20446), .Z(n20447) );
  OR U26799 ( .A(n20448), .B(n20447), .Z(n20449) );
  NAND U26800 ( .A(n28265), .B(n20449), .Z(n20450) );
  NANDN U26801 ( .A(n20451), .B(n20450), .Z(n20452) );
  ANDN U26802 ( .B(y[2836]), .A(x[2836]), .Z(n28267) );
  OR U26803 ( .A(n20452), .B(n28267), .Z(n20453) );
  AND U26804 ( .A(n20454), .B(n20453), .Z(n20455) );
  OR U26805 ( .A(n20456), .B(n20455), .Z(n20457) );
  NAND U26806 ( .A(n28277), .B(n20457), .Z(n20458) );
  NANDN U26807 ( .A(n28279), .B(n20458), .Z(n20462) );
  IV U26808 ( .A(n20459), .Z(n28280) );
  AND U26809 ( .A(n20460), .B(n28280), .Z(n20461) );
  NAND U26810 ( .A(n20462), .B(n20461), .Z(n20463) );
  NANDN U26811 ( .A(n20464), .B(n20463), .Z(n20466) );
  IV U26812 ( .A(n20465), .Z(n28282) );
  OR U26813 ( .A(n20466), .B(n28282), .Z(n20467) );
  NAND U26814 ( .A(n20468), .B(n20467), .Z(n20469) );
  NANDN U26815 ( .A(n20470), .B(n20469), .Z(n20471) );
  OR U26816 ( .A(n20471), .B(n28290), .Z(n20472) );
  AND U26817 ( .A(n20473), .B(n20472), .Z(n20477) );
  NANDN U26818 ( .A(n20477), .B(n28295), .Z(n20478) );
  AND U26819 ( .A(n20479), .B(n20478), .Z(n20480) );
  OR U26820 ( .A(n20481), .B(n20480), .Z(n20482) );
  NAND U26821 ( .A(n20483), .B(n20482), .Z(n20484) );
  NANDN U26822 ( .A(n20485), .B(n20484), .Z(n20489) );
  AND U26823 ( .A(n20487), .B(n20486), .Z(n20488) );
  NAND U26824 ( .A(n20489), .B(n20488), .Z(n20490) );
  NANDN U26825 ( .A(n20491), .B(n20490), .Z(n20492) );
  OR U26826 ( .A(n20493), .B(n20492), .Z(n20494) );
  AND U26827 ( .A(n20495), .B(n20494), .Z(n20496) );
  NANDN U26828 ( .A(n28304), .B(n20496), .Z(n20497) );
  AND U26829 ( .A(n20498), .B(n20497), .Z(n20499) );
  OR U26830 ( .A(n28306), .B(n20499), .Z(n20500) );
  NAND U26831 ( .A(n28307), .B(n20500), .Z(n20501) );
  NANDN U26832 ( .A(n28308), .B(n20501), .Z(n20502) );
  NAND U26833 ( .A(n28309), .B(n20502), .Z(n20503) );
  AND U26834 ( .A(n28310), .B(n20503), .Z(n20506) );
  NANDN U26835 ( .A(n20506), .B(n28311), .Z(n20507) );
  NAND U26836 ( .A(n20508), .B(n20507), .Z(n20509) );
  NANDN U26837 ( .A(n20510), .B(n20509), .Z(n20511) );
  OR U26838 ( .A(n20511), .B(n28312), .Z(n20512) );
  AND U26839 ( .A(n20513), .B(n20512), .Z(n20516) );
  NAND U26840 ( .A(n28317), .B(n20514), .Z(n20515) );
  OR U26841 ( .A(n20516), .B(n20515), .Z(n20517) );
  AND U26842 ( .A(n20518), .B(n20517), .Z(n20519) );
  OR U26843 ( .A(n28319), .B(n20519), .Z(n20520) );
  NAND U26844 ( .A(n20521), .B(n20520), .Z(n20522) );
  NANDN U26845 ( .A(n20523), .B(n20522), .Z(n20525) );
  IV U26846 ( .A(n20524), .Z(n28321) );
  OR U26847 ( .A(n20525), .B(n28321), .Z(n20526) );
  AND U26848 ( .A(n20527), .B(n20526), .Z(n20531) );
  NAND U26849 ( .A(n20529), .B(n20528), .Z(n20530) );
  OR U26850 ( .A(n20531), .B(n20530), .Z(n20532) );
  AND U26851 ( .A(n20533), .B(n20532), .Z(n20534) );
  OR U26852 ( .A(n20535), .B(n20534), .Z(n20536) );
  NAND U26853 ( .A(n20537), .B(n20536), .Z(n20541) );
  AND U26854 ( .A(n20539), .B(n20538), .Z(n20540) );
  NAND U26855 ( .A(n20541), .B(n20540), .Z(n20542) );
  NANDN U26856 ( .A(n28329), .B(n20542), .Z(n20543) );
  OR U26857 ( .A(n20544), .B(n20543), .Z(n20545) );
  AND U26858 ( .A(n20546), .B(n20545), .Z(n20547) );
  NANDN U26859 ( .A(n24148), .B(n20547), .Z(n20548) );
  AND U26860 ( .A(n28331), .B(n20548), .Z(n20549) );
  OR U26861 ( .A(n28332), .B(n20549), .Z(n20550) );
  NAND U26862 ( .A(n28333), .B(n20550), .Z(n20551) );
  NANDN U26863 ( .A(n28334), .B(n20551), .Z(n20552) );
  AND U26864 ( .A(n28335), .B(n20552), .Z(n20554) );
  IV U26865 ( .A(n20553), .Z(n28336) );
  OR U26866 ( .A(n20554), .B(n28336), .Z(n20555) );
  NAND U26867 ( .A(n28337), .B(n20555), .Z(n20556) );
  NANDN U26868 ( .A(n28338), .B(n20556), .Z(n20560) );
  IV U26869 ( .A(n20557), .Z(n28339) );
  AND U26870 ( .A(n20558), .B(n28339), .Z(n20559) );
  NAND U26871 ( .A(n20560), .B(n20559), .Z(n20561) );
  NANDN U26872 ( .A(n28340), .B(n20561), .Z(n20562) );
  OR U26873 ( .A(n20563), .B(n20562), .Z(n20564) );
  AND U26874 ( .A(n28342), .B(n20564), .Z(n20566) );
  NAND U26875 ( .A(n20566), .B(n20565), .Z(n20567) );
  NANDN U26876 ( .A(n20568), .B(n20567), .Z(n20569) );
  AND U26877 ( .A(n20569), .B(n28344), .Z(n20570) );
  OR U26878 ( .A(n28345), .B(n20570), .Z(n20571) );
  NAND U26879 ( .A(n20572), .B(n20571), .Z(n20573) );
  NANDN U26880 ( .A(n20574), .B(n20573), .Z(n20576) );
  IV U26881 ( .A(n20575), .Z(n28347) );
  OR U26882 ( .A(n20576), .B(n28347), .Z(n20577) );
  NAND U26883 ( .A(n20578), .B(n20577), .Z(n20582) );
  AND U26884 ( .A(n20580), .B(n20579), .Z(n20581) );
  NAND U26885 ( .A(n20582), .B(n20581), .Z(n20583) );
  NANDN U26886 ( .A(n28351), .B(n20583), .Z(n20585) );
  OR U26887 ( .A(n20585), .B(n20584), .Z(n20586) );
  NAND U26888 ( .A(n20587), .B(n20586), .Z(n20588) );
  NANDN U26889 ( .A(n28353), .B(n20588), .Z(n20590) );
  AND U26890 ( .A(n20590), .B(n20589), .Z(n20591) );
  NANDN U26891 ( .A(x[2898]), .B(y[2898]), .Z(n28354) );
  AND U26892 ( .A(n20591), .B(n28354), .Z(n20592) );
  OR U26893 ( .A(n20593), .B(n20592), .Z(n20594) );
  NAND U26894 ( .A(n20595), .B(n20594), .Z(n20596) );
  NANDN U26895 ( .A(n28357), .B(n20596), .Z(n20597) );
  AND U26896 ( .A(n20598), .B(n20597), .Z(n20599) );
  NAND U26897 ( .A(n28358), .B(n20599), .Z(n20600) );
  NANDN U26898 ( .A(n28359), .B(n20600), .Z(n20602) );
  IV U26899 ( .A(n20601), .Z(n28363) );
  OR U26900 ( .A(n20602), .B(n28363), .Z(n20603) );
  AND U26901 ( .A(n20604), .B(n20603), .Z(n20605) );
  NANDN U26902 ( .A(n28364), .B(n20605), .Z(n20606) );
  AND U26903 ( .A(n28365), .B(n20606), .Z(n20608) );
  NANDN U26904 ( .A(n20608), .B(n28366), .Z(n20609) );
  AND U26905 ( .A(n20610), .B(n20609), .Z(n20611) );
  NAND U26906 ( .A(n20611), .B(n28367), .Z(n20612) );
  ANDN U26907 ( .B(n20612), .A(n28370), .Z(n20613) );
  NANDN U26908 ( .A(n28368), .B(n20613), .Z(n20614) );
  NAND U26909 ( .A(n20615), .B(n20614), .Z(n20616) );
  NAND U26910 ( .A(n28371), .B(n20616), .Z(n20617) );
  AND U26911 ( .A(n20618), .B(n20617), .Z(n20619) );
  NAND U26912 ( .A(n24142), .B(n20619), .Z(n20620) );
  NANDN U26913 ( .A(n24141), .B(n20620), .Z(n20621) );
  AND U26914 ( .A(n20621), .B(n24140), .Z(n20622) );
  OR U26915 ( .A(n20622), .B(n28376), .Z(n20623) );
  NAND U26916 ( .A(n28378), .B(n20623), .Z(n20624) );
  NAND U26917 ( .A(n28379), .B(n20624), .Z(n20625) );
  NAND U26918 ( .A(n28380), .B(n20625), .Z(n20626) );
  ANDN U26919 ( .B(n20626), .A(n24139), .Z(n20627) );
  NANDN U26920 ( .A(n20628), .B(n20627), .Z(n20630) );
  IV U26921 ( .A(n20629), .Z(n28383) );
  AND U26922 ( .A(n20630), .B(n28383), .Z(n20631) );
  NAND U26923 ( .A(n28381), .B(n20631), .Z(n20632) );
  AND U26924 ( .A(n20633), .B(n20632), .Z(n20634) );
  NANDN U26925 ( .A(n28384), .B(n20634), .Z(n20635) );
  AND U26926 ( .A(n28385), .B(n20635), .Z(n20636) );
  NOR U26927 ( .A(n28386), .B(n20636), .Z(n20637) );
  NAND U26928 ( .A(n20638), .B(n20637), .Z(n20639) );
  NANDN U26929 ( .A(n24138), .B(n20639), .Z(n20640) );
  OR U26930 ( .A(n20640), .B(n28387), .Z(n20641) );
  AND U26931 ( .A(n20642), .B(n20641), .Z(n20643) );
  NANDN U26932 ( .A(n28388), .B(n20643), .Z(n20644) );
  AND U26933 ( .A(n28390), .B(n20644), .Z(n20647) );
  NANDN U26934 ( .A(x[2928]), .B(y[2928]), .Z(n20646) );
  NAND U26935 ( .A(n20646), .B(n20645), .Z(n28391) );
  OR U26936 ( .A(n20647), .B(n28391), .Z(n20648) );
  AND U26937 ( .A(n20649), .B(n20648), .Z(n20650) );
  NANDN U26938 ( .A(n28392), .B(n20650), .Z(n20651) );
  AND U26939 ( .A(n20652), .B(n20651), .Z(n20653) );
  OR U26940 ( .A(n20654), .B(n20653), .Z(n20655) );
  NAND U26941 ( .A(n20656), .B(n20655), .Z(n20657) );
  NANDN U26942 ( .A(n20658), .B(n20657), .Z(n20659) );
  OR U26943 ( .A(n20660), .B(n20659), .Z(n20661) );
  AND U26944 ( .A(n24135), .B(n20661), .Z(n20662) );
  ANDN U26945 ( .B(n20663), .A(n20662), .Z(n20664) );
  NAND U26946 ( .A(n24134), .B(n20664), .Z(n20665) );
  NANDN U26947 ( .A(n20666), .B(n20665), .Z(n20667) );
  OR U26948 ( .A(n20667), .B(n24136), .Z(n20668) );
  NAND U26949 ( .A(n20669), .B(n20668), .Z(n20670) );
  NANDN U26950 ( .A(n20671), .B(n20670), .Z(n20673) );
  OR U26951 ( .A(n20673), .B(n20672), .Z(n20674) );
  AND U26952 ( .A(n20675), .B(n20674), .Z(n20676) );
  OR U26953 ( .A(n20677), .B(n20676), .Z(n20678) );
  NAND U26954 ( .A(n20679), .B(n20678), .Z(n20682) );
  AND U26955 ( .A(n28406), .B(n20680), .Z(n20681) );
  NAND U26956 ( .A(n20682), .B(n20681), .Z(n20683) );
  NANDN U26957 ( .A(n20684), .B(n20683), .Z(n20685) );
  NANDN U26958 ( .A(n20686), .B(n20685), .Z(n20687) );
  AND U26959 ( .A(n24130), .B(n20687), .Z(n20688) );
  ANDN U26960 ( .B(n20689), .A(n20688), .Z(n20690) );
  NAND U26961 ( .A(n20691), .B(n20690), .Z(n20692) );
  NANDN U26962 ( .A(n24131), .B(n20692), .Z(n20694) );
  OR U26963 ( .A(n20694), .B(n20693), .Z(n20695) );
  NAND U26964 ( .A(n20696), .B(n20695), .Z(n20697) );
  NANDN U26965 ( .A(n20698), .B(n20697), .Z(n20700) );
  OR U26966 ( .A(n20700), .B(n20699), .Z(n20701) );
  NANDN U26967 ( .A(n28415), .B(n20701), .Z(n20702) );
  NANDN U26968 ( .A(n28414), .B(n20702), .Z(n20703) );
  OR U26969 ( .A(n20704), .B(n20703), .Z(n20705) );
  AND U26970 ( .A(n20705), .B(n24127), .Z(n20706) );
  NAND U26971 ( .A(n20706), .B(x[2953]), .Z(n20709) );
  XOR U26972 ( .A(n20706), .B(x[2953]), .Z(n20707) );
  NANDN U26973 ( .A(y[2953]), .B(n20707), .Z(n20708) );
  NAND U26974 ( .A(n20709), .B(n20708), .Z(n20711) );
  OR U26975 ( .A(n20711), .B(n20710), .Z(n20712) );
  AND U26976 ( .A(n20713), .B(n20712), .Z(n20714) );
  OR U26977 ( .A(n20715), .B(n20714), .Z(n20716) );
  NAND U26978 ( .A(n28421), .B(n20716), .Z(n20717) );
  NANDN U26979 ( .A(n20718), .B(n20717), .Z(n20719) );
  NANDN U26980 ( .A(n20719), .B(n28422), .Z(n20720) );
  AND U26981 ( .A(n20721), .B(n20720), .Z(n20723) );
  NOR U26982 ( .A(n20723), .B(n20722), .Z(n20724) );
  NANDN U26983 ( .A(n20725), .B(n20724), .Z(n20726) );
  AND U26984 ( .A(n20727), .B(n20726), .Z(n20728) );
  NAND U26985 ( .A(n28423), .B(n20728), .Z(n20729) );
  NANDN U26986 ( .A(n20730), .B(n20729), .Z(n20731) );
  AND U26987 ( .A(n20731), .B(n28426), .Z(n20734) );
  OR U26988 ( .A(n20734), .B(n28427), .Z(n20735) );
  AND U26989 ( .A(n28428), .B(n20735), .Z(n20737) );
  NAND U26990 ( .A(n20737), .B(n20736), .Z(n20738) );
  NANDN U26991 ( .A(n28429), .B(n20738), .Z(n20739) );
  AND U26992 ( .A(n20740), .B(n20739), .Z(n20741) );
  OR U26993 ( .A(n28433), .B(n20741), .Z(n20742) );
  NAND U26994 ( .A(n20743), .B(n20742), .Z(n20744) );
  NANDN U26995 ( .A(n20745), .B(n20744), .Z(n20746) );
  OR U26996 ( .A(n20746), .B(n28435), .Z(n20747) );
  NAND U26997 ( .A(n20748), .B(n20747), .Z(n20749) );
  NAND U26998 ( .A(n20750), .B(n20749), .Z(n20751) );
  NAND U26999 ( .A(n28440), .B(n20751), .Z(n20753) );
  IV U27000 ( .A(n20752), .Z(n28441) );
  AND U27001 ( .A(n20753), .B(n28441), .Z(n20755) );
  IV U27002 ( .A(n20754), .Z(n28444) );
  OR U27003 ( .A(n20755), .B(n28444), .Z(n20756) );
  AND U27004 ( .A(n24122), .B(n20756), .Z(n20757) );
  ANDN U27005 ( .B(n20758), .A(n20757), .Z(n20760) );
  OR U27006 ( .A(n20760), .B(n20759), .Z(n20761) );
  NAND U27007 ( .A(n28447), .B(n20761), .Z(n20762) );
  NANDN U27008 ( .A(n20763), .B(n20762), .Z(n20767) );
  IV U27009 ( .A(n20764), .Z(n28446) );
  AND U27010 ( .A(n20765), .B(n28446), .Z(n20766) );
  NAND U27011 ( .A(n20767), .B(n20766), .Z(n20768) );
  NANDN U27012 ( .A(n20769), .B(n20768), .Z(n20771) );
  OR U27013 ( .A(n20771), .B(n20770), .Z(n20772) );
  AND U27014 ( .A(n20773), .B(n20772), .Z(n20777) );
  NAND U27015 ( .A(n20775), .B(n20774), .Z(n20776) );
  OR U27016 ( .A(n20777), .B(n20776), .Z(n20778) );
  AND U27017 ( .A(n20779), .B(n20778), .Z(n20783) );
  NAND U27018 ( .A(n20781), .B(n20780), .Z(n20782) );
  OR U27019 ( .A(n20783), .B(n20782), .Z(n20784) );
  AND U27020 ( .A(n20785), .B(n20784), .Z(n20786) );
  NOR U27021 ( .A(n20787), .B(n20786), .Z(n20788) );
  NANDN U27022 ( .A(n20789), .B(n20788), .Z(n20790) );
  AND U27023 ( .A(n20791), .B(n20790), .Z(n20793) );
  NAND U27024 ( .A(n20793), .B(n20792), .Z(n20794) );
  NAND U27025 ( .A(n24116), .B(n20794), .Z(n20795) );
  AND U27026 ( .A(n20796), .B(n20795), .Z(n20797) );
  ANDN U27027 ( .B(n20798), .A(n20797), .Z(n20799) );
  NAND U27028 ( .A(n24118), .B(n20799), .Z(n20800) );
  NANDN U27029 ( .A(n20801), .B(n20800), .Z(n20803) );
  IV U27030 ( .A(n20802), .Z(n28459) );
  OR U27031 ( .A(n20803), .B(n28459), .Z(n20805) );
  IV U27032 ( .A(n20804), .Z(n28460) );
  AND U27033 ( .A(n20805), .B(n28460), .Z(n20807) );
  NAND U27034 ( .A(n20807), .B(n20806), .Z(n20808) );
  NANDN U27035 ( .A(n28461), .B(n20808), .Z(n20809) );
  AND U27036 ( .A(n28463), .B(n20809), .Z(n20812) );
  AND U27037 ( .A(n20812), .B(n28462), .Z(n20813) );
  OR U27038 ( .A(n28464), .B(n20813), .Z(n20814) );
  NAND U27039 ( .A(n20815), .B(n20814), .Z(n20816) );
  NANDN U27040 ( .A(n20817), .B(n20816), .Z(n20818) );
  NAND U27041 ( .A(n20819), .B(n20818), .Z(n20820) );
  NAND U27042 ( .A(n28470), .B(n20820), .Z(n20823) );
  AND U27043 ( .A(n20822), .B(n20821), .Z(n28471) );
  AND U27044 ( .A(n20823), .B(n28471), .Z(n20826) );
  NANDN U27045 ( .A(n20826), .B(n28472), .Z(n20827) );
  NAND U27046 ( .A(n24113), .B(n20827), .Z(n20828) );
  NANDN U27047 ( .A(n28474), .B(n20828), .Z(n20829) );
  NAND U27048 ( .A(n28475), .B(n20829), .Z(n20832) );
  AND U27049 ( .A(n20831), .B(n20830), .Z(n28476) );
  AND U27050 ( .A(n20832), .B(n28476), .Z(n20835) );
  NANDN U27051 ( .A(n20835), .B(n28477), .Z(n20836) );
  AND U27052 ( .A(n20837), .B(n20836), .Z(n20838) );
  NAND U27053 ( .A(n24112), .B(n20838), .Z(n20839) );
  NANDN U27054 ( .A(n20840), .B(n20839), .Z(n20841) );
  AND U27055 ( .A(n20842), .B(n20841), .Z(n20845) );
  AND U27056 ( .A(n20844), .B(n20843), .Z(n28481) );
  NANDN U27057 ( .A(n20845), .B(n28481), .Z(n20846) );
  NAND U27058 ( .A(n28482), .B(n20846), .Z(n20847) );
  NANDN U27059 ( .A(n20848), .B(n20847), .Z(n20852) );
  IV U27060 ( .A(n20849), .Z(n28484) );
  AND U27061 ( .A(n20850), .B(n28484), .Z(n20851) );
  NAND U27062 ( .A(n20852), .B(n20851), .Z(n20853) );
  NANDN U27063 ( .A(n20854), .B(n20853), .Z(n20856) );
  OR U27064 ( .A(n20856), .B(n20855), .Z(n20857) );
  NAND U27065 ( .A(n20858), .B(n20857), .Z(n20859) );
  NANDN U27066 ( .A(n20860), .B(n20859), .Z(n20862) );
  OR U27067 ( .A(n20862), .B(n20861), .Z(n20863) );
  NAND U27068 ( .A(n28492), .B(n20863), .Z(n20864) );
  NANDN U27069 ( .A(n28491), .B(n20864), .Z(n20865) );
  OR U27070 ( .A(n20866), .B(n20865), .Z(n20867) );
  AND U27071 ( .A(n20868), .B(n20867), .Z(n20869) );
  NAND U27072 ( .A(n20869), .B(n28490), .Z(n20871) );
  ANDN U27073 ( .B(n20871), .A(n20870), .Z(n20872) );
  NANDN U27074 ( .A(n20873), .B(n20872), .Z(n20874) );
  NAND U27075 ( .A(n20875), .B(n20874), .Z(n20876) );
  NANDN U27076 ( .A(n20877), .B(n20876), .Z(n20878) );
  AND U27077 ( .A(n20879), .B(n20878), .Z(n20880) );
  OR U27078 ( .A(n20881), .B(n20880), .Z(n20882) );
  NAND U27079 ( .A(n20883), .B(n20882), .Z(n20884) );
  NANDN U27080 ( .A(n20885), .B(n20884), .Z(n20886) );
  AND U27081 ( .A(n20887), .B(n20886), .Z(n20890) );
  AND U27082 ( .A(n20889), .B(n20888), .Z(n24107) );
  NANDN U27083 ( .A(n20890), .B(n24107), .Z(n20891) );
  AND U27084 ( .A(n20892), .B(n20891), .Z(n20893) );
  NAND U27085 ( .A(n24106), .B(n20893), .Z(n20895) );
  ANDN U27086 ( .B(n20895), .A(n20894), .Z(n20896) );
  NANDN U27087 ( .A(n24108), .B(n20896), .Z(n20897) );
  NAND U27088 ( .A(n20898), .B(n20897), .Z(n20899) );
  NANDN U27089 ( .A(n20900), .B(n20899), .Z(n20901) );
  AND U27090 ( .A(n20902), .B(n20901), .Z(n20903) );
  NAND U27091 ( .A(n20904), .B(n20903), .Z(n20905) );
  NAND U27092 ( .A(n28507), .B(n20905), .Z(n20906) );
  AND U27093 ( .A(n28508), .B(n20906), .Z(n20907) );
  OR U27094 ( .A(n28509), .B(n20907), .Z(n20908) );
  NAND U27095 ( .A(n28510), .B(n20908), .Z(n20909) );
  NANDN U27096 ( .A(n20910), .B(n20909), .Z(n20911) );
  NAND U27097 ( .A(n28515), .B(n20911), .Z(n20912) );
  ANDN U27098 ( .B(n20912), .A(n28514), .Z(n20913) );
  NANDN U27099 ( .A(n20914), .B(n20913), .Z(n20915) );
  AND U27100 ( .A(n20916), .B(n20915), .Z(n20917) );
  NAND U27101 ( .A(n28513), .B(n20917), .Z(n20921) );
  NAND U27102 ( .A(n20919), .B(n20918), .Z(n20920) );
  ANDN U27103 ( .B(n20921), .A(n20920), .Z(n20925) );
  NAND U27104 ( .A(n20923), .B(n20922), .Z(n20924) );
  OR U27105 ( .A(n20925), .B(n20924), .Z(n20926) );
  AND U27106 ( .A(n20927), .B(n20926), .Z(n20928) );
  OR U27107 ( .A(n20929), .B(n20928), .Z(n20930) );
  NAND U27108 ( .A(n20931), .B(n20930), .Z(n20935) );
  AND U27109 ( .A(n20933), .B(n20932), .Z(n20934) );
  NAND U27110 ( .A(n20935), .B(n20934), .Z(n20936) );
  NANDN U27111 ( .A(n20937), .B(n20936), .Z(n20939) );
  OR U27112 ( .A(n20939), .B(n20938), .Z(n20940) );
  NAND U27113 ( .A(n20941), .B(n20940), .Z(n20942) );
  NAND U27114 ( .A(n28526), .B(n20942), .Z(n20945) );
  AND U27115 ( .A(n20943), .B(n28525), .Z(n20944) );
  NAND U27116 ( .A(n20945), .B(n20944), .Z(n20946) );
  NANDN U27117 ( .A(n28524), .B(n20946), .Z(n20948) );
  OR U27118 ( .A(n20948), .B(n20947), .Z(n20949) );
  NAND U27119 ( .A(n20950), .B(n20949), .Z(n20951) );
  NANDN U27120 ( .A(n20952), .B(n20951), .Z(n20953) );
  OR U27121 ( .A(n20954), .B(n20953), .Z(n20955) );
  AND U27122 ( .A(n20956), .B(n20955), .Z(n20957) );
  OR U27123 ( .A(n20958), .B(n20957), .Z(n20959) );
  NAND U27124 ( .A(n24098), .B(n20959), .Z(n20960) );
  NANDN U27125 ( .A(n28531), .B(n20960), .Z(n20961) );
  AND U27126 ( .A(n28532), .B(n20961), .Z(n20962) );
  OR U27127 ( .A(n20963), .B(n20962), .Z(n20964) );
  NAND U27128 ( .A(n24097), .B(n20964), .Z(n20965) );
  NANDN U27129 ( .A(n20966), .B(n20965), .Z(n20967) );
  NANDN U27130 ( .A(n20967), .B(n24096), .Z(n20968) );
  NAND U27131 ( .A(n28534), .B(n20968), .Z(n20969) );
  NANDN U27132 ( .A(n20970), .B(n20969), .Z(n20972) );
  OR U27133 ( .A(n20972), .B(n20971), .Z(n20973) );
  AND U27134 ( .A(n20974), .B(n20973), .Z(n20978) );
  NAND U27135 ( .A(n20976), .B(n20975), .Z(n20977) );
  OR U27136 ( .A(n20978), .B(n20977), .Z(n20979) );
  AND U27137 ( .A(n20980), .B(n20979), .Z(n20981) );
  OR U27138 ( .A(n20982), .B(n20981), .Z(n20983) );
  NAND U27139 ( .A(n20984), .B(n20983), .Z(n20987) );
  AND U27140 ( .A(n20985), .B(n24095), .Z(n20986) );
  NAND U27141 ( .A(n20987), .B(n20986), .Z(n20988) );
  NANDN U27142 ( .A(n20989), .B(n20988), .Z(n20990) );
  OR U27143 ( .A(n20990), .B(n28544), .Z(n20991) );
  NAND U27144 ( .A(n28545), .B(n20991), .Z(n20992) );
  NANDN U27145 ( .A(n20993), .B(n20992), .Z(n20996) );
  AND U27146 ( .A(n20994), .B(n28547), .Z(n20995) );
  NAND U27147 ( .A(n20996), .B(n20995), .Z(n20997) );
  NANDN U27148 ( .A(n20998), .B(n20997), .Z(n20999) );
  OR U27149 ( .A(n28550), .B(n20999), .Z(n21000) );
  AND U27150 ( .A(n28551), .B(n21000), .Z(n21002) );
  NAND U27151 ( .A(n21002), .B(n21001), .Z(n21006) );
  NAND U27152 ( .A(n21006), .B(n28552), .Z(n21007) );
  AND U27153 ( .A(n28553), .B(n21007), .Z(n21008) );
  OR U27154 ( .A(n21008), .B(n28554), .Z(n21009) );
  AND U27155 ( .A(n21010), .B(n21009), .Z(n21011) );
  NAND U27156 ( .A(n21012), .B(n21011), .Z(n21013) );
  NAND U27157 ( .A(n28556), .B(n21013), .Z(n21014) );
  NANDN U27158 ( .A(n21015), .B(n21014), .Z(n21016) );
  NAND U27159 ( .A(n21017), .B(n21016), .Z(n21018) );
  NANDN U27160 ( .A(n21019), .B(n21018), .Z(n21021) );
  OR U27161 ( .A(n21021), .B(n21020), .Z(n21022) );
  NAND U27162 ( .A(n21023), .B(n21022), .Z(n21024) );
  NANDN U27163 ( .A(n21025), .B(n21024), .Z(n21027) );
  NAND U27164 ( .A(n21027), .B(n21026), .Z(n21029) );
  ANDN U27165 ( .B(n21029), .A(n21028), .Z(n21030) );
  NANDN U27166 ( .A(n21031), .B(n21030), .Z(n21035) );
  AND U27167 ( .A(n21033), .B(n21032), .Z(n21034) );
  NAND U27168 ( .A(n21035), .B(n21034), .Z(n21036) );
  NANDN U27169 ( .A(n21037), .B(n21036), .Z(n21039) );
  OR U27170 ( .A(n21039), .B(n21038), .Z(n21040) );
  NAND U27171 ( .A(n21041), .B(n21040), .Z(n21042) );
  NANDN U27172 ( .A(n21043), .B(n21042), .Z(n21044) );
  OR U27173 ( .A(n21045), .B(n21044), .Z(n21046) );
  AND U27174 ( .A(n21047), .B(n21046), .Z(n21049) );
  NAND U27175 ( .A(n21049), .B(n21048), .Z(n21051) );
  ANDN U27176 ( .B(n21051), .A(n21050), .Z(n21052) );
  NANDN U27177 ( .A(n21053), .B(n21052), .Z(n21057) );
  AND U27178 ( .A(n21055), .B(n21054), .Z(n21056) );
  NAND U27179 ( .A(n21057), .B(n21056), .Z(n21058) );
  NANDN U27180 ( .A(n21059), .B(n21058), .Z(n21061) );
  OR U27181 ( .A(n21061), .B(n21060), .Z(n21062) );
  NAND U27182 ( .A(n21063), .B(n21062), .Z(n21064) );
  NANDN U27183 ( .A(n21065), .B(n21064), .Z(n21066) );
  OR U27184 ( .A(n21067), .B(n21066), .Z(n21068) );
  AND U27185 ( .A(n21069), .B(n21068), .Z(n21071) );
  NAND U27186 ( .A(n21071), .B(n21070), .Z(n21073) );
  ANDN U27187 ( .B(n21073), .A(n21072), .Z(n21074) );
  NANDN U27188 ( .A(n21075), .B(n21074), .Z(n21079) );
  AND U27189 ( .A(n21077), .B(n21076), .Z(n21078) );
  NAND U27190 ( .A(n21079), .B(n21078), .Z(n21080) );
  NANDN U27191 ( .A(n21081), .B(n21080), .Z(n21083) );
  OR U27192 ( .A(n21083), .B(n21082), .Z(n21084) );
  NAND U27193 ( .A(n21085), .B(n21084), .Z(n21086) );
  NANDN U27194 ( .A(n21087), .B(n21086), .Z(n21088) );
  OR U27195 ( .A(n21089), .B(n21088), .Z(n21090) );
  AND U27196 ( .A(n21091), .B(n21090), .Z(n21093) );
  NAND U27197 ( .A(n21093), .B(n21092), .Z(n21095) );
  ANDN U27198 ( .B(n21095), .A(n21094), .Z(n21096) );
  NANDN U27199 ( .A(n21097), .B(n21096), .Z(n21101) );
  AND U27200 ( .A(n21099), .B(n21098), .Z(n21100) );
  NAND U27201 ( .A(n21101), .B(n21100), .Z(n21102) );
  NANDN U27202 ( .A(n21103), .B(n21102), .Z(n21105) );
  OR U27203 ( .A(n21105), .B(n21104), .Z(n21106) );
  NAND U27204 ( .A(n21107), .B(n21106), .Z(n21108) );
  NANDN U27205 ( .A(n21109), .B(n21108), .Z(n21110) );
  OR U27206 ( .A(n21111), .B(n21110), .Z(n21112) );
  AND U27207 ( .A(n21113), .B(n21112), .Z(n21115) );
  NAND U27208 ( .A(n21115), .B(n21114), .Z(n21117) );
  ANDN U27209 ( .B(n21117), .A(n21116), .Z(n21118) );
  NANDN U27210 ( .A(n21119), .B(n21118), .Z(n21123) );
  AND U27211 ( .A(n21121), .B(n21120), .Z(n21122) );
  NAND U27212 ( .A(n21123), .B(n21122), .Z(n21124) );
  NANDN U27213 ( .A(n21125), .B(n21124), .Z(n21127) );
  OR U27214 ( .A(n21127), .B(n21126), .Z(n21128) );
  NAND U27215 ( .A(n21129), .B(n21128), .Z(n21130) );
  NANDN U27216 ( .A(n21131), .B(n21130), .Z(n21132) );
  OR U27217 ( .A(n21133), .B(n21132), .Z(n21134) );
  AND U27218 ( .A(n21135), .B(n21134), .Z(n21137) );
  NAND U27219 ( .A(n21137), .B(n21136), .Z(n21139) );
  ANDN U27220 ( .B(n21139), .A(n21138), .Z(n21140) );
  NANDN U27221 ( .A(n21141), .B(n21140), .Z(n21145) );
  AND U27222 ( .A(n21143), .B(n21142), .Z(n21144) );
  NAND U27223 ( .A(n21145), .B(n21144), .Z(n21146) );
  NANDN U27224 ( .A(n21147), .B(n21146), .Z(n21149) );
  OR U27225 ( .A(n21149), .B(n21148), .Z(n21150) );
  NAND U27226 ( .A(n21151), .B(n21150), .Z(n21152) );
  NANDN U27227 ( .A(n21153), .B(n21152), .Z(n21154) );
  OR U27228 ( .A(n21155), .B(n21154), .Z(n21156) );
  AND U27229 ( .A(n21157), .B(n21156), .Z(n21159) );
  NAND U27230 ( .A(n21159), .B(n21158), .Z(n21161) );
  ANDN U27231 ( .B(n21161), .A(n21160), .Z(n21162) );
  NANDN U27232 ( .A(n21163), .B(n21162), .Z(n21167) );
  AND U27233 ( .A(n21165), .B(n21164), .Z(n21166) );
  NAND U27234 ( .A(n21167), .B(n21166), .Z(n21168) );
  NANDN U27235 ( .A(n21169), .B(n21168), .Z(n21171) );
  OR U27236 ( .A(n21171), .B(n21170), .Z(n21172) );
  NAND U27237 ( .A(n21173), .B(n21172), .Z(n21174) );
  NANDN U27238 ( .A(n21175), .B(n21174), .Z(n21176) );
  OR U27239 ( .A(n21177), .B(n21176), .Z(n21178) );
  AND U27240 ( .A(n21179), .B(n21178), .Z(n21181) );
  NAND U27241 ( .A(n21181), .B(n21180), .Z(n21183) );
  ANDN U27242 ( .B(n21183), .A(n21182), .Z(n21184) );
  NANDN U27243 ( .A(n21185), .B(n21184), .Z(n21189) );
  AND U27244 ( .A(n21187), .B(n21186), .Z(n21188) );
  NAND U27245 ( .A(n21189), .B(n21188), .Z(n21190) );
  NANDN U27246 ( .A(n21191), .B(n21190), .Z(n21193) );
  OR U27247 ( .A(n21193), .B(n21192), .Z(n21194) );
  NAND U27248 ( .A(n21195), .B(n21194), .Z(n21196) );
  NANDN U27249 ( .A(n21197), .B(n21196), .Z(n21198) );
  OR U27250 ( .A(n21199), .B(n21198), .Z(n21200) );
  AND U27251 ( .A(n21201), .B(n21200), .Z(n21202) );
  NANDN U27252 ( .A(n21203), .B(n21202), .Z(n21204) );
  AND U27253 ( .A(n21205), .B(n21204), .Z(n21210) );
  OR U27254 ( .A(n21207), .B(n21206), .Z(n21208) );
  AND U27255 ( .A(n28608), .B(n21208), .Z(n21209) );
  NANDN U27256 ( .A(n21210), .B(n21209), .Z(n21211) );
  NANDN U27257 ( .A(n28609), .B(n21211), .Z(n21212) );
  AND U27258 ( .A(n21212), .B(n28610), .Z(n21213) );
  OR U27259 ( .A(n21214), .B(n21213), .Z(n21215) );
  AND U27260 ( .A(n21216), .B(n21215), .Z(n21217) );
  ANDN U27261 ( .B(n21218), .A(n21217), .Z(n21219) );
  NAND U27262 ( .A(n21220), .B(n21219), .Z(n21221) );
  NANDN U27263 ( .A(n21222), .B(n21221), .Z(n21223) );
  OR U27264 ( .A(n21223), .B(n28613), .Z(n21229) );
  OR U27265 ( .A(n21225), .B(n21224), .Z(n21226) );
  AND U27266 ( .A(n21227), .B(n21226), .Z(n21228) );
  ANDN U27267 ( .B(n21229), .A(n21228), .Z(n21231) );
  XNOR U27268 ( .A(x[3151]), .B(y[3151]), .Z(n21230) );
  NANDN U27269 ( .A(n21231), .B(n21230), .Z(n21232) );
  NAND U27270 ( .A(n21233), .B(n21232), .Z(n21237) );
  AND U27271 ( .A(n21235), .B(n21234), .Z(n21236) );
  NAND U27272 ( .A(n21237), .B(n21236), .Z(n21238) );
  NANDN U27273 ( .A(n21239), .B(n21238), .Z(n21241) );
  OR U27274 ( .A(n21241), .B(n21240), .Z(n21242) );
  NAND U27275 ( .A(n21243), .B(n21242), .Z(n21244) );
  NANDN U27276 ( .A(n21245), .B(n21244), .Z(n21246) );
  OR U27277 ( .A(n21247), .B(n21246), .Z(n21248) );
  AND U27278 ( .A(n21249), .B(n21248), .Z(n21251) );
  NAND U27279 ( .A(n21251), .B(n21250), .Z(n21253) );
  ANDN U27280 ( .B(n21253), .A(n21252), .Z(n21254) );
  NANDN U27281 ( .A(n21255), .B(n21254), .Z(n21259) );
  AND U27282 ( .A(n21257), .B(n21256), .Z(n21258) );
  NAND U27283 ( .A(n21259), .B(n21258), .Z(n21260) );
  NANDN U27284 ( .A(n21261), .B(n21260), .Z(n21263) );
  OR U27285 ( .A(n21263), .B(n21262), .Z(n21264) );
  NAND U27286 ( .A(n21265), .B(n21264), .Z(n21266) );
  NANDN U27287 ( .A(n21267), .B(n21266), .Z(n21268) );
  OR U27288 ( .A(n21269), .B(n21268), .Z(n21270) );
  AND U27289 ( .A(n21271), .B(n21270), .Z(n21272) );
  NANDN U27290 ( .A(n21273), .B(n21272), .Z(n21274) );
  AND U27291 ( .A(n21275), .B(n21274), .Z(n21277) );
  NOR U27292 ( .A(n21277), .B(n21276), .Z(n21278) );
  NANDN U27293 ( .A(n21279), .B(n21278), .Z(n21280) );
  AND U27294 ( .A(n21281), .B(n21280), .Z(n21283) );
  AND U27295 ( .A(n21283), .B(n21282), .Z(n21287) );
  AND U27296 ( .A(n21285), .B(n21284), .Z(n21286) );
  NANDN U27297 ( .A(n21287), .B(n21286), .Z(n21288) );
  NANDN U27298 ( .A(n21289), .B(n21288), .Z(n21290) );
  AND U27299 ( .A(n21291), .B(n21290), .Z(n21293) );
  NAND U27300 ( .A(n21293), .B(n21292), .Z(n21294) );
  NANDN U27301 ( .A(n21295), .B(n21294), .Z(n21296) );
  AND U27302 ( .A(n21297), .B(n21296), .Z(n21299) );
  NAND U27303 ( .A(n21299), .B(n21298), .Z(n21300) );
  NANDN U27304 ( .A(n21301), .B(n21300), .Z(n21302) );
  AND U27305 ( .A(n21303), .B(n21302), .Z(n21305) );
  AND U27306 ( .A(n21305), .B(n21304), .Z(n21309) );
  NAND U27307 ( .A(n21307), .B(n21306), .Z(n21308) );
  OR U27308 ( .A(n21309), .B(n21308), .Z(n21310) );
  AND U27309 ( .A(n21311), .B(n21310), .Z(n21315) );
  NAND U27310 ( .A(n21313), .B(n21312), .Z(n21314) );
  OR U27311 ( .A(n21315), .B(n21314), .Z(n21316) );
  AND U27312 ( .A(n21317), .B(n21316), .Z(n21321) );
  NAND U27313 ( .A(n21319), .B(n21318), .Z(n21320) );
  OR U27314 ( .A(n21321), .B(n21320), .Z(n21322) );
  AND U27315 ( .A(n21323), .B(n21322), .Z(n21327) );
  NAND U27316 ( .A(n21325), .B(n21324), .Z(n21326) );
  OR U27317 ( .A(n21327), .B(n21326), .Z(n21328) );
  AND U27318 ( .A(n21329), .B(n21328), .Z(n21333) );
  NAND U27319 ( .A(n21331), .B(n21330), .Z(n21332) );
  OR U27320 ( .A(n21333), .B(n21332), .Z(n21334) );
  AND U27321 ( .A(n21335), .B(n21334), .Z(n21339) );
  NAND U27322 ( .A(n21337), .B(n21336), .Z(n21338) );
  OR U27323 ( .A(n21339), .B(n21338), .Z(n21340) );
  AND U27324 ( .A(n21341), .B(n21340), .Z(n21345) );
  NAND U27325 ( .A(n21343), .B(n21342), .Z(n21344) );
  OR U27326 ( .A(n21345), .B(n21344), .Z(n21346) );
  AND U27327 ( .A(n21347), .B(n21346), .Z(n21351) );
  NAND U27328 ( .A(n21349), .B(n21348), .Z(n21350) );
  OR U27329 ( .A(n21351), .B(n21350), .Z(n21352) );
  AND U27330 ( .A(n21353), .B(n21352), .Z(n21357) );
  NAND U27331 ( .A(n21355), .B(n21354), .Z(n21356) );
  OR U27332 ( .A(n21357), .B(n21356), .Z(n21358) );
  AND U27333 ( .A(n21359), .B(n21358), .Z(n21363) );
  NAND U27334 ( .A(n21361), .B(n21360), .Z(n21362) );
  OR U27335 ( .A(n21363), .B(n21362), .Z(n21364) );
  AND U27336 ( .A(n21365), .B(n21364), .Z(n21369) );
  NAND U27337 ( .A(n21367), .B(n21366), .Z(n21368) );
  OR U27338 ( .A(n21369), .B(n21368), .Z(n21370) );
  AND U27339 ( .A(n21371), .B(n21370), .Z(n21375) );
  NAND U27340 ( .A(n21373), .B(n21372), .Z(n21374) );
  OR U27341 ( .A(n21375), .B(n21374), .Z(n21376) );
  AND U27342 ( .A(n21377), .B(n21376), .Z(n21378) );
  NOR U27343 ( .A(n21379), .B(n21378), .Z(n21380) );
  NAND U27344 ( .A(n21381), .B(n21380), .Z(n21382) );
  NANDN U27345 ( .A(n21383), .B(n21382), .Z(n21384) );
  NAND U27346 ( .A(n21385), .B(n21384), .Z(n21386) );
  NANDN U27347 ( .A(n21387), .B(n21386), .Z(n21388) );
  AND U27348 ( .A(n21389), .B(n21388), .Z(n21391) );
  NAND U27349 ( .A(n21391), .B(n21390), .Z(n21392) );
  NANDN U27350 ( .A(n21393), .B(n21392), .Z(n21394) );
  AND U27351 ( .A(n21395), .B(n21394), .Z(n21397) );
  NAND U27352 ( .A(n21397), .B(n21396), .Z(n21398) );
  NANDN U27353 ( .A(n21399), .B(n21398), .Z(n21400) );
  AND U27354 ( .A(n21401), .B(n21400), .Z(n21402) );
  NANDN U27355 ( .A(n21403), .B(n21402), .Z(n21404) );
  NAND U27356 ( .A(n21405), .B(n21404), .Z(n21406) );
  NANDN U27357 ( .A(n21407), .B(n21406), .Z(n21409) );
  OR U27358 ( .A(n21409), .B(n21408), .Z(n21410) );
  NAND U27359 ( .A(n21411), .B(n21410), .Z(n21415) );
  NAND U27360 ( .A(n21413), .B(n21412), .Z(n21414) );
  ANDN U27361 ( .B(n21415), .A(n21414), .Z(n21419) );
  NAND U27362 ( .A(n21417), .B(n21416), .Z(n21418) );
  OR U27363 ( .A(n21419), .B(n21418), .Z(n21420) );
  AND U27364 ( .A(n21421), .B(n21420), .Z(n21425) );
  NAND U27365 ( .A(n21423), .B(n21422), .Z(n21424) );
  OR U27366 ( .A(n21425), .B(n21424), .Z(n21426) );
  AND U27367 ( .A(n21427), .B(n21426), .Z(n21428) );
  NOR U27368 ( .A(n21429), .B(n21428), .Z(n21430) );
  NAND U27369 ( .A(n21431), .B(n21430), .Z(n21432) );
  NANDN U27370 ( .A(n21433), .B(n21432), .Z(n21434) );
  NAND U27371 ( .A(n21435), .B(n21434), .Z(n21436) );
  NANDN U27372 ( .A(n21437), .B(n21436), .Z(n21438) );
  AND U27373 ( .A(n21439), .B(n21438), .Z(n21441) );
  NAND U27374 ( .A(n21441), .B(n21440), .Z(n21442) );
  NANDN U27375 ( .A(n21443), .B(n21442), .Z(n21444) );
  AND U27376 ( .A(n21445), .B(n21444), .Z(n21447) );
  NAND U27377 ( .A(n21447), .B(n21446), .Z(n21448) );
  NANDN U27378 ( .A(n21449), .B(n21448), .Z(n21450) );
  AND U27379 ( .A(n21451), .B(n21450), .Z(n21453) );
  AND U27380 ( .A(n21453), .B(n21452), .Z(n21457) );
  NAND U27381 ( .A(n21455), .B(n21454), .Z(n21456) );
  OR U27382 ( .A(n21457), .B(n21456), .Z(n21458) );
  AND U27383 ( .A(n21459), .B(n21458), .Z(n21463) );
  NAND U27384 ( .A(n21461), .B(n21460), .Z(n21462) );
  OR U27385 ( .A(n21463), .B(n21462), .Z(n21464) );
  AND U27386 ( .A(n21465), .B(n21464), .Z(n21469) );
  NAND U27387 ( .A(n21467), .B(n21466), .Z(n21468) );
  OR U27388 ( .A(n21469), .B(n21468), .Z(n21470) );
  AND U27389 ( .A(n21471), .B(n21470), .Z(n21475) );
  NAND U27390 ( .A(n21473), .B(n21472), .Z(n21474) );
  OR U27391 ( .A(n21475), .B(n21474), .Z(n21476) );
  AND U27392 ( .A(n21477), .B(n21476), .Z(n21481) );
  NAND U27393 ( .A(n21479), .B(n21478), .Z(n21480) );
  OR U27394 ( .A(n21481), .B(n21480), .Z(n21482) );
  AND U27395 ( .A(n21483), .B(n21482), .Z(n21487) );
  NAND U27396 ( .A(n21485), .B(n21484), .Z(n21486) );
  OR U27397 ( .A(n21487), .B(n21486), .Z(n21488) );
  AND U27398 ( .A(n21489), .B(n21488), .Z(n21493) );
  NAND U27399 ( .A(n21491), .B(n21490), .Z(n21492) );
  OR U27400 ( .A(n21493), .B(n21492), .Z(n21494) );
  AND U27401 ( .A(n21495), .B(n21494), .Z(n21499) );
  NAND U27402 ( .A(n21497), .B(n21496), .Z(n21498) );
  OR U27403 ( .A(n21499), .B(n21498), .Z(n21500) );
  AND U27404 ( .A(n21501), .B(n21500), .Z(n21505) );
  NAND U27405 ( .A(n21503), .B(n21502), .Z(n21504) );
  OR U27406 ( .A(n21505), .B(n21504), .Z(n21506) );
  AND U27407 ( .A(n21507), .B(n21506), .Z(n21511) );
  NAND U27408 ( .A(n21509), .B(n21508), .Z(n21510) );
  OR U27409 ( .A(n21511), .B(n21510), .Z(n21512) );
  AND U27410 ( .A(n21513), .B(n21512), .Z(n21517) );
  NAND U27411 ( .A(n21515), .B(n21514), .Z(n21516) );
  OR U27412 ( .A(n21517), .B(n21516), .Z(n21518) );
  AND U27413 ( .A(n21519), .B(n21518), .Z(n21523) );
  NAND U27414 ( .A(n21521), .B(n21520), .Z(n21522) );
  OR U27415 ( .A(n21523), .B(n21522), .Z(n21524) );
  AND U27416 ( .A(n21525), .B(n21524), .Z(n21526) );
  NOR U27417 ( .A(n21527), .B(n21526), .Z(n21528) );
  NAND U27418 ( .A(n21529), .B(n21528), .Z(n21533) );
  NAND U27419 ( .A(n21531), .B(n21530), .Z(n21532) );
  ANDN U27420 ( .B(n21533), .A(n21532), .Z(n21537) );
  NAND U27421 ( .A(n21535), .B(n21534), .Z(n21536) );
  OR U27422 ( .A(n21537), .B(n21536), .Z(n21538) );
  AND U27423 ( .A(n21539), .B(n21538), .Z(n21543) );
  NAND U27424 ( .A(n21541), .B(n21540), .Z(n21542) );
  OR U27425 ( .A(n21543), .B(n21542), .Z(n21544) );
  AND U27426 ( .A(n21545), .B(n21544), .Z(n21549) );
  NAND U27427 ( .A(n21547), .B(n21546), .Z(n21548) );
  OR U27428 ( .A(n21549), .B(n21548), .Z(n21550) );
  AND U27429 ( .A(n21551), .B(n21550), .Z(n21555) );
  NAND U27430 ( .A(n21553), .B(n21552), .Z(n21554) );
  OR U27431 ( .A(n21555), .B(n21554), .Z(n21556) );
  AND U27432 ( .A(n21557), .B(n21556), .Z(n21561) );
  NAND U27433 ( .A(n21559), .B(n21558), .Z(n21560) );
  OR U27434 ( .A(n21561), .B(n21560), .Z(n21562) );
  AND U27435 ( .A(n21563), .B(n21562), .Z(n21567) );
  NAND U27436 ( .A(n21565), .B(n21564), .Z(n21566) );
  OR U27437 ( .A(n21567), .B(n21566), .Z(n21568) );
  AND U27438 ( .A(n21569), .B(n21568), .Z(n21573) );
  NAND U27439 ( .A(n21571), .B(n21570), .Z(n21572) );
  OR U27440 ( .A(n21573), .B(n21572), .Z(n21574) );
  AND U27441 ( .A(n21575), .B(n21574), .Z(n21579) );
  NAND U27442 ( .A(n21577), .B(n21576), .Z(n21578) );
  OR U27443 ( .A(n21579), .B(n21578), .Z(n21580) );
  AND U27444 ( .A(n21581), .B(n21580), .Z(n21585) );
  NAND U27445 ( .A(n21583), .B(n21582), .Z(n21584) );
  OR U27446 ( .A(n21585), .B(n21584), .Z(n21586) );
  AND U27447 ( .A(n21587), .B(n21586), .Z(n21591) );
  NAND U27448 ( .A(n21589), .B(n21588), .Z(n21590) );
  OR U27449 ( .A(n21591), .B(n21590), .Z(n21592) );
  AND U27450 ( .A(n21593), .B(n21592), .Z(n21597) );
  NAND U27451 ( .A(n21595), .B(n21594), .Z(n21596) );
  OR U27452 ( .A(n21597), .B(n21596), .Z(n21598) );
  AND U27453 ( .A(n21599), .B(n21598), .Z(n21603) );
  NAND U27454 ( .A(n21601), .B(n21600), .Z(n21602) );
  OR U27455 ( .A(n21603), .B(n21602), .Z(n21604) );
  AND U27456 ( .A(n21605), .B(n21604), .Z(n21609) );
  NAND U27457 ( .A(n21607), .B(n21606), .Z(n21608) );
  OR U27458 ( .A(n21609), .B(n21608), .Z(n21610) );
  AND U27459 ( .A(n21611), .B(n21610), .Z(n21615) );
  NAND U27460 ( .A(n21613), .B(n21612), .Z(n21614) );
  OR U27461 ( .A(n21615), .B(n21614), .Z(n21616) );
  AND U27462 ( .A(n21617), .B(n21616), .Z(n21618) );
  NOR U27463 ( .A(n21619), .B(n21618), .Z(n21620) );
  NAND U27464 ( .A(n21621), .B(n21620), .Z(n21625) );
  NAND U27465 ( .A(n21623), .B(n21622), .Z(n21624) );
  ANDN U27466 ( .B(n21625), .A(n21624), .Z(n21629) );
  NAND U27467 ( .A(n21627), .B(n21626), .Z(n21628) );
  OR U27468 ( .A(n21629), .B(n21628), .Z(n21630) );
  AND U27469 ( .A(n21631), .B(n21630), .Z(n21635) );
  NAND U27470 ( .A(n21633), .B(n21632), .Z(n21634) );
  OR U27471 ( .A(n21635), .B(n21634), .Z(n21636) );
  AND U27472 ( .A(n21637), .B(n21636), .Z(n21641) );
  NAND U27473 ( .A(n21639), .B(n21638), .Z(n21640) );
  OR U27474 ( .A(n21641), .B(n21640), .Z(n21642) );
  AND U27475 ( .A(n21643), .B(n21642), .Z(n21644) );
  ANDN U27476 ( .B(n21645), .A(n21644), .Z(n21646) );
  NAND U27477 ( .A(n21647), .B(n21646), .Z(n21648) );
  NANDN U27478 ( .A(n21649), .B(n21648), .Z(n21650) );
  OR U27479 ( .A(n21651), .B(n21650), .Z(n21652) );
  AND U27480 ( .A(n21653), .B(n21652), .Z(n21655) );
  NAND U27481 ( .A(n21655), .B(n21654), .Z(n21656) );
  NANDN U27482 ( .A(n21657), .B(n21656), .Z(n21658) );
  AND U27483 ( .A(n21659), .B(n21658), .Z(n21661) );
  NAND U27484 ( .A(n21661), .B(n21660), .Z(n21662) );
  NANDN U27485 ( .A(n21663), .B(n21662), .Z(n21664) );
  AND U27486 ( .A(n21665), .B(n21664), .Z(n21667) );
  AND U27487 ( .A(n21667), .B(n21666), .Z(n21671) );
  NAND U27488 ( .A(n21669), .B(n21668), .Z(n21670) );
  OR U27489 ( .A(n21671), .B(n21670), .Z(n21672) );
  AND U27490 ( .A(n21673), .B(n21672), .Z(n21677) );
  NAND U27491 ( .A(n21675), .B(n21674), .Z(n21676) );
  OR U27492 ( .A(n21677), .B(n21676), .Z(n21678) );
  AND U27493 ( .A(n21679), .B(n21678), .Z(n21683) );
  NAND U27494 ( .A(n21681), .B(n21680), .Z(n21682) );
  OR U27495 ( .A(n21683), .B(n21682), .Z(n21684) );
  AND U27496 ( .A(n21685), .B(n21684), .Z(n21686) );
  OR U27497 ( .A(n21687), .B(n21686), .Z(n21688) );
  NAND U27498 ( .A(n21689), .B(n21688), .Z(n21690) );
  AND U27499 ( .A(n21691), .B(n21690), .Z(n21695) );
  AND U27500 ( .A(n21693), .B(n21692), .Z(n21694) );
  NANDN U27501 ( .A(n21695), .B(n21694), .Z(n21698) );
  NANDN U27502 ( .A(x[3302]), .B(y[3302]), .Z(n24044) );
  AND U27503 ( .A(n21696), .B(n24044), .Z(n21697) );
  NAND U27504 ( .A(n21698), .B(n21697), .Z(n21699) );
  NANDN U27505 ( .A(n21700), .B(n21699), .Z(n21701) );
  AND U27506 ( .A(n21702), .B(n21701), .Z(n21703) );
  OR U27507 ( .A(n21704), .B(n21703), .Z(n21705) );
  NAND U27508 ( .A(n21706), .B(n21705), .Z(n21710) );
  NAND U27509 ( .A(n21708), .B(n21707), .Z(n21709) );
  ANDN U27510 ( .B(n21710), .A(n21709), .Z(n21714) );
  NAND U27511 ( .A(n21712), .B(n21711), .Z(n21713) );
  OR U27512 ( .A(n21714), .B(n21713), .Z(n21715) );
  AND U27513 ( .A(n21716), .B(n21715), .Z(n21720) );
  NAND U27514 ( .A(n21718), .B(n21717), .Z(n21719) );
  OR U27515 ( .A(n21720), .B(n21719), .Z(n21721) );
  AND U27516 ( .A(n21722), .B(n21721), .Z(n21728) );
  OR U27517 ( .A(n21724), .B(n21723), .Z(n21725) );
  AND U27518 ( .A(n21726), .B(n21725), .Z(n21727) );
  OR U27519 ( .A(n21728), .B(n21727), .Z(n21729) );
  AND U27520 ( .A(n21730), .B(n21729), .Z(n21731) );
  OR U27521 ( .A(n21732), .B(n21731), .Z(n21733) );
  NAND U27522 ( .A(n21734), .B(n21733), .Z(n21735) );
  NANDN U27523 ( .A(n21736), .B(n21735), .Z(n21737) );
  ANDN U27524 ( .B(y[3316]), .A(x[3316]), .Z(n28755) );
  OR U27525 ( .A(n21737), .B(n28755), .Z(n21738) );
  NAND U27526 ( .A(n21739), .B(n21738), .Z(n21740) );
  NANDN U27527 ( .A(n21741), .B(n21740), .Z(n21743) );
  OR U27528 ( .A(n21743), .B(n21742), .Z(n21744) );
  NAND U27529 ( .A(n21745), .B(n21744), .Z(n21746) );
  NANDN U27530 ( .A(n21747), .B(n21746), .Z(n21748) );
  AND U27531 ( .A(n21749), .B(n21748), .Z(n21750) );
  NAND U27532 ( .A(n21751), .B(n21750), .Z(n21755) );
  NAND U27533 ( .A(n21753), .B(n21752), .Z(n21754) );
  ANDN U27534 ( .B(n21755), .A(n21754), .Z(n21759) );
  NAND U27535 ( .A(n21757), .B(n21756), .Z(n21758) );
  OR U27536 ( .A(n21759), .B(n21758), .Z(n21760) );
  AND U27537 ( .A(n21761), .B(n21760), .Z(n21765) );
  NAND U27538 ( .A(n21763), .B(n21762), .Z(n21764) );
  OR U27539 ( .A(n21765), .B(n21764), .Z(n21766) );
  AND U27540 ( .A(n21767), .B(n21766), .Z(n21771) );
  NAND U27541 ( .A(n21769), .B(n21768), .Z(n21770) );
  OR U27542 ( .A(n21771), .B(n21770), .Z(n21772) );
  AND U27543 ( .A(n21773), .B(n21772), .Z(n21777) );
  NAND U27544 ( .A(n21775), .B(n21774), .Z(n21776) );
  OR U27545 ( .A(n21777), .B(n21776), .Z(n21778) );
  AND U27546 ( .A(n21779), .B(n21778), .Z(n21783) );
  NAND U27547 ( .A(n21781), .B(n21780), .Z(n21782) );
  OR U27548 ( .A(n21783), .B(n21782), .Z(n21784) );
  AND U27549 ( .A(n21785), .B(n21784), .Z(n21789) );
  NAND U27550 ( .A(n21787), .B(n21786), .Z(n21788) );
  OR U27551 ( .A(n21789), .B(n21788), .Z(n21790) );
  AND U27552 ( .A(n21791), .B(n21790), .Z(n21792) );
  NOR U27553 ( .A(n21793), .B(n21792), .Z(n21794) );
  NAND U27554 ( .A(n21795), .B(n21794), .Z(n21799) );
  NAND U27555 ( .A(n21797), .B(n21796), .Z(n21798) );
  ANDN U27556 ( .B(n21799), .A(n21798), .Z(n21803) );
  NAND U27557 ( .A(n21801), .B(n21800), .Z(n21802) );
  OR U27558 ( .A(n21803), .B(n21802), .Z(n21804) );
  AND U27559 ( .A(n21805), .B(n21804), .Z(n21809) );
  NAND U27560 ( .A(n21807), .B(n21806), .Z(n21808) );
  OR U27561 ( .A(n21809), .B(n21808), .Z(n21810) );
  AND U27562 ( .A(n21811), .B(n21810), .Z(n21815) );
  NAND U27563 ( .A(n21813), .B(n21812), .Z(n21814) );
  OR U27564 ( .A(n21815), .B(n21814), .Z(n21816) );
  AND U27565 ( .A(n21817), .B(n21816), .Z(n21821) );
  NAND U27566 ( .A(n21819), .B(n21818), .Z(n21820) );
  OR U27567 ( .A(n21821), .B(n21820), .Z(n21822) );
  AND U27568 ( .A(n21823), .B(n21822), .Z(n21827) );
  NAND U27569 ( .A(n21825), .B(n21824), .Z(n21826) );
  OR U27570 ( .A(n21827), .B(n21826), .Z(n21828) );
  AND U27571 ( .A(n21829), .B(n21828), .Z(n21830) );
  OR U27572 ( .A(n21831), .B(n21830), .Z(n21832) );
  NAND U27573 ( .A(n21833), .B(n21832), .Z(n21834) );
  AND U27574 ( .A(n21835), .B(n21834), .Z(n21840) );
  OR U27575 ( .A(n21837), .B(n21836), .Z(n21838) );
  AND U27576 ( .A(n21838), .B(n24029), .Z(n21839) );
  NANDN U27577 ( .A(n21840), .B(n21839), .Z(n21841) );
  NANDN U27578 ( .A(n28786), .B(n21841), .Z(n21842) );
  AND U27579 ( .A(n21843), .B(n21842), .Z(n21844) );
  OR U27580 ( .A(n21845), .B(n21844), .Z(n21846) );
  NAND U27581 ( .A(n21847), .B(n21846), .Z(n21851) );
  NAND U27582 ( .A(n21849), .B(n21848), .Z(n21850) );
  ANDN U27583 ( .B(n21851), .A(n21850), .Z(n21855) );
  NAND U27584 ( .A(n21853), .B(n21852), .Z(n21854) );
  OR U27585 ( .A(n21855), .B(n21854), .Z(n21856) );
  AND U27586 ( .A(n21857), .B(n21856), .Z(n21861) );
  NAND U27587 ( .A(n21859), .B(n21858), .Z(n21860) );
  OR U27588 ( .A(n21861), .B(n21860), .Z(n21862) );
  AND U27589 ( .A(n21863), .B(n21862), .Z(n21867) );
  NAND U27590 ( .A(n21865), .B(n21864), .Z(n21866) );
  OR U27591 ( .A(n21867), .B(n21866), .Z(n21868) );
  AND U27592 ( .A(n21869), .B(n21868), .Z(n21870) );
  OR U27593 ( .A(n21871), .B(n21870), .Z(n21872) );
  NAND U27594 ( .A(n21873), .B(n21872), .Z(n21874) );
  NANDN U27595 ( .A(n28798), .B(n21874), .Z(n21875) );
  ANDN U27596 ( .B(y[3364]), .A(x[3364]), .Z(n24024) );
  OR U27597 ( .A(n21875), .B(n24024), .Z(n21876) );
  NAND U27598 ( .A(n21877), .B(n21876), .Z(n21878) );
  NANDN U27599 ( .A(n21879), .B(n21878), .Z(n21880) );
  ANDN U27600 ( .B(y[3366]), .A(x[3366]), .Z(n28799) );
  OR U27601 ( .A(n21880), .B(n28799), .Z(n21881) );
  NAND U27602 ( .A(n21882), .B(n21881), .Z(n21883) );
  NANDN U27603 ( .A(n21884), .B(n21883), .Z(n21886) );
  OR U27604 ( .A(n21886), .B(n21885), .Z(n21887) );
  NAND U27605 ( .A(n21888), .B(n21887), .Z(n21892) );
  NAND U27606 ( .A(n21890), .B(n21889), .Z(n21891) );
  ANDN U27607 ( .B(n21892), .A(n21891), .Z(n21896) );
  NAND U27608 ( .A(n21894), .B(n21893), .Z(n21895) );
  OR U27609 ( .A(n21896), .B(n21895), .Z(n21897) );
  AND U27610 ( .A(n21898), .B(n21897), .Z(n21902) );
  NAND U27611 ( .A(n21900), .B(n21899), .Z(n21901) );
  OR U27612 ( .A(n21902), .B(n21901), .Z(n21903) );
  AND U27613 ( .A(n21904), .B(n21903), .Z(n21908) );
  NAND U27614 ( .A(n21906), .B(n21905), .Z(n21907) );
  OR U27615 ( .A(n21908), .B(n21907), .Z(n21909) );
  AND U27616 ( .A(n21910), .B(n21909), .Z(n21914) );
  NAND U27617 ( .A(n21912), .B(n21911), .Z(n21913) );
  OR U27618 ( .A(n21914), .B(n21913), .Z(n21915) );
  AND U27619 ( .A(n21916), .B(n21915), .Z(n21920) );
  NAND U27620 ( .A(n21918), .B(n21917), .Z(n21919) );
  OR U27621 ( .A(n21920), .B(n21919), .Z(n21921) );
  AND U27622 ( .A(n21922), .B(n21921), .Z(n21926) );
  NAND U27623 ( .A(n21924), .B(n21923), .Z(n21925) );
  OR U27624 ( .A(n21926), .B(n21925), .Z(n21927) );
  AND U27625 ( .A(n21928), .B(n21927), .Z(n21932) );
  NAND U27626 ( .A(n21930), .B(n21929), .Z(n21931) );
  OR U27627 ( .A(n21932), .B(n21931), .Z(n21933) );
  AND U27628 ( .A(n21934), .B(n21933), .Z(n21938) );
  NAND U27629 ( .A(n21936), .B(n21935), .Z(n21937) );
  OR U27630 ( .A(n21938), .B(n21937), .Z(n21939) );
  AND U27631 ( .A(n21940), .B(n21939), .Z(n21941) );
  OR U27632 ( .A(n21942), .B(n21941), .Z(n21943) );
  NAND U27633 ( .A(n21944), .B(n21943), .Z(n21945) );
  NANDN U27634 ( .A(n21946), .B(n21945), .Z(n21947) );
  AND U27635 ( .A(n21947), .B(n24018), .Z(n21948) );
  OR U27636 ( .A(n21948), .B(n28822), .Z(n21949) );
  NAND U27637 ( .A(n28823), .B(n21949), .Z(n21950) );
  NANDN U27638 ( .A(n28824), .B(n21950), .Z(n21951) );
  AND U27639 ( .A(n21951), .B(n28825), .Z(n21952) );
  OR U27640 ( .A(n21953), .B(n21952), .Z(n21954) );
  NAND U27641 ( .A(n21955), .B(n21954), .Z(n21956) );
  NANDN U27642 ( .A(n21957), .B(n21956), .Z(n21959) );
  NANDN U27643 ( .A(n21959), .B(n21958), .Z(n21960) );
  AND U27644 ( .A(n21961), .B(n21960), .Z(n21962) );
  NOR U27645 ( .A(n21963), .B(n21962), .Z(n21965) );
  NAND U27646 ( .A(n21965), .B(n21964), .Z(n21966) );
  AND U27647 ( .A(n21966), .B(n28829), .Z(n21967) );
  NANDN U27648 ( .A(n24013), .B(n21967), .Z(n21968) );
  NAND U27649 ( .A(n21969), .B(n21968), .Z(n21970) );
  NANDN U27650 ( .A(n21971), .B(n21970), .Z(n21972) );
  ANDN U27651 ( .B(y[3400]), .A(x[3400]), .Z(n28830) );
  OR U27652 ( .A(n21972), .B(n28830), .Z(n21973) );
  NAND U27653 ( .A(n21974), .B(n21973), .Z(n21975) );
  NANDN U27654 ( .A(n21976), .B(n21975), .Z(n21978) );
  OR U27655 ( .A(n21978), .B(n21977), .Z(n21979) );
  NANDN U27656 ( .A(n21980), .B(n21979), .Z(n21981) );
  AND U27657 ( .A(n21982), .B(n21981), .Z(n21986) );
  NAND U27658 ( .A(n21984), .B(n21983), .Z(n21985) );
  OR U27659 ( .A(n21986), .B(n21985), .Z(n21987) );
  AND U27660 ( .A(n21988), .B(n21987), .Z(n21992) );
  NAND U27661 ( .A(n21990), .B(n21989), .Z(n21991) );
  OR U27662 ( .A(n21992), .B(n21991), .Z(n21993) );
  AND U27663 ( .A(n21994), .B(n21993), .Z(n21998) );
  NAND U27664 ( .A(n21996), .B(n21995), .Z(n21997) );
  OR U27665 ( .A(n21998), .B(n21997), .Z(n21999) );
  AND U27666 ( .A(n22000), .B(n21999), .Z(n22004) );
  NAND U27667 ( .A(n22002), .B(n22001), .Z(n22003) );
  OR U27668 ( .A(n22004), .B(n22003), .Z(n22005) );
  AND U27669 ( .A(n22006), .B(n22005), .Z(n22010) );
  NAND U27670 ( .A(n22008), .B(n22007), .Z(n22009) );
  OR U27671 ( .A(n22010), .B(n22009), .Z(n22011) );
  AND U27672 ( .A(n22012), .B(n22011), .Z(n22016) );
  NAND U27673 ( .A(n22014), .B(n22013), .Z(n22015) );
  OR U27674 ( .A(n22016), .B(n22015), .Z(n22017) );
  AND U27675 ( .A(n22018), .B(n22017), .Z(n22022) );
  NAND U27676 ( .A(n22020), .B(n22019), .Z(n22021) );
  OR U27677 ( .A(n22022), .B(n22021), .Z(n22023) );
  AND U27678 ( .A(n22024), .B(n22023), .Z(n22028) );
  NAND U27679 ( .A(n22026), .B(n22025), .Z(n22027) );
  OR U27680 ( .A(n22028), .B(n22027), .Z(n22029) );
  AND U27681 ( .A(n22030), .B(n22029), .Z(n22034) );
  NAND U27682 ( .A(n22032), .B(n22031), .Z(n22033) );
  OR U27683 ( .A(n22034), .B(n22033), .Z(n22035) );
  AND U27684 ( .A(n22036), .B(n22035), .Z(n22040) );
  NAND U27685 ( .A(n22038), .B(n22037), .Z(n22039) );
  OR U27686 ( .A(n22040), .B(n22039), .Z(n22041) );
  AND U27687 ( .A(n22042), .B(n22041), .Z(n22046) );
  NAND U27688 ( .A(n22044), .B(n22043), .Z(n22045) );
  OR U27689 ( .A(n22046), .B(n22045), .Z(n22047) );
  AND U27690 ( .A(n22048), .B(n22047), .Z(n22052) );
  NAND U27691 ( .A(n22050), .B(n22049), .Z(n22051) );
  OR U27692 ( .A(n22052), .B(n22051), .Z(n22053) );
  AND U27693 ( .A(n22054), .B(n22053), .Z(n22058) );
  NAND U27694 ( .A(n22056), .B(n22055), .Z(n22057) );
  OR U27695 ( .A(n22058), .B(n22057), .Z(n22059) );
  AND U27696 ( .A(n22060), .B(n22059), .Z(n22061) );
  OR U27697 ( .A(n22062), .B(n22061), .Z(n22063) );
  NAND U27698 ( .A(n22064), .B(n22063), .Z(n22065) );
  AND U27699 ( .A(n22066), .B(n22065), .Z(n22067) );
  NOR U27700 ( .A(n28856), .B(n22067), .Z(n22068) );
  NANDN U27701 ( .A(n22069), .B(n22068), .Z(n22070) );
  AND U27702 ( .A(n22071), .B(n22070), .Z(n22073) );
  NAND U27703 ( .A(n22073), .B(n22072), .Z(n22074) );
  NANDN U27704 ( .A(n22075), .B(n22074), .Z(n22076) );
  AND U27705 ( .A(n22077), .B(n22076), .Z(n22079) );
  NAND U27706 ( .A(n22079), .B(n22078), .Z(n22080) );
  NANDN U27707 ( .A(n22081), .B(n22080), .Z(n22082) );
  AND U27708 ( .A(n22083), .B(n22082), .Z(n22085) );
  NAND U27709 ( .A(n22085), .B(n22084), .Z(n22086) );
  NANDN U27710 ( .A(n22087), .B(n22086), .Z(n22088) );
  AND U27711 ( .A(n22089), .B(n22088), .Z(n22091) );
  AND U27712 ( .A(n22091), .B(n22090), .Z(n22095) );
  NAND U27713 ( .A(n22093), .B(n22092), .Z(n22094) );
  OR U27714 ( .A(n22095), .B(n22094), .Z(n22096) );
  AND U27715 ( .A(n22097), .B(n22096), .Z(n22101) );
  NAND U27716 ( .A(n22099), .B(n22098), .Z(n22100) );
  OR U27717 ( .A(n22101), .B(n22100), .Z(n22102) );
  AND U27718 ( .A(n22103), .B(n22102), .Z(n22104) );
  OR U27719 ( .A(n22105), .B(n22104), .Z(n22106) );
  NAND U27720 ( .A(n22107), .B(n22106), .Z(n22108) );
  AND U27721 ( .A(n22109), .B(n22108), .Z(n22113) );
  AND U27722 ( .A(n22111), .B(n22110), .Z(n22112) );
  NANDN U27723 ( .A(n22113), .B(n22112), .Z(n22116) );
  NANDN U27724 ( .A(x[3450]), .B(y[3450]), .Z(n23997) );
  AND U27725 ( .A(n22114), .B(n23997), .Z(n22115) );
  NAND U27726 ( .A(n22116), .B(n22115), .Z(n22117) );
  NANDN U27727 ( .A(n22118), .B(n22117), .Z(n22119) );
  NAND U27728 ( .A(n22120), .B(n22119), .Z(n22121) );
  NAND U27729 ( .A(n22122), .B(n22121), .Z(n22123) );
  NANDN U27730 ( .A(n22124), .B(n22123), .Z(n22126) );
  OR U27731 ( .A(n22126), .B(n22125), .Z(n22127) );
  NAND U27732 ( .A(n22128), .B(n22127), .Z(n22129) );
  NANDN U27733 ( .A(n28876), .B(n22129), .Z(n22133) );
  AND U27734 ( .A(n22131), .B(n22130), .Z(n22132) );
  OR U27735 ( .A(n22133), .B(n22132), .Z(n22134) );
  NAND U27736 ( .A(n28877), .B(n22134), .Z(n22135) );
  NANDN U27737 ( .A(n22136), .B(n22135), .Z(n22138) );
  NAND U27738 ( .A(n22138), .B(n22137), .Z(n22139) );
  NANDN U27739 ( .A(n22140), .B(n22139), .Z(n22141) );
  AND U27740 ( .A(n22142), .B(n22141), .Z(n22146) );
  NAND U27741 ( .A(n22144), .B(n22143), .Z(n22145) );
  OR U27742 ( .A(n22146), .B(n22145), .Z(n22147) );
  AND U27743 ( .A(n22148), .B(n22147), .Z(n22152) );
  NAND U27744 ( .A(n22150), .B(n22149), .Z(n22151) );
  OR U27745 ( .A(n22152), .B(n22151), .Z(n22153) );
  AND U27746 ( .A(n22154), .B(n22153), .Z(n22155) );
  OR U27747 ( .A(n22156), .B(n22155), .Z(n22157) );
  NAND U27748 ( .A(n22158), .B(n22157), .Z(n22159) );
  AND U27749 ( .A(n22160), .B(n22159), .Z(n22161) );
  NOR U27750 ( .A(n22162), .B(n22161), .Z(n22164) );
  NAND U27751 ( .A(n22164), .B(n22163), .Z(n22166) );
  AND U27752 ( .A(n22166), .B(n22165), .Z(n22167) );
  NAND U27753 ( .A(n28888), .B(n22167), .Z(n22168) );
  NANDN U27754 ( .A(n22169), .B(n22168), .Z(n22170) );
  AND U27755 ( .A(n22171), .B(n22170), .Z(n22173) );
  NAND U27756 ( .A(n22173), .B(n22172), .Z(n22174) );
  NANDN U27757 ( .A(n22175), .B(n22174), .Z(n22176) );
  AND U27758 ( .A(n22177), .B(n22176), .Z(n22179) );
  NAND U27759 ( .A(n22179), .B(n22178), .Z(n22180) );
  NANDN U27760 ( .A(n22181), .B(n22180), .Z(n22182) );
  AND U27761 ( .A(n22183), .B(n22182), .Z(n22185) );
  NAND U27762 ( .A(n22185), .B(n22184), .Z(n22186) );
  NANDN U27763 ( .A(n22187), .B(n22186), .Z(n22188) );
  AND U27764 ( .A(n22189), .B(n22188), .Z(n22190) );
  NANDN U27765 ( .A(n22191), .B(n22190), .Z(n22192) );
  NAND U27766 ( .A(n22193), .B(n22192), .Z(n22194) );
  NANDN U27767 ( .A(n22195), .B(n22194), .Z(n22196) );
  NAND U27768 ( .A(n22197), .B(n22196), .Z(n22198) );
  NANDN U27769 ( .A(n22199), .B(n22198), .Z(n22200) );
  AND U27770 ( .A(n22201), .B(n22200), .Z(n22203) );
  NAND U27771 ( .A(n22203), .B(n22202), .Z(n22204) );
  NANDN U27772 ( .A(n22205), .B(n22204), .Z(n22206) );
  AND U27773 ( .A(n22207), .B(n22206), .Z(n22208) );
  NANDN U27774 ( .A(n22209), .B(n22208), .Z(n22210) );
  NAND U27775 ( .A(n22211), .B(n22210), .Z(n22212) );
  NANDN U27776 ( .A(n22213), .B(n22212), .Z(n22214) );
  AND U27777 ( .A(n22215), .B(n22214), .Z(n22216) );
  NAND U27778 ( .A(n22217), .B(n22216), .Z(n22221) );
  NAND U27779 ( .A(n22219), .B(n22218), .Z(n22220) );
  ANDN U27780 ( .B(n22221), .A(n22220), .Z(n22225) );
  NAND U27781 ( .A(n22223), .B(n22222), .Z(n22224) );
  OR U27782 ( .A(n22225), .B(n22224), .Z(n22226) );
  AND U27783 ( .A(n22227), .B(n22226), .Z(n22231) );
  NAND U27784 ( .A(n22229), .B(n22228), .Z(n22230) );
  OR U27785 ( .A(n22231), .B(n22230), .Z(n22232) );
  AND U27786 ( .A(n22233), .B(n22232), .Z(n22237) );
  NAND U27787 ( .A(n22235), .B(n22234), .Z(n22236) );
  OR U27788 ( .A(n22237), .B(n22236), .Z(n22238) );
  AND U27789 ( .A(n22239), .B(n22238), .Z(n22243) );
  NAND U27790 ( .A(n22241), .B(n22240), .Z(n22242) );
  OR U27791 ( .A(n22243), .B(n22242), .Z(n22244) );
  AND U27792 ( .A(n22245), .B(n22244), .Z(n22249) );
  NAND U27793 ( .A(n22247), .B(n22246), .Z(n22248) );
  OR U27794 ( .A(n22249), .B(n22248), .Z(n22250) );
  AND U27795 ( .A(n22251), .B(n22250), .Z(n22255) );
  NAND U27796 ( .A(n22253), .B(n22252), .Z(n22254) );
  OR U27797 ( .A(n22255), .B(n22254), .Z(n22256) );
  AND U27798 ( .A(n22257), .B(n22256), .Z(n22261) );
  NAND U27799 ( .A(n22259), .B(n22258), .Z(n22260) );
  OR U27800 ( .A(n22261), .B(n22260), .Z(n22262) );
  AND U27801 ( .A(n22263), .B(n22262), .Z(n22267) );
  NAND U27802 ( .A(n22265), .B(n22264), .Z(n22266) );
  OR U27803 ( .A(n22267), .B(n22266), .Z(n22268) );
  AND U27804 ( .A(n22269), .B(n22268), .Z(n22273) );
  NAND U27805 ( .A(n22271), .B(n22270), .Z(n22272) );
  OR U27806 ( .A(n22273), .B(n22272), .Z(n22274) );
  AND U27807 ( .A(n22275), .B(n22274), .Z(n22279) );
  NAND U27808 ( .A(n22277), .B(n22276), .Z(n22278) );
  OR U27809 ( .A(n22279), .B(n22278), .Z(n22280) );
  AND U27810 ( .A(n22281), .B(n22280), .Z(n22282) );
  OR U27811 ( .A(n22283), .B(n22282), .Z(n22284) );
  NAND U27812 ( .A(n22285), .B(n22284), .Z(n22286) );
  NAND U27813 ( .A(n22287), .B(n22286), .Z(n22288) );
  NANDN U27814 ( .A(n22289), .B(n22288), .Z(n22290) );
  AND U27815 ( .A(n23982), .B(n22290), .Z(n22292) );
  NAND U27816 ( .A(n22292), .B(n22291), .Z(n22293) );
  NANDN U27817 ( .A(n22294), .B(n22293), .Z(n22295) );
  AND U27818 ( .A(n28930), .B(n22295), .Z(n22297) );
  NAND U27819 ( .A(n22297), .B(n22296), .Z(n22298) );
  NANDN U27820 ( .A(n22299), .B(n22298), .Z(n22300) );
  AND U27821 ( .A(n22301), .B(n22300), .Z(n22302) );
  NANDN U27822 ( .A(n28931), .B(n22302), .Z(n22303) );
  NAND U27823 ( .A(n22304), .B(n22303), .Z(n22308) );
  IV U27824 ( .A(n22305), .Z(n28934) );
  NAND U27825 ( .A(n28934), .B(n22306), .Z(n22307) );
  ANDN U27826 ( .B(n22308), .A(n22307), .Z(n22309) );
  OR U27827 ( .A(n22310), .B(n22309), .Z(n22311) );
  NAND U27828 ( .A(n22312), .B(n22311), .Z(n22313) );
  NAND U27829 ( .A(n22314), .B(n22313), .Z(n22315) );
  NANDN U27830 ( .A(n22316), .B(n22315), .Z(n22317) );
  AND U27831 ( .A(n22318), .B(n22317), .Z(n22320) );
  NAND U27832 ( .A(n22320), .B(n22319), .Z(n22321) );
  NANDN U27833 ( .A(n22322), .B(n22321), .Z(n22323) );
  AND U27834 ( .A(n22324), .B(n22323), .Z(n22326) );
  NAND U27835 ( .A(n22326), .B(n22325), .Z(n22327) );
  NANDN U27836 ( .A(n22328), .B(n22327), .Z(n22329) );
  NAND U27837 ( .A(n22330), .B(n22329), .Z(n22333) );
  NANDN U27838 ( .A(x[3530]), .B(y[3530]), .Z(n28943) );
  AND U27839 ( .A(n22331), .B(n28943), .Z(n22332) );
  NAND U27840 ( .A(n22333), .B(n22332), .Z(n22334) );
  NANDN U27841 ( .A(n22335), .B(n22334), .Z(n22336) );
  NAND U27842 ( .A(n22337), .B(n22336), .Z(n22338) );
  NAND U27843 ( .A(n22339), .B(n22338), .Z(n22340) );
  NANDN U27844 ( .A(n22341), .B(n22340), .Z(n22342) );
  ANDN U27845 ( .B(y[3534]), .A(x[3534]), .Z(n23973) );
  OR U27846 ( .A(n22342), .B(n23973), .Z(n22343) );
  NAND U27847 ( .A(n22344), .B(n22343), .Z(n22345) );
  NANDN U27848 ( .A(n22346), .B(n22345), .Z(n22348) );
  OR U27849 ( .A(n22348), .B(n22347), .Z(n22349) );
  NANDN U27850 ( .A(n22350), .B(n22349), .Z(n22351) );
  AND U27851 ( .A(n22352), .B(n22351), .Z(n22356) );
  NAND U27852 ( .A(n22354), .B(n22353), .Z(n22355) );
  OR U27853 ( .A(n22356), .B(n22355), .Z(n22357) );
  AND U27854 ( .A(n22358), .B(n22357), .Z(n22362) );
  NAND U27855 ( .A(n22360), .B(n22359), .Z(n22361) );
  OR U27856 ( .A(n22362), .B(n22361), .Z(n22363) );
  AND U27857 ( .A(n22364), .B(n22363), .Z(n22368) );
  NAND U27858 ( .A(n22366), .B(n22365), .Z(n22367) );
  OR U27859 ( .A(n22368), .B(n22367), .Z(n22369) );
  AND U27860 ( .A(n22370), .B(n22369), .Z(n22374) );
  NAND U27861 ( .A(n22372), .B(n22371), .Z(n22373) );
  OR U27862 ( .A(n22374), .B(n22373), .Z(n22375) );
  AND U27863 ( .A(n22376), .B(n22375), .Z(n22377) );
  NOR U27864 ( .A(n22378), .B(n22377), .Z(n22379) );
  NAND U27865 ( .A(n22380), .B(n22379), .Z(n22381) );
  NANDN U27866 ( .A(n22382), .B(n22381), .Z(n22383) );
  NAND U27867 ( .A(n22384), .B(n22383), .Z(n22385) );
  NANDN U27868 ( .A(n22386), .B(n22385), .Z(n22387) );
  AND U27869 ( .A(n22388), .B(n22387), .Z(n22390) );
  NAND U27870 ( .A(n22390), .B(n22389), .Z(n22391) );
  NANDN U27871 ( .A(n22392), .B(n22391), .Z(n22393) );
  AND U27872 ( .A(n22394), .B(n22393), .Z(n22396) );
  NAND U27873 ( .A(n22396), .B(n22395), .Z(n22397) );
  NANDN U27874 ( .A(n22398), .B(n22397), .Z(n22399) );
  NAND U27875 ( .A(n22400), .B(n22399), .Z(n22403) );
  NANDN U27876 ( .A(y[3556]), .B(n22403), .Z(n22402) );
  ANDN U27877 ( .B(n22402), .A(n22401), .Z(n22406) );
  XNOR U27878 ( .A(y[3556]), .B(n22403), .Z(n22404) );
  NAND U27879 ( .A(n22404), .B(x[3556]), .Z(n22405) );
  NAND U27880 ( .A(n22406), .B(n22405), .Z(n22407) );
  NAND U27881 ( .A(n28971), .B(n22407), .Z(n22408) );
  NAND U27882 ( .A(n28972), .B(n22408), .Z(n22409) );
  NANDN U27883 ( .A(n28973), .B(n22409), .Z(n22410) );
  AND U27884 ( .A(n28975), .B(n22410), .Z(n22411) );
  OR U27885 ( .A(n22411), .B(n28976), .Z(n22412) );
  NAND U27886 ( .A(n22413), .B(n22412), .Z(n22414) );
  NANDN U27887 ( .A(n22415), .B(n22414), .Z(n22416) );
  AND U27888 ( .A(n22417), .B(n22416), .Z(n22418) );
  OR U27889 ( .A(n22419), .B(n22418), .Z(n22420) );
  NAND U27890 ( .A(n22421), .B(n22420), .Z(n22425) );
  NAND U27891 ( .A(n22423), .B(n22422), .Z(n22424) );
  ANDN U27892 ( .B(n22425), .A(n22424), .Z(n22429) );
  NAND U27893 ( .A(n22427), .B(n22426), .Z(n22428) );
  OR U27894 ( .A(n22429), .B(n22428), .Z(n22430) );
  AND U27895 ( .A(n22431), .B(n22430), .Z(n22435) );
  NAND U27896 ( .A(n22433), .B(n22432), .Z(n22434) );
  OR U27897 ( .A(n22435), .B(n22434), .Z(n22436) );
  AND U27898 ( .A(n22437), .B(n22436), .Z(n22438) );
  NOR U27899 ( .A(n28986), .B(n22438), .Z(n22439) );
  NANDN U27900 ( .A(n22440), .B(n22439), .Z(n22441) );
  AND U27901 ( .A(n22442), .B(n22441), .Z(n22443) );
  NAND U27902 ( .A(n28987), .B(n22443), .Z(n22444) );
  NAND U27903 ( .A(n28989), .B(n22444), .Z(n22445) );
  NAND U27904 ( .A(n22446), .B(n22445), .Z(n22447) );
  NANDN U27905 ( .A(n22448), .B(n22447), .Z(n22449) );
  AND U27906 ( .A(n22450), .B(n22449), .Z(n22451) );
  NAND U27907 ( .A(n22452), .B(n22451), .Z(n22456) );
  NAND U27908 ( .A(n22454), .B(n22453), .Z(n22455) );
  ANDN U27909 ( .B(n22456), .A(n22455), .Z(n22460) );
  NAND U27910 ( .A(n22458), .B(n22457), .Z(n22459) );
  OR U27911 ( .A(n22460), .B(n22459), .Z(n22461) );
  AND U27912 ( .A(n22462), .B(n22461), .Z(n22466) );
  NAND U27913 ( .A(n22464), .B(n22463), .Z(n22465) );
  OR U27914 ( .A(n22466), .B(n22465), .Z(n22467) );
  AND U27915 ( .A(n22468), .B(n22467), .Z(n22472) );
  NAND U27916 ( .A(n22470), .B(n22469), .Z(n22471) );
  OR U27917 ( .A(n22472), .B(n22471), .Z(n22473) );
  AND U27918 ( .A(n22474), .B(n22473), .Z(n22475) );
  NOR U27919 ( .A(n22476), .B(n22475), .Z(n22477) );
  NAND U27920 ( .A(n22478), .B(n22477), .Z(n22482) );
  NAND U27921 ( .A(n22480), .B(n22479), .Z(n22481) );
  ANDN U27922 ( .B(n22482), .A(n22481), .Z(n22486) );
  NAND U27923 ( .A(n22484), .B(n22483), .Z(n22485) );
  OR U27924 ( .A(n22486), .B(n22485), .Z(n22487) );
  AND U27925 ( .A(n22488), .B(n22487), .Z(n22492) );
  NAND U27926 ( .A(n22490), .B(n22489), .Z(n22491) );
  OR U27927 ( .A(n22492), .B(n22491), .Z(n22493) );
  AND U27928 ( .A(n22494), .B(n22493), .Z(n22498) );
  NAND U27929 ( .A(n22496), .B(n22495), .Z(n22497) );
  OR U27930 ( .A(n22498), .B(n22497), .Z(n22499) );
  AND U27931 ( .A(n22500), .B(n22499), .Z(n22504) );
  NAND U27932 ( .A(n22502), .B(n22501), .Z(n22503) );
  OR U27933 ( .A(n22504), .B(n22503), .Z(n22505) );
  AND U27934 ( .A(n22506), .B(n22505), .Z(n22510) );
  NAND U27935 ( .A(n22508), .B(n22507), .Z(n22509) );
  OR U27936 ( .A(n22510), .B(n22509), .Z(n22511) );
  AND U27937 ( .A(n22512), .B(n22511), .Z(n22516) );
  NAND U27938 ( .A(n22514), .B(n22513), .Z(n22515) );
  OR U27939 ( .A(n22516), .B(n22515), .Z(n22517) );
  AND U27940 ( .A(n22518), .B(n22517), .Z(n22519) );
  NOR U27941 ( .A(n22520), .B(n22519), .Z(n22521) );
  NAND U27942 ( .A(n23965), .B(n22521), .Z(n22522) );
  NANDN U27943 ( .A(n22523), .B(n22522), .Z(n22525) );
  AND U27944 ( .A(n22525), .B(n22524), .Z(n22526) );
  NANDN U27945 ( .A(n23964), .B(n22526), .Z(n22527) );
  NAND U27946 ( .A(n22528), .B(n22527), .Z(n22529) );
  NANDN U27947 ( .A(n29015), .B(n22529), .Z(n22531) );
  OR U27948 ( .A(n22531), .B(n22530), .Z(n22532) );
  NAND U27949 ( .A(n22533), .B(n22532), .Z(n22534) );
  NANDN U27950 ( .A(n22535), .B(n22534), .Z(n22536) );
  NAND U27951 ( .A(n22537), .B(n22536), .Z(n22538) );
  ANDN U27952 ( .B(y[3606]), .A(x[3606]), .Z(n23963) );
  ANDN U27953 ( .B(n22538), .A(n23963), .Z(n22539) );
  NAND U27954 ( .A(n29022), .B(n22539), .Z(n22540) );
  AND U27955 ( .A(n22541), .B(n22540), .Z(n22542) );
  OR U27956 ( .A(n22543), .B(n22542), .Z(n22544) );
  AND U27957 ( .A(n22545), .B(n22544), .Z(n22547) );
  NAND U27958 ( .A(n22547), .B(n22546), .Z(n22548) );
  NANDN U27959 ( .A(n22549), .B(n22548), .Z(n22550) );
  AND U27960 ( .A(n22551), .B(n22550), .Z(n22552) );
  NANDN U27961 ( .A(n22553), .B(n22552), .Z(n22554) );
  NAND U27962 ( .A(n22555), .B(n22554), .Z(n22556) );
  NANDN U27963 ( .A(n22557), .B(n22556), .Z(n22558) );
  AND U27964 ( .A(n22559), .B(n22558), .Z(n22560) );
  OR U27965 ( .A(n22561), .B(n22560), .Z(n22562) );
  NAND U27966 ( .A(n22563), .B(n22562), .Z(n22564) );
  NANDN U27967 ( .A(n22565), .B(n22564), .Z(n22566) );
  NAND U27968 ( .A(n22567), .B(n22566), .Z(n22568) );
  NAND U27969 ( .A(n22569), .B(n22568), .Z(n22570) );
  NANDN U27970 ( .A(n29038), .B(n22570), .Z(n22571) );
  ANDN U27971 ( .B(y[3620]), .A(x[3620]), .Z(n23961) );
  OR U27972 ( .A(n22571), .B(n23961), .Z(n22572) );
  NAND U27973 ( .A(n22573), .B(n22572), .Z(n22574) );
  NANDN U27974 ( .A(n22575), .B(n22574), .Z(n22576) );
  ANDN U27975 ( .B(y[3622]), .A(x[3622]), .Z(n29039) );
  OR U27976 ( .A(n22576), .B(n29039), .Z(n22577) );
  NAND U27977 ( .A(n22578), .B(n22577), .Z(n22579) );
  NANDN U27978 ( .A(n22580), .B(n22579), .Z(n22582) );
  OR U27979 ( .A(n22582), .B(n22581), .Z(n22583) );
  NANDN U27980 ( .A(n22584), .B(n22583), .Z(n22585) );
  AND U27981 ( .A(n22586), .B(n22585), .Z(n22587) );
  OR U27982 ( .A(n22588), .B(n22587), .Z(n22589) );
  NAND U27983 ( .A(n22590), .B(n22589), .Z(n22591) );
  NAND U27984 ( .A(n22592), .B(n22591), .Z(n22593) );
  NANDN U27985 ( .A(n22594), .B(n22593), .Z(n22595) );
  AND U27986 ( .A(n22596), .B(n22595), .Z(n22598) );
  NAND U27987 ( .A(n22598), .B(n22597), .Z(n22599) );
  NANDN U27988 ( .A(n22600), .B(n22599), .Z(n22601) );
  AND U27989 ( .A(n22602), .B(n22601), .Z(n22603) );
  NANDN U27990 ( .A(n22604), .B(n22603), .Z(n22605) );
  NAND U27991 ( .A(n22606), .B(n22605), .Z(n22607) );
  NANDN U27992 ( .A(n22608), .B(n22607), .Z(n22609) );
  AND U27993 ( .A(n22610), .B(n22609), .Z(n22611) );
  NAND U27994 ( .A(n22612), .B(n22611), .Z(n22616) );
  NAND U27995 ( .A(n22614), .B(n22613), .Z(n22615) );
  ANDN U27996 ( .B(n22616), .A(n22615), .Z(n22620) );
  NAND U27997 ( .A(n22618), .B(n22617), .Z(n22619) );
  OR U27998 ( .A(n22620), .B(n22619), .Z(n22621) );
  AND U27999 ( .A(n22622), .B(n22621), .Z(n22626) );
  NAND U28000 ( .A(n22624), .B(n22623), .Z(n22625) );
  OR U28001 ( .A(n22626), .B(n22625), .Z(n22627) );
  AND U28002 ( .A(n22628), .B(n22627), .Z(n22632) );
  NAND U28003 ( .A(n22630), .B(n22629), .Z(n22631) );
  OR U28004 ( .A(n22632), .B(n22631), .Z(n22633) );
  AND U28005 ( .A(n22634), .B(n22633), .Z(n22638) );
  NAND U28006 ( .A(n22636), .B(n22635), .Z(n22637) );
  OR U28007 ( .A(n22638), .B(n22637), .Z(n22639) );
  AND U28008 ( .A(n22640), .B(n22639), .Z(n22644) );
  NAND U28009 ( .A(n22642), .B(n22641), .Z(n22643) );
  OR U28010 ( .A(n22644), .B(n22643), .Z(n22645) );
  AND U28011 ( .A(n22646), .B(n22645), .Z(n22647) );
  OR U28012 ( .A(n22648), .B(n22647), .Z(n22649) );
  NAND U28013 ( .A(n22650), .B(n22649), .Z(n22651) );
  AND U28014 ( .A(n22652), .B(n22651), .Z(n22653) );
  NOR U28015 ( .A(n22654), .B(n22653), .Z(n22656) );
  NAND U28016 ( .A(n22656), .B(n22655), .Z(n22658) );
  AND U28017 ( .A(n22658), .B(n22657), .Z(n22659) );
  NANDN U28018 ( .A(x[3652]), .B(y[3652]), .Z(n23956) );
  NAND U28019 ( .A(n22659), .B(n23956), .Z(n22660) );
  NANDN U28020 ( .A(n22661), .B(n22660), .Z(n22662) );
  AND U28021 ( .A(n22663), .B(n22662), .Z(n22665) );
  NAND U28022 ( .A(n22665), .B(n22664), .Z(n22666) );
  NANDN U28023 ( .A(n22667), .B(n22666), .Z(n22668) );
  AND U28024 ( .A(n22669), .B(n22668), .Z(n22671) );
  NAND U28025 ( .A(n22671), .B(n22670), .Z(n22672) );
  NANDN U28026 ( .A(n22673), .B(n22672), .Z(n22674) );
  AND U28027 ( .A(n22675), .B(n22674), .Z(n22677) );
  NAND U28028 ( .A(n22677), .B(n22676), .Z(n22678) );
  NANDN U28029 ( .A(n22679), .B(n22678), .Z(n22680) );
  AND U28030 ( .A(n22681), .B(n22680), .Z(n22683) );
  NAND U28031 ( .A(n22683), .B(n22682), .Z(n22684) );
  NANDN U28032 ( .A(n22685), .B(n22684), .Z(n22686) );
  AND U28033 ( .A(n22687), .B(n22686), .Z(n22688) );
  OR U28034 ( .A(n22689), .B(n22688), .Z(n22690) );
  NAND U28035 ( .A(n22691), .B(n22690), .Z(n22692) );
  NANDN U28036 ( .A(n22693), .B(n22692), .Z(n22694) );
  OR U28037 ( .A(n22695), .B(n22694), .Z(n22696) );
  NAND U28038 ( .A(n22697), .B(n22696), .Z(n22698) );
  NANDN U28039 ( .A(n22699), .B(n22698), .Z(n22701) );
  IV U28040 ( .A(n22700), .Z(n23949) );
  AND U28041 ( .A(n22701), .B(n23949), .Z(n22702) );
  NANDN U28042 ( .A(n29087), .B(n22702), .Z(n22703) );
  NAND U28043 ( .A(n22704), .B(n22703), .Z(n22705) );
  NANDN U28044 ( .A(n22706), .B(n22705), .Z(n22707) );
  NANDN U28045 ( .A(x[3670]), .B(y[3670]), .Z(n23950) );
  NANDN U28046 ( .A(n22707), .B(n23950), .Z(n22708) );
  NAND U28047 ( .A(n22709), .B(n22708), .Z(n22710) );
  NANDN U28048 ( .A(n29093), .B(n22710), .Z(n22711) );
  OR U28049 ( .A(n22712), .B(n22711), .Z(n22713) );
  AND U28050 ( .A(n22714), .B(n22713), .Z(n22716) );
  NAND U28051 ( .A(n22716), .B(n22715), .Z(n22717) );
  ANDN U28052 ( .B(y[3674]), .A(x[3674]), .Z(n29094) );
  ANDN U28053 ( .B(n22717), .A(n29094), .Z(n22718) );
  NANDN U28054 ( .A(n22719), .B(n22718), .Z(n22720) );
  NAND U28055 ( .A(n22721), .B(n22720), .Z(n22722) );
  NANDN U28056 ( .A(n22723), .B(n22722), .Z(n22724) );
  AND U28057 ( .A(n22725), .B(n22724), .Z(n22727) );
  NAND U28058 ( .A(n22727), .B(n22726), .Z(n22728) );
  NANDN U28059 ( .A(n22729), .B(n22728), .Z(n22730) );
  AND U28060 ( .A(n22731), .B(n22730), .Z(n22733) );
  NAND U28061 ( .A(n22733), .B(n22732), .Z(n22734) );
  NANDN U28062 ( .A(n22735), .B(n22734), .Z(n22736) );
  AND U28063 ( .A(n22737), .B(n22736), .Z(n22739) );
  NAND U28064 ( .A(n22739), .B(n22738), .Z(n22740) );
  AND U28065 ( .A(n22740), .B(n29103), .Z(n22741) );
  NANDN U28066 ( .A(x[3682]), .B(y[3682]), .Z(n23948) );
  AND U28067 ( .A(n22741), .B(n23948), .Z(n22745) );
  AND U28068 ( .A(n22743), .B(n22742), .Z(n22744) );
  NANDN U28069 ( .A(n22745), .B(n22744), .Z(n22748) );
  NANDN U28070 ( .A(x[3684]), .B(y[3684]), .Z(n29104) );
  AND U28071 ( .A(n22746), .B(n29104), .Z(n22747) );
  NAND U28072 ( .A(n22748), .B(n22747), .Z(n22749) );
  NANDN U28073 ( .A(n22750), .B(n22749), .Z(n22751) );
  NAND U28074 ( .A(n22752), .B(n22751), .Z(n22753) );
  NANDN U28075 ( .A(n22754), .B(n22753), .Z(n22755) );
  AND U28076 ( .A(n22756), .B(n22755), .Z(n22758) );
  NAND U28077 ( .A(n22758), .B(n22757), .Z(n22759) );
  NANDN U28078 ( .A(n22760), .B(n22759), .Z(n22761) );
  NAND U28079 ( .A(n22762), .B(n22761), .Z(n22764) );
  OR U28080 ( .A(n22764), .B(n22763), .Z(n22765) );
  NAND U28081 ( .A(n22766), .B(n22765), .Z(n22767) );
  NANDN U28082 ( .A(n22768), .B(n22767), .Z(n22770) );
  OR U28083 ( .A(n22770), .B(n22769), .Z(n22771) );
  NANDN U28084 ( .A(n22772), .B(n22771), .Z(n22773) );
  AND U28085 ( .A(n22774), .B(n22773), .Z(n22778) );
  NAND U28086 ( .A(n22776), .B(n22775), .Z(n22777) );
  OR U28087 ( .A(n22778), .B(n22777), .Z(n22779) );
  AND U28088 ( .A(n22780), .B(n22779), .Z(n22784) );
  NAND U28089 ( .A(n22782), .B(n22781), .Z(n22783) );
  OR U28090 ( .A(n22784), .B(n22783), .Z(n22785) );
  AND U28091 ( .A(n22786), .B(n22785), .Z(n22790) );
  NAND U28092 ( .A(n22788), .B(n22787), .Z(n22789) );
  OR U28093 ( .A(n22790), .B(n22789), .Z(n22791) );
  AND U28094 ( .A(n22792), .B(n22791), .Z(n22796) );
  NAND U28095 ( .A(n22794), .B(n22793), .Z(n22795) );
  OR U28096 ( .A(n22796), .B(n22795), .Z(n22797) );
  AND U28097 ( .A(n22798), .B(n22797), .Z(n22802) );
  NAND U28098 ( .A(n22800), .B(n22799), .Z(n22801) );
  OR U28099 ( .A(n22802), .B(n22801), .Z(n22803) );
  AND U28100 ( .A(n22804), .B(n22803), .Z(n22808) );
  NAND U28101 ( .A(n22806), .B(n22805), .Z(n22807) );
  OR U28102 ( .A(n22808), .B(n22807), .Z(n22809) );
  AND U28103 ( .A(n22810), .B(n22809), .Z(n22814) );
  NAND U28104 ( .A(n22812), .B(n22811), .Z(n22813) );
  OR U28105 ( .A(n22814), .B(n22813), .Z(n22815) );
  AND U28106 ( .A(n22816), .B(n22815), .Z(n22820) );
  NAND U28107 ( .A(n22818), .B(n22817), .Z(n22819) );
  OR U28108 ( .A(n22820), .B(n22819), .Z(n22821) );
  AND U28109 ( .A(n22822), .B(n22821), .Z(n22826) );
  NAND U28110 ( .A(n22824), .B(n22823), .Z(n22825) );
  OR U28111 ( .A(n22826), .B(n22825), .Z(n22827) );
  AND U28112 ( .A(n22828), .B(n22827), .Z(n22829) );
  NOR U28113 ( .A(n22830), .B(n22829), .Z(n22831) );
  NAND U28114 ( .A(n22832), .B(n22831), .Z(n22833) );
  NANDN U28115 ( .A(n22834), .B(n22833), .Z(n22835) );
  NAND U28116 ( .A(n22836), .B(n22835), .Z(n22837) );
  NANDN U28117 ( .A(n22838), .B(n22837), .Z(n22839) );
  AND U28118 ( .A(n22840), .B(n22839), .Z(n22842) );
  NAND U28119 ( .A(n22842), .B(n22841), .Z(n22843) );
  NANDN U28120 ( .A(n22844), .B(n22843), .Z(n22845) );
  AND U28121 ( .A(n22846), .B(n22845), .Z(n22848) );
  NAND U28122 ( .A(n22848), .B(n22847), .Z(n22849) );
  NANDN U28123 ( .A(n22850), .B(n22849), .Z(n22851) );
  AND U28124 ( .A(n22852), .B(n22851), .Z(n22853) );
  OR U28125 ( .A(n22854), .B(n22853), .Z(n22855) );
  NAND U28126 ( .A(n22856), .B(n22855), .Z(n22857) );
  AND U28127 ( .A(n22858), .B(n22857), .Z(n22862) );
  AND U28128 ( .A(n22860), .B(n22859), .Z(n22861) );
  NANDN U28129 ( .A(n22862), .B(n22861), .Z(n22865) );
  NANDN U28130 ( .A(x[3726]), .B(y[3726]), .Z(n29148) );
  AND U28131 ( .A(n22863), .B(n29148), .Z(n22864) );
  NAND U28132 ( .A(n22865), .B(n22864), .Z(n22866) );
  NANDN U28133 ( .A(n22867), .B(n22866), .Z(n22868) );
  NAND U28134 ( .A(n22869), .B(n22868), .Z(n22870) );
  NANDN U28135 ( .A(n22871), .B(n22870), .Z(n22872) );
  AND U28136 ( .A(n22873), .B(n22872), .Z(n22875) );
  NAND U28137 ( .A(n22875), .B(n22874), .Z(n22876) );
  NANDN U28138 ( .A(n22877), .B(n22876), .Z(n22878) );
  AND U28139 ( .A(n22879), .B(n22878), .Z(n22881) );
  NAND U28140 ( .A(n22881), .B(n22880), .Z(n22882) );
  NANDN U28141 ( .A(n22883), .B(n22882), .Z(n22884) );
  AND U28142 ( .A(n22885), .B(n22884), .Z(n22887) );
  NAND U28143 ( .A(n22887), .B(n22886), .Z(n22888) );
  NANDN U28144 ( .A(n22889), .B(n22888), .Z(n22890) );
  AND U28145 ( .A(n22891), .B(n22890), .Z(n22893) );
  AND U28146 ( .A(n22893), .B(n22892), .Z(n22897) );
  NAND U28147 ( .A(n22895), .B(n22894), .Z(n22896) );
  OR U28148 ( .A(n22897), .B(n22896), .Z(n22898) );
  AND U28149 ( .A(n22899), .B(n22898), .Z(n22903) );
  NAND U28150 ( .A(n22901), .B(n22900), .Z(n22902) );
  OR U28151 ( .A(n22903), .B(n22902), .Z(n22904) );
  AND U28152 ( .A(n22905), .B(n22904), .Z(n22909) );
  NAND U28153 ( .A(n22907), .B(n22906), .Z(n22908) );
  OR U28154 ( .A(n22909), .B(n22908), .Z(n22910) );
  AND U28155 ( .A(n22911), .B(n22910), .Z(n22912) );
  OR U28156 ( .A(n22913), .B(n22912), .Z(n22914) );
  NAND U28157 ( .A(n22915), .B(n22914), .Z(n22916) );
  AND U28158 ( .A(n22917), .B(n22916), .Z(n22918) );
  NOR U28159 ( .A(n29168), .B(n22918), .Z(n22919) );
  NANDN U28160 ( .A(n22920), .B(n22919), .Z(n22921) );
  AND U28161 ( .A(n22922), .B(n22921), .Z(n22924) );
  NAND U28162 ( .A(n22924), .B(n22923), .Z(n22925) );
  NANDN U28163 ( .A(n22926), .B(n22925), .Z(n22927) );
  AND U28164 ( .A(n22928), .B(n22927), .Z(n22930) );
  NAND U28165 ( .A(n22930), .B(n22929), .Z(n22931) );
  NANDN U28166 ( .A(n22932), .B(n22931), .Z(n22933) );
  AND U28167 ( .A(n22934), .B(n22933), .Z(n22936) );
  AND U28168 ( .A(n22936), .B(n22935), .Z(n22940) );
  NAND U28169 ( .A(n22938), .B(n22937), .Z(n22939) );
  OR U28170 ( .A(n22940), .B(n22939), .Z(n22941) );
  AND U28171 ( .A(n22942), .B(n22941), .Z(n22946) );
  NAND U28172 ( .A(n22944), .B(n22943), .Z(n22945) );
  OR U28173 ( .A(n22946), .B(n22945), .Z(n22947) );
  AND U28174 ( .A(n22948), .B(n22947), .Z(n22952) );
  NAND U28175 ( .A(n22950), .B(n22949), .Z(n22951) );
  OR U28176 ( .A(n22952), .B(n22951), .Z(n22953) );
  AND U28177 ( .A(n22954), .B(n22953), .Z(n22958) );
  NAND U28178 ( .A(n22956), .B(n22955), .Z(n22957) );
  OR U28179 ( .A(n22958), .B(n22957), .Z(n22959) );
  AND U28180 ( .A(n22960), .B(n22959), .Z(n22964) );
  NAND U28181 ( .A(n22962), .B(n22961), .Z(n22963) );
  OR U28182 ( .A(n22964), .B(n22963), .Z(n22965) );
  AND U28183 ( .A(n22966), .B(n22965), .Z(n22970) );
  NAND U28184 ( .A(n22968), .B(n22967), .Z(n22969) );
  OR U28185 ( .A(n22970), .B(n22969), .Z(n22971) );
  AND U28186 ( .A(n22972), .B(n22971), .Z(n22976) );
  NAND U28187 ( .A(n22974), .B(n22973), .Z(n22975) );
  OR U28188 ( .A(n22976), .B(n22975), .Z(n22977) );
  AND U28189 ( .A(n22978), .B(n22977), .Z(n22979) );
  OR U28190 ( .A(n22980), .B(n22979), .Z(n22981) );
  NAND U28191 ( .A(n22982), .B(n22981), .Z(n22985) );
  NANDN U28192 ( .A(x[3768]), .B(y[3768]), .Z(n29189) );
  AND U28193 ( .A(n22983), .B(n29189), .Z(n22984) );
  NAND U28194 ( .A(n22985), .B(n22984), .Z(n22986) );
  NANDN U28195 ( .A(n22987), .B(n22986), .Z(n22988) );
  NAND U28196 ( .A(n22989), .B(n22988), .Z(n22990) );
  NANDN U28197 ( .A(n22991), .B(n22990), .Z(n22992) );
  AND U28198 ( .A(n22993), .B(n22992), .Z(n22995) );
  NAND U28199 ( .A(n22995), .B(n22994), .Z(n22996) );
  NANDN U28200 ( .A(n22997), .B(n22996), .Z(n22998) );
  AND U28201 ( .A(n22999), .B(n22998), .Z(n23001) );
  NAND U28202 ( .A(n23001), .B(n23000), .Z(n23002) );
  NANDN U28203 ( .A(n23003), .B(n23002), .Z(n23004) );
  AND U28204 ( .A(n23005), .B(n23004), .Z(n23007) );
  AND U28205 ( .A(n23007), .B(n23006), .Z(n23011) );
  NAND U28206 ( .A(n23009), .B(n23008), .Z(n23010) );
  OR U28207 ( .A(n23011), .B(n23010), .Z(n23012) );
  AND U28208 ( .A(n23013), .B(n23012), .Z(n23017) );
  NAND U28209 ( .A(n23015), .B(n23014), .Z(n23016) );
  OR U28210 ( .A(n23017), .B(n23016), .Z(n23018) );
  AND U28211 ( .A(n23019), .B(n23018), .Z(n23023) );
  NAND U28212 ( .A(n23021), .B(n23020), .Z(n23022) );
  OR U28213 ( .A(n23023), .B(n23022), .Z(n23024) );
  AND U28214 ( .A(n23025), .B(n23024), .Z(n23026) );
  ANDN U28215 ( .B(n23027), .A(n23026), .Z(n23028) );
  NAND U28216 ( .A(n23029), .B(n23028), .Z(n23030) );
  NANDN U28217 ( .A(n23031), .B(n23030), .Z(n23032) );
  OR U28218 ( .A(n23033), .B(n23032), .Z(n23034) );
  AND U28219 ( .A(n23035), .B(n23034), .Z(n23037) );
  NAND U28220 ( .A(n23037), .B(n23036), .Z(n23038) );
  NANDN U28221 ( .A(n23039), .B(n23038), .Z(n23040) );
  AND U28222 ( .A(n23041), .B(n23040), .Z(n23043) );
  NAND U28223 ( .A(n23043), .B(n23042), .Z(n23044) );
  NANDN U28224 ( .A(n23045), .B(n23044), .Z(n23046) );
  AND U28225 ( .A(n23047), .B(n23046), .Z(n23049) );
  AND U28226 ( .A(n23049), .B(n23048), .Z(n23050) );
  OR U28227 ( .A(n23051), .B(n23050), .Z(n23052) );
  NAND U28228 ( .A(n23053), .B(n23052), .Z(n23054) );
  NANDN U28229 ( .A(n29217), .B(n23054), .Z(n23055) );
  ANDN U28230 ( .B(y[3792]), .A(x[3792]), .Z(n29213) );
  OR U28231 ( .A(n23055), .B(n29213), .Z(n23056) );
  NAND U28232 ( .A(n23057), .B(n23056), .Z(n23058) );
  NANDN U28233 ( .A(n23059), .B(n23058), .Z(n23060) );
  ANDN U28234 ( .B(y[3794]), .A(x[3794]), .Z(n23924) );
  OR U28235 ( .A(n23060), .B(n23924), .Z(n23061) );
  NAND U28236 ( .A(n23062), .B(n23061), .Z(n23063) );
  NANDN U28237 ( .A(n23064), .B(n23063), .Z(n23066) );
  OR U28238 ( .A(n23066), .B(n23065), .Z(n23067) );
  NAND U28239 ( .A(n23068), .B(n23067), .Z(n23072) );
  NAND U28240 ( .A(n23070), .B(n23069), .Z(n23071) );
  ANDN U28241 ( .B(n23072), .A(n23071), .Z(n23076) );
  NAND U28242 ( .A(n23074), .B(n23073), .Z(n23075) );
  OR U28243 ( .A(n23076), .B(n23075), .Z(n23077) );
  AND U28244 ( .A(n23078), .B(n23077), .Z(n23082) );
  NAND U28245 ( .A(n23080), .B(n23079), .Z(n23081) );
  OR U28246 ( .A(n23082), .B(n23081), .Z(n23083) );
  AND U28247 ( .A(n23084), .B(n23083), .Z(n23088) );
  NAND U28248 ( .A(n23086), .B(n23085), .Z(n23087) );
  OR U28249 ( .A(n23088), .B(n23087), .Z(n23089) );
  AND U28250 ( .A(n23090), .B(n23089), .Z(n23091) );
  OR U28251 ( .A(n23092), .B(n23091), .Z(n23093) );
  NAND U28252 ( .A(n23094), .B(n23093), .Z(n23095) );
  AND U28253 ( .A(n23096), .B(n23095), .Z(n23097) );
  ANDN U28254 ( .B(n23923), .A(n23097), .Z(n23098) );
  NANDN U28255 ( .A(n29235), .B(n23098), .Z(n23099) );
  AND U28256 ( .A(n23100), .B(n23099), .Z(n23102) );
  NAND U28257 ( .A(n23102), .B(n23101), .Z(n23103) );
  NANDN U28258 ( .A(n23104), .B(n23103), .Z(n23105) );
  AND U28259 ( .A(n23106), .B(n23105), .Z(n23107) );
  NANDN U28260 ( .A(n23108), .B(n23107), .Z(n23109) );
  NAND U28261 ( .A(n23110), .B(n23109), .Z(n23111) );
  NANDN U28262 ( .A(n23112), .B(n23111), .Z(n23114) );
  AND U28263 ( .A(n23114), .B(n23113), .Z(n23115) );
  NANDN U28264 ( .A(x[3814]), .B(y[3814]), .Z(n29241) );
  NAND U28265 ( .A(n23115), .B(n29241), .Z(n23116) );
  NANDN U28266 ( .A(n23117), .B(n23116), .Z(n23118) );
  AND U28267 ( .A(n29245), .B(n23118), .Z(n23120) );
  NAND U28268 ( .A(n23120), .B(n23119), .Z(n23121) );
  NANDN U28269 ( .A(n23122), .B(n23121), .Z(n23123) );
  AND U28270 ( .A(n29248), .B(n23123), .Z(n23124) );
  NANDN U28271 ( .A(x[3818]), .B(y[3818]), .Z(n29246) );
  AND U28272 ( .A(n23124), .B(n29246), .Z(n23125) );
  OR U28273 ( .A(n23126), .B(n23125), .Z(n23127) );
  AND U28274 ( .A(n23128), .B(n23127), .Z(n23132) );
  NAND U28275 ( .A(n23130), .B(n23129), .Z(n23131) );
  OR U28276 ( .A(n23132), .B(n23131), .Z(n23133) );
  AND U28277 ( .A(n23134), .B(n23133), .Z(n23138) );
  NAND U28278 ( .A(n23136), .B(n23135), .Z(n23137) );
  OR U28279 ( .A(n23138), .B(n23137), .Z(n23139) );
  AND U28280 ( .A(n23140), .B(n23139), .Z(n23141) );
  OR U28281 ( .A(n23142), .B(n23141), .Z(n23143) );
  NAND U28282 ( .A(n23144), .B(n23143), .Z(n23145) );
  AND U28283 ( .A(n23146), .B(n23145), .Z(n23147) );
  NOR U28284 ( .A(n23919), .B(n23147), .Z(n23148) );
  NANDN U28285 ( .A(n29260), .B(n23148), .Z(n23149) );
  AND U28286 ( .A(n23150), .B(n23149), .Z(n23152) );
  NAND U28287 ( .A(n23152), .B(n23151), .Z(n23153) );
  NANDN U28288 ( .A(n23154), .B(n23153), .Z(n23155) );
  AND U28289 ( .A(n23156), .B(n23155), .Z(n23157) );
  NANDN U28290 ( .A(n23158), .B(n23157), .Z(n23159) );
  NAND U28291 ( .A(n23160), .B(n23159), .Z(n23161) );
  NANDN U28292 ( .A(n23162), .B(n23161), .Z(n23163) );
  AND U28293 ( .A(n23164), .B(n23163), .Z(n23168) );
  AND U28294 ( .A(n23166), .B(n23165), .Z(n23167) );
  NANDN U28295 ( .A(n23168), .B(n23167), .Z(n23171) );
  NANDN U28296 ( .A(x[3836]), .B(y[3836]), .Z(n29267) );
  AND U28297 ( .A(n23169), .B(n29267), .Z(n23170) );
  NAND U28298 ( .A(n23171), .B(n23170), .Z(n23172) );
  NANDN U28299 ( .A(n23173), .B(n23172), .Z(n23174) );
  NAND U28300 ( .A(n23175), .B(n23174), .Z(n23176) );
  NANDN U28301 ( .A(n23177), .B(n23176), .Z(n23178) );
  AND U28302 ( .A(n23179), .B(n23178), .Z(n23181) );
  NAND U28303 ( .A(n23181), .B(n23180), .Z(n23182) );
  NANDN U28304 ( .A(n23183), .B(n23182), .Z(n23184) );
  AND U28305 ( .A(n29273), .B(n23184), .Z(n23186) );
  NAND U28306 ( .A(n23186), .B(n23185), .Z(n23187) );
  NANDN U28307 ( .A(n23188), .B(n23187), .Z(n23189) );
  AND U28308 ( .A(n23911), .B(n23189), .Z(n23190) );
  NANDN U28309 ( .A(x[3844]), .B(y[3844]), .Z(n29274) );
  AND U28310 ( .A(n23190), .B(n29274), .Z(n23194) );
  NAND U28311 ( .A(n23192), .B(n23191), .Z(n23193) );
  OR U28312 ( .A(n23194), .B(n23193), .Z(n23195) );
  AND U28313 ( .A(n23196), .B(n23195), .Z(n23197) );
  OR U28314 ( .A(n23198), .B(n23197), .Z(n23199) );
  NAND U28315 ( .A(n23200), .B(n23199), .Z(n23201) );
  AND U28316 ( .A(n23202), .B(n23201), .Z(n23203) );
  NOR U28317 ( .A(n29281), .B(n23203), .Z(n23204) );
  NANDN U28318 ( .A(n23909), .B(n23204), .Z(n23205) );
  AND U28319 ( .A(n23206), .B(n23205), .Z(n23208) );
  NAND U28320 ( .A(n23208), .B(n23207), .Z(n23209) );
  NANDN U28321 ( .A(n23210), .B(n23209), .Z(n23211) );
  AND U28322 ( .A(n23212), .B(n23211), .Z(n23214) );
  NAND U28323 ( .A(n23214), .B(n23213), .Z(n23215) );
  NANDN U28324 ( .A(n23216), .B(n23215), .Z(n23217) );
  AND U28325 ( .A(n23218), .B(n23217), .Z(n23220) );
  NAND U28326 ( .A(n23220), .B(n23219), .Z(n23221) );
  AND U28327 ( .A(n23222), .B(n23221), .Z(n23223) );
  NOR U28328 ( .A(n23224), .B(n23223), .Z(n23226) );
  NAND U28329 ( .A(n23226), .B(n23225), .Z(n23228) );
  AND U28330 ( .A(n23228), .B(n23227), .Z(n23229) );
  NANDN U28331 ( .A(x[3858]), .B(y[3858]), .Z(n23908) );
  AND U28332 ( .A(n23229), .B(n23908), .Z(n23230) );
  OR U28333 ( .A(n23231), .B(n23230), .Z(n23232) );
  NAND U28334 ( .A(n23233), .B(n23232), .Z(n23237) );
  NAND U28335 ( .A(n23235), .B(n23234), .Z(n23236) );
  ANDN U28336 ( .B(n23237), .A(n23236), .Z(n23241) );
  NAND U28337 ( .A(n23239), .B(n23238), .Z(n23240) );
  OR U28338 ( .A(n23241), .B(n23240), .Z(n23242) );
  AND U28339 ( .A(n23243), .B(n23242), .Z(n23247) );
  NAND U28340 ( .A(n23245), .B(n23244), .Z(n23246) );
  OR U28341 ( .A(n23247), .B(n23246), .Z(n23248) );
  AND U28342 ( .A(n23249), .B(n23248), .Z(n23253) );
  NAND U28343 ( .A(n23251), .B(n23250), .Z(n23252) );
  OR U28344 ( .A(n23253), .B(n23252), .Z(n23254) );
  AND U28345 ( .A(n23255), .B(n23254), .Z(n23259) );
  NAND U28346 ( .A(n23257), .B(n23256), .Z(n23258) );
  OR U28347 ( .A(n23259), .B(n23258), .Z(n23260) );
  AND U28348 ( .A(n23261), .B(n23260), .Z(n23262) );
  NOR U28349 ( .A(n23263), .B(n23262), .Z(n23264) );
  NAND U28350 ( .A(n23265), .B(n23264), .Z(n23266) );
  NANDN U28351 ( .A(n23267), .B(n23266), .Z(n23268) );
  AND U28352 ( .A(n23269), .B(n23268), .Z(n23270) );
  ANDN U28353 ( .B(n23271), .A(n23270), .Z(n23272) );
  OR U28354 ( .A(n23273), .B(n23272), .Z(n23274) );
  NAND U28355 ( .A(n23275), .B(n23274), .Z(n23276) );
  AND U28356 ( .A(n23277), .B(n23276), .Z(n23278) );
  NOR U28357 ( .A(n23279), .B(n23278), .Z(n23281) );
  NAND U28358 ( .A(n23281), .B(n23280), .Z(n23283) );
  NAND U28359 ( .A(n23283), .B(n23282), .Z(n23284) );
  ANDN U28360 ( .B(y[3878]), .A(x[3878]), .Z(n29306) );
  OR U28361 ( .A(n23284), .B(n29306), .Z(n23285) );
  NAND U28362 ( .A(n23286), .B(n23285), .Z(n23287) );
  NAND U28363 ( .A(n23288), .B(n23287), .Z(n23289) );
  NANDN U28364 ( .A(n23290), .B(n23289), .Z(n23291) );
  AND U28365 ( .A(n23904), .B(n23291), .Z(n23293) );
  NAND U28366 ( .A(n23293), .B(n23292), .Z(n23294) );
  NANDN U28367 ( .A(n23295), .B(n23294), .Z(n23296) );
  AND U28368 ( .A(n23297), .B(n23296), .Z(n23299) );
  NAND U28369 ( .A(n23299), .B(n23298), .Z(n23300) );
  NANDN U28370 ( .A(n23301), .B(n23300), .Z(n23302) );
  AND U28371 ( .A(n23303), .B(n23302), .Z(n23305) );
  NAND U28372 ( .A(n23305), .B(n23304), .Z(n23306) );
  NANDN U28373 ( .A(n23307), .B(n23306), .Z(n23308) );
  AND U28374 ( .A(n23308), .B(n29317), .Z(n23310) );
  AND U28375 ( .A(n23310), .B(n23309), .Z(n23314) );
  NAND U28376 ( .A(n23312), .B(n23311), .Z(n23313) );
  OR U28377 ( .A(n23314), .B(n23313), .Z(n23315) );
  AND U28378 ( .A(n23316), .B(n23315), .Z(n23317) );
  OR U28379 ( .A(n23318), .B(n23317), .Z(n23319) );
  NAND U28380 ( .A(n23320), .B(n23319), .Z(n23321) );
  NAND U28381 ( .A(n23322), .B(n23321), .Z(n23323) );
  NANDN U28382 ( .A(n23324), .B(n23323), .Z(n23325) );
  AND U28383 ( .A(n23326), .B(n23325), .Z(n23328) );
  NAND U28384 ( .A(n23328), .B(n23327), .Z(n23329) );
  NANDN U28385 ( .A(n23330), .B(n23329), .Z(n23331) );
  AND U28386 ( .A(n23332), .B(n23331), .Z(n23334) );
  NAND U28387 ( .A(n23334), .B(n23333), .Z(n23335) );
  NANDN U28388 ( .A(n23336), .B(n23335), .Z(n23337) );
  ANDN U28389 ( .B(y[3898]), .A(x[3898]), .Z(n23898) );
  OR U28390 ( .A(n23337), .B(n23898), .Z(n23338) );
  AND U28391 ( .A(n23339), .B(n23338), .Z(n23343) );
  NAND U28392 ( .A(n23341), .B(n23340), .Z(n23342) );
  OR U28393 ( .A(n23343), .B(n23342), .Z(n23344) );
  AND U28394 ( .A(n23345), .B(n23344), .Z(n23349) );
  NAND U28395 ( .A(n23347), .B(n23346), .Z(n23348) );
  OR U28396 ( .A(n23349), .B(n23348), .Z(n23350) );
  AND U28397 ( .A(n23351), .B(n23350), .Z(n23355) );
  NAND U28398 ( .A(n23353), .B(n23352), .Z(n23354) );
  OR U28399 ( .A(n23355), .B(n23354), .Z(n23356) );
  AND U28400 ( .A(n23357), .B(n23356), .Z(n23361) );
  NAND U28401 ( .A(n23359), .B(n23358), .Z(n23360) );
  OR U28402 ( .A(n23361), .B(n23360), .Z(n23362) );
  AND U28403 ( .A(n23363), .B(n23362), .Z(n23364) );
  OR U28404 ( .A(n23365), .B(n23364), .Z(n23366) );
  NAND U28405 ( .A(n23367), .B(n23366), .Z(n23368) );
  NANDN U28406 ( .A(n23369), .B(n23368), .Z(n23370) );
  ANDN U28407 ( .B(y[3910]), .A(x[3910]), .Z(n29341) );
  OR U28408 ( .A(n23370), .B(n29341), .Z(n23371) );
  NAND U28409 ( .A(n23372), .B(n23371), .Z(n23373) );
  NANDN U28410 ( .A(n23374), .B(n23373), .Z(n23376) );
  OR U28411 ( .A(n23376), .B(n23375), .Z(n23377) );
  NANDN U28412 ( .A(n23378), .B(n23377), .Z(n23379) );
  AND U28413 ( .A(n23380), .B(n23379), .Z(n23384) );
  NAND U28414 ( .A(n23382), .B(n23381), .Z(n23383) );
  OR U28415 ( .A(n23384), .B(n23383), .Z(n23385) );
  AND U28416 ( .A(n23386), .B(n23385), .Z(n23390) );
  NAND U28417 ( .A(n23388), .B(n23387), .Z(n23389) );
  OR U28418 ( .A(n23390), .B(n23389), .Z(n23391) );
  AND U28419 ( .A(n23392), .B(n23391), .Z(n23396) );
  NAND U28420 ( .A(n23394), .B(n23393), .Z(n23395) );
  OR U28421 ( .A(n23396), .B(n23395), .Z(n23397) );
  AND U28422 ( .A(n23398), .B(n23397), .Z(n23399) );
  OR U28423 ( .A(n23400), .B(n23399), .Z(n23401) );
  NAND U28424 ( .A(n23402), .B(n23401), .Z(n23403) );
  AND U28425 ( .A(n23404), .B(n23403), .Z(n23405) );
  ANDN U28426 ( .B(n23406), .A(n23405), .Z(n23407) );
  OR U28427 ( .A(n23408), .B(n23407), .Z(n23409) );
  NAND U28428 ( .A(n23410), .B(n23409), .Z(n23411) );
  AND U28429 ( .A(n23412), .B(n23411), .Z(n23413) );
  NAND U28430 ( .A(n23414), .B(n23413), .Z(n23415) );
  NANDN U28431 ( .A(n23416), .B(n23415), .Z(n23417) );
  AND U28432 ( .A(n23418), .B(n23417), .Z(n23419) );
  OR U28433 ( .A(n23420), .B(n23419), .Z(n23421) );
  NAND U28434 ( .A(n23422), .B(n23421), .Z(n23426) );
  NAND U28435 ( .A(n23424), .B(n23423), .Z(n23425) );
  ANDN U28436 ( .B(n23426), .A(n23425), .Z(n23430) );
  NAND U28437 ( .A(n23428), .B(n23427), .Z(n23429) );
  OR U28438 ( .A(n23430), .B(n23429), .Z(n23431) );
  AND U28439 ( .A(n23432), .B(n23431), .Z(n23436) );
  NAND U28440 ( .A(n23434), .B(n23433), .Z(n23435) );
  OR U28441 ( .A(n23436), .B(n23435), .Z(n23437) );
  AND U28442 ( .A(n23438), .B(n23437), .Z(n23439) );
  OR U28443 ( .A(n23440), .B(n23439), .Z(n23441) );
  NAND U28444 ( .A(n23442), .B(n23441), .Z(n23443) );
  AND U28445 ( .A(n23444), .B(n23443), .Z(n23445) );
  OR U28446 ( .A(n23446), .B(n23445), .Z(n23447) );
  NAND U28447 ( .A(n23448), .B(n23447), .Z(n23452) );
  NAND U28448 ( .A(n23450), .B(n23449), .Z(n23451) );
  ANDN U28449 ( .B(n23452), .A(n23451), .Z(n23456) );
  NAND U28450 ( .A(n23454), .B(n23453), .Z(n23455) );
  OR U28451 ( .A(n23456), .B(n23455), .Z(n23457) );
  AND U28452 ( .A(n23458), .B(n23457), .Z(n23462) );
  NAND U28453 ( .A(n23460), .B(n23459), .Z(n23461) );
  OR U28454 ( .A(n23462), .B(n23461), .Z(n23463) );
  AND U28455 ( .A(n23464), .B(n23463), .Z(n23468) );
  NAND U28456 ( .A(n23466), .B(n23465), .Z(n23467) );
  OR U28457 ( .A(n23468), .B(n23467), .Z(n23469) );
  AND U28458 ( .A(n23470), .B(n23469), .Z(n23474) );
  NAND U28459 ( .A(n23472), .B(n23471), .Z(n23473) );
  OR U28460 ( .A(n23474), .B(n23473), .Z(n23475) );
  AND U28461 ( .A(n23476), .B(n23475), .Z(n23477) );
  NOR U28462 ( .A(n23478), .B(n23477), .Z(n23479) );
  NAND U28463 ( .A(n23480), .B(n23479), .Z(n23481) );
  NANDN U28464 ( .A(n23482), .B(n23481), .Z(n23483) );
  NAND U28465 ( .A(n23484), .B(n23483), .Z(n23485) );
  NANDN U28466 ( .A(n23486), .B(n23485), .Z(n23487) );
  AND U28467 ( .A(n23488), .B(n23487), .Z(n23490) );
  NAND U28468 ( .A(n23490), .B(n23489), .Z(n23491) );
  NANDN U28469 ( .A(n23492), .B(n23491), .Z(n23493) );
  AND U28470 ( .A(n23494), .B(n23493), .Z(n23496) );
  NAND U28471 ( .A(n23496), .B(n23495), .Z(n23497) );
  NANDN U28472 ( .A(n23498), .B(n23497), .Z(n23499) );
  AND U28473 ( .A(n23500), .B(n23499), .Z(n23502) );
  AND U28474 ( .A(n23502), .B(n23501), .Z(n23506) );
  NAND U28475 ( .A(n23504), .B(n23503), .Z(n23505) );
  OR U28476 ( .A(n23506), .B(n23505), .Z(n23507) );
  AND U28477 ( .A(n23508), .B(n23507), .Z(n23512) );
  NAND U28478 ( .A(n23510), .B(n23509), .Z(n23511) );
  OR U28479 ( .A(n23512), .B(n23511), .Z(n23513) );
  AND U28480 ( .A(n23514), .B(n23513), .Z(n23515) );
  OR U28481 ( .A(n23516), .B(n23515), .Z(n23517) );
  NAND U28482 ( .A(n23518), .B(n23517), .Z(n23519) );
  AND U28483 ( .A(n23520), .B(n23519), .Z(n23521) );
  NOR U28484 ( .A(n23522), .B(n23521), .Z(n23524) );
  XNOR U28485 ( .A(x[3968]), .B(y[3968]), .Z(n23523) );
  NAND U28486 ( .A(n23524), .B(n23523), .Z(n23527) );
  NANDN U28487 ( .A(x[3968]), .B(y[3968]), .Z(n29401) );
  AND U28488 ( .A(n23525), .B(n29401), .Z(n23526) );
  NAND U28489 ( .A(n23527), .B(n23526), .Z(n23528) );
  NANDN U28490 ( .A(n23529), .B(n23528), .Z(n23530) );
  NAND U28491 ( .A(n23531), .B(n23530), .Z(n23532) );
  NANDN U28492 ( .A(n23533), .B(n23532), .Z(n23534) );
  AND U28493 ( .A(n23535), .B(n23534), .Z(n23537) );
  NAND U28494 ( .A(n23537), .B(n23536), .Z(n23538) );
  NANDN U28495 ( .A(n23539), .B(n23538), .Z(n23540) );
  AND U28496 ( .A(n23541), .B(n23540), .Z(n23543) );
  NAND U28497 ( .A(n23543), .B(n23542), .Z(n23544) );
  NANDN U28498 ( .A(n23545), .B(n23544), .Z(n23546) );
  AND U28499 ( .A(n23547), .B(n23546), .Z(n23549) );
  AND U28500 ( .A(n23549), .B(n23548), .Z(n23553) );
  NAND U28501 ( .A(n23551), .B(n23550), .Z(n23552) );
  OR U28502 ( .A(n23553), .B(n23552), .Z(n23554) );
  AND U28503 ( .A(n23555), .B(n23554), .Z(n23559) );
  NAND U28504 ( .A(n23557), .B(n23556), .Z(n23558) );
  OR U28505 ( .A(n23559), .B(n23558), .Z(n23560) );
  AND U28506 ( .A(n23561), .B(n23560), .Z(n23562) );
  NOR U28507 ( .A(n23563), .B(n23562), .Z(n23564) );
  NAND U28508 ( .A(n23565), .B(n23564), .Z(n23566) );
  NANDN U28509 ( .A(n23567), .B(n23566), .Z(n23568) );
  NAND U28510 ( .A(n23569), .B(n23568), .Z(n23570) );
  NANDN U28511 ( .A(n23571), .B(n23570), .Z(n23572) );
  AND U28512 ( .A(n23573), .B(n23572), .Z(n23575) );
  NAND U28513 ( .A(n23575), .B(n23574), .Z(n23576) );
  NANDN U28514 ( .A(n23577), .B(n23576), .Z(n23578) );
  AND U28515 ( .A(n23579), .B(n23578), .Z(n23581) );
  NAND U28516 ( .A(n23581), .B(n23580), .Z(n23582) );
  NANDN U28517 ( .A(n23583), .B(n23582), .Z(n23584) );
  AND U28518 ( .A(n23585), .B(n23584), .Z(n23587) );
  NAND U28519 ( .A(n23587), .B(n23586), .Z(n23588) );
  AND U28520 ( .A(n23588), .B(n23880), .Z(n23589) );
  NANDN U28521 ( .A(n29425), .B(n23589), .Z(n23590) );
  NAND U28522 ( .A(n23591), .B(n23590), .Z(n23592) );
  NANDN U28523 ( .A(n29429), .B(n23592), .Z(n23593) );
  ANDN U28524 ( .B(y[3992]), .A(x[3992]), .Z(n23881) );
  OR U28525 ( .A(n23593), .B(n23881), .Z(n23594) );
  NAND U28526 ( .A(n23595), .B(n23594), .Z(n23596) );
  NANDN U28527 ( .A(n23597), .B(n23596), .Z(n23598) );
  ANDN U28528 ( .B(y[3994]), .A(x[3994]), .Z(n29428) );
  OR U28529 ( .A(n23598), .B(n29428), .Z(n23599) );
  NAND U28530 ( .A(n23600), .B(n23599), .Z(n23601) );
  NANDN U28531 ( .A(n23602), .B(n23601), .Z(n23604) );
  OR U28532 ( .A(n23604), .B(n23603), .Z(n23605) );
  NAND U28533 ( .A(n23606), .B(n23605), .Z(n23610) );
  NAND U28534 ( .A(n23608), .B(n23607), .Z(n23609) );
  ANDN U28535 ( .B(n23610), .A(n23609), .Z(n23614) );
  NAND U28536 ( .A(n23612), .B(n23611), .Z(n23613) );
  OR U28537 ( .A(n23614), .B(n23613), .Z(n23615) );
  AND U28538 ( .A(n23616), .B(n23615), .Z(n23620) );
  NAND U28539 ( .A(n23618), .B(n23617), .Z(n23619) );
  OR U28540 ( .A(n23620), .B(n23619), .Z(n23621) );
  AND U28541 ( .A(n23622), .B(n23621), .Z(n23626) );
  NAND U28542 ( .A(n23624), .B(n23623), .Z(n23625) );
  OR U28543 ( .A(n23626), .B(n23625), .Z(n23627) );
  AND U28544 ( .A(n23628), .B(n23627), .Z(n23632) );
  NAND U28545 ( .A(n23630), .B(n23629), .Z(n23631) );
  OR U28546 ( .A(n23632), .B(n23631), .Z(n23633) );
  AND U28547 ( .A(n23634), .B(n23633), .Z(n23638) );
  NAND U28548 ( .A(n23636), .B(n23635), .Z(n23637) );
  OR U28549 ( .A(n23638), .B(n23637), .Z(n23639) );
  AND U28550 ( .A(n23640), .B(n23639), .Z(n23644) );
  NAND U28551 ( .A(n23642), .B(n23641), .Z(n23643) );
  OR U28552 ( .A(n23644), .B(n23643), .Z(n23645) );
  AND U28553 ( .A(n23646), .B(n23645), .Z(n23647) );
  OR U28554 ( .A(n23648), .B(n23647), .Z(n23649) );
  NAND U28555 ( .A(n23650), .B(n23649), .Z(n23651) );
  AND U28556 ( .A(n23652), .B(n23651), .Z(n23653) );
  NOR U28557 ( .A(n29450), .B(n23653), .Z(n23654) );
  NANDN U28558 ( .A(n23655), .B(n23654), .Z(n23656) );
  AND U28559 ( .A(n23657), .B(n23656), .Z(n23659) );
  NAND U28560 ( .A(n23659), .B(n23658), .Z(n23660) );
  NANDN U28561 ( .A(n23661), .B(n23660), .Z(n23662) );
  AND U28562 ( .A(n23663), .B(n23662), .Z(n23665) );
  NAND U28563 ( .A(n23665), .B(n23664), .Z(n23666) );
  NANDN U28564 ( .A(n23667), .B(n23666), .Z(n23668) );
  AND U28565 ( .A(n23669), .B(n23668), .Z(n23671) );
  AND U28566 ( .A(n23671), .B(n23670), .Z(n23675) );
  NAND U28567 ( .A(n23673), .B(n23672), .Z(n23674) );
  OR U28568 ( .A(n23675), .B(n23674), .Z(n23676) );
  AND U28569 ( .A(n23677), .B(n23676), .Z(n23678) );
  OR U28570 ( .A(n23679), .B(n23678), .Z(n23680) );
  NAND U28571 ( .A(n23681), .B(n23680), .Z(n23684) );
  NANDN U28572 ( .A(x[4024]), .B(y[4024]), .Z(n29461) );
  AND U28573 ( .A(n23682), .B(n29461), .Z(n23683) );
  NAND U28574 ( .A(n23684), .B(n23683), .Z(n23685) );
  NANDN U28575 ( .A(n23686), .B(n23685), .Z(n23687) );
  NAND U28576 ( .A(n23688), .B(n23687), .Z(n23689) );
  NANDN U28577 ( .A(n23690), .B(n23689), .Z(n23691) );
  AND U28578 ( .A(n23692), .B(n23691), .Z(n23694) );
  NAND U28579 ( .A(n23694), .B(n23693), .Z(n23695) );
  NANDN U28580 ( .A(n23696), .B(n23695), .Z(n23697) );
  AND U28581 ( .A(n23698), .B(n23697), .Z(n23700) );
  NAND U28582 ( .A(n23700), .B(n23699), .Z(n23701) );
  NANDN U28583 ( .A(n23702), .B(n23701), .Z(n23703) );
  AND U28584 ( .A(n23704), .B(n23703), .Z(n23706) );
  AND U28585 ( .A(n23706), .B(n23705), .Z(n23710) );
  NAND U28586 ( .A(n23708), .B(n23707), .Z(n23709) );
  OR U28587 ( .A(n23710), .B(n23709), .Z(n23711) );
  AND U28588 ( .A(n23712), .B(n23711), .Z(n23716) );
  NAND U28589 ( .A(n23714), .B(n23713), .Z(n23715) );
  OR U28590 ( .A(n23716), .B(n23715), .Z(n23717) );
  AND U28591 ( .A(n23718), .B(n23717), .Z(n23722) );
  NAND U28592 ( .A(n23720), .B(n23719), .Z(n23721) );
  OR U28593 ( .A(n23722), .B(n23721), .Z(n23723) );
  AND U28594 ( .A(n23724), .B(n23723), .Z(n23728) );
  NAND U28595 ( .A(n23726), .B(n23725), .Z(n23727) );
  OR U28596 ( .A(n23728), .B(n23727), .Z(n23729) );
  AND U28597 ( .A(n23730), .B(n23729), .Z(n23734) );
  NAND U28598 ( .A(n23732), .B(n23731), .Z(n23733) );
  OR U28599 ( .A(n23734), .B(n23733), .Z(n23735) );
  AND U28600 ( .A(n23736), .B(n23735), .Z(n23737) );
  ANDN U28601 ( .B(n23738), .A(n23737), .Z(n23739) );
  NAND U28602 ( .A(n23740), .B(n23739), .Z(n23741) );
  NANDN U28603 ( .A(n23742), .B(n23741), .Z(n23743) );
  OR U28604 ( .A(n23744), .B(n23743), .Z(n23745) );
  AND U28605 ( .A(n23746), .B(n23745), .Z(n23748) );
  NAND U28606 ( .A(n23748), .B(n23747), .Z(n23749) );
  NANDN U28607 ( .A(n23750), .B(n23749), .Z(n23751) );
  AND U28608 ( .A(n23752), .B(n23751), .Z(n23754) );
  NAND U28609 ( .A(n23754), .B(n23753), .Z(n23755) );
  NANDN U28610 ( .A(n23756), .B(n23755), .Z(n23757) );
  AND U28611 ( .A(n23758), .B(n23757), .Z(n23760) );
  NAND U28612 ( .A(n23760), .B(n23759), .Z(n23761) );
  NANDN U28613 ( .A(n23762), .B(n23761), .Z(n23763) );
  AND U28614 ( .A(n23764), .B(n23763), .Z(n23766) );
  XNOR U28615 ( .A(x[4052]), .B(y[4052]), .Z(n23765) );
  NAND U28616 ( .A(n23766), .B(n23765), .Z(n23767) );
  NANDN U28617 ( .A(n29486), .B(n23767), .Z(n23768) );
  ANDN U28618 ( .B(y[4052]), .A(x[4052]), .Z(n29483) );
  OR U28619 ( .A(n23768), .B(n29483), .Z(n23769) );
  NAND U28620 ( .A(n23770), .B(n23769), .Z(n23771) );
  NANDN U28621 ( .A(n23772), .B(n23771), .Z(n23773) );
  ANDN U28622 ( .B(y[4054]), .A(x[4054]), .Z(n29487) );
  OR U28623 ( .A(n23773), .B(n29487), .Z(n23774) );
  NAND U28624 ( .A(n23775), .B(n23774), .Z(n23776) );
  NANDN U28625 ( .A(n23777), .B(n23776), .Z(n23778) );
  ANDN U28626 ( .B(n23861), .A(n23778), .Z(n23779) );
  OR U28627 ( .A(n23780), .B(n23779), .Z(n23781) );
  NAND U28628 ( .A(n23782), .B(n23781), .Z(n23783) );
  NAND U28629 ( .A(n23784), .B(n23783), .Z(n23785) );
  NANDN U28630 ( .A(n23786), .B(n23785), .Z(n23787) );
  AND U28631 ( .A(n23788), .B(n23787), .Z(n23790) );
  NAND U28632 ( .A(n23790), .B(n23789), .Z(n23791) );
  NANDN U28633 ( .A(n23792), .B(n23791), .Z(n23793) );
  AND U28634 ( .A(n23794), .B(n23793), .Z(n23796) );
  NAND U28635 ( .A(n23796), .B(n23795), .Z(n23797) );
  NANDN U28636 ( .A(n23798), .B(n23797), .Z(n23799) );
  AND U28637 ( .A(n23800), .B(n23799), .Z(n23801) );
  NANDN U28638 ( .A(n23802), .B(n23801), .Z(n23803) );
  NAND U28639 ( .A(n23804), .B(n23803), .Z(n23808) );
  NAND U28640 ( .A(n23806), .B(n23805), .Z(n23807) );
  ANDN U28641 ( .B(n23808), .A(n23807), .Z(n23809) );
  OR U28642 ( .A(n23810), .B(n23809), .Z(n23811) );
  NAND U28643 ( .A(n23812), .B(n23811), .Z(n23813) );
  NANDN U28644 ( .A(n29507), .B(n23813), .Z(n23814) );
  ANDN U28645 ( .B(y[4070]), .A(x[4070]), .Z(n23857) );
  OR U28646 ( .A(n23814), .B(n23857), .Z(n23815) );
  NAND U28647 ( .A(n23816), .B(n23815), .Z(n23817) );
  NANDN U28648 ( .A(n23818), .B(n23817), .Z(n23819) );
  ANDN U28649 ( .B(y[4072]), .A(x[4072]), .Z(n29506) );
  OR U28650 ( .A(n23819), .B(n29506), .Z(n23820) );
  NAND U28651 ( .A(n23821), .B(n23820), .Z(n23822) );
  NANDN U28652 ( .A(n23823), .B(n23822), .Z(n23824) );
  AND U28653 ( .A(n23825), .B(n23824), .Z(n23826) );
  NOR U28654 ( .A(n23856), .B(n23826), .Z(n23827) );
  NANDN U28655 ( .A(n29514), .B(n23827), .Z(n23828) );
  AND U28656 ( .A(n23829), .B(n23828), .Z(n23831) );
  NAND U28657 ( .A(n23831), .B(n23830), .Z(n23832) );
  NANDN U28658 ( .A(n23833), .B(n23832), .Z(n23834) );
  AND U28659 ( .A(n23835), .B(n23834), .Z(n23837) );
  NAND U28660 ( .A(n23837), .B(n23836), .Z(n23838) );
  NANDN U28661 ( .A(n23839), .B(n23838), .Z(n23840) );
  AND U28662 ( .A(n23841), .B(n23840), .Z(n23843) );
  AND U28663 ( .A(n23843), .B(n23842), .Z(n23844) );
  OR U28664 ( .A(n23845), .B(n23844), .Z(n23846) );
  NAND U28665 ( .A(n23847), .B(n23846), .Z(n23848) );
  NAND U28666 ( .A(n23849), .B(n23848), .Z(n29531) );
  NANDN U28667 ( .A(n29531), .B(e), .Z(n5) );
  IV U28668 ( .A(n23879), .Z(n29433) );
  IV U28669 ( .A(n23886), .Z(n29406) );
  IV U28670 ( .A(n23897), .Z(n29333) );
  AND U28671 ( .A(n23923), .B(n23922), .Z(n29233) );
  IV U28672 ( .A(n23929), .Z(n29185) );
  IV U28673 ( .A(n23953), .Z(n29079) );
  IV U28674 ( .A(n23969), .Z(n29007) );
  IV U28675 ( .A(n24015), .Z(n28827) );
  IV U28676 ( .A(n24020), .Z(n28818) );
  IV U28677 ( .A(n24052), .Z(n28720) );
  IV U28678 ( .A(n24062), .Z(n28685) );
  IV U28679 ( .A(n24072), .Z(n28668) );
  IV U28680 ( .A(n24079), .Z(n28642) );
  IV U28681 ( .A(n24100), .Z(n28529) );
  NANDN U28682 ( .A(n24116), .B(n24115), .Z(n24117) );
  AND U28683 ( .A(n24118), .B(n24117), .Z(n28457) );
  IV U28684 ( .A(n24127), .Z(n28413) );
  IV U28685 ( .A(n24140), .Z(n28375) );
  AND U28686 ( .A(n24163), .B(n24162), .Z(n28212) );
  NANDN U28687 ( .A(n24177), .B(n24176), .Z(n28153) );
  IV U28688 ( .A(n24188), .Z(n24190) );
  IV U28689 ( .A(n24191), .Z(n24192) );
  NANDN U28690 ( .A(n24214), .B(n24213), .Z(n24215) );
  IV U28691 ( .A(n24221), .Z(n27969) );
  IV U28692 ( .A(n24295), .Z(n27438) );
  IV U28693 ( .A(n24311), .Z(n27374) );
  IV U28694 ( .A(n24322), .Z(n27293) );
  IV U28695 ( .A(n24326), .Z(n27279) );
  IV U28696 ( .A(n24341), .Z(n27112) );
  IV U28697 ( .A(n24355), .Z(n27021) );
  IV U28698 ( .A(n24435), .Z(n26479) );
  IV U28699 ( .A(n24444), .Z(n26393) );
  IV U28700 ( .A(n24455), .Z(n26332) );
  IV U28701 ( .A(n24467), .Z(n26276) );
  IV U28702 ( .A(n24472), .Z(n26247) );
  IV U28703 ( .A(n24486), .Z(n26151) );
  IV U28704 ( .A(n24496), .Z(n26109) );
  IV U28705 ( .A(n24515), .Z(n25925) );
  OR U28706 ( .A(n24541), .B(n24540), .Z(n24542) );
  NAND U28707 ( .A(n24543), .B(n24542), .Z(n24544) );
  NANDN U28708 ( .A(n24545), .B(n24544), .Z(n24546) );
  NAND U28709 ( .A(n24547), .B(n24546), .Z(n24548) );
  NANDN U28710 ( .A(n24549), .B(n24548), .Z(n24550) );
  AND U28711 ( .A(n24551), .B(n24550), .Z(n24552) );
  OR U28712 ( .A(n24553), .B(n24552), .Z(n24554) );
  NAND U28713 ( .A(n24555), .B(n24554), .Z(n24556) );
  NANDN U28714 ( .A(n24557), .B(n24556), .Z(n24558) );
  NAND U28715 ( .A(n24559), .B(n24558), .Z(n24560) );
  NANDN U28716 ( .A(n24561), .B(n24560), .Z(n24562) );
  AND U28717 ( .A(n24563), .B(n24562), .Z(n24564) );
  OR U28718 ( .A(n24565), .B(n24564), .Z(n24566) );
  NAND U28719 ( .A(n24567), .B(n24566), .Z(n24568) );
  NANDN U28720 ( .A(n24569), .B(n24568), .Z(n24570) );
  NAND U28721 ( .A(n24571), .B(n24570), .Z(n24572) );
  NANDN U28722 ( .A(n24573), .B(n24572), .Z(n24574) );
  AND U28723 ( .A(n24575), .B(n24574), .Z(n24576) );
  OR U28724 ( .A(n24577), .B(n24576), .Z(n24578) );
  NAND U28725 ( .A(n24579), .B(n24578), .Z(n24580) );
  NANDN U28726 ( .A(n24581), .B(n24580), .Z(n24582) );
  NAND U28727 ( .A(n24583), .B(n24582), .Z(n24584) );
  NANDN U28728 ( .A(n24585), .B(n24584), .Z(n24586) );
  AND U28729 ( .A(n24587), .B(n24586), .Z(n24588) );
  OR U28730 ( .A(n24589), .B(n24588), .Z(n24590) );
  NAND U28731 ( .A(n24591), .B(n24590), .Z(n24592) );
  NANDN U28732 ( .A(n24593), .B(n24592), .Z(n24594) );
  NAND U28733 ( .A(n24595), .B(n24594), .Z(n24596) );
  NANDN U28734 ( .A(n24597), .B(n24596), .Z(n24598) );
  AND U28735 ( .A(n24599), .B(n24598), .Z(n24600) );
  OR U28736 ( .A(n24601), .B(n24600), .Z(n24602) );
  NAND U28737 ( .A(n24603), .B(n24602), .Z(n24604) );
  NANDN U28738 ( .A(n24605), .B(n24604), .Z(n24606) );
  NAND U28739 ( .A(n24607), .B(n24606), .Z(n24608) );
  NANDN U28740 ( .A(n24609), .B(n24608), .Z(n24610) );
  AND U28741 ( .A(n24611), .B(n24610), .Z(n24612) );
  OR U28742 ( .A(n24613), .B(n24612), .Z(n24614) );
  NAND U28743 ( .A(n24615), .B(n24614), .Z(n24616) );
  NANDN U28744 ( .A(n24617), .B(n24616), .Z(n24618) );
  NAND U28745 ( .A(n24619), .B(n24618), .Z(n24620) );
  NANDN U28746 ( .A(n24621), .B(n24620), .Z(n24622) );
  AND U28747 ( .A(n24623), .B(n24622), .Z(n24624) );
  OR U28748 ( .A(n24625), .B(n24624), .Z(n24626) );
  NAND U28749 ( .A(n24627), .B(n24626), .Z(n24628) );
  NANDN U28750 ( .A(n24629), .B(n24628), .Z(n24630) );
  NAND U28751 ( .A(n24631), .B(n24630), .Z(n24632) );
  NANDN U28752 ( .A(n24633), .B(n24632), .Z(n24634) );
  AND U28753 ( .A(n24635), .B(n24634), .Z(n24636) );
  OR U28754 ( .A(n24637), .B(n24636), .Z(n24638) );
  NAND U28755 ( .A(n24639), .B(n24638), .Z(n24640) );
  NANDN U28756 ( .A(n24641), .B(n24640), .Z(n24642) );
  NAND U28757 ( .A(n24643), .B(n24642), .Z(n24644) );
  NANDN U28758 ( .A(n24645), .B(n24644), .Z(n24646) );
  AND U28759 ( .A(n24647), .B(n24646), .Z(n24648) );
  OR U28760 ( .A(n24649), .B(n24648), .Z(n24650) );
  NAND U28761 ( .A(n24651), .B(n24650), .Z(n24652) );
  NANDN U28762 ( .A(n24653), .B(n24652), .Z(n24654) );
  NAND U28763 ( .A(n24655), .B(n24654), .Z(n24656) );
  NANDN U28764 ( .A(n24657), .B(n24656), .Z(n24658) );
  AND U28765 ( .A(n24659), .B(n24658), .Z(n24660) );
  OR U28766 ( .A(n24661), .B(n24660), .Z(n24662) );
  NAND U28767 ( .A(n24663), .B(n24662), .Z(n24664) );
  NANDN U28768 ( .A(n24665), .B(n24664), .Z(n24666) );
  NAND U28769 ( .A(n24667), .B(n24666), .Z(n24668) );
  NANDN U28770 ( .A(n24669), .B(n24668), .Z(n24670) );
  AND U28771 ( .A(n24671), .B(n24670), .Z(n24673) );
  NANDN U28772 ( .A(n24673), .B(n24672), .Z(n24674) );
  NAND U28773 ( .A(n24675), .B(n24674), .Z(n24676) );
  NANDN U28774 ( .A(n24677), .B(n24676), .Z(n24678) );
  NAND U28775 ( .A(n24679), .B(n24678), .Z(n24680) );
  NANDN U28776 ( .A(n24681), .B(n24680), .Z(n24682) );
  AND U28777 ( .A(n24683), .B(n24682), .Z(n24684) );
  OR U28778 ( .A(n24685), .B(n24684), .Z(n24686) );
  NAND U28779 ( .A(n24687), .B(n24686), .Z(n24688) );
  NANDN U28780 ( .A(n24689), .B(n24688), .Z(n24690) );
  NAND U28781 ( .A(n24691), .B(n24690), .Z(n24692) );
  NANDN U28782 ( .A(n24693), .B(n24692), .Z(n24694) );
  AND U28783 ( .A(n24695), .B(n24694), .Z(n24696) );
  OR U28784 ( .A(n24697), .B(n24696), .Z(n24698) );
  NAND U28785 ( .A(n24699), .B(n24698), .Z(n24700) );
  NANDN U28786 ( .A(n24701), .B(n24700), .Z(n24702) );
  NAND U28787 ( .A(n24703), .B(n24702), .Z(n24704) );
  NANDN U28788 ( .A(n24705), .B(n24704), .Z(n24706) );
  AND U28789 ( .A(n24707), .B(n24706), .Z(n24708) );
  OR U28790 ( .A(n24709), .B(n24708), .Z(n24710) );
  NAND U28791 ( .A(n24711), .B(n24710), .Z(n24712) );
  NANDN U28792 ( .A(n24713), .B(n24712), .Z(n24714) );
  NAND U28793 ( .A(n24715), .B(n24714), .Z(n24716) );
  NANDN U28794 ( .A(n24717), .B(n24716), .Z(n24718) );
  AND U28795 ( .A(n24719), .B(n24718), .Z(n24720) );
  OR U28796 ( .A(n24721), .B(n24720), .Z(n24722) );
  NAND U28797 ( .A(n24723), .B(n24722), .Z(n24724) );
  NANDN U28798 ( .A(n24725), .B(n24724), .Z(n24726) );
  NAND U28799 ( .A(n24727), .B(n24726), .Z(n24728) );
  NANDN U28800 ( .A(n24729), .B(n24728), .Z(n24730) );
  AND U28801 ( .A(n24731), .B(n24730), .Z(n24732) );
  OR U28802 ( .A(n24733), .B(n24732), .Z(n24734) );
  NAND U28803 ( .A(n24735), .B(n24734), .Z(n24736) );
  NANDN U28804 ( .A(n24737), .B(n24736), .Z(n24738) );
  NAND U28805 ( .A(n24739), .B(n24738), .Z(n24740) );
  NANDN U28806 ( .A(n24741), .B(n24740), .Z(n24742) );
  AND U28807 ( .A(n24743), .B(n24742), .Z(n24744) );
  OR U28808 ( .A(n24745), .B(n24744), .Z(n24746) );
  NAND U28809 ( .A(n24747), .B(n24746), .Z(n24748) );
  NANDN U28810 ( .A(n24749), .B(n24748), .Z(n24750) );
  NAND U28811 ( .A(n24751), .B(n24750), .Z(n24752) );
  NANDN U28812 ( .A(n24753), .B(n24752), .Z(n24754) );
  AND U28813 ( .A(n24755), .B(n24754), .Z(n24756) );
  OR U28814 ( .A(n24757), .B(n24756), .Z(n24758) );
  NAND U28815 ( .A(n24759), .B(n24758), .Z(n24760) );
  NANDN U28816 ( .A(n24761), .B(n24760), .Z(n24762) );
  NAND U28817 ( .A(n24763), .B(n24762), .Z(n24764) );
  NANDN U28818 ( .A(n24765), .B(n24764), .Z(n24766) );
  AND U28819 ( .A(n24767), .B(n24766), .Z(n24768) );
  OR U28820 ( .A(n24769), .B(n24768), .Z(n24770) );
  NAND U28821 ( .A(n24771), .B(n24770), .Z(n24772) );
  NANDN U28822 ( .A(n24773), .B(n24772), .Z(n24774) );
  NAND U28823 ( .A(n24775), .B(n24774), .Z(n24776) );
  NANDN U28824 ( .A(n24777), .B(n24776), .Z(n24778) );
  AND U28825 ( .A(n24779), .B(n24778), .Z(n24780) );
  OR U28826 ( .A(n24781), .B(n24780), .Z(n24782) );
  NAND U28827 ( .A(n24783), .B(n24782), .Z(n24784) );
  NANDN U28828 ( .A(n24785), .B(n24784), .Z(n24786) );
  NAND U28829 ( .A(n24787), .B(n24786), .Z(n24788) );
  NANDN U28830 ( .A(n24789), .B(n24788), .Z(n24790) );
  AND U28831 ( .A(n24791), .B(n24790), .Z(n24792) );
  OR U28832 ( .A(n24793), .B(n24792), .Z(n24794) );
  NAND U28833 ( .A(n24795), .B(n24794), .Z(n24796) );
  NANDN U28834 ( .A(n24797), .B(n24796), .Z(n24798) );
  NAND U28835 ( .A(n24799), .B(n24798), .Z(n24800) );
  NANDN U28836 ( .A(n24801), .B(n24800), .Z(n24802) );
  AND U28837 ( .A(n24803), .B(n24802), .Z(n24804) );
  OR U28838 ( .A(n24805), .B(n24804), .Z(n24806) );
  NAND U28839 ( .A(n24807), .B(n24806), .Z(n24808) );
  NANDN U28840 ( .A(n24809), .B(n24808), .Z(n24810) );
  NAND U28841 ( .A(n24811), .B(n24810), .Z(n24812) );
  NANDN U28842 ( .A(n24813), .B(n24812), .Z(n24814) );
  AND U28843 ( .A(n24815), .B(n24814), .Z(n24817) );
  NANDN U28844 ( .A(n24817), .B(n24816), .Z(n24818) );
  NAND U28845 ( .A(n24819), .B(n24818), .Z(n24820) );
  NANDN U28846 ( .A(n24821), .B(n24820), .Z(n24822) );
  NAND U28847 ( .A(n24823), .B(n24822), .Z(n24824) );
  NANDN U28848 ( .A(n24825), .B(n24824), .Z(n24826) );
  AND U28849 ( .A(n24827), .B(n24826), .Z(n24828) );
  OR U28850 ( .A(n24829), .B(n24828), .Z(n24830) );
  NAND U28851 ( .A(n24831), .B(n24830), .Z(n24832) );
  NANDN U28852 ( .A(n24833), .B(n24832), .Z(n24834) );
  NAND U28853 ( .A(n24835), .B(n24834), .Z(n24836) );
  NANDN U28854 ( .A(n24837), .B(n24836), .Z(n24838) );
  AND U28855 ( .A(n24839), .B(n24838), .Z(n24840) );
  OR U28856 ( .A(n24841), .B(n24840), .Z(n24842) );
  NAND U28857 ( .A(n24843), .B(n24842), .Z(n24844) );
  NANDN U28858 ( .A(n24845), .B(n24844), .Z(n24846) );
  NAND U28859 ( .A(n24847), .B(n24846), .Z(n24848) );
  NANDN U28860 ( .A(n24849), .B(n24848), .Z(n24850) );
  AND U28861 ( .A(n24851), .B(n24850), .Z(n24852) );
  OR U28862 ( .A(n24853), .B(n24852), .Z(n24854) );
  NAND U28863 ( .A(n24855), .B(n24854), .Z(n24856) );
  NANDN U28864 ( .A(n24857), .B(n24856), .Z(n24858) );
  NAND U28865 ( .A(n24859), .B(n24858), .Z(n24860) );
  NANDN U28866 ( .A(n24861), .B(n24860), .Z(n24862) );
  AND U28867 ( .A(n24863), .B(n24862), .Z(n24864) );
  OR U28868 ( .A(n24865), .B(n24864), .Z(n24866) );
  NAND U28869 ( .A(n24867), .B(n24866), .Z(n24868) );
  NANDN U28870 ( .A(n24869), .B(n24868), .Z(n24870) );
  NAND U28871 ( .A(n24871), .B(n24870), .Z(n24872) );
  NANDN U28872 ( .A(n24873), .B(n24872), .Z(n24874) );
  AND U28873 ( .A(n24875), .B(n24874), .Z(n24876) );
  OR U28874 ( .A(n24877), .B(n24876), .Z(n24878) );
  NAND U28875 ( .A(n24879), .B(n24878), .Z(n24880) );
  NANDN U28876 ( .A(n24881), .B(n24880), .Z(n24882) );
  NAND U28877 ( .A(n24883), .B(n24882), .Z(n24884) );
  NANDN U28878 ( .A(n24885), .B(n24884), .Z(n24886) );
  AND U28879 ( .A(n24887), .B(n24886), .Z(n24888) );
  OR U28880 ( .A(n24889), .B(n24888), .Z(n24890) );
  NAND U28881 ( .A(n24891), .B(n24890), .Z(n24892) );
  NANDN U28882 ( .A(n24893), .B(n24892), .Z(n24894) );
  NAND U28883 ( .A(n24895), .B(n24894), .Z(n24896) );
  NANDN U28884 ( .A(n24897), .B(n24896), .Z(n24898) );
  AND U28885 ( .A(n24899), .B(n24898), .Z(n24900) );
  OR U28886 ( .A(n24901), .B(n24900), .Z(n24902) );
  NAND U28887 ( .A(n24903), .B(n24902), .Z(n24904) );
  NANDN U28888 ( .A(n24905), .B(n24904), .Z(n24906) );
  NAND U28889 ( .A(n24907), .B(n24906), .Z(n24908) );
  NANDN U28890 ( .A(n24909), .B(n24908), .Z(n24910) );
  AND U28891 ( .A(n24911), .B(n24910), .Z(n24912) );
  OR U28892 ( .A(n24913), .B(n24912), .Z(n24914) );
  NAND U28893 ( .A(n24915), .B(n24914), .Z(n24916) );
  NANDN U28894 ( .A(n24917), .B(n24916), .Z(n24918) );
  NAND U28895 ( .A(n24919), .B(n24918), .Z(n24920) );
  NANDN U28896 ( .A(n24921), .B(n24920), .Z(n24922) );
  AND U28897 ( .A(n24923), .B(n24922), .Z(n24924) );
  OR U28898 ( .A(n24925), .B(n24924), .Z(n24926) );
  NAND U28899 ( .A(n24927), .B(n24926), .Z(n24928) );
  NANDN U28900 ( .A(n24929), .B(n24928), .Z(n24930) );
  NAND U28901 ( .A(n24931), .B(n24930), .Z(n24932) );
  NANDN U28902 ( .A(n24933), .B(n24932), .Z(n24934) );
  AND U28903 ( .A(n24935), .B(n24934), .Z(n24936) );
  OR U28904 ( .A(n24937), .B(n24936), .Z(n24938) );
  NAND U28905 ( .A(n24939), .B(n24938), .Z(n24940) );
  NANDN U28906 ( .A(n24941), .B(n24940), .Z(n24942) );
  NAND U28907 ( .A(n24943), .B(n24942), .Z(n24944) );
  NANDN U28908 ( .A(n24945), .B(n24944), .Z(n24946) );
  AND U28909 ( .A(n24947), .B(n24946), .Z(n24948) );
  OR U28910 ( .A(n24949), .B(n24948), .Z(n24950) );
  NAND U28911 ( .A(n24951), .B(n24950), .Z(n24952) );
  NANDN U28912 ( .A(n24953), .B(n24952), .Z(n24954) );
  NAND U28913 ( .A(n24955), .B(n24954), .Z(n24956) );
  NANDN U28914 ( .A(n24957), .B(n24956), .Z(n24958) );
  AND U28915 ( .A(n24959), .B(n24958), .Z(n24960) );
  OR U28916 ( .A(n24961), .B(n24960), .Z(n24962) );
  NAND U28917 ( .A(n24963), .B(n24962), .Z(n24964) );
  NANDN U28918 ( .A(n24965), .B(n24964), .Z(n24966) );
  NAND U28919 ( .A(n24967), .B(n24966), .Z(n24968) );
  NANDN U28920 ( .A(n24969), .B(n24968), .Z(n24970) );
  AND U28921 ( .A(n24971), .B(n24970), .Z(n24972) );
  OR U28922 ( .A(n24973), .B(n24972), .Z(n24974) );
  NAND U28923 ( .A(n24975), .B(n24974), .Z(n24976) );
  NANDN U28924 ( .A(n24977), .B(n24976), .Z(n24978) );
  NAND U28925 ( .A(n24979), .B(n24978), .Z(n24980) );
  NANDN U28926 ( .A(n24981), .B(n24980), .Z(n24982) );
  AND U28927 ( .A(n24983), .B(n24982), .Z(n24984) );
  OR U28928 ( .A(n24985), .B(n24984), .Z(n24986) );
  NAND U28929 ( .A(n24987), .B(n24986), .Z(n24988) );
  NANDN U28930 ( .A(n24989), .B(n24988), .Z(n24990) );
  NAND U28931 ( .A(n24991), .B(n24990), .Z(n24992) );
  NANDN U28932 ( .A(n24993), .B(n24992), .Z(n24994) );
  AND U28933 ( .A(n24995), .B(n24994), .Z(n24996) );
  OR U28934 ( .A(n24997), .B(n24996), .Z(n24998) );
  NAND U28935 ( .A(n24999), .B(n24998), .Z(n25000) );
  NANDN U28936 ( .A(n25001), .B(n25000), .Z(n25002) );
  NAND U28937 ( .A(n25003), .B(n25002), .Z(n25004) );
  NANDN U28938 ( .A(n25005), .B(n25004), .Z(n25006) );
  AND U28939 ( .A(n25007), .B(n25006), .Z(n25008) );
  OR U28940 ( .A(n25009), .B(n25008), .Z(n25010) );
  NAND U28941 ( .A(n25011), .B(n25010), .Z(n25012) );
  NANDN U28942 ( .A(n25013), .B(n25012), .Z(n25014) );
  NAND U28943 ( .A(n25015), .B(n25014), .Z(n25016) );
  NANDN U28944 ( .A(n25017), .B(n25016), .Z(n25018) );
  AND U28945 ( .A(n25019), .B(n25018), .Z(n25020) );
  OR U28946 ( .A(n25021), .B(n25020), .Z(n25022) );
  NAND U28947 ( .A(n25023), .B(n25022), .Z(n25024) );
  NANDN U28948 ( .A(n25025), .B(n25024), .Z(n25026) );
  NAND U28949 ( .A(n25027), .B(n25026), .Z(n25028) );
  NANDN U28950 ( .A(n25029), .B(n25028), .Z(n25030) );
  AND U28951 ( .A(n25031), .B(n25030), .Z(n25032) );
  OR U28952 ( .A(n25033), .B(n25032), .Z(n25034) );
  NAND U28953 ( .A(n25035), .B(n25034), .Z(n25036) );
  NANDN U28954 ( .A(n25037), .B(n25036), .Z(n25038) );
  NAND U28955 ( .A(n25039), .B(n25038), .Z(n25040) );
  NANDN U28956 ( .A(n25041), .B(n25040), .Z(n25042) );
  AND U28957 ( .A(n25043), .B(n25042), .Z(n25044) );
  OR U28958 ( .A(n25045), .B(n25044), .Z(n25046) );
  NAND U28959 ( .A(n25047), .B(n25046), .Z(n25048) );
  NANDN U28960 ( .A(n25049), .B(n25048), .Z(n25050) );
  NAND U28961 ( .A(n25051), .B(n25050), .Z(n25052) );
  NANDN U28962 ( .A(n25053), .B(n25052), .Z(n25054) );
  AND U28963 ( .A(n25055), .B(n25054), .Z(n25056) );
  OR U28964 ( .A(n25057), .B(n25056), .Z(n25058) );
  NAND U28965 ( .A(n25059), .B(n25058), .Z(n25060) );
  NANDN U28966 ( .A(n25061), .B(n25060), .Z(n25062) );
  NAND U28967 ( .A(n25063), .B(n25062), .Z(n25064) );
  NANDN U28968 ( .A(n25065), .B(n25064), .Z(n25067) );
  AND U28969 ( .A(n25067), .B(n25066), .Z(n25069) );
  OR U28970 ( .A(n25069), .B(n25068), .Z(n25070) );
  NAND U28971 ( .A(n25071), .B(n25070), .Z(n25072) );
  NANDN U28972 ( .A(n25073), .B(n25072), .Z(n25074) );
  NAND U28973 ( .A(n25075), .B(n25074), .Z(n25076) );
  NANDN U28974 ( .A(n25077), .B(n25076), .Z(n25078) );
  AND U28975 ( .A(n25079), .B(n25078), .Z(n25080) );
  OR U28976 ( .A(n25081), .B(n25080), .Z(n25082) );
  NAND U28977 ( .A(n25083), .B(n25082), .Z(n25084) );
  NANDN U28978 ( .A(n25085), .B(n25084), .Z(n25086) );
  NAND U28979 ( .A(n25087), .B(n25086), .Z(n25088) );
  NANDN U28980 ( .A(n25089), .B(n25088), .Z(n25090) );
  AND U28981 ( .A(n25091), .B(n25090), .Z(n25092) );
  OR U28982 ( .A(n25093), .B(n25092), .Z(n25094) );
  NAND U28983 ( .A(n25095), .B(n25094), .Z(n25096) );
  NANDN U28984 ( .A(n25097), .B(n25096), .Z(n25098) );
  NAND U28985 ( .A(n25099), .B(n25098), .Z(n25100) );
  NANDN U28986 ( .A(n25101), .B(n25100), .Z(n25102) );
  AND U28987 ( .A(n25103), .B(n25102), .Z(n25104) );
  OR U28988 ( .A(n25105), .B(n25104), .Z(n25106) );
  NAND U28989 ( .A(n25107), .B(n25106), .Z(n25108) );
  NANDN U28990 ( .A(n25109), .B(n25108), .Z(n25110) );
  NAND U28991 ( .A(n25111), .B(n25110), .Z(n25112) );
  NANDN U28992 ( .A(n25113), .B(n25112), .Z(n25114) );
  AND U28993 ( .A(n25115), .B(n25114), .Z(n25116) );
  OR U28994 ( .A(n25117), .B(n25116), .Z(n25118) );
  NAND U28995 ( .A(n25119), .B(n25118), .Z(n25120) );
  NANDN U28996 ( .A(n25121), .B(n25120), .Z(n25122) );
  NAND U28997 ( .A(n25123), .B(n25122), .Z(n25124) );
  NANDN U28998 ( .A(n25125), .B(n25124), .Z(n25126) );
  AND U28999 ( .A(n25127), .B(n25126), .Z(n25128) );
  OR U29000 ( .A(n25129), .B(n25128), .Z(n25130) );
  NAND U29001 ( .A(n25131), .B(n25130), .Z(n25132) );
  NANDN U29002 ( .A(n25133), .B(n25132), .Z(n25134) );
  NAND U29003 ( .A(n25135), .B(n25134), .Z(n25136) );
  NANDN U29004 ( .A(n25137), .B(n25136), .Z(n25138) );
  AND U29005 ( .A(n25139), .B(n25138), .Z(n25140) );
  OR U29006 ( .A(n25141), .B(n25140), .Z(n25142) );
  NAND U29007 ( .A(n25143), .B(n25142), .Z(n25144) );
  NANDN U29008 ( .A(n25145), .B(n25144), .Z(n25146) );
  NAND U29009 ( .A(n25147), .B(n25146), .Z(n25148) );
  NANDN U29010 ( .A(n25149), .B(n25148), .Z(n25150) );
  AND U29011 ( .A(n25151), .B(n25150), .Z(n25152) );
  OR U29012 ( .A(n25153), .B(n25152), .Z(n25154) );
  NAND U29013 ( .A(n25155), .B(n25154), .Z(n25156) );
  NANDN U29014 ( .A(n25157), .B(n25156), .Z(n25158) );
  NAND U29015 ( .A(n25159), .B(n25158), .Z(n25160) );
  NANDN U29016 ( .A(n25161), .B(n25160), .Z(n25162) );
  AND U29017 ( .A(n25163), .B(n25162), .Z(n25164) );
  OR U29018 ( .A(n25165), .B(n25164), .Z(n25166) );
  NAND U29019 ( .A(n25167), .B(n25166), .Z(n25168) );
  NANDN U29020 ( .A(n25169), .B(n25168), .Z(n25170) );
  NAND U29021 ( .A(n25171), .B(n25170), .Z(n25172) );
  NANDN U29022 ( .A(n25173), .B(n25172), .Z(n25174) );
  AND U29023 ( .A(n25175), .B(n25174), .Z(n25176) );
  OR U29024 ( .A(n25177), .B(n25176), .Z(n25178) );
  NAND U29025 ( .A(n25179), .B(n25178), .Z(n25180) );
  NANDN U29026 ( .A(n25181), .B(n25180), .Z(n25182) );
  NAND U29027 ( .A(n25183), .B(n25182), .Z(n25184) );
  NANDN U29028 ( .A(n25185), .B(n25184), .Z(n25186) );
  AND U29029 ( .A(n25187), .B(n25186), .Z(n25188) );
  OR U29030 ( .A(n25189), .B(n25188), .Z(n25190) );
  NAND U29031 ( .A(n25191), .B(n25190), .Z(n25192) );
  NANDN U29032 ( .A(n25193), .B(n25192), .Z(n25194) );
  NAND U29033 ( .A(n25195), .B(n25194), .Z(n25196) );
  NANDN U29034 ( .A(n25197), .B(n25196), .Z(n25198) );
  AND U29035 ( .A(n25199), .B(n25198), .Z(n25200) );
  OR U29036 ( .A(n25201), .B(n25200), .Z(n25202) );
  NAND U29037 ( .A(n25203), .B(n25202), .Z(n25204) );
  NANDN U29038 ( .A(n25205), .B(n25204), .Z(n25206) );
  NAND U29039 ( .A(n25207), .B(n25206), .Z(n25208) );
  NAND U29040 ( .A(n25209), .B(n25208), .Z(n25210) );
  AND U29041 ( .A(n25211), .B(n25210), .Z(n25212) );
  OR U29042 ( .A(n25213), .B(n25212), .Z(n25214) );
  NAND U29043 ( .A(n25215), .B(n25214), .Z(n25216) );
  NANDN U29044 ( .A(n25217), .B(n25216), .Z(n25218) );
  NAND U29045 ( .A(n25219), .B(n25218), .Z(n25220) );
  NANDN U29046 ( .A(n25221), .B(n25220), .Z(n25222) );
  AND U29047 ( .A(n25223), .B(n25222), .Z(n25224) );
  OR U29048 ( .A(n25225), .B(n25224), .Z(n25226) );
  NAND U29049 ( .A(n25227), .B(n25226), .Z(n25228) );
  NANDN U29050 ( .A(n25229), .B(n25228), .Z(n25230) );
  NAND U29051 ( .A(n25231), .B(n25230), .Z(n25232) );
  NANDN U29052 ( .A(n25253), .B(n25252), .Z(n25254) );
  NAND U29053 ( .A(n25255), .B(n25254), .Z(n25256) );
  NANDN U29054 ( .A(n25257), .B(n25256), .Z(n25258) );
  AND U29055 ( .A(n25259), .B(n25258), .Z(n25260) );
  OR U29056 ( .A(n25261), .B(n25260), .Z(n25262) );
  NAND U29057 ( .A(n25263), .B(n25262), .Z(n25264) );
  NANDN U29058 ( .A(n25265), .B(n25264), .Z(n25266) );
  NAND U29059 ( .A(n25267), .B(n25266), .Z(n25268) );
  NANDN U29060 ( .A(n25269), .B(n25268), .Z(n25270) );
  AND U29061 ( .A(n25271), .B(n25270), .Z(n25272) );
  OR U29062 ( .A(n25273), .B(n25272), .Z(n25274) );
  NAND U29063 ( .A(n25275), .B(n25274), .Z(n25276) );
  NANDN U29064 ( .A(n25277), .B(n25276), .Z(n25278) );
  NAND U29065 ( .A(n25279), .B(n25278), .Z(n25280) );
  NANDN U29066 ( .A(n25281), .B(n25280), .Z(n25282) );
  AND U29067 ( .A(n25283), .B(n25282), .Z(n25284) );
  OR U29068 ( .A(n25285), .B(n25284), .Z(n25286) );
  NAND U29069 ( .A(n25287), .B(n25286), .Z(n25288) );
  NANDN U29070 ( .A(n25289), .B(n25288), .Z(n25290) );
  NAND U29071 ( .A(n25291), .B(n25290), .Z(n25292) );
  NANDN U29072 ( .A(n25293), .B(n25292), .Z(n25294) );
  AND U29073 ( .A(n25295), .B(n25294), .Z(n25296) );
  OR U29074 ( .A(n25297), .B(n25296), .Z(n25298) );
  NAND U29075 ( .A(n25299), .B(n25298), .Z(n25300) );
  NANDN U29076 ( .A(n25301), .B(n25300), .Z(n25302) );
  NAND U29077 ( .A(n25303), .B(n25302), .Z(n25304) );
  NANDN U29078 ( .A(n25305), .B(n25304), .Z(n25306) );
  AND U29079 ( .A(n25307), .B(n25306), .Z(n25308) );
  OR U29080 ( .A(n25309), .B(n25308), .Z(n25310) );
  NAND U29081 ( .A(n25311), .B(n25310), .Z(n25312) );
  NANDN U29082 ( .A(n25313), .B(n25312), .Z(n25314) );
  NAND U29083 ( .A(n25315), .B(n25314), .Z(n25316) );
  NANDN U29084 ( .A(n25317), .B(n25316), .Z(n25318) );
  AND U29085 ( .A(n25319), .B(n25318), .Z(n25320) );
  OR U29086 ( .A(n25321), .B(n25320), .Z(n25322) );
  NAND U29087 ( .A(n25323), .B(n25322), .Z(n25324) );
  NANDN U29088 ( .A(n25325), .B(n25324), .Z(n25326) );
  NAND U29089 ( .A(n25327), .B(n25326), .Z(n25328) );
  NANDN U29090 ( .A(n25329), .B(n25328), .Z(n25330) );
  AND U29091 ( .A(n25331), .B(n25330), .Z(n25332) );
  OR U29092 ( .A(n25333), .B(n25332), .Z(n25334) );
  NAND U29093 ( .A(n25335), .B(n25334), .Z(n25336) );
  NANDN U29094 ( .A(n25337), .B(n25336), .Z(n25338) );
  NAND U29095 ( .A(n25339), .B(n25338), .Z(n25340) );
  NANDN U29096 ( .A(n25341), .B(n25340), .Z(n25342) );
  AND U29097 ( .A(n25343), .B(n25342), .Z(n25344) );
  OR U29098 ( .A(n25345), .B(n25344), .Z(n25346) );
  NAND U29099 ( .A(n25347), .B(n25346), .Z(n25348) );
  NANDN U29100 ( .A(n25349), .B(n25348), .Z(n25350) );
  NAND U29101 ( .A(n25351), .B(n25350), .Z(n25352) );
  NANDN U29102 ( .A(n25353), .B(n25352), .Z(n25354) );
  AND U29103 ( .A(n25355), .B(n25354), .Z(n25356) );
  OR U29104 ( .A(n25357), .B(n25356), .Z(n25358) );
  NAND U29105 ( .A(n25359), .B(n25358), .Z(n25360) );
  NANDN U29106 ( .A(n25361), .B(n25360), .Z(n25362) );
  NAND U29107 ( .A(n25363), .B(n25362), .Z(n25364) );
  NANDN U29108 ( .A(n25365), .B(n25364), .Z(n25366) );
  AND U29109 ( .A(n25367), .B(n25366), .Z(n25368) );
  OR U29110 ( .A(n25369), .B(n25368), .Z(n25370) );
  NAND U29111 ( .A(n25371), .B(n25370), .Z(n25372) );
  NANDN U29112 ( .A(n25373), .B(n25372), .Z(n25374) );
  NAND U29113 ( .A(n25375), .B(n25374), .Z(n25376) );
  NANDN U29114 ( .A(n25377), .B(n25376), .Z(n25378) );
  AND U29115 ( .A(n25379), .B(n25378), .Z(n25380) );
  OR U29116 ( .A(n25381), .B(n25380), .Z(n25382) );
  NAND U29117 ( .A(n25383), .B(n25382), .Z(n25384) );
  NANDN U29118 ( .A(n25385), .B(n25384), .Z(n25386) );
  NAND U29119 ( .A(n25387), .B(n25386), .Z(n25388) );
  NANDN U29120 ( .A(n25389), .B(n25388), .Z(n25390) );
  AND U29121 ( .A(n25391), .B(n25390), .Z(n25392) );
  OR U29122 ( .A(n25393), .B(n25392), .Z(n25394) );
  NAND U29123 ( .A(n25395), .B(n25394), .Z(n25396) );
  NANDN U29124 ( .A(n25397), .B(n25396), .Z(n25398) );
  NAND U29125 ( .A(n25399), .B(n25398), .Z(n25400) );
  NANDN U29126 ( .A(n25401), .B(n25400), .Z(n25402) );
  AND U29127 ( .A(n25403), .B(n25402), .Z(n25404) );
  OR U29128 ( .A(n25405), .B(n25404), .Z(n25406) );
  NAND U29129 ( .A(n25407), .B(n25406), .Z(n25408) );
  NANDN U29130 ( .A(n25409), .B(n25408), .Z(n25410) );
  NAND U29131 ( .A(n25411), .B(n25410), .Z(n25412) );
  NANDN U29132 ( .A(n25413), .B(n25412), .Z(n25414) );
  AND U29133 ( .A(n25415), .B(n25414), .Z(n25416) );
  OR U29134 ( .A(n25417), .B(n25416), .Z(n25418) );
  NAND U29135 ( .A(n25419), .B(n25418), .Z(n25420) );
  NANDN U29136 ( .A(n25421), .B(n25420), .Z(n25422) );
  NAND U29137 ( .A(n25423), .B(n25422), .Z(n25424) );
  NANDN U29138 ( .A(n25425), .B(n25424), .Z(n25426) );
  AND U29139 ( .A(n25427), .B(n25426), .Z(n25428) );
  OR U29140 ( .A(n25429), .B(n25428), .Z(n25430) );
  NAND U29141 ( .A(n25431), .B(n25430), .Z(n25432) );
  NANDN U29142 ( .A(n25433), .B(n25432), .Z(n25434) );
  NAND U29143 ( .A(n25435), .B(n25434), .Z(n25436) );
  NANDN U29144 ( .A(n25437), .B(n25436), .Z(n25438) );
  AND U29145 ( .A(n25439), .B(n25438), .Z(n25440) );
  OR U29146 ( .A(n25441), .B(n25440), .Z(n25442) );
  NAND U29147 ( .A(n25443), .B(n25442), .Z(n25444) );
  NANDN U29148 ( .A(n25445), .B(n25444), .Z(n25446) );
  NAND U29149 ( .A(n25447), .B(n25446), .Z(n25448) );
  NANDN U29150 ( .A(n25449), .B(n25448), .Z(n25450) );
  AND U29151 ( .A(n25451), .B(n25450), .Z(n25452) );
  OR U29152 ( .A(n25453), .B(n25452), .Z(n25454) );
  NAND U29153 ( .A(n25455), .B(n25454), .Z(n25456) );
  NANDN U29154 ( .A(n25457), .B(n25456), .Z(n25458) );
  NAND U29155 ( .A(n25459), .B(n25458), .Z(n25460) );
  NANDN U29156 ( .A(n25461), .B(n25460), .Z(n25462) );
  AND U29157 ( .A(n25463), .B(n25462), .Z(n25464) );
  OR U29158 ( .A(n25465), .B(n25464), .Z(n25466) );
  NAND U29159 ( .A(n25467), .B(n25466), .Z(n25468) );
  NANDN U29160 ( .A(n25469), .B(n25468), .Z(n25470) );
  NAND U29161 ( .A(n25471), .B(n25470), .Z(n25472) );
  NANDN U29162 ( .A(n25473), .B(n25472), .Z(n25474) );
  AND U29163 ( .A(n25475), .B(n25474), .Z(n25476) );
  OR U29164 ( .A(n25477), .B(n25476), .Z(n25478) );
  NAND U29165 ( .A(n25479), .B(n25478), .Z(n25480) );
  NANDN U29166 ( .A(n25481), .B(n25480), .Z(n25482) );
  NAND U29167 ( .A(n25483), .B(n25482), .Z(n25484) );
  NANDN U29168 ( .A(n25485), .B(n25484), .Z(n25486) );
  AND U29169 ( .A(n25487), .B(n25486), .Z(n25488) );
  OR U29170 ( .A(n25489), .B(n25488), .Z(n25490) );
  NAND U29171 ( .A(n25491), .B(n25490), .Z(n25492) );
  NANDN U29172 ( .A(n25493), .B(n25492), .Z(n25494) );
  NAND U29173 ( .A(n25495), .B(n25494), .Z(n25496) );
  NANDN U29174 ( .A(n25497), .B(n25496), .Z(n25498) );
  AND U29175 ( .A(n25499), .B(n25498), .Z(n25500) );
  OR U29176 ( .A(n25501), .B(n25500), .Z(n25502) );
  NAND U29177 ( .A(n25503), .B(n25502), .Z(n25504) );
  NANDN U29178 ( .A(n25505), .B(n25504), .Z(n25506) );
  NAND U29179 ( .A(n25507), .B(n25506), .Z(n25508) );
  NANDN U29180 ( .A(n25509), .B(n25508), .Z(n25510) );
  AND U29181 ( .A(n25511), .B(n25510), .Z(n25512) );
  OR U29182 ( .A(n25513), .B(n25512), .Z(n25514) );
  NAND U29183 ( .A(n25515), .B(n25514), .Z(n25516) );
  NANDN U29184 ( .A(n25517), .B(n25516), .Z(n25518) );
  NAND U29185 ( .A(n25519), .B(n25518), .Z(n25520) );
  NANDN U29186 ( .A(n25521), .B(n25520), .Z(n25522) );
  AND U29187 ( .A(n25523), .B(n25522), .Z(n25524) );
  OR U29188 ( .A(n25525), .B(n25524), .Z(n25526) );
  NAND U29189 ( .A(n25527), .B(n25526), .Z(n25528) );
  NANDN U29190 ( .A(n25529), .B(n25528), .Z(n25530) );
  NAND U29191 ( .A(n25531), .B(n25530), .Z(n25533) );
  NANDN U29192 ( .A(n25552), .B(n25551), .Z(n25553) );
  NAND U29193 ( .A(n25554), .B(n25553), .Z(n25555) );
  NANDN U29194 ( .A(n25556), .B(n25555), .Z(n25557) );
  AND U29195 ( .A(n25558), .B(n25557), .Z(n25559) );
  OR U29196 ( .A(n25560), .B(n25559), .Z(n25561) );
  NAND U29197 ( .A(n25562), .B(n25561), .Z(n25563) );
  NANDN U29198 ( .A(n25564), .B(n25563), .Z(n25565) );
  NAND U29199 ( .A(n25566), .B(n25565), .Z(n25567) );
  NANDN U29200 ( .A(n25568), .B(n25567), .Z(n25569) );
  AND U29201 ( .A(n25570), .B(n25569), .Z(n25571) );
  OR U29202 ( .A(n25572), .B(n25571), .Z(n25573) );
  NAND U29203 ( .A(n25574), .B(n25573), .Z(n25575) );
  NANDN U29204 ( .A(n25576), .B(n25575), .Z(n25577) );
  NAND U29205 ( .A(n25578), .B(n25577), .Z(n25579) );
  NANDN U29206 ( .A(n25580), .B(n25579), .Z(n25581) );
  AND U29207 ( .A(n25582), .B(n25581), .Z(n25583) );
  OR U29208 ( .A(n25584), .B(n25583), .Z(n25585) );
  NAND U29209 ( .A(n25586), .B(n25585), .Z(n25587) );
  NANDN U29210 ( .A(n25588), .B(n25587), .Z(n25589) );
  NAND U29211 ( .A(n25590), .B(n25589), .Z(n25591) );
  NANDN U29212 ( .A(n25592), .B(n25591), .Z(n25593) );
  AND U29213 ( .A(n25594), .B(n25593), .Z(n25595) );
  OR U29214 ( .A(n25596), .B(n25595), .Z(n25597) );
  NAND U29215 ( .A(n25598), .B(n25597), .Z(n25599) );
  NANDN U29216 ( .A(n25600), .B(n25599), .Z(n25601) );
  NAND U29217 ( .A(n25602), .B(n25601), .Z(n25603) );
  NANDN U29218 ( .A(n25604), .B(n25603), .Z(n25605) );
  AND U29219 ( .A(n25606), .B(n25605), .Z(n25607) );
  OR U29220 ( .A(n25608), .B(n25607), .Z(n25609) );
  NAND U29221 ( .A(n25610), .B(n25609), .Z(n25611) );
  NANDN U29222 ( .A(n25612), .B(n25611), .Z(n25613) );
  NAND U29223 ( .A(n25614), .B(n25613), .Z(n25615) );
  NANDN U29224 ( .A(n25616), .B(n25615), .Z(n25617) );
  AND U29225 ( .A(n25618), .B(n25617), .Z(n25619) );
  OR U29226 ( .A(n25620), .B(n25619), .Z(n25621) );
  NAND U29227 ( .A(n25622), .B(n25621), .Z(n25623) );
  NANDN U29228 ( .A(n25624), .B(n25623), .Z(n25625) );
  NAND U29229 ( .A(n25626), .B(n25625), .Z(n25627) );
  NANDN U29230 ( .A(n25628), .B(n25627), .Z(n25629) );
  AND U29231 ( .A(n25630), .B(n25629), .Z(n25631) );
  OR U29232 ( .A(n25650), .B(n25649), .Z(n25651) );
  NAND U29233 ( .A(n25652), .B(n25651), .Z(n25653) );
  NANDN U29234 ( .A(n25654), .B(n25653), .Z(n25655) );
  NAND U29235 ( .A(n25656), .B(n25655), .Z(n25657) );
  NANDN U29236 ( .A(n25658), .B(n25657), .Z(n25659) );
  AND U29237 ( .A(n25660), .B(n25659), .Z(n25661) );
  OR U29238 ( .A(n25662), .B(n25661), .Z(n25663) );
  NAND U29239 ( .A(n25664), .B(n25663), .Z(n25665) );
  NANDN U29240 ( .A(n25666), .B(n25665), .Z(n25667) );
  NAND U29241 ( .A(n25668), .B(n25667), .Z(n25669) );
  NANDN U29242 ( .A(n25670), .B(n25669), .Z(n25671) );
  AND U29243 ( .A(n25672), .B(n25671), .Z(n25673) );
  OR U29244 ( .A(n25674), .B(n25673), .Z(n25675) );
  NAND U29245 ( .A(n25676), .B(n25675), .Z(n25677) );
  NANDN U29246 ( .A(n25678), .B(n25677), .Z(n25679) );
  NAND U29247 ( .A(n25680), .B(n25679), .Z(n25681) );
  NANDN U29248 ( .A(n25682), .B(n25681), .Z(n25683) );
  AND U29249 ( .A(n25684), .B(n25683), .Z(n25685) );
  OR U29250 ( .A(n25686), .B(n25685), .Z(n25687) );
  NAND U29251 ( .A(n25688), .B(n25687), .Z(n25689) );
  NANDN U29252 ( .A(n25690), .B(n25689), .Z(n25691) );
  NAND U29253 ( .A(n25692), .B(n25691), .Z(n25693) );
  NANDN U29254 ( .A(n25694), .B(n25693), .Z(n25695) );
  AND U29255 ( .A(n25696), .B(n25695), .Z(n25697) );
  OR U29256 ( .A(n25698), .B(n25697), .Z(n25699) );
  NAND U29257 ( .A(n25700), .B(n25699), .Z(n25701) );
  NANDN U29258 ( .A(n25702), .B(n25701), .Z(n25703) );
  NAND U29259 ( .A(n25704), .B(n25703), .Z(n25705) );
  NANDN U29260 ( .A(n25706), .B(n25705), .Z(n25707) );
  AND U29261 ( .A(n25708), .B(n25707), .Z(n25709) );
  OR U29262 ( .A(n25710), .B(n25709), .Z(n25711) );
  NAND U29263 ( .A(n25712), .B(n25711), .Z(n25713) );
  NANDN U29264 ( .A(n25714), .B(n25713), .Z(n25715) );
  NAND U29265 ( .A(n25716), .B(n25715), .Z(n25717) );
  NANDN U29266 ( .A(n25718), .B(n25717), .Z(n25719) );
  AND U29267 ( .A(n25720), .B(n25719), .Z(n25721) );
  OR U29268 ( .A(n25722), .B(n25721), .Z(n25723) );
  NAND U29269 ( .A(n25724), .B(n25723), .Z(n25725) );
  NANDN U29270 ( .A(n25726), .B(n25725), .Z(n25727) );
  NAND U29271 ( .A(n25728), .B(n25727), .Z(n25729) );
  NANDN U29272 ( .A(n25730), .B(n25729), .Z(n25731) );
  AND U29273 ( .A(n25732), .B(n25731), .Z(n25733) );
  OR U29274 ( .A(n25734), .B(n25733), .Z(n25735) );
  NAND U29275 ( .A(n25736), .B(n25735), .Z(n25737) );
  NANDN U29276 ( .A(n25738), .B(n25737), .Z(n25739) );
  NAND U29277 ( .A(n25740), .B(n25739), .Z(n25741) );
  NANDN U29278 ( .A(n25742), .B(n25741), .Z(n25743) );
  AND U29279 ( .A(n25744), .B(n25743), .Z(n25745) );
  OR U29280 ( .A(n25746), .B(n25745), .Z(n25747) );
  NAND U29281 ( .A(n25748), .B(n25747), .Z(n25749) );
  NANDN U29282 ( .A(n25750), .B(n25749), .Z(n25751) );
  NAND U29283 ( .A(n25752), .B(n25751), .Z(n25753) );
  NANDN U29284 ( .A(n25754), .B(n25753), .Z(n25755) );
  AND U29285 ( .A(n25756), .B(n25755), .Z(n25757) );
  OR U29286 ( .A(n25758), .B(n25757), .Z(n25759) );
  NAND U29287 ( .A(n25760), .B(n25759), .Z(n25761) );
  NANDN U29288 ( .A(n25762), .B(n25761), .Z(n25763) );
  NAND U29289 ( .A(n25764), .B(n25763), .Z(n25765) );
  NANDN U29290 ( .A(n25766), .B(n25765), .Z(n25767) );
  AND U29291 ( .A(n25768), .B(n25767), .Z(n25769) );
  OR U29292 ( .A(n25770), .B(n25769), .Z(n25771) );
  NAND U29293 ( .A(n25772), .B(n25771), .Z(n25773) );
  NANDN U29294 ( .A(n25774), .B(n25773), .Z(n25775) );
  NAND U29295 ( .A(n25776), .B(n25775), .Z(n25777) );
  NANDN U29296 ( .A(n25778), .B(n25777), .Z(n25779) );
  AND U29297 ( .A(n25780), .B(n25779), .Z(n25781) );
  OR U29298 ( .A(n25782), .B(n25781), .Z(n25783) );
  NAND U29299 ( .A(n25784), .B(n25783), .Z(n25785) );
  NANDN U29300 ( .A(n25786), .B(n25785), .Z(n25787) );
  NAND U29301 ( .A(n25788), .B(n25787), .Z(n25789) );
  NANDN U29302 ( .A(n25790), .B(n25789), .Z(n25791) );
  AND U29303 ( .A(n25792), .B(n25791), .Z(n25793) );
  OR U29304 ( .A(n25794), .B(n25793), .Z(n25795) );
  NAND U29305 ( .A(n25796), .B(n25795), .Z(n25797) );
  NANDN U29306 ( .A(n25798), .B(n25797), .Z(n25799) );
  NAND U29307 ( .A(n25800), .B(n25799), .Z(n25801) );
  NANDN U29308 ( .A(n25802), .B(n25801), .Z(n25803) );
  AND U29309 ( .A(n25804), .B(n25803), .Z(n25805) );
  OR U29310 ( .A(n25806), .B(n25805), .Z(n25807) );
  NAND U29311 ( .A(n25808), .B(n25807), .Z(n25809) );
  NANDN U29312 ( .A(n25810), .B(n25809), .Z(n25811) );
  NAND U29313 ( .A(n25812), .B(n25811), .Z(n25813) );
  NANDN U29314 ( .A(n25814), .B(n25813), .Z(n25815) );
  AND U29315 ( .A(n25816), .B(n25815), .Z(n25817) );
  OR U29316 ( .A(n25818), .B(n25817), .Z(n25819) );
  NAND U29317 ( .A(n25820), .B(n25819), .Z(n25821) );
  NANDN U29318 ( .A(n25822), .B(n25821), .Z(n25823) );
  NAND U29319 ( .A(n25824), .B(n25823), .Z(n25825) );
  NANDN U29320 ( .A(n25826), .B(n25825), .Z(n25827) );
  AND U29321 ( .A(n25828), .B(n25827), .Z(n25829) );
  OR U29322 ( .A(n25830), .B(n25829), .Z(n25831) );
  NAND U29323 ( .A(n25832), .B(n25831), .Z(n25833) );
  NANDN U29324 ( .A(n25834), .B(n25833), .Z(n25835) );
  NAND U29325 ( .A(n25836), .B(n25835), .Z(n25837) );
  NANDN U29326 ( .A(n25838), .B(n25837), .Z(n25839) );
  AND U29327 ( .A(n25840), .B(n25839), .Z(n25841) );
  OR U29328 ( .A(n25842), .B(n25841), .Z(n25843) );
  NAND U29329 ( .A(n25844), .B(n25843), .Z(n25845) );
  NANDN U29330 ( .A(n25846), .B(n25845), .Z(n25847) );
  NAND U29331 ( .A(n25848), .B(n25847), .Z(n25849) );
  IV U29332 ( .A(n25909), .Z(n25910) );
  AND U29333 ( .A(n25953), .B(n25952), .Z(n25954) );
  OR U29334 ( .A(n25955), .B(n25954), .Z(n25956) );
  NAND U29335 ( .A(n25957), .B(n25956), .Z(n25958) );
  NANDN U29336 ( .A(n25959), .B(n25958), .Z(n25960) );
  NAND U29337 ( .A(n25961), .B(n25960), .Z(n25962) );
  NANDN U29338 ( .A(n25963), .B(n25962), .Z(n25964) );
  AND U29339 ( .A(n25965), .B(n25964), .Z(n25966) );
  OR U29340 ( .A(n25967), .B(n25966), .Z(n25968) );
  NAND U29341 ( .A(n25969), .B(n25968), .Z(n25970) );
  NANDN U29342 ( .A(n25971), .B(n25970), .Z(n25972) );
  NAND U29343 ( .A(n25973), .B(n25972), .Z(n25974) );
  NANDN U29344 ( .A(n25975), .B(n25974), .Z(n25976) );
  AND U29345 ( .A(n25977), .B(n25976), .Z(n25978) );
  OR U29346 ( .A(n25979), .B(n25978), .Z(n25980) );
  NAND U29347 ( .A(n25981), .B(n25980), .Z(n25982) );
  NANDN U29348 ( .A(n25983), .B(n25982), .Z(n25984) );
  NAND U29349 ( .A(n25985), .B(n25984), .Z(n25986) );
  NANDN U29350 ( .A(n25987), .B(n25986), .Z(n25988) );
  AND U29351 ( .A(n25989), .B(n25988), .Z(n25991) );
  OR U29352 ( .A(n25991), .B(n25990), .Z(n25992) );
  AND U29353 ( .A(n25993), .B(n25992), .Z(n25994) );
  OR U29354 ( .A(n25995), .B(n25994), .Z(n25996) );
  NAND U29355 ( .A(n25997), .B(n25996), .Z(n25998) );
  NANDN U29356 ( .A(n25999), .B(n25998), .Z(n26001) );
  NAND U29357 ( .A(n26001), .B(n26000), .Z(n26002) );
  NANDN U29358 ( .A(n26003), .B(n26002), .Z(n26004) );
  AND U29359 ( .A(n26005), .B(n26004), .Z(n26007) );
  OR U29360 ( .A(n26007), .B(n26006), .Z(n26008) );
  NAND U29361 ( .A(n26009), .B(n26008), .Z(n26010) );
  NAND U29362 ( .A(n26011), .B(n26010), .Z(n26013) );
  NAND U29363 ( .A(n26013), .B(n26012), .Z(n26014) );
  NAND U29364 ( .A(n26015), .B(n26014), .Z(n26016) );
  AND U29365 ( .A(n26017), .B(n26016), .Z(n26018) );
  OR U29366 ( .A(n26019), .B(n26018), .Z(n26020) );
  NAND U29367 ( .A(n26021), .B(n26020), .Z(n26022) );
  NANDN U29368 ( .A(n26023), .B(n26022), .Z(n26024) );
  NAND U29369 ( .A(n26025), .B(n26024), .Z(n26026) );
  NANDN U29370 ( .A(n26027), .B(n26026), .Z(n26028) );
  AND U29371 ( .A(n26029), .B(n26028), .Z(n26030) );
  OR U29372 ( .A(n26031), .B(n26030), .Z(n26032) );
  IV U29373 ( .A(n26079), .Z(n26080) );
  IV U29374 ( .A(n26093), .Z(n26094) );
  IV U29375 ( .A(n26187), .Z(n26188) );
  IV U29376 ( .A(n26229), .Z(n26230) );
  IV U29377 ( .A(n26303), .Z(n26304) );
  IV U29378 ( .A(n26355), .Z(n26356) );
  IV U29379 ( .A(n26394), .Z(n26395) );
  NAND U29380 ( .A(n26406), .B(n26405), .Z(n26407) );
  NANDN U29381 ( .A(n26408), .B(n26407), .Z(n26410) );
  NAND U29382 ( .A(n26410), .B(n26409), .Z(n26411) );
  NANDN U29383 ( .A(n26412), .B(n26411), .Z(n26413) );
  AND U29384 ( .A(n26414), .B(n26413), .Z(n26415) );
  OR U29385 ( .A(n26416), .B(n26415), .Z(n26417) );
  NAND U29386 ( .A(n26418), .B(n26417), .Z(n26419) );
  NANDN U29387 ( .A(n26420), .B(n26419), .Z(n26421) );
  NAND U29388 ( .A(n26422), .B(n26421), .Z(n26423) );
  NANDN U29389 ( .A(n26424), .B(n26423), .Z(n26426) );
  AND U29390 ( .A(n26426), .B(n26425), .Z(n26428) );
  OR U29391 ( .A(n26428), .B(n26427), .Z(n26429) );
  NAND U29392 ( .A(n26430), .B(n26429), .Z(n26431) );
  NANDN U29393 ( .A(n26432), .B(n26431), .Z(n26433) );
  NAND U29394 ( .A(n26434), .B(n26433), .Z(n26435) );
  AND U29395 ( .A(n26436), .B(n26435), .Z(n26438) );
  NANDN U29396 ( .A(n26438), .B(n26437), .Z(n26439) );
  NAND U29397 ( .A(n26440), .B(n26439), .Z(n26441) );
  NAND U29398 ( .A(n26442), .B(n26441), .Z(n26444) );
  NAND U29399 ( .A(n26444), .B(n26443), .Z(n26445) );
  IV U29400 ( .A(n26517), .Z(n26518) );
  IV U29401 ( .A(n26573), .Z(n26574) );
  NANDN U29402 ( .A(n26605), .B(n26604), .Z(n26607) );
  AND U29403 ( .A(n26607), .B(n26606), .Z(n26609) );
  NANDN U29404 ( .A(n26609), .B(n26608), .Z(n26610) );
  NAND U29405 ( .A(n26611), .B(n26610), .Z(n26612) );
  NANDN U29406 ( .A(n26613), .B(n26612), .Z(n26615) );
  NAND U29407 ( .A(n26615), .B(n26614), .Z(n26616) );
  NANDN U29408 ( .A(n26617), .B(n26616), .Z(n26618) );
  AND U29409 ( .A(n26619), .B(n26618), .Z(n26620) );
  OR U29410 ( .A(n26621), .B(n26620), .Z(n26622) );
  NAND U29411 ( .A(n26623), .B(n26622), .Z(n26624) );
  NANDN U29412 ( .A(n26625), .B(n26624), .Z(n26626) );
  NANDN U29413 ( .A(n26627), .B(n26626), .Z(n26628) );
  AND U29414 ( .A(n26629), .B(n26628), .Z(n26631) );
  NANDN U29415 ( .A(n26631), .B(n26630), .Z(n26632) );
  NAND U29416 ( .A(n26633), .B(n26632), .Z(n26634) );
  NAND U29417 ( .A(n26635), .B(n26634), .Z(n26636) );
  NANDN U29418 ( .A(n26637), .B(n26636), .Z(n26638) );
  AND U29419 ( .A(n26639), .B(n26638), .Z(n26640) );
  OR U29420 ( .A(n26641), .B(n26640), .Z(n26642) );
  NAND U29421 ( .A(n26643), .B(n26642), .Z(n26644) );
  IV U29422 ( .A(n26881), .Z(n26882) );
  IV U29423 ( .A(n26884), .Z(n26885) );
  IV U29424 ( .A(n27037), .Z(n27038) );
  IV U29425 ( .A(n27054), .Z(n27055) );
  IV U29426 ( .A(n27084), .Z(n27085) );
  AND U29427 ( .A(n27129), .B(n27128), .Z(n27130) );
  OR U29428 ( .A(n27131), .B(n27130), .Z(n27132) );
  NAND U29429 ( .A(n27133), .B(n27132), .Z(n27134) );
  NANDN U29430 ( .A(n27135), .B(n27134), .Z(n27137) );
  NAND U29431 ( .A(n27137), .B(n27136), .Z(n27138) );
  NANDN U29432 ( .A(n27139), .B(n27138), .Z(n27140) );
  AND U29433 ( .A(n27141), .B(n27140), .Z(n27142) );
  OR U29434 ( .A(n27143), .B(n27142), .Z(n27144) );
  NAND U29435 ( .A(n27145), .B(n27144), .Z(n27146) );
  NANDN U29436 ( .A(n27147), .B(n27146), .Z(n27148) );
  NAND U29437 ( .A(n27149), .B(n27148), .Z(n27151) );
  AND U29438 ( .A(n27151), .B(n27150), .Z(n27153) );
  NANDN U29439 ( .A(n27153), .B(n27152), .Z(n27155) );
  ANDN U29440 ( .B(n27155), .A(n27154), .Z(n27157) );
  OR U29441 ( .A(n27157), .B(n27156), .Z(n27158) );
  AND U29442 ( .A(n27159), .B(n27158), .Z(n27161) );
  NANDN U29443 ( .A(n27161), .B(n27160), .Z(n27162) );
  AND U29444 ( .A(n27163), .B(n27162), .Z(n27165) );
  OR U29445 ( .A(n27165), .B(n27164), .Z(n27166) );
  AND U29446 ( .A(n27167), .B(n27166), .Z(n27168) );
  IV U29447 ( .A(n27207), .Z(n27208) );
  IV U29448 ( .A(n27235), .Z(n27236) );
  IV U29449 ( .A(n27454), .Z(n27455) );
  IV U29450 ( .A(n27471), .Z(n27472) );
  IV U29451 ( .A(n27530), .Z(n27531) );
  IV U29452 ( .A(n27570), .Z(n27571) );
  IV U29453 ( .A(n27627), .Z(n27628) );
  IV U29454 ( .A(n27647), .Z(n27648) );
  AND U29455 ( .A(n27674), .B(n27673), .Z(n27680) );
  NANDN U29456 ( .A(n27676), .B(n27675), .Z(n27678) );
  ANDN U29457 ( .B(n27678), .A(n27677), .Z(n27679) );
  NANDN U29458 ( .A(n27680), .B(n27679), .Z(n27681) );
  NAND U29459 ( .A(n27682), .B(n27681), .Z(n27683) );
  NANDN U29460 ( .A(n27684), .B(n27683), .Z(n27686) );
  AND U29461 ( .A(n27686), .B(n27685), .Z(n27688) );
  OR U29462 ( .A(n27688), .B(n27687), .Z(n27689) );
  NANDN U29463 ( .A(n27690), .B(n27689), .Z(n27691) );
  AND U29464 ( .A(n27692), .B(n27691), .Z(n27694) );
  NANDN U29465 ( .A(n27694), .B(n27693), .Z(n27696) );
  AND U29466 ( .A(n27696), .B(n27695), .Z(n27698) );
  OR U29467 ( .A(n27698), .B(n27697), .Z(n27699) );
  AND U29468 ( .A(n27700), .B(n27699), .Z(n27701) );
  OR U29469 ( .A(n27702), .B(n27701), .Z(n27703) );
  NAND U29470 ( .A(n27704), .B(n27703), .Z(n27705) );
  NANDN U29471 ( .A(n27706), .B(n27705), .Z(n27707) );
  NANDN U29472 ( .A(n27708), .B(n27707), .Z(n27709) );
  AND U29473 ( .A(n27710), .B(n27709), .Z(n27711) );
  OR U29474 ( .A(n27712), .B(n27711), .Z(n27713) );
  NAND U29475 ( .A(n27714), .B(n27713), .Z(n27715) );
  NANDN U29476 ( .A(n27716), .B(n27715), .Z(n27717) );
  IV U29477 ( .A(n27719), .Z(n27720) );
  IV U29478 ( .A(n27775), .Z(n27776) );
  IV U29479 ( .A(n27778), .Z(n27779) );
  XNOR U29480 ( .A(x[2450]), .B(n27823), .Z(n27824) );
  IV U29481 ( .A(n27861), .Z(n27863) );
  IV U29482 ( .A(n27956), .Z(n27958) );
  IV U29483 ( .A(n28005), .Z(n28007) );
  OR U29484 ( .A(n28025), .B(n28024), .Z(n28028) );
  IV U29485 ( .A(n28026), .Z(n28027) );
  IV U29486 ( .A(n28127), .Z(n28128) );
  IV U29487 ( .A(n28182), .Z(n28183) );
  IV U29488 ( .A(n28185), .Z(n28186) );
  IV U29489 ( .A(n28224), .Z(n28225) );
  IV U29490 ( .A(n28227), .Z(n28228) );
  NAND U29491 ( .A(n28257), .B(n28256), .Z(n28258) );
  NAND U29492 ( .A(n28259), .B(n28258), .Z(n28263) );
  NAND U29493 ( .A(n28261), .B(n28260), .Z(n28262) );
  NANDN U29494 ( .A(n28263), .B(n28262), .Z(n28264) );
  AND U29495 ( .A(n28265), .B(n28264), .Z(n28266) );
  OR U29496 ( .A(n28267), .B(n28266), .Z(n28268) );
  NAND U29497 ( .A(n28269), .B(n28268), .Z(n28270) );
  NANDN U29498 ( .A(n28271), .B(n28270), .Z(n28272) );
  AND U29499 ( .A(n28273), .B(n28272), .Z(n28275) );
  NANDN U29500 ( .A(n28275), .B(n28274), .Z(n28276) );
  NAND U29501 ( .A(n28277), .B(n28276), .Z(n28278) );
  NANDN U29502 ( .A(n28279), .B(n28278), .Z(n28281) );
  AND U29503 ( .A(n28281), .B(n28280), .Z(n28283) );
  OR U29504 ( .A(n28283), .B(n28282), .Z(n28284) );
  NANDN U29505 ( .A(n28285), .B(n28284), .Z(n28286) );
  AND U29506 ( .A(n28287), .B(n28286), .Z(n28289) );
  OR U29507 ( .A(n28289), .B(n28288), .Z(n28291) );
  ANDN U29508 ( .B(n28291), .A(n28290), .Z(n28293) );
  NANDN U29509 ( .A(n28293), .B(n28292), .Z(n28294) );
  NAND U29510 ( .A(n28295), .B(n28294), .Z(n28296) );
  IV U29511 ( .A(n28361), .Z(n28362) );
  IV U29512 ( .A(n28376), .Z(n28377) );
  OR U29513 ( .A(n28515), .B(n28514), .Z(n28516) );
  IV U29514 ( .A(n28628), .Z(n28629) );
  IV U29515 ( .A(n28733), .Z(n28734) );
  IV U29516 ( .A(n28757), .Z(n28758) );
  IV U29517 ( .A(n28770), .Z(n28771) );
  IV U29518 ( .A(n28790), .Z(n28791) );
  IV U29519 ( .A(n28793), .Z(n28794) );
  IV U29520 ( .A(n28819), .Z(n28820) );
  IV U29521 ( .A(n28976), .Z(n28977) );
  IV U29522 ( .A(n29018), .Z(n29019) );
  IV U29523 ( .A(n29066), .Z(n29067) );
  IV U29524 ( .A(n29105), .Z(n29106) );
  IV U29525 ( .A(n29133), .Z(n29134) );
  IV U29526 ( .A(n29175), .Z(n29176) );
  IV U29527 ( .A(n29186), .Z(n29187) );
  IV U29528 ( .A(n29263), .Z(n29264) );
  IV U29529 ( .A(n29374), .Z(n29375) );
  IV U29530 ( .A(n29407), .Z(n29408) );
  IV U29531 ( .A(n29418), .Z(n29419) );
  IV U29532 ( .A(n29421), .Z(n29422) );
  IV U29533 ( .A(n29466), .Z(n29467) );
  IV U29534 ( .A(n29474), .Z(n29475) );
  IV U29535 ( .A(n29497), .Z(n29498) );
  IV U29536 ( .A(n29511), .Z(n29512) );
endmodule

