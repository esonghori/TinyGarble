
module mult_N64_CC4 ( clk, rst, a, b, c );
  input [63:0] a;
  input [15:0] b;
  output [127:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153;
  wire   [127:0] sreg;

  DFF \sreg_reg[111]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(sreg[111]) );
  DFF \sreg_reg[110]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(sreg[110]) );
  DFF \sreg_reg[109]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(sreg[109]) );
  DFF \sreg_reg[108]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(sreg[108]) );
  DFF \sreg_reg[107]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(sreg[107]) );
  DFF \sreg_reg[106]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(sreg[106]) );
  DFF \sreg_reg[105]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(sreg[105]) );
  DFF \sreg_reg[104]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(sreg[104]) );
  DFF \sreg_reg[103]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(sreg[103]) );
  DFF \sreg_reg[102]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(sreg[102]) );
  DFF \sreg_reg[101]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(sreg[101]) );
  DFF \sreg_reg[100]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(sreg[100]) );
  DFF \sreg_reg[99]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(sreg[99]) );
  DFF \sreg_reg[98]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(sreg[98]) );
  DFF \sreg_reg[97]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(sreg[97]) );
  DFF \sreg_reg[96]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(sreg[96]) );
  DFF \sreg_reg[95]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(sreg[95]) );
  DFF \sreg_reg[94]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(sreg[94]) );
  DFF \sreg_reg[93]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(sreg[93]) );
  DFF \sreg_reg[92]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(sreg[92]) );
  DFF \sreg_reg[91]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(sreg[91]) );
  DFF \sreg_reg[90]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(sreg[90]) );
  DFF \sreg_reg[89]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(sreg[89]) );
  DFF \sreg_reg[88]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(sreg[88]) );
  DFF \sreg_reg[87]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(sreg[87]) );
  DFF \sreg_reg[86]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(sreg[86]) );
  DFF \sreg_reg[85]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(sreg[85]) );
  DFF \sreg_reg[84]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(sreg[84]) );
  DFF \sreg_reg[83]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(sreg[83]) );
  DFF \sreg_reg[82]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(sreg[82]) );
  DFF \sreg_reg[81]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(sreg[81]) );
  DFF \sreg_reg[80]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(sreg[80]) );
  DFF \sreg_reg[79]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(sreg[79]) );
  DFF \sreg_reg[78]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(sreg[78]) );
  DFF \sreg_reg[77]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(sreg[77]) );
  DFF \sreg_reg[76]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(sreg[76]) );
  DFF \sreg_reg[75]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(sreg[75]) );
  DFF \sreg_reg[74]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(sreg[74]) );
  DFF \sreg_reg[73]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(sreg[73]) );
  DFF \sreg_reg[72]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(sreg[72]) );
  DFF \sreg_reg[71]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(sreg[71]) );
  DFF \sreg_reg[70]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(sreg[70]) );
  DFF \sreg_reg[69]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(sreg[69]) );
  DFF \sreg_reg[68]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(sreg[68]) );
  DFF \sreg_reg[67]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(sreg[67]) );
  DFF \sreg_reg[66]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(sreg[66]) );
  DFF \sreg_reg[65]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(sreg[65]) );
  DFF \sreg_reg[64]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(sreg[64]) );
  DFF \sreg_reg[63]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(sreg[63]) );
  DFF \sreg_reg[62]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(sreg[62]) );
  DFF \sreg_reg[61]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(sreg[61]) );
  DFF \sreg_reg[60]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(sreg[60]) );
  DFF \sreg_reg[59]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(sreg[59]) );
  DFF \sreg_reg[58]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(sreg[58]) );
  DFF \sreg_reg[57]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(sreg[57]) );
  DFF \sreg_reg[56]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(sreg[56]) );
  DFF \sreg_reg[55]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(sreg[55]) );
  DFF \sreg_reg[54]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(sreg[54]) );
  DFF \sreg_reg[53]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(sreg[53]) );
  DFF \sreg_reg[52]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(sreg[52]) );
  DFF \sreg_reg[51]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(sreg[51]) );
  DFF \sreg_reg[50]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(sreg[50]) );
  DFF \sreg_reg[49]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(sreg[49]) );
  DFF \sreg_reg[48]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(sreg[48]) );
  DFF \sreg_reg[47]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[0]) );
  OR U19 ( .A(n4691), .B(n4692), .Z(n1) );
  NANDN U20 ( .A(n4693), .B(n4694), .Z(n2) );
  NAND U21 ( .A(n1), .B(n2), .Z(n4761) );
  NANDN U22 ( .A(n1363), .B(n1362), .Z(n3) );
  NANDN U23 ( .A(n1364), .B(n1365), .Z(n4) );
  NAND U24 ( .A(n3), .B(n4), .Z(n1402) );
  NANDN U25 ( .A(n3741), .B(n3740), .Z(n5) );
  NANDN U26 ( .A(n3742), .B(n3743), .Z(n6) );
  NAND U27 ( .A(n5), .B(n6), .Z(n3829) );
  OR U28 ( .A(n4760), .B(n4759), .Z(n7) );
  NANDN U29 ( .A(n4761), .B(n4762), .Z(n8) );
  AND U30 ( .A(n7), .B(n8), .Z(n4775) );
  NANDN U31 ( .A(n820), .B(n819), .Z(n9) );
  NANDN U32 ( .A(n817), .B(n818), .Z(n10) );
  NAND U33 ( .A(n9), .B(n10), .Z(n931) );
  OR U34 ( .A(n1366), .B(n1367), .Z(n11) );
  NANDN U35 ( .A(n1368), .B(n1369), .Z(n12) );
  NAND U36 ( .A(n11), .B(n12), .Z(n1403) );
  OR U37 ( .A(n1583), .B(n1584), .Z(n13) );
  NANDN U38 ( .A(n1585), .B(n1586), .Z(n14) );
  NAND U39 ( .A(n13), .B(n14), .Z(n1622) );
  OR U40 ( .A(n3830), .B(n3831), .Z(n15) );
  OR U41 ( .A(n3828), .B(n3829), .Z(n16) );
  AND U42 ( .A(n15), .B(n16), .Z(n3906) );
  NANDN U43 ( .A(n4169), .B(n4168), .Z(n17) );
  NANDN U44 ( .A(n4170), .B(n4171), .Z(n18) );
  NAND U45 ( .A(n17), .B(n18), .Z(n4225) );
  NANDN U46 ( .A(n4752), .B(n4787), .Z(n19) );
  NANDN U47 ( .A(n4753), .B(n4754), .Z(n20) );
  NAND U48 ( .A(n19), .B(n20), .Z(n4780) );
  NANDN U49 ( .A(n1248), .B(n1247), .Z(n21) );
  NANDN U50 ( .A(n1249), .B(n1250), .Z(n22) );
  NAND U51 ( .A(n21), .B(n22), .Z(n1324) );
  OR U52 ( .A(n4755), .B(n4756), .Z(n23) );
  NANDN U53 ( .A(n4757), .B(n4758), .Z(n24) );
  NAND U54 ( .A(n23), .B(n24), .Z(n4776) );
  XOR U55 ( .A(n1495), .B(n1496), .Z(n1498) );
  XOR U56 ( .A(n1713), .B(n1714), .Z(n1716) );
  XOR U57 ( .A(n1786), .B(n1787), .Z(n1789) );
  XOR U58 ( .A(n2387), .B(n2388), .Z(n2390) );
  XOR U59 ( .A(n2461), .B(n2462), .Z(n2464) );
  XOR U60 ( .A(n2535), .B(n2536), .Z(n2538) );
  XOR U61 ( .A(n2746), .B(n2747), .Z(n2749) );
  NANDN U62 ( .A(n788), .B(n787), .Z(n25) );
  NANDN U63 ( .A(n789), .B(n790), .Z(n26) );
  NAND U64 ( .A(n25), .B(n26), .Z(n860) );
  NANDN U65 ( .A(n899), .B(n900), .Z(n27) );
  NANDN U66 ( .A(n898), .B(n897), .Z(n28) );
  AND U67 ( .A(n27), .B(n28), .Z(n962) );
  NANDN U68 ( .A(n1580), .B(n1579), .Z(n29) );
  NANDN U69 ( .A(n1581), .B(n1582), .Z(n30) );
  NAND U70 ( .A(n29), .B(n30), .Z(n1621) );
  OR U71 ( .A(n3744), .B(n3745), .Z(n31) );
  NANDN U72 ( .A(n3746), .B(n3747), .Z(n32) );
  NAND U73 ( .A(n31), .B(n32), .Z(n3830) );
  XOR U74 ( .A(n4457), .B(n4458), .Z(n4460) );
  XNOR U75 ( .A(n651), .B(n652), .Z(n653) );
  NANDN U76 ( .A(n868), .B(n869), .Z(n33) );
  NANDN U77 ( .A(n867), .B(n866), .Z(n34) );
  AND U78 ( .A(n33), .B(n34), .Z(n877) );
  OR U79 ( .A(n928), .B(n929), .Z(n35) );
  NANDN U80 ( .A(n931), .B(n930), .Z(n36) );
  NAND U81 ( .A(n35), .B(n36), .Z(n949) );
  OR U82 ( .A(n1403), .B(n1404), .Z(n37) );
  OR U83 ( .A(n1401), .B(n1402), .Z(n38) );
  AND U84 ( .A(n37), .B(n38), .Z(n1526) );
  NANDN U85 ( .A(n4319), .B(n4318), .Z(n39) );
  NANDN U86 ( .A(n4320), .B(n4321), .Z(n40) );
  NAND U87 ( .A(n39), .B(n40), .Z(n4372) );
  XNOR U88 ( .A(n4516), .B(n4517), .Z(n4511) );
  OR U89 ( .A(n372), .B(n373), .Z(n41) );
  NAND U90 ( .A(n375), .B(n374), .Z(n42) );
  NAND U91 ( .A(n41), .B(n42), .Z(n430) );
  NANDN U92 ( .A(n1673), .B(n1672), .Z(n43) );
  NANDN U93 ( .A(n1674), .B(n1675), .Z(n44) );
  NAND U94 ( .A(n43), .B(n44), .Z(n1682) );
  NANDN U95 ( .A(n4231), .B(n4230), .Z(n45) );
  NANDN U96 ( .A(n4232), .B(n4233), .Z(n46) );
  NAND U97 ( .A(n45), .B(n46), .Z(n4292) );
  NANDN U98 ( .A(n4551), .B(n4550), .Z(n47) );
  NANDN U99 ( .A(n4552), .B(n4553), .Z(n48) );
  NAND U100 ( .A(n47), .B(n48), .Z(n4634) );
  XOR U101 ( .A(n5062), .B(n5061), .Z(n5066) );
  NANDN U102 ( .A(n1322), .B(n1321), .Z(n49) );
  NANDN U103 ( .A(n1323), .B(n1324), .Z(n50) );
  NAND U104 ( .A(n49), .B(n50), .Z(n1396) );
  NANDN U105 ( .A(n2729), .B(n2728), .Z(n51) );
  NANDN U106 ( .A(n2730), .B(n2731), .Z(n52) );
  NAND U107 ( .A(n51), .B(n52), .Z(n2803) );
  OR U108 ( .A(n2949), .B(n2950), .Z(n53) );
  NAND U109 ( .A(n2952), .B(n2951), .Z(n54) );
  NAND U110 ( .A(n53), .B(n54), .Z(n3026) );
  OR U111 ( .A(n3325), .B(n3326), .Z(n55) );
  NAND U112 ( .A(n3328), .B(n3327), .Z(n56) );
  NAND U113 ( .A(n55), .B(n56), .Z(n3402) );
  NANDN U114 ( .A(n3625), .B(n3624), .Z(n57) );
  NANDN U115 ( .A(n3626), .B(n3627), .Z(n58) );
  NAND U116 ( .A(n57), .B(n58), .Z(n3700) );
  NANDN U117 ( .A(n3844), .B(n3843), .Z(n59) );
  NANDN U118 ( .A(n3845), .B(n3846), .Z(n60) );
  NAND U119 ( .A(n59), .B(n60), .Z(n3920) );
  OR U120 ( .A(n4214), .B(n4215), .Z(n61) );
  NAND U121 ( .A(n4217), .B(n4216), .Z(n62) );
  NAND U122 ( .A(n61), .B(n62), .Z(n4290) );
  NANDN U123 ( .A(n4777), .B(n4778), .Z(n63) );
  NANDN U124 ( .A(n4776), .B(n4775), .Z(n64) );
  AND U125 ( .A(n63), .B(n64), .Z(n4832) );
  OR U126 ( .A(n4927), .B(n4928), .Z(n65) );
  NAND U127 ( .A(n4929), .B(n4930), .Z(n66) );
  AND U128 ( .A(n65), .B(n66), .Z(n4971) );
  XOR U129 ( .A(n746), .B(n747), .Z(n792) );
  XOR U130 ( .A(n981), .B(n982), .Z(n984) );
  XOR U131 ( .A(n1051), .B(n1052), .Z(n1054) );
  XOR U132 ( .A(n1197), .B(n1198), .Z(n1200) );
  XOR U133 ( .A(n1265), .B(n1266), .Z(n1268) );
  XOR U134 ( .A(n1420), .B(n1421), .Z(n1423) );
  XNOR U135 ( .A(n1639), .B(n1640), .Z(n1641) );
  XNOR U136 ( .A(n1860), .B(n1861), .Z(n1862) );
  XOR U137 ( .A(n1935), .B(n1936), .Z(n1938) );
  XOR U138 ( .A(n2011), .B(n2012), .Z(n2014) );
  XOR U139 ( .A(n2086), .B(n2087), .Z(n2089) );
  XOR U140 ( .A(n2161), .B(n2162), .Z(n2164) );
  XOR U141 ( .A(n2236), .B(n2237), .Z(n2239) );
  XOR U142 ( .A(n2311), .B(n2312), .Z(n2314) );
  XOR U143 ( .A(n2608), .B(n2609), .Z(n2611) );
  XOR U144 ( .A(n2672), .B(n2673), .Z(n2675) );
  XNOR U145 ( .A(n2830), .B(n2831), .Z(n2832) );
  XOR U146 ( .A(n2893), .B(n2894), .Z(n2896) );
  XOR U147 ( .A(n2979), .B(n2980), .Z(n2982) );
  XOR U148 ( .A(n3043), .B(n3044), .Z(n3046) );
  XNOR U149 ( .A(n3129), .B(n3130), .Z(n3131) );
  XOR U150 ( .A(n3205), .B(n3206), .Z(n3208) );
  XOR U151 ( .A(n3281), .B(n3282), .Z(n3284) );
  XOR U152 ( .A(n3355), .B(n3356), .Z(n3358) );
  XOR U153 ( .A(n3418), .B(n3419), .Z(n3421) );
  XOR U154 ( .A(n3504), .B(n3505), .Z(n3507) );
  XOR U155 ( .A(n3568), .B(n3569), .Z(n3571) );
  XNOR U156 ( .A(n3653), .B(n3654), .Z(n3655) );
  XOR U157 ( .A(n3791), .B(n3792), .Z(n3794) );
  XNOR U158 ( .A(n3873), .B(n3874), .Z(n3875) );
  XOR U159 ( .A(n3936), .B(n3937), .Z(n3939) );
  XOR U160 ( .A(n4021), .B(n4022), .Z(n4024) );
  XOR U161 ( .A(n4097), .B(n4098), .Z(n4100) );
  NANDN U162 ( .A(n1048), .B(n1047), .Z(n67) );
  NANDN U163 ( .A(n1049), .B(n1050), .Z(n68) );
  NAND U164 ( .A(n67), .B(n68), .Z(n1108) );
  NANDN U165 ( .A(n1124), .B(n1123), .Z(n69) );
  NANDN U166 ( .A(n1125), .B(n1126), .Z(n70) );
  NAND U167 ( .A(n69), .B(n70), .Z(n1231) );
  NANDN U168 ( .A(n1194), .B(n1193), .Z(n71) );
  NANDN U169 ( .A(n1195), .B(n1196), .Z(n72) );
  NAND U170 ( .A(n71), .B(n72), .Z(n1299) );
  NANDN U171 ( .A(n1262), .B(n1261), .Z(n73) );
  NANDN U172 ( .A(n1263), .B(n1264), .Z(n74) );
  NAND U173 ( .A(n73), .B(n74), .Z(n1371) );
  NANDN U174 ( .A(n1492), .B(n1491), .Z(n75) );
  NANDN U175 ( .A(n1493), .B(n1494), .Z(n76) );
  NAND U176 ( .A(n75), .B(n76), .Z(n1594) );
  NANDN U177 ( .A(n1502), .B(n1501), .Z(n77) );
  NANDN U178 ( .A(n1503), .B(n1504), .Z(n78) );
  NAND U179 ( .A(n77), .B(n78), .Z(n1588) );
  NANDN U180 ( .A(n1710), .B(n1709), .Z(n79) );
  NANDN U181 ( .A(n1711), .B(n1712), .Z(n80) );
  NAND U182 ( .A(n79), .B(n80), .Z(n1768) );
  NANDN U183 ( .A(n1741), .B(n1740), .Z(n81) );
  NANDN U184 ( .A(n1742), .B(n1743), .Z(n82) );
  NAND U185 ( .A(n81), .B(n82), .Z(n1762) );
  NANDN U186 ( .A(n1783), .B(n1782), .Z(n83) );
  NANDN U187 ( .A(n1784), .B(n1785), .Z(n84) );
  NAND U188 ( .A(n83), .B(n84), .Z(n1841) );
  NANDN U189 ( .A(n1814), .B(n1813), .Z(n85) );
  NANDN U190 ( .A(n1815), .B(n1816), .Z(n86) );
  NAND U191 ( .A(n85), .B(n86), .Z(n1835) );
  NANDN U192 ( .A(n1857), .B(n1856), .Z(n87) );
  NANDN U193 ( .A(n1858), .B(n1859), .Z(n88) );
  NAND U194 ( .A(n87), .B(n88), .Z(n1917) );
  NANDN U195 ( .A(n1932), .B(n1931), .Z(n89) );
  NANDN U196 ( .A(n1933), .B(n1934), .Z(n90) );
  NAND U197 ( .A(n89), .B(n90), .Z(n1992) );
  NANDN U198 ( .A(n2008), .B(n2007), .Z(n91) );
  NANDN U199 ( .A(n2009), .B(n2010), .Z(n92) );
  NAND U200 ( .A(n91), .B(n92), .Z(n2068) );
  NANDN U201 ( .A(n2083), .B(n2082), .Z(n93) );
  NANDN U202 ( .A(n2084), .B(n2085), .Z(n94) );
  NAND U203 ( .A(n93), .B(n94), .Z(n2143) );
  NANDN U204 ( .A(n2158), .B(n2157), .Z(n95) );
  NANDN U205 ( .A(n2159), .B(n2160), .Z(n96) );
  NAND U206 ( .A(n95), .B(n96), .Z(n2218) );
  NANDN U207 ( .A(n2233), .B(n2232), .Z(n97) );
  NANDN U208 ( .A(n2234), .B(n2235), .Z(n98) );
  NAND U209 ( .A(n97), .B(n98), .Z(n2293) );
  NANDN U210 ( .A(n2308), .B(n2307), .Z(n99) );
  NANDN U211 ( .A(n2309), .B(n2310), .Z(n100) );
  NAND U212 ( .A(n99), .B(n100), .Z(n2368) );
  NANDN U213 ( .A(n2384), .B(n2383), .Z(n101) );
  NANDN U214 ( .A(n2385), .B(n2386), .Z(n102) );
  NAND U215 ( .A(n101), .B(n102), .Z(n2442) );
  NANDN U216 ( .A(n2415), .B(n2414), .Z(n103) );
  NANDN U217 ( .A(n2416), .B(n2417), .Z(n104) );
  NAND U218 ( .A(n103), .B(n104), .Z(n2436) );
  NANDN U219 ( .A(n2458), .B(n2457), .Z(n105) );
  NANDN U220 ( .A(n2459), .B(n2460), .Z(n106) );
  NAND U221 ( .A(n105), .B(n106), .Z(n2516) );
  NANDN U222 ( .A(n2489), .B(n2488), .Z(n107) );
  NANDN U223 ( .A(n2490), .B(n2491), .Z(n108) );
  NAND U224 ( .A(n107), .B(n108), .Z(n2510) );
  NANDN U225 ( .A(n2532), .B(n2531), .Z(n109) );
  NANDN U226 ( .A(n2533), .B(n2534), .Z(n110) );
  NAND U227 ( .A(n109), .B(n110), .Z(n2590) );
  NANDN U228 ( .A(n2564), .B(n2565), .Z(n111) );
  NANDN U229 ( .A(n2563), .B(n2562), .Z(n112) );
  AND U230 ( .A(n111), .B(n112), .Z(n2583) );
  NANDN U231 ( .A(n2605), .B(n2604), .Z(n113) );
  NANDN U232 ( .A(n2606), .B(n2607), .Z(n114) );
  NAND U233 ( .A(n113), .B(n114), .Z(n2712) );
  NANDN U234 ( .A(n2669), .B(n2668), .Z(n115) );
  NANDN U235 ( .A(n2670), .B(n2671), .Z(n116) );
  NAND U236 ( .A(n115), .B(n116), .Z(n2778) );
  OR U237 ( .A(n2773), .B(n2774), .Z(n117) );
  NAND U238 ( .A(n2775), .B(n2776), .Z(n118) );
  AND U239 ( .A(n117), .B(n118), .Z(n2810) );
  NANDN U240 ( .A(n2743), .B(n2742), .Z(n119) );
  NANDN U241 ( .A(n2744), .B(n2745), .Z(n120) );
  NAND U242 ( .A(n119), .B(n120), .Z(n2805) );
  NANDN U243 ( .A(n2827), .B(n2826), .Z(n121) );
  NANDN U244 ( .A(n2828), .B(n2829), .Z(n122) );
  NAND U245 ( .A(n121), .B(n122), .Z(n2933) );
  NANDN U246 ( .A(n2890), .B(n2889), .Z(n123) );
  NANDN U247 ( .A(n2891), .B(n2892), .Z(n124) );
  NAND U248 ( .A(n123), .B(n124), .Z(n2960) );
  NANDN U249 ( .A(n2976), .B(n2975), .Z(n125) );
  NANDN U250 ( .A(n2977), .B(n2978), .Z(n126) );
  NAND U251 ( .A(n125), .B(n126), .Z(n3083) );
  NANDN U252 ( .A(n3040), .B(n3039), .Z(n127) );
  NANDN U253 ( .A(n3041), .B(n3042), .Z(n128) );
  NAND U254 ( .A(n127), .B(n128), .Z(n3104) );
  NANDN U255 ( .A(n3126), .B(n3125), .Z(n129) );
  NANDN U256 ( .A(n3127), .B(n3128), .Z(n130) );
  NAND U257 ( .A(n129), .B(n130), .Z(n3186) );
  NANDN U258 ( .A(n3202), .B(n3201), .Z(n131) );
  NANDN U259 ( .A(n3203), .B(n3204), .Z(n132) );
  NAND U260 ( .A(n131), .B(n132), .Z(n3262) );
  NANDN U261 ( .A(n3278), .B(n3277), .Z(n133) );
  NANDN U262 ( .A(n3279), .B(n3280), .Z(n134) );
  NAND U263 ( .A(n133), .B(n134), .Z(n3336) );
  NANDN U264 ( .A(n3352), .B(n3351), .Z(n135) );
  NANDN U265 ( .A(n3353), .B(n3354), .Z(n136) );
  NAND U266 ( .A(n135), .B(n136), .Z(n3458) );
  NANDN U267 ( .A(n3415), .B(n3414), .Z(n137) );
  NANDN U268 ( .A(n3416), .B(n3417), .Z(n138) );
  NAND U269 ( .A(n137), .B(n138), .Z(n3479) );
  NANDN U270 ( .A(n3501), .B(n3500), .Z(n139) );
  NANDN U271 ( .A(n3502), .B(n3503), .Z(n140) );
  NAND U272 ( .A(n139), .B(n140), .Z(n3608) );
  NANDN U273 ( .A(n3565), .B(n3564), .Z(n141) );
  NANDN U274 ( .A(n3566), .B(n3567), .Z(n142) );
  NAND U275 ( .A(n141), .B(n142), .Z(n3629) );
  NANDN U276 ( .A(n3650), .B(n3649), .Z(n143) );
  NANDN U277 ( .A(n3651), .B(n3652), .Z(n144) );
  NAND U278 ( .A(n143), .B(n144), .Z(n3755) );
  NANDN U279 ( .A(n3870), .B(n3869), .Z(n145) );
  NANDN U280 ( .A(n3871), .B(n3872), .Z(n146) );
  NAND U281 ( .A(n145), .B(n146), .Z(n3976) );
  NANDN U282 ( .A(n3933), .B(n3932), .Z(n147) );
  NANDN U283 ( .A(n3934), .B(n3935), .Z(n148) );
  NAND U284 ( .A(n147), .B(n148), .Z(n4003) );
  NANDN U285 ( .A(n4018), .B(n4017), .Z(n149) );
  NANDN U286 ( .A(n4019), .B(n4020), .Z(n150) );
  NAND U287 ( .A(n149), .B(n150), .Z(n4078) );
  NANDN U288 ( .A(n4094), .B(n4093), .Z(n151) );
  NANDN U289 ( .A(n4095), .B(n4096), .Z(n152) );
  NAND U290 ( .A(n151), .B(n152), .Z(n4154) );
  XOR U291 ( .A(n4255), .B(n4256), .Z(n4258) );
  OR U292 ( .A(b[0]), .B(n5094), .Z(n153) );
  AND U293 ( .A(b[1]), .B(n153), .Z(n4494) );
  NANDN U294 ( .A(n1398), .B(n1397), .Z(n154) );
  NANDN U295 ( .A(n1399), .B(n1400), .Z(n155) );
  NAND U296 ( .A(n154), .B(n155), .Z(n1527) );
  OR U297 ( .A(n1622), .B(n1623), .Z(n156) );
  OR U298 ( .A(n1620), .B(n1621), .Z(n157) );
  AND U299 ( .A(n156), .B(n157), .Z(n1744) );
  NANDN U300 ( .A(n3825), .B(n3824), .Z(n158) );
  NANDN U301 ( .A(n3826), .B(n3827), .Z(n159) );
  NAND U302 ( .A(n158), .B(n159), .Z(n3907) );
  NANDN U303 ( .A(n4175), .B(n4174), .Z(n160) );
  NANDN U304 ( .A(n4172), .B(n4173), .Z(n161) );
  NAND U305 ( .A(n160), .B(n161), .Z(n4226) );
  XOR U306 ( .A(n4398), .B(n4399), .Z(n4401) );
  NANDN U307 ( .A(n648), .B(n647), .Z(n162) );
  NANDN U308 ( .A(n649), .B(n650), .Z(n163) );
  NAND U309 ( .A(n162), .B(n163), .Z(n720) );
  NANDN U310 ( .A(n950), .B(n949), .Z(n164) );
  NANDN U311 ( .A(n951), .B(n952), .Z(n165) );
  NAND U312 ( .A(n164), .B(n165), .Z(n1019) );
  NANDN U313 ( .A(n4385), .B(n4384), .Z(n166) );
  NANDN U314 ( .A(n4386), .B(n4387), .Z(n167) );
  NAND U315 ( .A(n166), .B(n167), .Z(n4452) );
  OR U316 ( .A(n4562), .B(n4563), .Z(n168) );
  NANDN U317 ( .A(n4560), .B(n4561), .Z(n169) );
  AND U318 ( .A(n168), .B(n169), .Z(n4639) );
  XOR U319 ( .A(n4635), .B(n4636), .Z(n4630) );
  OR U320 ( .A(n4677), .B(n4678), .Z(n170) );
  NANDN U321 ( .A(n4675), .B(n4676), .Z(n171) );
  NAND U322 ( .A(n170), .B(n171), .Z(n4755) );
  NANDN U323 ( .A(n4873), .B(n4872), .Z(n172) );
  NANDN U324 ( .A(n4874), .B(n4875), .Z(n173) );
  NAND U325 ( .A(n172), .B(n173), .Z(n4891) );
  NANDN U326 ( .A(n5030), .B(n5062), .Z(n174) );
  NANDN U327 ( .A(n5031), .B(n5032), .Z(n175) );
  NAND U328 ( .A(n174), .B(n175), .Z(n5071) );
  OR U329 ( .A(n280), .B(n281), .Z(n176) );
  NANDN U330 ( .A(n283), .B(n282), .Z(n177) );
  AND U331 ( .A(n176), .B(n177), .Z(n292) );
  NANDN U332 ( .A(n814), .B(n813), .Z(n178) );
  NANDN U333 ( .A(n815), .B(n816), .Z(n179) );
  NAND U334 ( .A(n178), .B(n179), .Z(n870) );
  NANDN U335 ( .A(n1394), .B(n1393), .Z(n180) );
  NANDN U336 ( .A(n1395), .B(n1396), .Z(n181) );
  NAND U337 ( .A(n180), .B(n181), .Z(n1467) );
  NANDN U338 ( .A(n1611), .B(n1610), .Z(n182) );
  NANDN U339 ( .A(n1612), .B(n1613), .Z(n183) );
  NAND U340 ( .A(n182), .B(n183), .Z(n1684) );
  NANDN U341 ( .A(n2801), .B(n2800), .Z(n184) );
  NANDN U342 ( .A(n2802), .B(n2803), .Z(n185) );
  NAND U343 ( .A(n184), .B(n185), .Z(n2877) );
  NANDN U344 ( .A(n3100), .B(n3099), .Z(n186) );
  NANDN U345 ( .A(n3101), .B(n3102), .Z(n187) );
  NAND U346 ( .A(n186), .B(n187), .Z(n3176) );
  NANDN U347 ( .A(n3475), .B(n3474), .Z(n188) );
  NANDN U348 ( .A(n3476), .B(n3477), .Z(n189) );
  NAND U349 ( .A(n188), .B(n189), .Z(n3551) );
  NANDN U350 ( .A(n3772), .B(n3771), .Z(n190) );
  NANDN U351 ( .A(n3773), .B(n3774), .Z(n191) );
  NAND U352 ( .A(n190), .B(n191), .Z(n3846) );
  OR U353 ( .A(n3992), .B(n3993), .Z(n192) );
  NAND U354 ( .A(n3995), .B(n3994), .Z(n193) );
  NAND U355 ( .A(n192), .B(n193), .Z(n4068) );
  NANDN U356 ( .A(n4288), .B(n4287), .Z(n194) );
  NANDN U357 ( .A(n4289), .B(n4290), .Z(n195) );
  NAND U358 ( .A(n194), .B(n195), .Z(n4363) );
  OR U359 ( .A(n4443), .B(n4444), .Z(n196) );
  NANDN U360 ( .A(n4441), .B(n4442), .Z(n197) );
  NAND U361 ( .A(n196), .B(n197), .Z(n4504) );
  NANDN U362 ( .A(n444), .B(n443), .Z(n198) );
  NANDN U363 ( .A(n445), .B(n446), .Z(n199) );
  NAND U364 ( .A(n198), .B(n199), .Z(n485) );
  NAND U365 ( .A(n4833), .B(n4831), .Z(n200) );
  XOR U366 ( .A(n4831), .B(n4833), .Z(n201) );
  NANDN U367 ( .A(n4832), .B(n201), .Z(n202) );
  NAND U368 ( .A(n200), .B(n202), .Z(n4880) );
  NAND U369 ( .A(n4971), .B(n4972), .Z(n203) );
  XOR U370 ( .A(n4972), .B(n4971), .Z(n204) );
  NANDN U371 ( .A(n4973), .B(n204), .Z(n205) );
  NAND U372 ( .A(n203), .B(n205), .Z(n5014) );
  IV U373 ( .A(b[0]), .Z(n206) );
  IV U374 ( .A(b[1]), .Z(n207) );
  IV U375 ( .A(b[3]), .Z(n208) );
  IV U376 ( .A(b[5]), .Z(n209) );
  IV U377 ( .A(b[15]), .Z(n210) );
  NAND U378 ( .A(b[0]), .B(a[0]), .Z(n212) );
  XNOR U379 ( .A(n212), .B(sreg[48]), .Z(c[48]) );
  NAND U380 ( .A(b[0]), .B(a[1]), .Z(n217) );
  NAND U381 ( .A(b[1]), .B(a[0]), .Z(n211) );
  XOR U382 ( .A(n217), .B(n211), .Z(n220) );
  XNOR U383 ( .A(sreg[49]), .B(n220), .Z(n222) );
  NANDN U384 ( .A(n212), .B(sreg[48]), .Z(n221) );
  XOR U385 ( .A(n222), .B(n221), .Z(c[49]) );
  NAND U386 ( .A(b[0]), .B(a[2]), .Z(n213) );
  XNOR U387 ( .A(b[1]), .B(n213), .Z(n215) );
  NAND U388 ( .A(a[1]), .B(n206), .Z(n214) );
  AND U389 ( .A(n215), .B(n214), .Z(n226) );
  NAND U390 ( .A(a[0]), .B(b[2]), .Z(n216) );
  XNOR U391 ( .A(b[1]), .B(n216), .Z(n219) );
  IV U392 ( .A(a[0]), .Z(n760) );
  NANDN U393 ( .A(n217), .B(n760), .Z(n218) );
  AND U394 ( .A(n219), .B(n218), .Z(n225) );
  XNOR U395 ( .A(n226), .B(n225), .Z(n238) );
  NAND U396 ( .A(n220), .B(sreg[49]), .Z(n224) );
  OR U397 ( .A(n222), .B(n221), .Z(n223) );
  NAND U398 ( .A(n224), .B(n223), .Z(n236) );
  XNOR U399 ( .A(n236), .B(sreg[50]), .Z(n237) );
  XOR U400 ( .A(n238), .B(n237), .Z(c[50]) );
  NAND U401 ( .A(n226), .B(n225), .Z(n249) );
  XOR U402 ( .A(n207), .B(b[2]), .Z(n4488) );
  NOR U403 ( .A(n208), .B(n4488), .Z(n4523) );
  NAND U404 ( .A(n760), .B(n4523), .Z(n228) );
  NOR U405 ( .A(n208), .B(b[2]), .Z(n4606) );
  NAND U406 ( .A(n207), .B(n4606), .Z(n227) );
  NAND U407 ( .A(n228), .B(n227), .Z(n247) );
  XOR U408 ( .A(b[3]), .B(b[2]), .Z(n258) );
  XOR U409 ( .A(b[3]), .B(a[0]), .Z(n229) );
  NAND U410 ( .A(n258), .B(n229), .Z(n230) );
  XNOR U411 ( .A(n208), .B(n207), .Z(n257) );
  OR U412 ( .A(n230), .B(n257), .Z(n232) );
  IV U413 ( .A(a[1]), .Z(n770) );
  XNOR U414 ( .A(n208), .B(n770), .Z(n259) );
  OR U415 ( .A(n259), .B(n4488), .Z(n231) );
  NAND U416 ( .A(n232), .B(n231), .Z(n253) );
  NAND U417 ( .A(b[0]), .B(a[3]), .Z(n233) );
  XNOR U418 ( .A(b[1]), .B(n233), .Z(n235) );
  NAND U419 ( .A(a[2]), .B(n206), .Z(n234) );
  AND U420 ( .A(n235), .B(n234), .Z(n252) );
  XOR U421 ( .A(n253), .B(n252), .Z(n246) );
  XOR U422 ( .A(n247), .B(n246), .Z(n248) );
  XNOR U423 ( .A(n249), .B(n248), .Z(n241) );
  XNOR U424 ( .A(sreg[51]), .B(n241), .Z(n243) );
  NAND U425 ( .A(n236), .B(sreg[50]), .Z(n240) );
  OR U426 ( .A(n238), .B(n237), .Z(n239) );
  AND U427 ( .A(n240), .B(n239), .Z(n242) );
  XOR U428 ( .A(n243), .B(n242), .Z(c[51]) );
  NAND U429 ( .A(sreg[51]), .B(n241), .Z(n245) );
  OR U430 ( .A(n243), .B(n242), .Z(n244) );
  NAND U431 ( .A(n245), .B(n244), .Z(n284) );
  XNOR U432 ( .A(n284), .B(sreg[52]), .Z(n286) );
  NAND U433 ( .A(n247), .B(n246), .Z(n251) );
  NANDN U434 ( .A(n249), .B(n248), .Z(n250) );
  NAND U435 ( .A(n251), .B(n250), .Z(n283) );
  AND U436 ( .A(n253), .B(n252), .Z(n280) );
  XOR U437 ( .A(b[4]), .B(n208), .Z(n4612) );
  OR U438 ( .A(n4612), .B(n760), .Z(n277) );
  NAND U439 ( .A(b[0]), .B(a[4]), .Z(n254) );
  XNOR U440 ( .A(b[1]), .B(n254), .Z(n256) );
  NAND U441 ( .A(n206), .B(a[3]), .Z(n255) );
  AND U442 ( .A(n256), .B(n255), .Z(n275) );
  ANDN U443 ( .B(n258), .A(n257), .Z(n4521) );
  NANDN U444 ( .A(n259), .B(n4521), .Z(n261) );
  IV U445 ( .A(a[2]), .Z(n839) );
  XNOR U446 ( .A(n208), .B(n839), .Z(n271) );
  OR U447 ( .A(n271), .B(n4488), .Z(n260) );
  AND U448 ( .A(n261), .B(n260), .Z(n274) );
  XNOR U449 ( .A(n275), .B(n274), .Z(n276) );
  XNOR U450 ( .A(n277), .B(n276), .Z(n281) );
  XOR U451 ( .A(n280), .B(n281), .Z(n282) );
  XNOR U452 ( .A(n283), .B(n282), .Z(n285) );
  XOR U453 ( .A(n286), .B(n285), .Z(c[52]) );
  NAND U454 ( .A(b[0]), .B(a[5]), .Z(n262) );
  XNOR U455 ( .A(b[1]), .B(n262), .Z(n264) );
  NAND U456 ( .A(a[4]), .B(n206), .Z(n263) );
  AND U457 ( .A(n264), .B(n263), .Z(n295) );
  XNOR U458 ( .A(b[5]), .B(n770), .Z(n303) );
  NANDN U459 ( .A(n4612), .B(n303), .Z(n268) );
  XOR U460 ( .A(b[5]), .B(a[0]), .Z(n342) );
  XNOR U461 ( .A(n209), .B(b[4]), .Z(n266) );
  XOR U462 ( .A(b[5]), .B(b[3]), .Z(n265) );
  AND U463 ( .A(n266), .B(n265), .Z(n4669) );
  NAND U464 ( .A(n342), .B(n4669), .Z(n267) );
  NAND U465 ( .A(n268), .B(n267), .Z(n296) );
  XNOR U466 ( .A(n295), .B(n296), .Z(n309) );
  ANDN U467 ( .B(b[5]), .A(b[4]), .Z(n4751) );
  NAND U468 ( .A(n208), .B(n4751), .Z(n270) );
  NOR U469 ( .A(n209), .B(n4612), .Z(n4750) );
  NAND U470 ( .A(n760), .B(n4750), .Z(n269) );
  NAND U471 ( .A(n270), .B(n269), .Z(n307) );
  NANDN U472 ( .A(n271), .B(n4521), .Z(n273) );
  XOR U473 ( .A(b[3]), .B(a[3]), .Z(n297) );
  NANDN U474 ( .A(n4488), .B(n297), .Z(n272) );
  AND U475 ( .A(n273), .B(n272), .Z(n306) );
  XNOR U476 ( .A(n307), .B(n306), .Z(n308) );
  XOR U477 ( .A(n309), .B(n308), .Z(n289) );
  NANDN U478 ( .A(n275), .B(n274), .Z(n279) );
  NAND U479 ( .A(n277), .B(n276), .Z(n278) );
  NAND U480 ( .A(n279), .B(n278), .Z(n290) );
  XOR U481 ( .A(n289), .B(n290), .Z(n291) );
  XOR U482 ( .A(n291), .B(n292), .Z(n312) );
  XNOR U483 ( .A(sreg[53]), .B(n312), .Z(n314) );
  NAND U484 ( .A(n284), .B(sreg[52]), .Z(n288) );
  OR U485 ( .A(n286), .B(n285), .Z(n287) );
  AND U486 ( .A(n288), .B(n287), .Z(n313) );
  XOR U487 ( .A(n314), .B(n313), .Z(c[53]) );
  OR U488 ( .A(n290), .B(n289), .Z(n294) );
  NAND U489 ( .A(n292), .B(n291), .Z(n293) );
  NAND U490 ( .A(n294), .B(n293), .Z(n320) );
  AND U491 ( .A(n296), .B(n295), .Z(n326) );
  NAND U492 ( .A(n297), .B(n4521), .Z(n299) );
  XOR U493 ( .A(b[3]), .B(a[4]), .Z(n334) );
  NANDN U494 ( .A(n4488), .B(n334), .Z(n298) );
  NAND U495 ( .A(n299), .B(n298), .Z(n331) );
  XOR U496 ( .A(n209), .B(b[6]), .Z(n343) );
  ANDN U497 ( .B(a[0]), .A(n343), .Z(n346) );
  NAND U498 ( .A(b[0]), .B(a[6]), .Z(n300) );
  XNOR U499 ( .A(b[1]), .B(n300), .Z(n302) );
  NAND U500 ( .A(a[5]), .B(n206), .Z(n301) );
  AND U501 ( .A(n302), .B(n301), .Z(n329) );
  XOR U502 ( .A(n346), .B(n329), .Z(n330) );
  XNOR U503 ( .A(n331), .B(n330), .Z(n323) );
  NAND U504 ( .A(n4669), .B(n303), .Z(n305) );
  XOR U505 ( .A(b[5]), .B(a[2]), .Z(n337) );
  NANDN U506 ( .A(n4612), .B(n337), .Z(n304) );
  NAND U507 ( .A(n305), .B(n304), .Z(n324) );
  XNOR U508 ( .A(n323), .B(n324), .Z(n325) );
  XOR U509 ( .A(n326), .B(n325), .Z(n317) );
  NANDN U510 ( .A(n307), .B(n306), .Z(n311) );
  NAND U511 ( .A(n309), .B(n308), .Z(n310) );
  NAND U512 ( .A(n311), .B(n310), .Z(n318) );
  XNOR U513 ( .A(n317), .B(n318), .Z(n319) );
  XNOR U514 ( .A(n320), .B(n319), .Z(n352) );
  NAND U515 ( .A(sreg[53]), .B(n312), .Z(n316) );
  OR U516 ( .A(n314), .B(n313), .Z(n315) );
  NAND U517 ( .A(n316), .B(n315), .Z(n350) );
  XNOR U518 ( .A(n350), .B(sreg[54]), .Z(n351) );
  XOR U519 ( .A(n352), .B(n351), .Z(c[54]) );
  NANDN U520 ( .A(n318), .B(n317), .Z(n322) );
  NAND U521 ( .A(n320), .B(n319), .Z(n321) );
  NAND U522 ( .A(n322), .B(n321), .Z(n363) );
  NANDN U523 ( .A(n324), .B(n323), .Z(n328) );
  NANDN U524 ( .A(n326), .B(n325), .Z(n327) );
  NAND U525 ( .A(n328), .B(n327), .Z(n361) );
  NAND U526 ( .A(n346), .B(n329), .Z(n333) );
  NAND U527 ( .A(n331), .B(n330), .Z(n332) );
  NAND U528 ( .A(n333), .B(n332), .Z(n367) );
  NAND U529 ( .A(n334), .B(n4521), .Z(n336) );
  XOR U530 ( .A(b[3]), .B(a[5]), .Z(n379) );
  NANDN U531 ( .A(n4488), .B(n379), .Z(n335) );
  AND U532 ( .A(n336), .B(n335), .Z(n366) );
  XNOR U533 ( .A(n367), .B(n366), .Z(n368) );
  XOR U534 ( .A(b[5]), .B(a[3]), .Z(n387) );
  NANDN U535 ( .A(n4612), .B(n387), .Z(n339) );
  NAND U536 ( .A(n337), .B(n4669), .Z(n338) );
  NAND U537 ( .A(n339), .B(n338), .Z(n383) );
  XOR U538 ( .A(b[7]), .B(b[5]), .Z(n341) );
  XOR U539 ( .A(b[7]), .B(b[6]), .Z(n340) );
  AND U540 ( .A(n341), .B(n340), .Z(n4746) );
  NANDN U541 ( .A(n342), .B(n4746), .Z(n345) );
  IV U542 ( .A(b[7]), .Z(n4744) );
  XNOR U543 ( .A(n4744), .B(n770), .Z(n376) );
  IV U544 ( .A(n343), .Z(n4745) );
  NANDN U545 ( .A(n376), .B(n4745), .Z(n344) );
  NAND U546 ( .A(n345), .B(n344), .Z(n382) );
  XNOR U547 ( .A(n383), .B(n382), .Z(n375) );
  NAND U548 ( .A(b[5]), .B(b[6]), .Z(n4812) );
  ANDN U549 ( .B(n4812), .A(n4744), .Z(n4903) );
  ANDN U550 ( .B(n4903), .A(n346), .Z(n372) );
  NAND U551 ( .A(b[0]), .B(a[7]), .Z(n347) );
  XNOR U552 ( .A(b[1]), .B(n347), .Z(n349) );
  NAND U553 ( .A(a[6]), .B(n206), .Z(n348) );
  AND U554 ( .A(n349), .B(n348), .Z(n373) );
  XOR U555 ( .A(n372), .B(n373), .Z(n374) );
  XOR U556 ( .A(n375), .B(n374), .Z(n369) );
  XOR U557 ( .A(n368), .B(n369), .Z(n360) );
  XNOR U558 ( .A(n361), .B(n360), .Z(n362) );
  XNOR U559 ( .A(n363), .B(n362), .Z(n355) );
  XNOR U560 ( .A(n355), .B(sreg[55]), .Z(n357) );
  NAND U561 ( .A(n350), .B(sreg[54]), .Z(n354) );
  OR U562 ( .A(n352), .B(n351), .Z(n353) );
  AND U563 ( .A(n354), .B(n353), .Z(n356) );
  XOR U564 ( .A(n357), .B(n356), .Z(c[55]) );
  NAND U565 ( .A(n355), .B(sreg[55]), .Z(n359) );
  OR U566 ( .A(n357), .B(n356), .Z(n358) );
  NAND U567 ( .A(n359), .B(n358), .Z(n433) );
  XNOR U568 ( .A(n433), .B(sreg[56]), .Z(n435) );
  NAND U569 ( .A(n361), .B(n360), .Z(n365) );
  OR U570 ( .A(n363), .B(n362), .Z(n364) );
  NAND U571 ( .A(n365), .B(n364), .Z(n393) );
  NANDN U572 ( .A(n367), .B(n366), .Z(n371) );
  NAND U573 ( .A(n369), .B(n368), .Z(n370) );
  NAND U574 ( .A(n371), .B(n370), .Z(n390) );
  XNOR U575 ( .A(n4744), .B(n839), .Z(n408) );
  NANDN U576 ( .A(n408), .B(n4745), .Z(n378) );
  NANDN U577 ( .A(n376), .B(n4746), .Z(n377) );
  NAND U578 ( .A(n378), .B(n377), .Z(n396) );
  NAND U579 ( .A(n379), .B(n4521), .Z(n381) );
  IV U580 ( .A(a[6]), .Z(n1119) );
  XNOR U581 ( .A(n208), .B(n1119), .Z(n405) );
  OR U582 ( .A(n405), .B(n4488), .Z(n380) );
  AND U583 ( .A(n381), .B(n380), .Z(n397) );
  XNOR U584 ( .A(n396), .B(n397), .Z(n398) );
  NAND U585 ( .A(n383), .B(n382), .Z(n399) );
  XOR U586 ( .A(n398), .B(n399), .Z(n427) );
  XOR U587 ( .A(b[8]), .B(n4744), .Z(n4860) );
  OR U588 ( .A(n4860), .B(n760), .Z(n424) );
  AND U589 ( .A(a[8]), .B(b[0]), .Z(n384) );
  XOR U590 ( .A(b[1]), .B(n384), .Z(n386) );
  NAND U591 ( .A(a[7]), .B(n206), .Z(n385) );
  NAND U592 ( .A(n386), .B(n385), .Z(n421) );
  NAND U593 ( .A(n4669), .B(n387), .Z(n389) );
  XOR U594 ( .A(b[5]), .B(a[4]), .Z(n418) );
  NANDN U595 ( .A(n4612), .B(n418), .Z(n388) );
  NAND U596 ( .A(n389), .B(n388), .Z(n422) );
  XNOR U597 ( .A(n421), .B(n422), .Z(n423) );
  XNOR U598 ( .A(n424), .B(n423), .Z(n428) );
  XNOR U599 ( .A(n427), .B(n428), .Z(n429) );
  XNOR U600 ( .A(n430), .B(n429), .Z(n391) );
  XNOR U601 ( .A(n390), .B(n391), .Z(n392) );
  XOR U602 ( .A(n393), .B(n392), .Z(n434) );
  XOR U603 ( .A(n435), .B(n434), .Z(c[56]) );
  NANDN U604 ( .A(n391), .B(n390), .Z(n395) );
  NAND U605 ( .A(n393), .B(n392), .Z(n394) );
  NAND U606 ( .A(n395), .B(n394), .Z(n446) );
  NANDN U607 ( .A(n397), .B(n396), .Z(n401) );
  NANDN U608 ( .A(n399), .B(n398), .Z(n400) );
  NAND U609 ( .A(n401), .B(n400), .Z(n450) );
  NAND U610 ( .A(b[0]), .B(a[9]), .Z(n402) );
  XNOR U611 ( .A(b[1]), .B(n402), .Z(n404) );
  NAND U612 ( .A(a[8]), .B(n206), .Z(n403) );
  AND U613 ( .A(n404), .B(n403), .Z(n460) );
  NANDN U614 ( .A(n405), .B(n4521), .Z(n407) );
  IV U615 ( .A(a[7]), .Z(n1189) );
  XNOR U616 ( .A(n208), .B(n1189), .Z(n473) );
  OR U617 ( .A(n473), .B(n4488), .Z(n406) );
  AND U618 ( .A(n407), .B(n406), .Z(n459) );
  XNOR U619 ( .A(n460), .B(n459), .Z(n461) );
  XOR U620 ( .A(b[7]), .B(a[3]), .Z(n479) );
  NAND U621 ( .A(n4745), .B(n479), .Z(n410) );
  NANDN U622 ( .A(n408), .B(n4746), .Z(n409) );
  NAND U623 ( .A(n410), .B(n409), .Z(n465) );
  XOR U624 ( .A(b[9]), .B(a[0]), .Z(n413) );
  IV U625 ( .A(b[9]), .Z(n4859) );
  XNOR U626 ( .A(n4859), .B(b[8]), .Z(n412) );
  XOR U627 ( .A(b[9]), .B(b[7]), .Z(n411) );
  AND U628 ( .A(n412), .B(n411), .Z(n4915) );
  NAND U629 ( .A(n413), .B(n4915), .Z(n415) );
  XNOR U630 ( .A(b[9]), .B(n770), .Z(n467) );
  ANDN U631 ( .B(n467), .A(n4860), .Z(n414) );
  ANDN U632 ( .B(n415), .A(n414), .Z(n466) );
  XNOR U633 ( .A(n465), .B(n466), .Z(n456) );
  ANDN U634 ( .B(b[9]), .A(b[8]), .Z(n4957) );
  NAND U635 ( .A(n4744), .B(n4957), .Z(n417) );
  NOR U636 ( .A(n4859), .B(n4860), .Z(n4956) );
  NAND U637 ( .A(n760), .B(n4956), .Z(n416) );
  NAND U638 ( .A(n417), .B(n416), .Z(n454) );
  IV U639 ( .A(a[5]), .Z(n1043) );
  XNOR U640 ( .A(b[5]), .B(n1043), .Z(n470) );
  NANDN U641 ( .A(n4612), .B(n470), .Z(n420) );
  NAND U642 ( .A(n418), .B(n4669), .Z(n419) );
  NAND U643 ( .A(n420), .B(n419), .Z(n453) );
  XOR U644 ( .A(n454), .B(n453), .Z(n455) );
  XOR U645 ( .A(n456), .B(n455), .Z(n462) );
  XOR U646 ( .A(n461), .B(n462), .Z(n447) );
  NANDN U647 ( .A(n422), .B(n421), .Z(n426) );
  NAND U648 ( .A(n424), .B(n423), .Z(n425) );
  NAND U649 ( .A(n426), .B(n425), .Z(n448) );
  XNOR U650 ( .A(n447), .B(n448), .Z(n449) );
  XNOR U651 ( .A(n450), .B(n449), .Z(n443) );
  NANDN U652 ( .A(n428), .B(n427), .Z(n432) );
  NAND U653 ( .A(n430), .B(n429), .Z(n431) );
  AND U654 ( .A(n432), .B(n431), .Z(n444) );
  XOR U655 ( .A(n443), .B(n444), .Z(n445) );
  XOR U656 ( .A(n446), .B(n445), .Z(n438) );
  XNOR U657 ( .A(n438), .B(sreg[57]), .Z(n440) );
  NAND U658 ( .A(n433), .B(sreg[56]), .Z(n437) );
  OR U659 ( .A(n435), .B(n434), .Z(n436) );
  AND U660 ( .A(n437), .B(n436), .Z(n439) );
  XOR U661 ( .A(n440), .B(n439), .Z(c[57]) );
  NAND U662 ( .A(n438), .B(sreg[57]), .Z(n442) );
  OR U663 ( .A(n440), .B(n439), .Z(n441) );
  NAND U664 ( .A(n442), .B(n441), .Z(n536) );
  XNOR U665 ( .A(n536), .B(sreg[58]), .Z(n538) );
  NANDN U666 ( .A(n448), .B(n447), .Z(n452) );
  NAND U667 ( .A(n450), .B(n449), .Z(n451) );
  NAND U668 ( .A(n452), .B(n451), .Z(n483) );
  OR U669 ( .A(n454), .B(n453), .Z(n458) );
  NANDN U670 ( .A(n456), .B(n455), .Z(n457) );
  NAND U671 ( .A(n458), .B(n457), .Z(n490) );
  NANDN U672 ( .A(n460), .B(n459), .Z(n464) );
  NANDN U673 ( .A(n462), .B(n461), .Z(n463) );
  NAND U674 ( .A(n464), .B(n463), .Z(n489) );
  NANDN U675 ( .A(n466), .B(n465), .Z(n509) );
  NAND U676 ( .A(n4915), .B(n467), .Z(n469) );
  XOR U677 ( .A(b[9]), .B(a[2]), .Z(n522) );
  NANDN U678 ( .A(n4860), .B(n522), .Z(n468) );
  NAND U679 ( .A(n469), .B(n468), .Z(n507) );
  NAND U680 ( .A(n4669), .B(n470), .Z(n472) );
  XNOR U681 ( .A(b[5]), .B(n1119), .Z(n533) );
  NANDN U682 ( .A(n4612), .B(n533), .Z(n471) );
  AND U683 ( .A(n472), .B(n471), .Z(n506) );
  XNOR U684 ( .A(n507), .B(n506), .Z(n508) );
  XNOR U685 ( .A(n509), .B(n508), .Z(n495) );
  NANDN U686 ( .A(n473), .B(n4521), .Z(n475) );
  XOR U687 ( .A(b[3]), .B(a[8]), .Z(n519) );
  NANDN U688 ( .A(n4488), .B(n519), .Z(n474) );
  AND U689 ( .A(n475), .B(n474), .Z(n494) );
  XNOR U690 ( .A(n495), .B(n494), .Z(n496) );
  IV U691 ( .A(b[10]), .Z(n5033) );
  XNOR U692 ( .A(n5033), .B(n4859), .Z(n4986) );
  ANDN U693 ( .B(a[0]), .A(n4986), .Z(n503) );
  NAND U694 ( .A(b[0]), .B(a[10]), .Z(n476) );
  XNOR U695 ( .A(b[1]), .B(n476), .Z(n478) );
  NAND U696 ( .A(a[9]), .B(n206), .Z(n477) );
  AND U697 ( .A(n478), .B(n477), .Z(n501) );
  IV U698 ( .A(a[4]), .Z(n971) );
  XNOR U699 ( .A(n4744), .B(n971), .Z(n512) );
  NANDN U700 ( .A(n512), .B(n4745), .Z(n481) );
  NAND U701 ( .A(n479), .B(n4746), .Z(n480) );
  AND U702 ( .A(n481), .B(n480), .Z(n500) );
  XNOR U703 ( .A(n501), .B(n500), .Z(n502) );
  XOR U704 ( .A(n503), .B(n502), .Z(n497) );
  XNOR U705 ( .A(n496), .B(n497), .Z(n488) );
  XNOR U706 ( .A(n489), .B(n488), .Z(n491) );
  XNOR U707 ( .A(n490), .B(n491), .Z(n482) );
  XNOR U708 ( .A(n483), .B(n482), .Z(n484) );
  XOR U709 ( .A(n485), .B(n484), .Z(n537) );
  XOR U710 ( .A(n538), .B(n537), .Z(c[58]) );
  NANDN U711 ( .A(n483), .B(n482), .Z(n487) );
  NAND U712 ( .A(n485), .B(n484), .Z(n486) );
  NAND U713 ( .A(n487), .B(n486), .Z(n549) );
  NAND U714 ( .A(n489), .B(n488), .Z(n493) );
  NANDN U715 ( .A(n491), .B(n490), .Z(n492) );
  NAND U716 ( .A(n493), .B(n492), .Z(n547) );
  NANDN U717 ( .A(n495), .B(n494), .Z(n499) );
  NANDN U718 ( .A(n497), .B(n496), .Z(n498) );
  NAND U719 ( .A(n499), .B(n498), .Z(n554) );
  NANDN U720 ( .A(n501), .B(n500), .Z(n505) );
  NANDN U721 ( .A(n503), .B(n502), .Z(n504) );
  NAND U722 ( .A(n505), .B(n504), .Z(n553) );
  NANDN U723 ( .A(n507), .B(n506), .Z(n511) );
  NAND U724 ( .A(n509), .B(n508), .Z(n510) );
  NAND U725 ( .A(n511), .B(n510), .Z(n592) );
  XNOR U726 ( .A(n4744), .B(n1043), .Z(n574) );
  NANDN U727 ( .A(n574), .B(n4745), .Z(n514) );
  NANDN U728 ( .A(n512), .B(n4746), .Z(n513) );
  NAND U729 ( .A(n514), .B(n513), .Z(n561) );
  AND U730 ( .A(n760), .B(n4859), .Z(n517) );
  AND U731 ( .A(a[0]), .B(b[9]), .Z(n515) );
  NANDN U732 ( .A(n515), .B(n5033), .Z(n516) );
  NANDN U733 ( .A(n517), .B(n516), .Z(n518) );
  NAND U734 ( .A(b[11]), .B(n518), .Z(n558) );
  NAND U735 ( .A(n519), .B(n4521), .Z(n521) );
  IV U736 ( .A(a[9]), .Z(n1358) );
  XNOR U737 ( .A(n208), .B(n1358), .Z(n577) );
  OR U738 ( .A(n577), .B(n4488), .Z(n520) );
  NAND U739 ( .A(n521), .B(n520), .Z(n559) );
  XOR U740 ( .A(n558), .B(n559), .Z(n560) );
  XNOR U741 ( .A(n561), .B(n560), .Z(n593) );
  XNOR U742 ( .A(n592), .B(n593), .Z(n594) );
  XOR U743 ( .A(n4859), .B(a[3]), .Z(n583) );
  OR U744 ( .A(n583), .B(n4860), .Z(n524) );
  NAND U745 ( .A(n522), .B(n4915), .Z(n523) );
  NAND U746 ( .A(n524), .B(n523), .Z(n573) );
  XOR U747 ( .A(b[11]), .B(a[0]), .Z(n527) );
  XNOR U748 ( .A(b[11]), .B(n5033), .Z(n525) );
  XOR U749 ( .A(b[11]), .B(b[9]), .Z(n564) );
  AND U750 ( .A(n525), .B(n564), .Z(n526) );
  NAND U751 ( .A(n527), .B(n526), .Z(n529) );
  IV U752 ( .A(b[11]), .Z(n4909) );
  XNOR U753 ( .A(n4909), .B(n770), .Z(n566) );
  OR U754 ( .A(n566), .B(n4986), .Z(n528) );
  NAND U755 ( .A(n529), .B(n528), .Z(n572) );
  XNOR U756 ( .A(n573), .B(n572), .Z(n589) );
  NAND U757 ( .A(b[0]), .B(a[11]), .Z(n530) );
  XNOR U758 ( .A(b[1]), .B(n530), .Z(n532) );
  NAND U759 ( .A(n206), .B(a[10]), .Z(n531) );
  AND U760 ( .A(n532), .B(n531), .Z(n587) );
  NAND U761 ( .A(n4669), .B(n533), .Z(n535) );
  XNOR U762 ( .A(n209), .B(n1189), .Z(n569) );
  OR U763 ( .A(n569), .B(n4612), .Z(n534) );
  AND U764 ( .A(n535), .B(n534), .Z(n586) );
  XNOR U765 ( .A(n587), .B(n586), .Z(n588) );
  XOR U766 ( .A(n589), .B(n588), .Z(n595) );
  XOR U767 ( .A(n594), .B(n595), .Z(n552) );
  XNOR U768 ( .A(n553), .B(n552), .Z(n555) );
  XNOR U769 ( .A(n554), .B(n555), .Z(n546) );
  XOR U770 ( .A(n547), .B(n546), .Z(n548) );
  XNOR U771 ( .A(n549), .B(n548), .Z(n541) );
  XNOR U772 ( .A(n541), .B(sreg[59]), .Z(n543) );
  NAND U773 ( .A(n536), .B(sreg[58]), .Z(n540) );
  OR U774 ( .A(n538), .B(n537), .Z(n539) );
  AND U775 ( .A(n540), .B(n539), .Z(n542) );
  XOR U776 ( .A(n543), .B(n542), .Z(c[59]) );
  NAND U777 ( .A(n541), .B(sreg[59]), .Z(n545) );
  OR U778 ( .A(n543), .B(n542), .Z(n544) );
  NAND U779 ( .A(n545), .B(n544), .Z(n657) );
  XNOR U780 ( .A(n657), .B(sreg[60]), .Z(n659) );
  NAND U781 ( .A(n547), .B(n546), .Z(n551) );
  NAND U782 ( .A(n549), .B(n548), .Z(n550) );
  NAND U783 ( .A(n551), .B(n550), .Z(n601) );
  NAND U784 ( .A(n553), .B(n552), .Z(n557) );
  NANDN U785 ( .A(n555), .B(n554), .Z(n556) );
  NAND U786 ( .A(n557), .B(n556), .Z(n598) );
  NANDN U787 ( .A(n559), .B(n558), .Z(n563) );
  OR U788 ( .A(n561), .B(n560), .Z(n562) );
  NAND U789 ( .A(n563), .B(n562), .Z(n607) );
  XOR U790 ( .A(b[11]), .B(b[10]), .Z(n565) );
  AND U791 ( .A(n565), .B(n564), .Z(n4987) );
  NANDN U792 ( .A(n566), .B(n4987), .Z(n568) );
  XNOR U793 ( .A(n4909), .B(n839), .Z(n633) );
  OR U794 ( .A(n633), .B(n4986), .Z(n567) );
  NAND U795 ( .A(n568), .B(n567), .Z(n652) );
  NANDN U796 ( .A(n569), .B(n4669), .Z(n571) );
  XOR U797 ( .A(b[5]), .B(a[8]), .Z(n630) );
  NANDN U798 ( .A(n4612), .B(n630), .Z(n570) );
  AND U799 ( .A(n571), .B(n570), .Z(n651) );
  NAND U800 ( .A(n573), .B(n572), .Z(n613) );
  XNOR U801 ( .A(n4744), .B(n1119), .Z(n644) );
  NANDN U802 ( .A(n644), .B(n4745), .Z(n576) );
  NANDN U803 ( .A(n574), .B(n4746), .Z(n575) );
  NAND U804 ( .A(n576), .B(n575), .Z(n611) );
  NANDN U805 ( .A(n577), .B(n4521), .Z(n579) );
  XOR U806 ( .A(n208), .B(a[10]), .Z(n624) );
  OR U807 ( .A(n624), .B(n4488), .Z(n578) );
  AND U808 ( .A(n579), .B(n578), .Z(n610) );
  XNOR U809 ( .A(n611), .B(n610), .Z(n612) );
  XNOR U810 ( .A(n613), .B(n612), .Z(n654) );
  XOR U811 ( .A(n653), .B(n654), .Z(n650) );
  XNOR U812 ( .A(b[12]), .B(b[11]), .Z(n5041) );
  ANDN U813 ( .B(a[0]), .A(n5041), .Z(n619) );
  NAND U814 ( .A(b[0]), .B(a[12]), .Z(n580) );
  XNOR U815 ( .A(b[1]), .B(n580), .Z(n582) );
  NAND U816 ( .A(n206), .B(a[11]), .Z(n581) );
  AND U817 ( .A(n582), .B(n581), .Z(n617) );
  NANDN U818 ( .A(n583), .B(n4915), .Z(n585) );
  XNOR U819 ( .A(b[9]), .B(n971), .Z(n627) );
  NANDN U820 ( .A(n4860), .B(n627), .Z(n584) );
  AND U821 ( .A(n585), .B(n584), .Z(n616) );
  XNOR U822 ( .A(n617), .B(n616), .Z(n618) );
  XOR U823 ( .A(n619), .B(n618), .Z(n647) );
  NANDN U824 ( .A(n587), .B(n586), .Z(n591) );
  NAND U825 ( .A(n589), .B(n588), .Z(n590) );
  NAND U826 ( .A(n591), .B(n590), .Z(n648) );
  XOR U827 ( .A(n647), .B(n648), .Z(n649) );
  XOR U828 ( .A(n650), .B(n649), .Z(n604) );
  NANDN U829 ( .A(n593), .B(n592), .Z(n597) );
  NAND U830 ( .A(n595), .B(n594), .Z(n596) );
  AND U831 ( .A(n597), .B(n596), .Z(n605) );
  XNOR U832 ( .A(n604), .B(n605), .Z(n606) );
  XNOR U833 ( .A(n607), .B(n606), .Z(n599) );
  XNOR U834 ( .A(n598), .B(n599), .Z(n600) );
  XOR U835 ( .A(n601), .B(n600), .Z(n658) );
  XOR U836 ( .A(n659), .B(n658), .Z(c[60]) );
  NANDN U837 ( .A(n599), .B(n598), .Z(n603) );
  NAND U838 ( .A(n601), .B(n600), .Z(n602) );
  NAND U839 ( .A(n603), .B(n602), .Z(n670) );
  NANDN U840 ( .A(n605), .B(n604), .Z(n609) );
  NAND U841 ( .A(n607), .B(n606), .Z(n608) );
  NAND U842 ( .A(n609), .B(n608), .Z(n667) );
  NANDN U843 ( .A(n611), .B(n610), .Z(n615) );
  NAND U844 ( .A(n613), .B(n612), .Z(n614) );
  NAND U845 ( .A(n615), .B(n614), .Z(n708) );
  NANDN U846 ( .A(n617), .B(n616), .Z(n621) );
  NANDN U847 ( .A(n619), .B(n618), .Z(n620) );
  AND U848 ( .A(n621), .B(n620), .Z(n709) );
  XNOR U849 ( .A(n708), .B(n709), .Z(n710) );
  ANDN U850 ( .B(b[13]), .A(b[12]), .Z(n5085) );
  NAND U851 ( .A(n4909), .B(n5085), .Z(n623) );
  IV U852 ( .A(b[13]), .Z(n5129) );
  NOR U853 ( .A(n5129), .B(n5041), .Z(n5086) );
  NAND U854 ( .A(n760), .B(n5086), .Z(n622) );
  NAND U855 ( .A(n623), .B(n622), .Z(n703) );
  NANDN U856 ( .A(n624), .B(n4521), .Z(n626) );
  XOR U857 ( .A(b[3]), .B(a[11]), .Z(n696) );
  NANDN U858 ( .A(n4488), .B(n696), .Z(n625) );
  AND U859 ( .A(n626), .B(n625), .Z(n702) );
  XNOR U860 ( .A(n703), .B(n702), .Z(n704) );
  NAND U861 ( .A(n4915), .B(n627), .Z(n629) );
  XNOR U862 ( .A(b[9]), .B(n1043), .Z(n675) );
  NANDN U863 ( .A(n4860), .B(n675), .Z(n628) );
  AND U864 ( .A(n629), .B(n628), .Z(n705) );
  XNOR U865 ( .A(n704), .B(n705), .Z(n715) );
  XNOR U866 ( .A(b[5]), .B(n1358), .Z(n699) );
  NANDN U867 ( .A(n4612), .B(n699), .Z(n632) );
  NAND U868 ( .A(n630), .B(n4669), .Z(n631) );
  NAND U869 ( .A(n632), .B(n631), .Z(n714) );
  XOR U870 ( .A(n715), .B(n714), .Z(n717) );
  NANDN U871 ( .A(n633), .B(n4987), .Z(n635) );
  XOR U872 ( .A(b[11]), .B(a[3]), .Z(n687) );
  NANDN U873 ( .A(n4986), .B(n687), .Z(n634) );
  NAND U874 ( .A(n635), .B(n634), .Z(n673) );
  XNOR U875 ( .A(b[13]), .B(n770), .Z(n678) );
  ANDN U876 ( .B(n678), .A(n5041), .Z(n640) );
  XOR U877 ( .A(b[13]), .B(a[0]), .Z(n638) );
  XOR U878 ( .A(b[13]), .B(b[12]), .Z(n637) );
  XOR U879 ( .A(b[13]), .B(b[11]), .Z(n636) );
  AND U880 ( .A(n637), .B(n636), .Z(n5052) );
  NAND U881 ( .A(n638), .B(n5052), .Z(n639) );
  NANDN U882 ( .A(n640), .B(n639), .Z(n674) );
  XNOR U883 ( .A(n673), .B(n674), .Z(n684) );
  NAND U884 ( .A(b[0]), .B(a[13]), .Z(n641) );
  XNOR U885 ( .A(b[1]), .B(n641), .Z(n643) );
  NAND U886 ( .A(n206), .B(a[12]), .Z(n642) );
  AND U887 ( .A(n643), .B(n642), .Z(n682) );
  XNOR U888 ( .A(n4744), .B(n1189), .Z(n693) );
  NANDN U889 ( .A(n693), .B(n4745), .Z(n646) );
  NANDN U890 ( .A(n644), .B(n4746), .Z(n645) );
  AND U891 ( .A(n646), .B(n645), .Z(n681) );
  XNOR U892 ( .A(n682), .B(n681), .Z(n683) );
  XOR U893 ( .A(n684), .B(n683), .Z(n716) );
  XNOR U894 ( .A(n717), .B(n716), .Z(n711) );
  XOR U895 ( .A(n710), .B(n711), .Z(n723) );
  NANDN U896 ( .A(n652), .B(n651), .Z(n656) );
  NANDN U897 ( .A(n654), .B(n653), .Z(n655) );
  NAND U898 ( .A(n656), .B(n655), .Z(n721) );
  XNOR U899 ( .A(n720), .B(n721), .Z(n722) );
  XOR U900 ( .A(n723), .B(n722), .Z(n668) );
  XNOR U901 ( .A(n667), .B(n668), .Z(n669) );
  XNOR U902 ( .A(n670), .B(n669), .Z(n662) );
  XNOR U903 ( .A(n662), .B(sreg[61]), .Z(n664) );
  NAND U904 ( .A(n657), .B(sreg[60]), .Z(n661) );
  OR U905 ( .A(n659), .B(n658), .Z(n660) );
  AND U906 ( .A(n661), .B(n660), .Z(n663) );
  XOR U907 ( .A(n664), .B(n663), .Z(c[61]) );
  NAND U908 ( .A(n662), .B(sreg[61]), .Z(n666) );
  OR U909 ( .A(n664), .B(n663), .Z(n665) );
  NAND U910 ( .A(n666), .B(n665), .Z(n797) );
  XNOR U911 ( .A(n797), .B(sreg[62]), .Z(n799) );
  NANDN U912 ( .A(n668), .B(n667), .Z(n672) );
  NAND U913 ( .A(n670), .B(n669), .Z(n671) );
  NAND U914 ( .A(n672), .B(n671), .Z(n729) );
  AND U915 ( .A(n674), .B(n673), .Z(n789) );
  NAND U916 ( .A(n4915), .B(n675), .Z(n677) );
  XNOR U917 ( .A(b[9]), .B(n1119), .Z(n778) );
  NANDN U918 ( .A(n4860), .B(n778), .Z(n676) );
  NAND U919 ( .A(n677), .B(n676), .Z(n788) );
  NAND U920 ( .A(n5052), .B(n678), .Z(n680) );
  XOR U921 ( .A(b[13]), .B(a[2]), .Z(n767) );
  NANDN U922 ( .A(n5041), .B(n767), .Z(n679) );
  AND U923 ( .A(n680), .B(n679), .Z(n787) );
  XNOR U924 ( .A(n788), .B(n787), .Z(n790) );
  XOR U925 ( .A(n789), .B(n790), .Z(n738) );
  NANDN U926 ( .A(n682), .B(n681), .Z(n686) );
  NAND U927 ( .A(n684), .B(n683), .Z(n685) );
  NAND U928 ( .A(n686), .B(n685), .Z(n739) );
  XOR U929 ( .A(n738), .B(n739), .Z(n741) );
  NAND U930 ( .A(n687), .B(n4987), .Z(n689) );
  XNOR U931 ( .A(n4909), .B(n971), .Z(n750) );
  OR U932 ( .A(n750), .B(n4986), .Z(n688) );
  NAND U933 ( .A(n689), .B(n688), .Z(n782) );
  NAND U934 ( .A(b[0]), .B(a[14]), .Z(n690) );
  XNOR U935 ( .A(b[1]), .B(n690), .Z(n692) );
  NAND U936 ( .A(n206), .B(a[13]), .Z(n691) );
  AND U937 ( .A(n692), .B(n691), .Z(n781) );
  XNOR U938 ( .A(n782), .B(n781), .Z(n784) );
  XOR U939 ( .A(n5129), .B(b[14]), .Z(n5095) );
  ANDN U940 ( .B(a[0]), .A(n5095), .Z(n783) );
  XOR U941 ( .A(n784), .B(n783), .Z(n791) );
  IV U942 ( .A(a[8]), .Z(n1257) );
  XNOR U943 ( .A(n4744), .B(n1257), .Z(n764) );
  NANDN U944 ( .A(n764), .B(n4745), .Z(n695) );
  NANDN U945 ( .A(n693), .B(n4746), .Z(n694) );
  AND U946 ( .A(n695), .B(n694), .Z(n744) );
  NAND U947 ( .A(n696), .B(n4521), .Z(n698) );
  XOR U948 ( .A(n208), .B(a[12]), .Z(n756) );
  OR U949 ( .A(n756), .B(n4488), .Z(n697) );
  AND U950 ( .A(n698), .B(n697), .Z(n745) );
  XOR U951 ( .A(n744), .B(n745), .Z(n746) );
  NAND U952 ( .A(n4669), .B(n699), .Z(n701) );
  XOR U953 ( .A(b[5]), .B(a[10]), .Z(n753) );
  NANDN U954 ( .A(n4612), .B(n753), .Z(n700) );
  AND U955 ( .A(n701), .B(n700), .Z(n747) );
  XOR U956 ( .A(n791), .B(n792), .Z(n793) );
  NANDN U957 ( .A(n703), .B(n702), .Z(n707) );
  NAND U958 ( .A(n705), .B(n704), .Z(n706) );
  AND U959 ( .A(n707), .B(n706), .Z(n794) );
  XNOR U960 ( .A(n793), .B(n794), .Z(n740) );
  XNOR U961 ( .A(n741), .B(n740), .Z(n735) );
  NANDN U962 ( .A(n709), .B(n708), .Z(n713) );
  NANDN U963 ( .A(n711), .B(n710), .Z(n712) );
  NAND U964 ( .A(n713), .B(n712), .Z(n732) );
  OR U965 ( .A(n715), .B(n714), .Z(n719) );
  NAND U966 ( .A(n717), .B(n716), .Z(n718) );
  AND U967 ( .A(n719), .B(n718), .Z(n733) );
  XNOR U968 ( .A(n732), .B(n733), .Z(n734) );
  XNOR U969 ( .A(n735), .B(n734), .Z(n727) );
  NANDN U970 ( .A(n721), .B(n720), .Z(n725) );
  NAND U971 ( .A(n723), .B(n722), .Z(n724) );
  AND U972 ( .A(n725), .B(n724), .Z(n726) );
  XNOR U973 ( .A(n727), .B(n726), .Z(n728) );
  XOR U974 ( .A(n729), .B(n728), .Z(n798) );
  XOR U975 ( .A(n799), .B(n798), .Z(c[62]) );
  NANDN U976 ( .A(n727), .B(n726), .Z(n731) );
  NAND U977 ( .A(n729), .B(n728), .Z(n730) );
  NAND U978 ( .A(n731), .B(n730), .Z(n810) );
  NANDN U979 ( .A(n733), .B(n732), .Z(n737) );
  NAND U980 ( .A(n735), .B(n734), .Z(n736) );
  NAND U981 ( .A(n737), .B(n736), .Z(n808) );
  NANDN U982 ( .A(n739), .B(n738), .Z(n743) );
  OR U983 ( .A(n741), .B(n740), .Z(n742) );
  NAND U984 ( .A(n743), .B(n742), .Z(n814) );
  OR U985 ( .A(n745), .B(n744), .Z(n749) );
  NANDN U986 ( .A(n747), .B(n746), .Z(n748) );
  NAND U987 ( .A(n749), .B(n748), .Z(n867) );
  NANDN U988 ( .A(n750), .B(n4987), .Z(n752) );
  XNOR U989 ( .A(n4909), .B(n1043), .Z(n836) );
  OR U990 ( .A(n836), .B(n4986), .Z(n751) );
  NAND U991 ( .A(n752), .B(n751), .Z(n819) );
  NAND U992 ( .A(n4669), .B(n753), .Z(n755) );
  XOR U993 ( .A(b[5]), .B(a[11]), .Z(n833) );
  NANDN U994 ( .A(n4612), .B(n833), .Z(n754) );
  AND U995 ( .A(n755), .B(n754), .Z(n817) );
  NANDN U996 ( .A(n756), .B(n4521), .Z(n758) );
  XOR U997 ( .A(n208), .B(a[13]), .Z(n848) );
  OR U998 ( .A(n848), .B(n4488), .Z(n757) );
  NAND U999 ( .A(n758), .B(n757), .Z(n818) );
  XOR U1000 ( .A(n817), .B(n818), .Z(n820) );
  XOR U1001 ( .A(n819), .B(n820), .Z(n857) );
  AND U1002 ( .A(a[0]), .B(b[13]), .Z(n759) );
  OR U1003 ( .A(n759), .B(b[14]), .Z(n762) );
  NAND U1004 ( .A(n760), .B(n5129), .Z(n761) );
  NAND U1005 ( .A(n762), .B(n761), .Z(n763) );
  ANDN U1006 ( .B(n763), .A(n210), .Z(n854) );
  XNOR U1007 ( .A(n4744), .B(n1358), .Z(n843) );
  NANDN U1008 ( .A(n843), .B(n4745), .Z(n766) );
  NANDN U1009 ( .A(n764), .B(n4746), .Z(n765) );
  NAND U1010 ( .A(n766), .B(n765), .Z(n855) );
  XOR U1011 ( .A(n854), .B(n855), .Z(n856) );
  XOR U1012 ( .A(n857), .B(n856), .Z(n866) );
  XOR U1013 ( .A(n867), .B(n866), .Z(n868) );
  XOR U1014 ( .A(n5129), .B(a[3]), .Z(n830) );
  OR U1015 ( .A(n830), .B(n5041), .Z(n769) );
  NAND U1016 ( .A(n767), .B(n5052), .Z(n768) );
  NAND U1017 ( .A(n769), .B(n768), .Z(n847) );
  XNOR U1018 ( .A(b[15]), .B(n770), .Z(n840) );
  ANDN U1019 ( .B(n840), .A(n5095), .Z(n774) );
  XOR U1020 ( .A(b[15]), .B(a[0]), .Z(n772) );
  XOR U1021 ( .A(b[15]), .B(b[13]), .Z(n5131) );
  XOR U1022 ( .A(b[15]), .B(b[14]), .Z(n771) );
  AND U1023 ( .A(n5131), .B(n771), .Z(n5092) );
  NAND U1024 ( .A(n772), .B(n5092), .Z(n773) );
  NANDN U1025 ( .A(n774), .B(n773), .Z(n846) );
  XNOR U1026 ( .A(n847), .B(n846), .Z(n824) );
  NAND U1027 ( .A(b[0]), .B(a[15]), .Z(n775) );
  XNOR U1028 ( .A(b[1]), .B(n775), .Z(n777) );
  NAND U1029 ( .A(a[14]), .B(n206), .Z(n776) );
  AND U1030 ( .A(n777), .B(n776), .Z(n822) );
  NAND U1031 ( .A(n4915), .B(n778), .Z(n780) );
  XNOR U1032 ( .A(b[9]), .B(n1189), .Z(n851) );
  NANDN U1033 ( .A(n4860), .B(n851), .Z(n779) );
  AND U1034 ( .A(n780), .B(n779), .Z(n821) );
  XNOR U1035 ( .A(n822), .B(n821), .Z(n823) );
  XOR U1036 ( .A(n824), .B(n823), .Z(n869) );
  XNOR U1037 ( .A(n868), .B(n869), .Z(n813) );
  XOR U1038 ( .A(n814), .B(n813), .Z(n815) );
  OR U1039 ( .A(n782), .B(n781), .Z(n786) );
  OR U1040 ( .A(n784), .B(n783), .Z(n785) );
  NAND U1041 ( .A(n786), .B(n785), .Z(n863) );
  OR U1042 ( .A(n792), .B(n791), .Z(n796) );
  NAND U1043 ( .A(n794), .B(n793), .Z(n795) );
  NAND U1044 ( .A(n796), .B(n795), .Z(n861) );
  XNOR U1045 ( .A(n860), .B(n861), .Z(n862) );
  XOR U1046 ( .A(n863), .B(n862), .Z(n816) );
  XNOR U1047 ( .A(n815), .B(n816), .Z(n807) );
  XOR U1048 ( .A(n808), .B(n807), .Z(n809) );
  XNOR U1049 ( .A(n810), .B(n809), .Z(n802) );
  XNOR U1050 ( .A(n802), .B(sreg[63]), .Z(n804) );
  NAND U1051 ( .A(n797), .B(sreg[62]), .Z(n801) );
  OR U1052 ( .A(n799), .B(n798), .Z(n800) );
  AND U1053 ( .A(n801), .B(n800), .Z(n803) );
  XOR U1054 ( .A(n804), .B(n803), .Z(c[63]) );
  NAND U1055 ( .A(n802), .B(sreg[63]), .Z(n806) );
  OR U1056 ( .A(n804), .B(n803), .Z(n805) );
  NAND U1057 ( .A(n806), .B(n805), .Z(n938) );
  XNOR U1058 ( .A(n938), .B(sreg[64]), .Z(n940) );
  NAND U1059 ( .A(n808), .B(n807), .Z(n812) );
  NAND U1060 ( .A(n810), .B(n809), .Z(n811) );
  NAND U1061 ( .A(n812), .B(n811), .Z(n873) );
  NANDN U1062 ( .A(n822), .B(n821), .Z(n826) );
  NAND U1063 ( .A(n824), .B(n823), .Z(n825) );
  AND U1064 ( .A(n826), .B(n825), .Z(n928) );
  NAND U1065 ( .A(b[0]), .B(a[16]), .Z(n827) );
  XNOR U1066 ( .A(b[1]), .B(n827), .Z(n829) );
  NAND U1067 ( .A(n206), .B(a[15]), .Z(n828) );
  AND U1068 ( .A(n829), .B(n828), .Z(n907) );
  XNOR U1069 ( .A(n5129), .B(n971), .Z(n916) );
  OR U1070 ( .A(n916), .B(n5041), .Z(n832) );
  NANDN U1071 ( .A(n830), .B(n5052), .Z(n831) );
  AND U1072 ( .A(n832), .B(n831), .Z(n908) );
  XOR U1073 ( .A(n907), .B(n908), .Z(n910) );
  NAND U1074 ( .A(b[15]), .B(a[0]), .Z(n909) );
  XOR U1075 ( .A(n910), .B(n909), .Z(n929) );
  XOR U1076 ( .A(n928), .B(n929), .Z(n930) );
  XNOR U1077 ( .A(n931), .B(n930), .Z(n935) );
  XOR U1078 ( .A(n209), .B(a[12]), .Z(n922) );
  OR U1079 ( .A(n922), .B(n4612), .Z(n835) );
  NAND U1080 ( .A(n833), .B(n4669), .Z(n834) );
  NAND U1081 ( .A(n835), .B(n834), .Z(n900) );
  NANDN U1082 ( .A(n836), .B(n4987), .Z(n838) );
  XNOR U1083 ( .A(n4909), .B(n1119), .Z(n891) );
  OR U1084 ( .A(n891), .B(n4986), .Z(n837) );
  NAND U1085 ( .A(n838), .B(n837), .Z(n897) );
  XNOR U1086 ( .A(n210), .B(n839), .Z(n894) );
  OR U1087 ( .A(n894), .B(n5095), .Z(n842) );
  NAND U1088 ( .A(n840), .B(n5092), .Z(n841) );
  AND U1089 ( .A(n842), .B(n841), .Z(n898) );
  XOR U1090 ( .A(n897), .B(n898), .Z(n899) );
  XOR U1091 ( .A(n900), .B(n899), .Z(n901) );
  XOR U1092 ( .A(b[7]), .B(a[10]), .Z(n925) );
  NAND U1093 ( .A(n4745), .B(n925), .Z(n845) );
  NANDN U1094 ( .A(n843), .B(n4746), .Z(n844) );
  NAND U1095 ( .A(n845), .B(n844), .Z(n902) );
  XOR U1096 ( .A(n901), .B(n902), .Z(n904) );
  NAND U1097 ( .A(n847), .B(n846), .Z(n885) );
  NANDN U1098 ( .A(n848), .B(n4521), .Z(n850) );
  XOR U1099 ( .A(b[3]), .B(a[14]), .Z(n919) );
  NANDN U1100 ( .A(n4488), .B(n919), .Z(n849) );
  NAND U1101 ( .A(n850), .B(n849), .Z(n883) );
  NAND U1102 ( .A(n4915), .B(n851), .Z(n853) );
  XOR U1103 ( .A(b[9]), .B(a[8]), .Z(n888) );
  NANDN U1104 ( .A(n4860), .B(n888), .Z(n852) );
  AND U1105 ( .A(n853), .B(n852), .Z(n882) );
  XNOR U1106 ( .A(n883), .B(n882), .Z(n884) );
  XNOR U1107 ( .A(n885), .B(n884), .Z(n903) );
  XNOR U1108 ( .A(n904), .B(n903), .Z(n932) );
  OR U1109 ( .A(n855), .B(n854), .Z(n859) );
  NAND U1110 ( .A(n857), .B(n856), .Z(n858) );
  NAND U1111 ( .A(n859), .B(n858), .Z(n933) );
  XNOR U1112 ( .A(n932), .B(n933), .Z(n934) );
  XNOR U1113 ( .A(n935), .B(n934), .Z(n879) );
  NANDN U1114 ( .A(n861), .B(n860), .Z(n865) );
  NAND U1115 ( .A(n863), .B(n862), .Z(n864) );
  NAND U1116 ( .A(n865), .B(n864), .Z(n876) );
  XNOR U1117 ( .A(n876), .B(n877), .Z(n878) );
  XOR U1118 ( .A(n879), .B(n878), .Z(n871) );
  XNOR U1119 ( .A(n870), .B(n871), .Z(n872) );
  XOR U1120 ( .A(n873), .B(n872), .Z(n939) );
  XOR U1121 ( .A(n940), .B(n939), .Z(c[64]) );
  NANDN U1122 ( .A(n871), .B(n870), .Z(n875) );
  NAND U1123 ( .A(n873), .B(n872), .Z(n874) );
  NAND U1124 ( .A(n875), .B(n874), .Z(n946) );
  NANDN U1125 ( .A(n877), .B(n876), .Z(n881) );
  NANDN U1126 ( .A(n879), .B(n878), .Z(n880) );
  NAND U1127 ( .A(n881), .B(n880), .Z(n944) );
  NANDN U1128 ( .A(n883), .B(n882), .Z(n887) );
  NAND U1129 ( .A(n885), .B(n884), .Z(n886) );
  NAND U1130 ( .A(n887), .B(n886), .Z(n959) );
  XNOR U1131 ( .A(n4859), .B(n1358), .Z(n965) );
  OR U1132 ( .A(n965), .B(n4860), .Z(n890) );
  NAND U1133 ( .A(n888), .B(n4915), .Z(n889) );
  NAND U1134 ( .A(n890), .B(n889), .Z(n978) );
  NANDN U1135 ( .A(n891), .B(n4987), .Z(n893) );
  XNOR U1136 ( .A(n4909), .B(n1189), .Z(n968) );
  OR U1137 ( .A(n968), .B(n4986), .Z(n892) );
  NAND U1138 ( .A(n893), .B(n892), .Z(n975) );
  XOR U1139 ( .A(n210), .B(a[3]), .Z(n972) );
  OR U1140 ( .A(n972), .B(n5095), .Z(n896) );
  NANDN U1141 ( .A(n894), .B(n5092), .Z(n895) );
  AND U1142 ( .A(n896), .B(n895), .Z(n976) );
  XNOR U1143 ( .A(n975), .B(n976), .Z(n977) );
  XOR U1144 ( .A(n978), .B(n977), .Z(n960) );
  XNOR U1145 ( .A(n959), .B(n960), .Z(n961) );
  XNOR U1146 ( .A(n961), .B(n962), .Z(n956) );
  NANDN U1147 ( .A(n902), .B(n901), .Z(n906) );
  OR U1148 ( .A(n904), .B(n903), .Z(n905) );
  NAND U1149 ( .A(n906), .B(n905), .Z(n953) );
  NANDN U1150 ( .A(n908), .B(n907), .Z(n912) );
  OR U1151 ( .A(n910), .B(n909), .Z(n911) );
  NAND U1152 ( .A(n912), .B(n911), .Z(n990) );
  NAND U1153 ( .A(b[0]), .B(a[17]), .Z(n913) );
  XNOR U1154 ( .A(b[1]), .B(n913), .Z(n915) );
  NAND U1155 ( .A(a[16]), .B(n206), .Z(n914) );
  AND U1156 ( .A(n915), .B(n914), .Z(n993) );
  XNOR U1157 ( .A(n5129), .B(n1043), .Z(n999) );
  OR U1158 ( .A(n999), .B(n5041), .Z(n918) );
  NANDN U1159 ( .A(n916), .B(n5052), .Z(n917) );
  AND U1160 ( .A(n918), .B(n917), .Z(n994) );
  XOR U1161 ( .A(n993), .B(n994), .Z(n996) );
  NAND U1162 ( .A(a[1]), .B(b[15]), .Z(n995) );
  XOR U1163 ( .A(n996), .B(n995), .Z(n987) );
  NAND U1164 ( .A(n919), .B(n4521), .Z(n921) );
  XOR U1165 ( .A(b[3]), .B(a[15]), .Z(n1005) );
  NANDN U1166 ( .A(n4488), .B(n1005), .Z(n920) );
  NAND U1167 ( .A(n921), .B(n920), .Z(n983) );
  XOR U1168 ( .A(n209), .B(a[13]), .Z(n1008) );
  OR U1169 ( .A(n1008), .B(n4612), .Z(n924) );
  NANDN U1170 ( .A(n922), .B(n4669), .Z(n923) );
  NAND U1171 ( .A(n924), .B(n923), .Z(n981) );
  XOR U1172 ( .A(n4744), .B(a[11]), .Z(n1011) );
  NANDN U1173 ( .A(n1011), .B(n4745), .Z(n927) );
  NAND U1174 ( .A(n925), .B(n4746), .Z(n926) );
  AND U1175 ( .A(n927), .B(n926), .Z(n982) );
  XOR U1176 ( .A(n983), .B(n984), .Z(n988) );
  XNOR U1177 ( .A(n987), .B(n988), .Z(n989) );
  XOR U1178 ( .A(n990), .B(n989), .Z(n954) );
  XNOR U1179 ( .A(n953), .B(n954), .Z(n955) );
  XOR U1180 ( .A(n956), .B(n955), .Z(n951) );
  NANDN U1181 ( .A(n933), .B(n932), .Z(n937) );
  NANDN U1182 ( .A(n935), .B(n934), .Z(n936) );
  NAND U1183 ( .A(n937), .B(n936), .Z(n950) );
  XNOR U1184 ( .A(n949), .B(n950), .Z(n952) );
  XNOR U1185 ( .A(n951), .B(n952), .Z(n943) );
  XOR U1186 ( .A(n944), .B(n943), .Z(n945) );
  XNOR U1187 ( .A(n946), .B(n945), .Z(n1014) );
  XNOR U1188 ( .A(n1014), .B(sreg[65]), .Z(n1016) );
  NAND U1189 ( .A(n938), .B(sreg[64]), .Z(n942) );
  OR U1190 ( .A(n940), .B(n939), .Z(n941) );
  AND U1191 ( .A(n942), .B(n941), .Z(n1015) );
  XOR U1192 ( .A(n1016), .B(n1015), .Z(c[65]) );
  NAND U1193 ( .A(n944), .B(n943), .Z(n948) );
  NAND U1194 ( .A(n946), .B(n945), .Z(n947) );
  NAND U1195 ( .A(n948), .B(n947), .Z(n1022) );
  NANDN U1196 ( .A(n954), .B(n953), .Z(n958) );
  NANDN U1197 ( .A(n956), .B(n955), .Z(n957) );
  NAND U1198 ( .A(n958), .B(n957), .Z(n1086) );
  NANDN U1199 ( .A(n960), .B(n959), .Z(n964) );
  NAND U1200 ( .A(n962), .B(n961), .Z(n963) );
  NAND U1201 ( .A(n964), .B(n963), .Z(n1085) );
  XOR U1202 ( .A(n4859), .B(a[10]), .Z(n1037) );
  OR U1203 ( .A(n1037), .B(n4860), .Z(n967) );
  NANDN U1204 ( .A(n965), .B(n4915), .Z(n966) );
  NAND U1205 ( .A(n967), .B(n966), .Z(n1050) );
  NANDN U1206 ( .A(n968), .B(n4987), .Z(n970) );
  XNOR U1207 ( .A(n4909), .B(n1257), .Z(n1040) );
  OR U1208 ( .A(n1040), .B(n4986), .Z(n969) );
  NAND U1209 ( .A(n970), .B(n969), .Z(n1047) );
  XNOR U1210 ( .A(n210), .B(n971), .Z(n1044) );
  OR U1211 ( .A(n1044), .B(n5095), .Z(n974) );
  NANDN U1212 ( .A(n972), .B(n5092), .Z(n973) );
  AND U1213 ( .A(n974), .B(n973), .Z(n1048) );
  XOR U1214 ( .A(n1047), .B(n1048), .Z(n1049) );
  XOR U1215 ( .A(n1050), .B(n1049), .Z(n1031) );
  NANDN U1216 ( .A(n976), .B(n975), .Z(n980) );
  NAND U1217 ( .A(n978), .B(n977), .Z(n979) );
  NAND U1218 ( .A(n980), .B(n979), .Z(n1032) );
  XNOR U1219 ( .A(n1031), .B(n1032), .Z(n1033) );
  NANDN U1220 ( .A(n982), .B(n981), .Z(n986) );
  NANDN U1221 ( .A(n984), .B(n983), .Z(n985) );
  NAND U1222 ( .A(n986), .B(n985), .Z(n1034) );
  XOR U1223 ( .A(n1033), .B(n1034), .Z(n1028) );
  NANDN U1224 ( .A(n988), .B(n987), .Z(n992) );
  NAND U1225 ( .A(n990), .B(n989), .Z(n991) );
  NAND U1226 ( .A(n992), .B(n991), .Z(n1025) );
  NANDN U1227 ( .A(n994), .B(n993), .Z(n998) );
  OR U1228 ( .A(n996), .B(n995), .Z(n997) );
  NAND U1229 ( .A(n998), .B(n997), .Z(n1081) );
  XNOR U1230 ( .A(n5129), .B(n1119), .Z(n1060) );
  OR U1231 ( .A(n1060), .B(n5041), .Z(n1001) );
  NANDN U1232 ( .A(n999), .B(n5052), .Z(n1000) );
  AND U1233 ( .A(n1001), .B(n1000), .Z(n1073) );
  NAND U1234 ( .A(b[0]), .B(a[18]), .Z(n1002) );
  XNOR U1235 ( .A(b[1]), .B(n1002), .Z(n1004) );
  NAND U1236 ( .A(n206), .B(a[17]), .Z(n1003) );
  AND U1237 ( .A(n1004), .B(n1003), .Z(n1072) );
  XOR U1238 ( .A(n1073), .B(n1072), .Z(n1075) );
  NAND U1239 ( .A(a[2]), .B(b[15]), .Z(n1074) );
  XOR U1240 ( .A(n1075), .B(n1074), .Z(n1078) );
  NAND U1241 ( .A(n4521), .B(n1005), .Z(n1007) );
  IV U1242 ( .A(a[16]), .Z(n1852) );
  XNOR U1243 ( .A(b[3]), .B(n1852), .Z(n1063) );
  NANDN U1244 ( .A(n4488), .B(n1063), .Z(n1006) );
  NAND U1245 ( .A(n1007), .B(n1006), .Z(n1053) );
  IV U1246 ( .A(a[14]), .Z(n1705) );
  XNOR U1247 ( .A(n209), .B(n1705), .Z(n1066) );
  OR U1248 ( .A(n1066), .B(n4612), .Z(n1010) );
  NANDN U1249 ( .A(n1008), .B(n4669), .Z(n1009) );
  NAND U1250 ( .A(n1010), .B(n1009), .Z(n1051) );
  XOR U1251 ( .A(n4744), .B(a[12]), .Z(n1069) );
  NANDN U1252 ( .A(n1069), .B(n4745), .Z(n1013) );
  NANDN U1253 ( .A(n1011), .B(n4746), .Z(n1012) );
  AND U1254 ( .A(n1013), .B(n1012), .Z(n1052) );
  XOR U1255 ( .A(n1053), .B(n1054), .Z(n1079) );
  XNOR U1256 ( .A(n1078), .B(n1079), .Z(n1080) );
  XNOR U1257 ( .A(n1081), .B(n1080), .Z(n1026) );
  XNOR U1258 ( .A(n1025), .B(n1026), .Z(n1027) );
  XOR U1259 ( .A(n1028), .B(n1027), .Z(n1084) );
  XOR U1260 ( .A(n1085), .B(n1084), .Z(n1087) );
  XOR U1261 ( .A(n1086), .B(n1087), .Z(n1020) );
  XNOR U1262 ( .A(n1019), .B(n1020), .Z(n1021) );
  XNOR U1263 ( .A(n1022), .B(n1021), .Z(n1090) );
  XNOR U1264 ( .A(n1090), .B(sreg[66]), .Z(n1092) );
  NAND U1265 ( .A(n1014), .B(sreg[65]), .Z(n1018) );
  OR U1266 ( .A(n1016), .B(n1015), .Z(n1017) );
  AND U1267 ( .A(n1018), .B(n1017), .Z(n1091) );
  XOR U1268 ( .A(n1092), .B(n1091), .Z(c[66]) );
  NANDN U1269 ( .A(n1020), .B(n1019), .Z(n1024) );
  NAND U1270 ( .A(n1022), .B(n1021), .Z(n1023) );
  NAND U1271 ( .A(n1024), .B(n1023), .Z(n1098) );
  NANDN U1272 ( .A(n1026), .B(n1025), .Z(n1030) );
  NAND U1273 ( .A(n1028), .B(n1027), .Z(n1029) );
  NAND U1274 ( .A(n1030), .B(n1029), .Z(n1160) );
  NANDN U1275 ( .A(n1032), .B(n1031), .Z(n1036) );
  NANDN U1276 ( .A(n1034), .B(n1033), .Z(n1035) );
  NAND U1277 ( .A(n1036), .B(n1035), .Z(n1161) );
  XNOR U1278 ( .A(n1160), .B(n1161), .Z(n1162) );
  XOR U1279 ( .A(n4859), .B(a[11]), .Z(n1113) );
  OR U1280 ( .A(n1113), .B(n4860), .Z(n1039) );
  NANDN U1281 ( .A(n1037), .B(n4915), .Z(n1038) );
  NAND U1282 ( .A(n1039), .B(n1038), .Z(n1126) );
  NANDN U1283 ( .A(n1040), .B(n4987), .Z(n1042) );
  XNOR U1284 ( .A(n4909), .B(n1358), .Z(n1116) );
  OR U1285 ( .A(n1116), .B(n4986), .Z(n1041) );
  NAND U1286 ( .A(n1042), .B(n1041), .Z(n1123) );
  XNOR U1287 ( .A(n210), .B(n1043), .Z(n1120) );
  OR U1288 ( .A(n1120), .B(n5095), .Z(n1046) );
  NANDN U1289 ( .A(n1044), .B(n5092), .Z(n1045) );
  AND U1290 ( .A(n1046), .B(n1045), .Z(n1124) );
  XOR U1291 ( .A(n1123), .B(n1124), .Z(n1125) );
  XOR U1292 ( .A(n1126), .B(n1125), .Z(n1107) );
  XNOR U1293 ( .A(n1107), .B(n1108), .Z(n1109) );
  NANDN U1294 ( .A(n1052), .B(n1051), .Z(n1056) );
  NANDN U1295 ( .A(n1054), .B(n1053), .Z(n1055) );
  NAND U1296 ( .A(n1056), .B(n1055), .Z(n1110) );
  XOR U1297 ( .A(n1109), .B(n1110), .Z(n1104) );
  NAND U1298 ( .A(b[0]), .B(a[19]), .Z(n1057) );
  XNOR U1299 ( .A(b[1]), .B(n1057), .Z(n1059) );
  NAND U1300 ( .A(a[18]), .B(n206), .Z(n1058) );
  AND U1301 ( .A(n1059), .B(n1058), .Z(n1139) );
  XNOR U1302 ( .A(n5129), .B(n1189), .Z(n1145) );
  OR U1303 ( .A(n1145), .B(n5041), .Z(n1062) );
  NANDN U1304 ( .A(n1060), .B(n5052), .Z(n1061) );
  AND U1305 ( .A(n1062), .B(n1061), .Z(n1140) );
  XOR U1306 ( .A(n1139), .B(n1140), .Z(n1142) );
  NAND U1307 ( .A(b[15]), .B(a[3]), .Z(n1141) );
  XNOR U1308 ( .A(n1142), .B(n1141), .Z(n1133) );
  NAND U1309 ( .A(n4521), .B(n1063), .Z(n1065) );
  XOR U1310 ( .A(b[3]), .B(a[17]), .Z(n1151) );
  NANDN U1311 ( .A(n4488), .B(n1151), .Z(n1064) );
  NAND U1312 ( .A(n1065), .B(n1064), .Z(n1130) );
  XOR U1313 ( .A(n209), .B(a[15]), .Z(n1154) );
  OR U1314 ( .A(n1154), .B(n4612), .Z(n1068) );
  NANDN U1315 ( .A(n1066), .B(n4669), .Z(n1067) );
  NAND U1316 ( .A(n1068), .B(n1067), .Z(n1127) );
  XOR U1317 ( .A(n4744), .B(a[13]), .Z(n1157) );
  NANDN U1318 ( .A(n1157), .B(n4745), .Z(n1071) );
  NANDN U1319 ( .A(n1069), .B(n4746), .Z(n1070) );
  AND U1320 ( .A(n1071), .B(n1070), .Z(n1128) );
  XNOR U1321 ( .A(n1127), .B(n1128), .Z(n1129) );
  XOR U1322 ( .A(n1130), .B(n1129), .Z(n1134) );
  XNOR U1323 ( .A(n1133), .B(n1134), .Z(n1135) );
  NANDN U1324 ( .A(n1073), .B(n1072), .Z(n1077) );
  OR U1325 ( .A(n1075), .B(n1074), .Z(n1076) );
  NAND U1326 ( .A(n1077), .B(n1076), .Z(n1136) );
  XOR U1327 ( .A(n1135), .B(n1136), .Z(n1101) );
  NANDN U1328 ( .A(n1079), .B(n1078), .Z(n1083) );
  NAND U1329 ( .A(n1081), .B(n1080), .Z(n1082) );
  AND U1330 ( .A(n1083), .B(n1082), .Z(n1102) );
  XNOR U1331 ( .A(n1101), .B(n1102), .Z(n1103) );
  XNOR U1332 ( .A(n1104), .B(n1103), .Z(n1163) );
  XOR U1333 ( .A(n1162), .B(n1163), .Z(n1095) );
  NANDN U1334 ( .A(n1085), .B(n1084), .Z(n1089) );
  OR U1335 ( .A(n1087), .B(n1086), .Z(n1088) );
  NAND U1336 ( .A(n1089), .B(n1088), .Z(n1096) );
  XNOR U1337 ( .A(n1095), .B(n1096), .Z(n1097) );
  XNOR U1338 ( .A(n1098), .B(n1097), .Z(n1166) );
  XNOR U1339 ( .A(n1166), .B(sreg[67]), .Z(n1168) );
  NAND U1340 ( .A(n1090), .B(sreg[66]), .Z(n1094) );
  OR U1341 ( .A(n1092), .B(n1091), .Z(n1093) );
  AND U1342 ( .A(n1094), .B(n1093), .Z(n1167) );
  XOR U1343 ( .A(n1168), .B(n1167), .Z(c[67]) );
  NANDN U1344 ( .A(n1096), .B(n1095), .Z(n1100) );
  NAND U1345 ( .A(n1098), .B(n1097), .Z(n1099) );
  NAND U1346 ( .A(n1100), .B(n1099), .Z(n1174) );
  NANDN U1347 ( .A(n1102), .B(n1101), .Z(n1106) );
  NAND U1348 ( .A(n1104), .B(n1103), .Z(n1105) );
  NAND U1349 ( .A(n1106), .B(n1105), .Z(n1236) );
  NANDN U1350 ( .A(n1108), .B(n1107), .Z(n1112) );
  NANDN U1351 ( .A(n1110), .B(n1109), .Z(n1111) );
  NAND U1352 ( .A(n1112), .B(n1111), .Z(n1237) );
  XNOR U1353 ( .A(n1236), .B(n1237), .Z(n1238) );
  XOR U1354 ( .A(n4859), .B(a[12]), .Z(n1183) );
  OR U1355 ( .A(n1183), .B(n4860), .Z(n1115) );
  NANDN U1356 ( .A(n1113), .B(n4915), .Z(n1114) );
  NAND U1357 ( .A(n1115), .B(n1114), .Z(n1196) );
  NANDN U1358 ( .A(n1116), .B(n4987), .Z(n1118) );
  XOR U1359 ( .A(n4909), .B(a[10]), .Z(n1186) );
  OR U1360 ( .A(n1186), .B(n4986), .Z(n1117) );
  NAND U1361 ( .A(n1118), .B(n1117), .Z(n1193) );
  XNOR U1362 ( .A(n210), .B(n1119), .Z(n1190) );
  OR U1363 ( .A(n1190), .B(n5095), .Z(n1122) );
  NANDN U1364 ( .A(n1120), .B(n5092), .Z(n1121) );
  AND U1365 ( .A(n1122), .B(n1121), .Z(n1194) );
  XOR U1366 ( .A(n1193), .B(n1194), .Z(n1195) );
  XOR U1367 ( .A(n1196), .B(n1195), .Z(n1230) );
  XOR U1368 ( .A(n1230), .B(n1231), .Z(n1233) );
  NANDN U1369 ( .A(n1128), .B(n1127), .Z(n1132) );
  NAND U1370 ( .A(n1130), .B(n1129), .Z(n1131) );
  NAND U1371 ( .A(n1132), .B(n1131), .Z(n1232) );
  XNOR U1372 ( .A(n1233), .B(n1232), .Z(n1180) );
  NANDN U1373 ( .A(n1134), .B(n1133), .Z(n1138) );
  NANDN U1374 ( .A(n1136), .B(n1135), .Z(n1137) );
  NAND U1375 ( .A(n1138), .B(n1137), .Z(n1178) );
  NANDN U1376 ( .A(n1140), .B(n1139), .Z(n1144) );
  OR U1377 ( .A(n1142), .B(n1141), .Z(n1143) );
  NAND U1378 ( .A(n1144), .B(n1143), .Z(n1227) );
  XNOR U1379 ( .A(n5129), .B(n1257), .Z(n1212) );
  OR U1380 ( .A(n1212), .B(n5041), .Z(n1147) );
  NANDN U1381 ( .A(n1145), .B(n5052), .Z(n1146) );
  AND U1382 ( .A(n1147), .B(n1146), .Z(n1204) );
  NAND U1383 ( .A(b[0]), .B(a[20]), .Z(n1148) );
  XNOR U1384 ( .A(b[1]), .B(n1148), .Z(n1150) );
  NAND U1385 ( .A(n206), .B(a[19]), .Z(n1149) );
  AND U1386 ( .A(n1150), .B(n1149), .Z(n1203) );
  XOR U1387 ( .A(n1204), .B(n1203), .Z(n1206) );
  NAND U1388 ( .A(a[4]), .B(b[15]), .Z(n1205) );
  XOR U1389 ( .A(n1206), .B(n1205), .Z(n1224) );
  NAND U1390 ( .A(n4521), .B(n1151), .Z(n1153) );
  IV U1391 ( .A(a[18]), .Z(n2003) );
  XNOR U1392 ( .A(b[3]), .B(n2003), .Z(n1215) );
  NANDN U1393 ( .A(n4488), .B(n1215), .Z(n1152) );
  NAND U1394 ( .A(n1153), .B(n1152), .Z(n1199) );
  XNOR U1395 ( .A(n209), .B(n1852), .Z(n1218) );
  OR U1396 ( .A(n1218), .B(n4612), .Z(n1156) );
  NANDN U1397 ( .A(n1154), .B(n4669), .Z(n1155) );
  NAND U1398 ( .A(n1156), .B(n1155), .Z(n1197) );
  XNOR U1399 ( .A(n4744), .B(n1705), .Z(n1221) );
  NANDN U1400 ( .A(n1221), .B(n4745), .Z(n1159) );
  NANDN U1401 ( .A(n1157), .B(n4746), .Z(n1158) );
  AND U1402 ( .A(n1159), .B(n1158), .Z(n1198) );
  XOR U1403 ( .A(n1199), .B(n1200), .Z(n1225) );
  XNOR U1404 ( .A(n1224), .B(n1225), .Z(n1226) );
  XOR U1405 ( .A(n1227), .B(n1226), .Z(n1177) );
  XNOR U1406 ( .A(n1178), .B(n1177), .Z(n1179) );
  XNOR U1407 ( .A(n1180), .B(n1179), .Z(n1239) );
  XOR U1408 ( .A(n1238), .B(n1239), .Z(n1171) );
  NANDN U1409 ( .A(n1161), .B(n1160), .Z(n1165) );
  NANDN U1410 ( .A(n1163), .B(n1162), .Z(n1164) );
  NAND U1411 ( .A(n1165), .B(n1164), .Z(n1172) );
  XNOR U1412 ( .A(n1171), .B(n1172), .Z(n1173) );
  XNOR U1413 ( .A(n1174), .B(n1173), .Z(n1242) );
  XNOR U1414 ( .A(n1242), .B(sreg[68]), .Z(n1244) );
  NAND U1415 ( .A(n1166), .B(sreg[67]), .Z(n1170) );
  OR U1416 ( .A(n1168), .B(n1167), .Z(n1169) );
  AND U1417 ( .A(n1170), .B(n1169), .Z(n1243) );
  XOR U1418 ( .A(n1244), .B(n1243), .Z(c[68]) );
  NANDN U1419 ( .A(n1172), .B(n1171), .Z(n1176) );
  NAND U1420 ( .A(n1174), .B(n1173), .Z(n1175) );
  NAND U1421 ( .A(n1176), .B(n1175), .Z(n1250) );
  NANDN U1422 ( .A(n1178), .B(n1177), .Z(n1182) );
  NAND U1423 ( .A(n1180), .B(n1179), .Z(n1181) );
  NAND U1424 ( .A(n1182), .B(n1181), .Z(n1313) );
  XOR U1425 ( .A(n4859), .B(a[13]), .Z(n1251) );
  OR U1426 ( .A(n1251), .B(n4860), .Z(n1185) );
  NANDN U1427 ( .A(n1183), .B(n4915), .Z(n1184) );
  NAND U1428 ( .A(n1185), .B(n1184), .Z(n1264) );
  NANDN U1429 ( .A(n1186), .B(n4987), .Z(n1188) );
  XOR U1430 ( .A(n4909), .B(a[11]), .Z(n1254) );
  OR U1431 ( .A(n1254), .B(n4986), .Z(n1187) );
  NAND U1432 ( .A(n1188), .B(n1187), .Z(n1261) );
  XNOR U1433 ( .A(n210), .B(n1189), .Z(n1258) );
  OR U1434 ( .A(n1258), .B(n5095), .Z(n1192) );
  NANDN U1435 ( .A(n1190), .B(n5092), .Z(n1191) );
  AND U1436 ( .A(n1192), .B(n1191), .Z(n1262) );
  XOR U1437 ( .A(n1261), .B(n1262), .Z(n1263) );
  XOR U1438 ( .A(n1264), .B(n1263), .Z(n1298) );
  XOR U1439 ( .A(n1298), .B(n1299), .Z(n1301) );
  NANDN U1440 ( .A(n1198), .B(n1197), .Z(n1202) );
  NANDN U1441 ( .A(n1200), .B(n1199), .Z(n1201) );
  AND U1442 ( .A(n1202), .B(n1201), .Z(n1300) );
  XOR U1443 ( .A(n1301), .B(n1300), .Z(n1306) );
  NANDN U1444 ( .A(n1204), .B(n1203), .Z(n1208) );
  OR U1445 ( .A(n1206), .B(n1205), .Z(n1207) );
  NAND U1446 ( .A(n1208), .B(n1207), .Z(n1295) );
  NAND U1447 ( .A(b[0]), .B(a[21]), .Z(n1209) );
  XNOR U1448 ( .A(b[1]), .B(n1209), .Z(n1211) );
  NAND U1449 ( .A(n206), .B(a[20]), .Z(n1210) );
  AND U1450 ( .A(n1211), .B(n1210), .Z(n1271) );
  XNOR U1451 ( .A(n5129), .B(n1358), .Z(n1280) );
  OR U1452 ( .A(n1280), .B(n5041), .Z(n1214) );
  NANDN U1453 ( .A(n1212), .B(n5052), .Z(n1213) );
  AND U1454 ( .A(n1214), .B(n1213), .Z(n1272) );
  XOR U1455 ( .A(n1271), .B(n1272), .Z(n1274) );
  NAND U1456 ( .A(a[5]), .B(b[15]), .Z(n1273) );
  XOR U1457 ( .A(n1274), .B(n1273), .Z(n1292) );
  NAND U1458 ( .A(n4521), .B(n1215), .Z(n1217) );
  XOR U1459 ( .A(n208), .B(a[19]), .Z(n1283) );
  OR U1460 ( .A(n1283), .B(n4488), .Z(n1216) );
  NAND U1461 ( .A(n1217), .B(n1216), .Z(n1267) );
  XOR U1462 ( .A(b[5]), .B(a[17]), .Z(n1286) );
  NANDN U1463 ( .A(n4612), .B(n1286), .Z(n1220) );
  NANDN U1464 ( .A(n1218), .B(n4669), .Z(n1219) );
  NAND U1465 ( .A(n1220), .B(n1219), .Z(n1265) );
  XOR U1466 ( .A(n4744), .B(a[15]), .Z(n1289) );
  NANDN U1467 ( .A(n1289), .B(n4745), .Z(n1223) );
  NANDN U1468 ( .A(n1221), .B(n4746), .Z(n1222) );
  AND U1469 ( .A(n1223), .B(n1222), .Z(n1266) );
  XOR U1470 ( .A(n1267), .B(n1268), .Z(n1293) );
  XNOR U1471 ( .A(n1292), .B(n1293), .Z(n1294) );
  XNOR U1472 ( .A(n1295), .B(n1294), .Z(n1304) );
  NANDN U1473 ( .A(n1225), .B(n1224), .Z(n1229) );
  NAND U1474 ( .A(n1227), .B(n1226), .Z(n1228) );
  NAND U1475 ( .A(n1229), .B(n1228), .Z(n1305) );
  XOR U1476 ( .A(n1304), .B(n1305), .Z(n1307) );
  XNOR U1477 ( .A(n1306), .B(n1307), .Z(n1310) );
  NANDN U1478 ( .A(n1231), .B(n1230), .Z(n1235) );
  OR U1479 ( .A(n1233), .B(n1232), .Z(n1234) );
  NAND U1480 ( .A(n1235), .B(n1234), .Z(n1311) );
  XNOR U1481 ( .A(n1310), .B(n1311), .Z(n1312) );
  XNOR U1482 ( .A(n1313), .B(n1312), .Z(n1247) );
  NANDN U1483 ( .A(n1237), .B(n1236), .Z(n1241) );
  NANDN U1484 ( .A(n1239), .B(n1238), .Z(n1240) );
  NAND U1485 ( .A(n1241), .B(n1240), .Z(n1248) );
  XOR U1486 ( .A(n1247), .B(n1248), .Z(n1249) );
  XOR U1487 ( .A(n1250), .B(n1249), .Z(n1316) );
  XNOR U1488 ( .A(n1316), .B(sreg[69]), .Z(n1318) );
  NAND U1489 ( .A(n1242), .B(sreg[68]), .Z(n1246) );
  OR U1490 ( .A(n1244), .B(n1243), .Z(n1245) );
  AND U1491 ( .A(n1246), .B(n1245), .Z(n1317) );
  XOR U1492 ( .A(n1318), .B(n1317), .Z(c[69]) );
  XNOR U1493 ( .A(n4859), .B(n1705), .Z(n1352) );
  OR U1494 ( .A(n1352), .B(n4860), .Z(n1253) );
  NANDN U1495 ( .A(n1251), .B(n4915), .Z(n1252) );
  NAND U1496 ( .A(n1253), .B(n1252), .Z(n1365) );
  NANDN U1497 ( .A(n1254), .B(n4987), .Z(n1256) );
  XOR U1498 ( .A(n4909), .B(a[12]), .Z(n1355) );
  OR U1499 ( .A(n1355), .B(n4986), .Z(n1255) );
  NAND U1500 ( .A(n1256), .B(n1255), .Z(n1362) );
  XNOR U1501 ( .A(n210), .B(n1257), .Z(n1359) );
  OR U1502 ( .A(n1359), .B(n5095), .Z(n1260) );
  NANDN U1503 ( .A(n1258), .B(n5092), .Z(n1259) );
  AND U1504 ( .A(n1260), .B(n1259), .Z(n1363) );
  XOR U1505 ( .A(n1362), .B(n1363), .Z(n1364) );
  XOR U1506 ( .A(n1365), .B(n1364), .Z(n1370) );
  XOR U1507 ( .A(n1370), .B(n1371), .Z(n1373) );
  NANDN U1508 ( .A(n1266), .B(n1265), .Z(n1270) );
  NANDN U1509 ( .A(n1268), .B(n1267), .Z(n1269) );
  AND U1510 ( .A(n1270), .B(n1269), .Z(n1372) );
  XOR U1511 ( .A(n1373), .B(n1372), .Z(n1378) );
  NANDN U1512 ( .A(n1272), .B(n1271), .Z(n1276) );
  OR U1513 ( .A(n1274), .B(n1273), .Z(n1275) );
  NAND U1514 ( .A(n1276), .B(n1275), .Z(n1349) );
  NAND U1515 ( .A(b[0]), .B(a[22]), .Z(n1277) );
  XNOR U1516 ( .A(b[1]), .B(n1277), .Z(n1279) );
  NAND U1517 ( .A(n206), .B(a[21]), .Z(n1278) );
  AND U1518 ( .A(n1279), .B(n1278), .Z(n1325) );
  XOR U1519 ( .A(n5129), .B(a[10]), .Z(n1331) );
  OR U1520 ( .A(n1331), .B(n5041), .Z(n1282) );
  NANDN U1521 ( .A(n1280), .B(n5052), .Z(n1281) );
  AND U1522 ( .A(n1282), .B(n1281), .Z(n1326) );
  XOR U1523 ( .A(n1325), .B(n1326), .Z(n1328) );
  NAND U1524 ( .A(a[6]), .B(b[15]), .Z(n1327) );
  XOR U1525 ( .A(n1328), .B(n1327), .Z(n1346) );
  NANDN U1526 ( .A(n1283), .B(n4521), .Z(n1285) );
  XOR U1527 ( .A(b[3]), .B(a[20]), .Z(n1337) );
  NANDN U1528 ( .A(n4488), .B(n1337), .Z(n1284) );
  AND U1529 ( .A(n1285), .B(n1284), .Z(n1368) );
  NAND U1530 ( .A(n4669), .B(n1286), .Z(n1288) );
  XOR U1531 ( .A(b[5]), .B(a[18]), .Z(n1340) );
  NANDN U1532 ( .A(n4612), .B(n1340), .Z(n1287) );
  AND U1533 ( .A(n1288), .B(n1287), .Z(n1366) );
  XNOR U1534 ( .A(n4744), .B(n1852), .Z(n1343) );
  NANDN U1535 ( .A(n1343), .B(n4745), .Z(n1291) );
  NANDN U1536 ( .A(n1289), .B(n4746), .Z(n1290) );
  AND U1537 ( .A(n1291), .B(n1290), .Z(n1367) );
  XOR U1538 ( .A(n1366), .B(n1367), .Z(n1369) );
  XOR U1539 ( .A(n1368), .B(n1369), .Z(n1347) );
  XNOR U1540 ( .A(n1346), .B(n1347), .Z(n1348) );
  XNOR U1541 ( .A(n1349), .B(n1348), .Z(n1376) );
  NANDN U1542 ( .A(n1293), .B(n1292), .Z(n1297) );
  NAND U1543 ( .A(n1295), .B(n1294), .Z(n1296) );
  NAND U1544 ( .A(n1297), .B(n1296), .Z(n1377) );
  XOR U1545 ( .A(n1376), .B(n1377), .Z(n1379) );
  XNOR U1546 ( .A(n1378), .B(n1379), .Z(n1385) );
  NANDN U1547 ( .A(n1299), .B(n1298), .Z(n1303) );
  NANDN U1548 ( .A(n1301), .B(n1300), .Z(n1302) );
  NAND U1549 ( .A(n1303), .B(n1302), .Z(n1383) );
  NANDN U1550 ( .A(n1305), .B(n1304), .Z(n1309) );
  OR U1551 ( .A(n1307), .B(n1306), .Z(n1308) );
  AND U1552 ( .A(n1309), .B(n1308), .Z(n1382) );
  XNOR U1553 ( .A(n1383), .B(n1382), .Z(n1384) );
  XNOR U1554 ( .A(n1385), .B(n1384), .Z(n1321) );
  NANDN U1555 ( .A(n1311), .B(n1310), .Z(n1315) );
  NAND U1556 ( .A(n1313), .B(n1312), .Z(n1314) );
  NAND U1557 ( .A(n1315), .B(n1314), .Z(n1322) );
  XOR U1558 ( .A(n1321), .B(n1322), .Z(n1323) );
  XOR U1559 ( .A(n1324), .B(n1323), .Z(n1388) );
  XNOR U1560 ( .A(n1388), .B(sreg[70]), .Z(n1390) );
  NAND U1561 ( .A(n1316), .B(sreg[69]), .Z(n1320) );
  OR U1562 ( .A(n1318), .B(n1317), .Z(n1319) );
  AND U1563 ( .A(n1320), .B(n1319), .Z(n1389) );
  XOR U1564 ( .A(n1390), .B(n1389), .Z(c[70]) );
  NANDN U1565 ( .A(n1326), .B(n1325), .Z(n1330) );
  OR U1566 ( .A(n1328), .B(n1327), .Z(n1329) );
  NAND U1567 ( .A(n1330), .B(n1329), .Z(n1450) );
  XOR U1568 ( .A(n5129), .B(a[11]), .Z(n1429) );
  OR U1569 ( .A(n1429), .B(n5041), .Z(n1333) );
  NANDN U1570 ( .A(n1331), .B(n5052), .Z(n1332) );
  AND U1571 ( .A(n1333), .B(n1332), .Z(n1442) );
  NAND U1572 ( .A(b[0]), .B(a[23]), .Z(n1334) );
  XNOR U1573 ( .A(b[1]), .B(n1334), .Z(n1336) );
  NAND U1574 ( .A(n206), .B(a[22]), .Z(n1335) );
  AND U1575 ( .A(n1336), .B(n1335), .Z(n1441) );
  XOR U1576 ( .A(n1442), .B(n1441), .Z(n1444) );
  NAND U1577 ( .A(a[7]), .B(b[15]), .Z(n1443) );
  XOR U1578 ( .A(n1444), .B(n1443), .Z(n1447) );
  NAND U1579 ( .A(n1337), .B(n4521), .Z(n1339) );
  XOR U1580 ( .A(b[3]), .B(a[21]), .Z(n1432) );
  NANDN U1581 ( .A(n4488), .B(n1432), .Z(n1338) );
  NAND U1582 ( .A(n1339), .B(n1338), .Z(n1422) );
  XOR U1583 ( .A(n209), .B(a[19]), .Z(n1435) );
  OR U1584 ( .A(n1435), .B(n4612), .Z(n1342) );
  NAND U1585 ( .A(n1340), .B(n4669), .Z(n1341) );
  NAND U1586 ( .A(n1342), .B(n1341), .Z(n1420) );
  XOR U1587 ( .A(n4744), .B(a[17]), .Z(n1438) );
  NANDN U1588 ( .A(n1438), .B(n4745), .Z(n1345) );
  NANDN U1589 ( .A(n1343), .B(n4746), .Z(n1344) );
  AND U1590 ( .A(n1345), .B(n1344), .Z(n1421) );
  XOR U1591 ( .A(n1422), .B(n1423), .Z(n1448) );
  XNOR U1592 ( .A(n1447), .B(n1448), .Z(n1449) );
  XNOR U1593 ( .A(n1450), .B(n1449), .Z(n1397) );
  NANDN U1594 ( .A(n1347), .B(n1346), .Z(n1351) );
  NAND U1595 ( .A(n1349), .B(n1348), .Z(n1350) );
  NAND U1596 ( .A(n1351), .B(n1350), .Z(n1398) );
  XOR U1597 ( .A(n1397), .B(n1398), .Z(n1399) );
  XOR U1598 ( .A(n4859), .B(a[15]), .Z(n1405) );
  OR U1599 ( .A(n1405), .B(n4860), .Z(n1354) );
  NANDN U1600 ( .A(n1352), .B(n4915), .Z(n1353) );
  NAND U1601 ( .A(n1354), .B(n1353), .Z(n1417) );
  NANDN U1602 ( .A(n1355), .B(n4987), .Z(n1357) );
  XOR U1603 ( .A(n4909), .B(a[13]), .Z(n1408) );
  OR U1604 ( .A(n1408), .B(n4986), .Z(n1356) );
  NAND U1605 ( .A(n1357), .B(n1356), .Z(n1414) );
  XNOR U1606 ( .A(n210), .B(n1358), .Z(n1411) );
  OR U1607 ( .A(n1411), .B(n5095), .Z(n1361) );
  NANDN U1608 ( .A(n1359), .B(n5092), .Z(n1360) );
  AND U1609 ( .A(n1361), .B(n1360), .Z(n1415) );
  XNOR U1610 ( .A(n1414), .B(n1415), .Z(n1416) );
  XOR U1611 ( .A(n1417), .B(n1416), .Z(n1401) );
  XNOR U1612 ( .A(n1401), .B(n1402), .Z(n1404) );
  XOR U1613 ( .A(n1404), .B(n1403), .Z(n1400) );
  XNOR U1614 ( .A(n1399), .B(n1400), .Z(n1456) );
  NANDN U1615 ( .A(n1371), .B(n1370), .Z(n1375) );
  NANDN U1616 ( .A(n1373), .B(n1372), .Z(n1374) );
  NAND U1617 ( .A(n1375), .B(n1374), .Z(n1454) );
  NANDN U1618 ( .A(n1377), .B(n1376), .Z(n1381) );
  OR U1619 ( .A(n1379), .B(n1378), .Z(n1380) );
  AND U1620 ( .A(n1381), .B(n1380), .Z(n1453) );
  XNOR U1621 ( .A(n1454), .B(n1453), .Z(n1455) );
  XOR U1622 ( .A(n1456), .B(n1455), .Z(n1393) );
  NANDN U1623 ( .A(n1383), .B(n1382), .Z(n1387) );
  NAND U1624 ( .A(n1385), .B(n1384), .Z(n1386) );
  NAND U1625 ( .A(n1387), .B(n1386), .Z(n1394) );
  XOR U1626 ( .A(n1393), .B(n1394), .Z(n1395) );
  XOR U1627 ( .A(n1396), .B(n1395), .Z(n1459) );
  XNOR U1628 ( .A(n1459), .B(sreg[71]), .Z(n1461) );
  NAND U1629 ( .A(n1388), .B(sreg[70]), .Z(n1392) );
  OR U1630 ( .A(n1390), .B(n1389), .Z(n1391) );
  AND U1631 ( .A(n1392), .B(n1391), .Z(n1460) );
  XOR U1632 ( .A(n1461), .B(n1460), .Z(c[71]) );
  XNOR U1633 ( .A(n1527), .B(n1526), .Z(n1528) );
  XNOR U1634 ( .A(n4859), .B(n1852), .Z(n1482) );
  OR U1635 ( .A(n1482), .B(n4860), .Z(n1407) );
  NANDN U1636 ( .A(n1405), .B(n4915), .Z(n1406) );
  NAND U1637 ( .A(n1407), .B(n1406), .Z(n1494) );
  NANDN U1638 ( .A(n1408), .B(n4987), .Z(n1410) );
  XNOR U1639 ( .A(n4909), .B(n1705), .Z(n1485) );
  OR U1640 ( .A(n1485), .B(n4986), .Z(n1409) );
  NAND U1641 ( .A(n1410), .B(n1409), .Z(n1491) );
  XOR U1642 ( .A(n210), .B(a[10]), .Z(n1488) );
  OR U1643 ( .A(n1488), .B(n5095), .Z(n1413) );
  NANDN U1644 ( .A(n1411), .B(n5092), .Z(n1412) );
  AND U1645 ( .A(n1413), .B(n1412), .Z(n1492) );
  XOR U1646 ( .A(n1491), .B(n1492), .Z(n1493) );
  XOR U1647 ( .A(n1494), .B(n1493), .Z(n1476) );
  NANDN U1648 ( .A(n1415), .B(n1414), .Z(n1419) );
  NAND U1649 ( .A(n1417), .B(n1416), .Z(n1418) );
  NAND U1650 ( .A(n1419), .B(n1418), .Z(n1477) );
  XNOR U1651 ( .A(n1476), .B(n1477), .Z(n1478) );
  NANDN U1652 ( .A(n1421), .B(n1420), .Z(n1425) );
  NANDN U1653 ( .A(n1423), .B(n1422), .Z(n1424) );
  NAND U1654 ( .A(n1425), .B(n1424), .Z(n1479) );
  XOR U1655 ( .A(n1478), .B(n1479), .Z(n1473) );
  NAND U1656 ( .A(b[0]), .B(a[24]), .Z(n1426) );
  XNOR U1657 ( .A(b[1]), .B(n1426), .Z(n1428) );
  NAND U1658 ( .A(a[23]), .B(n206), .Z(n1427) );
  AND U1659 ( .A(n1428), .B(n1427), .Z(n1505) );
  XOR U1660 ( .A(n5129), .B(a[12]), .Z(n1511) );
  OR U1661 ( .A(n1511), .B(n5041), .Z(n1431) );
  NANDN U1662 ( .A(n1429), .B(n5052), .Z(n1430) );
  AND U1663 ( .A(n1431), .B(n1430), .Z(n1506) );
  XOR U1664 ( .A(n1505), .B(n1506), .Z(n1508) );
  NAND U1665 ( .A(b[15]), .B(a[8]), .Z(n1507) );
  XNOR U1666 ( .A(n1508), .B(n1507), .Z(n1504) );
  NAND U1667 ( .A(n4521), .B(n1432), .Z(n1434) );
  XOR U1668 ( .A(n208), .B(a[22]), .Z(n1517) );
  OR U1669 ( .A(n1517), .B(n4488), .Z(n1433) );
  NAND U1670 ( .A(n1434), .B(n1433), .Z(n1497) );
  XOR U1671 ( .A(b[5]), .B(a[20]), .Z(n1520) );
  NANDN U1672 ( .A(n4612), .B(n1520), .Z(n1437) );
  NANDN U1673 ( .A(n1435), .B(n4669), .Z(n1436) );
  NAND U1674 ( .A(n1437), .B(n1436), .Z(n1495) );
  XNOR U1675 ( .A(n4744), .B(n2003), .Z(n1523) );
  NANDN U1676 ( .A(n1523), .B(n4745), .Z(n1440) );
  NANDN U1677 ( .A(n1438), .B(n4746), .Z(n1439) );
  AND U1678 ( .A(n1440), .B(n1439), .Z(n1496) );
  XOR U1679 ( .A(n1497), .B(n1498), .Z(n1501) );
  NANDN U1680 ( .A(n1442), .B(n1441), .Z(n1446) );
  OR U1681 ( .A(n1444), .B(n1443), .Z(n1445) );
  NAND U1682 ( .A(n1446), .B(n1445), .Z(n1502) );
  XOR U1683 ( .A(n1501), .B(n1502), .Z(n1503) );
  XOR U1684 ( .A(n1504), .B(n1503), .Z(n1470) );
  NANDN U1685 ( .A(n1448), .B(n1447), .Z(n1452) );
  NAND U1686 ( .A(n1450), .B(n1449), .Z(n1451) );
  AND U1687 ( .A(n1452), .B(n1451), .Z(n1471) );
  XNOR U1688 ( .A(n1470), .B(n1471), .Z(n1472) );
  XNOR U1689 ( .A(n1473), .B(n1472), .Z(n1529) );
  XOR U1690 ( .A(n1528), .B(n1529), .Z(n1464) );
  NANDN U1691 ( .A(n1454), .B(n1453), .Z(n1458) );
  NANDN U1692 ( .A(n1456), .B(n1455), .Z(n1457) );
  NAND U1693 ( .A(n1458), .B(n1457), .Z(n1465) );
  XNOR U1694 ( .A(n1464), .B(n1465), .Z(n1466) );
  XNOR U1695 ( .A(n1467), .B(n1466), .Z(n1532) );
  XNOR U1696 ( .A(n1532), .B(sreg[72]), .Z(n1534) );
  NAND U1697 ( .A(n1459), .B(sreg[71]), .Z(n1463) );
  OR U1698 ( .A(n1461), .B(n1460), .Z(n1462) );
  AND U1699 ( .A(n1463), .B(n1462), .Z(n1533) );
  XOR U1700 ( .A(n1534), .B(n1533), .Z(c[72]) );
  NANDN U1701 ( .A(n1465), .B(n1464), .Z(n1469) );
  NAND U1702 ( .A(n1467), .B(n1466), .Z(n1468) );
  NAND U1703 ( .A(n1469), .B(n1468), .Z(n1540) );
  NANDN U1704 ( .A(n1471), .B(n1470), .Z(n1475) );
  NAND U1705 ( .A(n1473), .B(n1472), .Z(n1474) );
  NAND U1706 ( .A(n1475), .B(n1474), .Z(n1599) );
  NANDN U1707 ( .A(n1477), .B(n1476), .Z(n1481) );
  NANDN U1708 ( .A(n1479), .B(n1478), .Z(n1480) );
  NAND U1709 ( .A(n1481), .B(n1480), .Z(n1600) );
  XNOR U1710 ( .A(n1599), .B(n1600), .Z(n1601) );
  XOR U1711 ( .A(n4859), .B(a[17]), .Z(n1570) );
  OR U1712 ( .A(n1570), .B(n4860), .Z(n1484) );
  NANDN U1713 ( .A(n1482), .B(n4915), .Z(n1483) );
  NAND U1714 ( .A(n1484), .B(n1483), .Z(n1582) );
  NANDN U1715 ( .A(n1485), .B(n4987), .Z(n1487) );
  XOR U1716 ( .A(n4909), .B(a[15]), .Z(n1573) );
  OR U1717 ( .A(n1573), .B(n4986), .Z(n1486) );
  NAND U1718 ( .A(n1487), .B(n1486), .Z(n1579) );
  XOR U1719 ( .A(n210), .B(a[11]), .Z(n1576) );
  OR U1720 ( .A(n1576), .B(n5095), .Z(n1490) );
  NANDN U1721 ( .A(n1488), .B(n5092), .Z(n1489) );
  AND U1722 ( .A(n1490), .B(n1489), .Z(n1580) );
  XOR U1723 ( .A(n1579), .B(n1580), .Z(n1581) );
  XOR U1724 ( .A(n1582), .B(n1581), .Z(n1593) );
  XNOR U1725 ( .A(n1593), .B(n1594), .Z(n1595) );
  NANDN U1726 ( .A(n1496), .B(n1495), .Z(n1500) );
  NANDN U1727 ( .A(n1498), .B(n1497), .Z(n1499) );
  NAND U1728 ( .A(n1500), .B(n1499), .Z(n1596) );
  XOR U1729 ( .A(n1595), .B(n1596), .Z(n1590) );
  NANDN U1730 ( .A(n1506), .B(n1505), .Z(n1510) );
  OR U1731 ( .A(n1508), .B(n1507), .Z(n1509) );
  NAND U1732 ( .A(n1510), .B(n1509), .Z(n1567) );
  XOR U1733 ( .A(n5129), .B(a[13]), .Z(n1546) );
  OR U1734 ( .A(n1546), .B(n5041), .Z(n1513) );
  NANDN U1735 ( .A(n1511), .B(n5052), .Z(n1512) );
  AND U1736 ( .A(n1513), .B(n1512), .Z(n1559) );
  NAND U1737 ( .A(b[0]), .B(a[25]), .Z(n1514) );
  XNOR U1738 ( .A(b[1]), .B(n1514), .Z(n1516) );
  NAND U1739 ( .A(a[24]), .B(n206), .Z(n1515) );
  AND U1740 ( .A(n1516), .B(n1515), .Z(n1558) );
  XOR U1741 ( .A(n1559), .B(n1558), .Z(n1561) );
  NAND U1742 ( .A(a[9]), .B(b[15]), .Z(n1560) );
  XOR U1743 ( .A(n1561), .B(n1560), .Z(n1564) );
  NANDN U1744 ( .A(n1517), .B(n4521), .Z(n1519) );
  XOR U1745 ( .A(b[3]), .B(a[23]), .Z(n1549) );
  NANDN U1746 ( .A(n4488), .B(n1549), .Z(n1518) );
  AND U1747 ( .A(n1519), .B(n1518), .Z(n1585) );
  NAND U1748 ( .A(n4669), .B(n1520), .Z(n1522) );
  XOR U1749 ( .A(b[5]), .B(a[21]), .Z(n1552) );
  NANDN U1750 ( .A(n4612), .B(n1552), .Z(n1521) );
  AND U1751 ( .A(n1522), .B(n1521), .Z(n1583) );
  XOR U1752 ( .A(n4744), .B(a[19]), .Z(n1555) );
  NANDN U1753 ( .A(n1555), .B(n4745), .Z(n1525) );
  NANDN U1754 ( .A(n1523), .B(n4746), .Z(n1524) );
  AND U1755 ( .A(n1525), .B(n1524), .Z(n1584) );
  XOR U1756 ( .A(n1583), .B(n1584), .Z(n1586) );
  XOR U1757 ( .A(n1585), .B(n1586), .Z(n1565) );
  XNOR U1758 ( .A(n1564), .B(n1565), .Z(n1566) );
  XOR U1759 ( .A(n1567), .B(n1566), .Z(n1587) );
  XNOR U1760 ( .A(n1588), .B(n1587), .Z(n1589) );
  XNOR U1761 ( .A(n1590), .B(n1589), .Z(n1602) );
  XOR U1762 ( .A(n1601), .B(n1602), .Z(n1537) );
  NANDN U1763 ( .A(n1527), .B(n1526), .Z(n1531) );
  NANDN U1764 ( .A(n1529), .B(n1528), .Z(n1530) );
  NAND U1765 ( .A(n1531), .B(n1530), .Z(n1538) );
  XNOR U1766 ( .A(n1537), .B(n1538), .Z(n1539) );
  XNOR U1767 ( .A(n1540), .B(n1539), .Z(n1605) );
  XNOR U1768 ( .A(n1605), .B(sreg[73]), .Z(n1607) );
  NAND U1769 ( .A(n1532), .B(sreg[72]), .Z(n1536) );
  OR U1770 ( .A(n1534), .B(n1533), .Z(n1535) );
  AND U1771 ( .A(n1536), .B(n1535), .Z(n1606) );
  XOR U1772 ( .A(n1607), .B(n1606), .Z(c[73]) );
  NANDN U1773 ( .A(n1538), .B(n1537), .Z(n1542) );
  NAND U1774 ( .A(n1540), .B(n1539), .Z(n1541) );
  NAND U1775 ( .A(n1542), .B(n1541), .Z(n1613) );
  NAND U1776 ( .A(b[0]), .B(a[26]), .Z(n1543) );
  XNOR U1777 ( .A(b[1]), .B(n1543), .Z(n1545) );
  NAND U1778 ( .A(a[25]), .B(n206), .Z(n1544) );
  AND U1779 ( .A(n1545), .B(n1544), .Z(n1660) );
  XNOR U1780 ( .A(n5129), .B(n1705), .Z(n1648) );
  OR U1781 ( .A(n1648), .B(n5041), .Z(n1548) );
  NANDN U1782 ( .A(n1546), .B(n5052), .Z(n1547) );
  AND U1783 ( .A(n1548), .B(n1547), .Z(n1661) );
  XOR U1784 ( .A(n1660), .B(n1661), .Z(n1663) );
  NAND U1785 ( .A(b[15]), .B(a[10]), .Z(n1662) );
  XNOR U1786 ( .A(n1663), .B(n1662), .Z(n1666) );
  NAND U1787 ( .A(n1549), .B(n4521), .Z(n1551) );
  IV U1788 ( .A(a[24]), .Z(n2453) );
  XNOR U1789 ( .A(b[3]), .B(n2453), .Z(n1651) );
  NANDN U1790 ( .A(n4488), .B(n1651), .Z(n1550) );
  NAND U1791 ( .A(n1551), .B(n1550), .Z(n1642) );
  XOR U1792 ( .A(n209), .B(a[22]), .Z(n1654) );
  OR U1793 ( .A(n1654), .B(n4612), .Z(n1554) );
  NAND U1794 ( .A(n1552), .B(n4669), .Z(n1553) );
  NAND U1795 ( .A(n1554), .B(n1553), .Z(n1639) );
  XOR U1796 ( .A(n4744), .B(a[20]), .Z(n1657) );
  NANDN U1797 ( .A(n1657), .B(n4745), .Z(n1557) );
  NANDN U1798 ( .A(n1555), .B(n4746), .Z(n1556) );
  AND U1799 ( .A(n1557), .B(n1556), .Z(n1640) );
  XOR U1800 ( .A(n1642), .B(n1641), .Z(n1667) );
  XNOR U1801 ( .A(n1666), .B(n1667), .Z(n1668) );
  NANDN U1802 ( .A(n1559), .B(n1558), .Z(n1563) );
  OR U1803 ( .A(n1561), .B(n1560), .Z(n1562) );
  AND U1804 ( .A(n1563), .B(n1562), .Z(n1669) );
  XNOR U1805 ( .A(n1668), .B(n1669), .Z(n1615) );
  NANDN U1806 ( .A(n1565), .B(n1564), .Z(n1569) );
  NAND U1807 ( .A(n1567), .B(n1566), .Z(n1568) );
  AND U1808 ( .A(n1569), .B(n1568), .Z(n1614) );
  XNOR U1809 ( .A(n1615), .B(n1614), .Z(n1616) );
  XNOR U1810 ( .A(n4859), .B(n2003), .Z(n1624) );
  OR U1811 ( .A(n1624), .B(n4860), .Z(n1572) );
  NANDN U1812 ( .A(n1570), .B(n4915), .Z(n1571) );
  NAND U1813 ( .A(n1572), .B(n1571), .Z(n1636) );
  NANDN U1814 ( .A(n1573), .B(n4987), .Z(n1575) );
  XNOR U1815 ( .A(n4909), .B(n1852), .Z(n1627) );
  OR U1816 ( .A(n1627), .B(n4986), .Z(n1574) );
  NAND U1817 ( .A(n1575), .B(n1574), .Z(n1633) );
  XOR U1818 ( .A(n210), .B(a[12]), .Z(n1630) );
  OR U1819 ( .A(n1630), .B(n5095), .Z(n1578) );
  NANDN U1820 ( .A(n1576), .B(n5092), .Z(n1577) );
  AND U1821 ( .A(n1578), .B(n1577), .Z(n1634) );
  XNOR U1822 ( .A(n1633), .B(n1634), .Z(n1635) );
  XOR U1823 ( .A(n1636), .B(n1635), .Z(n1620) );
  XNOR U1824 ( .A(n1620), .B(n1621), .Z(n1623) );
  XOR U1825 ( .A(n1623), .B(n1622), .Z(n1617) );
  XOR U1826 ( .A(n1616), .B(n1617), .Z(n1674) );
  NANDN U1827 ( .A(n1588), .B(n1587), .Z(n1592) );
  NAND U1828 ( .A(n1590), .B(n1589), .Z(n1591) );
  NAND U1829 ( .A(n1592), .B(n1591), .Z(n1672) );
  NANDN U1830 ( .A(n1594), .B(n1593), .Z(n1598) );
  NANDN U1831 ( .A(n1596), .B(n1595), .Z(n1597) );
  NAND U1832 ( .A(n1598), .B(n1597), .Z(n1673) );
  XNOR U1833 ( .A(n1672), .B(n1673), .Z(n1675) );
  XOR U1834 ( .A(n1674), .B(n1675), .Z(n1610) );
  NANDN U1835 ( .A(n1600), .B(n1599), .Z(n1604) );
  NANDN U1836 ( .A(n1602), .B(n1601), .Z(n1603) );
  NAND U1837 ( .A(n1604), .B(n1603), .Z(n1611) );
  XOR U1838 ( .A(n1610), .B(n1611), .Z(n1612) );
  XOR U1839 ( .A(n1613), .B(n1612), .Z(n1676) );
  XNOR U1840 ( .A(n1676), .B(sreg[74]), .Z(n1678) );
  NAND U1841 ( .A(n1605), .B(sreg[73]), .Z(n1609) );
  OR U1842 ( .A(n1607), .B(n1606), .Z(n1608) );
  AND U1843 ( .A(n1609), .B(n1608), .Z(n1677) );
  XOR U1844 ( .A(n1678), .B(n1677), .Z(c[74]) );
  NANDN U1845 ( .A(n1615), .B(n1614), .Z(n1619) );
  NAND U1846 ( .A(n1617), .B(n1616), .Z(n1618) );
  NAND U1847 ( .A(n1619), .B(n1618), .Z(n1745) );
  XNOR U1848 ( .A(n1745), .B(n1744), .Z(n1746) );
  XOR U1849 ( .A(n4859), .B(a[19]), .Z(n1699) );
  OR U1850 ( .A(n1699), .B(n4860), .Z(n1626) );
  NANDN U1851 ( .A(n1624), .B(n4915), .Z(n1625) );
  NAND U1852 ( .A(n1626), .B(n1625), .Z(n1712) );
  NANDN U1853 ( .A(n1627), .B(n4987), .Z(n1629) );
  XOR U1854 ( .A(n4909), .B(a[17]), .Z(n1702) );
  OR U1855 ( .A(n1702), .B(n4986), .Z(n1628) );
  NAND U1856 ( .A(n1629), .B(n1628), .Z(n1709) );
  XOR U1857 ( .A(n210), .B(a[13]), .Z(n1706) );
  OR U1858 ( .A(n1706), .B(n5095), .Z(n1632) );
  NANDN U1859 ( .A(n1630), .B(n5092), .Z(n1631) );
  AND U1860 ( .A(n1632), .B(n1631), .Z(n1710) );
  XOR U1861 ( .A(n1709), .B(n1710), .Z(n1711) );
  XOR U1862 ( .A(n1712), .B(n1711), .Z(n1693) );
  NANDN U1863 ( .A(n1634), .B(n1633), .Z(n1638) );
  NAND U1864 ( .A(n1636), .B(n1635), .Z(n1637) );
  NAND U1865 ( .A(n1638), .B(n1637), .Z(n1694) );
  XNOR U1866 ( .A(n1693), .B(n1694), .Z(n1695) );
  NANDN U1867 ( .A(n1640), .B(n1639), .Z(n1644) );
  NAND U1868 ( .A(n1642), .B(n1641), .Z(n1643) );
  NAND U1869 ( .A(n1644), .B(n1643), .Z(n1696) );
  XOR U1870 ( .A(n1695), .B(n1696), .Z(n1690) );
  NAND U1871 ( .A(b[0]), .B(a[27]), .Z(n1645) );
  XNOR U1872 ( .A(b[1]), .B(n1645), .Z(n1647) );
  NAND U1873 ( .A(n206), .B(a[26]), .Z(n1646) );
  AND U1874 ( .A(n1647), .B(n1646), .Z(n1734) );
  XOR U1875 ( .A(n5129), .B(a[15]), .Z(n1722) );
  OR U1876 ( .A(n1722), .B(n5041), .Z(n1650) );
  NANDN U1877 ( .A(n1648), .B(n5052), .Z(n1649) );
  AND U1878 ( .A(n1650), .B(n1649), .Z(n1735) );
  XOR U1879 ( .A(n1734), .B(n1735), .Z(n1737) );
  NAND U1880 ( .A(b[15]), .B(a[11]), .Z(n1736) );
  XNOR U1881 ( .A(n1737), .B(n1736), .Z(n1743) );
  NAND U1882 ( .A(n4521), .B(n1651), .Z(n1653) );
  IV U1883 ( .A(a[25]), .Z(n2527) );
  XNOR U1884 ( .A(b[3]), .B(n2527), .Z(n1725) );
  NANDN U1885 ( .A(n4488), .B(n1725), .Z(n1652) );
  NAND U1886 ( .A(n1653), .B(n1652), .Z(n1715) );
  IV U1887 ( .A(a[23]), .Z(n2379) );
  XNOR U1888 ( .A(n209), .B(n2379), .Z(n1728) );
  OR U1889 ( .A(n1728), .B(n4612), .Z(n1656) );
  NANDN U1890 ( .A(n1654), .B(n4669), .Z(n1655) );
  NAND U1891 ( .A(n1656), .B(n1655), .Z(n1713) );
  XOR U1892 ( .A(n4744), .B(a[21]), .Z(n1731) );
  NANDN U1893 ( .A(n1731), .B(n4745), .Z(n1659) );
  NANDN U1894 ( .A(n1657), .B(n4746), .Z(n1658) );
  AND U1895 ( .A(n1659), .B(n1658), .Z(n1714) );
  XOR U1896 ( .A(n1715), .B(n1716), .Z(n1740) );
  NANDN U1897 ( .A(n1661), .B(n1660), .Z(n1665) );
  OR U1898 ( .A(n1663), .B(n1662), .Z(n1664) );
  NAND U1899 ( .A(n1665), .B(n1664), .Z(n1741) );
  XOR U1900 ( .A(n1740), .B(n1741), .Z(n1742) );
  XOR U1901 ( .A(n1743), .B(n1742), .Z(n1687) );
  NANDN U1902 ( .A(n1667), .B(n1666), .Z(n1671) );
  NAND U1903 ( .A(n1669), .B(n1668), .Z(n1670) );
  NAND U1904 ( .A(n1671), .B(n1670), .Z(n1688) );
  XNOR U1905 ( .A(n1687), .B(n1688), .Z(n1689) );
  XNOR U1906 ( .A(n1690), .B(n1689), .Z(n1747) );
  XOR U1907 ( .A(n1746), .B(n1747), .Z(n1681) );
  XNOR U1908 ( .A(n1681), .B(n1682), .Z(n1683) );
  XNOR U1909 ( .A(n1684), .B(n1683), .Z(n1750) );
  XNOR U1910 ( .A(n1750), .B(sreg[75]), .Z(n1752) );
  NAND U1911 ( .A(n1676), .B(sreg[74]), .Z(n1680) );
  OR U1912 ( .A(n1678), .B(n1677), .Z(n1679) );
  AND U1913 ( .A(n1680), .B(n1679), .Z(n1751) );
  XOR U1914 ( .A(n1752), .B(n1751), .Z(c[75]) );
  NANDN U1915 ( .A(n1682), .B(n1681), .Z(n1686) );
  NAND U1916 ( .A(n1684), .B(n1683), .Z(n1685) );
  NAND U1917 ( .A(n1686), .B(n1685), .Z(n1758) );
  NANDN U1918 ( .A(n1688), .B(n1687), .Z(n1692) );
  NAND U1919 ( .A(n1690), .B(n1689), .Z(n1691) );
  NAND U1920 ( .A(n1692), .B(n1691), .Z(n1817) );
  NANDN U1921 ( .A(n1694), .B(n1693), .Z(n1698) );
  NANDN U1922 ( .A(n1696), .B(n1695), .Z(n1697) );
  NAND U1923 ( .A(n1698), .B(n1697), .Z(n1818) );
  XNOR U1924 ( .A(n1817), .B(n1818), .Z(n1819) );
  XOR U1925 ( .A(n4859), .B(a[20]), .Z(n1773) );
  OR U1926 ( .A(n1773), .B(n4860), .Z(n1701) );
  NANDN U1927 ( .A(n1699), .B(n4915), .Z(n1700) );
  NAND U1928 ( .A(n1701), .B(n1700), .Z(n1785) );
  NANDN U1929 ( .A(n1702), .B(n4987), .Z(n1704) );
  XNOR U1930 ( .A(n4909), .B(n2003), .Z(n1776) );
  OR U1931 ( .A(n1776), .B(n4986), .Z(n1703) );
  NAND U1932 ( .A(n1704), .B(n1703), .Z(n1782) );
  XNOR U1933 ( .A(n210), .B(n1705), .Z(n1779) );
  OR U1934 ( .A(n1779), .B(n5095), .Z(n1708) );
  NANDN U1935 ( .A(n1706), .B(n5092), .Z(n1707) );
  AND U1936 ( .A(n1708), .B(n1707), .Z(n1783) );
  XOR U1937 ( .A(n1782), .B(n1783), .Z(n1784) );
  XOR U1938 ( .A(n1785), .B(n1784), .Z(n1767) );
  XNOR U1939 ( .A(n1767), .B(n1768), .Z(n1769) );
  NANDN U1940 ( .A(n1714), .B(n1713), .Z(n1718) );
  NANDN U1941 ( .A(n1716), .B(n1715), .Z(n1717) );
  NAND U1942 ( .A(n1718), .B(n1717), .Z(n1770) );
  XOR U1943 ( .A(n1769), .B(n1770), .Z(n1764) );
  NAND U1944 ( .A(b[0]), .B(a[28]), .Z(n1719) );
  XNOR U1945 ( .A(b[1]), .B(n1719), .Z(n1721) );
  NAND U1946 ( .A(a[27]), .B(n206), .Z(n1720) );
  AND U1947 ( .A(n1721), .B(n1720), .Z(n1807) );
  XNOR U1948 ( .A(n5129), .B(n1852), .Z(n1795) );
  OR U1949 ( .A(n1795), .B(n5041), .Z(n1724) );
  NANDN U1950 ( .A(n1722), .B(n5052), .Z(n1723) );
  AND U1951 ( .A(n1724), .B(n1723), .Z(n1808) );
  XOR U1952 ( .A(n1807), .B(n1808), .Z(n1810) );
  NAND U1953 ( .A(b[15]), .B(a[12]), .Z(n1809) );
  XNOR U1954 ( .A(n1810), .B(n1809), .Z(n1816) );
  NAND U1955 ( .A(n4521), .B(n1725), .Z(n1727) );
  XOR U1956 ( .A(b[3]), .B(a[26]), .Z(n1798) );
  NANDN U1957 ( .A(n4488), .B(n1798), .Z(n1726) );
  NAND U1958 ( .A(n1727), .B(n1726), .Z(n1788) );
  XNOR U1959 ( .A(n209), .B(n2453), .Z(n1801) );
  OR U1960 ( .A(n1801), .B(n4612), .Z(n1730) );
  NANDN U1961 ( .A(n1728), .B(n4669), .Z(n1729) );
  NAND U1962 ( .A(n1730), .B(n1729), .Z(n1786) );
  XOR U1963 ( .A(n4744), .B(a[22]), .Z(n1804) );
  NANDN U1964 ( .A(n1804), .B(n4745), .Z(n1733) );
  NANDN U1965 ( .A(n1731), .B(n4746), .Z(n1732) );
  AND U1966 ( .A(n1733), .B(n1732), .Z(n1787) );
  XOR U1967 ( .A(n1788), .B(n1789), .Z(n1813) );
  NANDN U1968 ( .A(n1735), .B(n1734), .Z(n1739) );
  OR U1969 ( .A(n1737), .B(n1736), .Z(n1738) );
  NAND U1970 ( .A(n1739), .B(n1738), .Z(n1814) );
  XOR U1971 ( .A(n1813), .B(n1814), .Z(n1815) );
  XOR U1972 ( .A(n1816), .B(n1815), .Z(n1761) );
  XNOR U1973 ( .A(n1761), .B(n1762), .Z(n1763) );
  XNOR U1974 ( .A(n1764), .B(n1763), .Z(n1820) );
  XOR U1975 ( .A(n1819), .B(n1820), .Z(n1755) );
  NANDN U1976 ( .A(n1745), .B(n1744), .Z(n1749) );
  NANDN U1977 ( .A(n1747), .B(n1746), .Z(n1748) );
  NAND U1978 ( .A(n1749), .B(n1748), .Z(n1756) );
  XNOR U1979 ( .A(n1755), .B(n1756), .Z(n1757) );
  XNOR U1980 ( .A(n1758), .B(n1757), .Z(n1823) );
  XNOR U1981 ( .A(n1823), .B(sreg[76]), .Z(n1825) );
  NAND U1982 ( .A(n1750), .B(sreg[75]), .Z(n1754) );
  OR U1983 ( .A(n1752), .B(n1751), .Z(n1753) );
  AND U1984 ( .A(n1754), .B(n1753), .Z(n1824) );
  XOR U1985 ( .A(n1825), .B(n1824), .Z(c[76]) );
  NANDN U1986 ( .A(n1756), .B(n1755), .Z(n1760) );
  NAND U1987 ( .A(n1758), .B(n1757), .Z(n1759) );
  NAND U1988 ( .A(n1760), .B(n1759), .Z(n1831) );
  NANDN U1989 ( .A(n1762), .B(n1761), .Z(n1766) );
  NAND U1990 ( .A(n1764), .B(n1763), .Z(n1765) );
  NAND U1991 ( .A(n1766), .B(n1765), .Z(n1893) );
  NANDN U1992 ( .A(n1768), .B(n1767), .Z(n1772) );
  NANDN U1993 ( .A(n1770), .B(n1769), .Z(n1771) );
  NAND U1994 ( .A(n1772), .B(n1771), .Z(n1894) );
  XNOR U1995 ( .A(n1893), .B(n1894), .Z(n1895) );
  XOR U1996 ( .A(n4859), .B(a[21]), .Z(n1846) );
  OR U1997 ( .A(n1846), .B(n4860), .Z(n1775) );
  NANDN U1998 ( .A(n1773), .B(n4915), .Z(n1774) );
  NAND U1999 ( .A(n1775), .B(n1774), .Z(n1859) );
  NANDN U2000 ( .A(n1776), .B(n4987), .Z(n1778) );
  XOR U2001 ( .A(n4909), .B(a[19]), .Z(n1849) );
  OR U2002 ( .A(n1849), .B(n4986), .Z(n1777) );
  NAND U2003 ( .A(n1778), .B(n1777), .Z(n1856) );
  XOR U2004 ( .A(n210), .B(a[15]), .Z(n1853) );
  OR U2005 ( .A(n1853), .B(n5095), .Z(n1781) );
  NANDN U2006 ( .A(n1779), .B(n5092), .Z(n1780) );
  AND U2007 ( .A(n1781), .B(n1780), .Z(n1857) );
  XOR U2008 ( .A(n1856), .B(n1857), .Z(n1858) );
  XOR U2009 ( .A(n1859), .B(n1858), .Z(n1840) );
  XNOR U2010 ( .A(n1840), .B(n1841), .Z(n1842) );
  NANDN U2011 ( .A(n1787), .B(n1786), .Z(n1791) );
  NANDN U2012 ( .A(n1789), .B(n1788), .Z(n1790) );
  NAND U2013 ( .A(n1791), .B(n1790), .Z(n1843) );
  XOR U2014 ( .A(n1842), .B(n1843), .Z(n1837) );
  NAND U2015 ( .A(b[0]), .B(a[29]), .Z(n1792) );
  XNOR U2016 ( .A(b[1]), .B(n1792), .Z(n1794) );
  NAND U2017 ( .A(a[28]), .B(n206), .Z(n1793) );
  AND U2018 ( .A(n1794), .B(n1793), .Z(n1872) );
  XOR U2019 ( .A(n5129), .B(a[17]), .Z(n1881) );
  OR U2020 ( .A(n1881), .B(n5041), .Z(n1797) );
  NANDN U2021 ( .A(n1795), .B(n5052), .Z(n1796) );
  AND U2022 ( .A(n1797), .B(n1796), .Z(n1873) );
  XOR U2023 ( .A(n1872), .B(n1873), .Z(n1875) );
  NAND U2024 ( .A(b[15]), .B(a[13]), .Z(n1874) );
  XNOR U2025 ( .A(n1875), .B(n1874), .Z(n1866) );
  NAND U2026 ( .A(n4521), .B(n1798), .Z(n1800) );
  IV U2027 ( .A(a[27]), .Z(n2664) );
  XNOR U2028 ( .A(b[3]), .B(n2664), .Z(n1884) );
  NANDN U2029 ( .A(n4488), .B(n1884), .Z(n1799) );
  NAND U2030 ( .A(n1800), .B(n1799), .Z(n1863) );
  XNOR U2031 ( .A(n209), .B(n2527), .Z(n1887) );
  OR U2032 ( .A(n1887), .B(n4612), .Z(n1803) );
  NANDN U2033 ( .A(n1801), .B(n4669), .Z(n1802) );
  NAND U2034 ( .A(n1803), .B(n1802), .Z(n1860) );
  XNOR U2035 ( .A(n4744), .B(n2379), .Z(n1890) );
  NANDN U2036 ( .A(n1890), .B(n4745), .Z(n1806) );
  NANDN U2037 ( .A(n1804), .B(n4746), .Z(n1805) );
  AND U2038 ( .A(n1806), .B(n1805), .Z(n1861) );
  XOR U2039 ( .A(n1863), .B(n1862), .Z(n1867) );
  XNOR U2040 ( .A(n1866), .B(n1867), .Z(n1868) );
  NANDN U2041 ( .A(n1808), .B(n1807), .Z(n1812) );
  OR U2042 ( .A(n1810), .B(n1809), .Z(n1811) );
  NAND U2043 ( .A(n1812), .B(n1811), .Z(n1869) );
  XOR U2044 ( .A(n1868), .B(n1869), .Z(n1834) );
  XNOR U2045 ( .A(n1834), .B(n1835), .Z(n1836) );
  XNOR U2046 ( .A(n1837), .B(n1836), .Z(n1896) );
  XOR U2047 ( .A(n1895), .B(n1896), .Z(n1828) );
  NANDN U2048 ( .A(n1818), .B(n1817), .Z(n1822) );
  NANDN U2049 ( .A(n1820), .B(n1819), .Z(n1821) );
  NAND U2050 ( .A(n1822), .B(n1821), .Z(n1829) );
  XNOR U2051 ( .A(n1828), .B(n1829), .Z(n1830) );
  XNOR U2052 ( .A(n1831), .B(n1830), .Z(n1899) );
  XNOR U2053 ( .A(n1899), .B(sreg[77]), .Z(n1901) );
  NAND U2054 ( .A(n1823), .B(sreg[76]), .Z(n1827) );
  OR U2055 ( .A(n1825), .B(n1824), .Z(n1826) );
  AND U2056 ( .A(n1827), .B(n1826), .Z(n1900) );
  XOR U2057 ( .A(n1901), .B(n1900), .Z(c[77]) );
  NANDN U2058 ( .A(n1829), .B(n1828), .Z(n1833) );
  NAND U2059 ( .A(n1831), .B(n1830), .Z(n1832) );
  NAND U2060 ( .A(n1833), .B(n1832), .Z(n1907) );
  NANDN U2061 ( .A(n1835), .B(n1834), .Z(n1839) );
  NAND U2062 ( .A(n1837), .B(n1836), .Z(n1838) );
  NAND U2063 ( .A(n1839), .B(n1838), .Z(n1968) );
  NANDN U2064 ( .A(n1841), .B(n1840), .Z(n1845) );
  NANDN U2065 ( .A(n1843), .B(n1842), .Z(n1844) );
  NAND U2066 ( .A(n1845), .B(n1844), .Z(n1969) );
  XNOR U2067 ( .A(n1968), .B(n1969), .Z(n1970) );
  XOR U2068 ( .A(n4859), .B(a[22]), .Z(n1922) );
  OR U2069 ( .A(n1922), .B(n4860), .Z(n1848) );
  NANDN U2070 ( .A(n1846), .B(n4915), .Z(n1847) );
  NAND U2071 ( .A(n1848), .B(n1847), .Z(n1934) );
  NANDN U2072 ( .A(n1849), .B(n4987), .Z(n1851) );
  XOR U2073 ( .A(n4909), .B(a[20]), .Z(n1925) );
  OR U2074 ( .A(n1925), .B(n4986), .Z(n1850) );
  NAND U2075 ( .A(n1851), .B(n1850), .Z(n1931) );
  XNOR U2076 ( .A(n210), .B(n1852), .Z(n1928) );
  OR U2077 ( .A(n1928), .B(n5095), .Z(n1855) );
  NANDN U2078 ( .A(n1853), .B(n5092), .Z(n1854) );
  AND U2079 ( .A(n1855), .B(n1854), .Z(n1932) );
  XOR U2080 ( .A(n1931), .B(n1932), .Z(n1933) );
  XOR U2081 ( .A(n1934), .B(n1933), .Z(n1916) );
  XNOR U2082 ( .A(n1916), .B(n1917), .Z(n1918) );
  NANDN U2083 ( .A(n1861), .B(n1860), .Z(n1865) );
  NAND U2084 ( .A(n1863), .B(n1862), .Z(n1864) );
  NAND U2085 ( .A(n1865), .B(n1864), .Z(n1919) );
  XOR U2086 ( .A(n1918), .B(n1919), .Z(n1913) );
  NANDN U2087 ( .A(n1867), .B(n1866), .Z(n1871) );
  NANDN U2088 ( .A(n1869), .B(n1868), .Z(n1870) );
  NAND U2089 ( .A(n1871), .B(n1870), .Z(n1911) );
  NANDN U2090 ( .A(n1873), .B(n1872), .Z(n1877) );
  OR U2091 ( .A(n1875), .B(n1874), .Z(n1876) );
  NAND U2092 ( .A(n1877), .B(n1876), .Z(n1942) );
  NAND U2093 ( .A(b[0]), .B(a[30]), .Z(n1878) );
  XNOR U2094 ( .A(b[1]), .B(n1878), .Z(n1880) );
  NAND U2095 ( .A(a[29]), .B(n206), .Z(n1879) );
  AND U2096 ( .A(n1880), .B(n1879), .Z(n1962) );
  XNOR U2097 ( .A(n5129), .B(n2003), .Z(n1950) );
  OR U2098 ( .A(n1950), .B(n5041), .Z(n1883) );
  NANDN U2099 ( .A(n1881), .B(n5052), .Z(n1882) );
  AND U2100 ( .A(n1883), .B(n1882), .Z(n1963) );
  XOR U2101 ( .A(n1962), .B(n1963), .Z(n1965) );
  NAND U2102 ( .A(a[14]), .B(b[15]), .Z(n1964) );
  XOR U2103 ( .A(n1965), .B(n1964), .Z(n1941) );
  XNOR U2104 ( .A(n1942), .B(n1941), .Z(n1943) );
  NAND U2105 ( .A(n4521), .B(n1884), .Z(n1886) );
  IV U2106 ( .A(a[28]), .Z(n2738) );
  XNOR U2107 ( .A(b[3]), .B(n2738), .Z(n1953) );
  NANDN U2108 ( .A(n4488), .B(n1953), .Z(n1885) );
  NAND U2109 ( .A(n1886), .B(n1885), .Z(n1937) );
  XOR U2110 ( .A(n209), .B(a[26]), .Z(n1956) );
  OR U2111 ( .A(n1956), .B(n4612), .Z(n1889) );
  NANDN U2112 ( .A(n1887), .B(n4669), .Z(n1888) );
  NAND U2113 ( .A(n1889), .B(n1888), .Z(n1935) );
  XNOR U2114 ( .A(n4744), .B(n2453), .Z(n1959) );
  NANDN U2115 ( .A(n1959), .B(n4745), .Z(n1892) );
  NANDN U2116 ( .A(n1890), .B(n4746), .Z(n1891) );
  AND U2117 ( .A(n1892), .B(n1891), .Z(n1936) );
  XOR U2118 ( .A(n1937), .B(n1938), .Z(n1944) );
  XOR U2119 ( .A(n1943), .B(n1944), .Z(n1910) );
  XNOR U2120 ( .A(n1911), .B(n1910), .Z(n1912) );
  XNOR U2121 ( .A(n1913), .B(n1912), .Z(n1971) );
  XOR U2122 ( .A(n1970), .B(n1971), .Z(n1904) );
  NANDN U2123 ( .A(n1894), .B(n1893), .Z(n1898) );
  NANDN U2124 ( .A(n1896), .B(n1895), .Z(n1897) );
  NAND U2125 ( .A(n1898), .B(n1897), .Z(n1905) );
  XNOR U2126 ( .A(n1904), .B(n1905), .Z(n1906) );
  XNOR U2127 ( .A(n1907), .B(n1906), .Z(n1974) );
  XNOR U2128 ( .A(n1974), .B(sreg[78]), .Z(n1976) );
  NAND U2129 ( .A(n1899), .B(sreg[77]), .Z(n1903) );
  OR U2130 ( .A(n1901), .B(n1900), .Z(n1902) );
  AND U2131 ( .A(n1903), .B(n1902), .Z(n1975) );
  XOR U2132 ( .A(n1976), .B(n1975), .Z(c[78]) );
  NANDN U2133 ( .A(n1905), .B(n1904), .Z(n1909) );
  NAND U2134 ( .A(n1907), .B(n1906), .Z(n1908) );
  NAND U2135 ( .A(n1909), .B(n1908), .Z(n1982) );
  NANDN U2136 ( .A(n1911), .B(n1910), .Z(n1915) );
  NAND U2137 ( .A(n1913), .B(n1912), .Z(n1914) );
  NAND U2138 ( .A(n1915), .B(n1914), .Z(n2044) );
  NANDN U2139 ( .A(n1917), .B(n1916), .Z(n1921) );
  NANDN U2140 ( .A(n1919), .B(n1918), .Z(n1920) );
  NAND U2141 ( .A(n1921), .B(n1920), .Z(n2045) );
  XNOR U2142 ( .A(n2044), .B(n2045), .Z(n2046) );
  XNOR U2143 ( .A(n4859), .B(n2379), .Z(n1997) );
  OR U2144 ( .A(n1997), .B(n4860), .Z(n1924) );
  NANDN U2145 ( .A(n1922), .B(n4915), .Z(n1923) );
  NAND U2146 ( .A(n1924), .B(n1923), .Z(n2010) );
  NANDN U2147 ( .A(n1925), .B(n4987), .Z(n1927) );
  XOR U2148 ( .A(n4909), .B(a[21]), .Z(n2000) );
  OR U2149 ( .A(n2000), .B(n4986), .Z(n1926) );
  NAND U2150 ( .A(n1927), .B(n1926), .Z(n2007) );
  XOR U2151 ( .A(n210), .B(a[17]), .Z(n2004) );
  OR U2152 ( .A(n2004), .B(n5095), .Z(n1930) );
  NANDN U2153 ( .A(n1928), .B(n5092), .Z(n1929) );
  AND U2154 ( .A(n1930), .B(n1929), .Z(n2008) );
  XOR U2155 ( .A(n2007), .B(n2008), .Z(n2009) );
  XOR U2156 ( .A(n2010), .B(n2009), .Z(n1991) );
  XNOR U2157 ( .A(n1991), .B(n1992), .Z(n1993) );
  NANDN U2158 ( .A(n1936), .B(n1935), .Z(n1940) );
  NANDN U2159 ( .A(n1938), .B(n1937), .Z(n1939) );
  NAND U2160 ( .A(n1940), .B(n1939), .Z(n1994) );
  XOR U2161 ( .A(n1993), .B(n1994), .Z(n1988) );
  NAND U2162 ( .A(n1942), .B(n1941), .Z(n1946) );
  OR U2163 ( .A(n1944), .B(n1943), .Z(n1945) );
  NAND U2164 ( .A(n1946), .B(n1945), .Z(n1985) );
  NAND U2165 ( .A(b[0]), .B(a[31]), .Z(n1947) );
  XNOR U2166 ( .A(b[1]), .B(n1947), .Z(n1949) );
  NAND U2167 ( .A(n206), .B(a[30]), .Z(n1948) );
  AND U2168 ( .A(n1949), .B(n1948), .Z(n2023) );
  XOR U2169 ( .A(n5129), .B(a[19]), .Z(n2032) );
  OR U2170 ( .A(n2032), .B(n5041), .Z(n1952) );
  NANDN U2171 ( .A(n1950), .B(n5052), .Z(n1951) );
  AND U2172 ( .A(n1952), .B(n1951), .Z(n2024) );
  XOR U2173 ( .A(n2023), .B(n2024), .Z(n2026) );
  NAND U2174 ( .A(b[15]), .B(a[15]), .Z(n2025) );
  XNOR U2175 ( .A(n2026), .B(n2025), .Z(n2020) );
  NAND U2176 ( .A(n4521), .B(n1953), .Z(n1955) );
  IV U2177 ( .A(a[29]), .Z(n2822) );
  XNOR U2178 ( .A(b[3]), .B(n2822), .Z(n2035) );
  NANDN U2179 ( .A(n4488), .B(n2035), .Z(n1954) );
  NAND U2180 ( .A(n1955), .B(n1954), .Z(n2013) );
  XNOR U2181 ( .A(n209), .B(n2664), .Z(n2038) );
  OR U2182 ( .A(n2038), .B(n4612), .Z(n1958) );
  NANDN U2183 ( .A(n1956), .B(n4669), .Z(n1957) );
  NAND U2184 ( .A(n1958), .B(n1957), .Z(n2011) );
  XNOR U2185 ( .A(n4744), .B(n2527), .Z(n2041) );
  NANDN U2186 ( .A(n2041), .B(n4745), .Z(n1961) );
  NANDN U2187 ( .A(n1959), .B(n4746), .Z(n1960) );
  AND U2188 ( .A(n1961), .B(n1960), .Z(n2012) );
  XOR U2189 ( .A(n2013), .B(n2014), .Z(n2017) );
  NANDN U2190 ( .A(n1963), .B(n1962), .Z(n1967) );
  OR U2191 ( .A(n1965), .B(n1964), .Z(n1966) );
  NAND U2192 ( .A(n1967), .B(n1966), .Z(n2018) );
  XNOR U2193 ( .A(n2017), .B(n2018), .Z(n2019) );
  XOR U2194 ( .A(n2020), .B(n2019), .Z(n1986) );
  XNOR U2195 ( .A(n1985), .B(n1986), .Z(n1987) );
  XNOR U2196 ( .A(n1988), .B(n1987), .Z(n2047) );
  XOR U2197 ( .A(n2046), .B(n2047), .Z(n1979) );
  NANDN U2198 ( .A(n1969), .B(n1968), .Z(n1973) );
  NANDN U2199 ( .A(n1971), .B(n1970), .Z(n1972) );
  NAND U2200 ( .A(n1973), .B(n1972), .Z(n1980) );
  XNOR U2201 ( .A(n1979), .B(n1980), .Z(n1981) );
  XNOR U2202 ( .A(n1982), .B(n1981), .Z(n2050) );
  XNOR U2203 ( .A(n2050), .B(sreg[79]), .Z(n2052) );
  NAND U2204 ( .A(n1974), .B(sreg[78]), .Z(n1978) );
  OR U2205 ( .A(n1976), .B(n1975), .Z(n1977) );
  AND U2206 ( .A(n1978), .B(n1977), .Z(n2051) );
  XOR U2207 ( .A(n2052), .B(n2051), .Z(c[79]) );
  NANDN U2208 ( .A(n1980), .B(n1979), .Z(n1984) );
  NAND U2209 ( .A(n1982), .B(n1981), .Z(n1983) );
  NAND U2210 ( .A(n1984), .B(n1983), .Z(n2058) );
  NANDN U2211 ( .A(n1986), .B(n1985), .Z(n1990) );
  NAND U2212 ( .A(n1988), .B(n1987), .Z(n1989) );
  NAND U2213 ( .A(n1990), .B(n1989), .Z(n2119) );
  NANDN U2214 ( .A(n1992), .B(n1991), .Z(n1996) );
  NANDN U2215 ( .A(n1994), .B(n1993), .Z(n1995) );
  NAND U2216 ( .A(n1996), .B(n1995), .Z(n2120) );
  XNOR U2217 ( .A(n2119), .B(n2120), .Z(n2121) );
  XNOR U2218 ( .A(n4859), .B(n2453), .Z(n2073) );
  OR U2219 ( .A(n2073), .B(n4860), .Z(n1999) );
  NANDN U2220 ( .A(n1997), .B(n4915), .Z(n1998) );
  NAND U2221 ( .A(n1999), .B(n1998), .Z(n2085) );
  NANDN U2222 ( .A(n2000), .B(n4987), .Z(n2002) );
  XOR U2223 ( .A(n4909), .B(a[22]), .Z(n2076) );
  OR U2224 ( .A(n2076), .B(n4986), .Z(n2001) );
  NAND U2225 ( .A(n2002), .B(n2001), .Z(n2082) );
  XNOR U2226 ( .A(n210), .B(n2003), .Z(n2079) );
  OR U2227 ( .A(n2079), .B(n5095), .Z(n2006) );
  NANDN U2228 ( .A(n2004), .B(n5092), .Z(n2005) );
  AND U2229 ( .A(n2006), .B(n2005), .Z(n2083) );
  XOR U2230 ( .A(n2082), .B(n2083), .Z(n2084) );
  XOR U2231 ( .A(n2085), .B(n2084), .Z(n2067) );
  XNOR U2232 ( .A(n2067), .B(n2068), .Z(n2069) );
  NANDN U2233 ( .A(n2012), .B(n2011), .Z(n2016) );
  NANDN U2234 ( .A(n2014), .B(n2013), .Z(n2015) );
  NAND U2235 ( .A(n2016), .B(n2015), .Z(n2070) );
  XOR U2236 ( .A(n2069), .B(n2070), .Z(n2064) );
  NANDN U2237 ( .A(n2018), .B(n2017), .Z(n2022) );
  NAND U2238 ( .A(n2020), .B(n2019), .Z(n2021) );
  NAND U2239 ( .A(n2022), .B(n2021), .Z(n2062) );
  NANDN U2240 ( .A(n2024), .B(n2023), .Z(n2028) );
  OR U2241 ( .A(n2026), .B(n2025), .Z(n2027) );
  NAND U2242 ( .A(n2028), .B(n2027), .Z(n2095) );
  NAND U2243 ( .A(b[0]), .B(a[32]), .Z(n2029) );
  XNOR U2244 ( .A(b[1]), .B(n2029), .Z(n2031) );
  NAND U2245 ( .A(a[31]), .B(n206), .Z(n2030) );
  AND U2246 ( .A(n2031), .B(n2030), .Z(n2113) );
  XOR U2247 ( .A(n5129), .B(a[20]), .Z(n2101) );
  OR U2248 ( .A(n2101), .B(n5041), .Z(n2034) );
  NANDN U2249 ( .A(n2032), .B(n5052), .Z(n2033) );
  AND U2250 ( .A(n2034), .B(n2033), .Z(n2114) );
  XOR U2251 ( .A(n2113), .B(n2114), .Z(n2116) );
  NAND U2252 ( .A(a[16]), .B(b[15]), .Z(n2115) );
  XOR U2253 ( .A(n2116), .B(n2115), .Z(n2092) );
  NAND U2254 ( .A(n4521), .B(n2035), .Z(n2037) );
  XOR U2255 ( .A(b[3]), .B(a[30]), .Z(n2104) );
  NANDN U2256 ( .A(n4488), .B(n2104), .Z(n2036) );
  NAND U2257 ( .A(n2037), .B(n2036), .Z(n2088) );
  XNOR U2258 ( .A(n209), .B(n2738), .Z(n2107) );
  OR U2259 ( .A(n2107), .B(n4612), .Z(n2040) );
  NANDN U2260 ( .A(n2038), .B(n4669), .Z(n2039) );
  NAND U2261 ( .A(n2040), .B(n2039), .Z(n2086) );
  XOR U2262 ( .A(n4744), .B(a[26]), .Z(n2110) );
  NANDN U2263 ( .A(n2110), .B(n4745), .Z(n2043) );
  NANDN U2264 ( .A(n2041), .B(n4746), .Z(n2042) );
  AND U2265 ( .A(n2043), .B(n2042), .Z(n2087) );
  XOR U2266 ( .A(n2088), .B(n2089), .Z(n2093) );
  XNOR U2267 ( .A(n2092), .B(n2093), .Z(n2094) );
  XOR U2268 ( .A(n2095), .B(n2094), .Z(n2061) );
  XNOR U2269 ( .A(n2062), .B(n2061), .Z(n2063) );
  XNOR U2270 ( .A(n2064), .B(n2063), .Z(n2122) );
  XOR U2271 ( .A(n2121), .B(n2122), .Z(n2055) );
  NANDN U2272 ( .A(n2045), .B(n2044), .Z(n2049) );
  NANDN U2273 ( .A(n2047), .B(n2046), .Z(n2048) );
  NAND U2274 ( .A(n2049), .B(n2048), .Z(n2056) );
  XNOR U2275 ( .A(n2055), .B(n2056), .Z(n2057) );
  XNOR U2276 ( .A(n2058), .B(n2057), .Z(n2125) );
  XNOR U2277 ( .A(n2125), .B(sreg[80]), .Z(n2127) );
  NAND U2278 ( .A(n2050), .B(sreg[79]), .Z(n2054) );
  OR U2279 ( .A(n2052), .B(n2051), .Z(n2053) );
  AND U2280 ( .A(n2054), .B(n2053), .Z(n2126) );
  XOR U2281 ( .A(n2127), .B(n2126), .Z(c[80]) );
  NANDN U2282 ( .A(n2056), .B(n2055), .Z(n2060) );
  NAND U2283 ( .A(n2058), .B(n2057), .Z(n2059) );
  NAND U2284 ( .A(n2060), .B(n2059), .Z(n2133) );
  NANDN U2285 ( .A(n2062), .B(n2061), .Z(n2066) );
  NAND U2286 ( .A(n2064), .B(n2063), .Z(n2065) );
  NAND U2287 ( .A(n2066), .B(n2065), .Z(n2194) );
  NANDN U2288 ( .A(n2068), .B(n2067), .Z(n2072) );
  NANDN U2289 ( .A(n2070), .B(n2069), .Z(n2071) );
  NAND U2290 ( .A(n2072), .B(n2071), .Z(n2195) );
  XNOR U2291 ( .A(n2194), .B(n2195), .Z(n2196) );
  XNOR U2292 ( .A(n4859), .B(n2527), .Z(n2148) );
  OR U2293 ( .A(n2148), .B(n4860), .Z(n2075) );
  NANDN U2294 ( .A(n2073), .B(n4915), .Z(n2074) );
  NAND U2295 ( .A(n2075), .B(n2074), .Z(n2160) );
  NANDN U2296 ( .A(n2076), .B(n4987), .Z(n2078) );
  XNOR U2297 ( .A(n4909), .B(n2379), .Z(n2151) );
  OR U2298 ( .A(n2151), .B(n4986), .Z(n2077) );
  NAND U2299 ( .A(n2078), .B(n2077), .Z(n2157) );
  XOR U2300 ( .A(n210), .B(a[19]), .Z(n2154) );
  OR U2301 ( .A(n2154), .B(n5095), .Z(n2081) );
  NANDN U2302 ( .A(n2079), .B(n5092), .Z(n2080) );
  AND U2303 ( .A(n2081), .B(n2080), .Z(n2158) );
  XOR U2304 ( .A(n2157), .B(n2158), .Z(n2159) );
  XOR U2305 ( .A(n2160), .B(n2159), .Z(n2142) );
  XNOR U2306 ( .A(n2142), .B(n2143), .Z(n2144) );
  NANDN U2307 ( .A(n2087), .B(n2086), .Z(n2091) );
  NANDN U2308 ( .A(n2089), .B(n2088), .Z(n2090) );
  NAND U2309 ( .A(n2091), .B(n2090), .Z(n2145) );
  XOR U2310 ( .A(n2144), .B(n2145), .Z(n2139) );
  NANDN U2311 ( .A(n2093), .B(n2092), .Z(n2097) );
  NAND U2312 ( .A(n2095), .B(n2094), .Z(n2096) );
  NAND U2313 ( .A(n2097), .B(n2096), .Z(n2136) );
  NAND U2314 ( .A(b[0]), .B(a[33]), .Z(n2098) );
  XNOR U2315 ( .A(b[1]), .B(n2098), .Z(n2100) );
  NAND U2316 ( .A(a[32]), .B(n206), .Z(n2099) );
  AND U2317 ( .A(n2100), .B(n2099), .Z(n2167) );
  XOR U2318 ( .A(n5129), .B(a[21]), .Z(n2173) );
  OR U2319 ( .A(n2173), .B(n5041), .Z(n2103) );
  NANDN U2320 ( .A(n2101), .B(n5052), .Z(n2102) );
  AND U2321 ( .A(n2103), .B(n2102), .Z(n2168) );
  XOR U2322 ( .A(n2167), .B(n2168), .Z(n2170) );
  NAND U2323 ( .A(b[15]), .B(a[17]), .Z(n2169) );
  XNOR U2324 ( .A(n2170), .B(n2169), .Z(n2191) );
  NAND U2325 ( .A(n4521), .B(n2104), .Z(n2106) );
  IV U2326 ( .A(a[31]), .Z(n2971) );
  XNOR U2327 ( .A(b[3]), .B(n2971), .Z(n2179) );
  NANDN U2328 ( .A(n4488), .B(n2179), .Z(n2105) );
  NAND U2329 ( .A(n2106), .B(n2105), .Z(n2163) );
  XNOR U2330 ( .A(n209), .B(n2822), .Z(n2182) );
  OR U2331 ( .A(n2182), .B(n4612), .Z(n2109) );
  NANDN U2332 ( .A(n2107), .B(n4669), .Z(n2108) );
  NAND U2333 ( .A(n2109), .B(n2108), .Z(n2161) );
  XNOR U2334 ( .A(n4744), .B(n2664), .Z(n2185) );
  NANDN U2335 ( .A(n2185), .B(n4745), .Z(n2112) );
  NANDN U2336 ( .A(n2110), .B(n4746), .Z(n2111) );
  AND U2337 ( .A(n2112), .B(n2111), .Z(n2162) );
  XOR U2338 ( .A(n2163), .B(n2164), .Z(n2188) );
  NANDN U2339 ( .A(n2114), .B(n2113), .Z(n2118) );
  OR U2340 ( .A(n2116), .B(n2115), .Z(n2117) );
  NAND U2341 ( .A(n2118), .B(n2117), .Z(n2189) );
  XNOR U2342 ( .A(n2188), .B(n2189), .Z(n2190) );
  XOR U2343 ( .A(n2191), .B(n2190), .Z(n2137) );
  XNOR U2344 ( .A(n2136), .B(n2137), .Z(n2138) );
  XNOR U2345 ( .A(n2139), .B(n2138), .Z(n2197) );
  XOR U2346 ( .A(n2196), .B(n2197), .Z(n2130) );
  NANDN U2347 ( .A(n2120), .B(n2119), .Z(n2124) );
  NANDN U2348 ( .A(n2122), .B(n2121), .Z(n2123) );
  NAND U2349 ( .A(n2124), .B(n2123), .Z(n2131) );
  XNOR U2350 ( .A(n2130), .B(n2131), .Z(n2132) );
  XNOR U2351 ( .A(n2133), .B(n2132), .Z(n2200) );
  XNOR U2352 ( .A(n2200), .B(sreg[81]), .Z(n2202) );
  NAND U2353 ( .A(n2125), .B(sreg[80]), .Z(n2129) );
  OR U2354 ( .A(n2127), .B(n2126), .Z(n2128) );
  AND U2355 ( .A(n2129), .B(n2128), .Z(n2201) );
  XOR U2356 ( .A(n2202), .B(n2201), .Z(c[81]) );
  NANDN U2357 ( .A(n2131), .B(n2130), .Z(n2135) );
  NAND U2358 ( .A(n2133), .B(n2132), .Z(n2134) );
  NAND U2359 ( .A(n2135), .B(n2134), .Z(n2208) );
  NANDN U2360 ( .A(n2137), .B(n2136), .Z(n2141) );
  NAND U2361 ( .A(n2139), .B(n2138), .Z(n2140) );
  NAND U2362 ( .A(n2141), .B(n2140), .Z(n2269) );
  NANDN U2363 ( .A(n2143), .B(n2142), .Z(n2147) );
  NANDN U2364 ( .A(n2145), .B(n2144), .Z(n2146) );
  NAND U2365 ( .A(n2147), .B(n2146), .Z(n2270) );
  XNOR U2366 ( .A(n2269), .B(n2270), .Z(n2271) );
  XOR U2367 ( .A(n4859), .B(a[26]), .Z(n2223) );
  OR U2368 ( .A(n2223), .B(n4860), .Z(n2150) );
  NANDN U2369 ( .A(n2148), .B(n4915), .Z(n2149) );
  NAND U2370 ( .A(n2150), .B(n2149), .Z(n2235) );
  NANDN U2371 ( .A(n2151), .B(n4987), .Z(n2153) );
  XNOR U2372 ( .A(n4909), .B(n2453), .Z(n2226) );
  OR U2373 ( .A(n2226), .B(n4986), .Z(n2152) );
  NAND U2374 ( .A(n2153), .B(n2152), .Z(n2232) );
  XOR U2375 ( .A(n210), .B(a[20]), .Z(n2229) );
  OR U2376 ( .A(n2229), .B(n5095), .Z(n2156) );
  NANDN U2377 ( .A(n2154), .B(n5092), .Z(n2155) );
  AND U2378 ( .A(n2156), .B(n2155), .Z(n2233) );
  XOR U2379 ( .A(n2232), .B(n2233), .Z(n2234) );
  XOR U2380 ( .A(n2235), .B(n2234), .Z(n2217) );
  XNOR U2381 ( .A(n2217), .B(n2218), .Z(n2219) );
  NANDN U2382 ( .A(n2162), .B(n2161), .Z(n2166) );
  NANDN U2383 ( .A(n2164), .B(n2163), .Z(n2165) );
  NAND U2384 ( .A(n2166), .B(n2165), .Z(n2220) );
  XOR U2385 ( .A(n2219), .B(n2220), .Z(n2214) );
  NANDN U2386 ( .A(n2168), .B(n2167), .Z(n2172) );
  OR U2387 ( .A(n2170), .B(n2169), .Z(n2171) );
  NAND U2388 ( .A(n2172), .B(n2171), .Z(n2245) );
  XOR U2389 ( .A(n5129), .B(a[22]), .Z(n2251) );
  OR U2390 ( .A(n2251), .B(n5041), .Z(n2175) );
  NANDN U2391 ( .A(n2173), .B(n5052), .Z(n2174) );
  AND U2392 ( .A(n2175), .B(n2174), .Z(n2264) );
  NAND U2393 ( .A(b[0]), .B(a[34]), .Z(n2176) );
  XNOR U2394 ( .A(b[1]), .B(n2176), .Z(n2178) );
  NAND U2395 ( .A(a[33]), .B(n206), .Z(n2177) );
  AND U2396 ( .A(n2178), .B(n2177), .Z(n2263) );
  XOR U2397 ( .A(n2264), .B(n2263), .Z(n2266) );
  NAND U2398 ( .A(a[18]), .B(b[15]), .Z(n2265) );
  XOR U2399 ( .A(n2266), .B(n2265), .Z(n2242) );
  NAND U2400 ( .A(n4521), .B(n2179), .Z(n2181) );
  IV U2401 ( .A(a[32]), .Z(n3035) );
  XNOR U2402 ( .A(b[3]), .B(n3035), .Z(n2254) );
  NANDN U2403 ( .A(n4488), .B(n2254), .Z(n2180) );
  NAND U2404 ( .A(n2181), .B(n2180), .Z(n2238) );
  XOR U2405 ( .A(n209), .B(a[30]), .Z(n2257) );
  OR U2406 ( .A(n2257), .B(n4612), .Z(n2184) );
  NANDN U2407 ( .A(n2182), .B(n4669), .Z(n2183) );
  NAND U2408 ( .A(n2184), .B(n2183), .Z(n2236) );
  XNOR U2409 ( .A(n4744), .B(n2738), .Z(n2260) );
  NANDN U2410 ( .A(n2260), .B(n4745), .Z(n2187) );
  NANDN U2411 ( .A(n2185), .B(n4746), .Z(n2186) );
  AND U2412 ( .A(n2187), .B(n2186), .Z(n2237) );
  XOR U2413 ( .A(n2238), .B(n2239), .Z(n2243) );
  XNOR U2414 ( .A(n2242), .B(n2243), .Z(n2244) );
  XNOR U2415 ( .A(n2245), .B(n2244), .Z(n2212) );
  NANDN U2416 ( .A(n2189), .B(n2188), .Z(n2193) );
  NAND U2417 ( .A(n2191), .B(n2190), .Z(n2192) );
  AND U2418 ( .A(n2193), .B(n2192), .Z(n2211) );
  XNOR U2419 ( .A(n2212), .B(n2211), .Z(n2213) );
  XNOR U2420 ( .A(n2214), .B(n2213), .Z(n2272) );
  XOR U2421 ( .A(n2271), .B(n2272), .Z(n2205) );
  NANDN U2422 ( .A(n2195), .B(n2194), .Z(n2199) );
  NANDN U2423 ( .A(n2197), .B(n2196), .Z(n2198) );
  NAND U2424 ( .A(n2199), .B(n2198), .Z(n2206) );
  XNOR U2425 ( .A(n2205), .B(n2206), .Z(n2207) );
  XNOR U2426 ( .A(n2208), .B(n2207), .Z(n2275) );
  XNOR U2427 ( .A(n2275), .B(sreg[82]), .Z(n2277) );
  NAND U2428 ( .A(n2200), .B(sreg[81]), .Z(n2204) );
  OR U2429 ( .A(n2202), .B(n2201), .Z(n2203) );
  AND U2430 ( .A(n2204), .B(n2203), .Z(n2276) );
  XOR U2431 ( .A(n2277), .B(n2276), .Z(c[82]) );
  NANDN U2432 ( .A(n2206), .B(n2205), .Z(n2210) );
  NAND U2433 ( .A(n2208), .B(n2207), .Z(n2209) );
  NAND U2434 ( .A(n2210), .B(n2209), .Z(n2283) );
  NANDN U2435 ( .A(n2212), .B(n2211), .Z(n2216) );
  NAND U2436 ( .A(n2214), .B(n2213), .Z(n2215) );
  NAND U2437 ( .A(n2216), .B(n2215), .Z(n2344) );
  NANDN U2438 ( .A(n2218), .B(n2217), .Z(n2222) );
  NANDN U2439 ( .A(n2220), .B(n2219), .Z(n2221) );
  NAND U2440 ( .A(n2222), .B(n2221), .Z(n2345) );
  XNOR U2441 ( .A(n2344), .B(n2345), .Z(n2346) );
  XNOR U2442 ( .A(n4859), .B(n2664), .Z(n2298) );
  OR U2443 ( .A(n2298), .B(n4860), .Z(n2225) );
  NANDN U2444 ( .A(n2223), .B(n4915), .Z(n2224) );
  NAND U2445 ( .A(n2225), .B(n2224), .Z(n2310) );
  NANDN U2446 ( .A(n2226), .B(n4987), .Z(n2228) );
  XNOR U2447 ( .A(n4909), .B(n2527), .Z(n2301) );
  OR U2448 ( .A(n2301), .B(n4986), .Z(n2227) );
  NAND U2449 ( .A(n2228), .B(n2227), .Z(n2307) );
  XOR U2450 ( .A(n210), .B(a[21]), .Z(n2304) );
  OR U2451 ( .A(n2304), .B(n5095), .Z(n2231) );
  NANDN U2452 ( .A(n2229), .B(n5092), .Z(n2230) );
  AND U2453 ( .A(n2231), .B(n2230), .Z(n2308) );
  XOR U2454 ( .A(n2307), .B(n2308), .Z(n2309) );
  XOR U2455 ( .A(n2310), .B(n2309), .Z(n2292) );
  XNOR U2456 ( .A(n2292), .B(n2293), .Z(n2294) );
  NANDN U2457 ( .A(n2237), .B(n2236), .Z(n2241) );
  NANDN U2458 ( .A(n2239), .B(n2238), .Z(n2240) );
  NAND U2459 ( .A(n2241), .B(n2240), .Z(n2295) );
  XOR U2460 ( .A(n2294), .B(n2295), .Z(n2289) );
  NANDN U2461 ( .A(n2243), .B(n2242), .Z(n2247) );
  NAND U2462 ( .A(n2245), .B(n2244), .Z(n2246) );
  NAND U2463 ( .A(n2247), .B(n2246), .Z(n2286) );
  NAND U2464 ( .A(b[0]), .B(a[35]), .Z(n2248) );
  XNOR U2465 ( .A(b[1]), .B(n2248), .Z(n2250) );
  NAND U2466 ( .A(a[34]), .B(n206), .Z(n2249) );
  AND U2467 ( .A(n2250), .B(n2249), .Z(n2332) );
  XNOR U2468 ( .A(n5129), .B(n2379), .Z(n2320) );
  OR U2469 ( .A(n2320), .B(n5041), .Z(n2253) );
  NANDN U2470 ( .A(n2251), .B(n5052), .Z(n2252) );
  AND U2471 ( .A(n2253), .B(n2252), .Z(n2333) );
  XOR U2472 ( .A(n2332), .B(n2333), .Z(n2335) );
  NAND U2473 ( .A(b[15]), .B(a[19]), .Z(n2334) );
  XNOR U2474 ( .A(n2335), .B(n2334), .Z(n2341) );
  NAND U2475 ( .A(n4521), .B(n2254), .Z(n2256) );
  IV U2476 ( .A(a[33]), .Z(n3121) );
  XNOR U2477 ( .A(b[3]), .B(n3121), .Z(n2323) );
  NANDN U2478 ( .A(n4488), .B(n2323), .Z(n2255) );
  NAND U2479 ( .A(n2256), .B(n2255), .Z(n2313) );
  XNOR U2480 ( .A(n209), .B(n2971), .Z(n2326) );
  OR U2481 ( .A(n2326), .B(n4612), .Z(n2259) );
  NANDN U2482 ( .A(n2257), .B(n4669), .Z(n2258) );
  NAND U2483 ( .A(n2259), .B(n2258), .Z(n2311) );
  XNOR U2484 ( .A(n4744), .B(n2822), .Z(n2329) );
  NANDN U2485 ( .A(n2329), .B(n4745), .Z(n2262) );
  NANDN U2486 ( .A(n2260), .B(n4746), .Z(n2261) );
  AND U2487 ( .A(n2262), .B(n2261), .Z(n2312) );
  XOR U2488 ( .A(n2313), .B(n2314), .Z(n2338) );
  NANDN U2489 ( .A(n2264), .B(n2263), .Z(n2268) );
  OR U2490 ( .A(n2266), .B(n2265), .Z(n2267) );
  NAND U2491 ( .A(n2268), .B(n2267), .Z(n2339) );
  XNOR U2492 ( .A(n2338), .B(n2339), .Z(n2340) );
  XOR U2493 ( .A(n2341), .B(n2340), .Z(n2287) );
  XNOR U2494 ( .A(n2286), .B(n2287), .Z(n2288) );
  XNOR U2495 ( .A(n2289), .B(n2288), .Z(n2347) );
  XOR U2496 ( .A(n2346), .B(n2347), .Z(n2280) );
  NANDN U2497 ( .A(n2270), .B(n2269), .Z(n2274) );
  NANDN U2498 ( .A(n2272), .B(n2271), .Z(n2273) );
  NAND U2499 ( .A(n2274), .B(n2273), .Z(n2281) );
  XNOR U2500 ( .A(n2280), .B(n2281), .Z(n2282) );
  XNOR U2501 ( .A(n2283), .B(n2282), .Z(n2350) );
  XNOR U2502 ( .A(n2350), .B(sreg[83]), .Z(n2352) );
  NAND U2503 ( .A(n2275), .B(sreg[82]), .Z(n2279) );
  OR U2504 ( .A(n2277), .B(n2276), .Z(n2278) );
  AND U2505 ( .A(n2279), .B(n2278), .Z(n2351) );
  XOR U2506 ( .A(n2352), .B(n2351), .Z(c[83]) );
  NANDN U2507 ( .A(n2281), .B(n2280), .Z(n2285) );
  NAND U2508 ( .A(n2283), .B(n2282), .Z(n2284) );
  NAND U2509 ( .A(n2285), .B(n2284), .Z(n2358) );
  NANDN U2510 ( .A(n2287), .B(n2286), .Z(n2291) );
  NAND U2511 ( .A(n2289), .B(n2288), .Z(n2290) );
  NAND U2512 ( .A(n2291), .B(n2290), .Z(n2418) );
  NANDN U2513 ( .A(n2293), .B(n2292), .Z(n2297) );
  NANDN U2514 ( .A(n2295), .B(n2294), .Z(n2296) );
  NAND U2515 ( .A(n2297), .B(n2296), .Z(n2419) );
  XNOR U2516 ( .A(n2418), .B(n2419), .Z(n2420) );
  XNOR U2517 ( .A(n4859), .B(n2738), .Z(n2373) );
  OR U2518 ( .A(n2373), .B(n4860), .Z(n2300) );
  NANDN U2519 ( .A(n2298), .B(n4915), .Z(n2299) );
  NAND U2520 ( .A(n2300), .B(n2299), .Z(n2386) );
  NANDN U2521 ( .A(n2301), .B(n4987), .Z(n2303) );
  XOR U2522 ( .A(n4909), .B(a[26]), .Z(n2376) );
  OR U2523 ( .A(n2376), .B(n4986), .Z(n2302) );
  NAND U2524 ( .A(n2303), .B(n2302), .Z(n2383) );
  XOR U2525 ( .A(n210), .B(a[22]), .Z(n2380) );
  OR U2526 ( .A(n2380), .B(n5095), .Z(n2306) );
  NANDN U2527 ( .A(n2304), .B(n5092), .Z(n2305) );
  AND U2528 ( .A(n2306), .B(n2305), .Z(n2384) );
  XOR U2529 ( .A(n2383), .B(n2384), .Z(n2385) );
  XOR U2530 ( .A(n2386), .B(n2385), .Z(n2367) );
  XNOR U2531 ( .A(n2367), .B(n2368), .Z(n2369) );
  NANDN U2532 ( .A(n2312), .B(n2311), .Z(n2316) );
  NANDN U2533 ( .A(n2314), .B(n2313), .Z(n2315) );
  NAND U2534 ( .A(n2316), .B(n2315), .Z(n2370) );
  XOR U2535 ( .A(n2369), .B(n2370), .Z(n2364) );
  NAND U2536 ( .A(b[0]), .B(a[36]), .Z(n2317) );
  XNOR U2537 ( .A(b[1]), .B(n2317), .Z(n2319) );
  NAND U2538 ( .A(a[35]), .B(n206), .Z(n2318) );
  AND U2539 ( .A(n2319), .B(n2318), .Z(n2408) );
  XNOR U2540 ( .A(n5129), .B(n2453), .Z(n2393) );
  OR U2541 ( .A(n2393), .B(n5041), .Z(n2322) );
  NANDN U2542 ( .A(n2320), .B(n5052), .Z(n2321) );
  AND U2543 ( .A(n2322), .B(n2321), .Z(n2409) );
  XOR U2544 ( .A(n2408), .B(n2409), .Z(n2411) );
  NAND U2545 ( .A(b[15]), .B(a[20]), .Z(n2410) );
  XNOR U2546 ( .A(n2411), .B(n2410), .Z(n2417) );
  NAND U2547 ( .A(n4521), .B(n2323), .Z(n2325) );
  IV U2548 ( .A(a[34]), .Z(n3197) );
  XNOR U2549 ( .A(b[3]), .B(n3197), .Z(n2399) );
  NANDN U2550 ( .A(n4488), .B(n2399), .Z(n2324) );
  NAND U2551 ( .A(n2325), .B(n2324), .Z(n2389) );
  XNOR U2552 ( .A(n209), .B(n3035), .Z(n2402) );
  OR U2553 ( .A(n2402), .B(n4612), .Z(n2328) );
  NANDN U2554 ( .A(n2326), .B(n4669), .Z(n2327) );
  NAND U2555 ( .A(n2328), .B(n2327), .Z(n2387) );
  XOR U2556 ( .A(n4744), .B(a[30]), .Z(n2405) );
  NANDN U2557 ( .A(n2405), .B(n4745), .Z(n2331) );
  NANDN U2558 ( .A(n2329), .B(n4746), .Z(n2330) );
  AND U2559 ( .A(n2331), .B(n2330), .Z(n2388) );
  XOR U2560 ( .A(n2389), .B(n2390), .Z(n2414) );
  NANDN U2561 ( .A(n2333), .B(n2332), .Z(n2337) );
  OR U2562 ( .A(n2335), .B(n2334), .Z(n2336) );
  NAND U2563 ( .A(n2337), .B(n2336), .Z(n2415) );
  XOR U2564 ( .A(n2414), .B(n2415), .Z(n2416) );
  XOR U2565 ( .A(n2417), .B(n2416), .Z(n2361) );
  NANDN U2566 ( .A(n2339), .B(n2338), .Z(n2343) );
  NAND U2567 ( .A(n2341), .B(n2340), .Z(n2342) );
  NAND U2568 ( .A(n2343), .B(n2342), .Z(n2362) );
  XNOR U2569 ( .A(n2361), .B(n2362), .Z(n2363) );
  XNOR U2570 ( .A(n2364), .B(n2363), .Z(n2421) );
  XOR U2571 ( .A(n2420), .B(n2421), .Z(n2355) );
  NANDN U2572 ( .A(n2345), .B(n2344), .Z(n2349) );
  NANDN U2573 ( .A(n2347), .B(n2346), .Z(n2348) );
  NAND U2574 ( .A(n2349), .B(n2348), .Z(n2356) );
  XNOR U2575 ( .A(n2355), .B(n2356), .Z(n2357) );
  XNOR U2576 ( .A(n2358), .B(n2357), .Z(n2424) );
  XNOR U2577 ( .A(n2424), .B(sreg[84]), .Z(n2426) );
  NAND U2578 ( .A(n2350), .B(sreg[83]), .Z(n2354) );
  OR U2579 ( .A(n2352), .B(n2351), .Z(n2353) );
  AND U2580 ( .A(n2354), .B(n2353), .Z(n2425) );
  XOR U2581 ( .A(n2426), .B(n2425), .Z(c[84]) );
  NANDN U2582 ( .A(n2356), .B(n2355), .Z(n2360) );
  NAND U2583 ( .A(n2358), .B(n2357), .Z(n2359) );
  NAND U2584 ( .A(n2360), .B(n2359), .Z(n2432) );
  NANDN U2585 ( .A(n2362), .B(n2361), .Z(n2366) );
  NAND U2586 ( .A(n2364), .B(n2363), .Z(n2365) );
  NAND U2587 ( .A(n2366), .B(n2365), .Z(n2492) );
  NANDN U2588 ( .A(n2368), .B(n2367), .Z(n2372) );
  NANDN U2589 ( .A(n2370), .B(n2369), .Z(n2371) );
  NAND U2590 ( .A(n2372), .B(n2371), .Z(n2493) );
  XNOR U2591 ( .A(n2492), .B(n2493), .Z(n2494) );
  XNOR U2592 ( .A(n4859), .B(n2822), .Z(n2447) );
  OR U2593 ( .A(n2447), .B(n4860), .Z(n2375) );
  NANDN U2594 ( .A(n2373), .B(n4915), .Z(n2374) );
  NAND U2595 ( .A(n2375), .B(n2374), .Z(n2460) );
  NANDN U2596 ( .A(n2376), .B(n4987), .Z(n2378) );
  XNOR U2597 ( .A(n4909), .B(n2664), .Z(n2450) );
  OR U2598 ( .A(n2450), .B(n4986), .Z(n2377) );
  NAND U2599 ( .A(n2378), .B(n2377), .Z(n2457) );
  XNOR U2600 ( .A(n210), .B(n2379), .Z(n2454) );
  OR U2601 ( .A(n2454), .B(n5095), .Z(n2382) );
  NANDN U2602 ( .A(n2380), .B(n5092), .Z(n2381) );
  AND U2603 ( .A(n2382), .B(n2381), .Z(n2458) );
  XOR U2604 ( .A(n2457), .B(n2458), .Z(n2459) );
  XOR U2605 ( .A(n2460), .B(n2459), .Z(n2441) );
  XNOR U2606 ( .A(n2441), .B(n2442), .Z(n2443) );
  NANDN U2607 ( .A(n2388), .B(n2387), .Z(n2392) );
  NANDN U2608 ( .A(n2390), .B(n2389), .Z(n2391) );
  NAND U2609 ( .A(n2392), .B(n2391), .Z(n2444) );
  XOR U2610 ( .A(n2443), .B(n2444), .Z(n2438) );
  XNOR U2611 ( .A(n5129), .B(n2527), .Z(n2467) );
  OR U2612 ( .A(n2467), .B(n5041), .Z(n2395) );
  NANDN U2613 ( .A(n2393), .B(n5052), .Z(n2394) );
  AND U2614 ( .A(n2395), .B(n2394), .Z(n2483) );
  NAND U2615 ( .A(b[0]), .B(a[37]), .Z(n2396) );
  XNOR U2616 ( .A(b[1]), .B(n2396), .Z(n2398) );
  NAND U2617 ( .A(a[36]), .B(n206), .Z(n2397) );
  AND U2618 ( .A(n2398), .B(n2397), .Z(n2482) );
  XOR U2619 ( .A(n2483), .B(n2482), .Z(n2485) );
  NAND U2620 ( .A(b[15]), .B(a[21]), .Z(n2484) );
  XNOR U2621 ( .A(n2485), .B(n2484), .Z(n2491) );
  NAND U2622 ( .A(n4521), .B(n2399), .Z(n2401) );
  IV U2623 ( .A(a[35]), .Z(n3273) );
  XNOR U2624 ( .A(b[3]), .B(n3273), .Z(n2473) );
  NANDN U2625 ( .A(n4488), .B(n2473), .Z(n2400) );
  NAND U2626 ( .A(n2401), .B(n2400), .Z(n2463) );
  XNOR U2627 ( .A(n209), .B(n3121), .Z(n2476) );
  OR U2628 ( .A(n2476), .B(n4612), .Z(n2404) );
  NANDN U2629 ( .A(n2402), .B(n4669), .Z(n2403) );
  NAND U2630 ( .A(n2404), .B(n2403), .Z(n2461) );
  XNOR U2631 ( .A(n4744), .B(n2971), .Z(n2479) );
  NANDN U2632 ( .A(n2479), .B(n4745), .Z(n2407) );
  NANDN U2633 ( .A(n2405), .B(n4746), .Z(n2406) );
  AND U2634 ( .A(n2407), .B(n2406), .Z(n2462) );
  XOR U2635 ( .A(n2463), .B(n2464), .Z(n2488) );
  NANDN U2636 ( .A(n2409), .B(n2408), .Z(n2413) );
  OR U2637 ( .A(n2411), .B(n2410), .Z(n2412) );
  NAND U2638 ( .A(n2413), .B(n2412), .Z(n2489) );
  XOR U2639 ( .A(n2488), .B(n2489), .Z(n2490) );
  XOR U2640 ( .A(n2491), .B(n2490), .Z(n2435) );
  XNOR U2641 ( .A(n2435), .B(n2436), .Z(n2437) );
  XNOR U2642 ( .A(n2438), .B(n2437), .Z(n2495) );
  XOR U2643 ( .A(n2494), .B(n2495), .Z(n2429) );
  NANDN U2644 ( .A(n2419), .B(n2418), .Z(n2423) );
  NANDN U2645 ( .A(n2421), .B(n2420), .Z(n2422) );
  NAND U2646 ( .A(n2423), .B(n2422), .Z(n2430) );
  XNOR U2647 ( .A(n2429), .B(n2430), .Z(n2431) );
  XNOR U2648 ( .A(n2432), .B(n2431), .Z(n2498) );
  XNOR U2649 ( .A(n2498), .B(sreg[85]), .Z(n2500) );
  NAND U2650 ( .A(n2424), .B(sreg[84]), .Z(n2428) );
  OR U2651 ( .A(n2426), .B(n2425), .Z(n2427) );
  AND U2652 ( .A(n2428), .B(n2427), .Z(n2499) );
  XOR U2653 ( .A(n2500), .B(n2499), .Z(c[85]) );
  NANDN U2654 ( .A(n2430), .B(n2429), .Z(n2434) );
  NAND U2655 ( .A(n2432), .B(n2431), .Z(n2433) );
  NAND U2656 ( .A(n2434), .B(n2433), .Z(n2506) );
  NANDN U2657 ( .A(n2436), .B(n2435), .Z(n2440) );
  NAND U2658 ( .A(n2438), .B(n2437), .Z(n2439) );
  NAND U2659 ( .A(n2440), .B(n2439), .Z(n2566) );
  NANDN U2660 ( .A(n2442), .B(n2441), .Z(n2446) );
  NANDN U2661 ( .A(n2444), .B(n2443), .Z(n2445) );
  NAND U2662 ( .A(n2446), .B(n2445), .Z(n2567) );
  XNOR U2663 ( .A(n2566), .B(n2567), .Z(n2568) );
  XOR U2664 ( .A(n4859), .B(a[30]), .Z(n2521) );
  OR U2665 ( .A(n2521), .B(n4860), .Z(n2449) );
  NANDN U2666 ( .A(n2447), .B(n4915), .Z(n2448) );
  NAND U2667 ( .A(n2449), .B(n2448), .Z(n2534) );
  NANDN U2668 ( .A(n2450), .B(n4987), .Z(n2452) );
  XNOR U2669 ( .A(n4909), .B(n2738), .Z(n2524) );
  OR U2670 ( .A(n2524), .B(n4986), .Z(n2451) );
  NAND U2671 ( .A(n2452), .B(n2451), .Z(n2531) );
  XNOR U2672 ( .A(n210), .B(n2453), .Z(n2528) );
  OR U2673 ( .A(n2528), .B(n5095), .Z(n2456) );
  NANDN U2674 ( .A(n2454), .B(n5092), .Z(n2455) );
  AND U2675 ( .A(n2456), .B(n2455), .Z(n2532) );
  XOR U2676 ( .A(n2531), .B(n2532), .Z(n2533) );
  XOR U2677 ( .A(n2534), .B(n2533), .Z(n2515) );
  XNOR U2678 ( .A(n2515), .B(n2516), .Z(n2517) );
  NANDN U2679 ( .A(n2462), .B(n2461), .Z(n2466) );
  NANDN U2680 ( .A(n2464), .B(n2463), .Z(n2465) );
  NAND U2681 ( .A(n2466), .B(n2465), .Z(n2518) );
  XOR U2682 ( .A(n2517), .B(n2518), .Z(n2512) );
  XOR U2683 ( .A(n5129), .B(a[26]), .Z(n2550) );
  OR U2684 ( .A(n2550), .B(n5041), .Z(n2469) );
  NANDN U2685 ( .A(n2467), .B(n5052), .Z(n2468) );
  AND U2686 ( .A(n2469), .B(n2468), .Z(n2542) );
  NAND U2687 ( .A(b[0]), .B(a[38]), .Z(n2470) );
  XNOR U2688 ( .A(b[1]), .B(n2470), .Z(n2472) );
  NAND U2689 ( .A(n206), .B(a[37]), .Z(n2471) );
  AND U2690 ( .A(n2472), .B(n2471), .Z(n2541) );
  XOR U2691 ( .A(n2542), .B(n2541), .Z(n2544) );
  NAND U2692 ( .A(b[15]), .B(a[22]), .Z(n2543) );
  XNOR U2693 ( .A(n2544), .B(n2543), .Z(n2565) );
  NAND U2694 ( .A(n4521), .B(n2473), .Z(n2475) );
  IV U2695 ( .A(a[36]), .Z(n3347) );
  XNOR U2696 ( .A(b[3]), .B(n3347), .Z(n2553) );
  NANDN U2697 ( .A(n4488), .B(n2553), .Z(n2474) );
  NAND U2698 ( .A(n2475), .B(n2474), .Z(n2537) );
  XNOR U2699 ( .A(n209), .B(n3197), .Z(n2556) );
  OR U2700 ( .A(n2556), .B(n4612), .Z(n2478) );
  NANDN U2701 ( .A(n2476), .B(n4669), .Z(n2477) );
  NAND U2702 ( .A(n2478), .B(n2477), .Z(n2535) );
  XNOR U2703 ( .A(n4744), .B(n3035), .Z(n2559) );
  NANDN U2704 ( .A(n2559), .B(n4745), .Z(n2481) );
  NANDN U2705 ( .A(n2479), .B(n4746), .Z(n2480) );
  AND U2706 ( .A(n2481), .B(n2480), .Z(n2536) );
  XOR U2707 ( .A(n2537), .B(n2538), .Z(n2562) );
  NANDN U2708 ( .A(n2483), .B(n2482), .Z(n2487) );
  OR U2709 ( .A(n2485), .B(n2484), .Z(n2486) );
  NAND U2710 ( .A(n2487), .B(n2486), .Z(n2563) );
  XOR U2711 ( .A(n2562), .B(n2563), .Z(n2564) );
  XOR U2712 ( .A(n2565), .B(n2564), .Z(n2509) );
  XNOR U2713 ( .A(n2509), .B(n2510), .Z(n2511) );
  XNOR U2714 ( .A(n2512), .B(n2511), .Z(n2569) );
  XOR U2715 ( .A(n2568), .B(n2569), .Z(n2503) );
  NANDN U2716 ( .A(n2493), .B(n2492), .Z(n2497) );
  NANDN U2717 ( .A(n2495), .B(n2494), .Z(n2496) );
  NAND U2718 ( .A(n2497), .B(n2496), .Z(n2504) );
  XNOR U2719 ( .A(n2503), .B(n2504), .Z(n2505) );
  XNOR U2720 ( .A(n2506), .B(n2505), .Z(n2572) );
  XNOR U2721 ( .A(n2572), .B(sreg[86]), .Z(n2574) );
  NAND U2722 ( .A(n2498), .B(sreg[85]), .Z(n2502) );
  OR U2723 ( .A(n2500), .B(n2499), .Z(n2501) );
  AND U2724 ( .A(n2502), .B(n2501), .Z(n2573) );
  XOR U2725 ( .A(n2574), .B(n2573), .Z(c[86]) );
  NANDN U2726 ( .A(n2504), .B(n2503), .Z(n2508) );
  NAND U2727 ( .A(n2506), .B(n2505), .Z(n2507) );
  NAND U2728 ( .A(n2508), .B(n2507), .Z(n2580) );
  NANDN U2729 ( .A(n2510), .B(n2509), .Z(n2514) );
  NAND U2730 ( .A(n2512), .B(n2511), .Z(n2513) );
  NAND U2731 ( .A(n2514), .B(n2513), .Z(n2641) );
  NANDN U2732 ( .A(n2516), .B(n2515), .Z(n2520) );
  NANDN U2733 ( .A(n2518), .B(n2517), .Z(n2519) );
  NAND U2734 ( .A(n2520), .B(n2519), .Z(n2642) );
  XNOR U2735 ( .A(n2641), .B(n2642), .Z(n2643) );
  XNOR U2736 ( .A(n4859), .B(n2971), .Z(n2595) );
  OR U2737 ( .A(n2595), .B(n4860), .Z(n2523) );
  NANDN U2738 ( .A(n2521), .B(n4915), .Z(n2522) );
  NAND U2739 ( .A(n2523), .B(n2522), .Z(n2607) );
  NANDN U2740 ( .A(n2524), .B(n4987), .Z(n2526) );
  XNOR U2741 ( .A(n4909), .B(n2822), .Z(n2598) );
  OR U2742 ( .A(n2598), .B(n4986), .Z(n2525) );
  NAND U2743 ( .A(n2526), .B(n2525), .Z(n2604) );
  XNOR U2744 ( .A(n210), .B(n2527), .Z(n2601) );
  OR U2745 ( .A(n2601), .B(n5095), .Z(n2530) );
  NANDN U2746 ( .A(n2528), .B(n5092), .Z(n2529) );
  AND U2747 ( .A(n2530), .B(n2529), .Z(n2605) );
  XOR U2748 ( .A(n2604), .B(n2605), .Z(n2606) );
  XOR U2749 ( .A(n2607), .B(n2606), .Z(n2589) );
  XNOR U2750 ( .A(n2589), .B(n2590), .Z(n2591) );
  NANDN U2751 ( .A(n2536), .B(n2535), .Z(n2540) );
  NANDN U2752 ( .A(n2538), .B(n2537), .Z(n2539) );
  NAND U2753 ( .A(n2540), .B(n2539), .Z(n2592) );
  XOR U2754 ( .A(n2591), .B(n2592), .Z(n2586) );
  NANDN U2755 ( .A(n2542), .B(n2541), .Z(n2546) );
  OR U2756 ( .A(n2544), .B(n2543), .Z(n2545) );
  NAND U2757 ( .A(n2546), .B(n2545), .Z(n2617) );
  NAND U2758 ( .A(b[0]), .B(a[39]), .Z(n2547) );
  XNOR U2759 ( .A(b[1]), .B(n2547), .Z(n2549) );
  NAND U2760 ( .A(a[38]), .B(n206), .Z(n2548) );
  AND U2761 ( .A(n2549), .B(n2548), .Z(n2620) );
  XNOR U2762 ( .A(n5129), .B(n2664), .Z(n2629) );
  OR U2763 ( .A(n2629), .B(n5041), .Z(n2552) );
  NANDN U2764 ( .A(n2550), .B(n5052), .Z(n2551) );
  AND U2765 ( .A(n2552), .B(n2551), .Z(n2621) );
  XOR U2766 ( .A(n2620), .B(n2621), .Z(n2623) );
  NAND U2767 ( .A(a[23]), .B(b[15]), .Z(n2622) );
  XOR U2768 ( .A(n2623), .B(n2622), .Z(n2614) );
  NAND U2769 ( .A(n4521), .B(n2553), .Z(n2555) );
  XOR U2770 ( .A(b[3]), .B(a[37]), .Z(n2632) );
  NANDN U2771 ( .A(n4488), .B(n2632), .Z(n2554) );
  NAND U2772 ( .A(n2555), .B(n2554), .Z(n2610) );
  XNOR U2773 ( .A(n209), .B(n3273), .Z(n2635) );
  OR U2774 ( .A(n2635), .B(n4612), .Z(n2558) );
  NANDN U2775 ( .A(n2556), .B(n4669), .Z(n2557) );
  NAND U2776 ( .A(n2558), .B(n2557), .Z(n2608) );
  XNOR U2777 ( .A(n4744), .B(n3121), .Z(n2638) );
  NANDN U2778 ( .A(n2638), .B(n4745), .Z(n2561) );
  NANDN U2779 ( .A(n2559), .B(n4746), .Z(n2560) );
  AND U2780 ( .A(n2561), .B(n2560), .Z(n2609) );
  XOR U2781 ( .A(n2610), .B(n2611), .Z(n2615) );
  XNOR U2782 ( .A(n2614), .B(n2615), .Z(n2616) );
  XNOR U2783 ( .A(n2617), .B(n2616), .Z(n2584) );
  XNOR U2784 ( .A(n2584), .B(n2583), .Z(n2585) );
  XNOR U2785 ( .A(n2586), .B(n2585), .Z(n2644) );
  XOR U2786 ( .A(n2643), .B(n2644), .Z(n2577) );
  NANDN U2787 ( .A(n2567), .B(n2566), .Z(n2571) );
  NANDN U2788 ( .A(n2569), .B(n2568), .Z(n2570) );
  NAND U2789 ( .A(n2571), .B(n2570), .Z(n2578) );
  XNOR U2790 ( .A(n2577), .B(n2578), .Z(n2579) );
  XNOR U2791 ( .A(n2580), .B(n2579), .Z(n2647) );
  XNOR U2792 ( .A(n2647), .B(sreg[87]), .Z(n2649) );
  NAND U2793 ( .A(n2572), .B(sreg[86]), .Z(n2576) );
  OR U2794 ( .A(n2574), .B(n2573), .Z(n2575) );
  AND U2795 ( .A(n2576), .B(n2575), .Z(n2648) );
  XOR U2796 ( .A(n2649), .B(n2648), .Z(c[87]) );
  NANDN U2797 ( .A(n2578), .B(n2577), .Z(n2582) );
  NAND U2798 ( .A(n2580), .B(n2579), .Z(n2581) );
  NAND U2799 ( .A(n2582), .B(n2581), .Z(n2655) );
  NANDN U2800 ( .A(n2584), .B(n2583), .Z(n2588) );
  NAND U2801 ( .A(n2586), .B(n2585), .Z(n2587) );
  NAND U2802 ( .A(n2588), .B(n2587), .Z(n2717) );
  NANDN U2803 ( .A(n2590), .B(n2589), .Z(n2594) );
  NANDN U2804 ( .A(n2592), .B(n2591), .Z(n2593) );
  NAND U2805 ( .A(n2594), .B(n2593), .Z(n2718) );
  XNOR U2806 ( .A(n2717), .B(n2718), .Z(n2719) );
  XNOR U2807 ( .A(n4859), .B(n3035), .Z(n2658) );
  OR U2808 ( .A(n2658), .B(n4860), .Z(n2597) );
  NANDN U2809 ( .A(n2595), .B(n4915), .Z(n2596) );
  NAND U2810 ( .A(n2597), .B(n2596), .Z(n2671) );
  NANDN U2811 ( .A(n2598), .B(n4987), .Z(n2600) );
  XOR U2812 ( .A(n4909), .B(a[30]), .Z(n2661) );
  OR U2813 ( .A(n2661), .B(n4986), .Z(n2599) );
  NAND U2814 ( .A(n2600), .B(n2599), .Z(n2668) );
  XOR U2815 ( .A(n210), .B(a[26]), .Z(n2665) );
  OR U2816 ( .A(n2665), .B(n5095), .Z(n2603) );
  NANDN U2817 ( .A(n2601), .B(n5092), .Z(n2602) );
  AND U2818 ( .A(n2603), .B(n2602), .Z(n2669) );
  XOR U2819 ( .A(n2668), .B(n2669), .Z(n2670) );
  XOR U2820 ( .A(n2671), .B(n2670), .Z(n2711) );
  XNOR U2821 ( .A(n2711), .B(n2712), .Z(n2713) );
  NANDN U2822 ( .A(n2609), .B(n2608), .Z(n2613) );
  NANDN U2823 ( .A(n2611), .B(n2610), .Z(n2612) );
  NAND U2824 ( .A(n2613), .B(n2612), .Z(n2714) );
  XOR U2825 ( .A(n2713), .B(n2714), .Z(n2708) );
  NANDN U2826 ( .A(n2615), .B(n2614), .Z(n2619) );
  NAND U2827 ( .A(n2617), .B(n2616), .Z(n2618) );
  NAND U2828 ( .A(n2619), .B(n2618), .Z(n2705) );
  NANDN U2829 ( .A(n2621), .B(n2620), .Z(n2625) );
  OR U2830 ( .A(n2623), .B(n2622), .Z(n2624) );
  NAND U2831 ( .A(n2625), .B(n2624), .Z(n2702) );
  NAND U2832 ( .A(b[0]), .B(a[40]), .Z(n2626) );
  XNOR U2833 ( .A(b[1]), .B(n2626), .Z(n2628) );
  NAND U2834 ( .A(a[39]), .B(n206), .Z(n2627) );
  AND U2835 ( .A(n2628), .B(n2627), .Z(n2678) );
  XNOR U2836 ( .A(n5129), .B(n2738), .Z(n2684) );
  OR U2837 ( .A(n2684), .B(n5041), .Z(n2631) );
  NANDN U2838 ( .A(n2629), .B(n5052), .Z(n2630) );
  AND U2839 ( .A(n2631), .B(n2630), .Z(n2679) );
  XOR U2840 ( .A(n2678), .B(n2679), .Z(n2681) );
  NAND U2841 ( .A(a[24]), .B(b[15]), .Z(n2680) );
  XOR U2842 ( .A(n2681), .B(n2680), .Z(n2699) );
  NAND U2843 ( .A(n4521), .B(n2632), .Z(n2634) );
  IV U2844 ( .A(a[38]), .Z(n3496) );
  XNOR U2845 ( .A(b[3]), .B(n3496), .Z(n2690) );
  NANDN U2846 ( .A(n4488), .B(n2690), .Z(n2633) );
  NAND U2847 ( .A(n2634), .B(n2633), .Z(n2674) );
  XNOR U2848 ( .A(n209), .B(n3347), .Z(n2693) );
  OR U2849 ( .A(n2693), .B(n4612), .Z(n2637) );
  NANDN U2850 ( .A(n2635), .B(n4669), .Z(n2636) );
  NAND U2851 ( .A(n2637), .B(n2636), .Z(n2672) );
  XNOR U2852 ( .A(n4744), .B(n3197), .Z(n2696) );
  NANDN U2853 ( .A(n2696), .B(n4745), .Z(n2640) );
  NANDN U2854 ( .A(n2638), .B(n4746), .Z(n2639) );
  AND U2855 ( .A(n2640), .B(n2639), .Z(n2673) );
  XOR U2856 ( .A(n2674), .B(n2675), .Z(n2700) );
  XNOR U2857 ( .A(n2699), .B(n2700), .Z(n2701) );
  XNOR U2858 ( .A(n2702), .B(n2701), .Z(n2706) );
  XNOR U2859 ( .A(n2705), .B(n2706), .Z(n2707) );
  XNOR U2860 ( .A(n2708), .B(n2707), .Z(n2720) );
  XOR U2861 ( .A(n2719), .B(n2720), .Z(n2652) );
  NANDN U2862 ( .A(n2642), .B(n2641), .Z(n2646) );
  NANDN U2863 ( .A(n2644), .B(n2643), .Z(n2645) );
  NAND U2864 ( .A(n2646), .B(n2645), .Z(n2653) );
  XNOR U2865 ( .A(n2652), .B(n2653), .Z(n2654) );
  XNOR U2866 ( .A(n2655), .B(n2654), .Z(n2723) );
  XNOR U2867 ( .A(n2723), .B(sreg[88]), .Z(n2725) );
  NAND U2868 ( .A(n2647), .B(sreg[87]), .Z(n2651) );
  OR U2869 ( .A(n2649), .B(n2648), .Z(n2650) );
  AND U2870 ( .A(n2651), .B(n2650), .Z(n2724) );
  XOR U2871 ( .A(n2725), .B(n2724), .Z(c[88]) );
  NANDN U2872 ( .A(n2653), .B(n2652), .Z(n2657) );
  NAND U2873 ( .A(n2655), .B(n2654), .Z(n2656) );
  NAND U2874 ( .A(n2657), .B(n2656), .Z(n2731) );
  XNOR U2875 ( .A(n4859), .B(n3121), .Z(n2732) );
  OR U2876 ( .A(n2732), .B(n4860), .Z(n2660) );
  NANDN U2877 ( .A(n2658), .B(n4915), .Z(n2659) );
  NAND U2878 ( .A(n2660), .B(n2659), .Z(n2745) );
  NANDN U2879 ( .A(n2661), .B(n4987), .Z(n2663) );
  XNOR U2880 ( .A(n4909), .B(n2971), .Z(n2735) );
  OR U2881 ( .A(n2735), .B(n4986), .Z(n2662) );
  NAND U2882 ( .A(n2663), .B(n2662), .Z(n2742) );
  XNOR U2883 ( .A(n210), .B(n2664), .Z(n2739) );
  OR U2884 ( .A(n2739), .B(n5095), .Z(n2667) );
  NANDN U2885 ( .A(n2665), .B(n5092), .Z(n2666) );
  AND U2886 ( .A(n2667), .B(n2666), .Z(n2743) );
  XOR U2887 ( .A(n2742), .B(n2743), .Z(n2744) );
  XOR U2888 ( .A(n2745), .B(n2744), .Z(n2777) );
  XOR U2889 ( .A(n2777), .B(n2778), .Z(n2780) );
  NANDN U2890 ( .A(n2673), .B(n2672), .Z(n2677) );
  NANDN U2891 ( .A(n2675), .B(n2674), .Z(n2676) );
  AND U2892 ( .A(n2677), .B(n2676), .Z(n2779) );
  XOR U2893 ( .A(n2780), .B(n2779), .Z(n2785) );
  NANDN U2894 ( .A(n2679), .B(n2678), .Z(n2683) );
  OR U2895 ( .A(n2681), .B(n2680), .Z(n2682) );
  NAND U2896 ( .A(n2683), .B(n2682), .Z(n2776) );
  XNOR U2897 ( .A(n5129), .B(n2822), .Z(n2755) );
  OR U2898 ( .A(n2755), .B(n5041), .Z(n2686) );
  NANDN U2899 ( .A(n2684), .B(n5052), .Z(n2685) );
  NAND U2900 ( .A(n2686), .B(n2685), .Z(n2767) );
  AND U2901 ( .A(a[41]), .B(b[0]), .Z(n2687) );
  XOR U2902 ( .A(b[1]), .B(n2687), .Z(n2689) );
  NAND U2903 ( .A(n206), .B(a[40]), .Z(n2688) );
  NAND U2904 ( .A(n2689), .B(n2688), .Z(n2768) );
  XNOR U2905 ( .A(n2767), .B(n2768), .Z(n2769) );
  NAND U2906 ( .A(a[25]), .B(b[15]), .Z(n2770) );
  XOR U2907 ( .A(n2769), .B(n2770), .Z(n2773) );
  NAND U2908 ( .A(n4521), .B(n2690), .Z(n2692) );
  IV U2909 ( .A(a[39]), .Z(n3560) );
  XNOR U2910 ( .A(b[3]), .B(n3560), .Z(n2758) );
  NANDN U2911 ( .A(n4488), .B(n2758), .Z(n2691) );
  NAND U2912 ( .A(n2692), .B(n2691), .Z(n2748) );
  XOR U2913 ( .A(n209), .B(a[37]), .Z(n2761) );
  OR U2914 ( .A(n2761), .B(n4612), .Z(n2695) );
  NANDN U2915 ( .A(n2693), .B(n4669), .Z(n2694) );
  NAND U2916 ( .A(n2695), .B(n2694), .Z(n2746) );
  XNOR U2917 ( .A(n4744), .B(n3273), .Z(n2764) );
  NANDN U2918 ( .A(n2764), .B(n4745), .Z(n2698) );
  NANDN U2919 ( .A(n2696), .B(n4746), .Z(n2697) );
  AND U2920 ( .A(n2698), .B(n2697), .Z(n2747) );
  XOR U2921 ( .A(n2748), .B(n2749), .Z(n2774) );
  XOR U2922 ( .A(n2773), .B(n2774), .Z(n2775) );
  XNOR U2923 ( .A(n2776), .B(n2775), .Z(n2783) );
  NANDN U2924 ( .A(n2700), .B(n2699), .Z(n2704) );
  NAND U2925 ( .A(n2702), .B(n2701), .Z(n2703) );
  NAND U2926 ( .A(n2704), .B(n2703), .Z(n2784) );
  XOR U2927 ( .A(n2783), .B(n2784), .Z(n2786) );
  XNOR U2928 ( .A(n2785), .B(n2786), .Z(n2792) );
  NANDN U2929 ( .A(n2706), .B(n2705), .Z(n2710) );
  NAND U2930 ( .A(n2708), .B(n2707), .Z(n2709) );
  NAND U2931 ( .A(n2710), .B(n2709), .Z(n2789) );
  NANDN U2932 ( .A(n2712), .B(n2711), .Z(n2716) );
  NANDN U2933 ( .A(n2714), .B(n2713), .Z(n2715) );
  NAND U2934 ( .A(n2716), .B(n2715), .Z(n2790) );
  XNOR U2935 ( .A(n2789), .B(n2790), .Z(n2791) );
  XNOR U2936 ( .A(n2792), .B(n2791), .Z(n2728) );
  NANDN U2937 ( .A(n2718), .B(n2717), .Z(n2722) );
  NANDN U2938 ( .A(n2720), .B(n2719), .Z(n2721) );
  NAND U2939 ( .A(n2722), .B(n2721), .Z(n2729) );
  XOR U2940 ( .A(n2728), .B(n2729), .Z(n2730) );
  XOR U2941 ( .A(n2731), .B(n2730), .Z(n2795) );
  XNOR U2942 ( .A(n2795), .B(sreg[89]), .Z(n2797) );
  NAND U2943 ( .A(n2723), .B(sreg[88]), .Z(n2727) );
  OR U2944 ( .A(n2725), .B(n2724), .Z(n2726) );
  AND U2945 ( .A(n2727), .B(n2726), .Z(n2796) );
  XOR U2946 ( .A(n2797), .B(n2796), .Z(c[89]) );
  XNOR U2947 ( .A(n4859), .B(n3197), .Z(n2816) );
  OR U2948 ( .A(n2816), .B(n4860), .Z(n2734) );
  NANDN U2949 ( .A(n2732), .B(n4915), .Z(n2733) );
  NAND U2950 ( .A(n2734), .B(n2733), .Z(n2829) );
  NANDN U2951 ( .A(n2735), .B(n4987), .Z(n2737) );
  XNOR U2952 ( .A(n4909), .B(n3035), .Z(n2819) );
  OR U2953 ( .A(n2819), .B(n4986), .Z(n2736) );
  NAND U2954 ( .A(n2737), .B(n2736), .Z(n2826) );
  XNOR U2955 ( .A(n210), .B(n2738), .Z(n2823) );
  OR U2956 ( .A(n2823), .B(n5095), .Z(n2741) );
  NANDN U2957 ( .A(n2739), .B(n5092), .Z(n2740) );
  AND U2958 ( .A(n2741), .B(n2740), .Z(n2827) );
  XOR U2959 ( .A(n2826), .B(n2827), .Z(n2828) );
  XOR U2960 ( .A(n2829), .B(n2828), .Z(n2804) );
  XOR U2961 ( .A(n2804), .B(n2805), .Z(n2807) );
  NANDN U2962 ( .A(n2747), .B(n2746), .Z(n2751) );
  NANDN U2963 ( .A(n2749), .B(n2748), .Z(n2750) );
  AND U2964 ( .A(n2751), .B(n2750), .Z(n2806) );
  XOR U2965 ( .A(n2807), .B(n2806), .Z(n2813) );
  NAND U2966 ( .A(b[0]), .B(a[42]), .Z(n2752) );
  XNOR U2967 ( .A(b[1]), .B(n2752), .Z(n2754) );
  NAND U2968 ( .A(a[41]), .B(n206), .Z(n2753) );
  AND U2969 ( .A(n2754), .B(n2753), .Z(n2842) );
  XOR U2970 ( .A(n5129), .B(a[30]), .Z(n2851) );
  OR U2971 ( .A(n2851), .B(n5041), .Z(n2757) );
  NANDN U2972 ( .A(n2755), .B(n5052), .Z(n2756) );
  AND U2973 ( .A(n2757), .B(n2756), .Z(n2843) );
  XOR U2974 ( .A(n2842), .B(n2843), .Z(n2845) );
  NAND U2975 ( .A(b[15]), .B(a[26]), .Z(n2844) );
  XNOR U2976 ( .A(n2845), .B(n2844), .Z(n2836) );
  NAND U2977 ( .A(n4521), .B(n2758), .Z(n2760) );
  XOR U2978 ( .A(b[3]), .B(a[40]), .Z(n2854) );
  NANDN U2979 ( .A(n4488), .B(n2854), .Z(n2759) );
  NAND U2980 ( .A(n2760), .B(n2759), .Z(n2833) );
  XNOR U2981 ( .A(n209), .B(n3496), .Z(n2857) );
  OR U2982 ( .A(n2857), .B(n4612), .Z(n2763) );
  NANDN U2983 ( .A(n2761), .B(n4669), .Z(n2762) );
  NAND U2984 ( .A(n2763), .B(n2762), .Z(n2830) );
  XNOR U2985 ( .A(n4744), .B(n3347), .Z(n2860) );
  NANDN U2986 ( .A(n2860), .B(n4745), .Z(n2766) );
  NANDN U2987 ( .A(n2764), .B(n4746), .Z(n2765) );
  AND U2988 ( .A(n2766), .B(n2765), .Z(n2831) );
  XOR U2989 ( .A(n2833), .B(n2832), .Z(n2837) );
  XNOR U2990 ( .A(n2836), .B(n2837), .Z(n2838) );
  NANDN U2991 ( .A(n2768), .B(n2767), .Z(n2772) );
  NANDN U2992 ( .A(n2770), .B(n2769), .Z(n2771) );
  AND U2993 ( .A(n2772), .B(n2771), .Z(n2839) );
  XNOR U2994 ( .A(n2838), .B(n2839), .Z(n2811) );
  XNOR U2995 ( .A(n2811), .B(n2810), .Z(n2812) );
  XOR U2996 ( .A(n2813), .B(n2812), .Z(n2866) );
  NANDN U2997 ( .A(n2778), .B(n2777), .Z(n2782) );
  NANDN U2998 ( .A(n2780), .B(n2779), .Z(n2781) );
  NAND U2999 ( .A(n2782), .B(n2781), .Z(n2864) );
  NANDN U3000 ( .A(n2784), .B(n2783), .Z(n2788) );
  OR U3001 ( .A(n2786), .B(n2785), .Z(n2787) );
  AND U3002 ( .A(n2788), .B(n2787), .Z(n2863) );
  XNOR U3003 ( .A(n2864), .B(n2863), .Z(n2865) );
  XNOR U3004 ( .A(n2866), .B(n2865), .Z(n2800) );
  NANDN U3005 ( .A(n2790), .B(n2789), .Z(n2794) );
  NAND U3006 ( .A(n2792), .B(n2791), .Z(n2793) );
  NAND U3007 ( .A(n2794), .B(n2793), .Z(n2801) );
  XOR U3008 ( .A(n2800), .B(n2801), .Z(n2802) );
  XOR U3009 ( .A(n2803), .B(n2802), .Z(n2869) );
  XNOR U3010 ( .A(n2869), .B(sreg[90]), .Z(n2871) );
  NAND U3011 ( .A(n2795), .B(sreg[89]), .Z(n2799) );
  OR U3012 ( .A(n2797), .B(n2796), .Z(n2798) );
  AND U3013 ( .A(n2799), .B(n2798), .Z(n2870) );
  XOR U3014 ( .A(n2871), .B(n2870), .Z(c[90]) );
  NANDN U3015 ( .A(n2805), .B(n2804), .Z(n2809) );
  NANDN U3016 ( .A(n2807), .B(n2806), .Z(n2808) );
  NAND U3017 ( .A(n2809), .B(n2808), .Z(n2939) );
  NANDN U3018 ( .A(n2811), .B(n2810), .Z(n2815) );
  NANDN U3019 ( .A(n2813), .B(n2812), .Z(n2814) );
  AND U3020 ( .A(n2815), .B(n2814), .Z(n2938) );
  XNOR U3021 ( .A(n2939), .B(n2938), .Z(n2940) );
  XNOR U3022 ( .A(n4859), .B(n3273), .Z(n2880) );
  OR U3023 ( .A(n2880), .B(n4860), .Z(n2818) );
  NANDN U3024 ( .A(n2816), .B(n4915), .Z(n2817) );
  NAND U3025 ( .A(n2818), .B(n2817), .Z(n2892) );
  NANDN U3026 ( .A(n2819), .B(n4987), .Z(n2821) );
  XNOR U3027 ( .A(n4909), .B(n3121), .Z(n2883) );
  OR U3028 ( .A(n2883), .B(n4986), .Z(n2820) );
  NAND U3029 ( .A(n2821), .B(n2820), .Z(n2889) );
  XNOR U3030 ( .A(n210), .B(n2822), .Z(n2886) );
  OR U3031 ( .A(n2886), .B(n5095), .Z(n2825) );
  NANDN U3032 ( .A(n2823), .B(n5092), .Z(n2824) );
  AND U3033 ( .A(n2825), .B(n2824), .Z(n2890) );
  XOR U3034 ( .A(n2889), .B(n2890), .Z(n2891) );
  XOR U3035 ( .A(n2892), .B(n2891), .Z(n2932) );
  XNOR U3036 ( .A(n2932), .B(n2933), .Z(n2934) );
  NANDN U3037 ( .A(n2831), .B(n2830), .Z(n2835) );
  NAND U3038 ( .A(n2833), .B(n2832), .Z(n2834) );
  NAND U3039 ( .A(n2835), .B(n2834), .Z(n2935) );
  XOR U3040 ( .A(n2934), .B(n2935), .Z(n2929) );
  NANDN U3041 ( .A(n2837), .B(n2836), .Z(n2841) );
  NAND U3042 ( .A(n2839), .B(n2838), .Z(n2840) );
  NAND U3043 ( .A(n2841), .B(n2840), .Z(n2927) );
  NANDN U3044 ( .A(n2843), .B(n2842), .Z(n2847) );
  OR U3045 ( .A(n2845), .B(n2844), .Z(n2846) );
  NAND U3046 ( .A(n2847), .B(n2846), .Z(n2902) );
  NAND U3047 ( .A(b[0]), .B(a[43]), .Z(n2848) );
  XNOR U3048 ( .A(b[1]), .B(n2848), .Z(n2850) );
  NAND U3049 ( .A(a[42]), .B(n206), .Z(n2849) );
  AND U3050 ( .A(n2850), .B(n2849), .Z(n2905) );
  XNOR U3051 ( .A(n5129), .B(n2971), .Z(n2911) );
  OR U3052 ( .A(n2911), .B(n5041), .Z(n2853) );
  NANDN U3053 ( .A(n2851), .B(n5052), .Z(n2852) );
  AND U3054 ( .A(n2853), .B(n2852), .Z(n2906) );
  XOR U3055 ( .A(n2905), .B(n2906), .Z(n2908) );
  NAND U3056 ( .A(a[27]), .B(b[15]), .Z(n2907) );
  XOR U3057 ( .A(n2908), .B(n2907), .Z(n2899) );
  NAND U3058 ( .A(n4521), .B(n2854), .Z(n2856) );
  IV U3059 ( .A(a[41]), .Z(n3736) );
  XNOR U3060 ( .A(b[3]), .B(n3736), .Z(n2917) );
  NANDN U3061 ( .A(n4488), .B(n2917), .Z(n2855) );
  NAND U3062 ( .A(n2856), .B(n2855), .Z(n2895) );
  XNOR U3063 ( .A(n209), .B(n3560), .Z(n2920) );
  OR U3064 ( .A(n2920), .B(n4612), .Z(n2859) );
  NANDN U3065 ( .A(n2857), .B(n4669), .Z(n2858) );
  NAND U3066 ( .A(n2859), .B(n2858), .Z(n2893) );
  XOR U3067 ( .A(n4744), .B(a[37]), .Z(n2923) );
  NANDN U3068 ( .A(n2923), .B(n4745), .Z(n2862) );
  NANDN U3069 ( .A(n2860), .B(n4746), .Z(n2861) );
  AND U3070 ( .A(n2862), .B(n2861), .Z(n2894) );
  XOR U3071 ( .A(n2895), .B(n2896), .Z(n2900) );
  XNOR U3072 ( .A(n2899), .B(n2900), .Z(n2901) );
  XOR U3073 ( .A(n2902), .B(n2901), .Z(n2926) );
  XNOR U3074 ( .A(n2927), .B(n2926), .Z(n2928) );
  XNOR U3075 ( .A(n2929), .B(n2928), .Z(n2941) );
  XOR U3076 ( .A(n2940), .B(n2941), .Z(n2874) );
  NANDN U3077 ( .A(n2864), .B(n2863), .Z(n2868) );
  NAND U3078 ( .A(n2866), .B(n2865), .Z(n2867) );
  NAND U3079 ( .A(n2868), .B(n2867), .Z(n2875) );
  XNOR U3080 ( .A(n2874), .B(n2875), .Z(n2876) );
  XNOR U3081 ( .A(n2877), .B(n2876), .Z(n2944) );
  XNOR U3082 ( .A(n2944), .B(sreg[91]), .Z(n2946) );
  NAND U3083 ( .A(n2869), .B(sreg[90]), .Z(n2873) );
  OR U3084 ( .A(n2871), .B(n2870), .Z(n2872) );
  AND U3085 ( .A(n2873), .B(n2872), .Z(n2945) );
  XOR U3086 ( .A(n2946), .B(n2945), .Z(c[91]) );
  NANDN U3087 ( .A(n2875), .B(n2874), .Z(n2879) );
  NAND U3088 ( .A(n2877), .B(n2876), .Z(n2878) );
  NAND U3089 ( .A(n2879), .B(n2878), .Z(n2952) );
  XNOR U3090 ( .A(n4859), .B(n3347), .Z(n2965) );
  OR U3091 ( .A(n2965), .B(n4860), .Z(n2882) );
  NANDN U3092 ( .A(n2880), .B(n4915), .Z(n2881) );
  NAND U3093 ( .A(n2882), .B(n2881), .Z(n2978) );
  NANDN U3094 ( .A(n2883), .B(n4987), .Z(n2885) );
  XNOR U3095 ( .A(n4909), .B(n3197), .Z(n2968) );
  OR U3096 ( .A(n2968), .B(n4986), .Z(n2884) );
  NAND U3097 ( .A(n2885), .B(n2884), .Z(n2975) );
  XOR U3098 ( .A(n210), .B(a[30]), .Z(n2972) );
  OR U3099 ( .A(n2972), .B(n5095), .Z(n2888) );
  NANDN U3100 ( .A(n2886), .B(n5092), .Z(n2887) );
  AND U3101 ( .A(n2888), .B(n2887), .Z(n2976) );
  XOR U3102 ( .A(n2975), .B(n2976), .Z(n2977) );
  XOR U3103 ( .A(n2978), .B(n2977), .Z(n2959) );
  XNOR U3104 ( .A(n2959), .B(n2960), .Z(n2961) );
  NANDN U3105 ( .A(n2894), .B(n2893), .Z(n2898) );
  NANDN U3106 ( .A(n2896), .B(n2895), .Z(n2897) );
  NAND U3107 ( .A(n2898), .B(n2897), .Z(n2962) );
  XOR U3108 ( .A(n2961), .B(n2962), .Z(n2955) );
  NANDN U3109 ( .A(n2900), .B(n2899), .Z(n2904) );
  NAND U3110 ( .A(n2902), .B(n2901), .Z(n2903) );
  NAND U3111 ( .A(n2904), .B(n2903), .Z(n2954) );
  NANDN U3112 ( .A(n2906), .B(n2905), .Z(n2910) );
  OR U3113 ( .A(n2908), .B(n2907), .Z(n2909) );
  NAND U3114 ( .A(n2910), .B(n2909), .Z(n2986) );
  XNOR U3115 ( .A(n5129), .B(n3035), .Z(n3000) );
  OR U3116 ( .A(n3000), .B(n5041), .Z(n2913) );
  NANDN U3117 ( .A(n2911), .B(n5052), .Z(n2912) );
  AND U3118 ( .A(n2913), .B(n2912), .Z(n2992) );
  NAND U3119 ( .A(b[0]), .B(a[44]), .Z(n2914) );
  XNOR U3120 ( .A(b[1]), .B(n2914), .Z(n2916) );
  NAND U3121 ( .A(a[43]), .B(n206), .Z(n2915) );
  AND U3122 ( .A(n2916), .B(n2915), .Z(n2991) );
  XOR U3123 ( .A(n2992), .B(n2991), .Z(n2994) );
  NAND U3124 ( .A(a[28]), .B(b[15]), .Z(n2993) );
  XOR U3125 ( .A(n2994), .B(n2993), .Z(n2985) );
  XNOR U3126 ( .A(n2986), .B(n2985), .Z(n2987) );
  NAND U3127 ( .A(n4521), .B(n2917), .Z(n2919) );
  IV U3128 ( .A(a[42]), .Z(n3781) );
  XNOR U3129 ( .A(b[3]), .B(n3781), .Z(n3003) );
  NANDN U3130 ( .A(n4488), .B(n3003), .Z(n2918) );
  NAND U3131 ( .A(n2919), .B(n2918), .Z(n2981) );
  XOR U3132 ( .A(n209), .B(a[40]), .Z(n3006) );
  OR U3133 ( .A(n3006), .B(n4612), .Z(n2922) );
  NANDN U3134 ( .A(n2920), .B(n4669), .Z(n2921) );
  NAND U3135 ( .A(n2922), .B(n2921), .Z(n2979) );
  XNOR U3136 ( .A(n4744), .B(n3496), .Z(n3009) );
  NANDN U3137 ( .A(n3009), .B(n4745), .Z(n2925) );
  NANDN U3138 ( .A(n2923), .B(n4746), .Z(n2924) );
  AND U3139 ( .A(n2925), .B(n2924), .Z(n2980) );
  XOR U3140 ( .A(n2981), .B(n2982), .Z(n2988) );
  XOR U3141 ( .A(n2987), .B(n2988), .Z(n2953) );
  XNOR U3142 ( .A(n2954), .B(n2953), .Z(n2956) );
  XNOR U3143 ( .A(n2955), .B(n2956), .Z(n3014) );
  NANDN U3144 ( .A(n2927), .B(n2926), .Z(n2931) );
  NAND U3145 ( .A(n2929), .B(n2928), .Z(n2930) );
  NAND U3146 ( .A(n2931), .B(n2930), .Z(n3012) );
  NANDN U3147 ( .A(n2933), .B(n2932), .Z(n2937) );
  NANDN U3148 ( .A(n2935), .B(n2934), .Z(n2936) );
  NAND U3149 ( .A(n2937), .B(n2936), .Z(n3013) );
  XNOR U3150 ( .A(n3012), .B(n3013), .Z(n3015) );
  XOR U3151 ( .A(n3014), .B(n3015), .Z(n2949) );
  NANDN U3152 ( .A(n2939), .B(n2938), .Z(n2943) );
  NANDN U3153 ( .A(n2941), .B(n2940), .Z(n2942) );
  NAND U3154 ( .A(n2943), .B(n2942), .Z(n2950) );
  XOR U3155 ( .A(n2949), .B(n2950), .Z(n2951) );
  XNOR U3156 ( .A(n2952), .B(n2951), .Z(n3018) );
  XNOR U3157 ( .A(n3018), .B(sreg[92]), .Z(n3020) );
  NAND U3158 ( .A(n2944), .B(sreg[91]), .Z(n2948) );
  OR U3159 ( .A(n2946), .B(n2945), .Z(n2947) );
  AND U3160 ( .A(n2948), .B(n2947), .Z(n3019) );
  XOR U3161 ( .A(n3020), .B(n3019), .Z(c[92]) );
  NAND U3162 ( .A(n2954), .B(n2953), .Z(n2958) );
  NANDN U3163 ( .A(n2956), .B(n2955), .Z(n2957) );
  NAND U3164 ( .A(n2958), .B(n2957), .Z(n3088) );
  NANDN U3165 ( .A(n2960), .B(n2959), .Z(n2964) );
  NANDN U3166 ( .A(n2962), .B(n2961), .Z(n2963) );
  NAND U3167 ( .A(n2964), .B(n2963), .Z(n3089) );
  XNOR U3168 ( .A(n3088), .B(n3089), .Z(n3090) );
  XOR U3169 ( .A(n4859), .B(a[37]), .Z(n3029) );
  OR U3170 ( .A(n3029), .B(n4860), .Z(n2967) );
  NANDN U3171 ( .A(n2965), .B(n4915), .Z(n2966) );
  NAND U3172 ( .A(n2967), .B(n2966), .Z(n3042) );
  NANDN U3173 ( .A(n2968), .B(n4987), .Z(n2970) );
  XNOR U3174 ( .A(n4909), .B(n3273), .Z(n3032) );
  OR U3175 ( .A(n3032), .B(n4986), .Z(n2969) );
  NAND U3176 ( .A(n2970), .B(n2969), .Z(n3039) );
  XNOR U3177 ( .A(n210), .B(n2971), .Z(n3036) );
  OR U3178 ( .A(n3036), .B(n5095), .Z(n2974) );
  NANDN U3179 ( .A(n2972), .B(n5092), .Z(n2973) );
  AND U3180 ( .A(n2974), .B(n2973), .Z(n3040) );
  XOR U3181 ( .A(n3039), .B(n3040), .Z(n3041) );
  XOR U3182 ( .A(n3042), .B(n3041), .Z(n3082) );
  XNOR U3183 ( .A(n3082), .B(n3083), .Z(n3084) );
  NANDN U3184 ( .A(n2980), .B(n2979), .Z(n2984) );
  NANDN U3185 ( .A(n2982), .B(n2981), .Z(n2983) );
  NAND U3186 ( .A(n2984), .B(n2983), .Z(n3085) );
  XOR U3187 ( .A(n3084), .B(n3085), .Z(n3079) );
  NAND U3188 ( .A(n2986), .B(n2985), .Z(n2990) );
  OR U3189 ( .A(n2988), .B(n2987), .Z(n2989) );
  NAND U3190 ( .A(n2990), .B(n2989), .Z(n3076) );
  NANDN U3191 ( .A(n2992), .B(n2991), .Z(n2996) );
  OR U3192 ( .A(n2994), .B(n2993), .Z(n2995) );
  NAND U3193 ( .A(n2996), .B(n2995), .Z(n3073) );
  NAND U3194 ( .A(b[0]), .B(a[45]), .Z(n2997) );
  XNOR U3195 ( .A(b[1]), .B(n2997), .Z(n2999) );
  NAND U3196 ( .A(n206), .B(a[44]), .Z(n2998) );
  AND U3197 ( .A(n2999), .B(n2998), .Z(n3064) );
  XNOR U3198 ( .A(n5129), .B(n3121), .Z(n3052) );
  OR U3199 ( .A(n3052), .B(n5041), .Z(n3002) );
  NANDN U3200 ( .A(n3000), .B(n5052), .Z(n3001) );
  AND U3201 ( .A(n3002), .B(n3001), .Z(n3065) );
  XOR U3202 ( .A(n3064), .B(n3065), .Z(n3067) );
  NAND U3203 ( .A(a[29]), .B(b[15]), .Z(n3066) );
  XOR U3204 ( .A(n3067), .B(n3066), .Z(n3070) );
  NAND U3205 ( .A(n4521), .B(n3003), .Z(n3005) );
  IV U3206 ( .A(a[43]), .Z(n3865) );
  XNOR U3207 ( .A(b[3]), .B(n3865), .Z(n3055) );
  NANDN U3208 ( .A(n4488), .B(n3055), .Z(n3004) );
  NAND U3209 ( .A(n3005), .B(n3004), .Z(n3045) );
  XNOR U3210 ( .A(n209), .B(n3736), .Z(n3058) );
  OR U3211 ( .A(n3058), .B(n4612), .Z(n3008) );
  NANDN U3212 ( .A(n3006), .B(n4669), .Z(n3007) );
  NAND U3213 ( .A(n3008), .B(n3007), .Z(n3043) );
  XNOR U3214 ( .A(n4744), .B(n3560), .Z(n3061) );
  NANDN U3215 ( .A(n3061), .B(n4745), .Z(n3011) );
  NANDN U3216 ( .A(n3009), .B(n4746), .Z(n3010) );
  AND U3217 ( .A(n3011), .B(n3010), .Z(n3044) );
  XOR U3218 ( .A(n3045), .B(n3046), .Z(n3071) );
  XNOR U3219 ( .A(n3070), .B(n3071), .Z(n3072) );
  XNOR U3220 ( .A(n3073), .B(n3072), .Z(n3077) );
  XNOR U3221 ( .A(n3076), .B(n3077), .Z(n3078) );
  XNOR U3222 ( .A(n3079), .B(n3078), .Z(n3091) );
  XOR U3223 ( .A(n3090), .B(n3091), .Z(n3023) );
  NANDN U3224 ( .A(n3013), .B(n3012), .Z(n3017) );
  NAND U3225 ( .A(n3015), .B(n3014), .Z(n3016) );
  NAND U3226 ( .A(n3017), .B(n3016), .Z(n3024) );
  XNOR U3227 ( .A(n3023), .B(n3024), .Z(n3025) );
  XNOR U3228 ( .A(n3026), .B(n3025), .Z(n3094) );
  XNOR U3229 ( .A(n3094), .B(sreg[93]), .Z(n3096) );
  NAND U3230 ( .A(n3018), .B(sreg[92]), .Z(n3022) );
  OR U3231 ( .A(n3020), .B(n3019), .Z(n3021) );
  AND U3232 ( .A(n3022), .B(n3021), .Z(n3095) );
  XOR U3233 ( .A(n3096), .B(n3095), .Z(c[93]) );
  NANDN U3234 ( .A(n3024), .B(n3023), .Z(n3028) );
  NAND U3235 ( .A(n3026), .B(n3025), .Z(n3027) );
  NAND U3236 ( .A(n3028), .B(n3027), .Z(n3102) );
  XNOR U3237 ( .A(n4859), .B(n3496), .Z(n3115) );
  OR U3238 ( .A(n3115), .B(n4860), .Z(n3031) );
  NANDN U3239 ( .A(n3029), .B(n4915), .Z(n3030) );
  NAND U3240 ( .A(n3031), .B(n3030), .Z(n3128) );
  NANDN U3241 ( .A(n3032), .B(n4987), .Z(n3034) );
  XNOR U3242 ( .A(n4909), .B(n3347), .Z(n3118) );
  OR U3243 ( .A(n3118), .B(n4986), .Z(n3033) );
  NAND U3244 ( .A(n3034), .B(n3033), .Z(n3125) );
  XNOR U3245 ( .A(n210), .B(n3035), .Z(n3122) );
  OR U3246 ( .A(n3122), .B(n5095), .Z(n3038) );
  NANDN U3247 ( .A(n3036), .B(n5092), .Z(n3037) );
  AND U3248 ( .A(n3038), .B(n3037), .Z(n3126) );
  XOR U3249 ( .A(n3125), .B(n3126), .Z(n3127) );
  XOR U3250 ( .A(n3128), .B(n3127), .Z(n3103) );
  XOR U3251 ( .A(n3103), .B(n3104), .Z(n3106) );
  NANDN U3252 ( .A(n3044), .B(n3043), .Z(n3048) );
  NANDN U3253 ( .A(n3046), .B(n3045), .Z(n3047) );
  AND U3254 ( .A(n3048), .B(n3047), .Z(n3105) );
  XOR U3255 ( .A(n3106), .B(n3105), .Z(n3112) );
  NAND U3256 ( .A(b[0]), .B(a[46]), .Z(n3049) );
  XNOR U3257 ( .A(b[1]), .B(n3049), .Z(n3051) );
  NAND U3258 ( .A(n206), .B(a[45]), .Z(n3050) );
  AND U3259 ( .A(n3051), .B(n3050), .Z(n3135) );
  XNOR U3260 ( .A(n5129), .B(n3197), .Z(n3144) );
  OR U3261 ( .A(n3144), .B(n5041), .Z(n3054) );
  NANDN U3262 ( .A(n3052), .B(n5052), .Z(n3053) );
  AND U3263 ( .A(n3054), .B(n3053), .Z(n3136) );
  XOR U3264 ( .A(n3135), .B(n3136), .Z(n3138) );
  NAND U3265 ( .A(b[15]), .B(a[30]), .Z(n3137) );
  XNOR U3266 ( .A(n3138), .B(n3137), .Z(n3156) );
  NAND U3267 ( .A(n4521), .B(n3055), .Z(n3057) );
  XOR U3268 ( .A(b[3]), .B(a[44]), .Z(n3147) );
  NANDN U3269 ( .A(n4488), .B(n3147), .Z(n3056) );
  NAND U3270 ( .A(n3057), .B(n3056), .Z(n3132) );
  XNOR U3271 ( .A(n209), .B(n3781), .Z(n3150) );
  OR U3272 ( .A(n3150), .B(n4612), .Z(n3060) );
  NANDN U3273 ( .A(n3058), .B(n4669), .Z(n3059) );
  NAND U3274 ( .A(n3060), .B(n3059), .Z(n3129) );
  XOR U3275 ( .A(n4744), .B(a[40]), .Z(n3153) );
  NANDN U3276 ( .A(n3153), .B(n4745), .Z(n3063) );
  NANDN U3277 ( .A(n3061), .B(n4746), .Z(n3062) );
  AND U3278 ( .A(n3063), .B(n3062), .Z(n3130) );
  XOR U3279 ( .A(n3132), .B(n3131), .Z(n3157) );
  XNOR U3280 ( .A(n3156), .B(n3157), .Z(n3158) );
  NANDN U3281 ( .A(n3065), .B(n3064), .Z(n3069) );
  OR U3282 ( .A(n3067), .B(n3066), .Z(n3068) );
  AND U3283 ( .A(n3069), .B(n3068), .Z(n3159) );
  XNOR U3284 ( .A(n3158), .B(n3159), .Z(n3110) );
  NANDN U3285 ( .A(n3071), .B(n3070), .Z(n3075) );
  NAND U3286 ( .A(n3073), .B(n3072), .Z(n3074) );
  AND U3287 ( .A(n3075), .B(n3074), .Z(n3109) );
  XNOR U3288 ( .A(n3110), .B(n3109), .Z(n3111) );
  XOR U3289 ( .A(n3112), .B(n3111), .Z(n3165) );
  NANDN U3290 ( .A(n3077), .B(n3076), .Z(n3081) );
  NAND U3291 ( .A(n3079), .B(n3078), .Z(n3080) );
  NAND U3292 ( .A(n3081), .B(n3080), .Z(n3162) );
  NANDN U3293 ( .A(n3083), .B(n3082), .Z(n3087) );
  NANDN U3294 ( .A(n3085), .B(n3084), .Z(n3086) );
  NAND U3295 ( .A(n3087), .B(n3086), .Z(n3163) );
  XNOR U3296 ( .A(n3162), .B(n3163), .Z(n3164) );
  XNOR U3297 ( .A(n3165), .B(n3164), .Z(n3099) );
  NANDN U3298 ( .A(n3089), .B(n3088), .Z(n3093) );
  NANDN U3299 ( .A(n3091), .B(n3090), .Z(n3092) );
  NAND U3300 ( .A(n3093), .B(n3092), .Z(n3100) );
  XOR U3301 ( .A(n3099), .B(n3100), .Z(n3101) );
  XOR U3302 ( .A(n3102), .B(n3101), .Z(n3168) );
  XNOR U3303 ( .A(n3168), .B(sreg[94]), .Z(n3170) );
  NAND U3304 ( .A(n3094), .B(sreg[93]), .Z(n3098) );
  OR U3305 ( .A(n3096), .B(n3095), .Z(n3097) );
  AND U3306 ( .A(n3098), .B(n3097), .Z(n3169) );
  XOR U3307 ( .A(n3170), .B(n3169), .Z(c[94]) );
  NANDN U3308 ( .A(n3104), .B(n3103), .Z(n3108) );
  NANDN U3309 ( .A(n3106), .B(n3105), .Z(n3107) );
  NAND U3310 ( .A(n3108), .B(n3107), .Z(n3239) );
  NANDN U3311 ( .A(n3110), .B(n3109), .Z(n3114) );
  NANDN U3312 ( .A(n3112), .B(n3111), .Z(n3113) );
  AND U3313 ( .A(n3114), .B(n3113), .Z(n3238) );
  XNOR U3314 ( .A(n3239), .B(n3238), .Z(n3240) );
  XNOR U3315 ( .A(n4859), .B(n3560), .Z(n3191) );
  OR U3316 ( .A(n3191), .B(n4860), .Z(n3117) );
  NANDN U3317 ( .A(n3115), .B(n4915), .Z(n3116) );
  NAND U3318 ( .A(n3117), .B(n3116), .Z(n3204) );
  NANDN U3319 ( .A(n3118), .B(n4987), .Z(n3120) );
  XOR U3320 ( .A(n4909), .B(a[37]), .Z(n3194) );
  OR U3321 ( .A(n3194), .B(n4986), .Z(n3119) );
  NAND U3322 ( .A(n3120), .B(n3119), .Z(n3201) );
  XNOR U3323 ( .A(n210), .B(n3121), .Z(n3198) );
  OR U3324 ( .A(n3198), .B(n5095), .Z(n3124) );
  NANDN U3325 ( .A(n3122), .B(n5092), .Z(n3123) );
  AND U3326 ( .A(n3124), .B(n3123), .Z(n3202) );
  XOR U3327 ( .A(n3201), .B(n3202), .Z(n3203) );
  XOR U3328 ( .A(n3204), .B(n3203), .Z(n3185) );
  XNOR U3329 ( .A(n3185), .B(n3186), .Z(n3187) );
  NANDN U3330 ( .A(n3130), .B(n3129), .Z(n3134) );
  NAND U3331 ( .A(n3132), .B(n3131), .Z(n3133) );
  NAND U3332 ( .A(n3134), .B(n3133), .Z(n3188) );
  XOR U3333 ( .A(n3187), .B(n3188), .Z(n3182) );
  NANDN U3334 ( .A(n3136), .B(n3135), .Z(n3140) );
  OR U3335 ( .A(n3138), .B(n3137), .Z(n3139) );
  NAND U3336 ( .A(n3140), .B(n3139), .Z(n3214) );
  NAND U3337 ( .A(b[0]), .B(a[47]), .Z(n3141) );
  XNOR U3338 ( .A(b[1]), .B(n3141), .Z(n3143) );
  NAND U3339 ( .A(a[46]), .B(n206), .Z(n3142) );
  AND U3340 ( .A(n3143), .B(n3142), .Z(n3217) );
  XNOR U3341 ( .A(n5129), .B(n3273), .Z(n3226) );
  OR U3342 ( .A(n3226), .B(n5041), .Z(n3146) );
  NANDN U3343 ( .A(n3144), .B(n5052), .Z(n3145) );
  AND U3344 ( .A(n3146), .B(n3145), .Z(n3218) );
  XOR U3345 ( .A(n3217), .B(n3218), .Z(n3220) );
  NAND U3346 ( .A(a[31]), .B(b[15]), .Z(n3219) );
  XOR U3347 ( .A(n3220), .B(n3219), .Z(n3211) );
  NAND U3348 ( .A(n4521), .B(n3147), .Z(n3149) );
  XOR U3349 ( .A(b[3]), .B(a[45]), .Z(n3229) );
  NANDN U3350 ( .A(n4488), .B(n3229), .Z(n3148) );
  NAND U3351 ( .A(n3149), .B(n3148), .Z(n3207) );
  XNOR U3352 ( .A(n209), .B(n3865), .Z(n3232) );
  OR U3353 ( .A(n3232), .B(n4612), .Z(n3152) );
  NANDN U3354 ( .A(n3150), .B(n4669), .Z(n3151) );
  NAND U3355 ( .A(n3152), .B(n3151), .Z(n3205) );
  XNOR U3356 ( .A(n4744), .B(n3736), .Z(n3235) );
  NANDN U3357 ( .A(n3235), .B(n4745), .Z(n3155) );
  NANDN U3358 ( .A(n3153), .B(n4746), .Z(n3154) );
  AND U3359 ( .A(n3155), .B(n3154), .Z(n3206) );
  XOR U3360 ( .A(n3207), .B(n3208), .Z(n3212) );
  XNOR U3361 ( .A(n3211), .B(n3212), .Z(n3213) );
  XNOR U3362 ( .A(n3214), .B(n3213), .Z(n3180) );
  NANDN U3363 ( .A(n3157), .B(n3156), .Z(n3161) );
  NAND U3364 ( .A(n3159), .B(n3158), .Z(n3160) );
  AND U3365 ( .A(n3161), .B(n3160), .Z(n3179) );
  XNOR U3366 ( .A(n3180), .B(n3179), .Z(n3181) );
  XNOR U3367 ( .A(n3182), .B(n3181), .Z(n3241) );
  XOR U3368 ( .A(n3240), .B(n3241), .Z(n3173) );
  NANDN U3369 ( .A(n3163), .B(n3162), .Z(n3167) );
  NAND U3370 ( .A(n3165), .B(n3164), .Z(n3166) );
  NAND U3371 ( .A(n3167), .B(n3166), .Z(n3174) );
  XNOR U3372 ( .A(n3173), .B(n3174), .Z(n3175) );
  XNOR U3373 ( .A(n3176), .B(n3175), .Z(n3244) );
  XNOR U3374 ( .A(n3244), .B(sreg[95]), .Z(n3246) );
  NAND U3375 ( .A(n3168), .B(sreg[94]), .Z(n3172) );
  OR U3376 ( .A(n3170), .B(n3169), .Z(n3171) );
  AND U3377 ( .A(n3172), .B(n3171), .Z(n3245) );
  XOR U3378 ( .A(n3246), .B(n3245), .Z(c[95]) );
  NANDN U3379 ( .A(n3174), .B(n3173), .Z(n3178) );
  NAND U3380 ( .A(n3176), .B(n3175), .Z(n3177) );
  NAND U3381 ( .A(n3178), .B(n3177), .Z(n3252) );
  NANDN U3382 ( .A(n3180), .B(n3179), .Z(n3184) );
  NAND U3383 ( .A(n3182), .B(n3181), .Z(n3183) );
  NAND U3384 ( .A(n3184), .B(n3183), .Z(n3314) );
  NANDN U3385 ( .A(n3186), .B(n3185), .Z(n3190) );
  NANDN U3386 ( .A(n3188), .B(n3187), .Z(n3189) );
  NAND U3387 ( .A(n3190), .B(n3189), .Z(n3315) );
  XNOR U3388 ( .A(n3314), .B(n3315), .Z(n3316) );
  XOR U3389 ( .A(n4859), .B(a[40]), .Z(n3267) );
  OR U3390 ( .A(n3267), .B(n4860), .Z(n3193) );
  NANDN U3391 ( .A(n3191), .B(n4915), .Z(n3192) );
  NAND U3392 ( .A(n3193), .B(n3192), .Z(n3280) );
  NANDN U3393 ( .A(n3194), .B(n4987), .Z(n3196) );
  XNOR U3394 ( .A(n4909), .B(n3496), .Z(n3270) );
  OR U3395 ( .A(n3270), .B(n4986), .Z(n3195) );
  NAND U3396 ( .A(n3196), .B(n3195), .Z(n3277) );
  XNOR U3397 ( .A(n210), .B(n3197), .Z(n3274) );
  OR U3398 ( .A(n3274), .B(n5095), .Z(n3200) );
  NANDN U3399 ( .A(n3198), .B(n5092), .Z(n3199) );
  AND U3400 ( .A(n3200), .B(n3199), .Z(n3278) );
  XOR U3401 ( .A(n3277), .B(n3278), .Z(n3279) );
  XOR U3402 ( .A(n3280), .B(n3279), .Z(n3261) );
  XNOR U3403 ( .A(n3261), .B(n3262), .Z(n3263) );
  NANDN U3404 ( .A(n3206), .B(n3205), .Z(n3210) );
  NANDN U3405 ( .A(n3208), .B(n3207), .Z(n3209) );
  NAND U3406 ( .A(n3210), .B(n3209), .Z(n3264) );
  XOR U3407 ( .A(n3263), .B(n3264), .Z(n3258) );
  NANDN U3408 ( .A(n3212), .B(n3211), .Z(n3216) );
  NAND U3409 ( .A(n3214), .B(n3213), .Z(n3215) );
  NAND U3410 ( .A(n3216), .B(n3215), .Z(n3255) );
  NANDN U3411 ( .A(n3218), .B(n3217), .Z(n3222) );
  OR U3412 ( .A(n3220), .B(n3219), .Z(n3221) );
  NAND U3413 ( .A(n3222), .B(n3221), .Z(n3290) );
  NAND U3414 ( .A(b[0]), .B(a[48]), .Z(n3223) );
  XNOR U3415 ( .A(b[1]), .B(n3223), .Z(n3225) );
  NAND U3416 ( .A(n206), .B(a[47]), .Z(n3224) );
  AND U3417 ( .A(n3225), .B(n3224), .Z(n3293) );
  XNOR U3418 ( .A(n5129), .B(n3347), .Z(n3299) );
  OR U3419 ( .A(n3299), .B(n5041), .Z(n3228) );
  NANDN U3420 ( .A(n3226), .B(n5052), .Z(n3227) );
  AND U3421 ( .A(n3228), .B(n3227), .Z(n3294) );
  XOR U3422 ( .A(n3293), .B(n3294), .Z(n3296) );
  NAND U3423 ( .A(a[32]), .B(b[15]), .Z(n3295) );
  XOR U3424 ( .A(n3296), .B(n3295), .Z(n3287) );
  NAND U3425 ( .A(n4521), .B(n3229), .Z(n3231) );
  IV U3426 ( .A(a[46]), .Z(n4089) );
  XNOR U3427 ( .A(b[3]), .B(n4089), .Z(n3305) );
  NANDN U3428 ( .A(n4488), .B(n3305), .Z(n3230) );
  NAND U3429 ( .A(n3231), .B(n3230), .Z(n3283) );
  XOR U3430 ( .A(n209), .B(a[44]), .Z(n3308) );
  OR U3431 ( .A(n3308), .B(n4612), .Z(n3234) );
  NANDN U3432 ( .A(n3232), .B(n4669), .Z(n3233) );
  NAND U3433 ( .A(n3234), .B(n3233), .Z(n3281) );
  XNOR U3434 ( .A(n4744), .B(n3781), .Z(n3311) );
  NANDN U3435 ( .A(n3311), .B(n4745), .Z(n3237) );
  NANDN U3436 ( .A(n3235), .B(n4746), .Z(n3236) );
  AND U3437 ( .A(n3237), .B(n3236), .Z(n3282) );
  XOR U3438 ( .A(n3283), .B(n3284), .Z(n3288) );
  XNOR U3439 ( .A(n3287), .B(n3288), .Z(n3289) );
  XNOR U3440 ( .A(n3290), .B(n3289), .Z(n3256) );
  XNOR U3441 ( .A(n3255), .B(n3256), .Z(n3257) );
  XNOR U3442 ( .A(n3258), .B(n3257), .Z(n3317) );
  XOR U3443 ( .A(n3316), .B(n3317), .Z(n3249) );
  NANDN U3444 ( .A(n3239), .B(n3238), .Z(n3243) );
  NANDN U3445 ( .A(n3241), .B(n3240), .Z(n3242) );
  NAND U3446 ( .A(n3243), .B(n3242), .Z(n3250) );
  XNOR U3447 ( .A(n3249), .B(n3250), .Z(n3251) );
  XNOR U3448 ( .A(n3252), .B(n3251), .Z(n3320) );
  XNOR U3449 ( .A(n3320), .B(sreg[96]), .Z(n3322) );
  NAND U3450 ( .A(n3244), .B(sreg[95]), .Z(n3248) );
  OR U3451 ( .A(n3246), .B(n3245), .Z(n3247) );
  AND U3452 ( .A(n3248), .B(n3247), .Z(n3321) );
  XOR U3453 ( .A(n3322), .B(n3321), .Z(c[96]) );
  NANDN U3454 ( .A(n3250), .B(n3249), .Z(n3254) );
  NAND U3455 ( .A(n3252), .B(n3251), .Z(n3253) );
  NAND U3456 ( .A(n3254), .B(n3253), .Z(n3328) );
  NANDN U3457 ( .A(n3256), .B(n3255), .Z(n3260) );
  NAND U3458 ( .A(n3258), .B(n3257), .Z(n3259) );
  NAND U3459 ( .A(n3260), .B(n3259), .Z(n3388) );
  NANDN U3460 ( .A(n3262), .B(n3261), .Z(n3266) );
  NANDN U3461 ( .A(n3264), .B(n3263), .Z(n3265) );
  NAND U3462 ( .A(n3266), .B(n3265), .Z(n3389) );
  XNOR U3463 ( .A(n3388), .B(n3389), .Z(n3390) );
  XNOR U3464 ( .A(n4859), .B(n3736), .Z(n3341) );
  OR U3465 ( .A(n3341), .B(n4860), .Z(n3269) );
  NANDN U3466 ( .A(n3267), .B(n4915), .Z(n3268) );
  NAND U3467 ( .A(n3269), .B(n3268), .Z(n3354) );
  NANDN U3468 ( .A(n3270), .B(n4987), .Z(n3272) );
  XNOR U3469 ( .A(n4909), .B(n3560), .Z(n3344) );
  OR U3470 ( .A(n3344), .B(n4986), .Z(n3271) );
  NAND U3471 ( .A(n3272), .B(n3271), .Z(n3351) );
  XNOR U3472 ( .A(n210), .B(n3273), .Z(n3348) );
  OR U3473 ( .A(n3348), .B(n5095), .Z(n3276) );
  NANDN U3474 ( .A(n3274), .B(n5092), .Z(n3275) );
  AND U3475 ( .A(n3276), .B(n3275), .Z(n3352) );
  XOR U3476 ( .A(n3351), .B(n3352), .Z(n3353) );
  XOR U3477 ( .A(n3354), .B(n3353), .Z(n3335) );
  XNOR U3478 ( .A(n3335), .B(n3336), .Z(n3337) );
  NANDN U3479 ( .A(n3282), .B(n3281), .Z(n3286) );
  NANDN U3480 ( .A(n3284), .B(n3283), .Z(n3285) );
  NAND U3481 ( .A(n3286), .B(n3285), .Z(n3338) );
  XOR U3482 ( .A(n3337), .B(n3338), .Z(n3331) );
  NANDN U3483 ( .A(n3288), .B(n3287), .Z(n3292) );
  NAND U3484 ( .A(n3290), .B(n3289), .Z(n3291) );
  NAND U3485 ( .A(n3292), .B(n3291), .Z(n3330) );
  NANDN U3486 ( .A(n3294), .B(n3293), .Z(n3298) );
  OR U3487 ( .A(n3296), .B(n3295), .Z(n3297) );
  NAND U3488 ( .A(n3298), .B(n3297), .Z(n3362) );
  XOR U3489 ( .A(n5129), .B(a[37]), .Z(n3376) );
  OR U3490 ( .A(n3376), .B(n5041), .Z(n3301) );
  NANDN U3491 ( .A(n3299), .B(n5052), .Z(n3300) );
  AND U3492 ( .A(n3301), .B(n3300), .Z(n3368) );
  NAND U3493 ( .A(b[0]), .B(a[49]), .Z(n3302) );
  XNOR U3494 ( .A(b[1]), .B(n3302), .Z(n3304) );
  NAND U3495 ( .A(n206), .B(a[48]), .Z(n3303) );
  AND U3496 ( .A(n3304), .B(n3303), .Z(n3367) );
  XOR U3497 ( .A(n3368), .B(n3367), .Z(n3370) );
  NAND U3498 ( .A(a[33]), .B(b[15]), .Z(n3369) );
  XOR U3499 ( .A(n3370), .B(n3369), .Z(n3361) );
  XNOR U3500 ( .A(n3362), .B(n3361), .Z(n3363) );
  NAND U3501 ( .A(n4521), .B(n3305), .Z(n3307) );
  XOR U3502 ( .A(b[3]), .B(a[47]), .Z(n3379) );
  NANDN U3503 ( .A(n4488), .B(n3379), .Z(n3306) );
  NAND U3504 ( .A(n3307), .B(n3306), .Z(n3357) );
  XOR U3505 ( .A(n209), .B(a[45]), .Z(n3382) );
  OR U3506 ( .A(n3382), .B(n4612), .Z(n3310) );
  NANDN U3507 ( .A(n3308), .B(n4669), .Z(n3309) );
  NAND U3508 ( .A(n3310), .B(n3309), .Z(n3355) );
  XNOR U3509 ( .A(n4744), .B(n3865), .Z(n3385) );
  NANDN U3510 ( .A(n3385), .B(n4745), .Z(n3313) );
  NANDN U3511 ( .A(n3311), .B(n4746), .Z(n3312) );
  AND U3512 ( .A(n3313), .B(n3312), .Z(n3356) );
  XOR U3513 ( .A(n3357), .B(n3358), .Z(n3364) );
  XOR U3514 ( .A(n3363), .B(n3364), .Z(n3329) );
  XNOR U3515 ( .A(n3330), .B(n3329), .Z(n3332) );
  XNOR U3516 ( .A(n3331), .B(n3332), .Z(n3391) );
  XOR U3517 ( .A(n3390), .B(n3391), .Z(n3325) );
  NANDN U3518 ( .A(n3315), .B(n3314), .Z(n3319) );
  NANDN U3519 ( .A(n3317), .B(n3316), .Z(n3318) );
  NAND U3520 ( .A(n3319), .B(n3318), .Z(n3326) );
  XOR U3521 ( .A(n3325), .B(n3326), .Z(n3327) );
  XNOR U3522 ( .A(n3328), .B(n3327), .Z(n3394) );
  XNOR U3523 ( .A(n3394), .B(sreg[97]), .Z(n3396) );
  NAND U3524 ( .A(n3320), .B(sreg[96]), .Z(n3324) );
  OR U3525 ( .A(n3322), .B(n3321), .Z(n3323) );
  AND U3526 ( .A(n3324), .B(n3323), .Z(n3395) );
  XOR U3527 ( .A(n3396), .B(n3395), .Z(c[97]) );
  NAND U3528 ( .A(n3330), .B(n3329), .Z(n3334) );
  NANDN U3529 ( .A(n3332), .B(n3331), .Z(n3333) );
  NAND U3530 ( .A(n3334), .B(n3333), .Z(n3463) );
  NANDN U3531 ( .A(n3336), .B(n3335), .Z(n3340) );
  NANDN U3532 ( .A(n3338), .B(n3337), .Z(n3339) );
  NAND U3533 ( .A(n3340), .B(n3339), .Z(n3464) );
  XNOR U3534 ( .A(n3463), .B(n3464), .Z(n3465) );
  XNOR U3535 ( .A(n4859), .B(n3781), .Z(n3405) );
  OR U3536 ( .A(n3405), .B(n4860), .Z(n3343) );
  NANDN U3537 ( .A(n3341), .B(n4915), .Z(n3342) );
  NAND U3538 ( .A(n3343), .B(n3342), .Z(n3417) );
  NANDN U3539 ( .A(n3344), .B(n4987), .Z(n3346) );
  XOR U3540 ( .A(n4909), .B(a[40]), .Z(n3408) );
  OR U3541 ( .A(n3408), .B(n4986), .Z(n3345) );
  NAND U3542 ( .A(n3346), .B(n3345), .Z(n3414) );
  XNOR U3543 ( .A(n210), .B(n3347), .Z(n3411) );
  OR U3544 ( .A(n3411), .B(n5095), .Z(n3350) );
  NANDN U3545 ( .A(n3348), .B(n5092), .Z(n3349) );
  AND U3546 ( .A(n3350), .B(n3349), .Z(n3415) );
  XOR U3547 ( .A(n3414), .B(n3415), .Z(n3416) );
  XOR U3548 ( .A(n3417), .B(n3416), .Z(n3457) );
  XNOR U3549 ( .A(n3457), .B(n3458), .Z(n3459) );
  NANDN U3550 ( .A(n3356), .B(n3355), .Z(n3360) );
  NANDN U3551 ( .A(n3358), .B(n3357), .Z(n3359) );
  NAND U3552 ( .A(n3360), .B(n3359), .Z(n3460) );
  XOR U3553 ( .A(n3459), .B(n3460), .Z(n3454) );
  NAND U3554 ( .A(n3362), .B(n3361), .Z(n3366) );
  OR U3555 ( .A(n3364), .B(n3363), .Z(n3365) );
  NAND U3556 ( .A(n3366), .B(n3365), .Z(n3451) );
  NANDN U3557 ( .A(n3368), .B(n3367), .Z(n3372) );
  OR U3558 ( .A(n3370), .B(n3369), .Z(n3371) );
  NAND U3559 ( .A(n3372), .B(n3371), .Z(n3448) );
  NAND U3560 ( .A(b[0]), .B(a[50]), .Z(n3373) );
  XNOR U3561 ( .A(b[1]), .B(n3373), .Z(n3375) );
  NAND U3562 ( .A(n206), .B(a[49]), .Z(n3374) );
  AND U3563 ( .A(n3375), .B(n3374), .Z(n3424) );
  XNOR U3564 ( .A(n5129), .B(n3496), .Z(n3430) );
  OR U3565 ( .A(n3430), .B(n5041), .Z(n3378) );
  NANDN U3566 ( .A(n3376), .B(n5052), .Z(n3377) );
  AND U3567 ( .A(n3378), .B(n3377), .Z(n3425) );
  XOR U3568 ( .A(n3424), .B(n3425), .Z(n3427) );
  NAND U3569 ( .A(a[34]), .B(b[15]), .Z(n3426) );
  XOR U3570 ( .A(n3427), .B(n3426), .Z(n3445) );
  NAND U3571 ( .A(n4521), .B(n3379), .Z(n3381) );
  XOR U3572 ( .A(b[3]), .B(a[48]), .Z(n3436) );
  NANDN U3573 ( .A(n4488), .B(n3436), .Z(n3380) );
  NAND U3574 ( .A(n3381), .B(n3380), .Z(n3420) );
  XNOR U3575 ( .A(n209), .B(n4089), .Z(n3439) );
  OR U3576 ( .A(n3439), .B(n4612), .Z(n3384) );
  NANDN U3577 ( .A(n3382), .B(n4669), .Z(n3383) );
  NAND U3578 ( .A(n3384), .B(n3383), .Z(n3418) );
  XOR U3579 ( .A(n4744), .B(a[44]), .Z(n3442) );
  NANDN U3580 ( .A(n3442), .B(n4745), .Z(n3387) );
  NANDN U3581 ( .A(n3385), .B(n4746), .Z(n3386) );
  AND U3582 ( .A(n3387), .B(n3386), .Z(n3419) );
  XOR U3583 ( .A(n3420), .B(n3421), .Z(n3446) );
  XNOR U3584 ( .A(n3445), .B(n3446), .Z(n3447) );
  XNOR U3585 ( .A(n3448), .B(n3447), .Z(n3452) );
  XNOR U3586 ( .A(n3451), .B(n3452), .Z(n3453) );
  XNOR U3587 ( .A(n3454), .B(n3453), .Z(n3466) );
  XOR U3588 ( .A(n3465), .B(n3466), .Z(n3399) );
  NANDN U3589 ( .A(n3389), .B(n3388), .Z(n3393) );
  NAND U3590 ( .A(n3391), .B(n3390), .Z(n3392) );
  NAND U3591 ( .A(n3393), .B(n3392), .Z(n3400) );
  XNOR U3592 ( .A(n3399), .B(n3400), .Z(n3401) );
  XNOR U3593 ( .A(n3402), .B(n3401), .Z(n3469) );
  XNOR U3594 ( .A(n3469), .B(sreg[98]), .Z(n3471) );
  NAND U3595 ( .A(n3394), .B(sreg[97]), .Z(n3398) );
  OR U3596 ( .A(n3396), .B(n3395), .Z(n3397) );
  AND U3597 ( .A(n3398), .B(n3397), .Z(n3470) );
  XOR U3598 ( .A(n3471), .B(n3470), .Z(c[98]) );
  NANDN U3599 ( .A(n3400), .B(n3399), .Z(n3404) );
  NAND U3600 ( .A(n3402), .B(n3401), .Z(n3403) );
  NAND U3601 ( .A(n3404), .B(n3403), .Z(n3477) );
  XNOR U3602 ( .A(n4859), .B(n3865), .Z(n3490) );
  OR U3603 ( .A(n3490), .B(n4860), .Z(n3407) );
  NANDN U3604 ( .A(n3405), .B(n4915), .Z(n3406) );
  NAND U3605 ( .A(n3407), .B(n3406), .Z(n3503) );
  NANDN U3606 ( .A(n3408), .B(n4987), .Z(n3410) );
  XNOR U3607 ( .A(n4909), .B(n3736), .Z(n3493) );
  OR U3608 ( .A(n3493), .B(n4986), .Z(n3409) );
  NAND U3609 ( .A(n3410), .B(n3409), .Z(n3500) );
  XOR U3610 ( .A(n210), .B(a[37]), .Z(n3497) );
  OR U3611 ( .A(n3497), .B(n5095), .Z(n3413) );
  NANDN U3612 ( .A(n3411), .B(n5092), .Z(n3412) );
  AND U3613 ( .A(n3413), .B(n3412), .Z(n3501) );
  XOR U3614 ( .A(n3500), .B(n3501), .Z(n3502) );
  XOR U3615 ( .A(n3503), .B(n3502), .Z(n3478) );
  XOR U3616 ( .A(n3478), .B(n3479), .Z(n3481) );
  NANDN U3617 ( .A(n3419), .B(n3418), .Z(n3423) );
  NANDN U3618 ( .A(n3421), .B(n3420), .Z(n3422) );
  AND U3619 ( .A(n3423), .B(n3422), .Z(n3480) );
  XOR U3620 ( .A(n3481), .B(n3480), .Z(n3486) );
  NANDN U3621 ( .A(n3425), .B(n3424), .Z(n3429) );
  OR U3622 ( .A(n3427), .B(n3426), .Z(n3428) );
  NAND U3623 ( .A(n3429), .B(n3428), .Z(n3513) );
  XNOR U3624 ( .A(n5129), .B(n3560), .Z(n3525) );
  OR U3625 ( .A(n3525), .B(n5041), .Z(n3432) );
  NANDN U3626 ( .A(n3430), .B(n5052), .Z(n3431) );
  AND U3627 ( .A(n3432), .B(n3431), .Z(n3517) );
  NAND U3628 ( .A(b[0]), .B(a[51]), .Z(n3433) );
  XNOR U3629 ( .A(b[1]), .B(n3433), .Z(n3435) );
  NAND U3630 ( .A(a[50]), .B(n206), .Z(n3434) );
  AND U3631 ( .A(n3435), .B(n3434), .Z(n3516) );
  XOR U3632 ( .A(n3517), .B(n3516), .Z(n3519) );
  NAND U3633 ( .A(a[35]), .B(b[15]), .Z(n3518) );
  XOR U3634 ( .A(n3519), .B(n3518), .Z(n3510) );
  NAND U3635 ( .A(n4521), .B(n3436), .Z(n3438) );
  XOR U3636 ( .A(b[3]), .B(a[49]), .Z(n3528) );
  NANDN U3637 ( .A(n4488), .B(n3528), .Z(n3437) );
  NAND U3638 ( .A(n3438), .B(n3437), .Z(n3506) );
  XOR U3639 ( .A(n209), .B(a[47]), .Z(n3531) );
  OR U3640 ( .A(n3531), .B(n4612), .Z(n3441) );
  NANDN U3641 ( .A(n3439), .B(n4669), .Z(n3440) );
  NAND U3642 ( .A(n3441), .B(n3440), .Z(n3504) );
  XOR U3643 ( .A(n4744), .B(a[45]), .Z(n3534) );
  NANDN U3644 ( .A(n3534), .B(n4745), .Z(n3444) );
  NANDN U3645 ( .A(n3442), .B(n4746), .Z(n3443) );
  AND U3646 ( .A(n3444), .B(n3443), .Z(n3505) );
  XOR U3647 ( .A(n3506), .B(n3507), .Z(n3511) );
  XNOR U3648 ( .A(n3510), .B(n3511), .Z(n3512) );
  XNOR U3649 ( .A(n3513), .B(n3512), .Z(n3484) );
  NANDN U3650 ( .A(n3446), .B(n3445), .Z(n3450) );
  NAND U3651 ( .A(n3448), .B(n3447), .Z(n3449) );
  NAND U3652 ( .A(n3450), .B(n3449), .Z(n3485) );
  XOR U3653 ( .A(n3484), .B(n3485), .Z(n3487) );
  XNOR U3654 ( .A(n3486), .B(n3487), .Z(n3540) );
  NANDN U3655 ( .A(n3452), .B(n3451), .Z(n3456) );
  NAND U3656 ( .A(n3454), .B(n3453), .Z(n3455) );
  NAND U3657 ( .A(n3456), .B(n3455), .Z(n3537) );
  NANDN U3658 ( .A(n3458), .B(n3457), .Z(n3462) );
  NANDN U3659 ( .A(n3460), .B(n3459), .Z(n3461) );
  NAND U3660 ( .A(n3462), .B(n3461), .Z(n3538) );
  XNOR U3661 ( .A(n3537), .B(n3538), .Z(n3539) );
  XNOR U3662 ( .A(n3540), .B(n3539), .Z(n3474) );
  NANDN U3663 ( .A(n3464), .B(n3463), .Z(n3468) );
  NANDN U3664 ( .A(n3466), .B(n3465), .Z(n3467) );
  NAND U3665 ( .A(n3468), .B(n3467), .Z(n3475) );
  XOR U3666 ( .A(n3474), .B(n3475), .Z(n3476) );
  XOR U3667 ( .A(n3477), .B(n3476), .Z(n3543) );
  XNOR U3668 ( .A(n3543), .B(sreg[99]), .Z(n3545) );
  NAND U3669 ( .A(n3469), .B(sreg[98]), .Z(n3473) );
  OR U3670 ( .A(n3471), .B(n3470), .Z(n3472) );
  AND U3671 ( .A(n3473), .B(n3472), .Z(n3544) );
  XOR U3672 ( .A(n3545), .B(n3544), .Z(c[99]) );
  NANDN U3673 ( .A(n3479), .B(n3478), .Z(n3483) );
  NANDN U3674 ( .A(n3481), .B(n3480), .Z(n3482) );
  NAND U3675 ( .A(n3483), .B(n3482), .Z(n3614) );
  NANDN U3676 ( .A(n3485), .B(n3484), .Z(n3489) );
  OR U3677 ( .A(n3487), .B(n3486), .Z(n3488) );
  AND U3678 ( .A(n3489), .B(n3488), .Z(n3613) );
  XNOR U3679 ( .A(n3614), .B(n3613), .Z(n3615) );
  XOR U3680 ( .A(n4859), .B(a[44]), .Z(n3554) );
  OR U3681 ( .A(n3554), .B(n4860), .Z(n3492) );
  NANDN U3682 ( .A(n3490), .B(n4915), .Z(n3491) );
  NAND U3683 ( .A(n3492), .B(n3491), .Z(n3567) );
  NANDN U3684 ( .A(n3493), .B(n4987), .Z(n3495) );
  XNOR U3685 ( .A(n4909), .B(n3781), .Z(n3557) );
  OR U3686 ( .A(n3557), .B(n4986), .Z(n3494) );
  NAND U3687 ( .A(n3495), .B(n3494), .Z(n3564) );
  XNOR U3688 ( .A(n210), .B(n3496), .Z(n3561) );
  OR U3689 ( .A(n3561), .B(n5095), .Z(n3499) );
  NANDN U3690 ( .A(n3497), .B(n5092), .Z(n3498) );
  AND U3691 ( .A(n3499), .B(n3498), .Z(n3565) );
  XOR U3692 ( .A(n3564), .B(n3565), .Z(n3566) );
  XOR U3693 ( .A(n3567), .B(n3566), .Z(n3607) );
  XNOR U3694 ( .A(n3607), .B(n3608), .Z(n3609) );
  NANDN U3695 ( .A(n3505), .B(n3504), .Z(n3509) );
  NANDN U3696 ( .A(n3507), .B(n3506), .Z(n3508) );
  NAND U3697 ( .A(n3509), .B(n3508), .Z(n3610) );
  XOR U3698 ( .A(n3609), .B(n3610), .Z(n3604) );
  NANDN U3699 ( .A(n3511), .B(n3510), .Z(n3515) );
  NAND U3700 ( .A(n3513), .B(n3512), .Z(n3514) );
  NAND U3701 ( .A(n3515), .B(n3514), .Z(n3601) );
  NANDN U3702 ( .A(n3517), .B(n3516), .Z(n3521) );
  OR U3703 ( .A(n3519), .B(n3518), .Z(n3520) );
  NAND U3704 ( .A(n3521), .B(n3520), .Z(n3598) );
  NAND U3705 ( .A(b[0]), .B(a[52]), .Z(n3522) );
  XNOR U3706 ( .A(b[1]), .B(n3522), .Z(n3524) );
  NAND U3707 ( .A(n206), .B(a[51]), .Z(n3523) );
  AND U3708 ( .A(n3524), .B(n3523), .Z(n3589) );
  XOR U3709 ( .A(n5129), .B(a[40]), .Z(n3574) );
  OR U3710 ( .A(n3574), .B(n5041), .Z(n3527) );
  NANDN U3711 ( .A(n3525), .B(n5052), .Z(n3526) );
  AND U3712 ( .A(n3527), .B(n3526), .Z(n3590) );
  XOR U3713 ( .A(n3589), .B(n3590), .Z(n3592) );
  NAND U3714 ( .A(a[36]), .B(b[15]), .Z(n3591) );
  XOR U3715 ( .A(n3592), .B(n3591), .Z(n3595) );
  NAND U3716 ( .A(n4521), .B(n3528), .Z(n3530) );
  IV U3717 ( .A(a[50]), .Z(n4394) );
  XNOR U3718 ( .A(b[3]), .B(n4394), .Z(n3580) );
  NANDN U3719 ( .A(n4488), .B(n3580), .Z(n3529) );
  NAND U3720 ( .A(n3530), .B(n3529), .Z(n3570) );
  XOR U3721 ( .A(n209), .B(a[48]), .Z(n3583) );
  OR U3722 ( .A(n3583), .B(n4612), .Z(n3533) );
  NANDN U3723 ( .A(n3531), .B(n4669), .Z(n3532) );
  NAND U3724 ( .A(n3533), .B(n3532), .Z(n3568) );
  XNOR U3725 ( .A(n4744), .B(n4089), .Z(n3586) );
  NANDN U3726 ( .A(n3586), .B(n4745), .Z(n3536) );
  NANDN U3727 ( .A(n3534), .B(n4746), .Z(n3535) );
  AND U3728 ( .A(n3536), .B(n3535), .Z(n3569) );
  XOR U3729 ( .A(n3570), .B(n3571), .Z(n3596) );
  XNOR U3730 ( .A(n3595), .B(n3596), .Z(n3597) );
  XNOR U3731 ( .A(n3598), .B(n3597), .Z(n3602) );
  XNOR U3732 ( .A(n3601), .B(n3602), .Z(n3603) );
  XNOR U3733 ( .A(n3604), .B(n3603), .Z(n3616) );
  XOR U3734 ( .A(n3615), .B(n3616), .Z(n3548) );
  NANDN U3735 ( .A(n3538), .B(n3537), .Z(n3542) );
  NAND U3736 ( .A(n3540), .B(n3539), .Z(n3541) );
  NAND U3737 ( .A(n3542), .B(n3541), .Z(n3549) );
  XNOR U3738 ( .A(n3548), .B(n3549), .Z(n3550) );
  XNOR U3739 ( .A(n3551), .B(n3550), .Z(n3619) );
  XNOR U3740 ( .A(n3619), .B(sreg[100]), .Z(n3621) );
  NAND U3741 ( .A(n3543), .B(sreg[99]), .Z(n3547) );
  OR U3742 ( .A(n3545), .B(n3544), .Z(n3546) );
  AND U3743 ( .A(n3547), .B(n3546), .Z(n3620) );
  XOR U3744 ( .A(n3621), .B(n3620), .Z(c[100]) );
  NANDN U3745 ( .A(n3549), .B(n3548), .Z(n3553) );
  NAND U3746 ( .A(n3551), .B(n3550), .Z(n3552) );
  NAND U3747 ( .A(n3553), .B(n3552), .Z(n3627) );
  XOR U3748 ( .A(n4859), .B(a[45]), .Z(n3640) );
  OR U3749 ( .A(n3640), .B(n4860), .Z(n3556) );
  NANDN U3750 ( .A(n3554), .B(n4915), .Z(n3555) );
  NAND U3751 ( .A(n3556), .B(n3555), .Z(n3652) );
  NANDN U3752 ( .A(n3557), .B(n4987), .Z(n3559) );
  XNOR U3753 ( .A(n4909), .B(n3865), .Z(n3643) );
  OR U3754 ( .A(n3643), .B(n4986), .Z(n3558) );
  NAND U3755 ( .A(n3559), .B(n3558), .Z(n3649) );
  XNOR U3756 ( .A(n210), .B(n3560), .Z(n3646) );
  OR U3757 ( .A(n3646), .B(n5095), .Z(n3563) );
  NANDN U3758 ( .A(n3561), .B(n5092), .Z(n3562) );
  AND U3759 ( .A(n3563), .B(n3562), .Z(n3650) );
  XOR U3760 ( .A(n3649), .B(n3650), .Z(n3651) );
  XOR U3761 ( .A(n3652), .B(n3651), .Z(n3628) );
  XOR U3762 ( .A(n3628), .B(n3629), .Z(n3631) );
  NANDN U3763 ( .A(n3569), .B(n3568), .Z(n3573) );
  NANDN U3764 ( .A(n3571), .B(n3570), .Z(n3572) );
  AND U3765 ( .A(n3573), .B(n3572), .Z(n3630) );
  XOR U3766 ( .A(n3631), .B(n3630), .Z(n3637) );
  XNOR U3767 ( .A(n5129), .B(n3736), .Z(n3674) );
  OR U3768 ( .A(n3674), .B(n5041), .Z(n3576) );
  NANDN U3769 ( .A(n3574), .B(n5052), .Z(n3575) );
  AND U3770 ( .A(n3576), .B(n3575), .Z(n3666) );
  NAND U3771 ( .A(b[0]), .B(a[53]), .Z(n3577) );
  XNOR U3772 ( .A(b[1]), .B(n3577), .Z(n3579) );
  NAND U3773 ( .A(a[52]), .B(n206), .Z(n3578) );
  AND U3774 ( .A(n3579), .B(n3578), .Z(n3665) );
  XOR U3775 ( .A(n3666), .B(n3665), .Z(n3668) );
  NAND U3776 ( .A(b[15]), .B(a[37]), .Z(n3667) );
  XNOR U3777 ( .A(n3668), .B(n3667), .Z(n3659) );
  NAND U3778 ( .A(n4521), .B(n3580), .Z(n3582) );
  XOR U3779 ( .A(n208), .B(a[51]), .Z(n3677) );
  OR U3780 ( .A(n3677), .B(n4488), .Z(n3581) );
  NAND U3781 ( .A(n3582), .B(n3581), .Z(n3656) );
  XOR U3782 ( .A(b[5]), .B(a[49]), .Z(n3680) );
  NANDN U3783 ( .A(n4612), .B(n3680), .Z(n3585) );
  NANDN U3784 ( .A(n3583), .B(n4669), .Z(n3584) );
  NAND U3785 ( .A(n3585), .B(n3584), .Z(n3653) );
  XOR U3786 ( .A(n4744), .B(a[47]), .Z(n3683) );
  NANDN U3787 ( .A(n3683), .B(n4745), .Z(n3588) );
  NANDN U3788 ( .A(n3586), .B(n4746), .Z(n3587) );
  AND U3789 ( .A(n3588), .B(n3587), .Z(n3654) );
  XOR U3790 ( .A(n3656), .B(n3655), .Z(n3660) );
  XNOR U3791 ( .A(n3659), .B(n3660), .Z(n3661) );
  NANDN U3792 ( .A(n3590), .B(n3589), .Z(n3594) );
  OR U3793 ( .A(n3592), .B(n3591), .Z(n3593) );
  AND U3794 ( .A(n3594), .B(n3593), .Z(n3662) );
  XNOR U3795 ( .A(n3661), .B(n3662), .Z(n3635) );
  NANDN U3796 ( .A(n3596), .B(n3595), .Z(n3600) );
  NAND U3797 ( .A(n3598), .B(n3597), .Z(n3599) );
  AND U3798 ( .A(n3600), .B(n3599), .Z(n3634) );
  XNOR U3799 ( .A(n3635), .B(n3634), .Z(n3636) );
  XOR U3800 ( .A(n3637), .B(n3636), .Z(n3689) );
  NANDN U3801 ( .A(n3602), .B(n3601), .Z(n3606) );
  NAND U3802 ( .A(n3604), .B(n3603), .Z(n3605) );
  NAND U3803 ( .A(n3606), .B(n3605), .Z(n3686) );
  NANDN U3804 ( .A(n3608), .B(n3607), .Z(n3612) );
  NANDN U3805 ( .A(n3610), .B(n3609), .Z(n3611) );
  NAND U3806 ( .A(n3612), .B(n3611), .Z(n3687) );
  XNOR U3807 ( .A(n3686), .B(n3687), .Z(n3688) );
  XNOR U3808 ( .A(n3689), .B(n3688), .Z(n3624) );
  NANDN U3809 ( .A(n3614), .B(n3613), .Z(n3618) );
  NANDN U3810 ( .A(n3616), .B(n3615), .Z(n3617) );
  NAND U3811 ( .A(n3618), .B(n3617), .Z(n3625) );
  XOR U3812 ( .A(n3624), .B(n3625), .Z(n3626) );
  XOR U3813 ( .A(n3627), .B(n3626), .Z(n3692) );
  XNOR U3814 ( .A(n3692), .B(sreg[101]), .Z(n3694) );
  NAND U3815 ( .A(n3619), .B(sreg[100]), .Z(n3623) );
  OR U3816 ( .A(n3621), .B(n3620), .Z(n3622) );
  AND U3817 ( .A(n3623), .B(n3622), .Z(n3693) );
  XOR U3818 ( .A(n3694), .B(n3693), .Z(c[101]) );
  NANDN U3819 ( .A(n3629), .B(n3628), .Z(n3633) );
  NANDN U3820 ( .A(n3631), .B(n3630), .Z(n3632) );
  NAND U3821 ( .A(n3633), .B(n3632), .Z(n3761) );
  NANDN U3822 ( .A(n3635), .B(n3634), .Z(n3639) );
  NANDN U3823 ( .A(n3637), .B(n3636), .Z(n3638) );
  AND U3824 ( .A(n3639), .B(n3638), .Z(n3760) );
  XNOR U3825 ( .A(n3761), .B(n3760), .Z(n3762) );
  XNOR U3826 ( .A(n4859), .B(n4089), .Z(n3730) );
  OR U3827 ( .A(n3730), .B(n4860), .Z(n3642) );
  NANDN U3828 ( .A(n3640), .B(n4915), .Z(n3641) );
  NAND U3829 ( .A(n3642), .B(n3641), .Z(n3743) );
  NANDN U3830 ( .A(n3643), .B(n4987), .Z(n3645) );
  XOR U3831 ( .A(n4909), .B(a[44]), .Z(n3733) );
  OR U3832 ( .A(n3733), .B(n4986), .Z(n3644) );
  NAND U3833 ( .A(n3645), .B(n3644), .Z(n3740) );
  XOR U3834 ( .A(n210), .B(a[40]), .Z(n3737) );
  OR U3835 ( .A(n3737), .B(n5095), .Z(n3648) );
  NANDN U3836 ( .A(n3646), .B(n5092), .Z(n3647) );
  AND U3837 ( .A(n3648), .B(n3647), .Z(n3741) );
  XOR U3838 ( .A(n3740), .B(n3741), .Z(n3742) );
  XOR U3839 ( .A(n3743), .B(n3742), .Z(n3754) );
  XNOR U3840 ( .A(n3754), .B(n3755), .Z(n3756) );
  NANDN U3841 ( .A(n3654), .B(n3653), .Z(n3658) );
  NAND U3842 ( .A(n3656), .B(n3655), .Z(n3657) );
  NAND U3843 ( .A(n3658), .B(n3657), .Z(n3757) );
  XOR U3844 ( .A(n3756), .B(n3757), .Z(n3751) );
  NANDN U3845 ( .A(n3660), .B(n3659), .Z(n3664) );
  NAND U3846 ( .A(n3662), .B(n3661), .Z(n3663) );
  NAND U3847 ( .A(n3664), .B(n3663), .Z(n3749) );
  NANDN U3848 ( .A(n3666), .B(n3665), .Z(n3670) );
  OR U3849 ( .A(n3668), .B(n3667), .Z(n3669) );
  NAND U3850 ( .A(n3670), .B(n3669), .Z(n3727) );
  NAND U3851 ( .A(b[0]), .B(a[54]), .Z(n3671) );
  XNOR U3852 ( .A(b[1]), .B(n3671), .Z(n3673) );
  NAND U3853 ( .A(n206), .B(a[53]), .Z(n3672) );
  AND U3854 ( .A(n3673), .B(n3672), .Z(n3703) );
  XNOR U3855 ( .A(n5129), .B(n3781), .Z(n3712) );
  OR U3856 ( .A(n3712), .B(n5041), .Z(n3676) );
  NANDN U3857 ( .A(n3674), .B(n5052), .Z(n3675) );
  AND U3858 ( .A(n3676), .B(n3675), .Z(n3704) );
  XOR U3859 ( .A(n3703), .B(n3704), .Z(n3706) );
  NAND U3860 ( .A(a[38]), .B(b[15]), .Z(n3705) );
  XOR U3861 ( .A(n3706), .B(n3705), .Z(n3724) );
  NANDN U3862 ( .A(n3677), .B(n4521), .Z(n3679) );
  XOR U3863 ( .A(a[52]), .B(b[3]), .Z(n3715) );
  NANDN U3864 ( .A(n4488), .B(n3715), .Z(n3678) );
  AND U3865 ( .A(n3679), .B(n3678), .Z(n3746) );
  NAND U3866 ( .A(n4669), .B(n3680), .Z(n3682) );
  XOR U3867 ( .A(b[5]), .B(a[50]), .Z(n3718) );
  NANDN U3868 ( .A(n4612), .B(n3718), .Z(n3681) );
  AND U3869 ( .A(n3682), .B(n3681), .Z(n3744) );
  XOR U3870 ( .A(n4744), .B(a[48]), .Z(n3721) );
  NANDN U3871 ( .A(n3721), .B(n4745), .Z(n3685) );
  NANDN U3872 ( .A(n3683), .B(n4746), .Z(n3684) );
  AND U3873 ( .A(n3685), .B(n3684), .Z(n3745) );
  XOR U3874 ( .A(n3744), .B(n3745), .Z(n3747) );
  XOR U3875 ( .A(n3746), .B(n3747), .Z(n3725) );
  XNOR U3876 ( .A(n3724), .B(n3725), .Z(n3726) );
  XOR U3877 ( .A(n3727), .B(n3726), .Z(n3748) );
  XNOR U3878 ( .A(n3749), .B(n3748), .Z(n3750) );
  XNOR U3879 ( .A(n3751), .B(n3750), .Z(n3763) );
  XOR U3880 ( .A(n3762), .B(n3763), .Z(n3697) );
  NANDN U3881 ( .A(n3687), .B(n3686), .Z(n3691) );
  NAND U3882 ( .A(n3689), .B(n3688), .Z(n3690) );
  NAND U3883 ( .A(n3691), .B(n3690), .Z(n3698) );
  XNOR U3884 ( .A(n3697), .B(n3698), .Z(n3699) );
  XNOR U3885 ( .A(n3700), .B(n3699), .Z(n3766) );
  XNOR U3886 ( .A(n3766), .B(sreg[102]), .Z(n3768) );
  NAND U3887 ( .A(n3692), .B(sreg[101]), .Z(n3696) );
  OR U3888 ( .A(n3694), .B(n3693), .Z(n3695) );
  AND U3889 ( .A(n3696), .B(n3695), .Z(n3767) );
  XOR U3890 ( .A(n3768), .B(n3767), .Z(c[102]) );
  NANDN U3891 ( .A(n3698), .B(n3697), .Z(n3702) );
  NAND U3892 ( .A(n3700), .B(n3699), .Z(n3701) );
  NAND U3893 ( .A(n3702), .B(n3701), .Z(n3774) );
  NANDN U3894 ( .A(n3704), .B(n3703), .Z(n3708) );
  OR U3895 ( .A(n3706), .B(n3705), .Z(n3707) );
  NAND U3896 ( .A(n3708), .B(n3707), .Z(n3821) );
  NAND U3897 ( .A(b[0]), .B(a[55]), .Z(n3709) );
  XNOR U3898 ( .A(b[1]), .B(n3709), .Z(n3711) );
  NAND U3899 ( .A(a[54]), .B(n206), .Z(n3710) );
  AND U3900 ( .A(n3711), .B(n3710), .Z(n3812) );
  XNOR U3901 ( .A(n5129), .B(n3865), .Z(n3800) );
  OR U3902 ( .A(n3800), .B(n5041), .Z(n3714) );
  NANDN U3903 ( .A(n3712), .B(n5052), .Z(n3713) );
  AND U3904 ( .A(n3714), .B(n3713), .Z(n3813) );
  XOR U3905 ( .A(n3812), .B(n3813), .Z(n3815) );
  NAND U3906 ( .A(a[39]), .B(b[15]), .Z(n3814) );
  XOR U3907 ( .A(n3815), .B(n3814), .Z(n3818) );
  NAND U3908 ( .A(n3715), .B(n4521), .Z(n3717) );
  XOR U3909 ( .A(b[3]), .B(a[53]), .Z(n3803) );
  NANDN U3910 ( .A(n4488), .B(n3803), .Z(n3716) );
  NAND U3911 ( .A(n3717), .B(n3716), .Z(n3793) );
  XOR U3912 ( .A(n209), .B(a[51]), .Z(n3806) );
  OR U3913 ( .A(n3806), .B(n4612), .Z(n3720) );
  NAND U3914 ( .A(n3718), .B(n4669), .Z(n3719) );
  NAND U3915 ( .A(n3720), .B(n3719), .Z(n3791) );
  XOR U3916 ( .A(n4744), .B(a[49]), .Z(n3809) );
  NANDN U3917 ( .A(n3809), .B(n4745), .Z(n3723) );
  NANDN U3918 ( .A(n3721), .B(n4746), .Z(n3722) );
  AND U3919 ( .A(n3723), .B(n3722), .Z(n3792) );
  XOR U3920 ( .A(n3793), .B(n3794), .Z(n3819) );
  XNOR U3921 ( .A(n3818), .B(n3819), .Z(n3820) );
  XNOR U3922 ( .A(n3821), .B(n3820), .Z(n3824) );
  NANDN U3923 ( .A(n3725), .B(n3724), .Z(n3729) );
  NAND U3924 ( .A(n3727), .B(n3726), .Z(n3728) );
  NAND U3925 ( .A(n3729), .B(n3728), .Z(n3825) );
  XOR U3926 ( .A(n3824), .B(n3825), .Z(n3826) );
  XOR U3927 ( .A(n4859), .B(a[47]), .Z(n3775) );
  OR U3928 ( .A(n3775), .B(n4860), .Z(n3732) );
  NANDN U3929 ( .A(n3730), .B(n4915), .Z(n3731) );
  NAND U3930 ( .A(n3732), .B(n3731), .Z(n3788) );
  NANDN U3931 ( .A(n3733), .B(n4987), .Z(n3735) );
  XOR U3932 ( .A(n4909), .B(a[45]), .Z(n3778) );
  OR U3933 ( .A(n3778), .B(n4986), .Z(n3734) );
  NAND U3934 ( .A(n3735), .B(n3734), .Z(n3785) );
  XNOR U3935 ( .A(n210), .B(n3736), .Z(n3782) );
  OR U3936 ( .A(n3782), .B(n5095), .Z(n3739) );
  NANDN U3937 ( .A(n3737), .B(n5092), .Z(n3738) );
  AND U3938 ( .A(n3739), .B(n3738), .Z(n3786) );
  XNOR U3939 ( .A(n3785), .B(n3786), .Z(n3787) );
  XOR U3940 ( .A(n3788), .B(n3787), .Z(n3828) );
  XNOR U3941 ( .A(n3828), .B(n3829), .Z(n3831) );
  XOR U3942 ( .A(n3831), .B(n3830), .Z(n3827) );
  XNOR U3943 ( .A(n3826), .B(n3827), .Z(n3835) );
  NANDN U3944 ( .A(n3749), .B(n3748), .Z(n3753) );
  NAND U3945 ( .A(n3751), .B(n3750), .Z(n3752) );
  NAND U3946 ( .A(n3753), .B(n3752), .Z(n3832) );
  NANDN U3947 ( .A(n3755), .B(n3754), .Z(n3759) );
  NANDN U3948 ( .A(n3757), .B(n3756), .Z(n3758) );
  NAND U3949 ( .A(n3759), .B(n3758), .Z(n3833) );
  XNOR U3950 ( .A(n3832), .B(n3833), .Z(n3834) );
  XOR U3951 ( .A(n3835), .B(n3834), .Z(n3771) );
  NANDN U3952 ( .A(n3761), .B(n3760), .Z(n3765) );
  NANDN U3953 ( .A(n3763), .B(n3762), .Z(n3764) );
  NAND U3954 ( .A(n3765), .B(n3764), .Z(n3772) );
  XOR U3955 ( .A(n3771), .B(n3772), .Z(n3773) );
  XOR U3956 ( .A(n3774), .B(n3773), .Z(n3838) );
  XNOR U3957 ( .A(n3838), .B(sreg[103]), .Z(n3840) );
  NAND U3958 ( .A(n3766), .B(sreg[102]), .Z(n3770) );
  OR U3959 ( .A(n3768), .B(n3767), .Z(n3769) );
  AND U3960 ( .A(n3770), .B(n3769), .Z(n3839) );
  XOR U3961 ( .A(n3840), .B(n3839), .Z(c[103]) );
  XOR U3962 ( .A(n4859), .B(a[48]), .Z(n3859) );
  OR U3963 ( .A(n3859), .B(n4860), .Z(n3777) );
  NANDN U3964 ( .A(n3775), .B(n4915), .Z(n3776) );
  NAND U3965 ( .A(n3777), .B(n3776), .Z(n3872) );
  NANDN U3966 ( .A(n3778), .B(n4987), .Z(n3780) );
  XNOR U3967 ( .A(n4909), .B(n4089), .Z(n3862) );
  OR U3968 ( .A(n3862), .B(n4986), .Z(n3779) );
  NAND U3969 ( .A(n3780), .B(n3779), .Z(n3869) );
  XNOR U3970 ( .A(n210), .B(n3781), .Z(n3866) );
  OR U3971 ( .A(n3866), .B(n5095), .Z(n3784) );
  NANDN U3972 ( .A(n3782), .B(n5092), .Z(n3783) );
  AND U3973 ( .A(n3784), .B(n3783), .Z(n3870) );
  XOR U3974 ( .A(n3869), .B(n3870), .Z(n3871) );
  XOR U3975 ( .A(n3872), .B(n3871), .Z(n3847) );
  NANDN U3976 ( .A(n3786), .B(n3785), .Z(n3790) );
  NAND U3977 ( .A(n3788), .B(n3787), .Z(n3789) );
  NAND U3978 ( .A(n3790), .B(n3789), .Z(n3848) );
  XOR U3979 ( .A(n3847), .B(n3848), .Z(n3850) );
  NANDN U3980 ( .A(n3792), .B(n3791), .Z(n3796) );
  NANDN U3981 ( .A(n3794), .B(n3793), .Z(n3795) );
  AND U3982 ( .A(n3796), .B(n3795), .Z(n3849) );
  XOR U3983 ( .A(n3850), .B(n3849), .Z(n3856) );
  NAND U3984 ( .A(b[0]), .B(a[56]), .Z(n3797) );
  XNOR U3985 ( .A(b[1]), .B(n3797), .Z(n3799) );
  NAND U3986 ( .A(a[55]), .B(n206), .Z(n3798) );
  AND U3987 ( .A(n3799), .B(n3798), .Z(n3885) );
  XOR U3988 ( .A(n5129), .B(a[44]), .Z(n3894) );
  OR U3989 ( .A(n3894), .B(n5041), .Z(n3802) );
  NANDN U3990 ( .A(n3800), .B(n5052), .Z(n3801) );
  AND U3991 ( .A(n3802), .B(n3801), .Z(n3886) );
  XOR U3992 ( .A(n3885), .B(n3886), .Z(n3888) );
  NAND U3993 ( .A(b[15]), .B(a[40]), .Z(n3887) );
  XNOR U3994 ( .A(n3888), .B(n3887), .Z(n3879) );
  NAND U3995 ( .A(n4521), .B(n3803), .Z(n3805) );
  XNOR U3996 ( .A(a[54]), .B(n208), .Z(n3897) );
  NANDN U3997 ( .A(n4488), .B(n3897), .Z(n3804) );
  NAND U3998 ( .A(n3805), .B(n3804), .Z(n3876) );
  IV U3999 ( .A(a[52]), .Z(n4528) );
  XNOR U4000 ( .A(n209), .B(n4528), .Z(n3900) );
  OR U4001 ( .A(n3900), .B(n4612), .Z(n3808) );
  NANDN U4002 ( .A(n3806), .B(n4669), .Z(n3807) );
  NAND U4003 ( .A(n3808), .B(n3807), .Z(n3873) );
  XNOR U4004 ( .A(n4744), .B(n4394), .Z(n3903) );
  NANDN U4005 ( .A(n3903), .B(n4745), .Z(n3811) );
  NANDN U4006 ( .A(n3809), .B(n4746), .Z(n3810) );
  AND U4007 ( .A(n3811), .B(n3810), .Z(n3874) );
  XOR U4008 ( .A(n3876), .B(n3875), .Z(n3880) );
  XNOR U4009 ( .A(n3879), .B(n3880), .Z(n3881) );
  NANDN U4010 ( .A(n3813), .B(n3812), .Z(n3817) );
  OR U4011 ( .A(n3815), .B(n3814), .Z(n3816) );
  AND U4012 ( .A(n3817), .B(n3816), .Z(n3882) );
  XNOR U4013 ( .A(n3881), .B(n3882), .Z(n3854) );
  NANDN U4014 ( .A(n3819), .B(n3818), .Z(n3823) );
  NAND U4015 ( .A(n3821), .B(n3820), .Z(n3822) );
  AND U4016 ( .A(n3823), .B(n3822), .Z(n3853) );
  XNOR U4017 ( .A(n3854), .B(n3853), .Z(n3855) );
  XOR U4018 ( .A(n3856), .B(n3855), .Z(n3909) );
  XNOR U4019 ( .A(n3907), .B(n3906), .Z(n3908) );
  XNOR U4020 ( .A(n3909), .B(n3908), .Z(n3843) );
  NANDN U4021 ( .A(n3833), .B(n3832), .Z(n3837) );
  NANDN U4022 ( .A(n3835), .B(n3834), .Z(n3836) );
  NAND U4023 ( .A(n3837), .B(n3836), .Z(n3844) );
  XOR U4024 ( .A(n3843), .B(n3844), .Z(n3845) );
  XOR U4025 ( .A(n3846), .B(n3845), .Z(n3912) );
  XNOR U4026 ( .A(n3912), .B(sreg[104]), .Z(n3914) );
  NAND U4027 ( .A(n3838), .B(sreg[103]), .Z(n3842) );
  OR U4028 ( .A(n3840), .B(n3839), .Z(n3841) );
  AND U4029 ( .A(n3842), .B(n3841), .Z(n3913) );
  XOR U4030 ( .A(n3914), .B(n3913), .Z(c[104]) );
  NANDN U4031 ( .A(n3848), .B(n3847), .Z(n3852) );
  NANDN U4032 ( .A(n3850), .B(n3849), .Z(n3851) );
  NAND U4033 ( .A(n3852), .B(n3851), .Z(n3982) );
  NANDN U4034 ( .A(n3854), .B(n3853), .Z(n3858) );
  NANDN U4035 ( .A(n3856), .B(n3855), .Z(n3857) );
  AND U4036 ( .A(n3858), .B(n3857), .Z(n3981) );
  XNOR U4037 ( .A(n3982), .B(n3981), .Z(n3983) );
  XOR U4038 ( .A(n4859), .B(a[49]), .Z(n3923) );
  OR U4039 ( .A(n3923), .B(n4860), .Z(n3861) );
  NANDN U4040 ( .A(n3859), .B(n4915), .Z(n3860) );
  NAND U4041 ( .A(n3861), .B(n3860), .Z(n3935) );
  NANDN U4042 ( .A(n3862), .B(n4987), .Z(n3864) );
  XOR U4043 ( .A(n4909), .B(a[47]), .Z(n3926) );
  OR U4044 ( .A(n3926), .B(n4986), .Z(n3863) );
  NAND U4045 ( .A(n3864), .B(n3863), .Z(n3932) );
  XNOR U4046 ( .A(n210), .B(n3865), .Z(n3929) );
  OR U4047 ( .A(n3929), .B(n5095), .Z(n3868) );
  NANDN U4048 ( .A(n3866), .B(n5092), .Z(n3867) );
  AND U4049 ( .A(n3868), .B(n3867), .Z(n3933) );
  XOR U4050 ( .A(n3932), .B(n3933), .Z(n3934) );
  XOR U4051 ( .A(n3935), .B(n3934), .Z(n3975) );
  XNOR U4052 ( .A(n3975), .B(n3976), .Z(n3977) );
  NANDN U4053 ( .A(n3874), .B(n3873), .Z(n3878) );
  NAND U4054 ( .A(n3876), .B(n3875), .Z(n3877) );
  NAND U4055 ( .A(n3878), .B(n3877), .Z(n3978) );
  XOR U4056 ( .A(n3977), .B(n3978), .Z(n3972) );
  NANDN U4057 ( .A(n3880), .B(n3879), .Z(n3884) );
  NAND U4058 ( .A(n3882), .B(n3881), .Z(n3883) );
  NAND U4059 ( .A(n3884), .B(n3883), .Z(n3970) );
  NANDN U4060 ( .A(n3886), .B(n3885), .Z(n3890) );
  OR U4061 ( .A(n3888), .B(n3887), .Z(n3889) );
  NAND U4062 ( .A(n3890), .B(n3889), .Z(n3945) );
  NAND U4063 ( .A(b[0]), .B(a[57]), .Z(n3891) );
  XNOR U4064 ( .A(b[1]), .B(n3891), .Z(n3893) );
  NAND U4065 ( .A(a[56]), .B(n206), .Z(n3892) );
  AND U4066 ( .A(n3893), .B(n3892), .Z(n3948) );
  XOR U4067 ( .A(n5129), .B(a[45]), .Z(n3957) );
  OR U4068 ( .A(n3957), .B(n5041), .Z(n3896) );
  NANDN U4069 ( .A(n3894), .B(n5052), .Z(n3895) );
  AND U4070 ( .A(n3896), .B(n3895), .Z(n3949) );
  XOR U4071 ( .A(n3948), .B(n3949), .Z(n3951) );
  NAND U4072 ( .A(a[41]), .B(b[15]), .Z(n3950) );
  XOR U4073 ( .A(n3951), .B(n3950), .Z(n3942) );
  NAND U4074 ( .A(n4521), .B(n3897), .Z(n3899) );
  XNOR U4075 ( .A(a[55]), .B(n208), .Z(n3960) );
  NANDN U4076 ( .A(n4488), .B(n3960), .Z(n3898) );
  NAND U4077 ( .A(n3899), .B(n3898), .Z(n3938) );
  XOR U4078 ( .A(n209), .B(a[53]), .Z(n3963) );
  OR U4079 ( .A(n3963), .B(n4612), .Z(n3902) );
  NANDN U4080 ( .A(n3900), .B(n4669), .Z(n3901) );
  NAND U4081 ( .A(n3902), .B(n3901), .Z(n3936) );
  XOR U4082 ( .A(n4744), .B(a[51]), .Z(n3966) );
  NANDN U4083 ( .A(n3966), .B(n4745), .Z(n3905) );
  NANDN U4084 ( .A(n3903), .B(n4746), .Z(n3904) );
  AND U4085 ( .A(n3905), .B(n3904), .Z(n3937) );
  XOR U4086 ( .A(n3938), .B(n3939), .Z(n3943) );
  XNOR U4087 ( .A(n3942), .B(n3943), .Z(n3944) );
  XOR U4088 ( .A(n3945), .B(n3944), .Z(n3969) );
  XNOR U4089 ( .A(n3970), .B(n3969), .Z(n3971) );
  XNOR U4090 ( .A(n3972), .B(n3971), .Z(n3984) );
  XOR U4091 ( .A(n3983), .B(n3984), .Z(n3917) );
  NANDN U4092 ( .A(n3907), .B(n3906), .Z(n3911) );
  NAND U4093 ( .A(n3909), .B(n3908), .Z(n3910) );
  NAND U4094 ( .A(n3911), .B(n3910), .Z(n3918) );
  XNOR U4095 ( .A(n3917), .B(n3918), .Z(n3919) );
  XNOR U4096 ( .A(n3920), .B(n3919), .Z(n3987) );
  XNOR U4097 ( .A(n3987), .B(sreg[105]), .Z(n3989) );
  NAND U4098 ( .A(n3912), .B(sreg[104]), .Z(n3916) );
  OR U4099 ( .A(n3914), .B(n3913), .Z(n3915) );
  AND U4100 ( .A(n3916), .B(n3915), .Z(n3988) );
  XOR U4101 ( .A(n3989), .B(n3988), .Z(c[105]) );
  NANDN U4102 ( .A(n3918), .B(n3917), .Z(n3922) );
  NAND U4103 ( .A(n3920), .B(n3919), .Z(n3921) );
  NAND U4104 ( .A(n3922), .B(n3921), .Z(n3995) );
  XNOR U4105 ( .A(n4859), .B(n4394), .Z(n4008) );
  OR U4106 ( .A(n4008), .B(n4860), .Z(n3925) );
  NANDN U4107 ( .A(n3923), .B(n4915), .Z(n3924) );
  NAND U4108 ( .A(n3925), .B(n3924), .Z(n4020) );
  NANDN U4109 ( .A(n3926), .B(n4987), .Z(n3928) );
  XOR U4110 ( .A(n4909), .B(a[48]), .Z(n4011) );
  OR U4111 ( .A(n4011), .B(n4986), .Z(n3927) );
  NAND U4112 ( .A(n3928), .B(n3927), .Z(n4017) );
  XOR U4113 ( .A(n210), .B(a[44]), .Z(n4014) );
  OR U4114 ( .A(n4014), .B(n5095), .Z(n3931) );
  NANDN U4115 ( .A(n3929), .B(n5092), .Z(n3930) );
  AND U4116 ( .A(n3931), .B(n3930), .Z(n4018) );
  XOR U4117 ( .A(n4017), .B(n4018), .Z(n4019) );
  XOR U4118 ( .A(n4020), .B(n4019), .Z(n4002) );
  XNOR U4119 ( .A(n4002), .B(n4003), .Z(n4004) );
  NANDN U4120 ( .A(n3937), .B(n3936), .Z(n3941) );
  NANDN U4121 ( .A(n3939), .B(n3938), .Z(n3940) );
  NAND U4122 ( .A(n3941), .B(n3940), .Z(n4005) );
  XOR U4123 ( .A(n4004), .B(n4005), .Z(n3998) );
  NANDN U4124 ( .A(n3943), .B(n3942), .Z(n3947) );
  NAND U4125 ( .A(n3945), .B(n3944), .Z(n3946) );
  NAND U4126 ( .A(n3947), .B(n3946), .Z(n3997) );
  NANDN U4127 ( .A(n3949), .B(n3948), .Z(n3953) );
  OR U4128 ( .A(n3951), .B(n3950), .Z(n3952) );
  NAND U4129 ( .A(n3953), .B(n3952), .Z(n4028) );
  NAND U4130 ( .A(b[0]), .B(a[58]), .Z(n3954) );
  XNOR U4131 ( .A(b[1]), .B(n3954), .Z(n3956) );
  NAND U4132 ( .A(a[57]), .B(n206), .Z(n3955) );
  AND U4133 ( .A(n3956), .B(n3955), .Z(n4033) );
  XNOR U4134 ( .A(n5129), .B(n4089), .Z(n4039) );
  OR U4135 ( .A(n4039), .B(n5041), .Z(n3959) );
  NANDN U4136 ( .A(n3957), .B(n5052), .Z(n3958) );
  AND U4137 ( .A(n3959), .B(n3958), .Z(n4034) );
  XOR U4138 ( .A(n4033), .B(n4034), .Z(n4036) );
  NAND U4139 ( .A(a[42]), .B(b[15]), .Z(n4035) );
  XOR U4140 ( .A(n4036), .B(n4035), .Z(n4027) );
  XNOR U4141 ( .A(n4028), .B(n4027), .Z(n4029) );
  NAND U4142 ( .A(n4521), .B(n3960), .Z(n3962) );
  XNOR U4143 ( .A(a[56]), .B(n208), .Z(n4045) );
  NANDN U4144 ( .A(n4488), .B(n4045), .Z(n3961) );
  NAND U4145 ( .A(n3962), .B(n3961), .Z(n4023) );
  IV U4146 ( .A(a[54]), .Z(n4542) );
  XNOR U4147 ( .A(n209), .B(n4542), .Z(n4048) );
  OR U4148 ( .A(n4048), .B(n4612), .Z(n3965) );
  NANDN U4149 ( .A(n3963), .B(n4669), .Z(n3964) );
  NAND U4150 ( .A(n3965), .B(n3964), .Z(n4021) );
  XNOR U4151 ( .A(n4744), .B(n4528), .Z(n4051) );
  NANDN U4152 ( .A(n4051), .B(n4745), .Z(n3968) );
  NANDN U4153 ( .A(n3966), .B(n4746), .Z(n3967) );
  AND U4154 ( .A(n3968), .B(n3967), .Z(n4022) );
  XOR U4155 ( .A(n4023), .B(n4024), .Z(n4030) );
  XOR U4156 ( .A(n4029), .B(n4030), .Z(n3996) );
  XNOR U4157 ( .A(n3997), .B(n3996), .Z(n3999) );
  XNOR U4158 ( .A(n3998), .B(n3999), .Z(n4056) );
  NANDN U4159 ( .A(n3970), .B(n3969), .Z(n3974) );
  NAND U4160 ( .A(n3972), .B(n3971), .Z(n3973) );
  NAND U4161 ( .A(n3974), .B(n3973), .Z(n4054) );
  NANDN U4162 ( .A(n3976), .B(n3975), .Z(n3980) );
  NANDN U4163 ( .A(n3978), .B(n3977), .Z(n3979) );
  NAND U4164 ( .A(n3980), .B(n3979), .Z(n4055) );
  XNOR U4165 ( .A(n4054), .B(n4055), .Z(n4057) );
  XOR U4166 ( .A(n4056), .B(n4057), .Z(n3992) );
  NANDN U4167 ( .A(n3982), .B(n3981), .Z(n3986) );
  NANDN U4168 ( .A(n3984), .B(n3983), .Z(n3985) );
  NAND U4169 ( .A(n3986), .B(n3985), .Z(n3993) );
  XOR U4170 ( .A(n3992), .B(n3993), .Z(n3994) );
  XNOR U4171 ( .A(n3995), .B(n3994), .Z(n4060) );
  XNOR U4172 ( .A(n4060), .B(sreg[106]), .Z(n4062) );
  NAND U4173 ( .A(n3987), .B(sreg[105]), .Z(n3991) );
  OR U4174 ( .A(n3989), .B(n3988), .Z(n3990) );
  AND U4175 ( .A(n3991), .B(n3990), .Z(n4061) );
  XOR U4176 ( .A(n4062), .B(n4061), .Z(c[106]) );
  NAND U4177 ( .A(n3997), .B(n3996), .Z(n4001) );
  NANDN U4178 ( .A(n3999), .B(n3998), .Z(n4000) );
  NAND U4179 ( .A(n4001), .B(n4000), .Z(n4130) );
  NANDN U4180 ( .A(n4003), .B(n4002), .Z(n4007) );
  NANDN U4181 ( .A(n4005), .B(n4004), .Z(n4006) );
  NAND U4182 ( .A(n4007), .B(n4006), .Z(n4131) );
  XNOR U4183 ( .A(n4130), .B(n4131), .Z(n4132) );
  XOR U4184 ( .A(n4859), .B(a[51]), .Z(n4083) );
  OR U4185 ( .A(n4083), .B(n4860), .Z(n4010) );
  NANDN U4186 ( .A(n4008), .B(n4915), .Z(n4009) );
  NAND U4187 ( .A(n4010), .B(n4009), .Z(n4096) );
  NANDN U4188 ( .A(n4011), .B(n4987), .Z(n4013) );
  XOR U4189 ( .A(n4909), .B(a[49]), .Z(n4086) );
  OR U4190 ( .A(n4086), .B(n4986), .Z(n4012) );
  NAND U4191 ( .A(n4013), .B(n4012), .Z(n4093) );
  XOR U4192 ( .A(n210), .B(a[45]), .Z(n4090) );
  OR U4193 ( .A(n4090), .B(n5095), .Z(n4016) );
  NANDN U4194 ( .A(n4014), .B(n5092), .Z(n4015) );
  AND U4195 ( .A(n4016), .B(n4015), .Z(n4094) );
  XOR U4196 ( .A(n4093), .B(n4094), .Z(n4095) );
  XOR U4197 ( .A(n4096), .B(n4095), .Z(n4077) );
  XNOR U4198 ( .A(n4077), .B(n4078), .Z(n4079) );
  NANDN U4199 ( .A(n4022), .B(n4021), .Z(n4026) );
  NANDN U4200 ( .A(n4024), .B(n4023), .Z(n4025) );
  NAND U4201 ( .A(n4026), .B(n4025), .Z(n4080) );
  XOR U4202 ( .A(n4079), .B(n4080), .Z(n4074) );
  NAND U4203 ( .A(n4028), .B(n4027), .Z(n4032) );
  OR U4204 ( .A(n4030), .B(n4029), .Z(n4031) );
  NAND U4205 ( .A(n4032), .B(n4031), .Z(n4071) );
  NANDN U4206 ( .A(n4034), .B(n4033), .Z(n4038) );
  OR U4207 ( .A(n4036), .B(n4035), .Z(n4037) );
  NAND U4208 ( .A(n4038), .B(n4037), .Z(n4127) );
  XOR U4209 ( .A(n5129), .B(a[47]), .Z(n4106) );
  OR U4210 ( .A(n4106), .B(n5041), .Z(n4041) );
  NANDN U4211 ( .A(n4039), .B(n5052), .Z(n4040) );
  AND U4212 ( .A(n4041), .B(n4040), .Z(n4119) );
  NAND U4213 ( .A(b[0]), .B(a[59]), .Z(n4042) );
  XNOR U4214 ( .A(b[1]), .B(n4042), .Z(n4044) );
  NAND U4215 ( .A(a[58]), .B(n206), .Z(n4043) );
  AND U4216 ( .A(n4044), .B(n4043), .Z(n4118) );
  XOR U4217 ( .A(n4119), .B(n4118), .Z(n4121) );
  NAND U4218 ( .A(a[43]), .B(b[15]), .Z(n4120) );
  XOR U4219 ( .A(n4121), .B(n4120), .Z(n4124) );
  NAND U4220 ( .A(n4521), .B(n4045), .Z(n4047) );
  IV U4221 ( .A(a[57]), .Z(n4852) );
  XNOR U4222 ( .A(n4852), .B(n208), .Z(n4109) );
  OR U4223 ( .A(n4109), .B(n4488), .Z(n4046) );
  NAND U4224 ( .A(n4047), .B(n4046), .Z(n4099) );
  IV U4225 ( .A(a[55]), .Z(n4731) );
  XNOR U4226 ( .A(b[5]), .B(n4731), .Z(n4112) );
  NANDN U4227 ( .A(n4612), .B(n4112), .Z(n4050) );
  NANDN U4228 ( .A(n4048), .B(n4669), .Z(n4049) );
  NAND U4229 ( .A(n4050), .B(n4049), .Z(n4097) );
  XOR U4230 ( .A(n4744), .B(a[53]), .Z(n4115) );
  NANDN U4231 ( .A(n4115), .B(n4745), .Z(n4053) );
  NANDN U4232 ( .A(n4051), .B(n4746), .Z(n4052) );
  AND U4233 ( .A(n4053), .B(n4052), .Z(n4098) );
  XOR U4234 ( .A(n4099), .B(n4100), .Z(n4125) );
  XNOR U4235 ( .A(n4124), .B(n4125), .Z(n4126) );
  XNOR U4236 ( .A(n4127), .B(n4126), .Z(n4072) );
  XNOR U4237 ( .A(n4071), .B(n4072), .Z(n4073) );
  XNOR U4238 ( .A(n4074), .B(n4073), .Z(n4133) );
  XOR U4239 ( .A(n4132), .B(n4133), .Z(n4065) );
  NANDN U4240 ( .A(n4055), .B(n4054), .Z(n4059) );
  NAND U4241 ( .A(n4057), .B(n4056), .Z(n4058) );
  NAND U4242 ( .A(n4059), .B(n4058), .Z(n4066) );
  XNOR U4243 ( .A(n4065), .B(n4066), .Z(n4067) );
  XNOR U4244 ( .A(n4068), .B(n4067), .Z(n4136) );
  XNOR U4245 ( .A(n4136), .B(sreg[107]), .Z(n4138) );
  NAND U4246 ( .A(n4060), .B(sreg[106]), .Z(n4064) );
  OR U4247 ( .A(n4062), .B(n4061), .Z(n4063) );
  AND U4248 ( .A(n4064), .B(n4063), .Z(n4137) );
  XOR U4249 ( .A(n4138), .B(n4137), .Z(c[107]) );
  NANDN U4250 ( .A(n4066), .B(n4065), .Z(n4070) );
  NAND U4251 ( .A(n4068), .B(n4067), .Z(n4069) );
  NAND U4252 ( .A(n4070), .B(n4069), .Z(n4144) );
  NANDN U4253 ( .A(n4072), .B(n4071), .Z(n4076) );
  NAND U4254 ( .A(n4074), .B(n4073), .Z(n4075) );
  NAND U4255 ( .A(n4076), .B(n4075), .Z(n4203) );
  NANDN U4256 ( .A(n4078), .B(n4077), .Z(n4082) );
  NANDN U4257 ( .A(n4080), .B(n4079), .Z(n4081) );
  NAND U4258 ( .A(n4082), .B(n4081), .Z(n4204) );
  XNOR U4259 ( .A(n4203), .B(n4204), .Z(n4205) );
  XNOR U4260 ( .A(n4859), .B(n4528), .Z(n4159) );
  OR U4261 ( .A(n4159), .B(n4860), .Z(n4085) );
  NANDN U4262 ( .A(n4083), .B(n4915), .Z(n4084) );
  NAND U4263 ( .A(n4085), .B(n4084), .Z(n4171) );
  NANDN U4264 ( .A(n4086), .B(n4987), .Z(n4088) );
  XNOR U4265 ( .A(n4909), .B(n4394), .Z(n4162) );
  OR U4266 ( .A(n4162), .B(n4986), .Z(n4087) );
  NAND U4267 ( .A(n4088), .B(n4087), .Z(n4168) );
  XNOR U4268 ( .A(n210), .B(n4089), .Z(n4165) );
  OR U4269 ( .A(n4165), .B(n5095), .Z(n4092) );
  NANDN U4270 ( .A(n4090), .B(n5092), .Z(n4091) );
  AND U4271 ( .A(n4092), .B(n4091), .Z(n4169) );
  XOR U4272 ( .A(n4168), .B(n4169), .Z(n4170) );
  XOR U4273 ( .A(n4171), .B(n4170), .Z(n4153) );
  XNOR U4274 ( .A(n4153), .B(n4154), .Z(n4155) );
  NANDN U4275 ( .A(n4098), .B(n4097), .Z(n4102) );
  NANDN U4276 ( .A(n4100), .B(n4099), .Z(n4101) );
  NAND U4277 ( .A(n4102), .B(n4101), .Z(n4156) );
  XOR U4278 ( .A(n4155), .B(n4156), .Z(n4150) );
  NAND U4279 ( .A(b[0]), .B(a[60]), .Z(n4103) );
  XNOR U4280 ( .A(b[1]), .B(n4103), .Z(n4105) );
  NAND U4281 ( .A(a[59]), .B(n206), .Z(n4104) );
  AND U4282 ( .A(n4105), .B(n4104), .Z(n4182) );
  XOR U4283 ( .A(n5129), .B(a[48]), .Z(n4191) );
  OR U4284 ( .A(n4191), .B(n5041), .Z(n4108) );
  NANDN U4285 ( .A(n4106), .B(n5052), .Z(n4107) );
  AND U4286 ( .A(n4108), .B(n4107), .Z(n4183) );
  XOR U4287 ( .A(n4182), .B(n4183), .Z(n4185) );
  NAND U4288 ( .A(b[15]), .B(a[44]), .Z(n4184) );
  XNOR U4289 ( .A(n4185), .B(n4184), .Z(n4179) );
  NANDN U4290 ( .A(n4109), .B(n4521), .Z(n4111) );
  XOR U4291 ( .A(a[58]), .B(b[3]), .Z(n4194) );
  NANDN U4292 ( .A(n4488), .B(n4194), .Z(n4110) );
  NAND U4293 ( .A(n4111), .B(n4110), .Z(n4174) );
  NAND U4294 ( .A(n4669), .B(n4112), .Z(n4114) );
  XOR U4295 ( .A(a[56]), .B(b[5]), .Z(n4197) );
  NANDN U4296 ( .A(n4612), .B(n4197), .Z(n4113) );
  AND U4297 ( .A(n4114), .B(n4113), .Z(n4172) );
  XOR U4298 ( .A(b[7]), .B(a[54]), .Z(n4200) );
  NAND U4299 ( .A(n4745), .B(n4200), .Z(n4117) );
  NANDN U4300 ( .A(n4115), .B(n4746), .Z(n4116) );
  NAND U4301 ( .A(n4117), .B(n4116), .Z(n4173) );
  XOR U4302 ( .A(n4172), .B(n4173), .Z(n4175) );
  XOR U4303 ( .A(n4174), .B(n4175), .Z(n4176) );
  NANDN U4304 ( .A(n4119), .B(n4118), .Z(n4123) );
  OR U4305 ( .A(n4121), .B(n4120), .Z(n4122) );
  NAND U4306 ( .A(n4123), .B(n4122), .Z(n4177) );
  XNOR U4307 ( .A(n4176), .B(n4177), .Z(n4178) );
  XNOR U4308 ( .A(n4179), .B(n4178), .Z(n4147) );
  NANDN U4309 ( .A(n4125), .B(n4124), .Z(n4129) );
  NAND U4310 ( .A(n4127), .B(n4126), .Z(n4128) );
  AND U4311 ( .A(n4129), .B(n4128), .Z(n4148) );
  XNOR U4312 ( .A(n4147), .B(n4148), .Z(n4149) );
  XNOR U4313 ( .A(n4150), .B(n4149), .Z(n4206) );
  XOR U4314 ( .A(n4205), .B(n4206), .Z(n4141) );
  NANDN U4315 ( .A(n4131), .B(n4130), .Z(n4135) );
  NANDN U4316 ( .A(n4133), .B(n4132), .Z(n4134) );
  NAND U4317 ( .A(n4135), .B(n4134), .Z(n4142) );
  XNOR U4318 ( .A(n4141), .B(n4142), .Z(n4143) );
  XNOR U4319 ( .A(n4144), .B(n4143), .Z(n4209) );
  XNOR U4320 ( .A(n4209), .B(sreg[108]), .Z(n4211) );
  NAND U4321 ( .A(n4136), .B(sreg[107]), .Z(n4140) );
  OR U4322 ( .A(n4138), .B(n4137), .Z(n4139) );
  AND U4323 ( .A(n4140), .B(n4139), .Z(n4210) );
  XOR U4324 ( .A(n4211), .B(n4210), .Z(c[108]) );
  NANDN U4325 ( .A(n4142), .B(n4141), .Z(n4146) );
  NAND U4326 ( .A(n4144), .B(n4143), .Z(n4145) );
  NAND U4327 ( .A(n4146), .B(n4145), .Z(n4217) );
  NANDN U4328 ( .A(n4148), .B(n4147), .Z(n4152) );
  NAND U4329 ( .A(n4150), .B(n4149), .Z(n4151) );
  NAND U4330 ( .A(n4152), .B(n4151), .Z(n4218) );
  NANDN U4331 ( .A(n4154), .B(n4153), .Z(n4158) );
  NANDN U4332 ( .A(n4156), .B(n4155), .Z(n4157) );
  NAND U4333 ( .A(n4158), .B(n4157), .Z(n4219) );
  XNOR U4334 ( .A(n4218), .B(n4219), .Z(n4220) );
  XOR U4335 ( .A(n4859), .B(a[53]), .Z(n4267) );
  OR U4336 ( .A(n4267), .B(n4860), .Z(n4161) );
  NANDN U4337 ( .A(n4159), .B(n4915), .Z(n4160) );
  NAND U4338 ( .A(n4161), .B(n4160), .Z(n4264) );
  NANDN U4339 ( .A(n4162), .B(n4987), .Z(n4164) );
  XOR U4340 ( .A(n4909), .B(a[51]), .Z(n4270) );
  OR U4341 ( .A(n4270), .B(n4986), .Z(n4163) );
  NAND U4342 ( .A(n4164), .B(n4163), .Z(n4261) );
  XOR U4343 ( .A(n210), .B(a[47]), .Z(n4273) );
  OR U4344 ( .A(n4273), .B(n5095), .Z(n4167) );
  NANDN U4345 ( .A(n4165), .B(n5092), .Z(n4166) );
  AND U4346 ( .A(n4167), .B(n4166), .Z(n4262) );
  XNOR U4347 ( .A(n4261), .B(n4262), .Z(n4263) );
  XOR U4348 ( .A(n4264), .B(n4263), .Z(n4224) );
  XNOR U4349 ( .A(n4224), .B(n4225), .Z(n4227) );
  XNOR U4350 ( .A(n4227), .B(n4226), .Z(n4233) );
  NANDN U4351 ( .A(n4177), .B(n4176), .Z(n4181) );
  NAND U4352 ( .A(n4179), .B(n4178), .Z(n4180) );
  NAND U4353 ( .A(n4181), .B(n4180), .Z(n4231) );
  NANDN U4354 ( .A(n4183), .B(n4182), .Z(n4187) );
  OR U4355 ( .A(n4185), .B(n4184), .Z(n4186) );
  NAND U4356 ( .A(n4187), .B(n4186), .Z(n4279) );
  NAND U4357 ( .A(b[0]), .B(a[61]), .Z(n4188) );
  XNOR U4358 ( .A(b[1]), .B(n4188), .Z(n4190) );
  NAND U4359 ( .A(a[60]), .B(n206), .Z(n4189) );
  AND U4360 ( .A(n4190), .B(n4189), .Z(n4236) );
  XOR U4361 ( .A(b[13]), .B(a[49]), .Z(n4243) );
  NANDN U4362 ( .A(n5041), .B(n4243), .Z(n4193) );
  NANDN U4363 ( .A(n4191), .B(n5052), .Z(n4192) );
  NAND U4364 ( .A(n4193), .B(n4192), .Z(n4234) );
  NAND U4365 ( .A(b[15]), .B(a[45]), .Z(n4235) );
  XNOR U4366 ( .A(n4234), .B(n4235), .Z(n4237) );
  XOR U4367 ( .A(n4236), .B(n4237), .Z(n4276) );
  NAND U4368 ( .A(n4194), .B(n4521), .Z(n4196) );
  XNOR U4369 ( .A(a[59]), .B(n208), .Z(n4246) );
  NANDN U4370 ( .A(n4488), .B(n4246), .Z(n4195) );
  NAND U4371 ( .A(n4196), .B(n4195), .Z(n4257) );
  XNOR U4372 ( .A(n4852), .B(n209), .Z(n4249) );
  OR U4373 ( .A(n4249), .B(n4612), .Z(n4199) );
  NAND U4374 ( .A(n4197), .B(n4669), .Z(n4198) );
  NAND U4375 ( .A(n4199), .B(n4198), .Z(n4255) );
  XNOR U4376 ( .A(n4744), .B(n4731), .Z(n4252) );
  NANDN U4377 ( .A(n4252), .B(n4745), .Z(n4202) );
  NAND U4378 ( .A(n4200), .B(n4746), .Z(n4201) );
  AND U4379 ( .A(n4202), .B(n4201), .Z(n4256) );
  XOR U4380 ( .A(n4257), .B(n4258), .Z(n4277) );
  XNOR U4381 ( .A(n4276), .B(n4277), .Z(n4278) );
  XOR U4382 ( .A(n4279), .B(n4278), .Z(n4230) );
  XOR U4383 ( .A(n4231), .B(n4230), .Z(n4232) );
  XNOR U4384 ( .A(n4233), .B(n4232), .Z(n4221) );
  XOR U4385 ( .A(n4220), .B(n4221), .Z(n4214) );
  NANDN U4386 ( .A(n4204), .B(n4203), .Z(n4208) );
  NANDN U4387 ( .A(n4206), .B(n4205), .Z(n4207) );
  NAND U4388 ( .A(n4208), .B(n4207), .Z(n4215) );
  XOR U4389 ( .A(n4214), .B(n4215), .Z(n4216) );
  XNOR U4390 ( .A(n4217), .B(n4216), .Z(n4282) );
  XNOR U4391 ( .A(n4282), .B(sreg[109]), .Z(n4284) );
  NAND U4392 ( .A(n4209), .B(sreg[108]), .Z(n4213) );
  OR U4393 ( .A(n4211), .B(n4210), .Z(n4212) );
  AND U4394 ( .A(n4213), .B(n4212), .Z(n4283) );
  XOR U4395 ( .A(n4284), .B(n4283), .Z(c[109]) );
  NANDN U4396 ( .A(n4219), .B(n4218), .Z(n4223) );
  NAND U4397 ( .A(n4221), .B(n4220), .Z(n4222) );
  NAND U4398 ( .A(n4223), .B(n4222), .Z(n4288) );
  OR U4399 ( .A(n4225), .B(n4224), .Z(n4229) );
  OR U4400 ( .A(n4227), .B(n4226), .Z(n4228) );
  NAND U4401 ( .A(n4229), .B(n4228), .Z(n4291) );
  XNOR U4402 ( .A(n4291), .B(n4292), .Z(n4293) );
  NANDN U4403 ( .A(n4235), .B(n4234), .Z(n4239) );
  NAND U4404 ( .A(n4237), .B(n4236), .Z(n4238) );
  NAND U4405 ( .A(n4239), .B(n4238), .Z(n4321) );
  AND U4406 ( .A(b[15]), .B(a[46]), .Z(n4340) );
  NAND U4407 ( .A(a[62]), .B(b[0]), .Z(n4240) );
  XNOR U4408 ( .A(b[1]), .B(n4240), .Z(n4242) );
  NAND U4409 ( .A(a[61]), .B(n206), .Z(n4241) );
  AND U4410 ( .A(n4242), .B(n4241), .Z(n4338) );
  NAND U4411 ( .A(n5052), .B(n4243), .Z(n4245) );
  XOR U4412 ( .A(b[13]), .B(a[50]), .Z(n4325) );
  NANDN U4413 ( .A(n5041), .B(n4325), .Z(n4244) );
  AND U4414 ( .A(n4245), .B(n4244), .Z(n4337) );
  XNOR U4415 ( .A(n4338), .B(n4337), .Z(n4339) );
  XOR U4416 ( .A(n4340), .B(n4339), .Z(n4318) );
  NAND U4417 ( .A(n4521), .B(n4246), .Z(n4248) );
  XNOR U4418 ( .A(a[60]), .B(n208), .Z(n4328) );
  NANDN U4419 ( .A(n4488), .B(n4328), .Z(n4247) );
  NAND U4420 ( .A(n4248), .B(n4247), .Z(n4315) );
  IV U4421 ( .A(a[58]), .Z(n4990) );
  XNOR U4422 ( .A(n4990), .B(n209), .Z(n4331) );
  OR U4423 ( .A(n4331), .B(n4612), .Z(n4251) );
  NANDN U4424 ( .A(n4249), .B(n4669), .Z(n4250) );
  NAND U4425 ( .A(n4251), .B(n4250), .Z(n4312) );
  IV U4426 ( .A(a[56]), .Z(n4525) );
  XNOR U4427 ( .A(n4744), .B(n4525), .Z(n4334) );
  NANDN U4428 ( .A(n4334), .B(n4745), .Z(n4254) );
  NANDN U4429 ( .A(n4252), .B(n4746), .Z(n4253) );
  AND U4430 ( .A(n4254), .B(n4253), .Z(n4313) );
  XNOR U4431 ( .A(n4312), .B(n4313), .Z(n4314) );
  XNOR U4432 ( .A(n4315), .B(n4314), .Z(n4319) );
  XOR U4433 ( .A(n4318), .B(n4319), .Z(n4320) );
  XOR U4434 ( .A(n4321), .B(n4320), .Z(n4346) );
  NANDN U4435 ( .A(n4256), .B(n4255), .Z(n4260) );
  NANDN U4436 ( .A(n4258), .B(n4257), .Z(n4259) );
  NAND U4437 ( .A(n4260), .B(n4259), .Z(n4352) );
  NANDN U4438 ( .A(n4262), .B(n4261), .Z(n4266) );
  NAND U4439 ( .A(n4264), .B(n4263), .Z(n4265) );
  NAND U4440 ( .A(n4266), .B(n4265), .Z(n4350) );
  XNOR U4441 ( .A(n4859), .B(n4542), .Z(n4297) );
  OR U4442 ( .A(n4297), .B(n4860), .Z(n4269) );
  NANDN U4443 ( .A(n4267), .B(n4915), .Z(n4268) );
  NAND U4444 ( .A(n4269), .B(n4268), .Z(n4309) );
  NANDN U4445 ( .A(n4270), .B(n4987), .Z(n4272) );
  XNOR U4446 ( .A(n4909), .B(n4528), .Z(n4300) );
  OR U4447 ( .A(n4300), .B(n4986), .Z(n4271) );
  NAND U4448 ( .A(n4272), .B(n4271), .Z(n4306) );
  XOR U4449 ( .A(n210), .B(a[48]), .Z(n4303) );
  OR U4450 ( .A(n4303), .B(n5095), .Z(n4275) );
  NANDN U4451 ( .A(n4273), .B(n5092), .Z(n4274) );
  AND U4452 ( .A(n4275), .B(n4274), .Z(n4307) );
  XNOR U4453 ( .A(n4306), .B(n4307), .Z(n4308) );
  XOR U4454 ( .A(n4309), .B(n4308), .Z(n4349) );
  XNOR U4455 ( .A(n4350), .B(n4349), .Z(n4351) );
  XNOR U4456 ( .A(n4352), .B(n4351), .Z(n4344) );
  NANDN U4457 ( .A(n4277), .B(n4276), .Z(n4281) );
  NAND U4458 ( .A(n4279), .B(n4278), .Z(n4280) );
  AND U4459 ( .A(n4281), .B(n4280), .Z(n4343) );
  XNOR U4460 ( .A(n4344), .B(n4343), .Z(n4345) );
  XOR U4461 ( .A(n4346), .B(n4345), .Z(n4294) );
  XOR U4462 ( .A(n4293), .B(n4294), .Z(n4287) );
  XOR U4463 ( .A(n4288), .B(n4287), .Z(n4289) );
  XOR U4464 ( .A(n4290), .B(n4289), .Z(n4355) );
  XNOR U4465 ( .A(n4355), .B(sreg[110]), .Z(n4357) );
  NAND U4466 ( .A(n4282), .B(sreg[109]), .Z(n4286) );
  OR U4467 ( .A(n4284), .B(n4283), .Z(n4285) );
  AND U4468 ( .A(n4286), .B(n4285), .Z(n4356) );
  XOR U4469 ( .A(n4357), .B(n4356), .Z(c[110]) );
  NANDN U4470 ( .A(n4292), .B(n4291), .Z(n4296) );
  NAND U4471 ( .A(n4294), .B(n4293), .Z(n4295) );
  NAND U4472 ( .A(n4296), .B(n4295), .Z(n4361) );
  XNOR U4473 ( .A(n4859), .B(n4731), .Z(n4388) );
  OR U4474 ( .A(n4388), .B(n4860), .Z(n4299) );
  NANDN U4475 ( .A(n4297), .B(n4915), .Z(n4298) );
  NAND U4476 ( .A(n4299), .B(n4298), .Z(n4387) );
  NANDN U4477 ( .A(n4300), .B(n4987), .Z(n4302) );
  XOR U4478 ( .A(n4909), .B(a[53]), .Z(n4391) );
  OR U4479 ( .A(n4391), .B(n4986), .Z(n4301) );
  NAND U4480 ( .A(n4302), .B(n4301), .Z(n4384) );
  XOR U4481 ( .A(n210), .B(a[49]), .Z(n4395) );
  OR U4482 ( .A(n4395), .B(n5095), .Z(n4305) );
  NANDN U4483 ( .A(n4303), .B(n5092), .Z(n4304) );
  AND U4484 ( .A(n4305), .B(n4304), .Z(n4385) );
  XOR U4485 ( .A(n4384), .B(n4385), .Z(n4386) );
  XOR U4486 ( .A(n4387), .B(n4386), .Z(n4378) );
  NANDN U4487 ( .A(n4307), .B(n4306), .Z(n4311) );
  NAND U4488 ( .A(n4309), .B(n4308), .Z(n4310) );
  NAND U4489 ( .A(n4311), .B(n4310), .Z(n4379) );
  XOR U4490 ( .A(n4378), .B(n4379), .Z(n4381) );
  NANDN U4491 ( .A(n4313), .B(n4312), .Z(n4317) );
  NAND U4492 ( .A(n4315), .B(n4314), .Z(n4316) );
  NAND U4493 ( .A(n4317), .B(n4316), .Z(n4380) );
  XNOR U4494 ( .A(n4381), .B(n4380), .Z(n4375) );
  NAND U4495 ( .A(b[0]), .B(a[63]), .Z(n4322) );
  XNOR U4496 ( .A(b[1]), .B(n4322), .Z(n4324) );
  NAND U4497 ( .A(a[62]), .B(n206), .Z(n4323) );
  AND U4498 ( .A(n4324), .B(n4323), .Z(n4412) );
  XOR U4499 ( .A(n5129), .B(a[51]), .Z(n4425) );
  OR U4500 ( .A(n4425), .B(n5041), .Z(n4327) );
  NAND U4501 ( .A(n4325), .B(n5052), .Z(n4326) );
  NAND U4502 ( .A(n4327), .B(n4326), .Z(n4410) );
  NAND U4503 ( .A(b[15]), .B(a[47]), .Z(n4411) );
  XNOR U4504 ( .A(n4410), .B(n4411), .Z(n4413) );
  XOR U4505 ( .A(n4412), .B(n4413), .Z(n4404) );
  NAND U4506 ( .A(n4521), .B(n4328), .Z(n4330) );
  XNOR U4507 ( .A(a[61]), .B(n208), .Z(n4416) );
  NANDN U4508 ( .A(n4488), .B(n4416), .Z(n4329) );
  NAND U4509 ( .A(n4330), .B(n4329), .Z(n4400) );
  IV U4510 ( .A(a[59]), .Z(n4952) );
  XNOR U4511 ( .A(n4952), .B(n209), .Z(n4419) );
  OR U4512 ( .A(n4419), .B(n4612), .Z(n4333) );
  NANDN U4513 ( .A(n4331), .B(n4669), .Z(n4332) );
  NAND U4514 ( .A(n4333), .B(n4332), .Z(n4398) );
  XNOR U4515 ( .A(n4744), .B(n4852), .Z(n4422) );
  NANDN U4516 ( .A(n4422), .B(n4745), .Z(n4336) );
  NANDN U4517 ( .A(n4334), .B(n4746), .Z(n4335) );
  AND U4518 ( .A(n4336), .B(n4335), .Z(n4399) );
  XOR U4519 ( .A(n4400), .B(n4401), .Z(n4405) );
  XNOR U4520 ( .A(n4404), .B(n4405), .Z(n4406) );
  NANDN U4521 ( .A(n4338), .B(n4337), .Z(n4342) );
  NANDN U4522 ( .A(n4340), .B(n4339), .Z(n4341) );
  AND U4523 ( .A(n4342), .B(n4341), .Z(n4407) );
  XNOR U4524 ( .A(n4406), .B(n4407), .Z(n4373) );
  XNOR U4525 ( .A(n4372), .B(n4373), .Z(n4374) );
  XNOR U4526 ( .A(n4375), .B(n4374), .Z(n4369) );
  NANDN U4527 ( .A(n4344), .B(n4343), .Z(n4348) );
  NAND U4528 ( .A(n4346), .B(n4345), .Z(n4347) );
  NAND U4529 ( .A(n4348), .B(n4347), .Z(n4366) );
  OR U4530 ( .A(n4350), .B(n4349), .Z(n4354) );
  OR U4531 ( .A(n4352), .B(n4351), .Z(n4353) );
  AND U4532 ( .A(n4354), .B(n4353), .Z(n4367) );
  XNOR U4533 ( .A(n4366), .B(n4367), .Z(n4368) );
  XOR U4534 ( .A(n4369), .B(n4368), .Z(n4360) );
  XOR U4535 ( .A(n4361), .B(n4360), .Z(n4362) );
  XNOR U4536 ( .A(n4363), .B(n4362), .Z(n4428) );
  XNOR U4537 ( .A(n4428), .B(sreg[111]), .Z(n4430) );
  NAND U4538 ( .A(n4355), .B(sreg[110]), .Z(n4359) );
  OR U4539 ( .A(n4357), .B(n4356), .Z(n4358) );
  AND U4540 ( .A(n4359), .B(n4358), .Z(n4429) );
  XOR U4541 ( .A(n4430), .B(n4429), .Z(c[111]) );
  NAND U4542 ( .A(n4361), .B(n4360), .Z(n4365) );
  NAND U4543 ( .A(n4363), .B(n4362), .Z(n4364) );
  NAND U4544 ( .A(n4365), .B(n4364), .Z(n4438) );
  NANDN U4545 ( .A(n4367), .B(n4366), .Z(n4371) );
  NAND U4546 ( .A(n4369), .B(n4368), .Z(n4370) );
  NAND U4547 ( .A(n4371), .B(n4370), .Z(n4436) );
  NANDN U4548 ( .A(n4373), .B(n4372), .Z(n4377) );
  NAND U4549 ( .A(n4375), .B(n4374), .Z(n4376) );
  NAND U4550 ( .A(n4377), .B(n4376), .Z(n4443) );
  NANDN U4551 ( .A(n4379), .B(n4378), .Z(n4383) );
  OR U4552 ( .A(n4381), .B(n4380), .Z(n4382) );
  NAND U4553 ( .A(n4383), .B(n4382), .Z(n4442) );
  XNOR U4554 ( .A(n4859), .B(n4525), .Z(n4469) );
  OR U4555 ( .A(n4469), .B(n4860), .Z(n4390) );
  NANDN U4556 ( .A(n4388), .B(n4915), .Z(n4389) );
  NAND U4557 ( .A(n4390), .B(n4389), .Z(n4475) );
  NANDN U4558 ( .A(n4391), .B(n4987), .Z(n4393) );
  XNOR U4559 ( .A(n4909), .B(n4542), .Z(n4466) );
  OR U4560 ( .A(n4466), .B(n4986), .Z(n4392) );
  NAND U4561 ( .A(n4393), .B(n4392), .Z(n4472) );
  XNOR U4562 ( .A(b[15]), .B(n4394), .Z(n4497) );
  NANDN U4563 ( .A(n5095), .B(n4497), .Z(n4397) );
  NANDN U4564 ( .A(n4395), .B(n5092), .Z(n4396) );
  AND U4565 ( .A(n4397), .B(n4396), .Z(n4473) );
  XNOR U4566 ( .A(n4472), .B(n4473), .Z(n4474) );
  XOR U4567 ( .A(n4475), .B(n4474), .Z(n4451) );
  XNOR U4568 ( .A(n4452), .B(n4451), .Z(n4454) );
  NANDN U4569 ( .A(n4399), .B(n4398), .Z(n4403) );
  NANDN U4570 ( .A(n4401), .B(n4400), .Z(n4402) );
  NAND U4571 ( .A(n4403), .B(n4402), .Z(n4453) );
  XOR U4572 ( .A(n4454), .B(n4453), .Z(n4445) );
  NANDN U4573 ( .A(n4405), .B(n4404), .Z(n4409) );
  NAND U4574 ( .A(n4407), .B(n4406), .Z(n4408) );
  AND U4575 ( .A(n4409), .B(n4408), .Z(n4446) );
  XNOR U4576 ( .A(n4445), .B(n4446), .Z(n4448) );
  NANDN U4577 ( .A(n4411), .B(n4410), .Z(n4415) );
  NAND U4578 ( .A(n4413), .B(n4412), .Z(n4414) );
  NAND U4579 ( .A(n4415), .B(n4414), .Z(n4480) );
  NAND U4580 ( .A(n4521), .B(n4416), .Z(n4418) );
  XNOR U4581 ( .A(a[62]), .B(n208), .Z(n4487) );
  NANDN U4582 ( .A(n4488), .B(n4487), .Z(n4417) );
  NAND U4583 ( .A(n4418), .B(n4417), .Z(n4459) );
  IV U4584 ( .A(a[60]), .Z(n4992) );
  XNOR U4585 ( .A(n4992), .B(n209), .Z(n4484) );
  OR U4586 ( .A(n4484), .B(n4612), .Z(n4421) );
  NANDN U4587 ( .A(n4419), .B(n4669), .Z(n4420) );
  NAND U4588 ( .A(n4421), .B(n4420), .Z(n4457) );
  XNOR U4589 ( .A(n4990), .B(n4744), .Z(n4463) );
  NANDN U4590 ( .A(n4463), .B(n4745), .Z(n4424) );
  NANDN U4591 ( .A(n4422), .B(n4746), .Z(n4423) );
  AND U4592 ( .A(n4424), .B(n4423), .Z(n4458) );
  XOR U4593 ( .A(n4459), .B(n4460), .Z(n4478) );
  IV U4594 ( .A(a[63]), .Z(n5094) );
  XNOR U4595 ( .A(n5129), .B(n4528), .Z(n4500) );
  OR U4596 ( .A(n4500), .B(n5041), .Z(n4427) );
  NANDN U4597 ( .A(n4425), .B(n5052), .Z(n4426) );
  NAND U4598 ( .A(n4427), .B(n4426), .Z(n4491) );
  NAND U4599 ( .A(b[15]), .B(a[48]), .Z(n4492) );
  XNOR U4600 ( .A(n4491), .B(n4492), .Z(n4493) );
  XOR U4601 ( .A(n4494), .B(n4493), .Z(n4479) );
  XOR U4602 ( .A(n4478), .B(n4479), .Z(n4481) );
  XOR U4603 ( .A(n4480), .B(n4481), .Z(n4447) );
  XOR U4604 ( .A(n4448), .B(n4447), .Z(n4441) );
  XOR U4605 ( .A(n4442), .B(n4441), .Z(n4444) );
  XOR U4606 ( .A(n4443), .B(n4444), .Z(n4435) );
  XOR U4607 ( .A(n4436), .B(n4435), .Z(n4437) );
  XOR U4608 ( .A(n4438), .B(n4437), .Z(n4434) );
  NAND U4609 ( .A(n4428), .B(sreg[111]), .Z(n4432) );
  OR U4610 ( .A(n4430), .B(n4429), .Z(n4431) );
  AND U4611 ( .A(n4432), .B(n4431), .Z(n4433) );
  XOR U4612 ( .A(n4434), .B(n4433), .Z(c[112]) );
  OR U4613 ( .A(n4434), .B(n4433), .Z(n4572) );
  NAND U4614 ( .A(n4436), .B(n4435), .Z(n4440) );
  NAND U4615 ( .A(n4438), .B(n4437), .Z(n4439) );
  NAND U4616 ( .A(n4440), .B(n4439), .Z(n4506) );
  NAND U4617 ( .A(n4446), .B(n4445), .Z(n4450) );
  NANDN U4618 ( .A(n4448), .B(n4447), .Z(n4449) );
  NAND U4619 ( .A(n4450), .B(n4449), .Z(n4564) );
  OR U4620 ( .A(n4452), .B(n4451), .Z(n4456) );
  OR U4621 ( .A(n4454), .B(n4453), .Z(n4455) );
  AND U4622 ( .A(n4456), .B(n4455), .Z(n4565) );
  XNOR U4623 ( .A(n4564), .B(n4565), .Z(n4566) );
  NANDN U4624 ( .A(n4458), .B(n4457), .Z(n4462) );
  NANDN U4625 ( .A(n4460), .B(n4459), .Z(n4461) );
  NAND U4626 ( .A(n4462), .B(n4461), .Z(n4557) );
  XNOR U4627 ( .A(n4952), .B(n4744), .Z(n4535) );
  NANDN U4628 ( .A(n4535), .B(n4745), .Z(n4465) );
  NANDN U4629 ( .A(n4463), .B(n4746), .Z(n4464) );
  NAND U4630 ( .A(n4465), .B(n4464), .Z(n4553) );
  NANDN U4631 ( .A(n4466), .B(n4987), .Z(n4468) );
  XNOR U4632 ( .A(n4909), .B(n4731), .Z(n4524) );
  OR U4633 ( .A(n4524), .B(n4986), .Z(n4467) );
  NAND U4634 ( .A(n4468), .B(n4467), .Z(n4550) );
  XNOR U4635 ( .A(n4859), .B(n4852), .Z(n4532) );
  OR U4636 ( .A(n4532), .B(n4860), .Z(n4471) );
  NANDN U4637 ( .A(n4469), .B(n4915), .Z(n4470) );
  AND U4638 ( .A(n4471), .B(n4470), .Z(n4551) );
  XOR U4639 ( .A(n4550), .B(n4551), .Z(n4552) );
  XOR U4640 ( .A(n4553), .B(n4552), .Z(n4554) );
  NANDN U4641 ( .A(n4473), .B(n4472), .Z(n4477) );
  NAND U4642 ( .A(n4475), .B(n4474), .Z(n4476) );
  NAND U4643 ( .A(n4477), .B(n4476), .Z(n4555) );
  XNOR U4644 ( .A(n4554), .B(n4555), .Z(n4556) );
  XOR U4645 ( .A(n4557), .B(n4556), .Z(n4562) );
  NANDN U4646 ( .A(n4479), .B(n4478), .Z(n4483) );
  OR U4647 ( .A(n4481), .B(n4480), .Z(n4482) );
  NAND U4648 ( .A(n4483), .B(n4482), .Z(n4561) );
  IV U4649 ( .A(a[61]), .Z(n5037) );
  XNOR U4650 ( .A(n5037), .B(n209), .Z(n4538) );
  OR U4651 ( .A(n4538), .B(n4612), .Z(n4486) );
  NANDN U4652 ( .A(n4484), .B(n4669), .Z(n4485) );
  NAND U4653 ( .A(n4486), .B(n4485), .Z(n4545) );
  XNOR U4654 ( .A(n207), .B(n4545), .Z(n4547) );
  NAND U4655 ( .A(n4521), .B(n4487), .Z(n4490) );
  XNOR U4656 ( .A(a[63]), .B(n208), .Z(n4520) );
  NANDN U4657 ( .A(n4488), .B(n4520), .Z(n4489) );
  NAND U4658 ( .A(n4490), .B(n4489), .Z(n4546) );
  XOR U4659 ( .A(n4547), .B(n4546), .Z(n4509) );
  NANDN U4660 ( .A(n4492), .B(n4491), .Z(n4496) );
  NAND U4661 ( .A(n4494), .B(n4493), .Z(n4495) );
  AND U4662 ( .A(n4496), .B(n4495), .Z(n4510) );
  XNOR U4663 ( .A(n4509), .B(n4510), .Z(n4512) );
  NAND U4664 ( .A(n5092), .B(n4497), .Z(n4499) );
  XOR U4665 ( .A(b[15]), .B(a[51]), .Z(n4529) );
  NANDN U4666 ( .A(n5095), .B(n4529), .Z(n4498) );
  NAND U4667 ( .A(n4499), .B(n4498), .Z(n4517) );
  ANDN U4668 ( .B(a[49]), .A(n210), .Z(n4679) );
  IV U4669 ( .A(n4679), .Z(n4607) );
  NANDN U4670 ( .A(n4500), .B(n5052), .Z(n4502) );
  XOR U4671 ( .A(b[13]), .B(a[53]), .Z(n4541) );
  NANDN U4672 ( .A(n5041), .B(n4541), .Z(n4501) );
  NAND U4673 ( .A(n4502), .B(n4501), .Z(n4515) );
  XOR U4674 ( .A(n4607), .B(n4515), .Z(n4516) );
  XOR U4675 ( .A(n4512), .B(n4511), .Z(n4560) );
  XOR U4676 ( .A(n4561), .B(n4560), .Z(n4563) );
  XOR U4677 ( .A(n4562), .B(n4563), .Z(n4567) );
  XOR U4678 ( .A(n4566), .B(n4567), .Z(n4503) );
  XOR U4679 ( .A(n4504), .B(n4503), .Z(n4505) );
  XOR U4680 ( .A(n4506), .B(n4505), .Z(n4571) );
  XOR U4681 ( .A(n4572), .B(n4571), .Z(c[113]) );
  NAND U4682 ( .A(n4504), .B(n4503), .Z(n4508) );
  NAND U4683 ( .A(n4506), .B(n4505), .Z(n4507) );
  NAND U4684 ( .A(n4508), .B(n4507), .Z(n4579) );
  NAND U4685 ( .A(n4510), .B(n4509), .Z(n4514) );
  NANDN U4686 ( .A(n4512), .B(n4511), .Z(n4513) );
  NAND U4687 ( .A(n4514), .B(n4513), .Z(n4627) );
  NANDN U4688 ( .A(n4515), .B(n4679), .Z(n4519) );
  NANDN U4689 ( .A(n4517), .B(n4516), .Z(n4518) );
  AND U4690 ( .A(n4519), .B(n4518), .Z(n4628) );
  XNOR U4691 ( .A(n4627), .B(n4628), .Z(n4629) );
  NAND U4692 ( .A(a[50]), .B(b[15]), .Z(n4590) );
  NAND U4693 ( .A(n4521), .B(n4520), .Z(n4522) );
  NANDN U4694 ( .A(n4523), .B(n4522), .Z(n4588) );
  XOR U4695 ( .A(n4607), .B(n4588), .Z(n4589) );
  XNOR U4696 ( .A(n4590), .B(n4589), .Z(n4596) );
  NANDN U4697 ( .A(n4524), .B(n4987), .Z(n4527) );
  XNOR U4698 ( .A(n4909), .B(n4525), .Z(n4608) );
  OR U4699 ( .A(n4608), .B(n4986), .Z(n4526) );
  NAND U4700 ( .A(n4527), .B(n4526), .Z(n4593) );
  XNOR U4701 ( .A(n210), .B(n4528), .Z(n4615) );
  OR U4702 ( .A(n4615), .B(n5095), .Z(n4531) );
  NAND U4703 ( .A(n4529), .B(n5092), .Z(n4530) );
  AND U4704 ( .A(n4531), .B(n4530), .Z(n4594) );
  XNOR U4705 ( .A(n4593), .B(n4594), .Z(n4595) );
  XOR U4706 ( .A(n4596), .B(n4595), .Z(n4601) );
  XNOR U4707 ( .A(b[9]), .B(n4990), .Z(n4621) );
  NANDN U4708 ( .A(n4860), .B(n4621), .Z(n4534) );
  NANDN U4709 ( .A(n4532), .B(n4915), .Z(n4533) );
  NAND U4710 ( .A(n4534), .B(n4533), .Z(n4585) );
  XNOR U4711 ( .A(n4992), .B(n4744), .Z(n4624) );
  NANDN U4712 ( .A(n4624), .B(n4745), .Z(n4537) );
  NANDN U4713 ( .A(n4535), .B(n4746), .Z(n4536) );
  NAND U4714 ( .A(n4537), .B(n4536), .Z(n4582) );
  XNOR U4715 ( .A(a[62]), .B(n209), .Z(n4611) );
  NANDN U4716 ( .A(n4612), .B(n4611), .Z(n4540) );
  NANDN U4717 ( .A(n4538), .B(n4669), .Z(n4539) );
  AND U4718 ( .A(n4540), .B(n4539), .Z(n4583) );
  XNOR U4719 ( .A(n4582), .B(n4583), .Z(n4584) );
  XNOR U4720 ( .A(n4585), .B(n4584), .Z(n4599) );
  NAND U4721 ( .A(n5052), .B(n4541), .Z(n4544) );
  XNOR U4722 ( .A(b[13]), .B(n4542), .Z(n4618) );
  NANDN U4723 ( .A(n5041), .B(n4618), .Z(n4543) );
  NAND U4724 ( .A(n4544), .B(n4543), .Z(n4600) );
  XOR U4725 ( .A(n4599), .B(n4600), .Z(n4602) );
  XOR U4726 ( .A(n4601), .B(n4602), .Z(n4635) );
  NANDN U4727 ( .A(n4545), .B(b[1]), .Z(n4549) );
  OR U4728 ( .A(n4547), .B(n4546), .Z(n4548) );
  AND U4729 ( .A(n4549), .B(n4548), .Z(n4633) );
  XNOR U4730 ( .A(n4633), .B(n4634), .Z(n4636) );
  XOR U4731 ( .A(n4629), .B(n4630), .Z(n4642) );
  NANDN U4732 ( .A(n4555), .B(n4554), .Z(n4559) );
  NANDN U4733 ( .A(n4557), .B(n4556), .Z(n4558) );
  NAND U4734 ( .A(n4559), .B(n4558), .Z(n4640) );
  XNOR U4735 ( .A(n4640), .B(n4639), .Z(n4641) );
  XNOR U4736 ( .A(n4642), .B(n4641), .Z(n4577) );
  IV U4737 ( .A(n4577), .Z(n4575) );
  NANDN U4738 ( .A(n4565), .B(n4564), .Z(n4569) );
  NAND U4739 ( .A(n4567), .B(n4566), .Z(n4568) );
  AND U4740 ( .A(n4569), .B(n4568), .Z(n4576) );
  XNOR U4741 ( .A(n4575), .B(n4576), .Z(n4570) );
  XNOR U4742 ( .A(n4579), .B(n4570), .Z(n4574) );
  OR U4743 ( .A(n4572), .B(n4571), .Z(n4573) );
  XOR U4744 ( .A(n4574), .B(n4573), .Z(c[114]) );
  OR U4745 ( .A(n4574), .B(n4573), .Z(n4709) );
  NAND U4746 ( .A(n4575), .B(n4576), .Z(n4581) );
  ANDN U4747 ( .B(n4577), .A(n4576), .Z(n4578) );
  OR U4748 ( .A(n4579), .B(n4578), .Z(n4580) );
  NAND U4749 ( .A(n4581), .B(n4580), .Z(n4648) );
  NANDN U4750 ( .A(n4583), .B(n4582), .Z(n4587) );
  NAND U4751 ( .A(n4585), .B(n4584), .Z(n4586) );
  NAND U4752 ( .A(n4587), .B(n4586), .Z(n4698) );
  NANDN U4753 ( .A(n4588), .B(n4679), .Z(n4592) );
  NAND U4754 ( .A(n4590), .B(n4589), .Z(n4591) );
  NAND U4755 ( .A(n4592), .B(n4591), .Z(n4695) );
  NANDN U4756 ( .A(n4594), .B(n4593), .Z(n4598) );
  NAND U4757 ( .A(n4596), .B(n4595), .Z(n4597) );
  NAND U4758 ( .A(n4598), .B(n4597), .Z(n4696) );
  XNOR U4759 ( .A(n4695), .B(n4696), .Z(n4697) );
  XOR U4760 ( .A(n4698), .B(n4697), .Z(n4651) );
  NANDN U4761 ( .A(n4600), .B(n4599), .Z(n4604) );
  OR U4762 ( .A(n4602), .B(n4601), .Z(n4603) );
  NAND U4763 ( .A(n4604), .B(n4603), .Z(n4652) );
  XNOR U4764 ( .A(n4651), .B(n4652), .Z(n4653) );
  NAND U4765 ( .A(b[15]), .B(a[51]), .Z(n4682) );
  NAND U4766 ( .A(n207), .B(b[3]), .Z(n4605) );
  NANDN U4767 ( .A(n4606), .B(n4605), .Z(n4680) );
  XOR U4768 ( .A(n4607), .B(n4680), .Z(n4681) );
  XOR U4769 ( .A(n4682), .B(n4681), .Z(n4688) );
  NANDN U4770 ( .A(n4608), .B(n4987), .Z(n4610) );
  XNOR U4771 ( .A(n4909), .B(n4852), .Z(n4657) );
  OR U4772 ( .A(n4657), .B(n4986), .Z(n4609) );
  NAND U4773 ( .A(n4610), .B(n4609), .Z(n4686) );
  NAND U4774 ( .A(n4669), .B(n4611), .Z(n4614) );
  XNOR U4775 ( .A(n5094), .B(n209), .Z(n4670) );
  OR U4776 ( .A(n4670), .B(n4612), .Z(n4613) );
  NAND U4777 ( .A(n4614), .B(n4613), .Z(n4685) );
  XNOR U4778 ( .A(n4686), .B(n4685), .Z(n4687) );
  XNOR U4779 ( .A(n4688), .B(n4687), .Z(n4677) );
  XOR U4780 ( .A(b[15]), .B(a[53]), .Z(n4672) );
  NANDN U4781 ( .A(n5095), .B(n4672), .Z(n4617) );
  NANDN U4782 ( .A(n4615), .B(n5092), .Z(n4616) );
  NAND U4783 ( .A(n4617), .B(n4616), .Z(n4676) );
  NAND U4784 ( .A(n5052), .B(n4618), .Z(n4620) );
  XNOR U4785 ( .A(b[13]), .B(n4731), .Z(n4666) );
  NANDN U4786 ( .A(n5041), .B(n4666), .Z(n4619) );
  AND U4787 ( .A(n4620), .B(n4619), .Z(n4693) );
  NAND U4788 ( .A(n4915), .B(n4621), .Z(n4623) );
  XOR U4789 ( .A(b[9]), .B(a[59]), .Z(n4660) );
  NANDN U4790 ( .A(n4860), .B(n4660), .Z(n4622) );
  AND U4791 ( .A(n4623), .B(n4622), .Z(n4691) );
  XNOR U4792 ( .A(n5037), .B(n4744), .Z(n4663) );
  NANDN U4793 ( .A(n4663), .B(n4745), .Z(n4626) );
  NANDN U4794 ( .A(n4624), .B(n4746), .Z(n4625) );
  AND U4795 ( .A(n4626), .B(n4625), .Z(n4692) );
  XOR U4796 ( .A(n4691), .B(n4692), .Z(n4694) );
  XOR U4797 ( .A(n4693), .B(n4694), .Z(n4675) );
  XOR U4798 ( .A(n4676), .B(n4675), .Z(n4678) );
  XOR U4799 ( .A(n4677), .B(n4678), .Z(n4654) );
  XNOR U4800 ( .A(n4653), .B(n4654), .Z(n4704) );
  NANDN U4801 ( .A(n4628), .B(n4627), .Z(n4632) );
  NANDN U4802 ( .A(n4630), .B(n4629), .Z(n4631) );
  NAND U4803 ( .A(n4632), .B(n4631), .Z(n4701) );
  OR U4804 ( .A(n4634), .B(n4633), .Z(n4638) );
  NANDN U4805 ( .A(n4636), .B(n4635), .Z(n4637) );
  AND U4806 ( .A(n4638), .B(n4637), .Z(n4702) );
  XNOR U4807 ( .A(n4701), .B(n4702), .Z(n4703) );
  XNOR U4808 ( .A(n4704), .B(n4703), .Z(n4646) );
  NANDN U4809 ( .A(n4640), .B(n4639), .Z(n4644) );
  NAND U4810 ( .A(n4642), .B(n4641), .Z(n4643) );
  AND U4811 ( .A(n4644), .B(n4643), .Z(n4645) );
  XNOR U4812 ( .A(n4646), .B(n4645), .Z(n4647) );
  XNOR U4813 ( .A(n4648), .B(n4647), .Z(n4708) );
  XOR U4814 ( .A(n4709), .B(n4708), .Z(c[115]) );
  NANDN U4815 ( .A(n4646), .B(n4645), .Z(n4650) );
  NANDN U4816 ( .A(n4648), .B(n4647), .Z(n4649) );
  NAND U4817 ( .A(n4650), .B(n4649), .Z(n4716) );
  NANDN U4818 ( .A(n4652), .B(n4651), .Z(n4656) );
  NAND U4819 ( .A(n4654), .B(n4653), .Z(n4655) );
  NAND U4820 ( .A(n4656), .B(n4655), .Z(n4766) );
  NANDN U4821 ( .A(n4657), .B(n4987), .Z(n4659) );
  XNOR U4822 ( .A(n4909), .B(n4990), .Z(n4741) );
  OR U4823 ( .A(n4741), .B(n4986), .Z(n4658) );
  NAND U4824 ( .A(n4659), .B(n4658), .Z(n4727) );
  XNOR U4825 ( .A(n4992), .B(n4859), .Z(n4735) );
  OR U4826 ( .A(n4735), .B(n4860), .Z(n4662) );
  NAND U4827 ( .A(n4660), .B(n4915), .Z(n4661) );
  NAND U4828 ( .A(n4662), .B(n4661), .Z(n4725) );
  IV U4829 ( .A(a[62]), .Z(n5056) );
  XNOR U4830 ( .A(n5056), .B(n4744), .Z(n4747) );
  NANDN U4831 ( .A(n4747), .B(n4745), .Z(n4665) );
  NANDN U4832 ( .A(n4663), .B(n4746), .Z(n4664) );
  AND U4833 ( .A(n4665), .B(n4664), .Z(n4726) );
  XNOR U4834 ( .A(n4725), .B(n4726), .Z(n4728) );
  XOR U4835 ( .A(n4727), .B(n4728), .Z(n4722) );
  NAND U4836 ( .A(n5052), .B(n4666), .Z(n4668) );
  XOR U4837 ( .A(b[13]), .B(a[56]), .Z(n4738) );
  NANDN U4838 ( .A(n5041), .B(n4738), .Z(n4667) );
  NAND U4839 ( .A(n4668), .B(n4667), .Z(n4719) );
  NANDN U4840 ( .A(n4670), .B(n4669), .Z(n4671) );
  NANDN U4841 ( .A(n4750), .B(n4671), .Z(n4752) );
  ANDN U4842 ( .B(a[52]), .A(n210), .Z(n4787) );
  XOR U4843 ( .A(n4752), .B(n4787), .Z(n4753) );
  NAND U4844 ( .A(n5092), .B(n4672), .Z(n4674) );
  XOR U4845 ( .A(b[15]), .B(a[54]), .Z(n4732) );
  NANDN U4846 ( .A(n5095), .B(n4732), .Z(n4673) );
  AND U4847 ( .A(n4674), .B(n4673), .Z(n4754) );
  XOR U4848 ( .A(n4753), .B(n4754), .Z(n4720) );
  XOR U4849 ( .A(n4719), .B(n4720), .Z(n4721) );
  XOR U4850 ( .A(n4722), .B(n4721), .Z(n4757) );
  NANDN U4851 ( .A(n4680), .B(n4679), .Z(n4684) );
  NANDN U4852 ( .A(n4682), .B(n4681), .Z(n4683) );
  NAND U4853 ( .A(n4684), .B(n4683), .Z(n4760) );
  NAND U4854 ( .A(n4686), .B(n4685), .Z(n4690) );
  OR U4855 ( .A(n4688), .B(n4687), .Z(n4689) );
  NAND U4856 ( .A(n4690), .B(n4689), .Z(n4759) );
  XOR U4857 ( .A(n4760), .B(n4759), .Z(n4762) );
  XOR U4858 ( .A(n4762), .B(n4761), .Z(n4756) );
  XOR U4859 ( .A(n4755), .B(n4756), .Z(n4758) );
  XNOR U4860 ( .A(n4757), .B(n4758), .Z(n4763) );
  NANDN U4861 ( .A(n4696), .B(n4695), .Z(n4700) );
  NANDN U4862 ( .A(n4698), .B(n4697), .Z(n4699) );
  NAND U4863 ( .A(n4700), .B(n4699), .Z(n4764) );
  XOR U4864 ( .A(n4763), .B(n4764), .Z(n4765) );
  XNOR U4865 ( .A(n4766), .B(n4765), .Z(n4714) );
  IV U4866 ( .A(n4714), .Z(n4712) );
  NANDN U4867 ( .A(n4702), .B(n4701), .Z(n4706) );
  NAND U4868 ( .A(n4704), .B(n4703), .Z(n4705) );
  AND U4869 ( .A(n4706), .B(n4705), .Z(n4713) );
  XNOR U4870 ( .A(n4712), .B(n4713), .Z(n4707) );
  XNOR U4871 ( .A(n4716), .B(n4707), .Z(n4711) );
  OR U4872 ( .A(n4709), .B(n4708), .Z(n4710) );
  XOR U4873 ( .A(n4711), .B(n4710), .Z(c[116]) );
  OR U4874 ( .A(n4711), .B(n4710), .Z(n4828) );
  NAND U4875 ( .A(n4712), .B(n4713), .Z(n4718) );
  ANDN U4876 ( .B(n4714), .A(n4713), .Z(n4715) );
  OR U4877 ( .A(n4716), .B(n4715), .Z(n4717) );
  NAND U4878 ( .A(n4718), .B(n4717), .Z(n4772) );
  OR U4879 ( .A(n4720), .B(n4719), .Z(n4724) );
  NANDN U4880 ( .A(n4722), .B(n4721), .Z(n4723) );
  NAND U4881 ( .A(n4724), .B(n4723), .Z(n4782) );
  NANDN U4882 ( .A(n4726), .B(n4725), .Z(n4730) );
  NAND U4883 ( .A(n4728), .B(n4727), .Z(n4729) );
  NAND U4884 ( .A(n4730), .B(n4729), .Z(n4822) );
  XNOR U4885 ( .A(b[15]), .B(n4731), .Z(n4817) );
  NANDN U4886 ( .A(n5095), .B(n4817), .Z(n4734) );
  NAND U4887 ( .A(n4732), .B(n5092), .Z(n4733) );
  NAND U4888 ( .A(n4734), .B(n4733), .Z(n4800) );
  XNOR U4889 ( .A(n5037), .B(n4859), .Z(n4809) );
  OR U4890 ( .A(n4809), .B(n4860), .Z(n4737) );
  NANDN U4891 ( .A(n4735), .B(n4915), .Z(n4736) );
  NAND U4892 ( .A(n4737), .B(n4736), .Z(n4797) );
  XNOR U4893 ( .A(n5129), .B(n4852), .Z(n4803) );
  OR U4894 ( .A(n4803), .B(n5041), .Z(n4740) );
  NAND U4895 ( .A(n4738), .B(n5052), .Z(n4739) );
  AND U4896 ( .A(n4740), .B(n4739), .Z(n4798) );
  XNOR U4897 ( .A(n4797), .B(n4798), .Z(n4799) );
  XNOR U4898 ( .A(n4800), .B(n4799), .Z(n4820) );
  NANDN U4899 ( .A(n4741), .B(n4987), .Z(n4743) );
  XNOR U4900 ( .A(n4909), .B(n4952), .Z(n4806) );
  OR U4901 ( .A(n4806), .B(n4986), .Z(n4742) );
  NAND U4902 ( .A(n4743), .B(n4742), .Z(n4791) );
  XNOR U4903 ( .A(n5094), .B(n4744), .Z(n4813) );
  NANDN U4904 ( .A(n4813), .B(n4745), .Z(n4749) );
  NANDN U4905 ( .A(n4747), .B(n4746), .Z(n4748) );
  AND U4906 ( .A(n4749), .B(n4748), .Z(n4792) );
  XOR U4907 ( .A(n4791), .B(n4792), .Z(n4794) );
  OR U4908 ( .A(n4751), .B(n4750), .Z(n4786) );
  NAND U4909 ( .A(b[15]), .B(a[53]), .Z(n4785) );
  XNOR U4910 ( .A(n4786), .B(n4785), .Z(n4788) );
  XOR U4911 ( .A(n4787), .B(n4788), .Z(n4793) );
  XOR U4912 ( .A(n4794), .B(n4793), .Z(n4821) );
  XOR U4913 ( .A(n4820), .B(n4821), .Z(n4823) );
  XNOR U4914 ( .A(n4822), .B(n4823), .Z(n4779) );
  XNOR U4915 ( .A(n4779), .B(n4780), .Z(n4781) );
  XOR U4916 ( .A(n4782), .B(n4781), .Z(n4777) );
  XNOR U4917 ( .A(n4776), .B(n4775), .Z(n4778) );
  XNOR U4918 ( .A(n4777), .B(n4778), .Z(n4769) );
  OR U4919 ( .A(n4764), .B(n4763), .Z(n4768) );
  NAND U4920 ( .A(n4766), .B(n4765), .Z(n4767) );
  NAND U4921 ( .A(n4768), .B(n4767), .Z(n4770) );
  XOR U4922 ( .A(n4769), .B(n4770), .Z(n4771) );
  XNOR U4923 ( .A(n4772), .B(n4771), .Z(n4827) );
  XOR U4924 ( .A(n4828), .B(n4827), .Z(c[117]) );
  OR U4925 ( .A(n4770), .B(n4769), .Z(n4774) );
  NANDN U4926 ( .A(n4772), .B(n4771), .Z(n4773) );
  AND U4927 ( .A(n4774), .B(n4773), .Z(n4833) );
  NANDN U4928 ( .A(n4780), .B(n4779), .Z(n4784) );
  NANDN U4929 ( .A(n4782), .B(n4781), .Z(n4783) );
  NAND U4930 ( .A(n4784), .B(n4783), .Z(n4837) );
  OR U4931 ( .A(n4786), .B(n4785), .Z(n4790) );
  NANDN U4932 ( .A(n4788), .B(n4787), .Z(n4789) );
  NAND U4933 ( .A(n4790), .B(n4789), .Z(n4848) );
  NANDN U4934 ( .A(n4792), .B(n4791), .Z(n4796) );
  OR U4935 ( .A(n4794), .B(n4793), .Z(n4795) );
  NAND U4936 ( .A(n4796), .B(n4795), .Z(n4847) );
  NANDN U4937 ( .A(n4798), .B(n4797), .Z(n4802) );
  NAND U4938 ( .A(n4800), .B(n4799), .Z(n4801) );
  NAND U4939 ( .A(n4802), .B(n4801), .Z(n4842) );
  XNOR U4940 ( .A(n5129), .B(n4990), .Z(n4864) );
  OR U4941 ( .A(n4864), .B(n5041), .Z(n4805) );
  NANDN U4942 ( .A(n4803), .B(n5052), .Z(n4804) );
  NAND U4943 ( .A(n4805), .B(n4804), .Z(n4875) );
  NANDN U4944 ( .A(n4806), .B(n4987), .Z(n4808) );
  XNOR U4945 ( .A(n4909), .B(n4992), .Z(n4856) );
  OR U4946 ( .A(n4856), .B(n4986), .Z(n4807) );
  NAND U4947 ( .A(n4808), .B(n4807), .Z(n4872) );
  XNOR U4948 ( .A(n5056), .B(n4859), .Z(n4861) );
  OR U4949 ( .A(n4861), .B(n4860), .Z(n4811) );
  NANDN U4950 ( .A(n4809), .B(n4915), .Z(n4810) );
  AND U4951 ( .A(n4811), .B(n4810), .Z(n4873) );
  XOR U4952 ( .A(n4872), .B(n4873), .Z(n4874) );
  XOR U4953 ( .A(n4875), .B(n4874), .Z(n4840) );
  XNOR U4954 ( .A(b[7]), .B(n4812), .Z(n4816) );
  XNOR U4955 ( .A(b[6]), .B(b[5]), .Z(n4814) );
  NAND U4956 ( .A(n4814), .B(n4813), .Z(n4815) );
  AND U4957 ( .A(n4816), .B(n4815), .Z(n4867) );
  ANDN U4958 ( .B(a[54]), .A(n210), .Z(n4902) );
  XNOR U4959 ( .A(n4867), .B(n4902), .Z(n4868) );
  NAND U4960 ( .A(n5092), .B(n4817), .Z(n4819) );
  XOR U4961 ( .A(b[15]), .B(a[56]), .Z(n4853) );
  NANDN U4962 ( .A(n5095), .B(n4853), .Z(n4818) );
  AND U4963 ( .A(n4819), .B(n4818), .Z(n4869) );
  XNOR U4964 ( .A(n4868), .B(n4869), .Z(n4841) );
  XOR U4965 ( .A(n4840), .B(n4841), .Z(n4843) );
  XOR U4966 ( .A(n4842), .B(n4843), .Z(n4846) );
  XOR U4967 ( .A(n4847), .B(n4846), .Z(n4849) );
  XNOR U4968 ( .A(n4848), .B(n4849), .Z(n4834) );
  NANDN U4969 ( .A(n4821), .B(n4820), .Z(n4825) );
  OR U4970 ( .A(n4823), .B(n4822), .Z(n4824) );
  NAND U4971 ( .A(n4825), .B(n4824), .Z(n4835) );
  XNOR U4972 ( .A(n4834), .B(n4835), .Z(n4836) );
  XOR U4973 ( .A(n4837), .B(n4836), .Z(n4831) );
  XNOR U4974 ( .A(n4832), .B(n4831), .Z(n4826) );
  XOR U4975 ( .A(n4833), .B(n4826), .Z(n4829) );
  OR U4976 ( .A(n4828), .B(n4827), .Z(n4830) );
  XNOR U4977 ( .A(n4829), .B(n4830), .Z(c[118]) );
  NANDN U4978 ( .A(n4830), .B(n4829), .Z(n4877) );
  NANDN U4979 ( .A(n4835), .B(n4834), .Z(n4839) );
  NAND U4980 ( .A(n4837), .B(n4836), .Z(n4838) );
  NAND U4981 ( .A(n4839), .B(n4838), .Z(n4879) );
  NANDN U4982 ( .A(n4841), .B(n4840), .Z(n4845) );
  OR U4983 ( .A(n4843), .B(n4842), .Z(n4844) );
  NAND U4984 ( .A(n4845), .B(n4844), .Z(n4884) );
  NANDN U4985 ( .A(n4847), .B(n4846), .Z(n4851) );
  OR U4986 ( .A(n4849), .B(n4848), .Z(n4850) );
  AND U4987 ( .A(n4851), .B(n4850), .Z(n4885) );
  XNOR U4988 ( .A(n4884), .B(n4885), .Z(n4886) );
  XNOR U4989 ( .A(n210), .B(n4852), .Z(n4918) );
  OR U4990 ( .A(n4918), .B(n5095), .Z(n4855) );
  NAND U4991 ( .A(n4853), .B(n5092), .Z(n4854) );
  NAND U4992 ( .A(n4855), .B(n4854), .Z(n4924) );
  NANDN U4993 ( .A(n4856), .B(n4987), .Z(n4858) );
  XNOR U4994 ( .A(n4909), .B(n5037), .Z(n4908) );
  OR U4995 ( .A(n4908), .B(n4986), .Z(n4857) );
  NAND U4996 ( .A(n4858), .B(n4857), .Z(n4921) );
  XNOR U4997 ( .A(n5094), .B(n4859), .Z(n4916) );
  OR U4998 ( .A(n4916), .B(n4860), .Z(n4863) );
  NANDN U4999 ( .A(n4861), .B(n4915), .Z(n4862) );
  NAND U5000 ( .A(n4863), .B(n4862), .Z(n4896) );
  XNOR U5001 ( .A(n5129), .B(n4952), .Z(n4912) );
  OR U5002 ( .A(n4912), .B(n5041), .Z(n4866) );
  NANDN U5003 ( .A(n4864), .B(n5052), .Z(n4865) );
  AND U5004 ( .A(n4866), .B(n4865), .Z(n4897) );
  XNOR U5005 ( .A(n4896), .B(n4897), .Z(n4898) );
  XOR U5006 ( .A(n4903), .B(n4902), .Z(n4905) );
  NAND U5007 ( .A(a[55]), .B(b[15]), .Z(n4904) );
  XOR U5008 ( .A(n4905), .B(n4904), .Z(n4899) );
  XOR U5009 ( .A(n4898), .B(n4899), .Z(n4922) );
  XOR U5010 ( .A(n4921), .B(n4922), .Z(n4923) );
  XNOR U5011 ( .A(n4924), .B(n4923), .Z(n4893) );
  NANDN U5012 ( .A(n4867), .B(n4902), .Z(n4871) );
  NAND U5013 ( .A(n4869), .B(n4868), .Z(n4870) );
  NAND U5014 ( .A(n4871), .B(n4870), .Z(n4890) );
  XNOR U5015 ( .A(n4890), .B(n4891), .Z(n4892) );
  XOR U5016 ( .A(n4893), .B(n4892), .Z(n4887) );
  XOR U5017 ( .A(n4886), .B(n4887), .Z(n4878) );
  XOR U5018 ( .A(n4879), .B(n4878), .Z(n4881) );
  XOR U5019 ( .A(n4880), .B(n4881), .Z(n4876) );
  XOR U5020 ( .A(n4877), .B(n4876), .Z(c[119]) );
  OR U5021 ( .A(n4877), .B(n4876), .Z(n4968) );
  NANDN U5022 ( .A(n4879), .B(n4878), .Z(n4883) );
  OR U5023 ( .A(n4881), .B(n4880), .Z(n4882) );
  NAND U5024 ( .A(n4883), .B(n4882), .Z(n4934) );
  NANDN U5025 ( .A(n4885), .B(n4884), .Z(n4889) );
  NAND U5026 ( .A(n4887), .B(n4886), .Z(n4888) );
  NAND U5027 ( .A(n4889), .B(n4888), .Z(n4931) );
  NANDN U5028 ( .A(n4891), .B(n4890), .Z(n4895) );
  NAND U5029 ( .A(n4893), .B(n4892), .Z(n4894) );
  NAND U5030 ( .A(n4895), .B(n4894), .Z(n4930) );
  NANDN U5031 ( .A(n4897), .B(n4896), .Z(n4901) );
  NAND U5032 ( .A(n4899), .B(n4898), .Z(n4900) );
  NAND U5033 ( .A(n4901), .B(n4900), .Z(n4937) );
  NANDN U5034 ( .A(n4903), .B(n4902), .Z(n4907) );
  OR U5035 ( .A(n4905), .B(n4904), .Z(n4906) );
  NAND U5036 ( .A(n4907), .B(n4906), .Z(n4946) );
  NANDN U5037 ( .A(n4908), .B(n4987), .Z(n4911) );
  XNOR U5038 ( .A(n5056), .B(n4909), .Z(n4958) );
  OR U5039 ( .A(n4958), .B(n4986), .Z(n4910) );
  NAND U5040 ( .A(n4911), .B(n4910), .Z(n4943) );
  XNOR U5041 ( .A(b[13]), .B(n4992), .Z(n4949) );
  NANDN U5042 ( .A(n5041), .B(n4949), .Z(n4914) );
  NANDN U5043 ( .A(n4912), .B(n5052), .Z(n4913) );
  AND U5044 ( .A(n4914), .B(n4913), .Z(n4944) );
  XNOR U5045 ( .A(n4943), .B(n4944), .Z(n4945) );
  XNOR U5046 ( .A(n4946), .B(n4945), .Z(n4938) );
  XNOR U5047 ( .A(n4937), .B(n4938), .Z(n4939) );
  NANDN U5048 ( .A(n4916), .B(n4915), .Z(n4917) );
  ANDN U5049 ( .B(n4917), .A(n4956), .Z(n4963) );
  ANDN U5050 ( .B(a[56]), .A(n210), .Z(n4982) );
  XNOR U5051 ( .A(n210), .B(n4990), .Z(n4953) );
  OR U5052 ( .A(n4953), .B(n5095), .Z(n4920) );
  NANDN U5053 ( .A(n4918), .B(n5092), .Z(n4919) );
  AND U5054 ( .A(n4920), .B(n4919), .Z(n4961) );
  XOR U5055 ( .A(n4982), .B(n4961), .Z(n4962) );
  XNOR U5056 ( .A(n4963), .B(n4962), .Z(n4940) );
  XOR U5057 ( .A(n4939), .B(n4940), .Z(n4927) );
  NAND U5058 ( .A(n4922), .B(n4921), .Z(n4926) );
  NAND U5059 ( .A(n4924), .B(n4923), .Z(n4925) );
  NAND U5060 ( .A(n4926), .B(n4925), .Z(n4928) );
  XOR U5061 ( .A(n4927), .B(n4928), .Z(n4929) );
  XNOR U5062 ( .A(n4930), .B(n4929), .Z(n4932) );
  XNOR U5063 ( .A(n4931), .B(n4932), .Z(n4933) );
  XOR U5064 ( .A(n4934), .B(n4933), .Z(n4967) );
  XOR U5065 ( .A(n4968), .B(n4967), .Z(c[120]) );
  NANDN U5066 ( .A(n4932), .B(n4931), .Z(n4936) );
  NAND U5067 ( .A(n4934), .B(n4933), .Z(n4935) );
  NAND U5068 ( .A(n4936), .B(n4935), .Z(n4973) );
  NANDN U5069 ( .A(n4938), .B(n4937), .Z(n4942) );
  NAND U5070 ( .A(n4940), .B(n4939), .Z(n4941) );
  NAND U5071 ( .A(n4942), .B(n4941), .Z(n5007) );
  NANDN U5072 ( .A(n4944), .B(n4943), .Z(n4948) );
  NAND U5073 ( .A(n4946), .B(n4945), .Z(n4947) );
  NAND U5074 ( .A(n4948), .B(n4947), .Z(n5004) );
  NAND U5075 ( .A(n5052), .B(n4949), .Z(n4951) );
  XNOR U5076 ( .A(b[13]), .B(n5037), .Z(n4995) );
  NANDN U5077 ( .A(n5041), .B(n4995), .Z(n4950) );
  AND U5078 ( .A(n4951), .B(n4950), .Z(n4974) );
  XNOR U5079 ( .A(b[15]), .B(n4952), .Z(n4991) );
  NANDN U5080 ( .A(n5095), .B(n4991), .Z(n4955) );
  NANDN U5081 ( .A(n4953), .B(n5092), .Z(n4954) );
  AND U5082 ( .A(n4955), .B(n4954), .Z(n4975) );
  XOR U5083 ( .A(n4974), .B(n4975), .Z(n4976) );
  OR U5084 ( .A(n4957), .B(n4956), .Z(n4981) );
  NAND U5085 ( .A(a[57]), .B(b[15]), .Z(n4980) );
  XOR U5086 ( .A(n4981), .B(n4980), .Z(n4983) );
  XNOR U5087 ( .A(n4982), .B(n4983), .Z(n4977) );
  XNOR U5088 ( .A(n4976), .B(n4977), .Z(n5001) );
  NANDN U5089 ( .A(n4958), .B(n4987), .Z(n4960) );
  XNOR U5090 ( .A(b[11]), .B(a[63]), .Z(n4988) );
  OR U5091 ( .A(n4988), .B(n4986), .Z(n4959) );
  NAND U5092 ( .A(n4960), .B(n4959), .Z(n4999) );
  OR U5093 ( .A(n4982), .B(n4961), .Z(n4965) );
  NANDN U5094 ( .A(n4963), .B(n4962), .Z(n4964) );
  AND U5095 ( .A(n4965), .B(n4964), .Z(n4998) );
  XNOR U5096 ( .A(n4999), .B(n4998), .Z(n5000) );
  XNOR U5097 ( .A(n5001), .B(n5000), .Z(n5005) );
  XNOR U5098 ( .A(n5004), .B(n5005), .Z(n5006) );
  XOR U5099 ( .A(n5007), .B(n5006), .Z(n4972) );
  XNOR U5100 ( .A(n4973), .B(n4972), .Z(n4966) );
  XOR U5101 ( .A(n4971), .B(n4966), .Z(n4969) );
  OR U5102 ( .A(n4968), .B(n4967), .Z(n4970) );
  XNOR U5103 ( .A(n4969), .B(n4970), .Z(c[121]) );
  NANDN U5104 ( .A(n4970), .B(n4969), .Z(n5011) );
  OR U5105 ( .A(n4975), .B(n4974), .Z(n4979) );
  NANDN U5106 ( .A(n4977), .B(n4976), .Z(n4978) );
  NAND U5107 ( .A(n4979), .B(n4978), .Z(n5021) );
  OR U5108 ( .A(n4981), .B(n4980), .Z(n4985) );
  NAND U5109 ( .A(n4983), .B(n4982), .Z(n4984) );
  NAND U5110 ( .A(n4985), .B(n4984), .Z(n5024) );
  NANDN U5111 ( .A(n4986), .B(b[11]), .Z(n5034) );
  NANDN U5112 ( .A(n4988), .B(n4987), .Z(n4989) );
  NAND U5113 ( .A(n5034), .B(n4989), .Z(n5030) );
  NOR U5114 ( .A(n4990), .B(n210), .Z(n5062) );
  XOR U5115 ( .A(n5030), .B(n5062), .Z(n5031) );
  NAND U5116 ( .A(n5092), .B(n4991), .Z(n4994) );
  XNOR U5117 ( .A(b[15]), .B(n4992), .Z(n5036) );
  NANDN U5118 ( .A(n5095), .B(n5036), .Z(n4993) );
  AND U5119 ( .A(n4994), .B(n4993), .Z(n5032) );
  XOR U5120 ( .A(n5031), .B(n5032), .Z(n5025) );
  XOR U5121 ( .A(n5024), .B(n5025), .Z(n5026) );
  NAND U5122 ( .A(n5052), .B(n4995), .Z(n4997) );
  XNOR U5123 ( .A(a[62]), .B(n5129), .Z(n5040) );
  NANDN U5124 ( .A(n5041), .B(n5040), .Z(n4996) );
  NAND U5125 ( .A(n4997), .B(n4996), .Z(n5027) );
  XOR U5126 ( .A(n5026), .B(n5027), .Z(n5018) );
  NANDN U5127 ( .A(n4999), .B(n4998), .Z(n5003) );
  NANDN U5128 ( .A(n5001), .B(n5000), .Z(n5002) );
  NAND U5129 ( .A(n5003), .B(n5002), .Z(n5019) );
  XNOR U5130 ( .A(n5018), .B(n5019), .Z(n5020) );
  XNOR U5131 ( .A(n5021), .B(n5020), .Z(n5012) );
  NANDN U5132 ( .A(n5005), .B(n5004), .Z(n5009) );
  NAND U5133 ( .A(n5007), .B(n5006), .Z(n5008) );
  NAND U5134 ( .A(n5009), .B(n5008), .Z(n5013) );
  XOR U5135 ( .A(n5012), .B(n5013), .Z(n5015) );
  XOR U5136 ( .A(n5014), .B(n5015), .Z(n5010) );
  XOR U5137 ( .A(n5011), .B(n5010), .Z(c[122]) );
  OR U5138 ( .A(n5011), .B(n5010), .Z(n5045) );
  NANDN U5139 ( .A(n5013), .B(n5012), .Z(n5017) );
  OR U5140 ( .A(n5015), .B(n5014), .Z(n5016) );
  NAND U5141 ( .A(n5017), .B(n5016), .Z(n5049) );
  NANDN U5142 ( .A(n5019), .B(n5018), .Z(n5023) );
  NAND U5143 ( .A(n5021), .B(n5020), .Z(n5022) );
  NAND U5144 ( .A(n5023), .B(n5022), .Z(n5047) );
  OR U5145 ( .A(n5025), .B(n5024), .Z(n5029) );
  NANDN U5146 ( .A(n5027), .B(n5026), .Z(n5028) );
  NAND U5147 ( .A(n5029), .B(n5028), .Z(n5074) );
  NAND U5148 ( .A(n5033), .B(b[11]), .Z(n5035) );
  NAND U5149 ( .A(n5035), .B(n5034), .Z(n5060) );
  NAND U5150 ( .A(a[59]), .B(b[15]), .Z(n5059) );
  XOR U5151 ( .A(n5060), .B(n5059), .Z(n5061) );
  NAND U5152 ( .A(n5092), .B(n5036), .Z(n5039) );
  XNOR U5153 ( .A(b[15]), .B(n5037), .Z(n5055) );
  NANDN U5154 ( .A(n5095), .B(n5055), .Z(n5038) );
  NAND U5155 ( .A(n5039), .B(n5038), .Z(n5065) );
  XOR U5156 ( .A(n5066), .B(n5065), .Z(n5067) );
  NAND U5157 ( .A(n5052), .B(n5040), .Z(n5043) );
  XNOR U5158 ( .A(n5129), .B(n5094), .Z(n5053) );
  OR U5159 ( .A(n5053), .B(n5041), .Z(n5042) );
  AND U5160 ( .A(n5043), .B(n5042), .Z(n5068) );
  XNOR U5161 ( .A(n5067), .B(n5068), .Z(n5072) );
  XNOR U5162 ( .A(n5071), .B(n5072), .Z(n5073) );
  XOR U5163 ( .A(n5074), .B(n5073), .Z(n5046) );
  XNOR U5164 ( .A(n5047), .B(n5046), .Z(n5048) );
  XOR U5165 ( .A(n5049), .B(n5048), .Z(n5044) );
  XOR U5166 ( .A(n5045), .B(n5044), .Z(c[123]) );
  OR U5167 ( .A(n5045), .B(n5044), .Z(n5078) );
  NANDN U5168 ( .A(n5047), .B(n5046), .Z(n5051) );
  NAND U5169 ( .A(n5049), .B(n5048), .Z(n5050) );
  NAND U5170 ( .A(n5051), .B(n5050), .Z(n5082) );
  NANDN U5171 ( .A(n5053), .B(n5052), .Z(n5054) );
  NANDN U5172 ( .A(n5086), .B(n5054), .Z(n5087) );
  ANDN U5173 ( .B(a[60]), .A(n210), .Z(n5114) );
  XNOR U5174 ( .A(n5087), .B(n5114), .Z(n5088) );
  NAND U5175 ( .A(n5092), .B(n5055), .Z(n5058) );
  XNOR U5176 ( .A(n210), .B(n5056), .Z(n5093) );
  OR U5177 ( .A(n5093), .B(n5095), .Z(n5057) );
  NAND U5178 ( .A(n5058), .B(n5057), .Z(n5089) );
  XOR U5179 ( .A(n5088), .B(n5089), .Z(n5098) );
  OR U5180 ( .A(n5060), .B(n5059), .Z(n5064) );
  NAND U5181 ( .A(n5062), .B(n5061), .Z(n5063) );
  AND U5182 ( .A(n5064), .B(n5063), .Z(n5099) );
  XNOR U5183 ( .A(n5098), .B(n5099), .Z(n5100) );
  OR U5184 ( .A(n5066), .B(n5065), .Z(n5070) );
  NAND U5185 ( .A(n5068), .B(n5067), .Z(n5069) );
  NAND U5186 ( .A(n5070), .B(n5069), .Z(n5101) );
  XOR U5187 ( .A(n5100), .B(n5101), .Z(n5079) );
  NANDN U5188 ( .A(n5072), .B(n5071), .Z(n5076) );
  NAND U5189 ( .A(n5074), .B(n5073), .Z(n5075) );
  AND U5190 ( .A(n5076), .B(n5075), .Z(n5080) );
  XNOR U5191 ( .A(n5079), .B(n5080), .Z(n5081) );
  XOR U5192 ( .A(n5082), .B(n5081), .Z(n5077) );
  XOR U5193 ( .A(n5078), .B(n5077), .Z(c[124]) );
  OR U5194 ( .A(n5078), .B(n5077), .Z(n5105) );
  NANDN U5195 ( .A(n5080), .B(n5079), .Z(n5084) );
  NAND U5196 ( .A(n5082), .B(n5081), .Z(n5083) );
  NAND U5197 ( .A(n5084), .B(n5083), .Z(n5120) );
  OR U5198 ( .A(n5086), .B(n5085), .Z(n5112) );
  AND U5199 ( .A(b[15]), .B(a[61]), .Z(n5111) );
  XNOR U5200 ( .A(n5112), .B(n5111), .Z(n5113) );
  XOR U5201 ( .A(n5114), .B(n5113), .Z(n5126) );
  NANDN U5202 ( .A(n5087), .B(n5114), .Z(n5091) );
  NANDN U5203 ( .A(n5089), .B(n5088), .Z(n5090) );
  AND U5204 ( .A(n5091), .B(n5090), .Z(n5123) );
  NANDN U5205 ( .A(n5093), .B(n5092), .Z(n5097) );
  XNOR U5206 ( .A(n210), .B(n5094), .Z(n5107) );
  OR U5207 ( .A(n5107), .B(n5095), .Z(n5096) );
  NAND U5208 ( .A(n5097), .B(n5096), .Z(n5124) );
  XOR U5209 ( .A(n5123), .B(n5124), .Z(n5125) );
  XOR U5210 ( .A(n5126), .B(n5125), .Z(n5118) );
  NANDN U5211 ( .A(n5099), .B(n5098), .Z(n5103) );
  NANDN U5212 ( .A(n5101), .B(n5100), .Z(n5102) );
  AND U5213 ( .A(n5103), .B(n5102), .Z(n5117) );
  XNOR U5214 ( .A(n5118), .B(n5117), .Z(n5119) );
  XOR U5215 ( .A(n5120), .B(n5119), .Z(n5104) );
  XOR U5216 ( .A(n5105), .B(n5104), .Z(c[125]) );
  OR U5217 ( .A(n5105), .B(n5104), .Z(n5141) );
  NAND U5218 ( .A(b[13]), .B(b[14]), .Z(n5106) );
  XNOR U5219 ( .A(b[15]), .B(n5106), .Z(n5110) );
  XNOR U5220 ( .A(b[14]), .B(b[13]), .Z(n5108) );
  NAND U5221 ( .A(n5108), .B(n5107), .Z(n5109) );
  AND U5222 ( .A(n5110), .B(n5109), .Z(n5147) );
  NAND U5223 ( .A(b[15]), .B(a[62]), .Z(n5149) );
  NANDN U5224 ( .A(n5112), .B(n5111), .Z(n5116) );
  NAND U5225 ( .A(n5114), .B(n5113), .Z(n5115) );
  AND U5226 ( .A(n5116), .B(n5115), .Z(n5148) );
  XNOR U5227 ( .A(n5149), .B(n5148), .Z(n5146) );
  XNOR U5228 ( .A(n5147), .B(n5146), .Z(n5136) );
  NANDN U5229 ( .A(n5118), .B(n5117), .Z(n5122) );
  NAND U5230 ( .A(n5120), .B(n5119), .Z(n5121) );
  NAND U5231 ( .A(n5122), .B(n5121), .Z(n5135) );
  OR U5232 ( .A(n5124), .B(n5123), .Z(n5128) );
  NANDN U5233 ( .A(n5126), .B(n5125), .Z(n5127) );
  NAND U5234 ( .A(n5128), .B(n5127), .Z(n5134) );
  XOR U5235 ( .A(n5135), .B(n5134), .Z(n5137) );
  XOR U5236 ( .A(n5136), .B(n5137), .Z(n5140) );
  XOR U5237 ( .A(n5141), .B(n5140), .Z(c[126]) );
  NAND U5238 ( .A(n5129), .B(n210), .Z(n5130) );
  AND U5239 ( .A(n5130), .B(a[63]), .Z(n5133) );
  NANDN U5240 ( .A(b[14]), .B(n5131), .Z(n5132) );
  NAND U5241 ( .A(n5133), .B(n5132), .Z(n5145) );
  AND U5242 ( .A(n5135), .B(n5134), .Z(n5139) );
  AND U5243 ( .A(n5137), .B(n5136), .Z(n5138) );
  OR U5244 ( .A(n5139), .B(n5138), .Z(n5143) );
  OR U5245 ( .A(n5141), .B(n5140), .Z(n5142) );
  NAND U5246 ( .A(n5143), .B(n5142), .Z(n5144) );
  XNOR U5247 ( .A(n5145), .B(n5144), .Z(n5153) );
  OR U5248 ( .A(n5147), .B(n5146), .Z(n5151) );
  OR U5249 ( .A(n5149), .B(n5148), .Z(n5150) );
  NAND U5250 ( .A(n5151), .B(n5150), .Z(n5152) );
  XNOR U5251 ( .A(n5153), .B(n5152), .Z(c[127]) );
endmodule

