
module mult_N64_CC1 ( clk, rst, a, b, c );
  input [63:0] a;
  input [63:0] b;
  output [63:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375;

  XOR U1 ( .A(n6352), .B(n6583), .Z(n6356) );
  XOR U2 ( .A(n6125), .B(n6335), .Z(n6126) );
  XOR U3 ( .A(n5880), .B(n6082), .Z(n5884) );
  XOR U4 ( .A(n5370), .B(n5559), .Z(n5374) );
  XOR U5 ( .A(n4815), .B(n5020), .Z(n4816) );
  XOR U6 ( .A(n4207), .B(n4462), .Z(n4208) );
  XOR U7 ( .A(n3939), .B(n4161), .Z(n3940) );
  XOR U8 ( .A(n4561), .B(n4732), .Z(n4565) );
  XOR U9 ( .A(n3297), .B(n3567), .Z(n3298) );
  XOR U10 ( .A(n3997), .B(n4147), .Z(n3998) );
  XOR U11 ( .A(n1657), .B(n1958), .Z(n1658) );
  XOR U12 ( .A(n3413), .B(n3539), .Z(n3414) );
  XOR U13 ( .A(n4023), .B(n4142), .Z(n4018) );
  XOR U14 ( .A(n3127), .B(n3223), .Z(n3128) );
  XOR U15 ( .A(n1829), .B(n1916), .Z(n1833) );
  XOR U16 ( .A(n1844), .B(n1913), .Z(n1848) );
  XOR U17 ( .A(n11293), .B(n11319), .Z(n11297) );
  XOR U18 ( .A(n6600), .B(n6819), .Z(n6604) );
  XOR U19 ( .A(n6371), .B(n6580), .Z(n6366) );
  XOR U20 ( .A(n5851), .B(n6090), .Z(n5855) );
  XOR U21 ( .A(n5875), .B(n6083), .Z(n5879) );
  XOR U22 ( .A(n5066), .B(n5300), .Z(n5067) );
  XOR U23 ( .A(n5049), .B(n5304), .Z(n5053) );
  XOR U24 ( .A(n6142), .B(n6331), .Z(n6150) );
  XOR U25 ( .A(n5897), .B(n6078), .Z(n5898) );
  XOR U26 ( .A(n5078), .B(n5297), .Z(n5082) );
  XOR U27 ( .A(n4817), .B(n5019), .Z(n4821) );
  XOR U28 ( .A(n3910), .B(n4168), .Z(n3911) );
  XOR U29 ( .A(n4190), .B(n4466), .Z(n4194) );
  XOR U30 ( .A(n4236), .B(n4455), .Z(n4237) );
  XOR U31 ( .A(n5385), .B(n5556), .Z(n5393) );
  XOR U32 ( .A(n8695), .B(n8860), .Z(n8699) );
  XOR U33 ( .A(n8334), .B(n8495), .Z(n8342) );
  XOR U34 ( .A(n4265), .B(n4448), .Z(n4266) );
  XOR U35 ( .A(n4219), .B(n4459), .Z(n4223) );
  XOR U36 ( .A(n3280), .B(n3571), .Z(n3284) );
  XOR U37 ( .A(n3326), .B(n3560), .Z(n3327) );
  XOR U38 ( .A(n3304), .B(n3565), .Z(n3308) );
  XOR U39 ( .A(n3951), .B(n4158), .Z(n3955) );
  XOR U40 ( .A(n7760), .B(n7907), .Z(n7768) );
  XOR U41 ( .A(n3355), .B(n3553), .Z(n3356) );
  XOR U42 ( .A(n4870), .B(n5007), .Z(n4865) );
  XOR U43 ( .A(n3980), .B(n4151), .Z(n3984) );
  XOR U44 ( .A(n2332), .B(n2619), .Z(n2336) );
  XOR U45 ( .A(n2313), .B(n2625), .Z(n2317) );
  XOR U46 ( .A(n2359), .B(n2613), .Z(n2360) );
  XOR U47 ( .A(n4004), .B(n4145), .Z(n4008) );
  XOR U48 ( .A(n3384), .B(n3546), .Z(n3385) );
  XOR U49 ( .A(n8894), .B(n9028), .Z(n8895) );
  XOR U50 ( .A(n3023), .B(n3248), .Z(n3027) );
  XOR U51 ( .A(n9229), .B(n9354), .Z(n9224) );
  XOR U52 ( .A(n8724), .B(n8853), .Z(n8728) );
  XOR U53 ( .A(n8363), .B(n8488), .Z(n8371) );
  XOR U54 ( .A(n7566), .B(n7695), .Z(n7570) );
  XOR U55 ( .A(n7133), .B(n7258), .Z(n7141) );
  XOR U56 ( .A(n2388), .B(n2606), .Z(n2389) );
  XOR U57 ( .A(n1312), .B(n1618), .Z(n1313) );
  XOR U58 ( .A(n3415), .B(n3538), .Z(n3419) );
  XOR U59 ( .A(n3052), .B(n3241), .Z(n3056) );
  XOR U60 ( .A(n1295), .B(n1622), .Z(n1299) );
  XOR U61 ( .A(n1341), .B(n1611), .Z(n1342) );
  XOR U62 ( .A(n2417), .B(n2599), .Z(n2418) );
  XOR U63 ( .A(n4026), .B(n4140), .Z(n4027) );
  XOR U64 ( .A(n2038), .B(n2281), .Z(n2042) );
  XOR U65 ( .A(n3081), .B(n3234), .Z(n3085) );
  XOR U66 ( .A(n6919), .B(n7032), .Z(n6923) );
  XOR U67 ( .A(n2446), .B(n2592), .Z(n2447) );
  XOR U68 ( .A(n1370), .B(n1604), .Z(n1371) );
  XOR U69 ( .A(n9542), .B(n9650), .Z(n9546) );
  XOR U70 ( .A(n3110), .B(n3227), .Z(n3114) );
  XOR U71 ( .A(n2067), .B(n2274), .Z(n2071) );
  XOR U72 ( .A(n1399), .B(n1597), .Z(n1400) );
  XOR U73 ( .A(n7801), .B(n7897), .Z(n7802) );
  XOR U74 ( .A(n3739), .B(n3838), .Z(n3747) );
  XOR U75 ( .A(n2096), .B(n2267), .Z(n2100) );
  XOR U76 ( .A(n3442), .B(n3532), .Z(n3443) );
  XOR U77 ( .A(n1428), .B(n1590), .Z(n1429) );
  XOR U78 ( .A(n2482), .B(n2582), .Z(n2486) );
  XOR U79 ( .A(n9838), .B(n9925), .Z(n9842) );
  XOR U80 ( .A(n8930), .B(n9019), .Z(n8934) );
  XOR U81 ( .A(n2164), .B(n2251), .Z(n2168) );
  XOR U82 ( .A(n2125), .B(n2260), .Z(n2129) );
  XOR U83 ( .A(n1457), .B(n1583), .Z(n1458) );
  XOR U84 ( .A(n6943), .B(n7026), .Z(n6947) );
  XOR U85 ( .A(n4349), .B(n4429), .Z(n4344) );
  XOR U86 ( .A(n2822), .B(n2903), .Z(n2826) );
  XOR U87 ( .A(n6478), .B(n6553), .Z(n6486) );
  XOR U88 ( .A(n1131), .B(n1232), .Z(n1135) );
  XOR U89 ( .A(n10107), .B(n10176), .Z(n10111) );
  XOR U90 ( .A(n9273), .B(n9342), .Z(n9277) );
  XOR U91 ( .A(n8221), .B(n8290), .Z(n8225) );
  XOR U92 ( .A(n5986), .B(n6056), .Z(n5990) );
  XOR U93 ( .A(n1494), .B(n1575), .Z(n1498) );
  XOR U94 ( .A(n2837), .B(n2900), .Z(n2841) );
  XOR U95 ( .A(n1161), .B(n1226), .Z(n1165) );
  XOR U96 ( .A(n5739), .B(n5796), .Z(n5747) );
  XOR U97 ( .A(n5211), .B(n5265), .Z(n5212) );
  XOR U98 ( .A(n11033), .B(n11084), .Z(n11037) );
  XOR U99 ( .A(n10348), .B(n10404), .Z(n10356) );
  XOR U100 ( .A(n9586), .B(n9640), .Z(n9594) );
  XOR U101 ( .A(n8606), .B(n8660), .Z(n8614) );
  XOR U102 ( .A(n7421), .B(n7465), .Z(n7416) );
  XOR U103 ( .A(n1524), .B(n1569), .Z(n1528) );
  XOR U104 ( .A(n7847), .B(n7886), .Z(n7855) );
  XOR U105 ( .A(n7205), .B(n7240), .Z(n7209) );
  XOR U106 ( .A(n6745), .B(n6784), .Z(n6749) );
  XOR U107 ( .A(n11159), .B(n11200), .Z(n11163) );
  XOR U108 ( .A(n10578), .B(n10607), .Z(n10573) );
  XOR U109 ( .A(n9886), .B(n9915), .Z(n9881) );
  XOR U110 ( .A(n8978), .B(n9009), .Z(n8973) );
  XOR U111 ( .A(n1186), .B(n1221), .Z(n1190) );
  XOR U112 ( .A(n11260), .B(n11286), .Z(n11264) );
  XOR U113 ( .A(n5501), .B(n5528), .Z(n5505) );
  XOR U114 ( .A(n3798), .B(n3825), .Z(n3802) );
  XOR U115 ( .A(n7060), .B(n7275), .Z(n7064) );
  XOR U116 ( .A(n6108), .B(n6339), .Z(n6112) );
  XOR U117 ( .A(n5606), .B(n5829), .Z(n5607) );
  XOR U118 ( .A(n7508), .B(n7709), .Z(n7512) );
  XOR U119 ( .A(n7075), .B(n7272), .Z(n7083) );
  XOR U120 ( .A(n6617), .B(n6815), .Z(n6618) );
  XOR U121 ( .A(n6132), .B(n6333), .Z(n6136) );
  XOR U122 ( .A(n5322), .B(n5571), .Z(n5326) );
  XOR U123 ( .A(n4786), .B(n5027), .Z(n4787) );
  XOR U124 ( .A(n5095), .B(n5293), .Z(n5096) );
  XOR U125 ( .A(n5351), .B(n5564), .Z(n5355) );
  XOR U126 ( .A(n8319), .B(n8498), .Z(n8323) );
  XOR U127 ( .A(n7933), .B(n8116), .Z(n7937) );
  XOR U128 ( .A(n7527), .B(n7706), .Z(n7522) );
  XOR U129 ( .A(n7089), .B(n7268), .Z(n7093) );
  XOR U130 ( .A(n6629), .B(n6812), .Z(n6633) );
  XOR U131 ( .A(n6151), .B(n6330), .Z(n6146) );
  XOR U132 ( .A(n5637), .B(n5820), .Z(n5641) );
  XOR U133 ( .A(n4484), .B(n4751), .Z(n4488) );
  XOR U134 ( .A(n4822), .B(n5018), .Z(n4826) );
  XOR U135 ( .A(n4513), .B(n4744), .Z(n4517) );
  XOR U136 ( .A(n3912), .B(n4167), .Z(n3916) );
  XOR U137 ( .A(n4238), .B(n4454), .Z(n4242) );
  XOR U138 ( .A(n7950), .B(n8112), .Z(n7951) );
  XOR U139 ( .A(n7537), .B(n7702), .Z(n7541) );
  XOR U140 ( .A(n7104), .B(n7265), .Z(n7112) );
  XOR U141 ( .A(n6646), .B(n6808), .Z(n6647) );
  XOR U142 ( .A(n6161), .B(n6326), .Z(n6165) );
  XOR U143 ( .A(n5652), .B(n5817), .Z(n5660) );
  XOR U144 ( .A(n5124), .B(n5286), .Z(n5125) );
  XOR U145 ( .A(n3589), .B(n3875), .Z(n3593) );
  XOR U146 ( .A(n4566), .B(n4731), .Z(n4570) );
  XOR U147 ( .A(n3968), .B(n4154), .Z(n3969) );
  XOR U148 ( .A(n2982), .B(n3258), .Z(n2983) );
  XOR U149 ( .A(n4547), .B(n4736), .Z(n4555) );
  XOR U150 ( .A(n8705), .B(n8858), .Z(n8713) );
  XOR U151 ( .A(n3927), .B(n4164), .Z(n3935) );
  XOR U152 ( .A(n3642), .B(n3862), .Z(n3646) );
  XOR U153 ( .A(n3011), .B(n3251), .Z(n3012) );
  XOR U154 ( .A(n9050), .B(n9197), .Z(n9054) );
  XOR U155 ( .A(n8531), .B(n8678), .Z(n8532) );
  XOR U156 ( .A(n8158), .B(n8305), .Z(n8162) );
  XOR U157 ( .A(n7337), .B(n7484), .Z(n7338) );
  XOR U158 ( .A(n6890), .B(n7039), .Z(n6894) );
  XOR U159 ( .A(n6420), .B(n6567), .Z(n6428) );
  XOR U160 ( .A(n5926), .B(n6071), .Z(n5927) );
  XOR U161 ( .A(n5404), .B(n5551), .Z(n5408) );
  XOR U162 ( .A(n4861), .B(n5008), .Z(n4869) );
  XOR U163 ( .A(n4294), .B(n4441), .Z(n4295) );
  XOR U164 ( .A(n3309), .B(n3564), .Z(n3313) );
  XOR U165 ( .A(n2643), .B(n2947), .Z(n2647) );
  XOR U166 ( .A(n3671), .B(n3855), .Z(n3675) );
  XOR U167 ( .A(n3040), .B(n3244), .Z(n3041) );
  XOR U168 ( .A(n1997), .B(n2291), .Z(n1998) );
  XOR U169 ( .A(n9518), .B(n9656), .Z(n9522) );
  XOR U170 ( .A(n7976), .B(n8107), .Z(n7971) );
  XOR U171 ( .A(n2696), .B(n2934), .Z(n2700) );
  XOR U172 ( .A(n2026), .B(n2284), .Z(n2027) );
  XOR U173 ( .A(n3700), .B(n3848), .Z(n3704) );
  XOR U174 ( .A(n3069), .B(n3237), .Z(n3070) );
  XOR U175 ( .A(n6675), .B(n6801), .Z(n6676) );
  XOR U176 ( .A(n6190), .B(n6319), .Z(n6194) );
  XOR U177 ( .A(n5681), .B(n5810), .Z(n5689) );
  XOR U178 ( .A(n5153), .B(n5279), .Z(n5154) );
  XOR U179 ( .A(n4595), .B(n4724), .Z(n4599) );
  XOR U180 ( .A(n2677), .B(n2939), .Z(n2685) );
  XOR U181 ( .A(n1640), .B(n1962), .Z(n1644) );
  XOR U182 ( .A(n9232), .B(n9352), .Z(n9233) );
  XOR U183 ( .A(n3098), .B(n3230), .Z(n3099) );
  XOR U184 ( .A(n2725), .B(n2927), .Z(n2729) );
  XOR U185 ( .A(n2055), .B(n2277), .Z(n2056) );
  XOR U186 ( .A(n2009), .B(n2288), .Z(n2013) );
  XOR U187 ( .A(n1314), .B(n1617), .Z(n1318) );
  XOR U188 ( .A(n937), .B(n1278), .Z(n941) );
  XOR U189 ( .A(n9814), .B(n9931), .Z(n9818) );
  XOR U190 ( .A(n9074), .B(n9191), .Z(n9078) );
  XOR U191 ( .A(n8375), .B(n8485), .Z(n8376) );
  XOR U192 ( .A(n7986), .B(n8103), .Z(n7990) );
  XOR U193 ( .A(n7363), .B(n7479), .Z(n7358) );
  XOR U194 ( .A(n1693), .B(n1949), .Z(n1697) );
  XOR U195 ( .A(n988), .B(n1266), .Z(n989) );
  XOR U196 ( .A(n2754), .B(n2920), .Z(n2758) );
  XOR U197 ( .A(n2084), .B(n2270), .Z(n2085) );
  XOR U198 ( .A(n10191), .B(n10298), .Z(n10195) );
  XOR U199 ( .A(n8743), .B(n8850), .Z(n8738) );
  XOR U200 ( .A(n7789), .B(n7900), .Z(n7797) );
  XOR U201 ( .A(n6449), .B(n6560), .Z(n6457) );
  XOR U202 ( .A(n5955), .B(n6064), .Z(n5956) );
  XOR U203 ( .A(n5433), .B(n5544), .Z(n5437) );
  XOR U204 ( .A(n4890), .B(n5001), .Z(n4898) );
  XOR U205 ( .A(n4323), .B(n4434), .Z(n4324) );
  XOR U206 ( .A(n3729), .B(n3840), .Z(n3733) );
  XOR U207 ( .A(n2783), .B(n2913), .Z(n2787) );
  XOR U208 ( .A(n2113), .B(n2263), .Z(n2114) );
  XOR U209 ( .A(n1722), .B(n1942), .Z(n1726) );
  XOR U210 ( .A(n1017), .B(n1259), .Z(n1018) );
  XOR U211 ( .A(n971), .B(n1270), .Z(n975) );
  XOR U212 ( .A(n10083), .B(n10182), .Z(n10091) );
  XOR U213 ( .A(n9547), .B(n9649), .Z(n9551) );
  XOR U214 ( .A(n9249), .B(n9348), .Z(n9257) );
  XOR U215 ( .A(n8387), .B(n8482), .Z(n8391) );
  XOR U216 ( .A(n7373), .B(n7475), .Z(n7377) );
  XOR U217 ( .A(n3439), .B(n3534), .Z(n3434) );
  XOR U218 ( .A(n1000), .B(n1263), .Z(n1004) );
  XOR U219 ( .A(n1751), .B(n1935), .Z(n1755) );
  XOR U220 ( .A(n1046), .B(n1252), .Z(n1047) );
  XOR U221 ( .A(n2142), .B(n2256), .Z(n2143) );
  XOR U222 ( .A(n10425), .B(n10518), .Z(n10429) );
  XOR U223 ( .A(n8008), .B(n8098), .Z(n8009) );
  XOR U224 ( .A(n6938), .B(n7029), .Z(n6933) );
  XOR U225 ( .A(n6463), .B(n6556), .Z(n6467) );
  XOR U226 ( .A(n5967), .B(n6061), .Z(n5971) );
  XOR U227 ( .A(n5452), .B(n5541), .Z(n5447) );
  XOR U228 ( .A(n4904), .B(n4997), .Z(n4908) );
  XOR U229 ( .A(n4335), .B(n4431), .Z(n4339) );
  XOR U230 ( .A(n1780), .B(n1928), .Z(n1784) );
  XOR U231 ( .A(n1075), .B(n1245), .Z(n1076) );
  XOR U232 ( .A(n1029), .B(n1256), .Z(n1033) );
  XOR U233 ( .A(n2487), .B(n2581), .Z(n2491) );
  XOR U234 ( .A(n1479), .B(n1578), .Z(n1483) );
  XOR U235 ( .A(n10717), .B(n10798), .Z(n10721) );
  XOR U236 ( .A(n10328), .B(n10410), .Z(n10323) );
  XOR U237 ( .A(n9843), .B(n9924), .Z(n9847) );
  XOR U238 ( .A(n9566), .B(n9646), .Z(n9561) );
  XOR U239 ( .A(n8935), .B(n9018), .Z(n8939) );
  XOR U240 ( .A(n8586), .B(n8666), .Z(n8581) );
  XOR U241 ( .A(n7605), .B(n7686), .Z(n7613) );
  XOR U242 ( .A(n4055), .B(n4133), .Z(n4056) );
  XOR U243 ( .A(n3449), .B(n3530), .Z(n3453) );
  XOR U244 ( .A(n2169), .B(n2250), .Z(n2173) );
  XOR U245 ( .A(n1058), .B(n1249), .Z(n1062) );
  XOR U246 ( .A(n10634), .B(n10709), .Z(n10638) );
  XOR U247 ( .A(n7176), .B(n7247), .Z(n7180) );
  XOR U248 ( .A(n5984), .B(n6057), .Z(n5985) );
  XOR U249 ( .A(n5462), .B(n5537), .Z(n5466) );
  XOR U250 ( .A(n4919), .B(n4994), .Z(n4927) );
  XOR U251 ( .A(n1464), .B(n1581), .Z(n1468) );
  XOR U252 ( .A(n3149), .B(n3218), .Z(n3153) );
  XOR U253 ( .A(n1087), .B(n1242), .Z(n1091) );
  XOR U254 ( .A(n1136), .B(n1231), .Z(n1140) );
  XOR U255 ( .A(n10886), .B(n10952), .Z(n10890) );
  XOR U256 ( .A(n10552), .B(n10612), .Z(n10553) );
  XOR U257 ( .A(n10112), .B(n10175), .Z(n10120) );
  XOR U258 ( .A(n9860), .B(n9920), .Z(n9861) );
  XOR U259 ( .A(n9278), .B(n9341), .Z(n9286) );
  XOR U260 ( .A(n8952), .B(n9014), .Z(n8953) );
  XOR U261 ( .A(n8226), .B(n8289), .Z(n8234) );
  XOR U262 ( .A(n7830), .B(n7890), .Z(n7831) );
  XOR U263 ( .A(n6958), .B(n7023), .Z(n6966) );
  XOR U264 ( .A(n4359), .B(n4425), .Z(n4363) );
  XOR U265 ( .A(n3768), .B(n3831), .Z(n3772) );
  XOR U266 ( .A(n2184), .B(n2247), .Z(n2188) );
  XOR U267 ( .A(n1509), .B(n1572), .Z(n1513) );
  XOR U268 ( .A(n10819), .B(n10872), .Z(n10827) );
  XOR U269 ( .A(n7407), .B(n7467), .Z(n7411) );
  XOR U270 ( .A(n6733), .B(n6787), .Z(n6734) );
  XOR U271 ( .A(n6248), .B(n6305), .Z(n6252) );
  XOR U272 ( .A(n5213), .B(n5264), .Z(n5217) );
  XOR U273 ( .A(n3474), .B(n3525), .Z(n3478) );
  XOR U274 ( .A(n1171), .B(n1224), .Z(n1175) );
  XOR U275 ( .A(n11149), .B(n11204), .Z(n11153) );
  XOR U276 ( .A(n11038), .B(n11083), .Z(n11042) );
  XOR U277 ( .A(n10746), .B(n10791), .Z(n10750) );
  XOR U278 ( .A(n10357), .B(n10403), .Z(n10352) );
  XOR U279 ( .A(n10126), .B(n10171), .Z(n10130) );
  XOR U280 ( .A(n9595), .B(n9639), .Z(n9590) );
  XOR U281 ( .A(n9292), .B(n9337), .Z(n9296) );
  XOR U282 ( .A(n8615), .B(n8659), .Z(n8610) );
  XOR U283 ( .A(n8240), .B(n8285), .Z(n8244) );
  XOR U284 ( .A(n6010), .B(n6052), .Z(n6005) );
  XOR U285 ( .A(n4943), .B(n4988), .Z(n4947) );
  XOR U286 ( .A(n4374), .B(n4422), .Z(n4378) );
  XOR U287 ( .A(n3169), .B(n3214), .Z(n3173) );
  XOR U288 ( .A(n2527), .B(n2573), .Z(n2531) );
  XOR U289 ( .A(n10983), .B(n11018), .Z(n10978) );
  XOR U290 ( .A(n6507), .B(n6546), .Z(n6515) );
  XOR U291 ( .A(n7856), .B(n7885), .Z(n7851) );
  XOR U292 ( .A(n5758), .B(n5791), .Z(n5762) );
  XOR U293 ( .A(n4092), .B(n4125), .Z(n4096) );
  XOR U294 ( .A(n2209), .B(n2242), .Z(n2213) );
  XNOR U295 ( .A(n11266), .B(n11224), .Z(n11226) );
  XOR U296 ( .A(n11164), .B(n11198), .Z(n11172) );
  XOR U297 ( .A(n10915), .B(n10945), .Z(n10919) );
  XOR U298 ( .A(n10581), .B(n10605), .Z(n10582) );
  XOR U299 ( .A(n10367), .B(n10399), .Z(n10371) );
  XOR U300 ( .A(n9889), .B(n9913), .Z(n9890) );
  XOR U301 ( .A(n9605), .B(n9635), .Z(n9609) );
  XOR U302 ( .A(n8981), .B(n9007), .Z(n8982) );
  XOR U303 ( .A(n8625), .B(n8655), .Z(n8629) );
  XOR U304 ( .A(n7648), .B(n7675), .Z(n7652) );
  XOR U305 ( .A(n6272), .B(n6299), .Z(n6276) );
  XOR U306 ( .A(n5233), .B(n5260), .Z(n5237) );
  XOR U307 ( .A(n4678), .B(n4705), .Z(n4682) );
  XOR U308 ( .A(n3494), .B(n3521), .Z(n3498) );
  XOR U309 ( .A(n2867), .B(n2894), .Z(n2871) );
  XOR U310 ( .A(n1879), .B(n1906), .Z(n1883) );
  XOR U311 ( .A(n1191), .B(n1220), .Z(n1195) );
  XOR U312 ( .A(n11298), .B(n11318), .Z(n11302) );
  XOR U313 ( .A(n6595), .B(n6820), .Z(n6599) );
  XOR U314 ( .A(n7503), .B(n7710), .Z(n7507) );
  XOR U315 ( .A(n7070), .B(n7273), .Z(n7074) );
  XOR U316 ( .A(n6614), .B(n6817), .Z(n6609) );
  XOR U317 ( .A(n6127), .B(n6334), .Z(n6131) );
  XOR U318 ( .A(n5339), .B(n5567), .Z(n5340) );
  XOR U319 ( .A(n5589), .B(n5833), .Z(n5593) );
  XOR U320 ( .A(n5368), .B(n5560), .Z(n5369) );
  XOR U321 ( .A(n5618), .B(n5826), .Z(n5622) );
  XOR U322 ( .A(n7928), .B(n8117), .Z(n7932) );
  XOR U323 ( .A(n7518), .B(n7707), .Z(n7526) );
  XOR U324 ( .A(n7087), .B(n7269), .Z(n7088) );
  XOR U325 ( .A(n6624), .B(n6813), .Z(n6628) );
  XOR U326 ( .A(n5894), .B(n6080), .Z(n5889) );
  XOR U327 ( .A(n4501), .B(n4747), .Z(n4502) );
  XOR U328 ( .A(n4769), .B(n5031), .Z(n4773) );
  XOR U329 ( .A(n4530), .B(n4740), .Z(n4531) );
  XOR U330 ( .A(n5380), .B(n5557), .Z(n5384) );
  XOR U331 ( .A(n4798), .B(n5024), .Z(n4802) );
  XOR U332 ( .A(n8509), .B(n8683), .Z(n8513) );
  XOR U333 ( .A(n8139), .B(n8310), .Z(n8147) );
  XOR U334 ( .A(n7743), .B(n7911), .Z(n7744) );
  XOR U335 ( .A(n7315), .B(n7489), .Z(n7319) );
  XOR U336 ( .A(n6871), .B(n7044), .Z(n6879) );
  XOR U337 ( .A(n6403), .B(n6571), .Z(n6404) );
  XOR U338 ( .A(n5904), .B(n6076), .Z(n5908) );
  XOR U339 ( .A(n3606), .B(n3871), .Z(n3607) );
  XOR U340 ( .A(n3893), .B(n4172), .Z(n3897) );
  XOR U341 ( .A(n5121), .B(n5288), .Z(n5116) );
  XOR U342 ( .A(n4243), .B(n4453), .Z(n4247) );
  XOR U343 ( .A(n3635), .B(n3864), .Z(n3636) );
  XOR U344 ( .A(n4267), .B(n4447), .Z(n4271) );
  XOR U345 ( .A(n3922), .B(n4165), .Z(n3926) );
  XOR U346 ( .A(n9205), .B(n9358), .Z(n9209) );
  XOR U347 ( .A(n8877), .B(n9032), .Z(n8881) );
  XOR U348 ( .A(n8528), .B(n8680), .Z(n8523) );
  XOR U349 ( .A(n8153), .B(n8306), .Z(n8157) );
  XOR U350 ( .A(n7755), .B(n7908), .Z(n7759) );
  XOR U351 ( .A(n7334), .B(n7486), .Z(n7329) );
  XOR U352 ( .A(n6885), .B(n7040), .Z(n6889) );
  XOR U353 ( .A(n6415), .B(n6568), .Z(n6419) );
  XOR U354 ( .A(n5923), .B(n6073), .Z(n5918) );
  XOR U355 ( .A(n5399), .B(n5552), .Z(n5403) );
  XOR U356 ( .A(n4856), .B(n5009), .Z(n4860) );
  XOR U357 ( .A(n3664), .B(n3857), .Z(n3665) );
  XOR U358 ( .A(n2660), .B(n2943), .Z(n2661) );
  XOR U359 ( .A(n2965), .B(n3262), .Z(n2969) );
  XOR U360 ( .A(n3956), .B(n4157), .Z(n3964) );
  XOR U361 ( .A(n3333), .B(n3558), .Z(n3337) );
  XOR U362 ( .A(n2689), .B(n2936), .Z(n2690) );
  XOR U363 ( .A(n3693), .B(n3850), .Z(n3694) );
  XOR U364 ( .A(n4296), .B(n4440), .Z(n4300) );
  XOR U365 ( .A(n3314), .B(n3563), .Z(n3322) );
  XOR U366 ( .A(n1630), .B(n1964), .Z(n1634) );
  XOR U367 ( .A(n9663), .B(n9798), .Z(n9667) );
  XOR U368 ( .A(n9374), .B(n9505), .Z(n9378) );
  XOR U369 ( .A(n8719), .B(n8854), .Z(n8723) );
  XOR U370 ( .A(n8358), .B(n8489), .Z(n8362) );
  XOR U371 ( .A(n7772), .B(n7904), .Z(n7773) );
  XOR U372 ( .A(n7344), .B(n7482), .Z(n7348) );
  XOR U373 ( .A(n6900), .B(n7037), .Z(n6908) );
  XOR U374 ( .A(n6432), .B(n6564), .Z(n6433) );
  XOR U375 ( .A(n5933), .B(n6069), .Z(n5937) );
  XOR U376 ( .A(n5414), .B(n5549), .Z(n5422) );
  XOR U377 ( .A(n4873), .B(n5005), .Z(n4874) );
  XOR U378 ( .A(n3985), .B(n4150), .Z(n3993) );
  XOR U379 ( .A(n3362), .B(n3551), .Z(n3366) );
  XOR U380 ( .A(n2718), .B(n2929), .Z(n2719) );
  XOR U381 ( .A(n2672), .B(n2940), .Z(n2676) );
  XOR U382 ( .A(n1999), .B(n2290), .Z(n2003) );
  XOR U383 ( .A(n1980), .B(n2295), .Z(n1984) );
  XOR U384 ( .A(n3028), .B(n3247), .Z(n3036) );
  XOR U385 ( .A(n2366), .B(n2611), .Z(n2370) );
  XOR U386 ( .A(n1686), .B(n1951), .Z(n1687) );
  XOR U387 ( .A(n4014), .B(n4143), .Z(n4022) );
  XOR U388 ( .A(n3391), .B(n3544), .Z(n3395) );
  XOR U389 ( .A(n2747), .B(n2922), .Z(n2748) );
  XOR U390 ( .A(n4600), .B(n4723), .Z(n4604) );
  XOR U391 ( .A(n959), .B(n1273), .Z(n960) );
  XOR U392 ( .A(n9944), .B(n10061), .Z(n9948) );
  XOR U393 ( .A(n9678), .B(n9795), .Z(n9686) );
  XOR U394 ( .A(n9234), .B(n9351), .Z(n9238) );
  XOR U395 ( .A(n8906), .B(n9025), .Z(n8910) );
  XOR U396 ( .A(n8557), .B(n8673), .Z(n8552) );
  XOR U397 ( .A(n8182), .B(n8299), .Z(n8186) );
  XOR U398 ( .A(n7784), .B(n7901), .Z(n7788) );
  XOR U399 ( .A(n7145), .B(n7255), .Z(n7146) );
  XOR U400 ( .A(n6682), .B(n6799), .Z(n6686) );
  XOR U401 ( .A(n6200), .B(n6317), .Z(n6208) );
  XOR U402 ( .A(n5693), .B(n5807), .Z(n5694) );
  XOR U403 ( .A(n5160), .B(n5277), .Z(n5164) );
  XOR U404 ( .A(n2776), .B(n2915), .Z(n2777) );
  XOR U405 ( .A(n3057), .B(n3240), .Z(n3065) );
  XOR U406 ( .A(n2395), .B(n2604), .Z(n2399) );
  XOR U407 ( .A(n1715), .B(n1944), .Z(n1716) );
  XOR U408 ( .A(n2014), .B(n2287), .Z(n2022) );
  XOR U409 ( .A(n1319), .B(n1616), .Z(n1323) );
  XOR U410 ( .A(n942), .B(n1277), .Z(n946) );
  XOR U411 ( .A(n9540), .B(n9651), .Z(n9541) );
  XOR U412 ( .A(n4028), .B(n4139), .Z(n4032) );
  XOR U413 ( .A(n2043), .B(n2280), .Z(n2051) );
  XOR U414 ( .A(n1348), .B(n1609), .Z(n1352) );
  XOR U415 ( .A(n631), .B(n913), .Z(n632) );
  XOR U416 ( .A(n3086), .B(n3233), .Z(n3094) );
  XOR U417 ( .A(n2424), .B(n2597), .Z(n2428) );
  XOR U418 ( .A(n1744), .B(n1937), .Z(n1745) );
  XOR U419 ( .A(n10304), .B(n10414), .Z(n10308) );
  XOR U420 ( .A(n4899), .B(n5000), .Z(n4894) );
  XOR U421 ( .A(n3734), .B(n3839), .Z(n3738) );
  XOR U422 ( .A(n10201), .B(n10296), .Z(n10205) );
  XOR U423 ( .A(n9963), .B(n10058), .Z(n9958) );
  XOR U424 ( .A(n9403), .B(n9498), .Z(n9407) );
  XOR U425 ( .A(n9093), .B(n9188), .Z(n9088) );
  XOR U426 ( .A(n8567), .B(n8669), .Z(n8571) );
  XOR U427 ( .A(n8197), .B(n8296), .Z(n8205) );
  XOR U428 ( .A(n7590), .B(n7689), .Z(n7594) );
  XOR U429 ( .A(n7157), .B(n7252), .Z(n7161) );
  XOR U430 ( .A(n6701), .B(n6796), .Z(n6696) );
  XOR U431 ( .A(n6214), .B(n6313), .Z(n6218) );
  XOR U432 ( .A(n5705), .B(n5804), .Z(n5709) );
  XOR U433 ( .A(n2807), .B(n2906), .Z(n2811) );
  XOR U434 ( .A(n3115), .B(n3226), .Z(n3123) );
  XOR U435 ( .A(n2453), .B(n2590), .Z(n2457) );
  XOR U436 ( .A(n1773), .B(n1930), .Z(n1774) );
  XOR U437 ( .A(n2072), .B(n2273), .Z(n2080) );
  XOR U438 ( .A(n1377), .B(n1602), .Z(n1381) );
  XOR U439 ( .A(n660), .B(n906), .Z(n661) );
  XOR U440 ( .A(n976), .B(n1269), .Z(n984) );
  XOR U441 ( .A(n9833), .B(n9926), .Z(n9837) );
  XOR U442 ( .A(n8925), .B(n9020), .Z(n8929) );
  XOR U443 ( .A(n4624), .B(n4717), .Z(n4628) );
  XOR U444 ( .A(n1005), .B(n1262), .Z(n1013) );
  XOR U445 ( .A(n2101), .B(n2266), .Z(n2109) );
  XOR U446 ( .A(n1406), .B(n1595), .Z(n1410) );
  XOR U447 ( .A(n689), .B(n899), .Z(n690) );
  XOR U448 ( .A(n1802), .B(n1923), .Z(n1803) );
  XOR U449 ( .A(n10530), .B(n10617), .Z(n10534) );
  XOR U450 ( .A(n5455), .B(n5539), .Z(n5456) );
  XOR U451 ( .A(n4340), .B(n4430), .Z(n4348) );
  XOR U452 ( .A(n10435), .B(n10516), .Z(n10443) );
  XOR U453 ( .A(n10218), .B(n10292), .Z(n10219) );
  XOR U454 ( .A(n9707), .B(n9788), .Z(n9715) );
  XOR U455 ( .A(n9420), .B(n9494), .Z(n9421) );
  XOR U456 ( .A(n8763), .B(n8844), .Z(n8771) );
  XOR U457 ( .A(n8404), .B(n8478), .Z(n8405) );
  XOR U458 ( .A(n7813), .B(n7894), .Z(n7817) );
  XOR U459 ( .A(n7392), .B(n7472), .Z(n7387) );
  XOR U460 ( .A(n6711), .B(n6792), .Z(n6715) );
  XOR U461 ( .A(n6229), .B(n6310), .Z(n6237) );
  XOR U462 ( .A(n3753), .B(n3834), .Z(n3757) );
  XOR U463 ( .A(n3139), .B(n3220), .Z(n3143) );
  XOR U464 ( .A(n2497), .B(n2579), .Z(n2501) );
  XOR U465 ( .A(n2130), .B(n2259), .Z(n2138) );
  XOR U466 ( .A(n1435), .B(n1588), .Z(n1439) );
  XOR U467 ( .A(n718), .B(n892), .Z(n719) );
  XOR U468 ( .A(n1034), .B(n1255), .Z(n1042) );
  XOR U469 ( .A(n2154), .B(n2253), .Z(n2158) );
  XOR U470 ( .A(n1834), .B(n1915), .Z(n1838) );
  XOR U471 ( .A(n1126), .B(n1233), .Z(n1130) );
  XOR U472 ( .A(n10102), .B(n10177), .Z(n10106) );
  XOR U473 ( .A(n9268), .B(n9343), .Z(n9272) );
  XOR U474 ( .A(n8216), .B(n8291), .Z(n8220) );
  XOR U475 ( .A(n5194), .B(n5269), .Z(n5198) );
  XOR U476 ( .A(n1063), .B(n1248), .Z(n1071) );
  XOR U477 ( .A(n747), .B(n885), .Z(n748) );
  XOR U478 ( .A(n10881), .B(n10953), .Z(n10885) );
  XOR U479 ( .A(n10727), .B(n10796), .Z(n10731) );
  XOR U480 ( .A(n4928), .B(n4993), .Z(n4923) );
  XOR U481 ( .A(n1111), .B(n1236), .Z(n1115) );
  XOR U482 ( .A(n1156), .B(n1227), .Z(n1160) );
  XOR U483 ( .A(n10648), .B(n10707), .Z(n10643) );
  XOR U484 ( .A(n10449), .B(n10512), .Z(n10453) );
  XOR U485 ( .A(n9992), .B(n10051), .Z(n9987) );
  XOR U486 ( .A(n9721), .B(n9784), .Z(n9725) );
  XOR U487 ( .A(n9122), .B(n9181), .Z(n9117) );
  XOR U488 ( .A(n8777), .B(n8840), .Z(n8781) );
  XOR U489 ( .A(n8034), .B(n8093), .Z(n8029) );
  XOR U490 ( .A(n7619), .B(n7682), .Z(n7623) );
  XOR U491 ( .A(n6490), .B(n6550), .Z(n6491) );
  XOR U492 ( .A(n4648), .B(n4711), .Z(n4652) );
  XOR U493 ( .A(n4067), .B(n4130), .Z(n4071) );
  XOR U494 ( .A(n3464), .B(n3527), .Z(n3468) );
  XOR U495 ( .A(n2512), .B(n2576), .Z(n2516) );
  XOR U496 ( .A(n1092), .B(n1241), .Z(n1100) );
  XOR U497 ( .A(n1849), .B(n1912), .Z(n1853) );
  XOR U498 ( .A(n1141), .B(n1230), .Z(n1145) );
  XOR U499 ( .A(n10343), .B(n10405), .Z(n10347) );
  XOR U500 ( .A(n9581), .B(n9641), .Z(n9585) );
  XOR U501 ( .A(n8601), .B(n8661), .Z(n8605) );
  XOR U502 ( .A(n5996), .B(n6054), .Z(n6000) );
  XOR U503 ( .A(n10896), .B(n10950), .Z(n10904) );
  XOR U504 ( .A(n7412), .B(n7466), .Z(n7420) );
  XOR U505 ( .A(n5748), .B(n5795), .Z(n5743) );
  XOR U506 ( .A(n1519), .B(n1570), .Z(n1523) );
  XOR U507 ( .A(n10831), .B(n10869), .Z(n10832) );
  XOR U508 ( .A(n10658), .B(n10703), .Z(n10662) );
  XOR U509 ( .A(n10247), .B(n10285), .Z(n10248) );
  XOR U510 ( .A(n10002), .B(n10047), .Z(n10006) );
  XOR U511 ( .A(n9449), .B(n9487), .Z(n9450) );
  XOR U512 ( .A(n9132), .B(n9177), .Z(n9136) );
  XOR U513 ( .A(n8433), .B(n8471), .Z(n8434) );
  XOR U514 ( .A(n8044), .B(n8089), .Z(n8048) );
  XOR U515 ( .A(n7203), .B(n7241), .Z(n7204) );
  XOR U516 ( .A(n6740), .B(n6785), .Z(n6744) );
  XOR U517 ( .A(n5218), .B(n5263), .Z(n5222) );
  XOR U518 ( .A(n4663), .B(n4708), .Z(n4667) );
  XOR U519 ( .A(n4082), .B(n4127), .Z(n4086) );
  XOR U520 ( .A(n3479), .B(n3524), .Z(n3483) );
  XOR U521 ( .A(n2852), .B(n2897), .Z(n2856) );
  XOR U522 ( .A(n2199), .B(n2244), .Z(n2203) );
  XOR U523 ( .A(n1176), .B(n1223), .Z(n1180) );
  XNOR U524 ( .A(n11256), .B(n11214), .Z(n11216) );
  XOR U525 ( .A(n11154), .B(n11202), .Z(n11158) );
  XOR U526 ( .A(n10569), .B(n10608), .Z(n10577) );
  XOR U527 ( .A(n9877), .B(n9916), .Z(n9885) );
  XOR U528 ( .A(n8969), .B(n9010), .Z(n8977) );
  XOR U529 ( .A(n11052), .B(n11081), .Z(n11047) );
  XOR U530 ( .A(n6270), .B(n6300), .Z(n6271) );
  XOR U531 ( .A(n10988), .B(n11015), .Z(n10992) );
  XOR U532 ( .A(n10843), .B(n10866), .Z(n10847) );
  XOR U533 ( .A(n10478), .B(n10505), .Z(n10482) );
  XOR U534 ( .A(n10259), .B(n10282), .Z(n10263) );
  XOR U535 ( .A(n9750), .B(n9777), .Z(n9754) );
  XOR U536 ( .A(n9461), .B(n9484), .Z(n9465) );
  XOR U537 ( .A(n8806), .B(n8833), .Z(n8810) );
  XOR U538 ( .A(n8445), .B(n8468), .Z(n8449) );
  XOR U539 ( .A(n7859), .B(n7883), .Z(n7860) );
  XOR U540 ( .A(n7431), .B(n7461), .Z(n7435) );
  XOR U541 ( .A(n6759), .B(n6782), .Z(n6754) );
  XOR U542 ( .A(n6020), .B(n6048), .Z(n6024) );
  XOR U543 ( .A(n4958), .B(n4985), .Z(n4962) );
  XOR U544 ( .A(n4389), .B(n4419), .Z(n4393) );
  XOR U545 ( .A(n3184), .B(n3211), .Z(n3188) );
  XOR U546 ( .A(n2542), .B(n2570), .Z(n2546) );
  XOR U547 ( .A(n1539), .B(n1566), .Z(n1543) );
  XOR U548 ( .A(n839), .B(n866), .Z(n843) );
  XOR U549 ( .A(n11325), .B(n11345), .Z(n11329) );
  XOR U550 ( .A(n11265), .B(n11285), .Z(n11269) );
  XNOR U551 ( .A(n11271), .B(n11229), .Z(n11231) );
  XOR U552 ( .A(n10770), .B(n10787), .Z(n10765) );
  XOR U553 ( .A(n10150), .B(n10167), .Z(n10145) );
  XOR U554 ( .A(n9316), .B(n9333), .Z(n9311) );
  XOR U555 ( .A(n8264), .B(n8281), .Z(n8259) );
  XOR U556 ( .A(n7220), .B(n7237), .Z(n7228) );
  XOR U557 ( .A(n5768), .B(n5789), .Z(n5772) );
  XOR U558 ( .A(n4102), .B(n4123), .Z(n4106) );
  XOR U559 ( .A(n2219), .B(n2240), .Z(n2223) );
  XOR U560 ( .A(n6827), .B(n7054), .Z(n6831) );
  XOR U561 ( .A(n6357), .B(n6582), .Z(n6361) );
  XOR U562 ( .A(n5841), .B(n6092), .Z(n5845) );
  XOR U563 ( .A(n7286), .B(n7496), .Z(n7290) );
  XOR U564 ( .A(n6842), .B(n7051), .Z(n6850) );
  XOR U565 ( .A(n6374), .B(n6578), .Z(n6375) );
  XOR U566 ( .A(n5608), .B(n5828), .Z(n5612) );
  XOR U567 ( .A(n5856), .B(n6089), .Z(n5864) );
  XOR U568 ( .A(n5317), .B(n5572), .Z(n5321) );
  XOR U569 ( .A(n4759), .B(n5033), .Z(n4763) );
  XOR U570 ( .A(n8124), .B(n8313), .Z(n8128) );
  XOR U571 ( .A(n7726), .B(n7915), .Z(n7730) );
  XOR U572 ( .A(n7305), .B(n7493), .Z(n7300) );
  XOR U573 ( .A(n6856), .B(n7047), .Z(n6860) );
  XOR U574 ( .A(n6386), .B(n6575), .Z(n6390) );
  XOR U575 ( .A(n5623), .B(n5825), .Z(n5631) );
  XOR U576 ( .A(n5073), .B(n5298), .Z(n5077) );
  XOR U577 ( .A(n5336), .B(n5569), .Z(n5331) );
  XOR U578 ( .A(n4503), .B(n4746), .Z(n4507) );
  XOR U579 ( .A(n4774), .B(n5030), .Z(n4782) );
  XOR U580 ( .A(n4185), .B(n4467), .Z(n4189) );
  XOR U581 ( .A(n5102), .B(n5291), .Z(n5106) );
  XOR U582 ( .A(n3579), .B(n3877), .Z(n3583) );
  XOR U583 ( .A(n4532), .B(n4739), .Z(n4536) );
  XOR U584 ( .A(n8690), .B(n8861), .Z(n8694) );
  XOR U585 ( .A(n8329), .B(n8496), .Z(n8333) );
  XOR U586 ( .A(n7947), .B(n8114), .Z(n7942) );
  XOR U587 ( .A(n7532), .B(n7703), .Z(n7536) );
  XOR U588 ( .A(n7099), .B(n7266), .Z(n7103) );
  XOR U589 ( .A(n6643), .B(n6810), .Z(n6638) );
  XOR U590 ( .A(n6156), .B(n6327), .Z(n6160) );
  XOR U591 ( .A(n5647), .B(n5818), .Z(n5651) );
  XOR U592 ( .A(n4559), .B(n4733), .Z(n4560) );
  XOR U593 ( .A(n5092), .B(n5295), .Z(n5087) );
  XOR U594 ( .A(n4518), .B(n4743), .Z(n4526) );
  XOR U595 ( .A(n3917), .B(n4166), .Z(n3921) );
  XOR U596 ( .A(n4204), .B(n4464), .Z(n4199) );
  XOR U597 ( .A(n4832), .B(n5016), .Z(n4840) );
  XOR U598 ( .A(n3594), .B(n3874), .Z(n3602) );
  XOR U599 ( .A(n2960), .B(n3263), .Z(n2964) );
  XOR U600 ( .A(n4248), .B(n4452), .Z(n4252) );
  XOR U601 ( .A(n9045), .B(n9198), .Z(n9049) );
  XOR U602 ( .A(n8346), .B(n8492), .Z(n8347) );
  XOR U603 ( .A(n7957), .B(n8110), .Z(n7961) );
  XOR U604 ( .A(n7547), .B(n7700), .Z(n7555) );
  XOR U605 ( .A(n7116), .B(n7262), .Z(n7117) );
  XOR U606 ( .A(n6653), .B(n6806), .Z(n6657) );
  XOR U607 ( .A(n6171), .B(n6324), .Z(n6179) );
  XOR U608 ( .A(n5664), .B(n5814), .Z(n5665) );
  XOR U609 ( .A(n5131), .B(n5284), .Z(n5135) );
  XOR U610 ( .A(n4272), .B(n4446), .Z(n4276) );
  XOR U611 ( .A(n2303), .B(n2627), .Z(n2307) );
  XOR U612 ( .A(n3328), .B(n3559), .Z(n3332) );
  XOR U613 ( .A(n9364), .B(n9507), .Z(n9368) );
  XOR U614 ( .A(n8882), .B(n9031), .Z(n8890) );
  XOR U615 ( .A(n4576), .B(n4729), .Z(n4584) );
  XOR U616 ( .A(n3936), .B(n4163), .Z(n3931) );
  XOR U617 ( .A(n2662), .B(n2942), .Z(n2666) );
  XOR U618 ( .A(n3357), .B(n3552), .Z(n3361) );
  XOR U619 ( .A(n2994), .B(n3255), .Z(n2998) );
  XOR U620 ( .A(n2979), .B(n3260), .Z(n2974) );
  XOR U621 ( .A(n3965), .B(n4156), .Z(n3960) );
  XOR U622 ( .A(n8538), .B(n8676), .Z(n8542) );
  XOR U623 ( .A(n8168), .B(n8303), .Z(n8176) );
  XOR U624 ( .A(n7561), .B(n7696), .Z(n7565) );
  XOR U625 ( .A(n7128), .B(n7259), .Z(n7132) );
  XOR U626 ( .A(n6672), .B(n6803), .Z(n6667) );
  XOR U627 ( .A(n6185), .B(n6320), .Z(n6189) );
  XOR U628 ( .A(n5676), .B(n5811), .Z(n5680) );
  XOR U629 ( .A(n5150), .B(n5281), .Z(n5145) );
  XOR U630 ( .A(n4590), .B(n4725), .Z(n4594) );
  XOR U631 ( .A(n2318), .B(n2624), .Z(n2326) );
  XOR U632 ( .A(n1635), .B(n1963), .Z(n1639) );
  XOR U633 ( .A(n3343), .B(n3556), .Z(n3351) );
  XOR U634 ( .A(n4009), .B(n4144), .Z(n4013) );
  XOR U635 ( .A(n3386), .B(n3545), .Z(n3390) );
  XOR U636 ( .A(n9668), .B(n9797), .Z(n9672) );
  XOR U637 ( .A(n9379), .B(n9504), .Z(n9387) );
  XOR U638 ( .A(n9067), .B(n9193), .Z(n9068) );
  XOR U639 ( .A(n7979), .B(n8105), .Z(n7980) );
  XOR U640 ( .A(n3994), .B(n4149), .Z(n3989) );
  XOR U641 ( .A(n2004), .B(n2289), .Z(n2008) );
  XOR U642 ( .A(n3372), .B(n3549), .Z(n3380) );
  XOR U643 ( .A(n2686), .B(n2938), .Z(n2681) );
  XOR U644 ( .A(n2371), .B(n2610), .Z(n2375) );
  XOR U645 ( .A(n1688), .B(n1950), .Z(n1692) );
  XOR U646 ( .A(n10068), .B(n10185), .Z(n10072) );
  XOR U647 ( .A(n8734), .B(n8851), .Z(n8742) );
  XOR U648 ( .A(n7576), .B(n7693), .Z(n7584) );
  XOR U649 ( .A(n6914), .B(n7033), .Z(n6918) );
  XOR U650 ( .A(n6444), .B(n6561), .Z(n6448) );
  XOR U651 ( .A(n5952), .B(n6066), .Z(n5947) );
  XOR U652 ( .A(n5428), .B(n5545), .Z(n5432) );
  XOR U653 ( .A(n4885), .B(n5002), .Z(n4889) );
  XOR U654 ( .A(n4320), .B(n4436), .Z(n4315) );
  XOR U655 ( .A(n3724), .B(n3841), .Z(n3728) );
  XOR U656 ( .A(n602), .B(n920), .Z(n603) );
  XOR U657 ( .A(n1654), .B(n1960), .Z(n1649) );
  XOR U658 ( .A(n2715), .B(n2931), .Z(n2710) );
  XOR U659 ( .A(n3401), .B(n3542), .Z(n3409) );
  XOR U660 ( .A(n9949), .B(n10060), .Z(n9953) );
  XOR U661 ( .A(n9687), .B(n9794), .Z(n9682) );
  XOR U662 ( .A(n9393), .B(n9500), .Z(n9397) );
  XOR U663 ( .A(n9079), .B(n9190), .Z(n9083) );
  XOR U664 ( .A(n8560), .B(n8671), .Z(n8561) );
  XOR U665 ( .A(n8187), .B(n8298), .Z(n8191) );
  XOR U666 ( .A(n7366), .B(n7477), .Z(n7367) );
  XOR U667 ( .A(n3425), .B(n3536), .Z(n3429) );
  XOR U668 ( .A(n2400), .B(n2603), .Z(n2404) );
  XOR U669 ( .A(n1717), .B(n1943), .Z(n1721) );
  XOR U670 ( .A(n1674), .B(n1954), .Z(n1682) );
  XOR U671 ( .A(n966), .B(n1271), .Z(n970) );
  XOR U672 ( .A(n947), .B(n1276), .Z(n955) );
  XOR U673 ( .A(n2744), .B(n2924), .Z(n2739) );
  XOR U674 ( .A(n1703), .B(n1947), .Z(n1711) );
  XOR U675 ( .A(n995), .B(n1264), .Z(n999) );
  XOR U676 ( .A(n2429), .B(n2596), .Z(n2433) );
  XOR U677 ( .A(n1746), .B(n1936), .Z(n1750) );
  XOR U678 ( .A(n10309), .B(n10413), .Z(n10313) );
  XOR U679 ( .A(n8005), .B(n8100), .Z(n8000) );
  XOR U680 ( .A(n6929), .B(n7030), .Z(n6937) );
  XOR U681 ( .A(n6461), .B(n6557), .Z(n6462) );
  XOR U682 ( .A(n5962), .B(n6062), .Z(n5966) );
  XOR U683 ( .A(n5443), .B(n5542), .Z(n5451) );
  XOR U684 ( .A(n4902), .B(n4998), .Z(n4903) );
  XOR U685 ( .A(n4330), .B(n4432), .Z(n4334) );
  XOR U686 ( .A(n2773), .B(n2917), .Z(n2768) );
  XOR U687 ( .A(n10206), .B(n10295), .Z(n10214) );
  XOR U688 ( .A(n9966), .B(n10056), .Z(n9967) );
  XOR U689 ( .A(n9697), .B(n9790), .Z(n9701) );
  XOR U690 ( .A(n9408), .B(n9497), .Z(n9416) );
  XOR U691 ( .A(n9096), .B(n9186), .Z(n9097) );
  XOR U692 ( .A(n8753), .B(n8846), .Z(n8757) );
  XOR U693 ( .A(n8392), .B(n8481), .Z(n8400) );
  XOR U694 ( .A(n7803), .B(n7896), .Z(n7807) );
  XOR U695 ( .A(n7378), .B(n7474), .Z(n7382) );
  XOR U696 ( .A(n3748), .B(n3837), .Z(n3743) );
  XOR U697 ( .A(n3129), .B(n3222), .Z(n3133) );
  XOR U698 ( .A(n2458), .B(n2589), .Z(n2462) );
  XOR U699 ( .A(n1775), .B(n1929), .Z(n1779) );
  XOR U700 ( .A(n1732), .B(n1940), .Z(n1740) );
  XOR U701 ( .A(n1024), .B(n1257), .Z(n1028) );
  XOR U702 ( .A(n985), .B(n1268), .Z(n980) );
  XOR U703 ( .A(n2802), .B(n2910), .Z(n2797) );
  XOR U704 ( .A(n1014), .B(n1261), .Z(n1009) );
  XOR U705 ( .A(n1761), .B(n1933), .Z(n1769) );
  XOR U706 ( .A(n1053), .B(n1250), .Z(n1057) );
  XOR U707 ( .A(n2149), .B(n2254), .Z(n2153) );
  XOR U708 ( .A(n10535), .B(n10616), .Z(n10539) );
  XOR U709 ( .A(n7174), .B(n7248), .Z(n7175) );
  XOR U710 ( .A(n6473), .B(n6554), .Z(n6477) );
  XOR U711 ( .A(n5981), .B(n6059), .Z(n5976) );
  XOR U712 ( .A(n5457), .B(n5538), .Z(n5461) );
  XOR U713 ( .A(n4914), .B(n4995), .Z(n4918) );
  XOR U714 ( .A(n1459), .B(n1582), .Z(n1463) );
  XOR U715 ( .A(n10804), .B(n10875), .Z(n10808) );
  XOR U716 ( .A(n10444), .B(n10515), .Z(n10439) );
  XOR U717 ( .A(n10220), .B(n10291), .Z(n10224) );
  XOR U718 ( .A(n9978), .B(n10053), .Z(n9982) );
  XOR U719 ( .A(n9716), .B(n9787), .Z(n9711) );
  XOR U720 ( .A(n9422), .B(n9493), .Z(n9426) );
  XOR U721 ( .A(n9108), .B(n9183), .Z(n9112) );
  XOR U722 ( .A(n8772), .B(n8843), .Z(n8767) );
  XOR U723 ( .A(n8406), .B(n8477), .Z(n8410) );
  XOR U724 ( .A(n8020), .B(n8095), .Z(n8024) );
  XOR U725 ( .A(n7614), .B(n7685), .Z(n7609) );
  XOR U726 ( .A(n6948), .B(n7025), .Z(n6952) );
  XOR U727 ( .A(n4643), .B(n4714), .Z(n4638) );
  XOR U728 ( .A(n4057), .B(n4132), .Z(n4061) );
  XOR U729 ( .A(n3454), .B(n3529), .Z(n3458) );
  XOR U730 ( .A(n2827), .B(n2902), .Z(n2831) );
  XOR U731 ( .A(n2174), .B(n2249), .Z(n2178) );
  XOR U732 ( .A(n1790), .B(n1926), .Z(n1798) );
  XOR U733 ( .A(n1082), .B(n1243), .Z(n1086) );
  XOR U734 ( .A(n1043), .B(n1254), .Z(n1038) );
  XOR U735 ( .A(n769), .B(n880), .Z(n773) );
  XOR U736 ( .A(n1072), .B(n1247), .Z(n1067) );
  XOR U737 ( .A(n1819), .B(n1919), .Z(n1823) );
  XOR U738 ( .A(n10732), .B(n10795), .Z(n10740) );
  XOR U739 ( .A(n6730), .B(n6789), .Z(n6725) );
  XOR U740 ( .A(n6243), .B(n6306), .Z(n6247) );
  XOR U741 ( .A(n5734), .B(n5797), .Z(n5738) );
  XOR U742 ( .A(n1116), .B(n1235), .Z(n1120) );
  XOR U743 ( .A(n799), .B(n874), .Z(n803) );
  XOR U744 ( .A(n10964), .B(n11021), .Z(n10968) );
  XOR U745 ( .A(n10651), .B(n10705), .Z(n10652) );
  XOR U746 ( .A(n10454), .B(n10511), .Z(n10458) );
  XOR U747 ( .A(n10235), .B(n10288), .Z(n10243) );
  XOR U748 ( .A(n9995), .B(n10049), .Z(n9996) );
  XOR U749 ( .A(n9726), .B(n9783), .Z(n9730) );
  XOR U750 ( .A(n9437), .B(n9490), .Z(n9445) );
  XOR U751 ( .A(n9125), .B(n9179), .Z(n9126) );
  XOR U752 ( .A(n8782), .B(n8839), .Z(n8786) );
  XOR U753 ( .A(n8421), .B(n8474), .Z(n8429) );
  XOR U754 ( .A(n8037), .B(n8091), .Z(n8038) );
  XOR U755 ( .A(n7624), .B(n7681), .Z(n7628) );
  XOR U756 ( .A(n7191), .B(n7244), .Z(n7199) );
  XOR U757 ( .A(n5481), .B(n5534), .Z(n5476) );
  XOR U758 ( .A(n4933), .B(n4990), .Z(n4937) );
  XOR U759 ( .A(n4364), .B(n4424), .Z(n4368) );
  XOR U760 ( .A(n3773), .B(n3830), .Z(n3777) );
  XOR U761 ( .A(n3159), .B(n3216), .Z(n3163) );
  XOR U762 ( .A(n2517), .B(n2575), .Z(n2521) );
  XOR U763 ( .A(n1854), .B(n1911), .Z(n1858) );
  XOR U764 ( .A(n1101), .B(n1240), .Z(n1096) );
  XOR U765 ( .A(n1146), .B(n1229), .Z(n1150) );
  XOR U766 ( .A(n1166), .B(n1225), .Z(n1170) );
  XOR U767 ( .A(n10905), .B(n10949), .Z(n10900) );
  XOR U768 ( .A(n6972), .B(n7019), .Z(n6976) );
  XOR U769 ( .A(n6502), .B(n6547), .Z(n6506) );
  XOR U770 ( .A(n11211), .B(n11249), .Z(n11215) );
  XOR U771 ( .A(n11101), .B(n11141), .Z(n11105) );
  XOR U772 ( .A(n10833), .B(n10868), .Z(n10837) );
  XOR U773 ( .A(n10663), .B(n10702), .Z(n10667) );
  XOR U774 ( .A(n10473), .B(n10508), .Z(n10468) );
  XOR U775 ( .A(n10249), .B(n10284), .Z(n10253) );
  XOR U776 ( .A(n10007), .B(n10046), .Z(n10011) );
  XOR U777 ( .A(n9745), .B(n9780), .Z(n9740) );
  XOR U778 ( .A(n9451), .B(n9486), .Z(n9455) );
  XOR U779 ( .A(n9137), .B(n9176), .Z(n9141) );
  XOR U780 ( .A(n8801), .B(n8836), .Z(n8796) );
  XOR U781 ( .A(n8435), .B(n8470), .Z(n8439) );
  XOR U782 ( .A(n8049), .B(n8088), .Z(n8053) );
  XOR U783 ( .A(n7643), .B(n7678), .Z(n7638) );
  XOR U784 ( .A(n6267), .B(n6302), .Z(n6262) );
  XOR U785 ( .A(n5753), .B(n5792), .Z(n5757) );
  XOR U786 ( .A(n5223), .B(n5262), .Z(n5227) );
  XOR U787 ( .A(n4668), .B(n4707), .Z(n4672) );
  XOR U788 ( .A(n4087), .B(n4126), .Z(n4091) );
  XOR U789 ( .A(n3484), .B(n3523), .Z(n3488) );
  XOR U790 ( .A(n2857), .B(n2896), .Z(n2861) );
  XOR U791 ( .A(n2204), .B(n2243), .Z(n2208) );
  XOR U792 ( .A(n1529), .B(n1568), .Z(n1533) );
  XOR U793 ( .A(n829), .B(n868), .Z(n833) );
  XOR U794 ( .A(n11055), .B(n11079), .Z(n11056) );
  XOR U795 ( .A(n7215), .B(n7238), .Z(n7219) );
  XNOR U796 ( .A(n11352), .B(n11328), .Z(n11330) );
  XNOR U797 ( .A(n11331), .B(n11301), .Z(n11303) );
  XNOR U798 ( .A(n11304), .B(n11268), .Z(n11270) );
  XOR U799 ( .A(n11226), .B(n11246), .Z(n11230) );
  XOR U800 ( .A(n10993), .B(n11014), .Z(n10997) );
  XOR U801 ( .A(n10848), .B(n10865), .Z(n10856) );
  XOR U802 ( .A(n10680), .B(n10698), .Z(n10681) );
  XOR U803 ( .A(n10483), .B(n10504), .Z(n10487) );
  XOR U804 ( .A(n10264), .B(n10281), .Z(n10272) );
  XOR U805 ( .A(n10024), .B(n10042), .Z(n10025) );
  XOR U806 ( .A(n9755), .B(n9776), .Z(n9759) );
  XOR U807 ( .A(n9466), .B(n9483), .Z(n9474) );
  XOR U808 ( .A(n9154), .B(n9172), .Z(n9155) );
  XOR U809 ( .A(n8811), .B(n8832), .Z(n8815) );
  XOR U810 ( .A(n8450), .B(n8467), .Z(n8458) );
  XOR U811 ( .A(n8066), .B(n8084), .Z(n8067) );
  XOR U812 ( .A(n7653), .B(n7674), .Z(n7657) );
  XOR U813 ( .A(n6996), .B(n7015), .Z(n6991) );
  XOR U814 ( .A(n6521), .B(n6542), .Z(n6525) );
  XOR U815 ( .A(n6025), .B(n6047), .Z(n6029) );
  XOR U816 ( .A(n5506), .B(n5527), .Z(n5510) );
  XOR U817 ( .A(n4963), .B(n4984), .Z(n4967) );
  XOR U818 ( .A(n4394), .B(n4418), .Z(n4398) );
  XOR U819 ( .A(n3803), .B(n3824), .Z(n3807) );
  XOR U820 ( .A(n3189), .B(n3210), .Z(n3193) );
  XOR U821 ( .A(n2547), .B(n2569), .Z(n2551) );
  XOR U822 ( .A(n1884), .B(n1905), .Z(n1888) );
  XOR U823 ( .A(n1196), .B(n1219), .Z(n1200) );
  XNOR U824 ( .A(n11235), .B(n11234), .Z(n11192) );
  XNOR U825 ( .A(n11185), .B(n11184), .Z(n11179) );
  XOR U826 ( .A(n6347), .B(n6584), .Z(n6351) );
  XOR U827 ( .A(n6832), .B(n7053), .Z(n6836) );
  XOR U828 ( .A(n6362), .B(n6581), .Z(n6370) );
  XOR U829 ( .A(n5846), .B(n6091), .Z(n5850) );
  XOR U830 ( .A(n5312), .B(n5573), .Z(n5316) );
  XOR U831 ( .A(n7716), .B(n7917), .Z(n7720) );
  XOR U832 ( .A(n7291), .B(n7495), .Z(n7295) );
  XOR U833 ( .A(n6851), .B(n7050), .Z(n6846) );
  XOR U834 ( .A(n6376), .B(n6577), .Z(n6380) );
  XOR U835 ( .A(n5613), .B(n5827), .Z(n5617) );
  XOR U836 ( .A(n5865), .B(n6088), .Z(n5860) );
  XOR U837 ( .A(n5068), .B(n5299), .Z(n5072) );
  XOR U838 ( .A(n5327), .B(n5570), .Z(n5335) );
  XOR U839 ( .A(n4764), .B(n5032), .Z(n4768) );
  XOR U840 ( .A(n4180), .B(n4468), .Z(n4184) );
  XOR U841 ( .A(n8129), .B(n8312), .Z(n8133) );
  XOR U842 ( .A(n7731), .B(n7914), .Z(n7739) );
  XOR U843 ( .A(n7308), .B(n7491), .Z(n7309) );
  XOR U844 ( .A(n6861), .B(n7046), .Z(n6865) );
  XOR U845 ( .A(n6391), .B(n6574), .Z(n6399) );
  XOR U846 ( .A(n5375), .B(n5558), .Z(n5379) );
  XOR U847 ( .A(n5632), .B(n5824), .Z(n5627) );
  XOR U848 ( .A(n5083), .B(n5296), .Z(n5091) );
  XOR U849 ( .A(n4508), .B(n4745), .Z(n4512) );
  XOR U850 ( .A(n4783), .B(n5029), .Z(n4778) );
  XOR U851 ( .A(n4195), .B(n4465), .Z(n4203) );
  XOR U852 ( .A(n3584), .B(n3876), .Z(n3588) );
  XOR U853 ( .A(n4827), .B(n5017), .Z(n4831) );
  XOR U854 ( .A(n8867), .B(n9034), .Z(n8871) );
  XOR U855 ( .A(n8514), .B(n8682), .Z(n8518) );
  XOR U856 ( .A(n8148), .B(n8309), .Z(n8143) );
  XOR U857 ( .A(n7745), .B(n7910), .Z(n7749) );
  XOR U858 ( .A(n7320), .B(n7488), .Z(n7324) );
  XOR U859 ( .A(n6880), .B(n7043), .Z(n6875) );
  XOR U860 ( .A(n6405), .B(n6570), .Z(n6409) );
  XOR U861 ( .A(n5909), .B(n6075), .Z(n5913) );
  XOR U862 ( .A(n5394), .B(n5555), .Z(n5389) );
  XOR U863 ( .A(n4846), .B(n5011), .Z(n4850) );
  XOR U864 ( .A(n2955), .B(n3264), .Z(n2959) );
  XOR U865 ( .A(n4527), .B(n4742), .Z(n4522) );
  XOR U866 ( .A(n3299), .B(n3566), .Z(n3303) );
  XOR U867 ( .A(n3946), .B(n4159), .Z(n3950) );
  XOR U868 ( .A(n3618), .B(n3868), .Z(n3622) );
  XOR U869 ( .A(n3603), .B(n3873), .Z(n3598) );
  XOR U870 ( .A(n4556), .B(n4735), .Z(n4551) );
  XOR U871 ( .A(n9210), .B(n9357), .Z(n9214) );
  XOR U872 ( .A(n8714), .B(n8857), .Z(n8709) );
  XOR U873 ( .A(n8348), .B(n8491), .Z(n8352) );
  XOR U874 ( .A(n7962), .B(n8109), .Z(n7966) );
  XOR U875 ( .A(n7556), .B(n7699), .Z(n7551) );
  XOR U876 ( .A(n7118), .B(n7261), .Z(n7122) );
  XOR U877 ( .A(n6658), .B(n6805), .Z(n6662) );
  XOR U878 ( .A(n6180), .B(n6323), .Z(n6175) );
  XOR U879 ( .A(n5666), .B(n5813), .Z(n5670) );
  XOR U880 ( .A(n5136), .B(n5283), .Z(n5140) );
  XOR U881 ( .A(n4277), .B(n4445), .Z(n4281) );
  XOR U882 ( .A(n3666), .B(n3856), .Z(n3670) );
  XOR U883 ( .A(n2970), .B(n3261), .Z(n2978) );
  XOR U884 ( .A(n2308), .B(n2626), .Z(n2312) );
  XOR U885 ( .A(n9055), .B(n9196), .Z(n9063) );
  XOR U886 ( .A(n4585), .B(n4728), .Z(n4580) );
  XOR U887 ( .A(n2667), .B(n2941), .Z(n2671) );
  XOR U888 ( .A(n3652), .B(n3860), .Z(n3660) );
  XOR U889 ( .A(n3018), .B(n3249), .Z(n3022) );
  XOR U890 ( .A(n3695), .B(n3849), .Z(n3699) );
  XOR U891 ( .A(n3323), .B(n3562), .Z(n3318) );
  XOR U892 ( .A(n2361), .B(n2612), .Z(n2365) );
  XOR U893 ( .A(n9804), .B(n9933), .Z(n9808) );
  XOR U894 ( .A(n9523), .B(n9655), .Z(n9527) );
  XOR U895 ( .A(n8896), .B(n9027), .Z(n8900) );
  XOR U896 ( .A(n8543), .B(n8675), .Z(n8547) );
  XOR U897 ( .A(n8177), .B(n8302), .Z(n8172) );
  XOR U898 ( .A(n7774), .B(n7903), .Z(n7778) );
  XOR U899 ( .A(n7349), .B(n7481), .Z(n7353) );
  XOR U900 ( .A(n6909), .B(n7036), .Z(n6904) );
  XOR U901 ( .A(n6434), .B(n6563), .Z(n6438) );
  XOR U902 ( .A(n5938), .B(n6068), .Z(n5942) );
  XOR U903 ( .A(n5423), .B(n5548), .Z(n5418) );
  XOR U904 ( .A(n4875), .B(n5004), .Z(n4879) );
  XOR U905 ( .A(n4306), .B(n4438), .Z(n4310) );
  XOR U906 ( .A(n3681), .B(n3853), .Z(n3689) );
  XOR U907 ( .A(n3047), .B(n3242), .Z(n3051) );
  XOR U908 ( .A(n1659), .B(n1957), .Z(n1663) );
  XOR U909 ( .A(n2327), .B(n2623), .Z(n2322) );
  XOR U910 ( .A(n932), .B(n1279), .Z(n936) );
  XOR U911 ( .A(n9388), .B(n9503), .Z(n9383) );
  XOR U912 ( .A(n2390), .B(n2605), .Z(n2394) );
  XOR U913 ( .A(n2347), .B(n2616), .Z(n2355) );
  XOR U914 ( .A(n1645), .B(n1961), .Z(n1653) );
  XOR U915 ( .A(n3037), .B(n3246), .Z(n3032) );
  XOR U916 ( .A(n3710), .B(n3846), .Z(n3718) );
  XOR U917 ( .A(n3076), .B(n3235), .Z(n3080) );
  XOR U918 ( .A(n2376), .B(n2609), .Z(n2384) );
  XOR U919 ( .A(n2419), .B(n2598), .Z(n2423) );
  XOR U920 ( .A(n10073), .B(n10184), .Z(n10077) );
  XOR U921 ( .A(n9819), .B(n9930), .Z(n9827) );
  XOR U922 ( .A(n9239), .B(n9350), .Z(n9243) );
  XOR U923 ( .A(n8911), .B(n9024), .Z(n8919) );
  XOR U924 ( .A(n8377), .B(n8484), .Z(n8381) );
  XOR U925 ( .A(n7991), .B(n8102), .Z(n7995) );
  XOR U926 ( .A(n7585), .B(n7692), .Z(n7580) );
  XOR U927 ( .A(n7147), .B(n7254), .Z(n7151) );
  XOR U928 ( .A(n6687), .B(n6798), .Z(n6691) );
  XOR U929 ( .A(n6209), .B(n6316), .Z(n6204) );
  XOR U930 ( .A(n5695), .B(n5806), .Z(n5699) );
  XOR U931 ( .A(n5165), .B(n5276), .Z(n5169) );
  XOR U932 ( .A(n4614), .B(n4721), .Z(n4609) );
  XOR U933 ( .A(n3105), .B(n3228), .Z(n3109) );
  XOR U934 ( .A(n3066), .B(n3239), .Z(n3061) );
  XOR U935 ( .A(n1324), .B(n1615), .Z(n1328) );
  XOR U936 ( .A(n604), .B(n919), .Z(n608) );
  XOR U937 ( .A(n585), .B(n924), .Z(n589) );
  XOR U938 ( .A(n9690), .B(n9792), .Z(n9691) );
  XOR U939 ( .A(n8746), .B(n8848), .Z(n8747) );
  XOR U940 ( .A(n4325), .B(n4433), .Z(n4329) );
  XOR U941 ( .A(n2448), .B(n2591), .Z(n2452) );
  XOR U942 ( .A(n2405), .B(n2602), .Z(n2413) );
  XOR U943 ( .A(n1683), .B(n1953), .Z(n1678) );
  XOR U944 ( .A(n956), .B(n1275), .Z(n951) );
  XOR U945 ( .A(n1353), .B(n1608), .Z(n1357) );
  XOR U946 ( .A(n633), .B(n912), .Z(n637) );
  XOR U947 ( .A(n3095), .B(n3232), .Z(n3090) );
  XOR U948 ( .A(n1712), .B(n1946), .Z(n1707) );
  XOR U949 ( .A(n2434), .B(n2595), .Z(n2442) );
  XOR U950 ( .A(n10314), .B(n10412), .Z(n10318) );
  XOR U951 ( .A(n10092), .B(n10181), .Z(n10087) );
  XOR U952 ( .A(n9552), .B(n9648), .Z(n9556) );
  XOR U953 ( .A(n9258), .B(n9347), .Z(n9253) );
  XOR U954 ( .A(n8572), .B(n8668), .Z(n8576) );
  XOR U955 ( .A(n8206), .B(n8295), .Z(n8201) );
  XOR U956 ( .A(n7595), .B(n7688), .Z(n7599) );
  XOR U957 ( .A(n7162), .B(n7251), .Z(n7170) );
  XOR U958 ( .A(n6704), .B(n6794), .Z(n6705) );
  XOR U959 ( .A(n6219), .B(n6312), .Z(n6223) );
  XOR U960 ( .A(n5710), .B(n5803), .Z(n5718) );
  XOR U961 ( .A(n5182), .B(n5272), .Z(n5183) );
  XOR U962 ( .A(n4043), .B(n4136), .Z(n4051) );
  XOR U963 ( .A(n2812), .B(n2905), .Z(n2816) );
  XOR U964 ( .A(n3124), .B(n3225), .Z(n3119) );
  XOR U965 ( .A(n1382), .B(n1601), .Z(n1386) );
  XOR U966 ( .A(n662), .B(n905), .Z(n666) );
  XOR U967 ( .A(n619), .B(n916), .Z(n627) );
  XOR U968 ( .A(n2144), .B(n2255), .Z(n2148) );
  XOR U969 ( .A(n10624), .B(n10711), .Z(n10628) );
  XOR U970 ( .A(n9968), .B(n10055), .Z(n9972) );
  XOR U971 ( .A(n9098), .B(n9185), .Z(n9102) );
  XOR U972 ( .A(n8010), .B(n8097), .Z(n8014) );
  XOR U973 ( .A(n4909), .B(n4996), .Z(n4913) );
  XOR U974 ( .A(n2463), .B(n2588), .Z(n2471) );
  XOR U975 ( .A(n1741), .B(n1939), .Z(n1736) );
  XOR U976 ( .A(n648), .B(n909), .Z(n656) );
  XOR U977 ( .A(n1411), .B(n1594), .Z(n1415) );
  XOR U978 ( .A(n691), .B(n898), .Z(n695) );
  XOR U979 ( .A(n1770), .B(n1932), .Z(n1765) );
  XOR U980 ( .A(n1104), .B(n1238), .Z(n1105) );
  XOR U981 ( .A(n10540), .B(n10615), .Z(n10548) );
  XOR U982 ( .A(n10331), .B(n10408), .Z(n10332) );
  XOR U983 ( .A(n9848), .B(n9923), .Z(n9856) );
  XOR U984 ( .A(n9569), .B(n9644), .Z(n9570) );
  XOR U985 ( .A(n8940), .B(n9017), .Z(n8948) );
  XOR U986 ( .A(n8589), .B(n8664), .Z(n8590) );
  XOR U987 ( .A(n7818), .B(n7893), .Z(n7826) );
  XOR U988 ( .A(n7395), .B(n7470), .Z(n7396) );
  XOR U989 ( .A(n6716), .B(n6791), .Z(n6720) );
  XOR U990 ( .A(n6238), .B(n6309), .Z(n6233) );
  XOR U991 ( .A(n5724), .B(n5799), .Z(n5728) );
  XOR U992 ( .A(n4352), .B(n4427), .Z(n4353) );
  XOR U993 ( .A(n3758), .B(n3833), .Z(n3762) );
  XOR U994 ( .A(n3144), .B(n3219), .Z(n3148) );
  XOR U995 ( .A(n2502), .B(n2578), .Z(n2506) );
  XOR U996 ( .A(n1440), .B(n1587), .Z(n1444) );
  XOR U997 ( .A(n720), .B(n891), .Z(n724) );
  XOR U998 ( .A(n677), .B(n902), .Z(n685) );
  XOR U999 ( .A(n1814), .B(n1920), .Z(n1818) );
  XOR U1000 ( .A(n1839), .B(n1914), .Z(n1843) );
  XOR U1001 ( .A(n10809), .B(n10874), .Z(n10813) );
  XOR U1002 ( .A(n10225), .B(n10290), .Z(n10229) );
  XOR U1003 ( .A(n9427), .B(n9492), .Z(n9431) );
  XOR U1004 ( .A(n8411), .B(n8476), .Z(n8415) );
  XOR U1005 ( .A(n7181), .B(n7246), .Z(n7185) );
  XOR U1006 ( .A(n5467), .B(n5536), .Z(n5471) );
  XOR U1007 ( .A(n1799), .B(n1925), .Z(n1794) );
  XOR U1008 ( .A(n706), .B(n895), .Z(n714) );
  XOR U1009 ( .A(n5208), .B(n5267), .Z(n5203) );
  XOR U1010 ( .A(n754), .B(n883), .Z(n758) );
  XOR U1011 ( .A(n11028), .B(n11085), .Z(n11032) );
  XOR U1012 ( .A(n10741), .B(n10794), .Z(n10736) );
  XOR U1013 ( .A(n10554), .B(n10611), .Z(n10558) );
  XOR U1014 ( .A(n10121), .B(n10174), .Z(n10116) );
  XOR U1015 ( .A(n9862), .B(n9919), .Z(n9866) );
  XOR U1016 ( .A(n9287), .B(n9340), .Z(n9282) );
  XOR U1017 ( .A(n8954), .B(n9013), .Z(n8958) );
  XOR U1018 ( .A(n8235), .B(n8288), .Z(n8230) );
  XOR U1019 ( .A(n7832), .B(n7889), .Z(n7836) );
  XOR U1020 ( .A(n6967), .B(n7022), .Z(n6962) );
  XOR U1021 ( .A(n6492), .B(n6549), .Z(n6496) );
  XOR U1022 ( .A(n4653), .B(n4710), .Z(n4657) );
  XOR U1023 ( .A(n4072), .B(n4129), .Z(n4076) );
  XOR U1024 ( .A(n3469), .B(n3526), .Z(n3473) );
  XOR U1025 ( .A(n2842), .B(n2899), .Z(n2846) );
  XOR U1026 ( .A(n2189), .B(n2246), .Z(n2193) );
  XOR U1027 ( .A(n1514), .B(n1571), .Z(n1518) );
  XOR U1028 ( .A(n735), .B(n888), .Z(n743) );
  XOR U1029 ( .A(n1121), .B(n1234), .Z(n1125) );
  XOR U1030 ( .A(n784), .B(n877), .Z(n788) );
  XOR U1031 ( .A(n10969), .B(n11020), .Z(n10973) );
  XOR U1032 ( .A(n10459), .B(n10510), .Z(n10463) );
  XOR U1033 ( .A(n9731), .B(n9782), .Z(n9735) );
  XOR U1034 ( .A(n8787), .B(n8838), .Z(n8791) );
  XOR U1035 ( .A(n7629), .B(n7680), .Z(n7633) );
  XOR U1036 ( .A(n6253), .B(n6304), .Z(n6257) );
  XOR U1037 ( .A(n1151), .B(n1228), .Z(n1155) );
  XOR U1038 ( .A(n5751), .B(n5793), .Z(n5752) );
  XOR U1039 ( .A(n814), .B(n871), .Z(n818) );
  XOR U1040 ( .A(n10908), .B(n10947), .Z(n10909) );
  XOR U1041 ( .A(n10751), .B(n10790), .Z(n10755) );
  XOR U1042 ( .A(n10360), .B(n10401), .Z(n10361) );
  XOR U1043 ( .A(n10131), .B(n10170), .Z(n10135) );
  XOR U1044 ( .A(n9598), .B(n9637), .Z(n9599) );
  XOR U1045 ( .A(n9297), .B(n9336), .Z(n9301) );
  XOR U1046 ( .A(n8618), .B(n8657), .Z(n8619) );
  XOR U1047 ( .A(n8245), .B(n8284), .Z(n8249) );
  XOR U1048 ( .A(n7424), .B(n7463), .Z(n7425) );
  XOR U1049 ( .A(n6977), .B(n7018), .Z(n6981) );
  XOR U1050 ( .A(n5491), .B(n5530), .Z(n5495) );
  XOR U1051 ( .A(n4948), .B(n4987), .Z(n4952) );
  XOR U1052 ( .A(n4379), .B(n4421), .Z(n4383) );
  XOR U1053 ( .A(n3788), .B(n3827), .Z(n3792) );
  XOR U1054 ( .A(n3174), .B(n3213), .Z(n3178) );
  XOR U1055 ( .A(n2532), .B(n2572), .Z(n2536) );
  XOR U1056 ( .A(n1869), .B(n1908), .Z(n1873) );
  XOR U1057 ( .A(n1181), .B(n1222), .Z(n1185) );
  XOR U1058 ( .A(n11255), .B(n11287), .Z(n11259) );
  XNOR U1059 ( .A(n11261), .B(n11219), .Z(n11221) );
  XOR U1060 ( .A(n11106), .B(n11140), .Z(n11114) );
  XOR U1061 ( .A(n10668), .B(n10701), .Z(n10676) );
  XOR U1062 ( .A(n10012), .B(n10045), .Z(n10020) );
  XOR U1063 ( .A(n9142), .B(n9175), .Z(n9150) );
  XOR U1064 ( .A(n8054), .B(n8087), .Z(n8062) );
  XOR U1065 ( .A(n6750), .B(n6783), .Z(n6758) );
  XOR U1066 ( .A(n6519), .B(n6543), .Z(n6520) );
  XOR U1067 ( .A(n11057), .B(n11078), .Z(n11061) );
  XOR U1068 ( .A(n10920), .B(n10944), .Z(n10924) );
  XOR U1069 ( .A(n10583), .B(n10604), .Z(n10587) );
  XOR U1070 ( .A(n10372), .B(n10398), .Z(n10376) );
  XOR U1071 ( .A(n9891), .B(n9912), .Z(n9895) );
  XOR U1072 ( .A(n9610), .B(n9634), .Z(n9614) );
  XOR U1073 ( .A(n8983), .B(n9006), .Z(n8987) );
  XOR U1074 ( .A(n8630), .B(n8654), .Z(n8634) );
  XOR U1075 ( .A(n7861), .B(n7882), .Z(n7865) );
  XOR U1076 ( .A(n7436), .B(n7460), .Z(n7440) );
  XOR U1077 ( .A(n6277), .B(n6298), .Z(n6281) );
  XOR U1078 ( .A(n5238), .B(n5259), .Z(n5242) );
  XOR U1079 ( .A(n4683), .B(n4704), .Z(n4687) );
  XOR U1080 ( .A(n3499), .B(n3520), .Z(n3503) );
  XOR U1081 ( .A(n2872), .B(n2893), .Z(n2876) );
  XOR U1082 ( .A(n1544), .B(n1565), .Z(n1548) );
  XOR U1083 ( .A(n844), .B(n865), .Z(n848) );
  XOR U1084 ( .A(n11351), .B(n11356), .Z(n11340) );
  XNOR U1085 ( .A(n11334), .B(n11333), .Z(n11314) );
  XNOR U1086 ( .A(n11307), .B(n11306), .Z(n11281) );
  XOR U1087 ( .A(n11270), .B(n11275), .Z(n11241) );
  XOR U1088 ( .A(n11231), .B(n11236), .Z(n11191) );
  XOR U1089 ( .A(n11168), .B(n11186), .Z(n11178) );
  XOR U1090 ( .A(n10857), .B(n10864), .Z(n10851) );
  XOR U1091 ( .A(n10273), .B(n10280), .Z(n10267) );
  XOR U1092 ( .A(n9475), .B(n9482), .Z(n9469) );
  XOR U1093 ( .A(n8459), .B(n8466), .Z(n8453) );
  XOR U1094 ( .A(n7229), .B(n7236), .Z(n7223) );
  XNOR U1095 ( .A(n6030), .B(n6046), .Z(n6038) );
  XNOR U1096 ( .A(n4399), .B(n4417), .Z(n4407) );
  XNOR U1097 ( .A(n2552), .B(n2568), .Z(n2560) );
  XOR U1098 ( .A(n6590), .B(n6821), .Z(n6594) );
  XOR U1099 ( .A(n6103), .B(n6340), .Z(n6107) );
  XOR U1100 ( .A(n5579), .B(n5835), .Z(n5583) );
  XOR U1101 ( .A(n7065), .B(n7274), .Z(n7069) );
  XOR U1102 ( .A(n6605), .B(n6818), .Z(n6613) );
  XOR U1103 ( .A(n5870), .B(n6084), .Z(n5874) );
  XOR U1104 ( .A(n6122), .B(n6337), .Z(n6117) );
  XOR U1105 ( .A(n5594), .B(n5832), .Z(n5602) );
  XOR U1106 ( .A(n5044), .B(n5305), .Z(n5048) );
  XOR U1107 ( .A(n7721), .B(n7916), .Z(n7725) );
  XOR U1108 ( .A(n7296), .B(n7494), .Z(n7304) );
  XOR U1109 ( .A(n6854), .B(n7048), .Z(n6855) );
  XOR U1110 ( .A(n6381), .B(n6576), .Z(n6385) );
  XOR U1111 ( .A(n5885), .B(n6081), .Z(n5893) );
  XOR U1112 ( .A(n5346), .B(n5565), .Z(n5350) );
  XOR U1113 ( .A(n4474), .B(n4753), .Z(n4478) );
  XOR U1114 ( .A(n4788), .B(n5026), .Z(n4792) );
  XOR U1115 ( .A(n5063), .B(n5302), .Z(n5058) );
  XOR U1116 ( .A(n8504), .B(n8684), .Z(n8508) );
  XOR U1117 ( .A(n8134), .B(n8311), .Z(n8138) );
  XOR U1118 ( .A(n7740), .B(n7913), .Z(n7735) );
  XOR U1119 ( .A(n7310), .B(n7490), .Z(n7314) );
  XOR U1120 ( .A(n6866), .B(n7045), .Z(n6870) );
  XOR U1121 ( .A(n6400), .B(n6573), .Z(n6395) );
  XOR U1122 ( .A(n5899), .B(n6077), .Z(n5903) );
  XOR U1123 ( .A(n5365), .B(n5562), .Z(n5360) );
  XOR U1124 ( .A(n4489), .B(n4750), .Z(n4497) );
  XOR U1125 ( .A(n3888), .B(n4173), .Z(n3892) );
  XOR U1126 ( .A(n5107), .B(n5290), .Z(n5111) );
  XOR U1127 ( .A(n4803), .B(n5023), .Z(n4811) );
  XOR U1128 ( .A(n4214), .B(n4460), .Z(n4218) );
  XOR U1129 ( .A(n3270), .B(n3573), .Z(n3274) );
  XOR U1130 ( .A(n4537), .B(n4738), .Z(n4541) );
  XOR U1131 ( .A(n3608), .B(n3870), .Z(n3612) );
  XOR U1132 ( .A(n8872), .B(n9033), .Z(n8876) );
  XOR U1133 ( .A(n8519), .B(n8681), .Z(n8527) );
  XOR U1134 ( .A(n8151), .B(n8307), .Z(n8152) );
  XOR U1135 ( .A(n7750), .B(n7909), .Z(n7754) );
  XOR U1136 ( .A(n7325), .B(n7487), .Z(n7333) );
  XOR U1137 ( .A(n6883), .B(n7041), .Z(n6884) );
  XOR U1138 ( .A(n6410), .B(n6569), .Z(n6414) );
  XOR U1139 ( .A(n5914), .B(n6074), .Z(n5922) );
  XOR U1140 ( .A(n5397), .B(n5553), .Z(n5398) );
  XOR U1141 ( .A(n4851), .B(n5010), .Z(n4855) );
  XOR U1142 ( .A(n3907), .B(n4170), .Z(n3902) );
  XOR U1143 ( .A(n4841), .B(n5015), .Z(n4836) );
  XOR U1144 ( .A(n3637), .B(n3863), .Z(n3641) );
  XOR U1145 ( .A(n4233), .B(n4457), .Z(n4228) );
  XOR U1146 ( .A(n3285), .B(n3570), .Z(n3293) );
  XOR U1147 ( .A(n2638), .B(n2948), .Z(n2642) );
  XOR U1148 ( .A(n4253), .B(n4451), .Z(n4261) );
  XOR U1149 ( .A(n3975), .B(n4152), .Z(n3979) );
  XOR U1150 ( .A(n3623), .B(n3867), .Z(n3631) );
  XOR U1151 ( .A(n2989), .B(n3256), .Z(n2993) );
  XOR U1152 ( .A(n1970), .B(n2297), .Z(n1974) );
  XOR U1153 ( .A(n9369), .B(n9506), .Z(n9373) );
  XOR U1154 ( .A(n8891), .B(n9030), .Z(n8886) );
  XOR U1155 ( .A(n8533), .B(n8677), .Z(n8537) );
  XOR U1156 ( .A(n8163), .B(n8304), .Z(n8167) );
  XOR U1157 ( .A(n7769), .B(n7906), .Z(n7764) );
  XOR U1158 ( .A(n7339), .B(n7483), .Z(n7343) );
  XOR U1159 ( .A(n6895), .B(n7038), .Z(n6899) );
  XOR U1160 ( .A(n6429), .B(n6566), .Z(n6424) );
  XOR U1161 ( .A(n5928), .B(n6070), .Z(n5932) );
  XOR U1162 ( .A(n5409), .B(n5550), .Z(n5413) );
  XOR U1163 ( .A(n4588), .B(n4726), .Z(n4589) );
  XOR U1164 ( .A(n4282), .B(n4444), .Z(n4290) );
  XOR U1165 ( .A(n3338), .B(n3557), .Z(n3342) );
  XOR U1166 ( .A(n2691), .B(n2935), .Z(n2695) );
  XOR U1167 ( .A(n9220), .B(n9355), .Z(n9228) );
  XOR U1168 ( .A(n4301), .B(n4439), .Z(n4305) );
  XOR U1169 ( .A(n2657), .B(n2945), .Z(n2652) );
  XOR U1170 ( .A(n3661), .B(n3859), .Z(n3656) );
  XOR U1171 ( .A(n3367), .B(n3550), .Z(n3371) );
  XOR U1172 ( .A(n2720), .B(n2928), .Z(n2724) );
  XOR U1173 ( .A(n3008), .B(n3253), .Z(n3003) );
  XOR U1174 ( .A(n2342), .B(n2617), .Z(n2346) );
  XOR U1175 ( .A(n1985), .B(n2294), .Z(n1993) );
  XOR U1176 ( .A(n1290), .B(n1623), .Z(n1294) );
  XOR U1177 ( .A(n9939), .B(n10062), .Z(n9943) );
  XOR U1178 ( .A(n9673), .B(n9796), .Z(n9677) );
  XOR U1179 ( .A(n9069), .B(n9192), .Z(n9073) );
  XOR U1180 ( .A(n8729), .B(n8852), .Z(n8733) );
  XOR U1181 ( .A(n8372), .B(n8487), .Z(n8367) );
  XOR U1182 ( .A(n7981), .B(n8104), .Z(n7985) );
  XOR U1183 ( .A(n7571), .B(n7694), .Z(n7575) );
  XOR U1184 ( .A(n7142), .B(n7257), .Z(n7137) );
  XOR U1185 ( .A(n6677), .B(n6800), .Z(n6681) );
  XOR U1186 ( .A(n6195), .B(n6318), .Z(n6199) );
  XOR U1187 ( .A(n5690), .B(n5809), .Z(n5685) );
  XOR U1188 ( .A(n5155), .B(n5278), .Z(n5159) );
  XOR U1189 ( .A(n3690), .B(n3852), .Z(n3685) );
  XOR U1190 ( .A(n1664), .B(n1956), .Z(n1668) );
  XOR U1191 ( .A(n575), .B(n926), .Z(n579) );
  XOR U1192 ( .A(n2706), .B(n2932), .Z(n2714) );
  XOR U1193 ( .A(n2033), .B(n2282), .Z(n2037) );
  XOR U1194 ( .A(n3396), .B(n3543), .Z(n3400) );
  XOR U1195 ( .A(n2749), .B(n2921), .Z(n2753) );
  XOR U1196 ( .A(n9537), .B(n9653), .Z(n9532) );
  XOR U1197 ( .A(n4605), .B(n4722), .Z(n4613) );
  XOR U1198 ( .A(n3420), .B(n3537), .Z(n3424) );
  XOR U1199 ( .A(n1343), .B(n1610), .Z(n1347) );
  XOR U1200 ( .A(n3719), .B(n3845), .Z(n3714) );
  XOR U1201 ( .A(n2778), .B(n2914), .Z(n2782) );
  XOR U1202 ( .A(n2735), .B(n2925), .Z(n2743) );
  XOR U1203 ( .A(n2062), .B(n2275), .Z(n2066) );
  XOR U1204 ( .A(n2023), .B(n2286), .Z(n2018) );
  XOR U1205 ( .A(n1309), .B(n1620), .Z(n1304) );
  XOR U1206 ( .A(n10196), .B(n10297), .Z(n10200) );
  XOR U1207 ( .A(n9954), .B(n10059), .Z(n9962) );
  XOR U1208 ( .A(n9398), .B(n9499), .Z(n9402) );
  XOR U1209 ( .A(n9084), .B(n9189), .Z(n9092) );
  XOR U1210 ( .A(n8562), .B(n8670), .Z(n8566) );
  XOR U1211 ( .A(n8192), .B(n8297), .Z(n8196) );
  XOR U1212 ( .A(n7798), .B(n7899), .Z(n7793) );
  XOR U1213 ( .A(n7368), .B(n7476), .Z(n7372) );
  XOR U1214 ( .A(n6924), .B(n7031), .Z(n6928) );
  XOR U1215 ( .A(n6458), .B(n6559), .Z(n6453) );
  XOR U1216 ( .A(n5957), .B(n6063), .Z(n5961) );
  XOR U1217 ( .A(n5438), .B(n5543), .Z(n5442) );
  XOR U1218 ( .A(n1372), .B(n1603), .Z(n1376) );
  XOR U1219 ( .A(n1329), .B(n1614), .Z(n1337) );
  XOR U1220 ( .A(n609), .B(n918), .Z(n613) );
  XOR U1221 ( .A(n590), .B(n923), .Z(n598) );
  XOR U1222 ( .A(n2052), .B(n2279), .Z(n2047) );
  XOR U1223 ( .A(n2764), .B(n2918), .Z(n2772) );
  XOR U1224 ( .A(n2091), .B(n2268), .Z(n2095) );
  XOR U1225 ( .A(n9831), .B(n9927), .Z(n9832) );
  XOR U1226 ( .A(n8923), .B(n9021), .Z(n8924) );
  XOR U1227 ( .A(n5179), .B(n5274), .Z(n5174) );
  XOR U1228 ( .A(n4619), .B(n4718), .Z(n4623) );
  XOR U1229 ( .A(n4038), .B(n4137), .Z(n4042) );
  XOR U1230 ( .A(n1358), .B(n1607), .Z(n1366) );
  XOR U1231 ( .A(n638), .B(n911), .Z(n642) );
  XOR U1232 ( .A(n1401), .B(n1596), .Z(n1405) );
  XOR U1233 ( .A(n2477), .B(n2583), .Z(n2481) );
  XOR U1234 ( .A(n10525), .B(n10618), .Z(n10529) );
  XOR U1235 ( .A(n2793), .B(n2911), .Z(n2801) );
  XOR U1236 ( .A(n2120), .B(n2261), .Z(n2124) );
  XOR U1237 ( .A(n2081), .B(n2272), .Z(n2076) );
  XOR U1238 ( .A(n10430), .B(n10517), .Z(n10434) );
  XOR U1239 ( .A(n10215), .B(n10294), .Z(n10210) );
  XOR U1240 ( .A(n9702), .B(n9789), .Z(n9706) );
  XOR U1241 ( .A(n9417), .B(n9496), .Z(n9412) );
  XOR U1242 ( .A(n8758), .B(n8845), .Z(n8762) );
  XOR U1243 ( .A(n8401), .B(n8480), .Z(n8396) );
  XOR U1244 ( .A(n7808), .B(n7895), .Z(n7812) );
  XOR U1245 ( .A(n7383), .B(n7473), .Z(n7391) );
  XOR U1246 ( .A(n6941), .B(n7027), .Z(n6942) );
  XOR U1247 ( .A(n6468), .B(n6555), .Z(n6472) );
  XOR U1248 ( .A(n5972), .B(n6060), .Z(n5980) );
  XOR U1249 ( .A(n3751), .B(n3835), .Z(n3752) );
  XOR U1250 ( .A(n3134), .B(n3221), .Z(n3138) );
  XOR U1251 ( .A(n1430), .B(n1589), .Z(n1434) );
  XOR U1252 ( .A(n1387), .B(n1600), .Z(n1395) );
  XOR U1253 ( .A(n667), .B(n904), .Z(n671) );
  XOR U1254 ( .A(n628), .B(n915), .Z(n623) );
  XOR U1255 ( .A(n2110), .B(n2265), .Z(n2105) );
  XOR U1256 ( .A(n10097), .B(n10178), .Z(n10101) );
  XOR U1257 ( .A(n9263), .B(n9344), .Z(n9267) );
  XOR U1258 ( .A(n8211), .B(n8292), .Z(n8215) );
  XOR U1259 ( .A(n5722), .B(n5800), .Z(n5723) );
  XOR U1260 ( .A(n5189), .B(n5270), .Z(n5193) );
  XOR U1261 ( .A(n4634), .B(n4715), .Z(n4642) );
  XOR U1262 ( .A(n657), .B(n908), .Z(n652) );
  XOR U1263 ( .A(n1416), .B(n1593), .Z(n1424) );
  XOR U1264 ( .A(n696), .B(n897), .Z(n700) );
  XOR U1265 ( .A(n2492), .B(n2580), .Z(n2496) );
  XOR U1266 ( .A(n1809), .B(n1921), .Z(n1813) );
  XOR U1267 ( .A(n10722), .B(n10797), .Z(n10726) );
  XOR U1268 ( .A(n2139), .B(n2258), .Z(n2134) );
  XOR U1269 ( .A(n1106), .B(n1237), .Z(n1110) );
  XOR U1270 ( .A(n1489), .B(n1576), .Z(n1493) );
  XOR U1271 ( .A(n10639), .B(n10708), .Z(n10647) );
  XOR U1272 ( .A(n10447), .B(n10513), .Z(n10448) );
  XOR U1273 ( .A(n9983), .B(n10052), .Z(n9991) );
  XOR U1274 ( .A(n9719), .B(n9785), .Z(n9720) );
  XOR U1275 ( .A(n9113), .B(n9182), .Z(n9121) );
  XOR U1276 ( .A(n8775), .B(n8841), .Z(n8776) );
  XOR U1277 ( .A(n8025), .B(n8094), .Z(n8033) );
  XOR U1278 ( .A(n7617), .B(n7683), .Z(n7618) );
  XOR U1279 ( .A(n6953), .B(n7024), .Z(n6957) );
  XOR U1280 ( .A(n6487), .B(n6552), .Z(n6482) );
  XOR U1281 ( .A(n4354), .B(n4426), .Z(n4358) );
  XOR U1282 ( .A(n3763), .B(n3832), .Z(n3767) );
  XOR U1283 ( .A(n2507), .B(n2577), .Z(n2511) );
  XOR U1284 ( .A(n1445), .B(n1586), .Z(n1453) );
  XOR U1285 ( .A(n725), .B(n890), .Z(n729) );
  XOR U1286 ( .A(n686), .B(n901), .Z(n681) );
  XOR U1287 ( .A(n774), .B(n879), .Z(n778) );
  XOR U1288 ( .A(n10338), .B(n10406), .Z(n10342) );
  XOR U1289 ( .A(n9576), .B(n9642), .Z(n9580) );
  XOR U1290 ( .A(n8596), .B(n8662), .Z(n8600) );
  XOR U1291 ( .A(n7402), .B(n7468), .Z(n7406) );
  XOR U1292 ( .A(n5991), .B(n6055), .Z(n5995) );
  XOR U1293 ( .A(n5472), .B(n5535), .Z(n5480) );
  XOR U1294 ( .A(n4931), .B(n4991), .Z(n4932) );
  XOR U1295 ( .A(n3154), .B(n3217), .Z(n3158) );
  XOR U1296 ( .A(n715), .B(n894), .Z(n710) );
  XOR U1297 ( .A(n1474), .B(n1579), .Z(n1478) );
  XOR U1298 ( .A(n10891), .B(n10951), .Z(n10895) );
  XOR U1299 ( .A(n759), .B(n882), .Z(n763) );
  XOR U1300 ( .A(n1504), .B(n1573), .Z(n1508) );
  XOR U1301 ( .A(n804), .B(n873), .Z(n808) );
  XOR U1302 ( .A(n11091), .B(n11143), .Z(n11095) );
  XOR U1303 ( .A(n10828), .B(n10871), .Z(n10823) );
  XOR U1304 ( .A(n10653), .B(n10704), .Z(n10657) );
  XOR U1305 ( .A(n10244), .B(n10287), .Z(n10239) );
  XOR U1306 ( .A(n9997), .B(n10048), .Z(n10001) );
  XOR U1307 ( .A(n9446), .B(n9489), .Z(n9441) );
  XOR U1308 ( .A(n9127), .B(n9178), .Z(n9131) );
  XOR U1309 ( .A(n8430), .B(n8473), .Z(n8425) );
  XOR U1310 ( .A(n8039), .B(n8090), .Z(n8043) );
  XOR U1311 ( .A(n7200), .B(n7243), .Z(n7195) );
  XOR U1312 ( .A(n6735), .B(n6786), .Z(n6739) );
  XOR U1313 ( .A(n4658), .B(n4709), .Z(n4662) );
  XOR U1314 ( .A(n4077), .B(n4128), .Z(n4081) );
  XOR U1315 ( .A(n2847), .B(n2898), .Z(n2851) );
  XOR U1316 ( .A(n2194), .B(n2245), .Z(n2198) );
  XOR U1317 ( .A(n744), .B(n887), .Z(n739) );
  XOR U1318 ( .A(n789), .B(n876), .Z(n793) );
  XOR U1319 ( .A(n10564), .B(n10609), .Z(n10568) );
  XOR U1320 ( .A(n9872), .B(n9917), .Z(n9876) );
  XOR U1321 ( .A(n8964), .B(n9011), .Z(n8968) );
  XOR U1322 ( .A(n7842), .B(n7887), .Z(n7846) );
  XOR U1323 ( .A(n6258), .B(n6303), .Z(n6266) );
  XOR U1324 ( .A(n5486), .B(n5531), .Z(n5490) );
  XOR U1325 ( .A(n3783), .B(n3828), .Z(n3787) );
  XOR U1326 ( .A(n1864), .B(n1909), .Z(n1868) );
  XOR U1327 ( .A(n11043), .B(n11082), .Z(n11051) );
  XOR U1328 ( .A(n6013), .B(n6050), .Z(n6014) );
  XOR U1329 ( .A(n819), .B(n870), .Z(n823) );
  XNOR U1330 ( .A(n11294), .B(n11258), .Z(n11260) );
  XOR U1331 ( .A(n11216), .B(n11248), .Z(n11220) );
  XOR U1332 ( .A(n10986), .B(n11016), .Z(n10987) );
  XOR U1333 ( .A(n10838), .B(n10867), .Z(n10842) );
  XOR U1334 ( .A(n10476), .B(n10506), .Z(n10477) );
  XOR U1335 ( .A(n10254), .B(n10283), .Z(n10258) );
  XOR U1336 ( .A(n9748), .B(n9778), .Z(n9749) );
  XOR U1337 ( .A(n9456), .B(n9485), .Z(n9460) );
  XOR U1338 ( .A(n8804), .B(n8834), .Z(n8805) );
  XOR U1339 ( .A(n8440), .B(n8469), .Z(n8444) );
  XOR U1340 ( .A(n7646), .B(n7676), .Z(n7647) );
  XOR U1341 ( .A(n7210), .B(n7239), .Z(n7214) );
  XOR U1342 ( .A(n5228), .B(n5261), .Z(n5232) );
  XOR U1343 ( .A(n4673), .B(n4706), .Z(n4677) );
  XOR U1344 ( .A(n3489), .B(n3522), .Z(n3493) );
  XOR U1345 ( .A(n2862), .B(n2895), .Z(n2866) );
  XOR U1346 ( .A(n1534), .B(n1567), .Z(n1538) );
  XOR U1347 ( .A(n834), .B(n867), .Z(n838) );
  XOR U1348 ( .A(n10761), .B(n10788), .Z(n10769) );
  XOR U1349 ( .A(n10141), .B(n10168), .Z(n10149) );
  XOR U1350 ( .A(n9307), .B(n9334), .Z(n9315) );
  XOR U1351 ( .A(n8255), .B(n8282), .Z(n8263) );
  XOR U1352 ( .A(n6987), .B(n7016), .Z(n6995) );
  XOR U1353 ( .A(n5763), .B(n5790), .Z(n5767) );
  XOR U1354 ( .A(n4097), .B(n4124), .Z(n4101) );
  XOR U1355 ( .A(n2214), .B(n2241), .Z(n2218) );
  XOR U1356 ( .A(n11173), .B(n11196), .Z(n11167) );
  XOR U1357 ( .A(n6762), .B(n6780), .Z(n6763) );
  XNOR U1358 ( .A(n11355), .B(n11354), .Z(n11341) );
  XOR U1359 ( .A(n11330), .B(n11335), .Z(n11313) );
  XOR U1360 ( .A(n11303), .B(n11308), .Z(n11280) );
  XNOR U1361 ( .A(n11274), .B(n11273), .Z(n11242) );
  XOR U1362 ( .A(n11120), .B(n11135), .Z(n11129) );
  XOR U1363 ( .A(n10998), .B(n11013), .Z(n11007) );
  XOR U1364 ( .A(n10682), .B(n10697), .Z(n10691) );
  XOR U1365 ( .A(n10488), .B(n10503), .Z(n10497) );
  XOR U1366 ( .A(n10026), .B(n10041), .Z(n10035) );
  XOR U1367 ( .A(n9760), .B(n9775), .Z(n9769) );
  XOR U1368 ( .A(n9156), .B(n9171), .Z(n9165) );
  XOR U1369 ( .A(n8816), .B(n8831), .Z(n8825) );
  XOR U1370 ( .A(n8068), .B(n8083), .Z(n8077) );
  XOR U1371 ( .A(n7658), .B(n7673), .Z(n7667) );
  XOR U1372 ( .A(n6526), .B(n6541), .Z(n6535) );
  XOR U1373 ( .A(n5511), .B(n5526), .Z(n5520) );
  XOR U1374 ( .A(n4968), .B(n4983), .Z(n4977) );
  XOR U1375 ( .A(n3808), .B(n3823), .Z(n3817) );
  XOR U1376 ( .A(n3194), .B(n3209), .Z(n3203) );
  XOR U1377 ( .A(n1889), .B(n1904), .Z(n1898) );
  XOR U1378 ( .A(n1201), .B(n1218), .Z(n1210) );
  XNOR U1379 ( .A(n11192), .B(n11189), .Z(n11181) );
  XNOR U1380 ( .A(n10929), .B(n10939), .Z(n10937) );
  XNOR U1381 ( .A(n10381), .B(n10393), .Z(n10389) );
  XNOR U1382 ( .A(n9619), .B(n9629), .Z(n9627) );
  XNOR U1383 ( .A(n8639), .B(n8649), .Z(n8647) );
  XNOR U1384 ( .A(n7445), .B(n7455), .Z(n7453) );
  XOR U1385 ( .A(n6038), .B(n6042), .Z(n6034) );
  XOR U1386 ( .A(n4407), .B(n4413), .Z(n4403) );
  XOR U1387 ( .A(n2560), .B(n2564), .Z(n2556) );
  XOR U1388 ( .A(n6098), .B(n6341), .Z(n6102) );
  XOR U1389 ( .A(n7281), .B(n7497), .Z(n7285) );
  XOR U1390 ( .A(n6837), .B(n7052), .Z(n6841) );
  XOR U1391 ( .A(n6113), .B(n6338), .Z(n6121) );
  XOR U1392 ( .A(n5584), .B(n5834), .Z(n5588) );
  XOR U1393 ( .A(n5039), .B(n5306), .Z(n5043) );
  XOR U1394 ( .A(n5341), .B(n5566), .Z(n5345) );
  XOR U1395 ( .A(n7923), .B(n8118), .Z(n7927) );
  XOR U1396 ( .A(n7513), .B(n7708), .Z(n7517) );
  XOR U1397 ( .A(n7084), .B(n7271), .Z(n7079) );
  XOR U1398 ( .A(n6619), .B(n6814), .Z(n6623) );
  XOR U1399 ( .A(n6137), .B(n6332), .Z(n6141) );
  XOR U1400 ( .A(n5603), .B(n5831), .Z(n5598) );
  XOR U1401 ( .A(n5054), .B(n5303), .Z(n5062) );
  XOR U1402 ( .A(n4479), .B(n4752), .Z(n4483) );
  XOR U1403 ( .A(n5097), .B(n5292), .Z(n5101) );
  XOR U1404 ( .A(n5356), .B(n5563), .Z(n5364) );
  XOR U1405 ( .A(n4793), .B(n5025), .Z(n4797) );
  XOR U1406 ( .A(n3883), .B(n4174), .Z(n3887) );
  XOR U1407 ( .A(n8324), .B(n8497), .Z(n8328) );
  XOR U1408 ( .A(n7938), .B(n8115), .Z(n7946) );
  XOR U1409 ( .A(n7530), .B(n7704), .Z(n7531) );
  XOR U1410 ( .A(n7094), .B(n7267), .Z(n7098) );
  XOR U1411 ( .A(n6634), .B(n6811), .Z(n6642) );
  XOR U1412 ( .A(n6154), .B(n6328), .Z(n6155) );
  XOR U1413 ( .A(n5642), .B(n5819), .Z(n5646) );
  XOR U1414 ( .A(n4209), .B(n4461), .Z(n4213) );
  XOR U1415 ( .A(n4498), .B(n4749), .Z(n4493) );
  XOR U1416 ( .A(n5112), .B(n5289), .Z(n5120) );
  XOR U1417 ( .A(n4812), .B(n5022), .Z(n4807) );
  XOR U1418 ( .A(n3898), .B(n4171), .Z(n3906) );
  XOR U1419 ( .A(n3275), .B(n3572), .Z(n3279) );
  XOR U1420 ( .A(n4542), .B(n4737), .Z(n4546) );
  XOR U1421 ( .A(n3941), .B(n4160), .Z(n3945) );
  XOR U1422 ( .A(n9040), .B(n9199), .Z(n9044) );
  XOR U1423 ( .A(n8700), .B(n8859), .Z(n8704) );
  XOR U1424 ( .A(n8343), .B(n8494), .Z(n8338) );
  XOR U1425 ( .A(n7952), .B(n8111), .Z(n7956) );
  XOR U1426 ( .A(n7542), .B(n7701), .Z(n7546) );
  XOR U1427 ( .A(n7113), .B(n7264), .Z(n7108) );
  XOR U1428 ( .A(n6648), .B(n6807), .Z(n6652) );
  XOR U1429 ( .A(n6166), .B(n6325), .Z(n6170) );
  XOR U1430 ( .A(n5661), .B(n5816), .Z(n5656) );
  XOR U1431 ( .A(n5126), .B(n5285), .Z(n5130) );
  XOR U1432 ( .A(n4224), .B(n4458), .Z(n4232) );
  XOR U1433 ( .A(n3613), .B(n3869), .Z(n3617) );
  XOR U1434 ( .A(n2633), .B(n2949), .Z(n2637) );
  XOR U1435 ( .A(n4571), .B(n4730), .Z(n4575) );
  XOR U1436 ( .A(n3970), .B(n4153), .Z(n3974) );
  XOR U1437 ( .A(n2984), .B(n3257), .Z(n2988) );
  XOR U1438 ( .A(n3294), .B(n3569), .Z(n3289) );
  XOR U1439 ( .A(n4262), .B(n4450), .Z(n4257) );
  XOR U1440 ( .A(n3647), .B(n3861), .Z(n3651) );
  XOR U1441 ( .A(n3013), .B(n3250), .Z(n3017) );
  XOR U1442 ( .A(n3999), .B(n4146), .Z(n4003) );
  XOR U1443 ( .A(n9513), .B(n9657), .Z(n9517) );
  XOR U1444 ( .A(n9215), .B(n9356), .Z(n9219) );
  XOR U1445 ( .A(n8717), .B(n8855), .Z(n8718) );
  XOR U1446 ( .A(n8353), .B(n8490), .Z(n8357) );
  XOR U1447 ( .A(n7967), .B(n8108), .Z(n7975) );
  XOR U1448 ( .A(n7559), .B(n7697), .Z(n7560) );
  XOR U1449 ( .A(n7123), .B(n7260), .Z(n7127) );
  XOR U1450 ( .A(n6663), .B(n6804), .Z(n6671) );
  XOR U1451 ( .A(n6183), .B(n6321), .Z(n6184) );
  XOR U1452 ( .A(n5671), .B(n5812), .Z(n5675) );
  XOR U1453 ( .A(n5141), .B(n5282), .Z(n5149) );
  XOR U1454 ( .A(n3632), .B(n3866), .Z(n3627) );
  XOR U1455 ( .A(n2648), .B(n2946), .Z(n2656) );
  XOR U1456 ( .A(n1975), .B(n2296), .Z(n1979) );
  XOR U1457 ( .A(n9064), .B(n9195), .Z(n9059) );
  XOR U1458 ( .A(n4291), .B(n4443), .Z(n4286) );
  XOR U1459 ( .A(n3676), .B(n3854), .Z(n3680) );
  XOR U1460 ( .A(n3042), .B(n3243), .Z(n3046) );
  XOR U1461 ( .A(n2999), .B(n3254), .Z(n3007) );
  XOR U1462 ( .A(n2337), .B(n2618), .Z(n2341) );
  XOR U1463 ( .A(n1285), .B(n1624), .Z(n1289) );
  XOR U1464 ( .A(n3352), .B(n3555), .Z(n3347) );
  XOR U1465 ( .A(n2701), .B(n2933), .Z(n2705) );
  XOR U1466 ( .A(n2028), .B(n2283), .Z(n2032) );
  XOR U1467 ( .A(n3705), .B(n3847), .Z(n3709) );
  XOR U1468 ( .A(n3071), .B(n3236), .Z(n3075) );
  XOR U1469 ( .A(n9809), .B(n9932), .Z(n9813) );
  XOR U1470 ( .A(n9528), .B(n9654), .Z(n9536) );
  XOR U1471 ( .A(n8901), .B(n9026), .Z(n8905) );
  XOR U1472 ( .A(n8548), .B(n8674), .Z(n8556) );
  XOR U1473 ( .A(n8180), .B(n8300), .Z(n8181) );
  XOR U1474 ( .A(n7779), .B(n7902), .Z(n7783) );
  XOR U1475 ( .A(n7354), .B(n7480), .Z(n7362) );
  XOR U1476 ( .A(n6912), .B(n7034), .Z(n6913) );
  XOR U1477 ( .A(n6439), .B(n6562), .Z(n6443) );
  XOR U1478 ( .A(n5943), .B(n6067), .Z(n5951) );
  XOR U1479 ( .A(n5426), .B(n5546), .Z(n5427) );
  XOR U1480 ( .A(n4880), .B(n5003), .Z(n4884) );
  XOR U1481 ( .A(n4311), .B(n4437), .Z(n4319) );
  XOR U1482 ( .A(n1994), .B(n2293), .Z(n1989) );
  XOR U1483 ( .A(n9391), .B(n9501), .Z(n9392) );
  XOR U1484 ( .A(n3100), .B(n3229), .Z(n3104) );
  XOR U1485 ( .A(n3381), .B(n3548), .Z(n3376) );
  XOR U1486 ( .A(n2730), .B(n2926), .Z(n2734) );
  XOR U1487 ( .A(n2057), .B(n2276), .Z(n2061) );
  XOR U1488 ( .A(n2356), .B(n2615), .Z(n2351) );
  XOR U1489 ( .A(n1669), .B(n1955), .Z(n1673) );
  XOR U1490 ( .A(n961), .B(n1272), .Z(n965) );
  XOR U1491 ( .A(n1300), .B(n1621), .Z(n1308) );
  XOR U1492 ( .A(n580), .B(n925), .Z(n584) );
  XOR U1493 ( .A(n2385), .B(n2608), .Z(n2380) );
  XOR U1494 ( .A(n1698), .B(n1948), .Z(n1702) );
  XOR U1495 ( .A(n990), .B(n1265), .Z(n994) );
  XOR U1496 ( .A(n3410), .B(n3541), .Z(n3405) );
  XOR U1497 ( .A(n2759), .B(n2919), .Z(n2763) );
  XOR U1498 ( .A(n2086), .B(n2269), .Z(n2090) );
  XOR U1499 ( .A(n10078), .B(n10183), .Z(n10082) );
  XOR U1500 ( .A(n9828), .B(n9929), .Z(n9823) );
  XOR U1501 ( .A(n9244), .B(n9349), .Z(n9248) );
  XOR U1502 ( .A(n8920), .B(n9023), .Z(n8915) );
  XOR U1503 ( .A(n8382), .B(n8483), .Z(n8386) );
  XOR U1504 ( .A(n7996), .B(n8101), .Z(n8004) );
  XOR U1505 ( .A(n7588), .B(n7690), .Z(n7589) );
  XOR U1506 ( .A(n7152), .B(n7253), .Z(n7156) );
  XOR U1507 ( .A(n6692), .B(n6797), .Z(n6700) );
  XOR U1508 ( .A(n6212), .B(n6314), .Z(n6213) );
  XOR U1509 ( .A(n5700), .B(n5805), .Z(n5704) );
  XOR U1510 ( .A(n5170), .B(n5275), .Z(n5178) );
  XOR U1511 ( .A(n4617), .B(n4719), .Z(n4618) );
  XOR U1512 ( .A(n4033), .B(n4138), .Z(n4037) );
  XOR U1513 ( .A(n3430), .B(n3535), .Z(n3438) );
  XOR U1514 ( .A(n10420), .B(n10519), .Z(n10424) );
  XOR U1515 ( .A(n9692), .B(n9791), .Z(n9696) );
  XOR U1516 ( .A(n8748), .B(n8847), .Z(n8752) );
  XOR U1517 ( .A(n2788), .B(n2912), .Z(n2792) );
  XOR U1518 ( .A(n2115), .B(n2262), .Z(n2119) );
  XOR U1519 ( .A(n2414), .B(n2601), .Z(n2409) );
  XOR U1520 ( .A(n1727), .B(n1941), .Z(n1731) );
  XOR U1521 ( .A(n1019), .B(n1258), .Z(n1023) );
  XOR U1522 ( .A(n1338), .B(n1613), .Z(n1333) );
  XOR U1523 ( .A(n614), .B(n917), .Z(n618) );
  XOR U1524 ( .A(n599), .B(n922), .Z(n594) );
  XOR U1525 ( .A(n1367), .B(n1606), .Z(n1362) );
  XOR U1526 ( .A(n643), .B(n910), .Z(n647) );
  XOR U1527 ( .A(n2443), .B(n2594), .Z(n2438) );
  XOR U1528 ( .A(n1756), .B(n1934), .Z(n1760) );
  XOR U1529 ( .A(n1048), .B(n1251), .Z(n1052) );
  XOR U1530 ( .A(n10319), .B(n10411), .Z(n10327) );
  XOR U1531 ( .A(n10095), .B(n10179), .Z(n10096) );
  XOR U1532 ( .A(n9557), .B(n9647), .Z(n9565) );
  XOR U1533 ( .A(n9261), .B(n9345), .Z(n9262) );
  XOR U1534 ( .A(n8577), .B(n8667), .Z(n8585) );
  XOR U1535 ( .A(n8209), .B(n8293), .Z(n8210) );
  XOR U1536 ( .A(n7600), .B(n7687), .Z(n7604) );
  XOR U1537 ( .A(n7171), .B(n7250), .Z(n7166) );
  XOR U1538 ( .A(n6706), .B(n6793), .Z(n6710) );
  XOR U1539 ( .A(n6224), .B(n6311), .Z(n6228) );
  XOR U1540 ( .A(n5719), .B(n5802), .Z(n5714) );
  XOR U1541 ( .A(n5184), .B(n5271), .Z(n5188) );
  XOR U1542 ( .A(n4629), .B(n4716), .Z(n4633) );
  XOR U1543 ( .A(n4052), .B(n4135), .Z(n4047) );
  XOR U1544 ( .A(n3444), .B(n3531), .Z(n3448) );
  XOR U1545 ( .A(n2817), .B(n2904), .Z(n2821) );
  XOR U1546 ( .A(n1804), .B(n1922), .Z(n1808) );
  XOR U1547 ( .A(n10629), .B(n10710), .Z(n10633) );
  XOR U1548 ( .A(n9973), .B(n10054), .Z(n9977) );
  XOR U1549 ( .A(n9103), .B(n9184), .Z(n9107) );
  XOR U1550 ( .A(n8015), .B(n8096), .Z(n8019) );
  XOR U1551 ( .A(n2472), .B(n2587), .Z(n2467) );
  XOR U1552 ( .A(n1785), .B(n1927), .Z(n1789) );
  XOR U1553 ( .A(n1077), .B(n1244), .Z(n1081) );
  XOR U1554 ( .A(n1396), .B(n1599), .Z(n1391) );
  XOR U1555 ( .A(n672), .B(n903), .Z(n676) );
  XOR U1556 ( .A(n252), .B(n531), .Z(n282) );
  XOR U1557 ( .A(n1484), .B(n1577), .Z(n1488) );
  XOR U1558 ( .A(n236), .B(n512), .Z(n292) );
  XOR U1559 ( .A(n1425), .B(n1592), .Z(n1420) );
  XOR U1560 ( .A(n701), .B(n896), .Z(n705) );
  XOR U1561 ( .A(n2159), .B(n2252), .Z(n2163) );
  XOR U1562 ( .A(n10549), .B(n10614), .Z(n10544) );
  XOR U1563 ( .A(n10333), .B(n10407), .Z(n10337) );
  XOR U1564 ( .A(n9857), .B(n9922), .Z(n9852) );
  XOR U1565 ( .A(n9571), .B(n9643), .Z(n9575) );
  XOR U1566 ( .A(n8949), .B(n9016), .Z(n8944) );
  XOR U1567 ( .A(n8591), .B(n8663), .Z(n8595) );
  XOR U1568 ( .A(n7827), .B(n7892), .Z(n7822) );
  XOR U1569 ( .A(n7397), .B(n7469), .Z(n7401) );
  XOR U1570 ( .A(n6721), .B(n6790), .Z(n6729) );
  XOR U1571 ( .A(n6241), .B(n6307), .Z(n6242) );
  XOR U1572 ( .A(n5729), .B(n5798), .Z(n5733) );
  XOR U1573 ( .A(n5199), .B(n5268), .Z(n5207) );
  XOR U1574 ( .A(n4646), .B(n4712), .Z(n4647) );
  XOR U1575 ( .A(n4062), .B(n4131), .Z(n4066) );
  XOR U1576 ( .A(n3459), .B(n3528), .Z(n3463) );
  XOR U1577 ( .A(n2832), .B(n2901), .Z(n2836) );
  XOR U1578 ( .A(n2179), .B(n2248), .Z(n2183) );
  XOR U1579 ( .A(n1469), .B(n1580), .Z(n1473) );
  XOR U1580 ( .A(n749), .B(n884), .Z(n753) );
  XOR U1581 ( .A(n10959), .B(n11022), .Z(n10963) );
  XOR U1582 ( .A(n10814), .B(n10873), .Z(n10818) );
  XOR U1583 ( .A(n10230), .B(n10289), .Z(n10234) );
  XOR U1584 ( .A(n9432), .B(n9491), .Z(n9436) );
  XOR U1585 ( .A(n8416), .B(n8475), .Z(n8420) );
  XOR U1586 ( .A(n7186), .B(n7245), .Z(n7190) );
  XOR U1587 ( .A(n1454), .B(n1585), .Z(n1449) );
  XOR U1588 ( .A(n730), .B(n889), .Z(n734) );
  XOR U1589 ( .A(n220), .B(n493), .Z(n302) );
  XOR U1590 ( .A(n1499), .B(n1574), .Z(n1503) );
  XOR U1591 ( .A(n779), .B(n878), .Z(n783) );
  XOR U1592 ( .A(n204), .B(n474), .Z(n312) );
  XOR U1593 ( .A(n10744), .B(n10792), .Z(n10745) );
  XOR U1594 ( .A(n10559), .B(n10610), .Z(n10563) );
  XOR U1595 ( .A(n10124), .B(n10172), .Z(n10125) );
  XOR U1596 ( .A(n9867), .B(n9918), .Z(n9871) );
  XOR U1597 ( .A(n9290), .B(n9338), .Z(n9291) );
  XOR U1598 ( .A(n8959), .B(n9012), .Z(n8963) );
  XOR U1599 ( .A(n8238), .B(n8286), .Z(n8239) );
  XOR U1600 ( .A(n7837), .B(n7888), .Z(n7841) );
  XOR U1601 ( .A(n6970), .B(n7020), .Z(n6971) );
  XOR U1602 ( .A(n6497), .B(n6548), .Z(n6501) );
  XOR U1603 ( .A(n6001), .B(n6053), .Z(n6009) );
  XOR U1604 ( .A(n5484), .B(n5532), .Z(n5485) );
  XOR U1605 ( .A(n4938), .B(n4989), .Z(n4942) );
  XOR U1606 ( .A(n4369), .B(n4423), .Z(n4373) );
  XOR U1607 ( .A(n3778), .B(n3829), .Z(n3782) );
  XOR U1608 ( .A(n3164), .B(n3215), .Z(n3168) );
  XOR U1609 ( .A(n2522), .B(n2574), .Z(n2526) );
  XOR U1610 ( .A(n1859), .B(n1910), .Z(n1863) );
  XOR U1611 ( .A(n764), .B(n881), .Z(n768) );
  XOR U1612 ( .A(n809), .B(n872), .Z(n813) );
  XOR U1613 ( .A(n11096), .B(n11142), .Z(n11100) );
  XOR U1614 ( .A(n10974), .B(n11019), .Z(n10982) );
  XOR U1615 ( .A(n10464), .B(n10509), .Z(n10472) );
  XOR U1616 ( .A(n9736), .B(n9781), .Z(n9744) );
  XOR U1617 ( .A(n8792), .B(n8837), .Z(n8800) );
  XOR U1618 ( .A(n7634), .B(n7679), .Z(n7642) );
  XOR U1619 ( .A(n188), .B(n455), .Z(n322) );
  XOR U1620 ( .A(n794), .B(n875), .Z(n798) );
  XOR U1621 ( .A(n10910), .B(n10946), .Z(n10914) );
  XOR U1622 ( .A(n10756), .B(n10789), .Z(n10760) );
  XOR U1623 ( .A(n10362), .B(n10400), .Z(n10366) );
  XOR U1624 ( .A(n10136), .B(n10169), .Z(n10140) );
  XOR U1625 ( .A(n9600), .B(n9636), .Z(n9604) );
  XOR U1626 ( .A(n9302), .B(n9335), .Z(n9306) );
  XOR U1627 ( .A(n8620), .B(n8656), .Z(n8624) );
  XOR U1628 ( .A(n8250), .B(n8283), .Z(n8254) );
  XOR U1629 ( .A(n7426), .B(n7462), .Z(n7430) );
  XOR U1630 ( .A(n6982), .B(n7017), .Z(n6986) );
  XOR U1631 ( .A(n6516), .B(n6545), .Z(n6511) );
  XOR U1632 ( .A(n6015), .B(n6049), .Z(n6019) );
  XOR U1633 ( .A(n5496), .B(n5529), .Z(n5500) );
  XOR U1634 ( .A(n4953), .B(n4986), .Z(n4957) );
  XOR U1635 ( .A(n4384), .B(n4420), .Z(n4388) );
  XOR U1636 ( .A(n3793), .B(n3826), .Z(n3797) );
  XOR U1637 ( .A(n3179), .B(n3212), .Z(n3183) );
  XOR U1638 ( .A(n2537), .B(n2571), .Z(n2541) );
  XOR U1639 ( .A(n1874), .B(n1907), .Z(n1878) );
  XOR U1640 ( .A(n824), .B(n869), .Z(n828) );
  XNOR U1641 ( .A(n11326), .B(n11296), .Z(n11298) );
  XNOR U1642 ( .A(n11299), .B(n11263), .Z(n11265) );
  XOR U1643 ( .A(n11221), .B(n11247), .Z(n11225) );
  XOR U1644 ( .A(n11115), .B(n11139), .Z(n11109) );
  XOR U1645 ( .A(n10677), .B(n10700), .Z(n10672) );
  XOR U1646 ( .A(n10021), .B(n10044), .Z(n10016) );
  XOR U1647 ( .A(n9151), .B(n9174), .Z(n9146) );
  XOR U1648 ( .A(n8063), .B(n8086), .Z(n8058) );
  XOR U1649 ( .A(n11062), .B(n11077), .Z(n11071) );
  XNOR U1650 ( .A(n10925), .B(n10943), .Z(n10929) );
  XOR U1651 ( .A(n10588), .B(n10603), .Z(n10597) );
  XNOR U1652 ( .A(n10377), .B(n10397), .Z(n10381) );
  XOR U1653 ( .A(n9896), .B(n9911), .Z(n9905) );
  XNOR U1654 ( .A(n9615), .B(n9633), .Z(n9619) );
  XOR U1655 ( .A(n8988), .B(n9005), .Z(n8997) );
  XNOR U1656 ( .A(n8635), .B(n8653), .Z(n8639) );
  XOR U1657 ( .A(n7866), .B(n7881), .Z(n7875) );
  XNOR U1658 ( .A(n7441), .B(n7459), .Z(n7445) );
  XOR U1659 ( .A(n6764), .B(n6779), .Z(n6773) );
  XOR U1660 ( .A(n6282), .B(n6297), .Z(n6291) );
  XOR U1661 ( .A(n5773), .B(n5788), .Z(n5781) );
  XOR U1662 ( .A(n5243), .B(n5258), .Z(n5252) );
  XOR U1663 ( .A(n4688), .B(n4703), .Z(n4697) );
  XOR U1664 ( .A(n4107), .B(n4122), .Z(n4115) );
  XOR U1665 ( .A(n3504), .B(n3519), .Z(n3513) );
  XOR U1666 ( .A(n2877), .B(n2892), .Z(n2886) );
  XOR U1667 ( .A(n2224), .B(n2239), .Z(n2232) );
  XOR U1668 ( .A(n1549), .B(n1564), .Z(n1558) );
  XOR U1669 ( .A(n849), .B(n864), .Z(n858) );
  XNOR U1670 ( .A(n11362), .B(n11359), .Z(n11344) );
  XNOR U1671 ( .A(n11341), .B(n11338), .Z(n11317) );
  XNOR U1672 ( .A(n11314), .B(n11311), .Z(n11284) );
  XNOR U1673 ( .A(n11281), .B(n11278), .Z(n11245) );
  XNOR U1674 ( .A(n11242), .B(n11239), .Z(n11195) );
  XNOR U1675 ( .A(n11179), .B(n11177), .Z(n11134) );
  XOR U1676 ( .A(n10852), .B(n10863), .Z(n10860) );
  XOR U1677 ( .A(n10268), .B(n10279), .Z(n10276) );
  XOR U1678 ( .A(n9470), .B(n9481), .Z(n9478) );
  XOR U1679 ( .A(n8454), .B(n8465), .Z(n8462) );
  XOR U1680 ( .A(n7224), .B(n7235), .Z(n7232) );
  XNOR U1681 ( .A(n6034), .B(n6033), .Z(n5787) );
  XNOR U1682 ( .A(n4403), .B(n4402), .Z(n4121) );
  XNOR U1683 ( .A(n2556), .B(n2555), .Z(n2238) );
  XOR U1684 ( .A(n1), .B(n2), .Z(c[9]) );
  XNOR U1685 ( .A(n3), .B(n4), .Z(c[8]) );
  XNOR U1686 ( .A(n5), .B(n6), .Z(c[7]) );
  XNOR U1687 ( .A(n7), .B(n8), .Z(c[6]) );
  XOR U1688 ( .A(n9), .B(n10), .Z(c[63]) );
  XOR U1689 ( .A(n11), .B(n12), .Z(n10) );
  XOR U1690 ( .A(n13), .B(n14), .Z(n12) );
  XOR U1691 ( .A(n15), .B(n16), .Z(n14) );
  XOR U1692 ( .A(n17), .B(n18), .Z(n16) );
  XOR U1693 ( .A(n19), .B(n20), .Z(n18) );
  AND U1694 ( .A(b[3]), .B(a[60]), .Z(n20) );
  AND U1695 ( .A(b[4]), .B(a[59]), .Z(n19) );
  XOR U1696 ( .A(n21), .B(n22), .Z(n17) );
  XOR U1697 ( .A(n23), .B(n24), .Z(n22) );
  XOR U1698 ( .A(n25), .B(n26), .Z(n24) );
  AND U1699 ( .A(b[9]), .B(a[54]), .Z(n26) );
  AND U1700 ( .A(a[53]), .B(b[10]), .Z(n25) );
  XOR U1701 ( .A(n27), .B(n28), .Z(n23) );
  XOR U1702 ( .A(n29), .B(n30), .Z(n28) );
  XOR U1703 ( .A(n31), .B(n32), .Z(n30) );
  AND U1704 ( .A(b[15]), .B(a[48]), .Z(n32) );
  AND U1705 ( .A(a[47]), .B(b[16]), .Z(n31) );
  XOR U1706 ( .A(n33), .B(n34), .Z(n29) );
  XOR U1707 ( .A(n35), .B(n36), .Z(n34) );
  XOR U1708 ( .A(n37), .B(n38), .Z(n36) );
  AND U1709 ( .A(b[21]), .B(a[42]), .Z(n38) );
  AND U1710 ( .A(a[41]), .B(b[22]), .Z(n37) );
  XOR U1711 ( .A(n39), .B(n40), .Z(n35) );
  XOR U1712 ( .A(n41), .B(n42), .Z(n40) );
  XOR U1713 ( .A(n43), .B(n44), .Z(n42) );
  XOR U1714 ( .A(n45), .B(n46), .Z(n44) );
  XOR U1715 ( .A(n47), .B(n48), .Z(n46) );
  XOR U1716 ( .A(n49), .B(n50), .Z(n48) );
  XOR U1717 ( .A(n51), .B(n52), .Z(n50) );
  XOR U1718 ( .A(n53), .B(n54), .Z(n52) );
  XOR U1719 ( .A(n55), .B(n56), .Z(n54) );
  XOR U1720 ( .A(n57), .B(n58), .Z(n56) );
  XOR U1721 ( .A(n59), .B(n60), .Z(n58) );
  XOR U1722 ( .A(n61), .B(n62), .Z(n60) );
  AND U1723 ( .A(b[45]), .B(a[18]), .Z(n62) );
  AND U1724 ( .A(b[51]), .B(a[12]), .Z(n61) );
  XOR U1725 ( .A(n63), .B(n64), .Z(n59) );
  XOR U1726 ( .A(n65), .B(n66), .Z(n64) );
  XOR U1727 ( .A(n67), .B(n68), .Z(n66) );
  XOR U1728 ( .A(n69), .B(n70), .Z(n68) );
  AND U1729 ( .A(a[11]), .B(b[52]), .Z(n70) );
  AND U1730 ( .A(a[6]), .B(b[57]), .Z(n69) );
  XOR U1731 ( .A(n71), .B(n72), .Z(n67) );
  AND U1732 ( .A(a[5]), .B(b[58]), .Z(n72) );
  AND U1733 ( .A(a[4]), .B(b[59]), .Z(n71) );
  XOR U1734 ( .A(n73), .B(n74), .Z(n65) );
  XOR U1735 ( .A(n75), .B(n76), .Z(n74) );
  AND U1736 ( .A(a[3]), .B(b[60]), .Z(n76) );
  AND U1737 ( .A(a[2]), .B(b[61]), .Z(n75) );
  XOR U1738 ( .A(n77), .B(n78), .Z(n73) );
  AND U1739 ( .A(a[1]), .B(b[62]), .Z(n78) );
  AND U1740 ( .A(b[63]), .B(a[0]), .Z(n77) );
  AND U1741 ( .A(a[17]), .B(b[46]), .Z(n63) );
  XOR U1742 ( .A(n79), .B(n80), .Z(n57) );
  XOR U1743 ( .A(n81), .B(n82), .Z(n80) );
  AND U1744 ( .A(a[10]), .B(b[53]), .Z(n82) );
  AND U1745 ( .A(a[9]), .B(b[54]), .Z(n81) );
  XOR U1746 ( .A(n83), .B(n84), .Z(n79) );
  AND U1747 ( .A(a[8]), .B(b[55]), .Z(n84) );
  AND U1748 ( .A(a[7]), .B(b[56]), .Z(n83) );
  AND U1749 ( .A(a[23]), .B(b[40]), .Z(n55) );
  AND U1750 ( .A(b[39]), .B(a[24]), .Z(n53) );
  XOR U1751 ( .A(n85), .B(n86), .Z(n51) );
  XOR U1752 ( .A(n87), .B(n88), .Z(n86) );
  AND U1753 ( .A(a[16]), .B(b[47]), .Z(n88) );
  AND U1754 ( .A(a[15]), .B(b[48]), .Z(n87) );
  XOR U1755 ( .A(n89), .B(n90), .Z(n85) );
  AND U1756 ( .A(a[14]), .B(b[49]), .Z(n90) );
  AND U1757 ( .A(a[13]), .B(b[50]), .Z(n89) );
  AND U1758 ( .A(a[29]), .B(b[34]), .Z(n49) );
  AND U1759 ( .A(b[33]), .B(a[30]), .Z(n47) );
  XOR U1760 ( .A(n91), .B(n92), .Z(n45) );
  XOR U1761 ( .A(n93), .B(n94), .Z(n92) );
  AND U1762 ( .A(a[22]), .B(b[41]), .Z(n94) );
  AND U1763 ( .A(a[21]), .B(b[42]), .Z(n93) );
  XOR U1764 ( .A(n95), .B(n96), .Z(n91) );
  AND U1765 ( .A(a[20]), .B(b[43]), .Z(n96) );
  AND U1766 ( .A(a[19]), .B(b[44]), .Z(n95) );
  AND U1767 ( .A(a[35]), .B(b[28]), .Z(n43) );
  AND U1768 ( .A(b[27]), .B(a[36]), .Z(n41) );
  XOR U1769 ( .A(n97), .B(n98), .Z(n39) );
  XOR U1770 ( .A(n99), .B(n100), .Z(n98) );
  AND U1771 ( .A(a[28]), .B(b[35]), .Z(n100) );
  AND U1772 ( .A(a[27]), .B(b[36]), .Z(n99) );
  XOR U1773 ( .A(n101), .B(n102), .Z(n97) );
  AND U1774 ( .A(a[26]), .B(b[37]), .Z(n102) );
  AND U1775 ( .A(a[25]), .B(b[38]), .Z(n101) );
  XOR U1776 ( .A(n103), .B(n104), .Z(n33) );
  XOR U1777 ( .A(n105), .B(n106), .Z(n104) );
  AND U1778 ( .A(a[34]), .B(b[29]), .Z(n106) );
  AND U1779 ( .A(a[33]), .B(b[30]), .Z(n105) );
  XOR U1780 ( .A(n107), .B(n108), .Z(n103) );
  AND U1781 ( .A(a[32]), .B(b[31]), .Z(n108) );
  AND U1782 ( .A(a[31]), .B(b[32]), .Z(n107) );
  XOR U1783 ( .A(n109), .B(n110), .Z(n27) );
  XOR U1784 ( .A(n111), .B(n112), .Z(n110) );
  AND U1785 ( .A(a[40]), .B(b[23]), .Z(n112) );
  AND U1786 ( .A(a[39]), .B(b[24]), .Z(n111) );
  XOR U1787 ( .A(n113), .B(n114), .Z(n109) );
  AND U1788 ( .A(a[38]), .B(b[25]), .Z(n114) );
  AND U1789 ( .A(a[37]), .B(b[26]), .Z(n113) );
  XOR U1790 ( .A(n115), .B(n116), .Z(n21) );
  XOR U1791 ( .A(n117), .B(n118), .Z(n116) );
  AND U1792 ( .A(a[46]), .B(b[17]), .Z(n118) );
  AND U1793 ( .A(a[45]), .B(b[18]), .Z(n117) );
  XOR U1794 ( .A(n119), .B(n120), .Z(n115) );
  AND U1795 ( .A(a[44]), .B(b[19]), .Z(n120) );
  AND U1796 ( .A(a[43]), .B(b[20]), .Z(n119) );
  XOR U1797 ( .A(n121), .B(n122), .Z(n15) );
  XOR U1798 ( .A(n123), .B(n124), .Z(n122) );
  AND U1799 ( .A(a[52]), .B(b[11]), .Z(n124) );
  AND U1800 ( .A(a[51]), .B(b[12]), .Z(n123) );
  XOR U1801 ( .A(n125), .B(n126), .Z(n121) );
  AND U1802 ( .A(a[50]), .B(b[13]), .Z(n126) );
  AND U1803 ( .A(a[49]), .B(b[14]), .Z(n125) );
  AND U1804 ( .A(a[63]), .B(b[0]), .Z(n13) );
  XOR U1805 ( .A(n127), .B(n128), .Z(n11) );
  AND U1806 ( .A(b[1]), .B(a[62]), .Z(n128) );
  AND U1807 ( .A(b[2]), .B(a[61]), .Z(n127) );
  XOR U1808 ( .A(n129), .B(n130), .Z(n9) );
  XOR U1809 ( .A(n131), .B(n132), .Z(n130) );
  AND U1810 ( .A(b[5]), .B(a[58]), .Z(n132) );
  AND U1811 ( .A(b[6]), .B(a[57]), .Z(n131) );
  XOR U1812 ( .A(n133), .B(n134), .Z(n129) );
  AND U1813 ( .A(b[7]), .B(a[56]), .Z(n134) );
  AND U1814 ( .A(b[8]), .B(a[55]), .Z(n133) );
  XOR U1815 ( .A(n135), .B(n136), .Z(c[62]) );
  XOR U1816 ( .A(n137), .B(n138), .Z(n136) );
  XOR U1817 ( .A(n139), .B(n140), .Z(n138) );
  XOR U1818 ( .A(n141), .B(n142), .Z(n140) );
  XOR U1819 ( .A(n143), .B(n144), .Z(n142) );
  XOR U1820 ( .A(n145), .B(n146), .Z(n144) );
  AND U1821 ( .A(b[3]), .B(a[59]), .Z(n145) );
  XOR U1822 ( .A(n147), .B(n148), .Z(n143) );
  XOR U1823 ( .A(n149), .B(n150), .Z(n148) );
  XOR U1824 ( .A(n151), .B(n152), .Z(n150) );
  XOR U1825 ( .A(n153), .B(n154), .Z(n152) );
  AND U1826 ( .A(b[9]), .B(a[53]), .Z(n153) );
  XOR U1827 ( .A(n155), .B(n156), .Z(n151) );
  XOR U1828 ( .A(n157), .B(n158), .Z(n156) );
  XOR U1829 ( .A(n159), .B(n160), .Z(n158) );
  XOR U1830 ( .A(n161), .B(n162), .Z(n160) );
  AND U1831 ( .A(a[47]), .B(b[15]), .Z(n161) );
  XOR U1832 ( .A(n163), .B(n164), .Z(n159) );
  XOR U1833 ( .A(n165), .B(n166), .Z(n164) );
  XOR U1834 ( .A(n167), .B(n168), .Z(n166) );
  XOR U1835 ( .A(n169), .B(n167), .Z(n168) );
  AND U1836 ( .A(a[41]), .B(b[21]), .Z(n169) );
  XOR U1837 ( .A(n170), .B(n171), .Z(n167) );
  ANDN U1838 ( .B(n172), .A(n173), .Z(n170) );
  XOR U1839 ( .A(n174), .B(n175), .Z(n165) );
  XOR U1840 ( .A(n176), .B(n177), .Z(n175) );
  AND U1841 ( .A(b[26]), .B(a[36]), .Z(n176) );
  XOR U1842 ( .A(n177), .B(n178), .Z(n174) );
  XOR U1843 ( .A(n179), .B(n180), .Z(n178) );
  XOR U1844 ( .A(n181), .B(n182), .Z(n180) );
  XOR U1845 ( .A(n183), .B(n184), .Z(n182) );
  XOR U1846 ( .A(n185), .B(n183), .Z(n184) );
  AND U1847 ( .A(a[35]), .B(b[27]), .Z(n185) );
  XOR U1848 ( .A(n186), .B(n187), .Z(n183) );
  NOR U1849 ( .A(n188), .B(n189), .Z(n186) );
  XOR U1850 ( .A(n190), .B(n191), .Z(n181) );
  XOR U1851 ( .A(n192), .B(n193), .Z(n191) );
  AND U1852 ( .A(b[32]), .B(a[30]), .Z(n192) );
  XOR U1853 ( .A(n193), .B(n194), .Z(n190) );
  XOR U1854 ( .A(n195), .B(n196), .Z(n194) );
  XOR U1855 ( .A(n197), .B(n198), .Z(n196) );
  XOR U1856 ( .A(n199), .B(n200), .Z(n198) );
  XOR U1857 ( .A(n201), .B(n199), .Z(n200) );
  AND U1858 ( .A(a[29]), .B(b[33]), .Z(n201) );
  XOR U1859 ( .A(n202), .B(n203), .Z(n199) );
  NOR U1860 ( .A(n204), .B(n205), .Z(n202) );
  XOR U1861 ( .A(n206), .B(n207), .Z(n197) );
  XOR U1862 ( .A(n208), .B(n209), .Z(n207) );
  AND U1863 ( .A(b[38]), .B(a[24]), .Z(n208) );
  XOR U1864 ( .A(n209), .B(n210), .Z(n206) );
  XOR U1865 ( .A(n211), .B(n212), .Z(n210) );
  XOR U1866 ( .A(n213), .B(n214), .Z(n212) );
  XOR U1867 ( .A(n215), .B(n216), .Z(n214) );
  XOR U1868 ( .A(n217), .B(n215), .Z(n216) );
  AND U1869 ( .A(a[23]), .B(b[39]), .Z(n217) );
  XOR U1870 ( .A(n218), .B(n219), .Z(n215) );
  NOR U1871 ( .A(n220), .B(n221), .Z(n218) );
  XOR U1872 ( .A(n222), .B(n223), .Z(n213) );
  XOR U1873 ( .A(n224), .B(n225), .Z(n223) );
  AND U1874 ( .A(b[44]), .B(a[18]), .Z(n224) );
  XOR U1875 ( .A(n225), .B(n226), .Z(n222) );
  XOR U1876 ( .A(n227), .B(n228), .Z(n226) );
  XOR U1877 ( .A(n229), .B(n230), .Z(n228) );
  XOR U1878 ( .A(n231), .B(n232), .Z(n230) );
  XOR U1879 ( .A(n233), .B(n231), .Z(n232) );
  AND U1880 ( .A(a[17]), .B(b[45]), .Z(n233) );
  XOR U1881 ( .A(n234), .B(n235), .Z(n231) );
  NOR U1882 ( .A(n236), .B(n237), .Z(n234) );
  XOR U1883 ( .A(n238), .B(n239), .Z(n229) );
  XOR U1884 ( .A(n240), .B(n241), .Z(n239) );
  AND U1885 ( .A(b[50]), .B(a[12]), .Z(n240) );
  XOR U1886 ( .A(n241), .B(n242), .Z(n238) );
  XOR U1887 ( .A(n243), .B(n244), .Z(n242) );
  XOR U1888 ( .A(n245), .B(n246), .Z(n244) );
  XOR U1889 ( .A(n247), .B(n248), .Z(n246) );
  XOR U1890 ( .A(n249), .B(n247), .Z(n248) );
  AND U1891 ( .A(a[11]), .B(b[51]), .Z(n249) );
  XOR U1892 ( .A(n250), .B(n251), .Z(n247) );
  NOR U1893 ( .A(n252), .B(n253), .Z(n250) );
  XOR U1894 ( .A(n254), .B(n255), .Z(n245) );
  XOR U1895 ( .A(n256), .B(n257), .Z(n255) );
  AND U1896 ( .A(b[56]), .B(a[6]), .Z(n256) );
  XOR U1897 ( .A(n258), .B(n259), .Z(n254) );
  XOR U1898 ( .A(n257), .B(n260), .Z(n259) );
  XOR U1899 ( .A(n261), .B(n262), .Z(n260) );
  AND U1900 ( .A(b[57]), .B(a[5]), .Z(n262) );
  AND U1901 ( .A(b[58]), .B(a[4]), .Z(n261) );
  XOR U1902 ( .A(n263), .B(n264), .Z(n257) );
  ANDN U1903 ( .B(n265), .A(n266), .Z(n263) );
  XOR U1904 ( .A(n267), .B(n268), .Z(n258) );
  XOR U1905 ( .A(n269), .B(n270), .Z(n268) );
  AND U1906 ( .A(b[59]), .B(a[3]), .Z(n270) );
  AND U1907 ( .A(b[60]), .B(a[2]), .Z(n269) );
  XOR U1908 ( .A(n271), .B(n272), .Z(n267) );
  AND U1909 ( .A(b[61]), .B(a[1]), .Z(n272) );
  AND U1910 ( .A(b[62]), .B(a[0]), .Z(n271) );
  XOR U1911 ( .A(n273), .B(n274), .Z(n243) );
  XOR U1912 ( .A(n275), .B(n276), .Z(n274) );
  AND U1913 ( .A(b[52]), .B(a[10]), .Z(n276) );
  AND U1914 ( .A(b[53]), .B(a[9]), .Z(n275) );
  XOR U1915 ( .A(n277), .B(n278), .Z(n273) );
  AND U1916 ( .A(b[54]), .B(a[8]), .Z(n278) );
  AND U1917 ( .A(b[55]), .B(a[7]), .Z(n277) );
  XOR U1918 ( .A(n279), .B(n280), .Z(n241) );
  AND U1919 ( .A(n281), .B(n282), .Z(n279) );
  XOR U1920 ( .A(n283), .B(n284), .Z(n227) );
  XOR U1921 ( .A(n285), .B(n286), .Z(n284) );
  AND U1922 ( .A(a[16]), .B(b[46]), .Z(n286) );
  AND U1923 ( .A(a[15]), .B(b[47]), .Z(n285) );
  XOR U1924 ( .A(n287), .B(n288), .Z(n283) );
  AND U1925 ( .A(a[14]), .B(b[48]), .Z(n288) );
  AND U1926 ( .A(a[13]), .B(b[49]), .Z(n287) );
  XOR U1927 ( .A(n289), .B(n290), .Z(n225) );
  AND U1928 ( .A(n291), .B(n292), .Z(n289) );
  XOR U1929 ( .A(n293), .B(n294), .Z(n211) );
  XOR U1930 ( .A(n295), .B(n296), .Z(n294) );
  AND U1931 ( .A(a[22]), .B(b[40]), .Z(n296) );
  AND U1932 ( .A(a[21]), .B(b[41]), .Z(n295) );
  XOR U1933 ( .A(n297), .B(n298), .Z(n293) );
  AND U1934 ( .A(a[20]), .B(b[42]), .Z(n298) );
  AND U1935 ( .A(a[19]), .B(b[43]), .Z(n297) );
  XOR U1936 ( .A(n299), .B(n300), .Z(n209) );
  AND U1937 ( .A(n301), .B(n302), .Z(n299) );
  XOR U1938 ( .A(n303), .B(n304), .Z(n195) );
  XOR U1939 ( .A(n305), .B(n306), .Z(n304) );
  AND U1940 ( .A(a[28]), .B(b[34]), .Z(n306) );
  AND U1941 ( .A(a[27]), .B(b[35]), .Z(n305) );
  XOR U1942 ( .A(n307), .B(n308), .Z(n303) );
  AND U1943 ( .A(a[26]), .B(b[36]), .Z(n308) );
  AND U1944 ( .A(a[25]), .B(b[37]), .Z(n307) );
  XOR U1945 ( .A(n309), .B(n310), .Z(n193) );
  AND U1946 ( .A(n311), .B(n312), .Z(n309) );
  XOR U1947 ( .A(n313), .B(n314), .Z(n179) );
  XOR U1948 ( .A(n315), .B(n316), .Z(n314) );
  AND U1949 ( .A(a[34]), .B(b[28]), .Z(n316) );
  AND U1950 ( .A(a[33]), .B(b[29]), .Z(n315) );
  XOR U1951 ( .A(n317), .B(n318), .Z(n313) );
  AND U1952 ( .A(a[32]), .B(b[30]), .Z(n318) );
  AND U1953 ( .A(a[31]), .B(b[31]), .Z(n317) );
  XOR U1954 ( .A(n319), .B(n320), .Z(n177) );
  AND U1955 ( .A(n321), .B(n322), .Z(n319) );
  XOR U1956 ( .A(n323), .B(n324), .Z(n163) );
  XOR U1957 ( .A(n325), .B(n326), .Z(n324) );
  AND U1958 ( .A(a[40]), .B(b[22]), .Z(n326) );
  AND U1959 ( .A(a[39]), .B(b[23]), .Z(n325) );
  XOR U1960 ( .A(n327), .B(n328), .Z(n323) );
  AND U1961 ( .A(a[38]), .B(b[24]), .Z(n328) );
  AND U1962 ( .A(a[37]), .B(b[25]), .Z(n327) );
  XOR U1963 ( .A(n329), .B(n162), .Z(n157) );
  XOR U1964 ( .A(n330), .B(n331), .Z(n162) );
  ANDN U1965 ( .B(n332), .A(n333), .Z(n330) );
  AND U1966 ( .A(a[46]), .B(b[16]), .Z(n329) );
  XOR U1967 ( .A(n334), .B(n335), .Z(n155) );
  XOR U1968 ( .A(n336), .B(n337), .Z(n335) );
  AND U1969 ( .A(a[45]), .B(b[17]), .Z(n337) );
  AND U1970 ( .A(a[44]), .B(b[18]), .Z(n336) );
  XOR U1971 ( .A(n338), .B(n339), .Z(n334) );
  AND U1972 ( .A(a[43]), .B(b[19]), .Z(n339) );
  AND U1973 ( .A(b[20]), .B(a[42]), .Z(n338) );
  XOR U1974 ( .A(n340), .B(n154), .Z(n149) );
  XOR U1975 ( .A(n341), .B(n342), .Z(n154) );
  ANDN U1976 ( .B(n343), .A(n344), .Z(n341) );
  AND U1977 ( .A(a[52]), .B(b[10]), .Z(n340) );
  XOR U1978 ( .A(n345), .B(n346), .Z(n147) );
  XOR U1979 ( .A(n347), .B(n348), .Z(n346) );
  AND U1980 ( .A(a[51]), .B(b[11]), .Z(n348) );
  AND U1981 ( .A(a[50]), .B(b[12]), .Z(n347) );
  XOR U1982 ( .A(n349), .B(n350), .Z(n345) );
  AND U1983 ( .A(a[49]), .B(b[13]), .Z(n350) );
  AND U1984 ( .A(b[14]), .B(a[48]), .Z(n349) );
  XOR U1985 ( .A(n351), .B(n146), .Z(n141) );
  XNOR U1986 ( .A(n352), .B(n353), .Z(n146) );
  ANDN U1987 ( .B(n354), .A(n355), .Z(n352) );
  AND U1988 ( .A(b[4]), .B(a[58]), .Z(n351) );
  XOR U1989 ( .A(n356), .B(n357), .Z(n139) );
  XOR U1990 ( .A(n358), .B(n359), .Z(n357) );
  AND U1991 ( .A(b[5]), .B(a[57]), .Z(n359) );
  AND U1992 ( .A(b[6]), .B(a[56]), .Z(n358) );
  XOR U1993 ( .A(n360), .B(n361), .Z(n356) );
  AND U1994 ( .A(b[7]), .B(a[55]), .Z(n361) );
  AND U1995 ( .A(b[8]), .B(a[54]), .Z(n360) );
  AND U1996 ( .A(a[62]), .B(b[0]), .Z(n137) );
  XOR U1997 ( .A(n362), .B(n363), .Z(n135) );
  AND U1998 ( .A(b[1]), .B(a[61]), .Z(n363) );
  AND U1999 ( .A(b[2]), .B(a[60]), .Z(n362) );
  XOR U2000 ( .A(n364), .B(n365), .Z(c[61]) );
  XOR U2001 ( .A(n366), .B(n367), .Z(n365) );
  XNOR U2002 ( .A(n368), .B(n369), .Z(n367) );
  AND U2003 ( .A(b[1]), .B(a[60]), .Z(n369) );
  XNOR U2004 ( .A(n355), .B(n370), .Z(n366) );
  XNOR U2005 ( .A(n368), .B(n354), .Z(n370) );
  XNOR U2006 ( .A(n371), .B(n353), .Z(n354) );
  AND U2007 ( .A(b[2]), .B(a[59]), .Z(n371) );
  NANDN U2008 ( .A(n372), .B(n373), .Z(n368) );
  XOR U2009 ( .A(n374), .B(n375), .Z(n355) );
  XNOR U2010 ( .A(n353), .B(n376), .Z(n375) );
  XOR U2011 ( .A(n377), .B(n378), .Z(n376) );
  XOR U2012 ( .A(n379), .B(n380), .Z(n378) );
  XOR U2013 ( .A(n381), .B(n382), .Z(n380) );
  XOR U2014 ( .A(n383), .B(n384), .Z(n382) );
  XOR U2015 ( .A(n385), .B(n386), .Z(n384) );
  XOR U2016 ( .A(n387), .B(n388), .Z(n386) );
  XOR U2017 ( .A(n389), .B(n390), .Z(n388) );
  XOR U2018 ( .A(n391), .B(n392), .Z(n390) );
  XOR U2019 ( .A(n343), .B(n393), .Z(n392) );
  XOR U2020 ( .A(n394), .B(n344), .Z(n393) );
  XOR U2021 ( .A(n395), .B(n396), .Z(n344) );
  XOR U2022 ( .A(n342), .B(n397), .Z(n396) );
  XOR U2023 ( .A(n398), .B(n399), .Z(n397) );
  XOR U2024 ( .A(n400), .B(n401), .Z(n399) );
  XOR U2025 ( .A(n402), .B(n403), .Z(n401) );
  XOR U2026 ( .A(n404), .B(n405), .Z(n403) );
  XOR U2027 ( .A(n406), .B(n407), .Z(n405) );
  XOR U2028 ( .A(n408), .B(n409), .Z(n407) );
  XOR U2029 ( .A(n410), .B(n411), .Z(n409) );
  XOR U2030 ( .A(n412), .B(n413), .Z(n411) );
  XOR U2031 ( .A(n332), .B(n414), .Z(n413) );
  XOR U2032 ( .A(n415), .B(n333), .Z(n414) );
  XOR U2033 ( .A(n416), .B(n417), .Z(n333) );
  XOR U2034 ( .A(n331), .B(n418), .Z(n417) );
  XOR U2035 ( .A(n419), .B(n420), .Z(n418) );
  XOR U2036 ( .A(n421), .B(n422), .Z(n420) );
  XOR U2037 ( .A(n423), .B(n424), .Z(n422) );
  XOR U2038 ( .A(n425), .B(n426), .Z(n424) );
  XOR U2039 ( .A(n427), .B(n428), .Z(n426) );
  XOR U2040 ( .A(n429), .B(n430), .Z(n428) );
  XOR U2041 ( .A(n431), .B(n432), .Z(n430) );
  XOR U2042 ( .A(n433), .B(n434), .Z(n432) );
  XOR U2043 ( .A(n172), .B(n435), .Z(n434) );
  XOR U2044 ( .A(n436), .B(n173), .Z(n435) );
  XOR U2045 ( .A(n437), .B(n438), .Z(n173) );
  XOR U2046 ( .A(n171), .B(n439), .Z(n438) );
  XOR U2047 ( .A(n440), .B(n441), .Z(n439) );
  XOR U2048 ( .A(n442), .B(n443), .Z(n441) );
  XOR U2049 ( .A(n444), .B(n445), .Z(n443) );
  XOR U2050 ( .A(n446), .B(n447), .Z(n445) );
  XOR U2051 ( .A(n448), .B(n449), .Z(n447) );
  XOR U2052 ( .A(n450), .B(n451), .Z(n449) );
  XOR U2053 ( .A(n452), .B(n453), .Z(n451) );
  XNOR U2054 ( .A(n322), .B(n321), .Z(n453) );
  XOR U2055 ( .A(n454), .B(n320), .Z(n321) );
  AND U2056 ( .A(b[25]), .B(a[36]), .Z(n454) );
  XOR U2057 ( .A(n320), .B(n189), .Z(n455) );
  XOR U2058 ( .A(n456), .B(n457), .Z(n189) );
  XOR U2059 ( .A(n187), .B(n458), .Z(n457) );
  XOR U2060 ( .A(n459), .B(n460), .Z(n458) );
  XOR U2061 ( .A(n461), .B(n462), .Z(n460) );
  XOR U2062 ( .A(n463), .B(n464), .Z(n462) );
  XOR U2063 ( .A(n465), .B(n466), .Z(n464) );
  XOR U2064 ( .A(n467), .B(n468), .Z(n466) );
  XOR U2065 ( .A(n469), .B(n470), .Z(n468) );
  XOR U2066 ( .A(n471), .B(n472), .Z(n470) );
  XNOR U2067 ( .A(n312), .B(n311), .Z(n472) );
  XOR U2068 ( .A(n473), .B(n310), .Z(n311) );
  AND U2069 ( .A(b[31]), .B(a[30]), .Z(n473) );
  XOR U2070 ( .A(n310), .B(n205), .Z(n474) );
  XOR U2071 ( .A(n475), .B(n476), .Z(n205) );
  XOR U2072 ( .A(n203), .B(n477), .Z(n476) );
  XOR U2073 ( .A(n478), .B(n479), .Z(n477) );
  XOR U2074 ( .A(n480), .B(n481), .Z(n479) );
  XOR U2075 ( .A(n482), .B(n483), .Z(n481) );
  XOR U2076 ( .A(n484), .B(n485), .Z(n483) );
  XOR U2077 ( .A(n486), .B(n487), .Z(n485) );
  XOR U2078 ( .A(n488), .B(n489), .Z(n487) );
  XOR U2079 ( .A(n490), .B(n491), .Z(n489) );
  XNOR U2080 ( .A(n302), .B(n301), .Z(n491) );
  XOR U2081 ( .A(n492), .B(n300), .Z(n301) );
  AND U2082 ( .A(b[37]), .B(a[24]), .Z(n492) );
  XOR U2083 ( .A(n300), .B(n221), .Z(n493) );
  XOR U2084 ( .A(n494), .B(n495), .Z(n221) );
  XOR U2085 ( .A(n219), .B(n496), .Z(n495) );
  XOR U2086 ( .A(n497), .B(n498), .Z(n496) );
  XOR U2087 ( .A(n499), .B(n500), .Z(n498) );
  XOR U2088 ( .A(n501), .B(n502), .Z(n500) );
  XOR U2089 ( .A(n503), .B(n504), .Z(n502) );
  XOR U2090 ( .A(n505), .B(n506), .Z(n504) );
  XOR U2091 ( .A(n507), .B(n508), .Z(n506) );
  XOR U2092 ( .A(n509), .B(n510), .Z(n508) );
  XNOR U2093 ( .A(n292), .B(n291), .Z(n510) );
  XOR U2094 ( .A(n511), .B(n290), .Z(n291) );
  AND U2095 ( .A(b[43]), .B(a[18]), .Z(n511) );
  XOR U2096 ( .A(n290), .B(n237), .Z(n512) );
  XOR U2097 ( .A(n513), .B(n514), .Z(n237) );
  XOR U2098 ( .A(n235), .B(n515), .Z(n514) );
  XOR U2099 ( .A(n516), .B(n517), .Z(n515) );
  XOR U2100 ( .A(n518), .B(n519), .Z(n517) );
  XOR U2101 ( .A(n520), .B(n521), .Z(n519) );
  XOR U2102 ( .A(n522), .B(n523), .Z(n521) );
  XOR U2103 ( .A(n524), .B(n525), .Z(n523) );
  XOR U2104 ( .A(n526), .B(n527), .Z(n525) );
  XOR U2105 ( .A(n528), .B(n529), .Z(n527) );
  XNOR U2106 ( .A(n282), .B(n281), .Z(n529) );
  XOR U2107 ( .A(n530), .B(n280), .Z(n281) );
  AND U2108 ( .A(b[49]), .B(a[12]), .Z(n530) );
  XOR U2109 ( .A(n280), .B(n253), .Z(n531) );
  XOR U2110 ( .A(n532), .B(n533), .Z(n253) );
  XOR U2111 ( .A(n251), .B(n534), .Z(n533) );
  XOR U2112 ( .A(n535), .B(n536), .Z(n534) );
  XOR U2113 ( .A(n537), .B(n538), .Z(n536) );
  XOR U2114 ( .A(n539), .B(n540), .Z(n538) );
  XOR U2115 ( .A(n541), .B(n542), .Z(n540) );
  XOR U2116 ( .A(n543), .B(n544), .Z(n542) );
  XOR U2117 ( .A(n545), .B(n546), .Z(n544) );
  XOR U2118 ( .A(n547), .B(n548), .Z(n546) );
  XOR U2119 ( .A(n266), .B(n265), .Z(n548) );
  XOR U2120 ( .A(n549), .B(n264), .Z(n265) );
  AND U2121 ( .A(a[6]), .B(b[55]), .Z(n549) );
  XOR U2122 ( .A(n550), .B(n551), .Z(n266) );
  XOR U2123 ( .A(n264), .B(n552), .Z(n551) );
  XOR U2124 ( .A(n553), .B(n554), .Z(n552) );
  XOR U2125 ( .A(n555), .B(n556), .Z(n554) );
  XOR U2126 ( .A(n557), .B(n558), .Z(n556) );
  XOR U2127 ( .A(n559), .B(n560), .Z(n558) );
  XOR U2128 ( .A(n561), .B(n562), .Z(n560) );
  XOR U2129 ( .A(n563), .B(n564), .Z(n562) );
  XOR U2130 ( .A(n565), .B(n566), .Z(n564) );
  XOR U2131 ( .A(n567), .B(n568), .Z(n566) );
  XOR U2132 ( .A(n569), .B(n570), .Z(n568) );
  AND U2133 ( .A(a[0]), .B(b[61]), .Z(n569) );
  XNOR U2134 ( .A(n571), .B(n570), .Z(n565) );
  XNOR U2135 ( .A(n572), .B(n573), .Z(n570) );
  ANDN U2136 ( .B(n574), .A(n575), .Z(n572) );
  AND U2137 ( .A(a[1]), .B(b[60]), .Z(n571) );
  XOR U2138 ( .A(n576), .B(n567), .Z(n561) );
  XOR U2139 ( .A(n577), .B(n578), .Z(n567) );
  ANDN U2140 ( .B(n579), .A(n580), .Z(n577) );
  AND U2141 ( .A(a[2]), .B(b[59]), .Z(n576) );
  XOR U2142 ( .A(n581), .B(n563), .Z(n557) );
  XOR U2143 ( .A(n582), .B(n583), .Z(n563) );
  ANDN U2144 ( .B(n584), .A(n585), .Z(n582) );
  AND U2145 ( .A(a[3]), .B(b[58]), .Z(n581) );
  XOR U2146 ( .A(n586), .B(n559), .Z(n553) );
  XOR U2147 ( .A(n587), .B(n588), .Z(n559) );
  ANDN U2148 ( .B(n589), .A(n590), .Z(n587) );
  AND U2149 ( .A(a[4]), .B(b[57]), .Z(n586) );
  XOR U2150 ( .A(n591), .B(n592), .Z(n264) );
  AND U2151 ( .A(n593), .B(n594), .Z(n591) );
  XOR U2152 ( .A(n595), .B(n555), .Z(n550) );
  XOR U2153 ( .A(n596), .B(n597), .Z(n555) );
  ANDN U2154 ( .B(n598), .A(n599), .Z(n596) );
  AND U2155 ( .A(a[5]), .B(b[56]), .Z(n595) );
  XOR U2156 ( .A(n600), .B(n547), .Z(n543) );
  XNOR U2157 ( .A(n601), .B(n602), .Z(n547) );
  ANDN U2158 ( .B(n603), .A(n604), .Z(n601) );
  AND U2159 ( .A(a[7]), .B(b[54]), .Z(n600) );
  XOR U2160 ( .A(n605), .B(n545), .Z(n539) );
  XOR U2161 ( .A(n606), .B(n607), .Z(n545) );
  ANDN U2162 ( .B(n608), .A(n609), .Z(n606) );
  AND U2163 ( .A(a[8]), .B(b[53]), .Z(n605) );
  XOR U2164 ( .A(n610), .B(n541), .Z(n535) );
  XOR U2165 ( .A(n611), .B(n612), .Z(n541) );
  ANDN U2166 ( .B(n613), .A(n614), .Z(n611) );
  AND U2167 ( .A(a[9]), .B(b[52]), .Z(n610) );
  XOR U2168 ( .A(n615), .B(n537), .Z(n532) );
  XOR U2169 ( .A(n616), .B(n617), .Z(n537) );
  ANDN U2170 ( .B(n618), .A(n619), .Z(n616) );
  AND U2171 ( .A(a[10]), .B(b[51]), .Z(n615) );
  XOR U2172 ( .A(n620), .B(n621), .Z(n280) );
  AND U2173 ( .A(n622), .B(n623), .Z(n620) );
  XNOR U2174 ( .A(n624), .B(n251), .Z(n252) );
  XOR U2175 ( .A(n625), .B(n626), .Z(n251) );
  ANDN U2176 ( .B(n627), .A(n628), .Z(n625) );
  AND U2177 ( .A(b[50]), .B(a[11]), .Z(n624) );
  XOR U2178 ( .A(n629), .B(n528), .Z(n524) );
  XNOR U2179 ( .A(n630), .B(n631), .Z(n528) );
  ANDN U2180 ( .B(n632), .A(n633), .Z(n630) );
  AND U2181 ( .A(a[13]), .B(b[48]), .Z(n629) );
  XOR U2182 ( .A(n634), .B(n526), .Z(n520) );
  XOR U2183 ( .A(n635), .B(n636), .Z(n526) );
  ANDN U2184 ( .B(n637), .A(n638), .Z(n635) );
  AND U2185 ( .A(a[14]), .B(b[47]), .Z(n634) );
  XOR U2186 ( .A(n639), .B(n522), .Z(n516) );
  XOR U2187 ( .A(n640), .B(n641), .Z(n522) );
  ANDN U2188 ( .B(n642), .A(n643), .Z(n640) );
  AND U2189 ( .A(a[15]), .B(b[46]), .Z(n639) );
  XOR U2190 ( .A(n644), .B(n518), .Z(n513) );
  XOR U2191 ( .A(n645), .B(n646), .Z(n518) );
  ANDN U2192 ( .B(n647), .A(n648), .Z(n645) );
  AND U2193 ( .A(a[16]), .B(b[45]), .Z(n644) );
  XOR U2194 ( .A(n649), .B(n650), .Z(n290) );
  AND U2195 ( .A(n651), .B(n652), .Z(n649) );
  XNOR U2196 ( .A(n653), .B(n235), .Z(n236) );
  XOR U2197 ( .A(n654), .B(n655), .Z(n235) );
  ANDN U2198 ( .B(n656), .A(n657), .Z(n654) );
  AND U2199 ( .A(b[44]), .B(a[17]), .Z(n653) );
  XOR U2200 ( .A(n658), .B(n509), .Z(n505) );
  XNOR U2201 ( .A(n659), .B(n660), .Z(n509) );
  ANDN U2202 ( .B(n661), .A(n662), .Z(n659) );
  AND U2203 ( .A(a[19]), .B(b[42]), .Z(n658) );
  XOR U2204 ( .A(n663), .B(n507), .Z(n501) );
  XOR U2205 ( .A(n664), .B(n665), .Z(n507) );
  ANDN U2206 ( .B(n666), .A(n667), .Z(n664) );
  AND U2207 ( .A(a[20]), .B(b[41]), .Z(n663) );
  XOR U2208 ( .A(n668), .B(n503), .Z(n497) );
  XOR U2209 ( .A(n669), .B(n670), .Z(n503) );
  ANDN U2210 ( .B(n671), .A(n672), .Z(n669) );
  AND U2211 ( .A(a[21]), .B(b[40]), .Z(n668) );
  XOR U2212 ( .A(n673), .B(n499), .Z(n494) );
  XOR U2213 ( .A(n674), .B(n675), .Z(n499) );
  ANDN U2214 ( .B(n676), .A(n677), .Z(n674) );
  AND U2215 ( .A(a[22]), .B(b[39]), .Z(n673) );
  XOR U2216 ( .A(n678), .B(n679), .Z(n300) );
  AND U2217 ( .A(n680), .B(n681), .Z(n678) );
  XNOR U2218 ( .A(n682), .B(n219), .Z(n220) );
  XOR U2219 ( .A(n683), .B(n684), .Z(n219) );
  ANDN U2220 ( .B(n685), .A(n686), .Z(n683) );
  AND U2221 ( .A(b[38]), .B(a[23]), .Z(n682) );
  XOR U2222 ( .A(n687), .B(n490), .Z(n486) );
  XNOR U2223 ( .A(n688), .B(n689), .Z(n490) );
  ANDN U2224 ( .B(n690), .A(n691), .Z(n688) );
  AND U2225 ( .A(a[25]), .B(b[36]), .Z(n687) );
  XOR U2226 ( .A(n692), .B(n488), .Z(n482) );
  XOR U2227 ( .A(n693), .B(n694), .Z(n488) );
  ANDN U2228 ( .B(n695), .A(n696), .Z(n693) );
  AND U2229 ( .A(a[26]), .B(b[35]), .Z(n692) );
  XOR U2230 ( .A(n697), .B(n484), .Z(n478) );
  XOR U2231 ( .A(n698), .B(n699), .Z(n484) );
  ANDN U2232 ( .B(n700), .A(n701), .Z(n698) );
  AND U2233 ( .A(a[27]), .B(b[34]), .Z(n697) );
  XOR U2234 ( .A(n702), .B(n480), .Z(n475) );
  XOR U2235 ( .A(n703), .B(n704), .Z(n480) );
  ANDN U2236 ( .B(n705), .A(n706), .Z(n703) );
  AND U2237 ( .A(a[28]), .B(b[33]), .Z(n702) );
  XOR U2238 ( .A(n707), .B(n708), .Z(n310) );
  AND U2239 ( .A(n709), .B(n710), .Z(n707) );
  XNOR U2240 ( .A(n711), .B(n203), .Z(n204) );
  XOR U2241 ( .A(n712), .B(n713), .Z(n203) );
  ANDN U2242 ( .B(n714), .A(n715), .Z(n712) );
  AND U2243 ( .A(b[32]), .B(a[29]), .Z(n711) );
  XOR U2244 ( .A(n716), .B(n471), .Z(n467) );
  XNOR U2245 ( .A(n717), .B(n718), .Z(n471) );
  ANDN U2246 ( .B(n719), .A(n720), .Z(n717) );
  AND U2247 ( .A(a[31]), .B(b[30]), .Z(n716) );
  XOR U2248 ( .A(n721), .B(n469), .Z(n463) );
  XOR U2249 ( .A(n722), .B(n723), .Z(n469) );
  ANDN U2250 ( .B(n724), .A(n725), .Z(n722) );
  AND U2251 ( .A(a[32]), .B(b[29]), .Z(n721) );
  XOR U2252 ( .A(n726), .B(n465), .Z(n459) );
  XOR U2253 ( .A(n727), .B(n728), .Z(n465) );
  ANDN U2254 ( .B(n729), .A(n730), .Z(n727) );
  AND U2255 ( .A(a[33]), .B(b[28]), .Z(n726) );
  XOR U2256 ( .A(n731), .B(n461), .Z(n456) );
  XOR U2257 ( .A(n732), .B(n733), .Z(n461) );
  ANDN U2258 ( .B(n734), .A(n735), .Z(n732) );
  AND U2259 ( .A(a[34]), .B(b[27]), .Z(n731) );
  XOR U2260 ( .A(n736), .B(n737), .Z(n320) );
  AND U2261 ( .A(n738), .B(n739), .Z(n736) );
  XNOR U2262 ( .A(n740), .B(n187), .Z(n188) );
  XOR U2263 ( .A(n741), .B(n742), .Z(n187) );
  ANDN U2264 ( .B(n743), .A(n744), .Z(n741) );
  AND U2265 ( .A(b[26]), .B(a[35]), .Z(n740) );
  XOR U2266 ( .A(n745), .B(n452), .Z(n448) );
  XNOR U2267 ( .A(n746), .B(n747), .Z(n452) );
  ANDN U2268 ( .B(n748), .A(n749), .Z(n746) );
  AND U2269 ( .A(a[37]), .B(b[24]), .Z(n745) );
  XOR U2270 ( .A(n750), .B(n450), .Z(n444) );
  XOR U2271 ( .A(n751), .B(n752), .Z(n450) );
  ANDN U2272 ( .B(n753), .A(n754), .Z(n751) );
  AND U2273 ( .A(a[38]), .B(b[23]), .Z(n750) );
  XOR U2274 ( .A(n755), .B(n446), .Z(n440) );
  XOR U2275 ( .A(n756), .B(n757), .Z(n446) );
  ANDN U2276 ( .B(n758), .A(n759), .Z(n756) );
  AND U2277 ( .A(a[39]), .B(b[22]), .Z(n755) );
  XOR U2278 ( .A(n760), .B(n442), .Z(n437) );
  XOR U2279 ( .A(n761), .B(n762), .Z(n442) );
  ANDN U2280 ( .B(n763), .A(n764), .Z(n761) );
  AND U2281 ( .A(a[40]), .B(b[21]), .Z(n760) );
  XOR U2282 ( .A(n765), .B(n171), .Z(n172) );
  XOR U2283 ( .A(n766), .B(n767), .Z(n171) );
  ANDN U2284 ( .B(n768), .A(n769), .Z(n766) );
  AND U2285 ( .A(b[20]), .B(a[41]), .Z(n765) );
  XOR U2286 ( .A(n770), .B(n436), .Z(n431) );
  XOR U2287 ( .A(n771), .B(n772), .Z(n436) );
  ANDN U2288 ( .B(n773), .A(n774), .Z(n771) );
  AND U2289 ( .A(b[19]), .B(a[42]), .Z(n770) );
  XOR U2290 ( .A(n775), .B(n433), .Z(n427) );
  XOR U2291 ( .A(n776), .B(n777), .Z(n433) );
  ANDN U2292 ( .B(n778), .A(n779), .Z(n776) );
  AND U2293 ( .A(a[43]), .B(b[18]), .Z(n775) );
  XOR U2294 ( .A(n780), .B(n429), .Z(n423) );
  XOR U2295 ( .A(n781), .B(n782), .Z(n429) );
  ANDN U2296 ( .B(n783), .A(n784), .Z(n781) );
  AND U2297 ( .A(a[44]), .B(b[17]), .Z(n780) );
  XOR U2298 ( .A(n785), .B(n425), .Z(n419) );
  XOR U2299 ( .A(n786), .B(n787), .Z(n425) );
  ANDN U2300 ( .B(n788), .A(n789), .Z(n786) );
  AND U2301 ( .A(a[45]), .B(b[16]), .Z(n785) );
  XOR U2302 ( .A(n790), .B(n421), .Z(n416) );
  XOR U2303 ( .A(n791), .B(n792), .Z(n421) );
  ANDN U2304 ( .B(n793), .A(n794), .Z(n791) );
  AND U2305 ( .A(a[46]), .B(b[15]), .Z(n790) );
  XOR U2306 ( .A(n795), .B(n331), .Z(n332) );
  XOR U2307 ( .A(n796), .B(n797), .Z(n331) );
  ANDN U2308 ( .B(n798), .A(n799), .Z(n796) );
  AND U2309 ( .A(b[14]), .B(a[47]), .Z(n795) );
  XOR U2310 ( .A(n800), .B(n415), .Z(n410) );
  XOR U2311 ( .A(n801), .B(n802), .Z(n415) );
  ANDN U2312 ( .B(n803), .A(n804), .Z(n801) );
  AND U2313 ( .A(b[13]), .B(a[48]), .Z(n800) );
  XOR U2314 ( .A(n805), .B(n412), .Z(n406) );
  XOR U2315 ( .A(n806), .B(n807), .Z(n412) );
  ANDN U2316 ( .B(n808), .A(n809), .Z(n806) );
  AND U2317 ( .A(a[49]), .B(b[12]), .Z(n805) );
  XOR U2318 ( .A(n810), .B(n408), .Z(n402) );
  XOR U2319 ( .A(n811), .B(n812), .Z(n408) );
  ANDN U2320 ( .B(n813), .A(n814), .Z(n811) );
  AND U2321 ( .A(a[50]), .B(b[11]), .Z(n810) );
  XOR U2322 ( .A(n815), .B(n404), .Z(n398) );
  XOR U2323 ( .A(n816), .B(n817), .Z(n404) );
  ANDN U2324 ( .B(n818), .A(n819), .Z(n816) );
  AND U2325 ( .A(a[51]), .B(b[10]), .Z(n815) );
  XOR U2326 ( .A(n820), .B(n400), .Z(n395) );
  XOR U2327 ( .A(n821), .B(n822), .Z(n400) );
  ANDN U2328 ( .B(n823), .A(n824), .Z(n821) );
  AND U2329 ( .A(b[9]), .B(a[52]), .Z(n820) );
  XOR U2330 ( .A(n825), .B(n342), .Z(n343) );
  XOR U2331 ( .A(n826), .B(n827), .Z(n342) );
  ANDN U2332 ( .B(n828), .A(n829), .Z(n826) );
  AND U2333 ( .A(b[8]), .B(a[53]), .Z(n825) );
  XOR U2334 ( .A(n830), .B(n394), .Z(n389) );
  XOR U2335 ( .A(n831), .B(n832), .Z(n394) );
  ANDN U2336 ( .B(n833), .A(n834), .Z(n831) );
  AND U2337 ( .A(b[7]), .B(a[54]), .Z(n830) );
  XOR U2338 ( .A(n835), .B(n391), .Z(n385) );
  XOR U2339 ( .A(n836), .B(n837), .Z(n391) );
  ANDN U2340 ( .B(n838), .A(n839), .Z(n836) );
  AND U2341 ( .A(b[6]), .B(a[55]), .Z(n835) );
  XOR U2342 ( .A(n840), .B(n387), .Z(n381) );
  XOR U2343 ( .A(n841), .B(n842), .Z(n387) );
  ANDN U2344 ( .B(n843), .A(n844), .Z(n841) );
  AND U2345 ( .A(b[5]), .B(a[56]), .Z(n840) );
  XOR U2346 ( .A(n845), .B(n383), .Z(n377) );
  XOR U2347 ( .A(n846), .B(n847), .Z(n383) );
  ANDN U2348 ( .B(n848), .A(n849), .Z(n846) );
  AND U2349 ( .A(b[4]), .B(a[57]), .Z(n845) );
  XNOR U2350 ( .A(n850), .B(n851), .Z(n353) );
  NANDN U2351 ( .A(n852), .B(n853), .Z(n851) );
  XOR U2352 ( .A(n854), .B(n379), .Z(n374) );
  XNOR U2353 ( .A(n855), .B(n856), .Z(n379) );
  AND U2354 ( .A(n857), .B(n858), .Z(n855) );
  AND U2355 ( .A(b[3]), .B(a[58]), .Z(n854) );
  AND U2356 ( .A(a[61]), .B(b[0]), .Z(n364) );
  XNOR U2357 ( .A(n372), .B(n373), .Z(c[60]) );
  XNOR U2358 ( .A(n852), .B(n853), .Z(n373) );
  XOR U2359 ( .A(n850), .B(n859), .Z(n853) );
  NAND U2360 ( .A(b[1]), .B(a[59]), .Z(n859) );
  XOR U2361 ( .A(n858), .B(n860), .Z(n852) );
  XOR U2362 ( .A(n850), .B(n857), .Z(n860) );
  XNOR U2363 ( .A(n861), .B(n856), .Z(n857) );
  AND U2364 ( .A(b[2]), .B(a[58]), .Z(n861) );
  NANDN U2365 ( .A(n862), .B(n863), .Z(n850) );
  XOR U2366 ( .A(n856), .B(n848), .Z(n864) );
  XNOR U2367 ( .A(n847), .B(n843), .Z(n865) );
  XNOR U2368 ( .A(n842), .B(n838), .Z(n866) );
  XNOR U2369 ( .A(n837), .B(n833), .Z(n867) );
  XNOR U2370 ( .A(n832), .B(n828), .Z(n868) );
  XNOR U2371 ( .A(n827), .B(n823), .Z(n869) );
  XNOR U2372 ( .A(n822), .B(n818), .Z(n870) );
  XNOR U2373 ( .A(n817), .B(n813), .Z(n871) );
  XNOR U2374 ( .A(n812), .B(n808), .Z(n872) );
  XNOR U2375 ( .A(n807), .B(n803), .Z(n873) );
  XNOR U2376 ( .A(n802), .B(n798), .Z(n874) );
  XNOR U2377 ( .A(n797), .B(n793), .Z(n875) );
  XNOR U2378 ( .A(n792), .B(n788), .Z(n876) );
  XNOR U2379 ( .A(n787), .B(n783), .Z(n877) );
  XNOR U2380 ( .A(n782), .B(n778), .Z(n878) );
  XNOR U2381 ( .A(n777), .B(n773), .Z(n879) );
  XNOR U2382 ( .A(n772), .B(n768), .Z(n880) );
  XNOR U2383 ( .A(n767), .B(n763), .Z(n881) );
  XNOR U2384 ( .A(n762), .B(n758), .Z(n882) );
  XNOR U2385 ( .A(n757), .B(n753), .Z(n883) );
  XNOR U2386 ( .A(n752), .B(n748), .Z(n884) );
  XNOR U2387 ( .A(n739), .B(n738), .Z(n885) );
  XOR U2388 ( .A(n886), .B(n737), .Z(n738) );
  AND U2389 ( .A(b[24]), .B(a[36]), .Z(n886) );
  XNOR U2390 ( .A(n737), .B(n743), .Z(n887) );
  XNOR U2391 ( .A(n742), .B(n734), .Z(n888) );
  XNOR U2392 ( .A(n733), .B(n729), .Z(n889) );
  XNOR U2393 ( .A(n728), .B(n724), .Z(n890) );
  XNOR U2394 ( .A(n723), .B(n719), .Z(n891) );
  XNOR U2395 ( .A(n710), .B(n709), .Z(n892) );
  XOR U2396 ( .A(n893), .B(n708), .Z(n709) );
  AND U2397 ( .A(b[30]), .B(a[30]), .Z(n893) );
  XNOR U2398 ( .A(n708), .B(n714), .Z(n894) );
  XNOR U2399 ( .A(n713), .B(n705), .Z(n895) );
  XNOR U2400 ( .A(n704), .B(n700), .Z(n896) );
  XNOR U2401 ( .A(n699), .B(n695), .Z(n897) );
  XNOR U2402 ( .A(n694), .B(n690), .Z(n898) );
  XNOR U2403 ( .A(n681), .B(n680), .Z(n899) );
  XOR U2404 ( .A(n900), .B(n679), .Z(n680) );
  AND U2405 ( .A(b[36]), .B(a[24]), .Z(n900) );
  XNOR U2406 ( .A(n679), .B(n685), .Z(n901) );
  XNOR U2407 ( .A(n684), .B(n676), .Z(n902) );
  XNOR U2408 ( .A(n675), .B(n671), .Z(n903) );
  XNOR U2409 ( .A(n670), .B(n666), .Z(n904) );
  XNOR U2410 ( .A(n665), .B(n661), .Z(n905) );
  XNOR U2411 ( .A(n652), .B(n651), .Z(n906) );
  XOR U2412 ( .A(n907), .B(n650), .Z(n651) );
  AND U2413 ( .A(b[42]), .B(a[18]), .Z(n907) );
  XNOR U2414 ( .A(n650), .B(n656), .Z(n908) );
  XNOR U2415 ( .A(n655), .B(n647), .Z(n909) );
  XNOR U2416 ( .A(n646), .B(n642), .Z(n910) );
  XNOR U2417 ( .A(n641), .B(n637), .Z(n911) );
  XNOR U2418 ( .A(n636), .B(n632), .Z(n912) );
  XNOR U2419 ( .A(n623), .B(n622), .Z(n913) );
  XOR U2420 ( .A(n914), .B(n621), .Z(n622) );
  AND U2421 ( .A(b[48]), .B(a[12]), .Z(n914) );
  XNOR U2422 ( .A(n621), .B(n627), .Z(n915) );
  XNOR U2423 ( .A(n626), .B(n618), .Z(n916) );
  XNOR U2424 ( .A(n617), .B(n613), .Z(n917) );
  XNOR U2425 ( .A(n612), .B(n608), .Z(n918) );
  XNOR U2426 ( .A(n607), .B(n603), .Z(n919) );
  XNOR U2427 ( .A(n594), .B(n593), .Z(n920) );
  XOR U2428 ( .A(n921), .B(n592), .Z(n593) );
  AND U2429 ( .A(a[6]), .B(b[54]), .Z(n921) );
  XNOR U2430 ( .A(n592), .B(n598), .Z(n922) );
  XNOR U2431 ( .A(n597), .B(n589), .Z(n923) );
  XNOR U2432 ( .A(n588), .B(n584), .Z(n924) );
  XNOR U2433 ( .A(n583), .B(n579), .Z(n925) );
  XNOR U2434 ( .A(n578), .B(n574), .Z(n926) );
  XOR U2435 ( .A(n927), .B(n573), .Z(n574) );
  AND U2436 ( .A(a[0]), .B(b[60]), .Z(n927) );
  XNOR U2437 ( .A(n928), .B(n573), .Z(n575) );
  XNOR U2438 ( .A(n929), .B(n930), .Z(n573) );
  ANDN U2439 ( .B(n931), .A(n932), .Z(n929) );
  AND U2440 ( .A(a[1]), .B(b[59]), .Z(n928) );
  XNOR U2441 ( .A(n933), .B(n578), .Z(n580) );
  XOR U2442 ( .A(n934), .B(n935), .Z(n578) );
  ANDN U2443 ( .B(n936), .A(n937), .Z(n934) );
  AND U2444 ( .A(a[2]), .B(b[58]), .Z(n933) );
  XNOR U2445 ( .A(n938), .B(n583), .Z(n585) );
  XOR U2446 ( .A(n939), .B(n940), .Z(n583) );
  ANDN U2447 ( .B(n941), .A(n942), .Z(n939) );
  AND U2448 ( .A(a[3]), .B(b[57]), .Z(n938) );
  XNOR U2449 ( .A(n943), .B(n588), .Z(n590) );
  XOR U2450 ( .A(n944), .B(n945), .Z(n588) );
  ANDN U2451 ( .B(n946), .A(n947), .Z(n944) );
  AND U2452 ( .A(a[4]), .B(b[56]), .Z(n943) );
  XOR U2453 ( .A(n948), .B(n949), .Z(n592) );
  AND U2454 ( .A(n950), .B(n951), .Z(n948) );
  XNOR U2455 ( .A(n952), .B(n597), .Z(n599) );
  XOR U2456 ( .A(n953), .B(n954), .Z(n597) );
  ANDN U2457 ( .B(n955), .A(n956), .Z(n953) );
  AND U2458 ( .A(a[5]), .B(b[55]), .Z(n952) );
  XOR U2459 ( .A(n957), .B(n602), .Z(n604) );
  XOR U2460 ( .A(n958), .B(n959), .Z(n602) );
  ANDN U2461 ( .B(n960), .A(n961), .Z(n958) );
  AND U2462 ( .A(a[7]), .B(b[53]), .Z(n957) );
  XNOR U2463 ( .A(n962), .B(n607), .Z(n609) );
  XOR U2464 ( .A(n963), .B(n964), .Z(n607) );
  ANDN U2465 ( .B(n965), .A(n966), .Z(n963) );
  AND U2466 ( .A(a[8]), .B(b[52]), .Z(n962) );
  XNOR U2467 ( .A(n967), .B(n612), .Z(n614) );
  XOR U2468 ( .A(n968), .B(n969), .Z(n612) );
  ANDN U2469 ( .B(n970), .A(n971), .Z(n968) );
  AND U2470 ( .A(a[9]), .B(b[51]), .Z(n967) );
  XNOR U2471 ( .A(n972), .B(n617), .Z(n619) );
  XOR U2472 ( .A(n973), .B(n974), .Z(n617) );
  ANDN U2473 ( .B(n975), .A(n976), .Z(n973) );
  AND U2474 ( .A(b[50]), .B(a[10]), .Z(n972) );
  XOR U2475 ( .A(n977), .B(n978), .Z(n621) );
  AND U2476 ( .A(n979), .B(n980), .Z(n977) );
  XNOR U2477 ( .A(n981), .B(n626), .Z(n628) );
  XOR U2478 ( .A(n982), .B(n983), .Z(n626) );
  ANDN U2479 ( .B(n984), .A(n985), .Z(n982) );
  AND U2480 ( .A(b[49]), .B(a[11]), .Z(n981) );
  XOR U2481 ( .A(n986), .B(n631), .Z(n633) );
  XOR U2482 ( .A(n987), .B(n988), .Z(n631) );
  ANDN U2483 ( .B(n989), .A(n990), .Z(n987) );
  AND U2484 ( .A(a[13]), .B(b[47]), .Z(n986) );
  XNOR U2485 ( .A(n991), .B(n636), .Z(n638) );
  XOR U2486 ( .A(n992), .B(n993), .Z(n636) );
  ANDN U2487 ( .B(n994), .A(n995), .Z(n992) );
  AND U2488 ( .A(a[14]), .B(b[46]), .Z(n991) );
  XNOR U2489 ( .A(n996), .B(n641), .Z(n643) );
  XOR U2490 ( .A(n997), .B(n998), .Z(n641) );
  ANDN U2491 ( .B(n999), .A(n1000), .Z(n997) );
  AND U2492 ( .A(a[15]), .B(b[45]), .Z(n996) );
  XNOR U2493 ( .A(n1001), .B(n646), .Z(n648) );
  XOR U2494 ( .A(n1002), .B(n1003), .Z(n646) );
  ANDN U2495 ( .B(n1004), .A(n1005), .Z(n1002) );
  AND U2496 ( .A(b[44]), .B(a[16]), .Z(n1001) );
  XOR U2497 ( .A(n1006), .B(n1007), .Z(n650) );
  AND U2498 ( .A(n1008), .B(n1009), .Z(n1006) );
  XNOR U2499 ( .A(n1010), .B(n655), .Z(n657) );
  XOR U2500 ( .A(n1011), .B(n1012), .Z(n655) );
  ANDN U2501 ( .B(n1013), .A(n1014), .Z(n1011) );
  AND U2502 ( .A(b[43]), .B(a[17]), .Z(n1010) );
  XOR U2503 ( .A(n1015), .B(n660), .Z(n662) );
  XOR U2504 ( .A(n1016), .B(n1017), .Z(n660) );
  ANDN U2505 ( .B(n1018), .A(n1019), .Z(n1016) );
  AND U2506 ( .A(a[19]), .B(b[41]), .Z(n1015) );
  XNOR U2507 ( .A(n1020), .B(n665), .Z(n667) );
  XOR U2508 ( .A(n1021), .B(n1022), .Z(n665) );
  ANDN U2509 ( .B(n1023), .A(n1024), .Z(n1021) );
  AND U2510 ( .A(a[20]), .B(b[40]), .Z(n1020) );
  XNOR U2511 ( .A(n1025), .B(n670), .Z(n672) );
  XOR U2512 ( .A(n1026), .B(n1027), .Z(n670) );
  ANDN U2513 ( .B(n1028), .A(n1029), .Z(n1026) );
  AND U2514 ( .A(a[21]), .B(b[39]), .Z(n1025) );
  XNOR U2515 ( .A(n1030), .B(n675), .Z(n677) );
  XOR U2516 ( .A(n1031), .B(n1032), .Z(n675) );
  ANDN U2517 ( .B(n1033), .A(n1034), .Z(n1031) );
  AND U2518 ( .A(b[38]), .B(a[22]), .Z(n1030) );
  XOR U2519 ( .A(n1035), .B(n1036), .Z(n679) );
  AND U2520 ( .A(n1037), .B(n1038), .Z(n1035) );
  XNOR U2521 ( .A(n1039), .B(n684), .Z(n686) );
  XOR U2522 ( .A(n1040), .B(n1041), .Z(n684) );
  ANDN U2523 ( .B(n1042), .A(n1043), .Z(n1040) );
  AND U2524 ( .A(b[37]), .B(a[23]), .Z(n1039) );
  XOR U2525 ( .A(n1044), .B(n689), .Z(n691) );
  XOR U2526 ( .A(n1045), .B(n1046), .Z(n689) );
  ANDN U2527 ( .B(n1047), .A(n1048), .Z(n1045) );
  AND U2528 ( .A(a[25]), .B(b[35]), .Z(n1044) );
  XNOR U2529 ( .A(n1049), .B(n694), .Z(n696) );
  XOR U2530 ( .A(n1050), .B(n1051), .Z(n694) );
  ANDN U2531 ( .B(n1052), .A(n1053), .Z(n1050) );
  AND U2532 ( .A(a[26]), .B(b[34]), .Z(n1049) );
  XNOR U2533 ( .A(n1054), .B(n699), .Z(n701) );
  XOR U2534 ( .A(n1055), .B(n1056), .Z(n699) );
  ANDN U2535 ( .B(n1057), .A(n1058), .Z(n1055) );
  AND U2536 ( .A(a[27]), .B(b[33]), .Z(n1054) );
  XNOR U2537 ( .A(n1059), .B(n704), .Z(n706) );
  XOR U2538 ( .A(n1060), .B(n1061), .Z(n704) );
  ANDN U2539 ( .B(n1062), .A(n1063), .Z(n1060) );
  AND U2540 ( .A(b[32]), .B(a[28]), .Z(n1059) );
  XOR U2541 ( .A(n1064), .B(n1065), .Z(n708) );
  AND U2542 ( .A(n1066), .B(n1067), .Z(n1064) );
  XNOR U2543 ( .A(n1068), .B(n713), .Z(n715) );
  XOR U2544 ( .A(n1069), .B(n1070), .Z(n713) );
  ANDN U2545 ( .B(n1071), .A(n1072), .Z(n1069) );
  AND U2546 ( .A(b[31]), .B(a[29]), .Z(n1068) );
  XOR U2547 ( .A(n1073), .B(n718), .Z(n720) );
  XOR U2548 ( .A(n1074), .B(n1075), .Z(n718) );
  ANDN U2549 ( .B(n1076), .A(n1077), .Z(n1074) );
  AND U2550 ( .A(a[31]), .B(b[29]), .Z(n1073) );
  XNOR U2551 ( .A(n1078), .B(n723), .Z(n725) );
  XOR U2552 ( .A(n1079), .B(n1080), .Z(n723) );
  ANDN U2553 ( .B(n1081), .A(n1082), .Z(n1079) );
  AND U2554 ( .A(a[32]), .B(b[28]), .Z(n1078) );
  XNOR U2555 ( .A(n1083), .B(n728), .Z(n730) );
  XOR U2556 ( .A(n1084), .B(n1085), .Z(n728) );
  ANDN U2557 ( .B(n1086), .A(n1087), .Z(n1084) );
  AND U2558 ( .A(a[33]), .B(b[27]), .Z(n1083) );
  XNOR U2559 ( .A(n1088), .B(n733), .Z(n735) );
  XOR U2560 ( .A(n1089), .B(n1090), .Z(n733) );
  ANDN U2561 ( .B(n1091), .A(n1092), .Z(n1089) );
  AND U2562 ( .A(b[26]), .B(a[34]), .Z(n1088) );
  XOR U2563 ( .A(n1093), .B(n1094), .Z(n737) );
  AND U2564 ( .A(n1095), .B(n1096), .Z(n1093) );
  XNOR U2565 ( .A(n1097), .B(n742), .Z(n744) );
  XOR U2566 ( .A(n1098), .B(n1099), .Z(n742) );
  ANDN U2567 ( .B(n1100), .A(n1101), .Z(n1098) );
  AND U2568 ( .A(b[25]), .B(a[35]), .Z(n1097) );
  XOR U2569 ( .A(n1102), .B(n747), .Z(n749) );
  XOR U2570 ( .A(n1103), .B(n1104), .Z(n747) );
  ANDN U2571 ( .B(n1105), .A(n1106), .Z(n1103) );
  AND U2572 ( .A(a[37]), .B(b[23]), .Z(n1102) );
  XNOR U2573 ( .A(n1107), .B(n752), .Z(n754) );
  XOR U2574 ( .A(n1108), .B(n1109), .Z(n752) );
  ANDN U2575 ( .B(n1110), .A(n1111), .Z(n1108) );
  AND U2576 ( .A(a[38]), .B(b[22]), .Z(n1107) );
  XNOR U2577 ( .A(n1112), .B(n757), .Z(n759) );
  XOR U2578 ( .A(n1113), .B(n1114), .Z(n757) );
  ANDN U2579 ( .B(n1115), .A(n1116), .Z(n1113) );
  AND U2580 ( .A(a[39]), .B(b[21]), .Z(n1112) );
  XNOR U2581 ( .A(n1117), .B(n762), .Z(n764) );
  XOR U2582 ( .A(n1118), .B(n1119), .Z(n762) );
  ANDN U2583 ( .B(n1120), .A(n1121), .Z(n1118) );
  AND U2584 ( .A(b[20]), .B(a[40]), .Z(n1117) );
  XNOR U2585 ( .A(n1122), .B(n767), .Z(n769) );
  XOR U2586 ( .A(n1123), .B(n1124), .Z(n767) );
  ANDN U2587 ( .B(n1125), .A(n1126), .Z(n1123) );
  AND U2588 ( .A(b[19]), .B(a[41]), .Z(n1122) );
  XNOR U2589 ( .A(n1127), .B(n772), .Z(n774) );
  XOR U2590 ( .A(n1128), .B(n1129), .Z(n772) );
  ANDN U2591 ( .B(n1130), .A(n1131), .Z(n1128) );
  AND U2592 ( .A(b[18]), .B(a[42]), .Z(n1127) );
  XNOR U2593 ( .A(n1132), .B(n777), .Z(n779) );
  XOR U2594 ( .A(n1133), .B(n1134), .Z(n777) );
  ANDN U2595 ( .B(n1135), .A(n1136), .Z(n1133) );
  AND U2596 ( .A(a[43]), .B(b[17]), .Z(n1132) );
  XNOR U2597 ( .A(n1137), .B(n782), .Z(n784) );
  XOR U2598 ( .A(n1138), .B(n1139), .Z(n782) );
  ANDN U2599 ( .B(n1140), .A(n1141), .Z(n1138) );
  AND U2600 ( .A(a[44]), .B(b[16]), .Z(n1137) );
  XNOR U2601 ( .A(n1142), .B(n787), .Z(n789) );
  XOR U2602 ( .A(n1143), .B(n1144), .Z(n787) );
  ANDN U2603 ( .B(n1145), .A(n1146), .Z(n1143) );
  AND U2604 ( .A(a[45]), .B(b[15]), .Z(n1142) );
  XNOR U2605 ( .A(n1147), .B(n792), .Z(n794) );
  XOR U2606 ( .A(n1148), .B(n1149), .Z(n792) );
  ANDN U2607 ( .B(n1150), .A(n1151), .Z(n1148) );
  AND U2608 ( .A(b[14]), .B(a[46]), .Z(n1147) );
  XNOR U2609 ( .A(n1152), .B(n797), .Z(n799) );
  XOR U2610 ( .A(n1153), .B(n1154), .Z(n797) );
  ANDN U2611 ( .B(n1155), .A(n1156), .Z(n1153) );
  AND U2612 ( .A(b[13]), .B(a[47]), .Z(n1152) );
  XNOR U2613 ( .A(n1157), .B(n802), .Z(n804) );
  XOR U2614 ( .A(n1158), .B(n1159), .Z(n802) );
  ANDN U2615 ( .B(n1160), .A(n1161), .Z(n1158) );
  AND U2616 ( .A(b[12]), .B(a[48]), .Z(n1157) );
  XNOR U2617 ( .A(n1162), .B(n807), .Z(n809) );
  XOR U2618 ( .A(n1163), .B(n1164), .Z(n807) );
  ANDN U2619 ( .B(n1165), .A(n1166), .Z(n1163) );
  AND U2620 ( .A(a[49]), .B(b[11]), .Z(n1162) );
  XNOR U2621 ( .A(n1167), .B(n812), .Z(n814) );
  XOR U2622 ( .A(n1168), .B(n1169), .Z(n812) );
  ANDN U2623 ( .B(n1170), .A(n1171), .Z(n1168) );
  AND U2624 ( .A(a[50]), .B(b[10]), .Z(n1167) );
  XNOR U2625 ( .A(n1172), .B(n817), .Z(n819) );
  XOR U2626 ( .A(n1173), .B(n1174), .Z(n817) );
  ANDN U2627 ( .B(n1175), .A(n1176), .Z(n1173) );
  AND U2628 ( .A(b[9]), .B(a[51]), .Z(n1172) );
  XNOR U2629 ( .A(n1177), .B(n822), .Z(n824) );
  XOR U2630 ( .A(n1178), .B(n1179), .Z(n822) );
  ANDN U2631 ( .B(n1180), .A(n1181), .Z(n1178) );
  AND U2632 ( .A(b[8]), .B(a[52]), .Z(n1177) );
  XNOR U2633 ( .A(n1182), .B(n827), .Z(n829) );
  XOR U2634 ( .A(n1183), .B(n1184), .Z(n827) );
  ANDN U2635 ( .B(n1185), .A(n1186), .Z(n1183) );
  AND U2636 ( .A(b[7]), .B(a[53]), .Z(n1182) );
  XNOR U2637 ( .A(n1187), .B(n832), .Z(n834) );
  XOR U2638 ( .A(n1188), .B(n1189), .Z(n832) );
  ANDN U2639 ( .B(n1190), .A(n1191), .Z(n1188) );
  AND U2640 ( .A(b[6]), .B(a[54]), .Z(n1187) );
  XNOR U2641 ( .A(n1192), .B(n837), .Z(n839) );
  XOR U2642 ( .A(n1193), .B(n1194), .Z(n837) );
  ANDN U2643 ( .B(n1195), .A(n1196), .Z(n1193) );
  AND U2644 ( .A(b[5]), .B(a[55]), .Z(n1192) );
  XNOR U2645 ( .A(n1197), .B(n842), .Z(n844) );
  XOR U2646 ( .A(n1198), .B(n1199), .Z(n842) );
  ANDN U2647 ( .B(n1200), .A(n1201), .Z(n1198) );
  AND U2648 ( .A(b[4]), .B(a[56]), .Z(n1197) );
  XNOR U2649 ( .A(n1202), .B(n1203), .Z(n856) );
  NANDN U2650 ( .A(n1204), .B(n1205), .Z(n1203) );
  XNOR U2651 ( .A(n1206), .B(n847), .Z(n849) );
  XNOR U2652 ( .A(n1207), .B(n1208), .Z(n847) );
  AND U2653 ( .A(n1209), .B(n1210), .Z(n1207) );
  AND U2654 ( .A(b[3]), .B(a[57]), .Z(n1206) );
  NAND U2655 ( .A(a[60]), .B(b[0]), .Z(n372) );
  XNOR U2656 ( .A(n1211), .B(n1212), .Z(c[5]) );
  XNOR U2657 ( .A(n862), .B(n863), .Z(c[59]) );
  XNOR U2658 ( .A(n1204), .B(n1205), .Z(n863) );
  XOR U2659 ( .A(n1202), .B(n1213), .Z(n1205) );
  NAND U2660 ( .A(b[1]), .B(a[58]), .Z(n1213) );
  XOR U2661 ( .A(n1210), .B(n1214), .Z(n1204) );
  XOR U2662 ( .A(n1202), .B(n1209), .Z(n1214) );
  XNOR U2663 ( .A(n1215), .B(n1208), .Z(n1209) );
  AND U2664 ( .A(b[2]), .B(a[57]), .Z(n1215) );
  NANDN U2665 ( .A(n1216), .B(n1217), .Z(n1202) );
  XOR U2666 ( .A(n1208), .B(n1200), .Z(n1218) );
  XNOR U2667 ( .A(n1199), .B(n1195), .Z(n1219) );
  XNOR U2668 ( .A(n1194), .B(n1190), .Z(n1220) );
  XNOR U2669 ( .A(n1189), .B(n1185), .Z(n1221) );
  XNOR U2670 ( .A(n1184), .B(n1180), .Z(n1222) );
  XNOR U2671 ( .A(n1179), .B(n1175), .Z(n1223) );
  XNOR U2672 ( .A(n1174), .B(n1170), .Z(n1224) );
  XNOR U2673 ( .A(n1169), .B(n1165), .Z(n1225) );
  XNOR U2674 ( .A(n1164), .B(n1160), .Z(n1226) );
  XNOR U2675 ( .A(n1159), .B(n1155), .Z(n1227) );
  XNOR U2676 ( .A(n1154), .B(n1150), .Z(n1228) );
  XNOR U2677 ( .A(n1149), .B(n1145), .Z(n1229) );
  XNOR U2678 ( .A(n1144), .B(n1140), .Z(n1230) );
  XNOR U2679 ( .A(n1139), .B(n1135), .Z(n1231) );
  XNOR U2680 ( .A(n1134), .B(n1130), .Z(n1232) );
  XNOR U2681 ( .A(n1129), .B(n1125), .Z(n1233) );
  XNOR U2682 ( .A(n1124), .B(n1120), .Z(n1234) );
  XNOR U2683 ( .A(n1119), .B(n1115), .Z(n1235) );
  XNOR U2684 ( .A(n1114), .B(n1110), .Z(n1236) );
  XNOR U2685 ( .A(n1109), .B(n1105), .Z(n1237) );
  XNOR U2686 ( .A(n1096), .B(n1095), .Z(n1238) );
  XOR U2687 ( .A(n1239), .B(n1094), .Z(n1095) );
  AND U2688 ( .A(b[23]), .B(a[36]), .Z(n1239) );
  XNOR U2689 ( .A(n1094), .B(n1100), .Z(n1240) );
  XNOR U2690 ( .A(n1099), .B(n1091), .Z(n1241) );
  XNOR U2691 ( .A(n1090), .B(n1086), .Z(n1242) );
  XNOR U2692 ( .A(n1085), .B(n1081), .Z(n1243) );
  XNOR U2693 ( .A(n1080), .B(n1076), .Z(n1244) );
  XNOR U2694 ( .A(n1067), .B(n1066), .Z(n1245) );
  XOR U2695 ( .A(n1246), .B(n1065), .Z(n1066) );
  AND U2696 ( .A(b[29]), .B(a[30]), .Z(n1246) );
  XNOR U2697 ( .A(n1065), .B(n1071), .Z(n1247) );
  XNOR U2698 ( .A(n1070), .B(n1062), .Z(n1248) );
  XNOR U2699 ( .A(n1061), .B(n1057), .Z(n1249) );
  XNOR U2700 ( .A(n1056), .B(n1052), .Z(n1250) );
  XNOR U2701 ( .A(n1051), .B(n1047), .Z(n1251) );
  XNOR U2702 ( .A(n1038), .B(n1037), .Z(n1252) );
  XOR U2703 ( .A(n1253), .B(n1036), .Z(n1037) );
  AND U2704 ( .A(b[35]), .B(a[24]), .Z(n1253) );
  XNOR U2705 ( .A(n1036), .B(n1042), .Z(n1254) );
  XNOR U2706 ( .A(n1041), .B(n1033), .Z(n1255) );
  XNOR U2707 ( .A(n1032), .B(n1028), .Z(n1256) );
  XNOR U2708 ( .A(n1027), .B(n1023), .Z(n1257) );
  XNOR U2709 ( .A(n1022), .B(n1018), .Z(n1258) );
  XNOR U2710 ( .A(n1009), .B(n1008), .Z(n1259) );
  XOR U2711 ( .A(n1260), .B(n1007), .Z(n1008) );
  AND U2712 ( .A(b[41]), .B(a[18]), .Z(n1260) );
  XNOR U2713 ( .A(n1007), .B(n1013), .Z(n1261) );
  XNOR U2714 ( .A(n1012), .B(n1004), .Z(n1262) );
  XNOR U2715 ( .A(n1003), .B(n999), .Z(n1263) );
  XNOR U2716 ( .A(n998), .B(n994), .Z(n1264) );
  XNOR U2717 ( .A(n993), .B(n989), .Z(n1265) );
  XNOR U2718 ( .A(n980), .B(n979), .Z(n1266) );
  XOR U2719 ( .A(n1267), .B(n978), .Z(n979) );
  AND U2720 ( .A(b[47]), .B(a[12]), .Z(n1267) );
  XNOR U2721 ( .A(n978), .B(n984), .Z(n1268) );
  XNOR U2722 ( .A(n983), .B(n975), .Z(n1269) );
  XNOR U2723 ( .A(n974), .B(n970), .Z(n1270) );
  XNOR U2724 ( .A(n969), .B(n965), .Z(n1271) );
  XNOR U2725 ( .A(n964), .B(n960), .Z(n1272) );
  XNOR U2726 ( .A(n951), .B(n950), .Z(n1273) );
  XOR U2727 ( .A(n1274), .B(n949), .Z(n950) );
  AND U2728 ( .A(a[6]), .B(b[53]), .Z(n1274) );
  XNOR U2729 ( .A(n949), .B(n955), .Z(n1275) );
  XNOR U2730 ( .A(n954), .B(n946), .Z(n1276) );
  XNOR U2731 ( .A(n945), .B(n941), .Z(n1277) );
  XNOR U2732 ( .A(n940), .B(n936), .Z(n1278) );
  XNOR U2733 ( .A(n935), .B(n931), .Z(n1279) );
  XNOR U2734 ( .A(n1280), .B(n930), .Z(n931) );
  AND U2735 ( .A(a[0]), .B(b[59]), .Z(n1280) );
  XOR U2736 ( .A(n1281), .B(n930), .Z(n932) );
  XNOR U2737 ( .A(n1282), .B(n1283), .Z(n930) );
  ANDN U2738 ( .B(n1284), .A(n1285), .Z(n1282) );
  AND U2739 ( .A(a[1]), .B(b[58]), .Z(n1281) );
  XNOR U2740 ( .A(n1286), .B(n935), .Z(n937) );
  XOR U2741 ( .A(n1287), .B(n1288), .Z(n935) );
  ANDN U2742 ( .B(n1289), .A(n1290), .Z(n1287) );
  AND U2743 ( .A(a[2]), .B(b[57]), .Z(n1286) );
  XNOR U2744 ( .A(n1291), .B(n940), .Z(n942) );
  XOR U2745 ( .A(n1292), .B(n1293), .Z(n940) );
  ANDN U2746 ( .B(n1294), .A(n1295), .Z(n1292) );
  AND U2747 ( .A(a[3]), .B(b[56]), .Z(n1291) );
  XNOR U2748 ( .A(n1296), .B(n945), .Z(n947) );
  XOR U2749 ( .A(n1297), .B(n1298), .Z(n945) );
  ANDN U2750 ( .B(n1299), .A(n1300), .Z(n1297) );
  AND U2751 ( .A(a[4]), .B(b[55]), .Z(n1296) );
  XOR U2752 ( .A(n1301), .B(n1302), .Z(n949) );
  AND U2753 ( .A(n1303), .B(n1304), .Z(n1301) );
  XNOR U2754 ( .A(n1305), .B(n954), .Z(n956) );
  XOR U2755 ( .A(n1306), .B(n1307), .Z(n954) );
  ANDN U2756 ( .B(n1308), .A(n1309), .Z(n1306) );
  AND U2757 ( .A(a[5]), .B(b[54]), .Z(n1305) );
  XOR U2758 ( .A(n1310), .B(n959), .Z(n961) );
  XOR U2759 ( .A(n1311), .B(n1312), .Z(n959) );
  ANDN U2760 ( .B(n1313), .A(n1314), .Z(n1311) );
  AND U2761 ( .A(a[7]), .B(b[52]), .Z(n1310) );
  XNOR U2762 ( .A(n1315), .B(n964), .Z(n966) );
  XOR U2763 ( .A(n1316), .B(n1317), .Z(n964) );
  ANDN U2764 ( .B(n1318), .A(n1319), .Z(n1316) );
  AND U2765 ( .A(a[8]), .B(b[51]), .Z(n1315) );
  XNOR U2766 ( .A(n1320), .B(n969), .Z(n971) );
  XOR U2767 ( .A(n1321), .B(n1322), .Z(n969) );
  ANDN U2768 ( .B(n1323), .A(n1324), .Z(n1321) );
  AND U2769 ( .A(a[9]), .B(b[50]), .Z(n1320) );
  XNOR U2770 ( .A(n1325), .B(n974), .Z(n976) );
  XOR U2771 ( .A(n1326), .B(n1327), .Z(n974) );
  ANDN U2772 ( .B(n1328), .A(n1329), .Z(n1326) );
  AND U2773 ( .A(b[49]), .B(a[10]), .Z(n1325) );
  XOR U2774 ( .A(n1330), .B(n1331), .Z(n978) );
  AND U2775 ( .A(n1332), .B(n1333), .Z(n1330) );
  XNOR U2776 ( .A(n1334), .B(n983), .Z(n985) );
  XOR U2777 ( .A(n1335), .B(n1336), .Z(n983) );
  ANDN U2778 ( .B(n1337), .A(n1338), .Z(n1335) );
  AND U2779 ( .A(b[48]), .B(a[11]), .Z(n1334) );
  XOR U2780 ( .A(n1339), .B(n988), .Z(n990) );
  XOR U2781 ( .A(n1340), .B(n1341), .Z(n988) );
  ANDN U2782 ( .B(n1342), .A(n1343), .Z(n1340) );
  AND U2783 ( .A(a[13]), .B(b[46]), .Z(n1339) );
  XNOR U2784 ( .A(n1344), .B(n993), .Z(n995) );
  XOR U2785 ( .A(n1345), .B(n1346), .Z(n993) );
  ANDN U2786 ( .B(n1347), .A(n1348), .Z(n1345) );
  AND U2787 ( .A(a[14]), .B(b[45]), .Z(n1344) );
  XNOR U2788 ( .A(n1349), .B(n998), .Z(n1000) );
  XOR U2789 ( .A(n1350), .B(n1351), .Z(n998) );
  ANDN U2790 ( .B(n1352), .A(n1353), .Z(n1350) );
  AND U2791 ( .A(b[44]), .B(a[15]), .Z(n1349) );
  XNOR U2792 ( .A(n1354), .B(n1003), .Z(n1005) );
  XOR U2793 ( .A(n1355), .B(n1356), .Z(n1003) );
  ANDN U2794 ( .B(n1357), .A(n1358), .Z(n1355) );
  AND U2795 ( .A(b[43]), .B(a[16]), .Z(n1354) );
  XOR U2796 ( .A(n1359), .B(n1360), .Z(n1007) );
  AND U2797 ( .A(n1361), .B(n1362), .Z(n1359) );
  XNOR U2798 ( .A(n1363), .B(n1012), .Z(n1014) );
  XOR U2799 ( .A(n1364), .B(n1365), .Z(n1012) );
  ANDN U2800 ( .B(n1366), .A(n1367), .Z(n1364) );
  AND U2801 ( .A(b[42]), .B(a[17]), .Z(n1363) );
  XOR U2802 ( .A(n1368), .B(n1017), .Z(n1019) );
  XOR U2803 ( .A(n1369), .B(n1370), .Z(n1017) );
  ANDN U2804 ( .B(n1371), .A(n1372), .Z(n1369) );
  AND U2805 ( .A(a[19]), .B(b[40]), .Z(n1368) );
  XNOR U2806 ( .A(n1373), .B(n1022), .Z(n1024) );
  XOR U2807 ( .A(n1374), .B(n1375), .Z(n1022) );
  ANDN U2808 ( .B(n1376), .A(n1377), .Z(n1374) );
  AND U2809 ( .A(a[20]), .B(b[39]), .Z(n1373) );
  XNOR U2810 ( .A(n1378), .B(n1027), .Z(n1029) );
  XOR U2811 ( .A(n1379), .B(n1380), .Z(n1027) );
  ANDN U2812 ( .B(n1381), .A(n1382), .Z(n1379) );
  AND U2813 ( .A(b[38]), .B(a[21]), .Z(n1378) );
  XNOR U2814 ( .A(n1383), .B(n1032), .Z(n1034) );
  XOR U2815 ( .A(n1384), .B(n1385), .Z(n1032) );
  ANDN U2816 ( .B(n1386), .A(n1387), .Z(n1384) );
  AND U2817 ( .A(b[37]), .B(a[22]), .Z(n1383) );
  XOR U2818 ( .A(n1388), .B(n1389), .Z(n1036) );
  AND U2819 ( .A(n1390), .B(n1391), .Z(n1388) );
  XNOR U2820 ( .A(n1392), .B(n1041), .Z(n1043) );
  XOR U2821 ( .A(n1393), .B(n1394), .Z(n1041) );
  ANDN U2822 ( .B(n1395), .A(n1396), .Z(n1393) );
  AND U2823 ( .A(b[36]), .B(a[23]), .Z(n1392) );
  XOR U2824 ( .A(n1397), .B(n1046), .Z(n1048) );
  XOR U2825 ( .A(n1398), .B(n1399), .Z(n1046) );
  ANDN U2826 ( .B(n1400), .A(n1401), .Z(n1398) );
  AND U2827 ( .A(a[25]), .B(b[34]), .Z(n1397) );
  XNOR U2828 ( .A(n1402), .B(n1051), .Z(n1053) );
  XOR U2829 ( .A(n1403), .B(n1404), .Z(n1051) );
  ANDN U2830 ( .B(n1405), .A(n1406), .Z(n1403) );
  AND U2831 ( .A(a[26]), .B(b[33]), .Z(n1402) );
  XNOR U2832 ( .A(n1407), .B(n1056), .Z(n1058) );
  XOR U2833 ( .A(n1408), .B(n1409), .Z(n1056) );
  ANDN U2834 ( .B(n1410), .A(n1411), .Z(n1408) );
  AND U2835 ( .A(b[32]), .B(a[27]), .Z(n1407) );
  XNOR U2836 ( .A(n1412), .B(n1061), .Z(n1063) );
  XOR U2837 ( .A(n1413), .B(n1414), .Z(n1061) );
  ANDN U2838 ( .B(n1415), .A(n1416), .Z(n1413) );
  AND U2839 ( .A(b[31]), .B(a[28]), .Z(n1412) );
  XOR U2840 ( .A(n1417), .B(n1418), .Z(n1065) );
  AND U2841 ( .A(n1419), .B(n1420), .Z(n1417) );
  XNOR U2842 ( .A(n1421), .B(n1070), .Z(n1072) );
  XOR U2843 ( .A(n1422), .B(n1423), .Z(n1070) );
  ANDN U2844 ( .B(n1424), .A(n1425), .Z(n1422) );
  AND U2845 ( .A(b[30]), .B(a[29]), .Z(n1421) );
  XOR U2846 ( .A(n1426), .B(n1075), .Z(n1077) );
  XOR U2847 ( .A(n1427), .B(n1428), .Z(n1075) );
  ANDN U2848 ( .B(n1429), .A(n1430), .Z(n1427) );
  AND U2849 ( .A(a[31]), .B(b[28]), .Z(n1426) );
  XNOR U2850 ( .A(n1431), .B(n1080), .Z(n1082) );
  XOR U2851 ( .A(n1432), .B(n1433), .Z(n1080) );
  ANDN U2852 ( .B(n1434), .A(n1435), .Z(n1432) );
  AND U2853 ( .A(a[32]), .B(b[27]), .Z(n1431) );
  XNOR U2854 ( .A(n1436), .B(n1085), .Z(n1087) );
  XOR U2855 ( .A(n1437), .B(n1438), .Z(n1085) );
  ANDN U2856 ( .B(n1439), .A(n1440), .Z(n1437) );
  AND U2857 ( .A(b[26]), .B(a[33]), .Z(n1436) );
  XNOR U2858 ( .A(n1441), .B(n1090), .Z(n1092) );
  XOR U2859 ( .A(n1442), .B(n1443), .Z(n1090) );
  ANDN U2860 ( .B(n1444), .A(n1445), .Z(n1442) );
  AND U2861 ( .A(b[25]), .B(a[34]), .Z(n1441) );
  XOR U2862 ( .A(n1446), .B(n1447), .Z(n1094) );
  AND U2863 ( .A(n1448), .B(n1449), .Z(n1446) );
  XNOR U2864 ( .A(n1450), .B(n1099), .Z(n1101) );
  XOR U2865 ( .A(n1451), .B(n1452), .Z(n1099) );
  ANDN U2866 ( .B(n1453), .A(n1454), .Z(n1451) );
  AND U2867 ( .A(b[24]), .B(a[35]), .Z(n1450) );
  XOR U2868 ( .A(n1455), .B(n1104), .Z(n1106) );
  XOR U2869 ( .A(n1456), .B(n1457), .Z(n1104) );
  ANDN U2870 ( .B(n1458), .A(n1459), .Z(n1456) );
  AND U2871 ( .A(a[37]), .B(b[22]), .Z(n1455) );
  XNOR U2872 ( .A(n1460), .B(n1109), .Z(n1111) );
  XOR U2873 ( .A(n1461), .B(n1462), .Z(n1109) );
  ANDN U2874 ( .B(n1463), .A(n1464), .Z(n1461) );
  AND U2875 ( .A(a[38]), .B(b[21]), .Z(n1460) );
  XNOR U2876 ( .A(n1465), .B(n1114), .Z(n1116) );
  XOR U2877 ( .A(n1466), .B(n1467), .Z(n1114) );
  ANDN U2878 ( .B(n1468), .A(n1469), .Z(n1466) );
  AND U2879 ( .A(b[20]), .B(a[39]), .Z(n1465) );
  XNOR U2880 ( .A(n1470), .B(n1119), .Z(n1121) );
  XOR U2881 ( .A(n1471), .B(n1472), .Z(n1119) );
  ANDN U2882 ( .B(n1473), .A(n1474), .Z(n1471) );
  AND U2883 ( .A(b[19]), .B(a[40]), .Z(n1470) );
  XNOR U2884 ( .A(n1475), .B(n1124), .Z(n1126) );
  XOR U2885 ( .A(n1476), .B(n1477), .Z(n1124) );
  ANDN U2886 ( .B(n1478), .A(n1479), .Z(n1476) );
  AND U2887 ( .A(b[18]), .B(a[41]), .Z(n1475) );
  XNOR U2888 ( .A(n1480), .B(n1129), .Z(n1131) );
  XOR U2889 ( .A(n1481), .B(n1482), .Z(n1129) );
  ANDN U2890 ( .B(n1483), .A(n1484), .Z(n1481) );
  AND U2891 ( .A(b[17]), .B(a[42]), .Z(n1480) );
  XNOR U2892 ( .A(n1485), .B(n1134), .Z(n1136) );
  XOR U2893 ( .A(n1486), .B(n1487), .Z(n1134) );
  ANDN U2894 ( .B(n1488), .A(n1489), .Z(n1486) );
  AND U2895 ( .A(a[43]), .B(b[16]), .Z(n1485) );
  XNOR U2896 ( .A(n1490), .B(n1139), .Z(n1141) );
  XOR U2897 ( .A(n1491), .B(n1492), .Z(n1139) );
  ANDN U2898 ( .B(n1493), .A(n1494), .Z(n1491) );
  AND U2899 ( .A(a[44]), .B(b[15]), .Z(n1490) );
  XNOR U2900 ( .A(n1495), .B(n1144), .Z(n1146) );
  XOR U2901 ( .A(n1496), .B(n1497), .Z(n1144) );
  ANDN U2902 ( .B(n1498), .A(n1499), .Z(n1496) );
  AND U2903 ( .A(b[14]), .B(a[45]), .Z(n1495) );
  XNOR U2904 ( .A(n1500), .B(n1149), .Z(n1151) );
  XOR U2905 ( .A(n1501), .B(n1502), .Z(n1149) );
  ANDN U2906 ( .B(n1503), .A(n1504), .Z(n1501) );
  AND U2907 ( .A(b[13]), .B(a[46]), .Z(n1500) );
  XNOR U2908 ( .A(n1505), .B(n1154), .Z(n1156) );
  XOR U2909 ( .A(n1506), .B(n1507), .Z(n1154) );
  ANDN U2910 ( .B(n1508), .A(n1509), .Z(n1506) );
  AND U2911 ( .A(b[12]), .B(a[47]), .Z(n1505) );
  XNOR U2912 ( .A(n1510), .B(n1159), .Z(n1161) );
  XOR U2913 ( .A(n1511), .B(n1512), .Z(n1159) );
  ANDN U2914 ( .B(n1513), .A(n1514), .Z(n1511) );
  AND U2915 ( .A(b[11]), .B(a[48]), .Z(n1510) );
  XNOR U2916 ( .A(n1515), .B(n1164), .Z(n1166) );
  XOR U2917 ( .A(n1516), .B(n1517), .Z(n1164) );
  ANDN U2918 ( .B(n1518), .A(n1519), .Z(n1516) );
  AND U2919 ( .A(a[49]), .B(b[10]), .Z(n1515) );
  XNOR U2920 ( .A(n1520), .B(n1169), .Z(n1171) );
  XOR U2921 ( .A(n1521), .B(n1522), .Z(n1169) );
  ANDN U2922 ( .B(n1523), .A(n1524), .Z(n1521) );
  AND U2923 ( .A(b[9]), .B(a[50]), .Z(n1520) );
  XNOR U2924 ( .A(n1525), .B(n1174), .Z(n1176) );
  XOR U2925 ( .A(n1526), .B(n1527), .Z(n1174) );
  ANDN U2926 ( .B(n1528), .A(n1529), .Z(n1526) );
  AND U2927 ( .A(b[8]), .B(a[51]), .Z(n1525) );
  XNOR U2928 ( .A(n1530), .B(n1179), .Z(n1181) );
  XOR U2929 ( .A(n1531), .B(n1532), .Z(n1179) );
  ANDN U2930 ( .B(n1533), .A(n1534), .Z(n1531) );
  AND U2931 ( .A(b[7]), .B(a[52]), .Z(n1530) );
  XNOR U2932 ( .A(n1535), .B(n1184), .Z(n1186) );
  XOR U2933 ( .A(n1536), .B(n1537), .Z(n1184) );
  ANDN U2934 ( .B(n1538), .A(n1539), .Z(n1536) );
  AND U2935 ( .A(b[6]), .B(a[53]), .Z(n1535) );
  XNOR U2936 ( .A(n1540), .B(n1189), .Z(n1191) );
  XOR U2937 ( .A(n1541), .B(n1542), .Z(n1189) );
  ANDN U2938 ( .B(n1543), .A(n1544), .Z(n1541) );
  AND U2939 ( .A(b[5]), .B(a[54]), .Z(n1540) );
  XNOR U2940 ( .A(n1545), .B(n1194), .Z(n1196) );
  XOR U2941 ( .A(n1546), .B(n1547), .Z(n1194) );
  ANDN U2942 ( .B(n1548), .A(n1549), .Z(n1546) );
  AND U2943 ( .A(b[4]), .B(a[55]), .Z(n1545) );
  XNOR U2944 ( .A(n1550), .B(n1551), .Z(n1208) );
  NANDN U2945 ( .A(n1552), .B(n1553), .Z(n1551) );
  XNOR U2946 ( .A(n1554), .B(n1199), .Z(n1201) );
  XNOR U2947 ( .A(n1555), .B(n1556), .Z(n1199) );
  AND U2948 ( .A(n1557), .B(n1558), .Z(n1555) );
  AND U2949 ( .A(b[3]), .B(a[56]), .Z(n1554) );
  NAND U2950 ( .A(a[59]), .B(b[0]), .Z(n862) );
  XNOR U2951 ( .A(n1216), .B(n1217), .Z(c[58]) );
  XNOR U2952 ( .A(n1552), .B(n1553), .Z(n1217) );
  XOR U2953 ( .A(n1550), .B(n1559), .Z(n1553) );
  NAND U2954 ( .A(b[1]), .B(a[57]), .Z(n1559) );
  XOR U2955 ( .A(n1558), .B(n1560), .Z(n1552) );
  XOR U2956 ( .A(n1550), .B(n1557), .Z(n1560) );
  XNOR U2957 ( .A(n1561), .B(n1556), .Z(n1557) );
  AND U2958 ( .A(b[2]), .B(a[56]), .Z(n1561) );
  NANDN U2959 ( .A(n1562), .B(n1563), .Z(n1550) );
  XOR U2960 ( .A(n1556), .B(n1548), .Z(n1564) );
  XNOR U2961 ( .A(n1547), .B(n1543), .Z(n1565) );
  XNOR U2962 ( .A(n1542), .B(n1538), .Z(n1566) );
  XNOR U2963 ( .A(n1537), .B(n1533), .Z(n1567) );
  XNOR U2964 ( .A(n1532), .B(n1528), .Z(n1568) );
  XNOR U2965 ( .A(n1527), .B(n1523), .Z(n1569) );
  XNOR U2966 ( .A(n1522), .B(n1518), .Z(n1570) );
  XNOR U2967 ( .A(n1517), .B(n1513), .Z(n1571) );
  XNOR U2968 ( .A(n1512), .B(n1508), .Z(n1572) );
  XNOR U2969 ( .A(n1507), .B(n1503), .Z(n1573) );
  XNOR U2970 ( .A(n1502), .B(n1498), .Z(n1574) );
  XNOR U2971 ( .A(n1497), .B(n1493), .Z(n1575) );
  XNOR U2972 ( .A(n1492), .B(n1488), .Z(n1576) );
  XNOR U2973 ( .A(n1487), .B(n1483), .Z(n1577) );
  XNOR U2974 ( .A(n1482), .B(n1478), .Z(n1578) );
  XNOR U2975 ( .A(n1477), .B(n1473), .Z(n1579) );
  XNOR U2976 ( .A(n1472), .B(n1468), .Z(n1580) );
  XNOR U2977 ( .A(n1467), .B(n1463), .Z(n1581) );
  XNOR U2978 ( .A(n1462), .B(n1458), .Z(n1582) );
  XNOR U2979 ( .A(n1449), .B(n1448), .Z(n1583) );
  XOR U2980 ( .A(n1584), .B(n1447), .Z(n1448) );
  AND U2981 ( .A(b[22]), .B(a[36]), .Z(n1584) );
  XNOR U2982 ( .A(n1447), .B(n1453), .Z(n1585) );
  XNOR U2983 ( .A(n1452), .B(n1444), .Z(n1586) );
  XNOR U2984 ( .A(n1443), .B(n1439), .Z(n1587) );
  XNOR U2985 ( .A(n1438), .B(n1434), .Z(n1588) );
  XNOR U2986 ( .A(n1433), .B(n1429), .Z(n1589) );
  XNOR U2987 ( .A(n1420), .B(n1419), .Z(n1590) );
  XOR U2988 ( .A(n1591), .B(n1418), .Z(n1419) );
  AND U2989 ( .A(b[28]), .B(a[30]), .Z(n1591) );
  XNOR U2990 ( .A(n1418), .B(n1424), .Z(n1592) );
  XNOR U2991 ( .A(n1423), .B(n1415), .Z(n1593) );
  XNOR U2992 ( .A(n1414), .B(n1410), .Z(n1594) );
  XNOR U2993 ( .A(n1409), .B(n1405), .Z(n1595) );
  XNOR U2994 ( .A(n1404), .B(n1400), .Z(n1596) );
  XNOR U2995 ( .A(n1391), .B(n1390), .Z(n1597) );
  XOR U2996 ( .A(n1598), .B(n1389), .Z(n1390) );
  AND U2997 ( .A(b[34]), .B(a[24]), .Z(n1598) );
  XNOR U2998 ( .A(n1389), .B(n1395), .Z(n1599) );
  XNOR U2999 ( .A(n1394), .B(n1386), .Z(n1600) );
  XNOR U3000 ( .A(n1385), .B(n1381), .Z(n1601) );
  XNOR U3001 ( .A(n1380), .B(n1376), .Z(n1602) );
  XNOR U3002 ( .A(n1375), .B(n1371), .Z(n1603) );
  XNOR U3003 ( .A(n1362), .B(n1361), .Z(n1604) );
  XOR U3004 ( .A(n1605), .B(n1360), .Z(n1361) );
  AND U3005 ( .A(b[40]), .B(a[18]), .Z(n1605) );
  XNOR U3006 ( .A(n1360), .B(n1366), .Z(n1606) );
  XNOR U3007 ( .A(n1365), .B(n1357), .Z(n1607) );
  XNOR U3008 ( .A(n1356), .B(n1352), .Z(n1608) );
  XNOR U3009 ( .A(n1351), .B(n1347), .Z(n1609) );
  XNOR U3010 ( .A(n1346), .B(n1342), .Z(n1610) );
  XNOR U3011 ( .A(n1333), .B(n1332), .Z(n1611) );
  XOR U3012 ( .A(n1612), .B(n1331), .Z(n1332) );
  AND U3013 ( .A(b[46]), .B(a[12]), .Z(n1612) );
  XNOR U3014 ( .A(n1331), .B(n1337), .Z(n1613) );
  XNOR U3015 ( .A(n1336), .B(n1328), .Z(n1614) );
  XNOR U3016 ( .A(n1327), .B(n1323), .Z(n1615) );
  XNOR U3017 ( .A(n1322), .B(n1318), .Z(n1616) );
  XNOR U3018 ( .A(n1317), .B(n1313), .Z(n1617) );
  XNOR U3019 ( .A(n1304), .B(n1303), .Z(n1618) );
  XOR U3020 ( .A(n1619), .B(n1302), .Z(n1303) );
  AND U3021 ( .A(a[6]), .B(b[52]), .Z(n1619) );
  XNOR U3022 ( .A(n1302), .B(n1308), .Z(n1620) );
  XNOR U3023 ( .A(n1307), .B(n1299), .Z(n1621) );
  XNOR U3024 ( .A(n1298), .B(n1294), .Z(n1622) );
  XNOR U3025 ( .A(n1293), .B(n1289), .Z(n1623) );
  XNOR U3026 ( .A(n1288), .B(n1284), .Z(n1624) );
  XOR U3027 ( .A(n1625), .B(n1283), .Z(n1284) );
  AND U3028 ( .A(a[0]), .B(b[58]), .Z(n1625) );
  XNOR U3029 ( .A(n1626), .B(n1283), .Z(n1285) );
  XNOR U3030 ( .A(n1627), .B(n1628), .Z(n1283) );
  ANDN U3031 ( .B(n1629), .A(n1630), .Z(n1627) );
  AND U3032 ( .A(a[1]), .B(b[57]), .Z(n1626) );
  XNOR U3033 ( .A(n1631), .B(n1288), .Z(n1290) );
  XOR U3034 ( .A(n1632), .B(n1633), .Z(n1288) );
  ANDN U3035 ( .B(n1634), .A(n1635), .Z(n1632) );
  AND U3036 ( .A(a[2]), .B(b[56]), .Z(n1631) );
  XNOR U3037 ( .A(n1636), .B(n1293), .Z(n1295) );
  XOR U3038 ( .A(n1637), .B(n1638), .Z(n1293) );
  ANDN U3039 ( .B(n1639), .A(n1640), .Z(n1637) );
  AND U3040 ( .A(a[3]), .B(b[55]), .Z(n1636) );
  XNOR U3041 ( .A(n1641), .B(n1298), .Z(n1300) );
  XOR U3042 ( .A(n1642), .B(n1643), .Z(n1298) );
  ANDN U3043 ( .B(n1644), .A(n1645), .Z(n1642) );
  AND U3044 ( .A(a[4]), .B(b[54]), .Z(n1641) );
  XOR U3045 ( .A(n1646), .B(n1647), .Z(n1302) );
  AND U3046 ( .A(n1648), .B(n1649), .Z(n1646) );
  XNOR U3047 ( .A(n1650), .B(n1307), .Z(n1309) );
  XOR U3048 ( .A(n1651), .B(n1652), .Z(n1307) );
  ANDN U3049 ( .B(n1653), .A(n1654), .Z(n1651) );
  AND U3050 ( .A(a[5]), .B(b[53]), .Z(n1650) );
  XOR U3051 ( .A(n1655), .B(n1312), .Z(n1314) );
  XOR U3052 ( .A(n1656), .B(n1657), .Z(n1312) );
  ANDN U3053 ( .B(n1658), .A(n1659), .Z(n1656) );
  AND U3054 ( .A(a[7]), .B(b[51]), .Z(n1655) );
  XNOR U3055 ( .A(n1660), .B(n1317), .Z(n1319) );
  XOR U3056 ( .A(n1661), .B(n1662), .Z(n1317) );
  ANDN U3057 ( .B(n1663), .A(n1664), .Z(n1661) );
  AND U3058 ( .A(a[8]), .B(b[50]), .Z(n1660) );
  XNOR U3059 ( .A(n1665), .B(n1322), .Z(n1324) );
  XOR U3060 ( .A(n1666), .B(n1667), .Z(n1322) );
  ANDN U3061 ( .B(n1668), .A(n1669), .Z(n1666) );
  AND U3062 ( .A(a[9]), .B(b[49]), .Z(n1665) );
  XNOR U3063 ( .A(n1670), .B(n1327), .Z(n1329) );
  XOR U3064 ( .A(n1671), .B(n1672), .Z(n1327) );
  ANDN U3065 ( .B(n1673), .A(n1674), .Z(n1671) );
  AND U3066 ( .A(b[48]), .B(a[10]), .Z(n1670) );
  XOR U3067 ( .A(n1675), .B(n1676), .Z(n1331) );
  AND U3068 ( .A(n1677), .B(n1678), .Z(n1675) );
  XNOR U3069 ( .A(n1679), .B(n1336), .Z(n1338) );
  XOR U3070 ( .A(n1680), .B(n1681), .Z(n1336) );
  ANDN U3071 ( .B(n1682), .A(n1683), .Z(n1680) );
  AND U3072 ( .A(b[47]), .B(a[11]), .Z(n1679) );
  XOR U3073 ( .A(n1684), .B(n1341), .Z(n1343) );
  XOR U3074 ( .A(n1685), .B(n1686), .Z(n1341) );
  ANDN U3075 ( .B(n1687), .A(n1688), .Z(n1685) );
  AND U3076 ( .A(a[13]), .B(b[45]), .Z(n1684) );
  XNOR U3077 ( .A(n1689), .B(n1346), .Z(n1348) );
  XOR U3078 ( .A(n1690), .B(n1691), .Z(n1346) );
  ANDN U3079 ( .B(n1692), .A(n1693), .Z(n1690) );
  AND U3080 ( .A(b[44]), .B(a[14]), .Z(n1689) );
  XNOR U3081 ( .A(n1694), .B(n1351), .Z(n1353) );
  XOR U3082 ( .A(n1695), .B(n1696), .Z(n1351) );
  ANDN U3083 ( .B(n1697), .A(n1698), .Z(n1695) );
  AND U3084 ( .A(b[43]), .B(a[15]), .Z(n1694) );
  XNOR U3085 ( .A(n1699), .B(n1356), .Z(n1358) );
  XOR U3086 ( .A(n1700), .B(n1701), .Z(n1356) );
  ANDN U3087 ( .B(n1702), .A(n1703), .Z(n1700) );
  AND U3088 ( .A(b[42]), .B(a[16]), .Z(n1699) );
  XOR U3089 ( .A(n1704), .B(n1705), .Z(n1360) );
  AND U3090 ( .A(n1706), .B(n1707), .Z(n1704) );
  XNOR U3091 ( .A(n1708), .B(n1365), .Z(n1367) );
  XOR U3092 ( .A(n1709), .B(n1710), .Z(n1365) );
  ANDN U3093 ( .B(n1711), .A(n1712), .Z(n1709) );
  AND U3094 ( .A(b[41]), .B(a[17]), .Z(n1708) );
  XOR U3095 ( .A(n1713), .B(n1370), .Z(n1372) );
  XOR U3096 ( .A(n1714), .B(n1715), .Z(n1370) );
  ANDN U3097 ( .B(n1716), .A(n1717), .Z(n1714) );
  AND U3098 ( .A(a[19]), .B(b[39]), .Z(n1713) );
  XNOR U3099 ( .A(n1718), .B(n1375), .Z(n1377) );
  XOR U3100 ( .A(n1719), .B(n1720), .Z(n1375) );
  ANDN U3101 ( .B(n1721), .A(n1722), .Z(n1719) );
  AND U3102 ( .A(b[38]), .B(a[20]), .Z(n1718) );
  XNOR U3103 ( .A(n1723), .B(n1380), .Z(n1382) );
  XOR U3104 ( .A(n1724), .B(n1725), .Z(n1380) );
  ANDN U3105 ( .B(n1726), .A(n1727), .Z(n1724) );
  AND U3106 ( .A(b[37]), .B(a[21]), .Z(n1723) );
  XNOR U3107 ( .A(n1728), .B(n1385), .Z(n1387) );
  XOR U3108 ( .A(n1729), .B(n1730), .Z(n1385) );
  ANDN U3109 ( .B(n1731), .A(n1732), .Z(n1729) );
  AND U3110 ( .A(b[36]), .B(a[22]), .Z(n1728) );
  XOR U3111 ( .A(n1733), .B(n1734), .Z(n1389) );
  AND U3112 ( .A(n1735), .B(n1736), .Z(n1733) );
  XNOR U3113 ( .A(n1737), .B(n1394), .Z(n1396) );
  XOR U3114 ( .A(n1738), .B(n1739), .Z(n1394) );
  ANDN U3115 ( .B(n1740), .A(n1741), .Z(n1738) );
  AND U3116 ( .A(b[35]), .B(a[23]), .Z(n1737) );
  XOR U3117 ( .A(n1742), .B(n1399), .Z(n1401) );
  XOR U3118 ( .A(n1743), .B(n1744), .Z(n1399) );
  ANDN U3119 ( .B(n1745), .A(n1746), .Z(n1743) );
  AND U3120 ( .A(a[25]), .B(b[33]), .Z(n1742) );
  XNOR U3121 ( .A(n1747), .B(n1404), .Z(n1406) );
  XOR U3122 ( .A(n1748), .B(n1749), .Z(n1404) );
  ANDN U3123 ( .B(n1750), .A(n1751), .Z(n1748) );
  AND U3124 ( .A(b[32]), .B(a[26]), .Z(n1747) );
  XNOR U3125 ( .A(n1752), .B(n1409), .Z(n1411) );
  XOR U3126 ( .A(n1753), .B(n1754), .Z(n1409) );
  ANDN U3127 ( .B(n1755), .A(n1756), .Z(n1753) );
  AND U3128 ( .A(b[31]), .B(a[27]), .Z(n1752) );
  XNOR U3129 ( .A(n1757), .B(n1414), .Z(n1416) );
  XOR U3130 ( .A(n1758), .B(n1759), .Z(n1414) );
  ANDN U3131 ( .B(n1760), .A(n1761), .Z(n1758) );
  AND U3132 ( .A(b[30]), .B(a[28]), .Z(n1757) );
  XOR U3133 ( .A(n1762), .B(n1763), .Z(n1418) );
  AND U3134 ( .A(n1764), .B(n1765), .Z(n1762) );
  XNOR U3135 ( .A(n1766), .B(n1423), .Z(n1425) );
  XOR U3136 ( .A(n1767), .B(n1768), .Z(n1423) );
  ANDN U3137 ( .B(n1769), .A(n1770), .Z(n1767) );
  AND U3138 ( .A(b[29]), .B(a[29]), .Z(n1766) );
  XOR U3139 ( .A(n1771), .B(n1428), .Z(n1430) );
  XOR U3140 ( .A(n1772), .B(n1773), .Z(n1428) );
  ANDN U3141 ( .B(n1774), .A(n1775), .Z(n1772) );
  AND U3142 ( .A(a[31]), .B(b[27]), .Z(n1771) );
  XNOR U3143 ( .A(n1776), .B(n1433), .Z(n1435) );
  XOR U3144 ( .A(n1777), .B(n1778), .Z(n1433) );
  ANDN U3145 ( .B(n1779), .A(n1780), .Z(n1777) );
  AND U3146 ( .A(b[26]), .B(a[32]), .Z(n1776) );
  XNOR U3147 ( .A(n1781), .B(n1438), .Z(n1440) );
  XOR U3148 ( .A(n1782), .B(n1783), .Z(n1438) );
  ANDN U3149 ( .B(n1784), .A(n1785), .Z(n1782) );
  AND U3150 ( .A(b[25]), .B(a[33]), .Z(n1781) );
  XNOR U3151 ( .A(n1786), .B(n1443), .Z(n1445) );
  XOR U3152 ( .A(n1787), .B(n1788), .Z(n1443) );
  ANDN U3153 ( .B(n1789), .A(n1790), .Z(n1787) );
  AND U3154 ( .A(b[24]), .B(a[34]), .Z(n1786) );
  XOR U3155 ( .A(n1791), .B(n1792), .Z(n1447) );
  AND U3156 ( .A(n1793), .B(n1794), .Z(n1791) );
  XNOR U3157 ( .A(n1795), .B(n1452), .Z(n1454) );
  XOR U3158 ( .A(n1796), .B(n1797), .Z(n1452) );
  ANDN U3159 ( .B(n1798), .A(n1799), .Z(n1796) );
  AND U3160 ( .A(b[23]), .B(a[35]), .Z(n1795) );
  XOR U3161 ( .A(n1800), .B(n1457), .Z(n1459) );
  XOR U3162 ( .A(n1801), .B(n1802), .Z(n1457) );
  ANDN U3163 ( .B(n1803), .A(n1804), .Z(n1801) );
  AND U3164 ( .A(a[37]), .B(b[21]), .Z(n1800) );
  XNOR U3165 ( .A(n1805), .B(n1462), .Z(n1464) );
  XOR U3166 ( .A(n1806), .B(n1807), .Z(n1462) );
  ANDN U3167 ( .B(n1808), .A(n1809), .Z(n1806) );
  AND U3168 ( .A(b[20]), .B(a[38]), .Z(n1805) );
  XNOR U3169 ( .A(n1810), .B(n1467), .Z(n1469) );
  XOR U3170 ( .A(n1811), .B(n1812), .Z(n1467) );
  ANDN U3171 ( .B(n1813), .A(n1814), .Z(n1811) );
  AND U3172 ( .A(b[19]), .B(a[39]), .Z(n1810) );
  XNOR U3173 ( .A(n1815), .B(n1472), .Z(n1474) );
  XOR U3174 ( .A(n1816), .B(n1817), .Z(n1472) );
  ANDN U3175 ( .B(n1818), .A(n1819), .Z(n1816) );
  AND U3176 ( .A(b[18]), .B(a[40]), .Z(n1815) );
  XNOR U3177 ( .A(n1820), .B(n1477), .Z(n1479) );
  XOR U3178 ( .A(n1821), .B(n1822), .Z(n1477) );
  ANDN U3179 ( .B(n1823), .A(n1824), .Z(n1821) );
  AND U3180 ( .A(b[17]), .B(a[41]), .Z(n1820) );
  XNOR U3181 ( .A(n1825), .B(n1482), .Z(n1484) );
  XOR U3182 ( .A(n1826), .B(n1827), .Z(n1482) );
  ANDN U3183 ( .B(n1828), .A(n1829), .Z(n1826) );
  AND U3184 ( .A(b[16]), .B(a[42]), .Z(n1825) );
  XNOR U3185 ( .A(n1830), .B(n1487), .Z(n1489) );
  XOR U3186 ( .A(n1831), .B(n1832), .Z(n1487) );
  ANDN U3187 ( .B(n1833), .A(n1834), .Z(n1831) );
  AND U3188 ( .A(a[43]), .B(b[15]), .Z(n1830) );
  XNOR U3189 ( .A(n1835), .B(n1492), .Z(n1494) );
  XOR U3190 ( .A(n1836), .B(n1837), .Z(n1492) );
  ANDN U3191 ( .B(n1838), .A(n1839), .Z(n1836) );
  AND U3192 ( .A(b[14]), .B(a[44]), .Z(n1835) );
  XNOR U3193 ( .A(n1840), .B(n1497), .Z(n1499) );
  XOR U3194 ( .A(n1841), .B(n1842), .Z(n1497) );
  ANDN U3195 ( .B(n1843), .A(n1844), .Z(n1841) );
  AND U3196 ( .A(b[13]), .B(a[45]), .Z(n1840) );
  XNOR U3197 ( .A(n1845), .B(n1502), .Z(n1504) );
  XOR U3198 ( .A(n1846), .B(n1847), .Z(n1502) );
  ANDN U3199 ( .B(n1848), .A(n1849), .Z(n1846) );
  AND U3200 ( .A(b[12]), .B(a[46]), .Z(n1845) );
  XNOR U3201 ( .A(n1850), .B(n1507), .Z(n1509) );
  XOR U3202 ( .A(n1851), .B(n1852), .Z(n1507) );
  ANDN U3203 ( .B(n1853), .A(n1854), .Z(n1851) );
  AND U3204 ( .A(b[11]), .B(a[47]), .Z(n1850) );
  XNOR U3205 ( .A(n1855), .B(n1512), .Z(n1514) );
  XOR U3206 ( .A(n1856), .B(n1857), .Z(n1512) );
  ANDN U3207 ( .B(n1858), .A(n1859), .Z(n1856) );
  AND U3208 ( .A(b[10]), .B(a[48]), .Z(n1855) );
  XNOR U3209 ( .A(n1860), .B(n1517), .Z(n1519) );
  XOR U3210 ( .A(n1861), .B(n1862), .Z(n1517) );
  ANDN U3211 ( .B(n1863), .A(n1864), .Z(n1861) );
  AND U3212 ( .A(b[9]), .B(a[49]), .Z(n1860) );
  XNOR U3213 ( .A(n1865), .B(n1522), .Z(n1524) );
  XOR U3214 ( .A(n1866), .B(n1867), .Z(n1522) );
  ANDN U3215 ( .B(n1868), .A(n1869), .Z(n1866) );
  AND U3216 ( .A(b[8]), .B(a[50]), .Z(n1865) );
  XNOR U3217 ( .A(n1870), .B(n1527), .Z(n1529) );
  XOR U3218 ( .A(n1871), .B(n1872), .Z(n1527) );
  ANDN U3219 ( .B(n1873), .A(n1874), .Z(n1871) );
  AND U3220 ( .A(b[7]), .B(a[51]), .Z(n1870) );
  XNOR U3221 ( .A(n1875), .B(n1532), .Z(n1534) );
  XOR U3222 ( .A(n1876), .B(n1877), .Z(n1532) );
  ANDN U3223 ( .B(n1878), .A(n1879), .Z(n1876) );
  AND U3224 ( .A(b[6]), .B(a[52]), .Z(n1875) );
  XNOR U3225 ( .A(n1880), .B(n1537), .Z(n1539) );
  XOR U3226 ( .A(n1881), .B(n1882), .Z(n1537) );
  ANDN U3227 ( .B(n1883), .A(n1884), .Z(n1881) );
  AND U3228 ( .A(b[5]), .B(a[53]), .Z(n1880) );
  XNOR U3229 ( .A(n1885), .B(n1542), .Z(n1544) );
  XOR U3230 ( .A(n1886), .B(n1887), .Z(n1542) );
  ANDN U3231 ( .B(n1888), .A(n1889), .Z(n1886) );
  AND U3232 ( .A(b[4]), .B(a[54]), .Z(n1885) );
  XNOR U3233 ( .A(n1890), .B(n1891), .Z(n1556) );
  NANDN U3234 ( .A(n1892), .B(n1893), .Z(n1891) );
  XNOR U3235 ( .A(n1894), .B(n1547), .Z(n1549) );
  XNOR U3236 ( .A(n1895), .B(n1896), .Z(n1547) );
  AND U3237 ( .A(n1897), .B(n1898), .Z(n1895) );
  AND U3238 ( .A(b[3]), .B(a[55]), .Z(n1894) );
  NAND U3239 ( .A(a[58]), .B(b[0]), .Z(n1216) );
  XNOR U3240 ( .A(n1562), .B(n1563), .Z(c[57]) );
  XNOR U3241 ( .A(n1892), .B(n1893), .Z(n1563) );
  XOR U3242 ( .A(n1890), .B(n1899), .Z(n1893) );
  NAND U3243 ( .A(b[1]), .B(a[56]), .Z(n1899) );
  XOR U3244 ( .A(n1898), .B(n1900), .Z(n1892) );
  XOR U3245 ( .A(n1890), .B(n1897), .Z(n1900) );
  XNOR U3246 ( .A(n1901), .B(n1896), .Z(n1897) );
  AND U3247 ( .A(b[2]), .B(a[55]), .Z(n1901) );
  NANDN U3248 ( .A(n1902), .B(n1903), .Z(n1890) );
  XOR U3249 ( .A(n1896), .B(n1888), .Z(n1904) );
  XNOR U3250 ( .A(n1887), .B(n1883), .Z(n1905) );
  XNOR U3251 ( .A(n1882), .B(n1878), .Z(n1906) );
  XNOR U3252 ( .A(n1877), .B(n1873), .Z(n1907) );
  XNOR U3253 ( .A(n1872), .B(n1868), .Z(n1908) );
  XNOR U3254 ( .A(n1867), .B(n1863), .Z(n1909) );
  XNOR U3255 ( .A(n1862), .B(n1858), .Z(n1910) );
  XNOR U3256 ( .A(n1857), .B(n1853), .Z(n1911) );
  XNOR U3257 ( .A(n1852), .B(n1848), .Z(n1912) );
  XNOR U3258 ( .A(n1847), .B(n1843), .Z(n1913) );
  XNOR U3259 ( .A(n1842), .B(n1838), .Z(n1914) );
  XNOR U3260 ( .A(n1837), .B(n1833), .Z(n1915) );
  XNOR U3261 ( .A(n1832), .B(n1828), .Z(n1916) );
  XNOR U3262 ( .A(n1917), .B(n1918), .Z(n1828) );
  XNOR U3263 ( .A(n1827), .B(n1823), .Z(n1918) );
  XNOR U3264 ( .A(n1822), .B(n1818), .Z(n1919) );
  XNOR U3265 ( .A(n1817), .B(n1813), .Z(n1920) );
  XNOR U3266 ( .A(n1812), .B(n1808), .Z(n1921) );
  XNOR U3267 ( .A(n1807), .B(n1803), .Z(n1922) );
  XNOR U3268 ( .A(n1794), .B(n1793), .Z(n1923) );
  XOR U3269 ( .A(n1924), .B(n1792), .Z(n1793) );
  AND U3270 ( .A(b[21]), .B(a[36]), .Z(n1924) );
  XNOR U3271 ( .A(n1792), .B(n1798), .Z(n1925) );
  XNOR U3272 ( .A(n1797), .B(n1789), .Z(n1926) );
  XNOR U3273 ( .A(n1788), .B(n1784), .Z(n1927) );
  XNOR U3274 ( .A(n1783), .B(n1779), .Z(n1928) );
  XNOR U3275 ( .A(n1778), .B(n1774), .Z(n1929) );
  XNOR U3276 ( .A(n1765), .B(n1764), .Z(n1930) );
  XOR U3277 ( .A(n1931), .B(n1763), .Z(n1764) );
  AND U3278 ( .A(b[27]), .B(a[30]), .Z(n1931) );
  XNOR U3279 ( .A(n1763), .B(n1769), .Z(n1932) );
  XNOR U3280 ( .A(n1768), .B(n1760), .Z(n1933) );
  XNOR U3281 ( .A(n1759), .B(n1755), .Z(n1934) );
  XNOR U3282 ( .A(n1754), .B(n1750), .Z(n1935) );
  XNOR U3283 ( .A(n1749), .B(n1745), .Z(n1936) );
  XNOR U3284 ( .A(n1736), .B(n1735), .Z(n1937) );
  XOR U3285 ( .A(n1938), .B(n1734), .Z(n1735) );
  AND U3286 ( .A(b[33]), .B(a[24]), .Z(n1938) );
  XNOR U3287 ( .A(n1734), .B(n1740), .Z(n1939) );
  XNOR U3288 ( .A(n1739), .B(n1731), .Z(n1940) );
  XNOR U3289 ( .A(n1730), .B(n1726), .Z(n1941) );
  XNOR U3290 ( .A(n1725), .B(n1721), .Z(n1942) );
  XNOR U3291 ( .A(n1720), .B(n1716), .Z(n1943) );
  XNOR U3292 ( .A(n1707), .B(n1706), .Z(n1944) );
  XOR U3293 ( .A(n1945), .B(n1705), .Z(n1706) );
  AND U3294 ( .A(b[39]), .B(a[18]), .Z(n1945) );
  XNOR U3295 ( .A(n1705), .B(n1711), .Z(n1946) );
  XNOR U3296 ( .A(n1710), .B(n1702), .Z(n1947) );
  XNOR U3297 ( .A(n1701), .B(n1697), .Z(n1948) );
  XNOR U3298 ( .A(n1696), .B(n1692), .Z(n1949) );
  XNOR U3299 ( .A(n1691), .B(n1687), .Z(n1950) );
  XNOR U3300 ( .A(n1678), .B(n1677), .Z(n1951) );
  XOR U3301 ( .A(n1952), .B(n1676), .Z(n1677) );
  AND U3302 ( .A(b[45]), .B(a[12]), .Z(n1952) );
  XNOR U3303 ( .A(n1676), .B(n1682), .Z(n1953) );
  XNOR U3304 ( .A(n1681), .B(n1673), .Z(n1954) );
  XNOR U3305 ( .A(n1672), .B(n1668), .Z(n1955) );
  XNOR U3306 ( .A(n1667), .B(n1663), .Z(n1956) );
  XNOR U3307 ( .A(n1662), .B(n1658), .Z(n1957) );
  XNOR U3308 ( .A(n1649), .B(n1648), .Z(n1958) );
  XOR U3309 ( .A(n1959), .B(n1647), .Z(n1648) );
  AND U3310 ( .A(a[6]), .B(b[51]), .Z(n1959) );
  XNOR U3311 ( .A(n1647), .B(n1653), .Z(n1960) );
  XNOR U3312 ( .A(n1652), .B(n1644), .Z(n1961) );
  XNOR U3313 ( .A(n1643), .B(n1639), .Z(n1962) );
  XNOR U3314 ( .A(n1638), .B(n1634), .Z(n1963) );
  XNOR U3315 ( .A(n1633), .B(n1629), .Z(n1964) );
  XNOR U3316 ( .A(n1965), .B(n1628), .Z(n1629) );
  AND U3317 ( .A(a[0]), .B(b[57]), .Z(n1965) );
  XOR U3318 ( .A(n1966), .B(n1628), .Z(n1630) );
  XNOR U3319 ( .A(n1967), .B(n1968), .Z(n1628) );
  ANDN U3320 ( .B(n1969), .A(n1970), .Z(n1967) );
  AND U3321 ( .A(a[1]), .B(b[56]), .Z(n1966) );
  XNOR U3322 ( .A(n1971), .B(n1633), .Z(n1635) );
  XOR U3323 ( .A(n1972), .B(n1973), .Z(n1633) );
  ANDN U3324 ( .B(n1974), .A(n1975), .Z(n1972) );
  AND U3325 ( .A(a[2]), .B(b[55]), .Z(n1971) );
  XNOR U3326 ( .A(n1976), .B(n1638), .Z(n1640) );
  XOR U3327 ( .A(n1977), .B(n1978), .Z(n1638) );
  ANDN U3328 ( .B(n1979), .A(n1980), .Z(n1977) );
  AND U3329 ( .A(a[3]), .B(b[54]), .Z(n1976) );
  XNOR U3330 ( .A(n1981), .B(n1643), .Z(n1645) );
  XOR U3331 ( .A(n1982), .B(n1983), .Z(n1643) );
  ANDN U3332 ( .B(n1984), .A(n1985), .Z(n1982) );
  AND U3333 ( .A(a[4]), .B(b[53]), .Z(n1981) );
  XOR U3334 ( .A(n1986), .B(n1987), .Z(n1647) );
  AND U3335 ( .A(n1988), .B(n1989), .Z(n1986) );
  XNOR U3336 ( .A(n1990), .B(n1652), .Z(n1654) );
  XOR U3337 ( .A(n1991), .B(n1992), .Z(n1652) );
  ANDN U3338 ( .B(n1993), .A(n1994), .Z(n1991) );
  AND U3339 ( .A(a[5]), .B(b[52]), .Z(n1990) );
  XOR U3340 ( .A(n1995), .B(n1657), .Z(n1659) );
  XOR U3341 ( .A(n1996), .B(n1997), .Z(n1657) );
  ANDN U3342 ( .B(n1998), .A(n1999), .Z(n1996) );
  AND U3343 ( .A(a[7]), .B(b[50]), .Z(n1995) );
  XNOR U3344 ( .A(n2000), .B(n1662), .Z(n1664) );
  XOR U3345 ( .A(n2001), .B(n2002), .Z(n1662) );
  ANDN U3346 ( .B(n2003), .A(n2004), .Z(n2001) );
  AND U3347 ( .A(a[8]), .B(b[49]), .Z(n2000) );
  XNOR U3348 ( .A(n2005), .B(n1667), .Z(n1669) );
  XOR U3349 ( .A(n2006), .B(n2007), .Z(n1667) );
  ANDN U3350 ( .B(n2008), .A(n2009), .Z(n2006) );
  AND U3351 ( .A(a[9]), .B(b[48]), .Z(n2005) );
  XNOR U3352 ( .A(n2010), .B(n1672), .Z(n1674) );
  XOR U3353 ( .A(n2011), .B(n2012), .Z(n1672) );
  ANDN U3354 ( .B(n2013), .A(n2014), .Z(n2011) );
  AND U3355 ( .A(b[47]), .B(a[10]), .Z(n2010) );
  XOR U3356 ( .A(n2015), .B(n2016), .Z(n1676) );
  AND U3357 ( .A(n2017), .B(n2018), .Z(n2015) );
  XNOR U3358 ( .A(n2019), .B(n1681), .Z(n1683) );
  XOR U3359 ( .A(n2020), .B(n2021), .Z(n1681) );
  ANDN U3360 ( .B(n2022), .A(n2023), .Z(n2020) );
  AND U3361 ( .A(b[46]), .B(a[11]), .Z(n2019) );
  XOR U3362 ( .A(n2024), .B(n1686), .Z(n1688) );
  XOR U3363 ( .A(n2025), .B(n2026), .Z(n1686) );
  ANDN U3364 ( .B(n2027), .A(n2028), .Z(n2025) );
  AND U3365 ( .A(b[44]), .B(a[13]), .Z(n2024) );
  XNOR U3366 ( .A(n2029), .B(n1691), .Z(n1693) );
  XOR U3367 ( .A(n2030), .B(n2031), .Z(n1691) );
  ANDN U3368 ( .B(n2032), .A(n2033), .Z(n2030) );
  AND U3369 ( .A(b[43]), .B(a[14]), .Z(n2029) );
  XNOR U3370 ( .A(n2034), .B(n1696), .Z(n1698) );
  XOR U3371 ( .A(n2035), .B(n2036), .Z(n1696) );
  ANDN U3372 ( .B(n2037), .A(n2038), .Z(n2035) );
  AND U3373 ( .A(b[42]), .B(a[15]), .Z(n2034) );
  XNOR U3374 ( .A(n2039), .B(n1701), .Z(n1703) );
  XOR U3375 ( .A(n2040), .B(n2041), .Z(n1701) );
  ANDN U3376 ( .B(n2042), .A(n2043), .Z(n2040) );
  AND U3377 ( .A(b[41]), .B(a[16]), .Z(n2039) );
  XOR U3378 ( .A(n2044), .B(n2045), .Z(n1705) );
  AND U3379 ( .A(n2046), .B(n2047), .Z(n2044) );
  XNOR U3380 ( .A(n2048), .B(n1710), .Z(n1712) );
  XOR U3381 ( .A(n2049), .B(n2050), .Z(n1710) );
  ANDN U3382 ( .B(n2051), .A(n2052), .Z(n2049) );
  AND U3383 ( .A(b[40]), .B(a[17]), .Z(n2048) );
  XOR U3384 ( .A(n2053), .B(n1715), .Z(n1717) );
  XOR U3385 ( .A(n2054), .B(n2055), .Z(n1715) );
  ANDN U3386 ( .B(n2056), .A(n2057), .Z(n2054) );
  AND U3387 ( .A(b[38]), .B(a[19]), .Z(n2053) );
  XNOR U3388 ( .A(n2058), .B(n1720), .Z(n1722) );
  XOR U3389 ( .A(n2059), .B(n2060), .Z(n1720) );
  ANDN U3390 ( .B(n2061), .A(n2062), .Z(n2059) );
  AND U3391 ( .A(b[37]), .B(a[20]), .Z(n2058) );
  XNOR U3392 ( .A(n2063), .B(n1725), .Z(n1727) );
  XOR U3393 ( .A(n2064), .B(n2065), .Z(n1725) );
  ANDN U3394 ( .B(n2066), .A(n2067), .Z(n2064) );
  AND U3395 ( .A(b[36]), .B(a[21]), .Z(n2063) );
  XNOR U3396 ( .A(n2068), .B(n1730), .Z(n1732) );
  XOR U3397 ( .A(n2069), .B(n2070), .Z(n1730) );
  ANDN U3398 ( .B(n2071), .A(n2072), .Z(n2069) );
  AND U3399 ( .A(b[35]), .B(a[22]), .Z(n2068) );
  XOR U3400 ( .A(n2073), .B(n2074), .Z(n1734) );
  AND U3401 ( .A(n2075), .B(n2076), .Z(n2073) );
  XNOR U3402 ( .A(n2077), .B(n1739), .Z(n1741) );
  XOR U3403 ( .A(n2078), .B(n2079), .Z(n1739) );
  ANDN U3404 ( .B(n2080), .A(n2081), .Z(n2078) );
  AND U3405 ( .A(b[34]), .B(a[23]), .Z(n2077) );
  XOR U3406 ( .A(n2082), .B(n1744), .Z(n1746) );
  XOR U3407 ( .A(n2083), .B(n2084), .Z(n1744) );
  ANDN U3408 ( .B(n2085), .A(n2086), .Z(n2083) );
  AND U3409 ( .A(b[32]), .B(a[25]), .Z(n2082) );
  XNOR U3410 ( .A(n2087), .B(n1749), .Z(n1751) );
  XOR U3411 ( .A(n2088), .B(n2089), .Z(n1749) );
  ANDN U3412 ( .B(n2090), .A(n2091), .Z(n2088) );
  AND U3413 ( .A(b[31]), .B(a[26]), .Z(n2087) );
  XNOR U3414 ( .A(n2092), .B(n1754), .Z(n1756) );
  XOR U3415 ( .A(n2093), .B(n2094), .Z(n1754) );
  ANDN U3416 ( .B(n2095), .A(n2096), .Z(n2093) );
  AND U3417 ( .A(b[30]), .B(a[27]), .Z(n2092) );
  XNOR U3418 ( .A(n2097), .B(n1759), .Z(n1761) );
  XOR U3419 ( .A(n2098), .B(n2099), .Z(n1759) );
  ANDN U3420 ( .B(n2100), .A(n2101), .Z(n2098) );
  AND U3421 ( .A(b[29]), .B(a[28]), .Z(n2097) );
  XOR U3422 ( .A(n2102), .B(n2103), .Z(n1763) );
  AND U3423 ( .A(n2104), .B(n2105), .Z(n2102) );
  XNOR U3424 ( .A(n2106), .B(n1768), .Z(n1770) );
  XOR U3425 ( .A(n2107), .B(n2108), .Z(n1768) );
  ANDN U3426 ( .B(n2109), .A(n2110), .Z(n2107) );
  AND U3427 ( .A(b[28]), .B(a[29]), .Z(n2106) );
  XOR U3428 ( .A(n2111), .B(n1773), .Z(n1775) );
  XOR U3429 ( .A(n2112), .B(n2113), .Z(n1773) );
  ANDN U3430 ( .B(n2114), .A(n2115), .Z(n2112) );
  AND U3431 ( .A(b[26]), .B(a[31]), .Z(n2111) );
  XNOR U3432 ( .A(n2116), .B(n1778), .Z(n1780) );
  XOR U3433 ( .A(n2117), .B(n2118), .Z(n1778) );
  ANDN U3434 ( .B(n2119), .A(n2120), .Z(n2117) );
  AND U3435 ( .A(b[25]), .B(a[32]), .Z(n2116) );
  XNOR U3436 ( .A(n2121), .B(n1783), .Z(n1785) );
  XOR U3437 ( .A(n2122), .B(n2123), .Z(n1783) );
  ANDN U3438 ( .B(n2124), .A(n2125), .Z(n2122) );
  AND U3439 ( .A(b[24]), .B(a[33]), .Z(n2121) );
  XNOR U3440 ( .A(n2126), .B(n1788), .Z(n1790) );
  XOR U3441 ( .A(n2127), .B(n2128), .Z(n1788) );
  ANDN U3442 ( .B(n2129), .A(n2130), .Z(n2127) );
  AND U3443 ( .A(b[23]), .B(a[34]), .Z(n2126) );
  XOR U3444 ( .A(n2131), .B(n2132), .Z(n1792) );
  AND U3445 ( .A(n2133), .B(n2134), .Z(n2131) );
  XNOR U3446 ( .A(n2135), .B(n1797), .Z(n1799) );
  XOR U3447 ( .A(n2136), .B(n2137), .Z(n1797) );
  ANDN U3448 ( .B(n2138), .A(n2139), .Z(n2136) );
  AND U3449 ( .A(b[22]), .B(a[35]), .Z(n2135) );
  XOR U3450 ( .A(n2140), .B(n1802), .Z(n1804) );
  XOR U3451 ( .A(n2141), .B(n2142), .Z(n1802) );
  ANDN U3452 ( .B(n2143), .A(n2144), .Z(n2141) );
  AND U3453 ( .A(b[20]), .B(a[37]), .Z(n2140) );
  XNOR U3454 ( .A(n2145), .B(n1807), .Z(n1809) );
  XOR U3455 ( .A(n2146), .B(n2147), .Z(n1807) );
  ANDN U3456 ( .B(n2148), .A(n2149), .Z(n2146) );
  AND U3457 ( .A(b[19]), .B(a[38]), .Z(n2145) );
  XNOR U3458 ( .A(n2150), .B(n1812), .Z(n1814) );
  XOR U3459 ( .A(n2151), .B(n2152), .Z(n1812) );
  ANDN U3460 ( .B(n2153), .A(n2154), .Z(n2151) );
  AND U3461 ( .A(b[18]), .B(a[39]), .Z(n2150) );
  XNOR U3462 ( .A(n2155), .B(n1817), .Z(n1819) );
  XOR U3463 ( .A(n2156), .B(n2157), .Z(n1817) );
  ANDN U3464 ( .B(n2158), .A(n2159), .Z(n2156) );
  AND U3465 ( .A(b[17]), .B(a[40]), .Z(n2155) );
  IV U3466 ( .A(n1824), .Z(n1917) );
  XNOR U3467 ( .A(n2160), .B(n1822), .Z(n1824) );
  XOR U3468 ( .A(n2161), .B(n2162), .Z(n1822) );
  ANDN U3469 ( .B(n2163), .A(n2164), .Z(n2161) );
  AND U3470 ( .A(b[16]), .B(a[41]), .Z(n2160) );
  XNOR U3471 ( .A(n2165), .B(n1827), .Z(n1829) );
  XOR U3472 ( .A(n2166), .B(n2167), .Z(n1827) );
  ANDN U3473 ( .B(n2168), .A(n2169), .Z(n2166) );
  AND U3474 ( .A(b[15]), .B(a[42]), .Z(n2165) );
  XNOR U3475 ( .A(n2170), .B(n1832), .Z(n1834) );
  XOR U3476 ( .A(n2171), .B(n2172), .Z(n1832) );
  ANDN U3477 ( .B(n2173), .A(n2174), .Z(n2171) );
  AND U3478 ( .A(b[14]), .B(a[43]), .Z(n2170) );
  XNOR U3479 ( .A(n2175), .B(n1837), .Z(n1839) );
  XOR U3480 ( .A(n2176), .B(n2177), .Z(n1837) );
  ANDN U3481 ( .B(n2178), .A(n2179), .Z(n2176) );
  AND U3482 ( .A(b[13]), .B(a[44]), .Z(n2175) );
  XNOR U3483 ( .A(n2180), .B(n1842), .Z(n1844) );
  XOR U3484 ( .A(n2181), .B(n2182), .Z(n1842) );
  ANDN U3485 ( .B(n2183), .A(n2184), .Z(n2181) );
  AND U3486 ( .A(b[12]), .B(a[45]), .Z(n2180) );
  XNOR U3487 ( .A(n2185), .B(n1847), .Z(n1849) );
  XOR U3488 ( .A(n2186), .B(n2187), .Z(n1847) );
  ANDN U3489 ( .B(n2188), .A(n2189), .Z(n2186) );
  AND U3490 ( .A(b[11]), .B(a[46]), .Z(n2185) );
  XNOR U3491 ( .A(n2190), .B(n1852), .Z(n1854) );
  XOR U3492 ( .A(n2191), .B(n2192), .Z(n1852) );
  ANDN U3493 ( .B(n2193), .A(n2194), .Z(n2191) );
  AND U3494 ( .A(b[10]), .B(a[47]), .Z(n2190) );
  XNOR U3495 ( .A(n2195), .B(n1857), .Z(n1859) );
  XOR U3496 ( .A(n2196), .B(n2197), .Z(n1857) );
  ANDN U3497 ( .B(n2198), .A(n2199), .Z(n2196) );
  AND U3498 ( .A(b[9]), .B(a[48]), .Z(n2195) );
  XNOR U3499 ( .A(n2200), .B(n1862), .Z(n1864) );
  XOR U3500 ( .A(n2201), .B(n2202), .Z(n1862) );
  ANDN U3501 ( .B(n2203), .A(n2204), .Z(n2201) );
  AND U3502 ( .A(b[8]), .B(a[49]), .Z(n2200) );
  XNOR U3503 ( .A(n2205), .B(n1867), .Z(n1869) );
  XOR U3504 ( .A(n2206), .B(n2207), .Z(n1867) );
  ANDN U3505 ( .B(n2208), .A(n2209), .Z(n2206) );
  AND U3506 ( .A(b[7]), .B(a[50]), .Z(n2205) );
  XNOR U3507 ( .A(n2210), .B(n1872), .Z(n1874) );
  XOR U3508 ( .A(n2211), .B(n2212), .Z(n1872) );
  ANDN U3509 ( .B(n2213), .A(n2214), .Z(n2211) );
  AND U3510 ( .A(b[6]), .B(a[51]), .Z(n2210) );
  XNOR U3511 ( .A(n2215), .B(n1877), .Z(n1879) );
  XOR U3512 ( .A(n2216), .B(n2217), .Z(n1877) );
  ANDN U3513 ( .B(n2218), .A(n2219), .Z(n2216) );
  AND U3514 ( .A(b[5]), .B(a[52]), .Z(n2215) );
  XNOR U3515 ( .A(n2220), .B(n1882), .Z(n1884) );
  XOR U3516 ( .A(n2221), .B(n2222), .Z(n1882) );
  ANDN U3517 ( .B(n2223), .A(n2224), .Z(n2221) );
  AND U3518 ( .A(b[4]), .B(a[53]), .Z(n2220) );
  XNOR U3519 ( .A(n2225), .B(n2226), .Z(n1896) );
  NANDN U3520 ( .A(n2227), .B(n2228), .Z(n2226) );
  XNOR U3521 ( .A(n2229), .B(n1887), .Z(n1889) );
  XNOR U3522 ( .A(n2230), .B(n2231), .Z(n1887) );
  AND U3523 ( .A(n2232), .B(n2233), .Z(n2230) );
  AND U3524 ( .A(b[3]), .B(a[54]), .Z(n2229) );
  NAND U3525 ( .A(a[57]), .B(b[0]), .Z(n1562) );
  XNOR U3526 ( .A(n1902), .B(n1903), .Z(c[56]) );
  XNOR U3527 ( .A(n2227), .B(n2228), .Z(n1903) );
  XOR U3528 ( .A(n2225), .B(n2234), .Z(n2228) );
  NAND U3529 ( .A(b[1]), .B(a[55]), .Z(n2234) );
  XOR U3530 ( .A(n2232), .B(n2235), .Z(n2227) );
  XOR U3531 ( .A(n2225), .B(n2233), .Z(n2235) );
  XNOR U3532 ( .A(n2236), .B(n2231), .Z(n2233) );
  AND U3533 ( .A(b[2]), .B(a[54]), .Z(n2236) );
  NANDN U3534 ( .A(n2237), .B(n2238), .Z(n2225) );
  XOR U3535 ( .A(n2231), .B(n2223), .Z(n2239) );
  XNOR U3536 ( .A(n2222), .B(n2218), .Z(n2240) );
  XNOR U3537 ( .A(n2217), .B(n2213), .Z(n2241) );
  XNOR U3538 ( .A(n2212), .B(n2208), .Z(n2242) );
  XNOR U3539 ( .A(n2207), .B(n2203), .Z(n2243) );
  XNOR U3540 ( .A(n2202), .B(n2198), .Z(n2244) );
  XNOR U3541 ( .A(n2197), .B(n2193), .Z(n2245) );
  XNOR U3542 ( .A(n2192), .B(n2188), .Z(n2246) );
  XNOR U3543 ( .A(n2187), .B(n2183), .Z(n2247) );
  XNOR U3544 ( .A(n2182), .B(n2178), .Z(n2248) );
  XNOR U3545 ( .A(n2177), .B(n2173), .Z(n2249) );
  XNOR U3546 ( .A(n2172), .B(n2168), .Z(n2250) );
  XNOR U3547 ( .A(n2167), .B(n2163), .Z(n2251) );
  XNOR U3548 ( .A(n2162), .B(n2158), .Z(n2252) );
  XNOR U3549 ( .A(n2157), .B(n2153), .Z(n2253) );
  XNOR U3550 ( .A(n2152), .B(n2148), .Z(n2254) );
  XNOR U3551 ( .A(n2147), .B(n2143), .Z(n2255) );
  XNOR U3552 ( .A(n2134), .B(n2133), .Z(n2256) );
  XOR U3553 ( .A(n2257), .B(n2132), .Z(n2133) );
  AND U3554 ( .A(b[20]), .B(a[36]), .Z(n2257) );
  XNOR U3555 ( .A(n2132), .B(n2138), .Z(n2258) );
  XNOR U3556 ( .A(n2137), .B(n2129), .Z(n2259) );
  XNOR U3557 ( .A(n2128), .B(n2124), .Z(n2260) );
  XNOR U3558 ( .A(n2123), .B(n2119), .Z(n2261) );
  XNOR U3559 ( .A(n2118), .B(n2114), .Z(n2262) );
  XNOR U3560 ( .A(n2105), .B(n2104), .Z(n2263) );
  XOR U3561 ( .A(n2264), .B(n2103), .Z(n2104) );
  AND U3562 ( .A(b[26]), .B(a[30]), .Z(n2264) );
  XNOR U3563 ( .A(n2103), .B(n2109), .Z(n2265) );
  XNOR U3564 ( .A(n2108), .B(n2100), .Z(n2266) );
  XNOR U3565 ( .A(n2099), .B(n2095), .Z(n2267) );
  XNOR U3566 ( .A(n2094), .B(n2090), .Z(n2268) );
  XNOR U3567 ( .A(n2089), .B(n2085), .Z(n2269) );
  XNOR U3568 ( .A(n2076), .B(n2075), .Z(n2270) );
  XOR U3569 ( .A(n2271), .B(n2074), .Z(n2075) );
  AND U3570 ( .A(b[32]), .B(a[24]), .Z(n2271) );
  XNOR U3571 ( .A(n2074), .B(n2080), .Z(n2272) );
  XNOR U3572 ( .A(n2079), .B(n2071), .Z(n2273) );
  XNOR U3573 ( .A(n2070), .B(n2066), .Z(n2274) );
  XNOR U3574 ( .A(n2065), .B(n2061), .Z(n2275) );
  XNOR U3575 ( .A(n2060), .B(n2056), .Z(n2276) );
  XNOR U3576 ( .A(n2047), .B(n2046), .Z(n2277) );
  XOR U3577 ( .A(n2278), .B(n2045), .Z(n2046) );
  AND U3578 ( .A(b[38]), .B(a[18]), .Z(n2278) );
  XNOR U3579 ( .A(n2045), .B(n2051), .Z(n2279) );
  XNOR U3580 ( .A(n2050), .B(n2042), .Z(n2280) );
  XNOR U3581 ( .A(n2041), .B(n2037), .Z(n2281) );
  XNOR U3582 ( .A(n2036), .B(n2032), .Z(n2282) );
  XNOR U3583 ( .A(n2031), .B(n2027), .Z(n2283) );
  XNOR U3584 ( .A(n2018), .B(n2017), .Z(n2284) );
  XOR U3585 ( .A(n2285), .B(n2016), .Z(n2017) );
  AND U3586 ( .A(b[44]), .B(a[12]), .Z(n2285) );
  XNOR U3587 ( .A(n2016), .B(n2022), .Z(n2286) );
  XNOR U3588 ( .A(n2021), .B(n2013), .Z(n2287) );
  XNOR U3589 ( .A(n2012), .B(n2008), .Z(n2288) );
  XNOR U3590 ( .A(n2007), .B(n2003), .Z(n2289) );
  XNOR U3591 ( .A(n2002), .B(n1998), .Z(n2290) );
  XNOR U3592 ( .A(n1989), .B(n1988), .Z(n2291) );
  XOR U3593 ( .A(n2292), .B(n1987), .Z(n1988) );
  AND U3594 ( .A(a[6]), .B(b[50]), .Z(n2292) );
  XNOR U3595 ( .A(n1987), .B(n1993), .Z(n2293) );
  XNOR U3596 ( .A(n1992), .B(n1984), .Z(n2294) );
  XNOR U3597 ( .A(n1983), .B(n1979), .Z(n2295) );
  XNOR U3598 ( .A(n1978), .B(n1974), .Z(n2296) );
  XNOR U3599 ( .A(n1973), .B(n1969), .Z(n2297) );
  XOR U3600 ( .A(n2298), .B(n1968), .Z(n1969) );
  AND U3601 ( .A(a[0]), .B(b[56]), .Z(n2298) );
  XNOR U3602 ( .A(n2299), .B(n1968), .Z(n1970) );
  XNOR U3603 ( .A(n2300), .B(n2301), .Z(n1968) );
  ANDN U3604 ( .B(n2302), .A(n2303), .Z(n2300) );
  AND U3605 ( .A(a[1]), .B(b[55]), .Z(n2299) );
  XNOR U3606 ( .A(n2304), .B(n1973), .Z(n1975) );
  XOR U3607 ( .A(n2305), .B(n2306), .Z(n1973) );
  ANDN U3608 ( .B(n2307), .A(n2308), .Z(n2305) );
  AND U3609 ( .A(a[2]), .B(b[54]), .Z(n2304) );
  XNOR U3610 ( .A(n2309), .B(n1978), .Z(n1980) );
  XOR U3611 ( .A(n2310), .B(n2311), .Z(n1978) );
  ANDN U3612 ( .B(n2312), .A(n2313), .Z(n2310) );
  AND U3613 ( .A(a[3]), .B(b[53]), .Z(n2309) );
  XNOR U3614 ( .A(n2314), .B(n1983), .Z(n1985) );
  XOR U3615 ( .A(n2315), .B(n2316), .Z(n1983) );
  ANDN U3616 ( .B(n2317), .A(n2318), .Z(n2315) );
  AND U3617 ( .A(a[4]), .B(b[52]), .Z(n2314) );
  XOR U3618 ( .A(n2319), .B(n2320), .Z(n1987) );
  AND U3619 ( .A(n2321), .B(n2322), .Z(n2319) );
  XNOR U3620 ( .A(n2323), .B(n1992), .Z(n1994) );
  XOR U3621 ( .A(n2324), .B(n2325), .Z(n1992) );
  ANDN U3622 ( .B(n2326), .A(n2327), .Z(n2324) );
  AND U3623 ( .A(a[5]), .B(b[51]), .Z(n2323) );
  XOR U3624 ( .A(n2328), .B(n1997), .Z(n1999) );
  XOR U3625 ( .A(n2329), .B(n2330), .Z(n1997) );
  ANDN U3626 ( .B(n2331), .A(n2332), .Z(n2329) );
  AND U3627 ( .A(a[7]), .B(b[49]), .Z(n2328) );
  XNOR U3628 ( .A(n2333), .B(n2002), .Z(n2004) );
  XOR U3629 ( .A(n2334), .B(n2335), .Z(n2002) );
  ANDN U3630 ( .B(n2336), .A(n2337), .Z(n2334) );
  AND U3631 ( .A(a[8]), .B(b[48]), .Z(n2333) );
  XNOR U3632 ( .A(n2338), .B(n2007), .Z(n2009) );
  XOR U3633 ( .A(n2339), .B(n2340), .Z(n2007) );
  ANDN U3634 ( .B(n2341), .A(n2342), .Z(n2339) );
  AND U3635 ( .A(a[9]), .B(b[47]), .Z(n2338) );
  XNOR U3636 ( .A(n2343), .B(n2012), .Z(n2014) );
  XOR U3637 ( .A(n2344), .B(n2345), .Z(n2012) );
  ANDN U3638 ( .B(n2346), .A(n2347), .Z(n2344) );
  AND U3639 ( .A(b[46]), .B(a[10]), .Z(n2343) );
  XOR U3640 ( .A(n2348), .B(n2349), .Z(n2016) );
  AND U3641 ( .A(n2350), .B(n2351), .Z(n2348) );
  XNOR U3642 ( .A(n2352), .B(n2021), .Z(n2023) );
  XOR U3643 ( .A(n2353), .B(n2354), .Z(n2021) );
  ANDN U3644 ( .B(n2355), .A(n2356), .Z(n2353) );
  AND U3645 ( .A(a[11]), .B(b[45]), .Z(n2352) );
  XOR U3646 ( .A(n2357), .B(n2026), .Z(n2028) );
  XOR U3647 ( .A(n2358), .B(n2359), .Z(n2026) );
  ANDN U3648 ( .B(n2360), .A(n2361), .Z(n2358) );
  AND U3649 ( .A(b[43]), .B(a[13]), .Z(n2357) );
  XNOR U3650 ( .A(n2362), .B(n2031), .Z(n2033) );
  XOR U3651 ( .A(n2363), .B(n2364), .Z(n2031) );
  ANDN U3652 ( .B(n2365), .A(n2366), .Z(n2363) );
  AND U3653 ( .A(b[42]), .B(a[14]), .Z(n2362) );
  XNOR U3654 ( .A(n2367), .B(n2036), .Z(n2038) );
  XOR U3655 ( .A(n2368), .B(n2369), .Z(n2036) );
  ANDN U3656 ( .B(n2370), .A(n2371), .Z(n2368) );
  AND U3657 ( .A(b[41]), .B(a[15]), .Z(n2367) );
  XNOR U3658 ( .A(n2372), .B(n2041), .Z(n2043) );
  XOR U3659 ( .A(n2373), .B(n2374), .Z(n2041) );
  ANDN U3660 ( .B(n2375), .A(n2376), .Z(n2373) );
  AND U3661 ( .A(b[40]), .B(a[16]), .Z(n2372) );
  XOR U3662 ( .A(n2377), .B(n2378), .Z(n2045) );
  AND U3663 ( .A(n2379), .B(n2380), .Z(n2377) );
  XNOR U3664 ( .A(n2381), .B(n2050), .Z(n2052) );
  XOR U3665 ( .A(n2382), .B(n2383), .Z(n2050) );
  ANDN U3666 ( .B(n2384), .A(n2385), .Z(n2382) );
  AND U3667 ( .A(a[17]), .B(b[39]), .Z(n2381) );
  XOR U3668 ( .A(n2386), .B(n2055), .Z(n2057) );
  XOR U3669 ( .A(n2387), .B(n2388), .Z(n2055) );
  ANDN U3670 ( .B(n2389), .A(n2390), .Z(n2387) );
  AND U3671 ( .A(b[37]), .B(a[19]), .Z(n2386) );
  XNOR U3672 ( .A(n2391), .B(n2060), .Z(n2062) );
  XOR U3673 ( .A(n2392), .B(n2393), .Z(n2060) );
  ANDN U3674 ( .B(n2394), .A(n2395), .Z(n2392) );
  AND U3675 ( .A(b[36]), .B(a[20]), .Z(n2391) );
  XNOR U3676 ( .A(n2396), .B(n2065), .Z(n2067) );
  XOR U3677 ( .A(n2397), .B(n2398), .Z(n2065) );
  ANDN U3678 ( .B(n2399), .A(n2400), .Z(n2397) );
  AND U3679 ( .A(b[35]), .B(a[21]), .Z(n2396) );
  XNOR U3680 ( .A(n2401), .B(n2070), .Z(n2072) );
  XOR U3681 ( .A(n2402), .B(n2403), .Z(n2070) );
  ANDN U3682 ( .B(n2404), .A(n2405), .Z(n2402) );
  AND U3683 ( .A(b[34]), .B(a[22]), .Z(n2401) );
  XOR U3684 ( .A(n2406), .B(n2407), .Z(n2074) );
  AND U3685 ( .A(n2408), .B(n2409), .Z(n2406) );
  XNOR U3686 ( .A(n2410), .B(n2079), .Z(n2081) );
  XOR U3687 ( .A(n2411), .B(n2412), .Z(n2079) );
  ANDN U3688 ( .B(n2413), .A(n2414), .Z(n2411) );
  AND U3689 ( .A(a[23]), .B(b[33]), .Z(n2410) );
  XOR U3690 ( .A(n2415), .B(n2084), .Z(n2086) );
  XOR U3691 ( .A(n2416), .B(n2417), .Z(n2084) );
  ANDN U3692 ( .B(n2418), .A(n2419), .Z(n2416) );
  AND U3693 ( .A(b[31]), .B(a[25]), .Z(n2415) );
  XNOR U3694 ( .A(n2420), .B(n2089), .Z(n2091) );
  XOR U3695 ( .A(n2421), .B(n2422), .Z(n2089) );
  ANDN U3696 ( .B(n2423), .A(n2424), .Z(n2421) );
  AND U3697 ( .A(b[30]), .B(a[26]), .Z(n2420) );
  XNOR U3698 ( .A(n2425), .B(n2094), .Z(n2096) );
  XOR U3699 ( .A(n2426), .B(n2427), .Z(n2094) );
  ANDN U3700 ( .B(n2428), .A(n2429), .Z(n2426) );
  AND U3701 ( .A(b[29]), .B(a[27]), .Z(n2425) );
  XNOR U3702 ( .A(n2430), .B(n2099), .Z(n2101) );
  XOR U3703 ( .A(n2431), .B(n2432), .Z(n2099) );
  ANDN U3704 ( .B(n2433), .A(n2434), .Z(n2431) );
  AND U3705 ( .A(b[28]), .B(a[28]), .Z(n2430) );
  XOR U3706 ( .A(n2435), .B(n2436), .Z(n2103) );
  AND U3707 ( .A(n2437), .B(n2438), .Z(n2435) );
  XNOR U3708 ( .A(n2439), .B(n2108), .Z(n2110) );
  XOR U3709 ( .A(n2440), .B(n2441), .Z(n2108) );
  ANDN U3710 ( .B(n2442), .A(n2443), .Z(n2440) );
  AND U3711 ( .A(a[29]), .B(b[27]), .Z(n2439) );
  XOR U3712 ( .A(n2444), .B(n2113), .Z(n2115) );
  XOR U3713 ( .A(n2445), .B(n2446), .Z(n2113) );
  ANDN U3714 ( .B(n2447), .A(n2448), .Z(n2445) );
  AND U3715 ( .A(b[25]), .B(a[31]), .Z(n2444) );
  XNOR U3716 ( .A(n2449), .B(n2118), .Z(n2120) );
  XOR U3717 ( .A(n2450), .B(n2451), .Z(n2118) );
  ANDN U3718 ( .B(n2452), .A(n2453), .Z(n2450) );
  AND U3719 ( .A(b[24]), .B(a[32]), .Z(n2449) );
  XNOR U3720 ( .A(n2454), .B(n2123), .Z(n2125) );
  XOR U3721 ( .A(n2455), .B(n2456), .Z(n2123) );
  ANDN U3722 ( .B(n2457), .A(n2458), .Z(n2455) );
  AND U3723 ( .A(b[23]), .B(a[33]), .Z(n2454) );
  XNOR U3724 ( .A(n2459), .B(n2128), .Z(n2130) );
  XOR U3725 ( .A(n2460), .B(n2461), .Z(n2128) );
  ANDN U3726 ( .B(n2462), .A(n2463), .Z(n2460) );
  AND U3727 ( .A(b[22]), .B(a[34]), .Z(n2459) );
  XOR U3728 ( .A(n2464), .B(n2465), .Z(n2132) );
  AND U3729 ( .A(n2466), .B(n2467), .Z(n2464) );
  XNOR U3730 ( .A(n2468), .B(n2137), .Z(n2139) );
  XOR U3731 ( .A(n2469), .B(n2470), .Z(n2137) );
  ANDN U3732 ( .B(n2471), .A(n2472), .Z(n2469) );
  AND U3733 ( .A(a[35]), .B(b[21]), .Z(n2468) );
  XOR U3734 ( .A(n2473), .B(n2142), .Z(n2144) );
  XOR U3735 ( .A(n2474), .B(n2475), .Z(n2142) );
  ANDN U3736 ( .B(n2476), .A(n2477), .Z(n2474) );
  AND U3737 ( .A(b[19]), .B(a[37]), .Z(n2473) );
  XNOR U3738 ( .A(n2478), .B(n2147), .Z(n2149) );
  XOR U3739 ( .A(n2479), .B(n2480), .Z(n2147) );
  ANDN U3740 ( .B(n2481), .A(n2482), .Z(n2479) );
  AND U3741 ( .A(b[18]), .B(a[38]), .Z(n2478) );
  XNOR U3742 ( .A(n2483), .B(n2152), .Z(n2154) );
  XOR U3743 ( .A(n2484), .B(n2485), .Z(n2152) );
  ANDN U3744 ( .B(n2486), .A(n2487), .Z(n2484) );
  AND U3745 ( .A(b[17]), .B(a[39]), .Z(n2483) );
  XNOR U3746 ( .A(n2488), .B(n2157), .Z(n2159) );
  XOR U3747 ( .A(n2489), .B(n2490), .Z(n2157) );
  ANDN U3748 ( .B(n2491), .A(n2492), .Z(n2489) );
  AND U3749 ( .A(b[16]), .B(a[40]), .Z(n2488) );
  XNOR U3750 ( .A(n2493), .B(n2162), .Z(n2164) );
  XOR U3751 ( .A(n2494), .B(n2495), .Z(n2162) );
  ANDN U3752 ( .B(n2496), .A(n2497), .Z(n2494) );
  AND U3753 ( .A(a[41]), .B(b[15]), .Z(n2493) );
  XNOR U3754 ( .A(n2498), .B(n2167), .Z(n2169) );
  XOR U3755 ( .A(n2499), .B(n2500), .Z(n2167) );
  ANDN U3756 ( .B(n2501), .A(n2502), .Z(n2499) );
  AND U3757 ( .A(b[14]), .B(a[42]), .Z(n2498) );
  XNOR U3758 ( .A(n2503), .B(n2172), .Z(n2174) );
  XOR U3759 ( .A(n2504), .B(n2505), .Z(n2172) );
  ANDN U3760 ( .B(n2506), .A(n2507), .Z(n2504) );
  AND U3761 ( .A(b[13]), .B(a[43]), .Z(n2503) );
  XNOR U3762 ( .A(n2508), .B(n2177), .Z(n2179) );
  XOR U3763 ( .A(n2509), .B(n2510), .Z(n2177) );
  ANDN U3764 ( .B(n2511), .A(n2512), .Z(n2509) );
  AND U3765 ( .A(b[12]), .B(a[44]), .Z(n2508) );
  XNOR U3766 ( .A(n2513), .B(n2182), .Z(n2184) );
  XOR U3767 ( .A(n2514), .B(n2515), .Z(n2182) );
  ANDN U3768 ( .B(n2516), .A(n2517), .Z(n2514) );
  AND U3769 ( .A(b[11]), .B(a[45]), .Z(n2513) );
  XNOR U3770 ( .A(n2518), .B(n2187), .Z(n2189) );
  XOR U3771 ( .A(n2519), .B(n2520), .Z(n2187) );
  ANDN U3772 ( .B(n2521), .A(n2522), .Z(n2519) );
  AND U3773 ( .A(b[10]), .B(a[46]), .Z(n2518) );
  XNOR U3774 ( .A(n2523), .B(n2192), .Z(n2194) );
  XOR U3775 ( .A(n2524), .B(n2525), .Z(n2192) );
  ANDN U3776 ( .B(n2526), .A(n2527), .Z(n2524) );
  AND U3777 ( .A(b[9]), .B(a[47]), .Z(n2523) );
  XNOR U3778 ( .A(n2528), .B(n2197), .Z(n2199) );
  XOR U3779 ( .A(n2529), .B(n2530), .Z(n2197) );
  ANDN U3780 ( .B(n2531), .A(n2532), .Z(n2529) );
  AND U3781 ( .A(b[8]), .B(a[48]), .Z(n2528) );
  XNOR U3782 ( .A(n2533), .B(n2202), .Z(n2204) );
  XOR U3783 ( .A(n2534), .B(n2535), .Z(n2202) );
  ANDN U3784 ( .B(n2536), .A(n2537), .Z(n2534) );
  AND U3785 ( .A(b[7]), .B(a[49]), .Z(n2533) );
  XNOR U3786 ( .A(n2538), .B(n2207), .Z(n2209) );
  XOR U3787 ( .A(n2539), .B(n2540), .Z(n2207) );
  ANDN U3788 ( .B(n2541), .A(n2542), .Z(n2539) );
  AND U3789 ( .A(b[6]), .B(a[50]), .Z(n2538) );
  XNOR U3790 ( .A(n2543), .B(n2212), .Z(n2214) );
  XOR U3791 ( .A(n2544), .B(n2545), .Z(n2212) );
  ANDN U3792 ( .B(n2546), .A(n2547), .Z(n2544) );
  AND U3793 ( .A(b[5]), .B(a[51]), .Z(n2543) );
  XNOR U3794 ( .A(n2548), .B(n2217), .Z(n2219) );
  XOR U3795 ( .A(n2549), .B(n2550), .Z(n2217) );
  ANDN U3796 ( .B(n2551), .A(n2552), .Z(n2549) );
  AND U3797 ( .A(b[4]), .B(a[52]), .Z(n2548) );
  XNOR U3798 ( .A(n2553), .B(n2554), .Z(n2231) );
  NANDN U3799 ( .A(n2555), .B(n2556), .Z(n2554) );
  XNOR U3800 ( .A(n2557), .B(n2222), .Z(n2224) );
  XNOR U3801 ( .A(n2558), .B(n2559), .Z(n2222) );
  NOR U3802 ( .A(n2560), .B(n2561), .Z(n2558) );
  AND U3803 ( .A(b[3]), .B(a[53]), .Z(n2557) );
  NAND U3804 ( .A(a[56]), .B(b[0]), .Z(n1902) );
  XNOR U3805 ( .A(n2237), .B(n2238), .Z(c[55]) );
  XOR U3806 ( .A(n2562), .B(n2563), .Z(n2555) );
  NAND U3807 ( .A(b[1]), .B(a[54]), .Z(n2563) );
  XOR U3808 ( .A(n2562), .B(n2561), .Z(n2564) );
  XOR U3809 ( .A(n2565), .B(n2559), .Z(n2561) );
  AND U3810 ( .A(b[2]), .B(a[53]), .Z(n2565) );
  IV U3811 ( .A(n2553), .Z(n2562) );
  NANDN U3812 ( .A(n2566), .B(n2567), .Z(n2553) );
  XOR U3813 ( .A(n2559), .B(n2551), .Z(n2568) );
  XNOR U3814 ( .A(n2550), .B(n2546), .Z(n2569) );
  XNOR U3815 ( .A(n2545), .B(n2541), .Z(n2570) );
  XNOR U3816 ( .A(n2540), .B(n2536), .Z(n2571) );
  XNOR U3817 ( .A(n2535), .B(n2531), .Z(n2572) );
  XNOR U3818 ( .A(n2530), .B(n2526), .Z(n2573) );
  XNOR U3819 ( .A(n2525), .B(n2521), .Z(n2574) );
  XNOR U3820 ( .A(n2520), .B(n2516), .Z(n2575) );
  XNOR U3821 ( .A(n2515), .B(n2511), .Z(n2576) );
  XNOR U3822 ( .A(n2510), .B(n2506), .Z(n2577) );
  XNOR U3823 ( .A(n2505), .B(n2501), .Z(n2578) );
  XNOR U3824 ( .A(n2500), .B(n2496), .Z(n2579) );
  XNOR U3825 ( .A(n2495), .B(n2491), .Z(n2580) );
  XNOR U3826 ( .A(n2490), .B(n2486), .Z(n2581) );
  XNOR U3827 ( .A(n2485), .B(n2481), .Z(n2582) );
  XNOR U3828 ( .A(n2480), .B(n2476), .Z(n2583) );
  XNOR U3829 ( .A(n2584), .B(n2585), .Z(n2476) );
  XNOR U3830 ( .A(n2467), .B(n2466), .Z(n2585) );
  XOR U3831 ( .A(n2586), .B(n2465), .Z(n2466) );
  AND U3832 ( .A(b[19]), .B(a[36]), .Z(n2586) );
  XNOR U3833 ( .A(n2465), .B(n2471), .Z(n2587) );
  XNOR U3834 ( .A(n2470), .B(n2462), .Z(n2588) );
  XNOR U3835 ( .A(n2461), .B(n2457), .Z(n2589) );
  XNOR U3836 ( .A(n2456), .B(n2452), .Z(n2590) );
  XNOR U3837 ( .A(n2451), .B(n2447), .Z(n2591) );
  XNOR U3838 ( .A(n2438), .B(n2437), .Z(n2592) );
  XOR U3839 ( .A(n2593), .B(n2436), .Z(n2437) );
  AND U3840 ( .A(b[25]), .B(a[30]), .Z(n2593) );
  XNOR U3841 ( .A(n2436), .B(n2442), .Z(n2594) );
  XNOR U3842 ( .A(n2441), .B(n2433), .Z(n2595) );
  XNOR U3843 ( .A(n2432), .B(n2428), .Z(n2596) );
  XNOR U3844 ( .A(n2427), .B(n2423), .Z(n2597) );
  XNOR U3845 ( .A(n2422), .B(n2418), .Z(n2598) );
  XNOR U3846 ( .A(n2409), .B(n2408), .Z(n2599) );
  XOR U3847 ( .A(n2600), .B(n2407), .Z(n2408) );
  AND U3848 ( .A(b[31]), .B(a[24]), .Z(n2600) );
  XNOR U3849 ( .A(n2407), .B(n2413), .Z(n2601) );
  XNOR U3850 ( .A(n2412), .B(n2404), .Z(n2602) );
  XNOR U3851 ( .A(n2403), .B(n2399), .Z(n2603) );
  XNOR U3852 ( .A(n2398), .B(n2394), .Z(n2604) );
  XNOR U3853 ( .A(n2393), .B(n2389), .Z(n2605) );
  XNOR U3854 ( .A(n2380), .B(n2379), .Z(n2606) );
  XOR U3855 ( .A(n2607), .B(n2378), .Z(n2379) );
  AND U3856 ( .A(b[37]), .B(a[18]), .Z(n2607) );
  XNOR U3857 ( .A(n2378), .B(n2384), .Z(n2608) );
  XNOR U3858 ( .A(n2383), .B(n2375), .Z(n2609) );
  XNOR U3859 ( .A(n2374), .B(n2370), .Z(n2610) );
  XNOR U3860 ( .A(n2369), .B(n2365), .Z(n2611) );
  XNOR U3861 ( .A(n2364), .B(n2360), .Z(n2612) );
  XNOR U3862 ( .A(n2351), .B(n2350), .Z(n2613) );
  XOR U3863 ( .A(n2614), .B(n2349), .Z(n2350) );
  AND U3864 ( .A(b[43]), .B(a[12]), .Z(n2614) );
  XNOR U3865 ( .A(n2349), .B(n2355), .Z(n2615) );
  XNOR U3866 ( .A(n2354), .B(n2346), .Z(n2616) );
  XNOR U3867 ( .A(n2345), .B(n2341), .Z(n2617) );
  XNOR U3868 ( .A(n2340), .B(n2336), .Z(n2618) );
  XNOR U3869 ( .A(n2335), .B(n2331), .Z(n2619) );
  XNOR U3870 ( .A(n2620), .B(n2621), .Z(n2331) );
  XNOR U3871 ( .A(n2322), .B(n2321), .Z(n2621) );
  XOR U3872 ( .A(n2622), .B(n2320), .Z(n2321) );
  AND U3873 ( .A(a[6]), .B(b[49]), .Z(n2622) );
  XNOR U3874 ( .A(n2320), .B(n2326), .Z(n2623) );
  XNOR U3875 ( .A(n2325), .B(n2317), .Z(n2624) );
  XNOR U3876 ( .A(n2316), .B(n2312), .Z(n2625) );
  XNOR U3877 ( .A(n2311), .B(n2307), .Z(n2626) );
  XNOR U3878 ( .A(n2306), .B(n2302), .Z(n2627) );
  XNOR U3879 ( .A(n2628), .B(n2301), .Z(n2302) );
  AND U3880 ( .A(a[0]), .B(b[55]), .Z(n2628) );
  XOR U3881 ( .A(n2629), .B(n2301), .Z(n2303) );
  XNOR U3882 ( .A(n2630), .B(n2631), .Z(n2301) );
  ANDN U3883 ( .B(n2632), .A(n2633), .Z(n2630) );
  AND U3884 ( .A(a[1]), .B(b[54]), .Z(n2629) );
  XNOR U3885 ( .A(n2634), .B(n2306), .Z(n2308) );
  XOR U3886 ( .A(n2635), .B(n2636), .Z(n2306) );
  ANDN U3887 ( .B(n2637), .A(n2638), .Z(n2635) );
  AND U3888 ( .A(a[2]), .B(b[53]), .Z(n2634) );
  XNOR U3889 ( .A(n2639), .B(n2311), .Z(n2313) );
  XOR U3890 ( .A(n2640), .B(n2641), .Z(n2311) );
  ANDN U3891 ( .B(n2642), .A(n2643), .Z(n2640) );
  AND U3892 ( .A(a[3]), .B(b[52]), .Z(n2639) );
  XNOR U3893 ( .A(n2644), .B(n2316), .Z(n2318) );
  XOR U3894 ( .A(n2645), .B(n2646), .Z(n2316) );
  ANDN U3895 ( .B(n2647), .A(n2648), .Z(n2645) );
  AND U3896 ( .A(a[4]), .B(b[51]), .Z(n2644) );
  XOR U3897 ( .A(n2649), .B(n2650), .Z(n2320) );
  AND U3898 ( .A(n2651), .B(n2652), .Z(n2649) );
  XNOR U3899 ( .A(n2653), .B(n2325), .Z(n2327) );
  XOR U3900 ( .A(n2654), .B(n2655), .Z(n2325) );
  ANDN U3901 ( .B(n2656), .A(n2657), .Z(n2654) );
  AND U3902 ( .A(a[5]), .B(b[50]), .Z(n2653) );
  IV U3903 ( .A(n2330), .Z(n2620) );
  XOR U3904 ( .A(n2658), .B(n2330), .Z(n2332) );
  XOR U3905 ( .A(n2659), .B(n2660), .Z(n2330) );
  ANDN U3906 ( .B(n2661), .A(n2662), .Z(n2659) );
  AND U3907 ( .A(a[7]), .B(b[48]), .Z(n2658) );
  XNOR U3908 ( .A(n2663), .B(n2335), .Z(n2337) );
  XOR U3909 ( .A(n2664), .B(n2665), .Z(n2335) );
  ANDN U3910 ( .B(n2666), .A(n2667), .Z(n2664) );
  AND U3911 ( .A(a[8]), .B(b[47]), .Z(n2663) );
  XNOR U3912 ( .A(n2668), .B(n2340), .Z(n2342) );
  XOR U3913 ( .A(n2669), .B(n2670), .Z(n2340) );
  ANDN U3914 ( .B(n2671), .A(n2672), .Z(n2669) );
  AND U3915 ( .A(a[9]), .B(b[46]), .Z(n2668) );
  XNOR U3916 ( .A(n2673), .B(n2345), .Z(n2347) );
  XOR U3917 ( .A(n2674), .B(n2675), .Z(n2345) );
  ANDN U3918 ( .B(n2676), .A(n2677), .Z(n2674) );
  AND U3919 ( .A(a[10]), .B(b[45]), .Z(n2673) );
  XOR U3920 ( .A(n2678), .B(n2679), .Z(n2349) );
  AND U3921 ( .A(n2680), .B(n2681), .Z(n2678) );
  XNOR U3922 ( .A(n2682), .B(n2354), .Z(n2356) );
  XOR U3923 ( .A(n2683), .B(n2684), .Z(n2354) );
  ANDN U3924 ( .B(n2685), .A(n2686), .Z(n2683) );
  AND U3925 ( .A(b[44]), .B(a[11]), .Z(n2682) );
  XOR U3926 ( .A(n2687), .B(n2359), .Z(n2361) );
  XOR U3927 ( .A(n2688), .B(n2689), .Z(n2359) );
  ANDN U3928 ( .B(n2690), .A(n2691), .Z(n2688) );
  AND U3929 ( .A(b[42]), .B(a[13]), .Z(n2687) );
  XNOR U3930 ( .A(n2692), .B(n2364), .Z(n2366) );
  XOR U3931 ( .A(n2693), .B(n2694), .Z(n2364) );
  ANDN U3932 ( .B(n2695), .A(n2696), .Z(n2693) );
  AND U3933 ( .A(b[41]), .B(a[14]), .Z(n2692) );
  XNOR U3934 ( .A(n2697), .B(n2369), .Z(n2371) );
  XOR U3935 ( .A(n2698), .B(n2699), .Z(n2369) );
  ANDN U3936 ( .B(n2700), .A(n2701), .Z(n2698) );
  AND U3937 ( .A(b[40]), .B(a[15]), .Z(n2697) );
  XNOR U3938 ( .A(n2702), .B(n2374), .Z(n2376) );
  XOR U3939 ( .A(n2703), .B(n2704), .Z(n2374) );
  ANDN U3940 ( .B(n2705), .A(n2706), .Z(n2703) );
  AND U3941 ( .A(a[16]), .B(b[39]), .Z(n2702) );
  XOR U3942 ( .A(n2707), .B(n2708), .Z(n2378) );
  AND U3943 ( .A(n2709), .B(n2710), .Z(n2707) );
  XNOR U3944 ( .A(n2711), .B(n2383), .Z(n2385) );
  XOR U3945 ( .A(n2712), .B(n2713), .Z(n2383) );
  ANDN U3946 ( .B(n2714), .A(n2715), .Z(n2712) );
  AND U3947 ( .A(b[38]), .B(a[17]), .Z(n2711) );
  XOR U3948 ( .A(n2716), .B(n2388), .Z(n2390) );
  XOR U3949 ( .A(n2717), .B(n2718), .Z(n2388) );
  ANDN U3950 ( .B(n2719), .A(n2720), .Z(n2717) );
  AND U3951 ( .A(b[36]), .B(a[19]), .Z(n2716) );
  XNOR U3952 ( .A(n2721), .B(n2393), .Z(n2395) );
  XOR U3953 ( .A(n2722), .B(n2723), .Z(n2393) );
  ANDN U3954 ( .B(n2724), .A(n2725), .Z(n2722) );
  AND U3955 ( .A(b[35]), .B(a[20]), .Z(n2721) );
  XNOR U3956 ( .A(n2726), .B(n2398), .Z(n2400) );
  XOR U3957 ( .A(n2727), .B(n2728), .Z(n2398) );
  ANDN U3958 ( .B(n2729), .A(n2730), .Z(n2727) );
  AND U3959 ( .A(b[34]), .B(a[21]), .Z(n2726) );
  XNOR U3960 ( .A(n2731), .B(n2403), .Z(n2405) );
  XOR U3961 ( .A(n2732), .B(n2733), .Z(n2403) );
  ANDN U3962 ( .B(n2734), .A(n2735), .Z(n2732) );
  AND U3963 ( .A(a[22]), .B(b[33]), .Z(n2731) );
  XOR U3964 ( .A(n2736), .B(n2737), .Z(n2407) );
  AND U3965 ( .A(n2738), .B(n2739), .Z(n2736) );
  XNOR U3966 ( .A(n2740), .B(n2412), .Z(n2414) );
  XOR U3967 ( .A(n2741), .B(n2742), .Z(n2412) );
  ANDN U3968 ( .B(n2743), .A(n2744), .Z(n2741) );
  AND U3969 ( .A(b[32]), .B(a[23]), .Z(n2740) );
  XOR U3970 ( .A(n2745), .B(n2417), .Z(n2419) );
  XOR U3971 ( .A(n2746), .B(n2747), .Z(n2417) );
  ANDN U3972 ( .B(n2748), .A(n2749), .Z(n2746) );
  AND U3973 ( .A(b[30]), .B(a[25]), .Z(n2745) );
  XNOR U3974 ( .A(n2750), .B(n2422), .Z(n2424) );
  XOR U3975 ( .A(n2751), .B(n2752), .Z(n2422) );
  ANDN U3976 ( .B(n2753), .A(n2754), .Z(n2751) );
  AND U3977 ( .A(b[29]), .B(a[26]), .Z(n2750) );
  XNOR U3978 ( .A(n2755), .B(n2427), .Z(n2429) );
  XOR U3979 ( .A(n2756), .B(n2757), .Z(n2427) );
  ANDN U3980 ( .B(n2758), .A(n2759), .Z(n2756) );
  AND U3981 ( .A(b[28]), .B(a[27]), .Z(n2755) );
  XNOR U3982 ( .A(n2760), .B(n2432), .Z(n2434) );
  XOR U3983 ( .A(n2761), .B(n2762), .Z(n2432) );
  ANDN U3984 ( .B(n2763), .A(n2764), .Z(n2761) );
  AND U3985 ( .A(a[28]), .B(b[27]), .Z(n2760) );
  XOR U3986 ( .A(n2765), .B(n2766), .Z(n2436) );
  AND U3987 ( .A(n2767), .B(n2768), .Z(n2765) );
  XNOR U3988 ( .A(n2769), .B(n2441), .Z(n2443) );
  XOR U3989 ( .A(n2770), .B(n2771), .Z(n2441) );
  ANDN U3990 ( .B(n2772), .A(n2773), .Z(n2770) );
  AND U3991 ( .A(b[26]), .B(a[29]), .Z(n2769) );
  XOR U3992 ( .A(n2774), .B(n2446), .Z(n2448) );
  XOR U3993 ( .A(n2775), .B(n2776), .Z(n2446) );
  ANDN U3994 ( .B(n2777), .A(n2778), .Z(n2775) );
  AND U3995 ( .A(b[24]), .B(a[31]), .Z(n2774) );
  XNOR U3996 ( .A(n2779), .B(n2451), .Z(n2453) );
  XOR U3997 ( .A(n2780), .B(n2781), .Z(n2451) );
  ANDN U3998 ( .B(n2782), .A(n2783), .Z(n2780) );
  AND U3999 ( .A(b[23]), .B(a[32]), .Z(n2779) );
  XNOR U4000 ( .A(n2784), .B(n2456), .Z(n2458) );
  XOR U4001 ( .A(n2785), .B(n2786), .Z(n2456) );
  ANDN U4002 ( .B(n2787), .A(n2788), .Z(n2785) );
  AND U4003 ( .A(b[22]), .B(a[33]), .Z(n2784) );
  XNOR U4004 ( .A(n2789), .B(n2461), .Z(n2463) );
  XOR U4005 ( .A(n2790), .B(n2791), .Z(n2461) );
  ANDN U4006 ( .B(n2792), .A(n2793), .Z(n2790) );
  AND U4007 ( .A(a[34]), .B(b[21]), .Z(n2789) );
  XOR U4008 ( .A(n2794), .B(n2795), .Z(n2465) );
  AND U4009 ( .A(n2796), .B(n2797), .Z(n2794) );
  XNOR U4010 ( .A(n2798), .B(n2470), .Z(n2472) );
  XOR U4011 ( .A(n2799), .B(n2800), .Z(n2470) );
  ANDN U4012 ( .B(n2801), .A(n2802), .Z(n2799) );
  AND U4013 ( .A(b[20]), .B(a[35]), .Z(n2798) );
  IV U4014 ( .A(n2475), .Z(n2584) );
  XOR U4015 ( .A(n2803), .B(n2475), .Z(n2477) );
  XOR U4016 ( .A(n2804), .B(n2805), .Z(n2475) );
  ANDN U4017 ( .B(n2806), .A(n2807), .Z(n2804) );
  AND U4018 ( .A(b[18]), .B(a[37]), .Z(n2803) );
  XNOR U4019 ( .A(n2808), .B(n2480), .Z(n2482) );
  XOR U4020 ( .A(n2809), .B(n2810), .Z(n2480) );
  ANDN U4021 ( .B(n2811), .A(n2812), .Z(n2809) );
  AND U4022 ( .A(b[17]), .B(a[38]), .Z(n2808) );
  XNOR U4023 ( .A(n2813), .B(n2485), .Z(n2487) );
  XOR U4024 ( .A(n2814), .B(n2815), .Z(n2485) );
  ANDN U4025 ( .B(n2816), .A(n2817), .Z(n2814) );
  AND U4026 ( .A(b[16]), .B(a[39]), .Z(n2813) );
  XNOR U4027 ( .A(n2818), .B(n2490), .Z(n2492) );
  XOR U4028 ( .A(n2819), .B(n2820), .Z(n2490) );
  ANDN U4029 ( .B(n2821), .A(n2822), .Z(n2819) );
  AND U4030 ( .A(a[40]), .B(b[15]), .Z(n2818) );
  XNOR U4031 ( .A(n2823), .B(n2495), .Z(n2497) );
  XOR U4032 ( .A(n2824), .B(n2825), .Z(n2495) );
  ANDN U4033 ( .B(n2826), .A(n2827), .Z(n2824) );
  AND U4034 ( .A(b[14]), .B(a[41]), .Z(n2823) );
  XNOR U4035 ( .A(n2828), .B(n2500), .Z(n2502) );
  XOR U4036 ( .A(n2829), .B(n2830), .Z(n2500) );
  ANDN U4037 ( .B(n2831), .A(n2832), .Z(n2829) );
  AND U4038 ( .A(b[13]), .B(a[42]), .Z(n2828) );
  XNOR U4039 ( .A(n2833), .B(n2505), .Z(n2507) );
  XOR U4040 ( .A(n2834), .B(n2835), .Z(n2505) );
  ANDN U4041 ( .B(n2836), .A(n2837), .Z(n2834) );
  AND U4042 ( .A(b[12]), .B(a[43]), .Z(n2833) );
  XNOR U4043 ( .A(n2838), .B(n2510), .Z(n2512) );
  XOR U4044 ( .A(n2839), .B(n2840), .Z(n2510) );
  ANDN U4045 ( .B(n2841), .A(n2842), .Z(n2839) );
  AND U4046 ( .A(b[11]), .B(a[44]), .Z(n2838) );
  XNOR U4047 ( .A(n2843), .B(n2515), .Z(n2517) );
  XOR U4048 ( .A(n2844), .B(n2845), .Z(n2515) );
  ANDN U4049 ( .B(n2846), .A(n2847), .Z(n2844) );
  AND U4050 ( .A(b[10]), .B(a[45]), .Z(n2843) );
  XNOR U4051 ( .A(n2848), .B(n2520), .Z(n2522) );
  XOR U4052 ( .A(n2849), .B(n2850), .Z(n2520) );
  ANDN U4053 ( .B(n2851), .A(n2852), .Z(n2849) );
  AND U4054 ( .A(b[9]), .B(a[46]), .Z(n2848) );
  XNOR U4055 ( .A(n2853), .B(n2525), .Z(n2527) );
  XOR U4056 ( .A(n2854), .B(n2855), .Z(n2525) );
  ANDN U4057 ( .B(n2856), .A(n2857), .Z(n2854) );
  AND U4058 ( .A(b[8]), .B(a[47]), .Z(n2853) );
  XNOR U4059 ( .A(n2858), .B(n2530), .Z(n2532) );
  XOR U4060 ( .A(n2859), .B(n2860), .Z(n2530) );
  ANDN U4061 ( .B(n2861), .A(n2862), .Z(n2859) );
  AND U4062 ( .A(b[7]), .B(a[48]), .Z(n2858) );
  XNOR U4063 ( .A(n2863), .B(n2535), .Z(n2537) );
  XOR U4064 ( .A(n2864), .B(n2865), .Z(n2535) );
  ANDN U4065 ( .B(n2866), .A(n2867), .Z(n2864) );
  AND U4066 ( .A(b[6]), .B(a[49]), .Z(n2863) );
  XNOR U4067 ( .A(n2868), .B(n2540), .Z(n2542) );
  XOR U4068 ( .A(n2869), .B(n2870), .Z(n2540) );
  ANDN U4069 ( .B(n2871), .A(n2872), .Z(n2869) );
  AND U4070 ( .A(b[5]), .B(a[50]), .Z(n2868) );
  XNOR U4071 ( .A(n2873), .B(n2545), .Z(n2547) );
  XOR U4072 ( .A(n2874), .B(n2875), .Z(n2545) );
  ANDN U4073 ( .B(n2876), .A(n2877), .Z(n2874) );
  AND U4074 ( .A(b[4]), .B(a[51]), .Z(n2873) );
  XOR U4075 ( .A(n2878), .B(n2879), .Z(n2559) );
  NANDN U4076 ( .A(n2880), .B(n2881), .Z(n2879) );
  XNOR U4077 ( .A(n2882), .B(n2550), .Z(n2552) );
  XNOR U4078 ( .A(n2883), .B(n2884), .Z(n2550) );
  AND U4079 ( .A(n2885), .B(n2886), .Z(n2883) );
  AND U4080 ( .A(b[3]), .B(a[52]), .Z(n2882) );
  NAND U4081 ( .A(a[55]), .B(b[0]), .Z(n2237) );
  XNOR U4082 ( .A(n2566), .B(n2567), .Z(c[54]) );
  XNOR U4083 ( .A(n2881), .B(n2880), .Z(n2567) );
  XOR U4084 ( .A(n2878), .B(n2887), .Z(n2880) );
  NAND U4085 ( .A(b[1]), .B(a[53]), .Z(n2887) );
  XNOR U4086 ( .A(n2886), .B(n2888), .Z(n2881) );
  XNOR U4087 ( .A(n2878), .B(n2885), .Z(n2888) );
  XNOR U4088 ( .A(n2889), .B(n2884), .Z(n2885) );
  AND U4089 ( .A(b[2]), .B(a[52]), .Z(n2889) );
  ANDN U4090 ( .B(n2890), .A(n2891), .Z(n2878) );
  XOR U4091 ( .A(n2884), .B(n2876), .Z(n2892) );
  XNOR U4092 ( .A(n2875), .B(n2871), .Z(n2893) );
  XNOR U4093 ( .A(n2870), .B(n2866), .Z(n2894) );
  XNOR U4094 ( .A(n2865), .B(n2861), .Z(n2895) );
  XNOR U4095 ( .A(n2860), .B(n2856), .Z(n2896) );
  XNOR U4096 ( .A(n2855), .B(n2851), .Z(n2897) );
  XNOR U4097 ( .A(n2850), .B(n2846), .Z(n2898) );
  XNOR U4098 ( .A(n2845), .B(n2841), .Z(n2899) );
  XNOR U4099 ( .A(n2840), .B(n2836), .Z(n2900) );
  XNOR U4100 ( .A(n2835), .B(n2831), .Z(n2901) );
  XNOR U4101 ( .A(n2830), .B(n2826), .Z(n2902) );
  XNOR U4102 ( .A(n2825), .B(n2821), .Z(n2903) );
  XNOR U4103 ( .A(n2820), .B(n2816), .Z(n2904) );
  XNOR U4104 ( .A(n2815), .B(n2811), .Z(n2905) );
  XNOR U4105 ( .A(n2810), .B(n2806), .Z(n2906) );
  XNOR U4106 ( .A(n2907), .B(n2908), .Z(n2806) );
  XNOR U4107 ( .A(n2797), .B(n2796), .Z(n2908) );
  XOR U4108 ( .A(n2909), .B(n2795), .Z(n2796) );
  AND U4109 ( .A(b[18]), .B(a[36]), .Z(n2909) );
  XNOR U4110 ( .A(n2795), .B(n2801), .Z(n2910) );
  XNOR U4111 ( .A(n2800), .B(n2792), .Z(n2911) );
  XNOR U4112 ( .A(n2791), .B(n2787), .Z(n2912) );
  XNOR U4113 ( .A(n2786), .B(n2782), .Z(n2913) );
  XNOR U4114 ( .A(n2781), .B(n2777), .Z(n2914) );
  XNOR U4115 ( .A(n2768), .B(n2767), .Z(n2915) );
  XOR U4116 ( .A(n2916), .B(n2766), .Z(n2767) );
  AND U4117 ( .A(b[24]), .B(a[30]), .Z(n2916) );
  XNOR U4118 ( .A(n2766), .B(n2772), .Z(n2917) );
  XNOR U4119 ( .A(n2771), .B(n2763), .Z(n2918) );
  XNOR U4120 ( .A(n2762), .B(n2758), .Z(n2919) );
  XNOR U4121 ( .A(n2757), .B(n2753), .Z(n2920) );
  XNOR U4122 ( .A(n2752), .B(n2748), .Z(n2921) );
  XNOR U4123 ( .A(n2739), .B(n2738), .Z(n2922) );
  XOR U4124 ( .A(n2923), .B(n2737), .Z(n2738) );
  AND U4125 ( .A(b[30]), .B(a[24]), .Z(n2923) );
  XNOR U4126 ( .A(n2737), .B(n2743), .Z(n2924) );
  XNOR U4127 ( .A(n2742), .B(n2734), .Z(n2925) );
  XNOR U4128 ( .A(n2733), .B(n2729), .Z(n2926) );
  XNOR U4129 ( .A(n2728), .B(n2724), .Z(n2927) );
  XNOR U4130 ( .A(n2723), .B(n2719), .Z(n2928) );
  XNOR U4131 ( .A(n2710), .B(n2709), .Z(n2929) );
  XOR U4132 ( .A(n2930), .B(n2708), .Z(n2709) );
  AND U4133 ( .A(b[36]), .B(a[18]), .Z(n2930) );
  XNOR U4134 ( .A(n2708), .B(n2714), .Z(n2931) );
  XNOR U4135 ( .A(n2713), .B(n2705), .Z(n2932) );
  XNOR U4136 ( .A(n2704), .B(n2700), .Z(n2933) );
  XNOR U4137 ( .A(n2699), .B(n2695), .Z(n2934) );
  XNOR U4138 ( .A(n2694), .B(n2690), .Z(n2935) );
  XNOR U4139 ( .A(n2681), .B(n2680), .Z(n2936) );
  XOR U4140 ( .A(n2937), .B(n2679), .Z(n2680) );
  AND U4141 ( .A(b[42]), .B(a[12]), .Z(n2937) );
  XNOR U4142 ( .A(n2679), .B(n2685), .Z(n2938) );
  XNOR U4143 ( .A(n2684), .B(n2676), .Z(n2939) );
  XNOR U4144 ( .A(n2675), .B(n2671), .Z(n2940) );
  XNOR U4145 ( .A(n2670), .B(n2666), .Z(n2941) );
  XNOR U4146 ( .A(n2665), .B(n2661), .Z(n2942) );
  XNOR U4147 ( .A(n2652), .B(n2651), .Z(n2943) );
  XOR U4148 ( .A(n2944), .B(n2650), .Z(n2651) );
  AND U4149 ( .A(a[6]), .B(b[48]), .Z(n2944) );
  XNOR U4150 ( .A(n2650), .B(n2656), .Z(n2945) );
  XNOR U4151 ( .A(n2655), .B(n2647), .Z(n2946) );
  XNOR U4152 ( .A(n2646), .B(n2642), .Z(n2947) );
  XNOR U4153 ( .A(n2641), .B(n2637), .Z(n2948) );
  XNOR U4154 ( .A(n2636), .B(n2632), .Z(n2949) );
  XOR U4155 ( .A(n2950), .B(n2631), .Z(n2632) );
  AND U4156 ( .A(a[0]), .B(b[54]), .Z(n2950) );
  XNOR U4157 ( .A(n2951), .B(n2631), .Z(n2633) );
  XNOR U4158 ( .A(n2952), .B(n2953), .Z(n2631) );
  ANDN U4159 ( .B(n2954), .A(n2955), .Z(n2952) );
  AND U4160 ( .A(a[1]), .B(b[53]), .Z(n2951) );
  XNOR U4161 ( .A(n2956), .B(n2636), .Z(n2638) );
  XOR U4162 ( .A(n2957), .B(n2958), .Z(n2636) );
  ANDN U4163 ( .B(n2959), .A(n2960), .Z(n2957) );
  AND U4164 ( .A(a[2]), .B(b[52]), .Z(n2956) );
  XNOR U4165 ( .A(n2961), .B(n2641), .Z(n2643) );
  XOR U4166 ( .A(n2962), .B(n2963), .Z(n2641) );
  ANDN U4167 ( .B(n2964), .A(n2965), .Z(n2962) );
  AND U4168 ( .A(a[3]), .B(b[51]), .Z(n2961) );
  XNOR U4169 ( .A(n2966), .B(n2646), .Z(n2648) );
  XOR U4170 ( .A(n2967), .B(n2968), .Z(n2646) );
  ANDN U4171 ( .B(n2969), .A(n2970), .Z(n2967) );
  AND U4172 ( .A(a[4]), .B(b[50]), .Z(n2966) );
  XOR U4173 ( .A(n2971), .B(n2972), .Z(n2650) );
  AND U4174 ( .A(n2973), .B(n2974), .Z(n2971) );
  XNOR U4175 ( .A(n2975), .B(n2655), .Z(n2657) );
  XOR U4176 ( .A(n2976), .B(n2977), .Z(n2655) );
  ANDN U4177 ( .B(n2978), .A(n2979), .Z(n2976) );
  AND U4178 ( .A(a[5]), .B(b[49]), .Z(n2975) );
  XOR U4179 ( .A(n2980), .B(n2660), .Z(n2662) );
  XOR U4180 ( .A(n2981), .B(n2982), .Z(n2660) );
  ANDN U4181 ( .B(n2983), .A(n2984), .Z(n2981) );
  AND U4182 ( .A(a[7]), .B(b[47]), .Z(n2980) );
  XNOR U4183 ( .A(n2985), .B(n2665), .Z(n2667) );
  XOR U4184 ( .A(n2986), .B(n2987), .Z(n2665) );
  ANDN U4185 ( .B(n2988), .A(n2989), .Z(n2986) );
  AND U4186 ( .A(a[8]), .B(b[46]), .Z(n2985) );
  XNOR U4187 ( .A(n2990), .B(n2670), .Z(n2672) );
  XOR U4188 ( .A(n2991), .B(n2992), .Z(n2670) );
  ANDN U4189 ( .B(n2993), .A(n2994), .Z(n2991) );
  AND U4190 ( .A(a[9]), .B(b[45]), .Z(n2990) );
  XNOR U4191 ( .A(n2995), .B(n2675), .Z(n2677) );
  XOR U4192 ( .A(n2996), .B(n2997), .Z(n2675) );
  ANDN U4193 ( .B(n2998), .A(n2999), .Z(n2996) );
  AND U4194 ( .A(b[44]), .B(a[10]), .Z(n2995) );
  XOR U4195 ( .A(n3000), .B(n3001), .Z(n2679) );
  AND U4196 ( .A(n3002), .B(n3003), .Z(n3000) );
  XNOR U4197 ( .A(n3004), .B(n2684), .Z(n2686) );
  XOR U4198 ( .A(n3005), .B(n3006), .Z(n2684) );
  ANDN U4199 ( .B(n3007), .A(n3008), .Z(n3005) );
  AND U4200 ( .A(b[43]), .B(a[11]), .Z(n3004) );
  XOR U4201 ( .A(n3009), .B(n2689), .Z(n2691) );
  XOR U4202 ( .A(n3010), .B(n3011), .Z(n2689) );
  ANDN U4203 ( .B(n3012), .A(n3013), .Z(n3010) );
  AND U4204 ( .A(b[41]), .B(a[13]), .Z(n3009) );
  XNOR U4205 ( .A(n3014), .B(n2694), .Z(n2696) );
  XOR U4206 ( .A(n3015), .B(n3016), .Z(n2694) );
  ANDN U4207 ( .B(n3017), .A(n3018), .Z(n3015) );
  AND U4208 ( .A(b[40]), .B(a[14]), .Z(n3014) );
  XNOR U4209 ( .A(n3019), .B(n2699), .Z(n2701) );
  XOR U4210 ( .A(n3020), .B(n3021), .Z(n2699) );
  ANDN U4211 ( .B(n3022), .A(n3023), .Z(n3020) );
  AND U4212 ( .A(a[15]), .B(b[39]), .Z(n3019) );
  XNOR U4213 ( .A(n3024), .B(n2704), .Z(n2706) );
  XOR U4214 ( .A(n3025), .B(n3026), .Z(n2704) );
  ANDN U4215 ( .B(n3027), .A(n3028), .Z(n3025) );
  AND U4216 ( .A(b[38]), .B(a[16]), .Z(n3024) );
  XOR U4217 ( .A(n3029), .B(n3030), .Z(n2708) );
  AND U4218 ( .A(n3031), .B(n3032), .Z(n3029) );
  XNOR U4219 ( .A(n3033), .B(n2713), .Z(n2715) );
  XOR U4220 ( .A(n3034), .B(n3035), .Z(n2713) );
  ANDN U4221 ( .B(n3036), .A(n3037), .Z(n3034) );
  AND U4222 ( .A(b[37]), .B(a[17]), .Z(n3033) );
  XOR U4223 ( .A(n3038), .B(n2718), .Z(n2720) );
  XOR U4224 ( .A(n3039), .B(n3040), .Z(n2718) );
  ANDN U4225 ( .B(n3041), .A(n3042), .Z(n3039) );
  AND U4226 ( .A(b[35]), .B(a[19]), .Z(n3038) );
  XNOR U4227 ( .A(n3043), .B(n2723), .Z(n2725) );
  XOR U4228 ( .A(n3044), .B(n3045), .Z(n2723) );
  ANDN U4229 ( .B(n3046), .A(n3047), .Z(n3044) );
  AND U4230 ( .A(b[34]), .B(a[20]), .Z(n3043) );
  XNOR U4231 ( .A(n3048), .B(n2728), .Z(n2730) );
  XOR U4232 ( .A(n3049), .B(n3050), .Z(n2728) );
  ANDN U4233 ( .B(n3051), .A(n3052), .Z(n3049) );
  AND U4234 ( .A(a[21]), .B(b[33]), .Z(n3048) );
  XNOR U4235 ( .A(n3053), .B(n2733), .Z(n2735) );
  XOR U4236 ( .A(n3054), .B(n3055), .Z(n2733) );
  ANDN U4237 ( .B(n3056), .A(n3057), .Z(n3054) );
  AND U4238 ( .A(b[32]), .B(a[22]), .Z(n3053) );
  XOR U4239 ( .A(n3058), .B(n3059), .Z(n2737) );
  AND U4240 ( .A(n3060), .B(n3061), .Z(n3058) );
  XNOR U4241 ( .A(n3062), .B(n2742), .Z(n2744) );
  XOR U4242 ( .A(n3063), .B(n3064), .Z(n2742) );
  ANDN U4243 ( .B(n3065), .A(n3066), .Z(n3063) );
  AND U4244 ( .A(b[31]), .B(a[23]), .Z(n3062) );
  XOR U4245 ( .A(n3067), .B(n2747), .Z(n2749) );
  XOR U4246 ( .A(n3068), .B(n3069), .Z(n2747) );
  ANDN U4247 ( .B(n3070), .A(n3071), .Z(n3068) );
  AND U4248 ( .A(b[29]), .B(a[25]), .Z(n3067) );
  XNOR U4249 ( .A(n3072), .B(n2752), .Z(n2754) );
  XOR U4250 ( .A(n3073), .B(n3074), .Z(n2752) );
  ANDN U4251 ( .B(n3075), .A(n3076), .Z(n3073) );
  AND U4252 ( .A(b[28]), .B(a[26]), .Z(n3072) );
  XNOR U4253 ( .A(n3077), .B(n2757), .Z(n2759) );
  XOR U4254 ( .A(n3078), .B(n3079), .Z(n2757) );
  ANDN U4255 ( .B(n3080), .A(n3081), .Z(n3078) );
  AND U4256 ( .A(a[27]), .B(b[27]), .Z(n3077) );
  XNOR U4257 ( .A(n3082), .B(n2762), .Z(n2764) );
  XOR U4258 ( .A(n3083), .B(n3084), .Z(n2762) );
  ANDN U4259 ( .B(n3085), .A(n3086), .Z(n3083) );
  AND U4260 ( .A(b[26]), .B(a[28]), .Z(n3082) );
  XOR U4261 ( .A(n3087), .B(n3088), .Z(n2766) );
  AND U4262 ( .A(n3089), .B(n3090), .Z(n3087) );
  XNOR U4263 ( .A(n3091), .B(n2771), .Z(n2773) );
  XOR U4264 ( .A(n3092), .B(n3093), .Z(n2771) );
  ANDN U4265 ( .B(n3094), .A(n3095), .Z(n3092) );
  AND U4266 ( .A(b[25]), .B(a[29]), .Z(n3091) );
  XOR U4267 ( .A(n3096), .B(n2776), .Z(n2778) );
  XOR U4268 ( .A(n3097), .B(n3098), .Z(n2776) );
  ANDN U4269 ( .B(n3099), .A(n3100), .Z(n3097) );
  AND U4270 ( .A(b[23]), .B(a[31]), .Z(n3096) );
  XNOR U4271 ( .A(n3101), .B(n2781), .Z(n2783) );
  XOR U4272 ( .A(n3102), .B(n3103), .Z(n2781) );
  ANDN U4273 ( .B(n3104), .A(n3105), .Z(n3102) );
  AND U4274 ( .A(b[22]), .B(a[32]), .Z(n3101) );
  XNOR U4275 ( .A(n3106), .B(n2786), .Z(n2788) );
  XOR U4276 ( .A(n3107), .B(n3108), .Z(n2786) );
  ANDN U4277 ( .B(n3109), .A(n3110), .Z(n3107) );
  AND U4278 ( .A(a[33]), .B(b[21]), .Z(n3106) );
  XNOR U4279 ( .A(n3111), .B(n2791), .Z(n2793) );
  XOR U4280 ( .A(n3112), .B(n3113), .Z(n2791) );
  ANDN U4281 ( .B(n3114), .A(n3115), .Z(n3112) );
  AND U4282 ( .A(b[20]), .B(a[34]), .Z(n3111) );
  XOR U4283 ( .A(n3116), .B(n3117), .Z(n2795) );
  AND U4284 ( .A(n3118), .B(n3119), .Z(n3116) );
  XNOR U4285 ( .A(n3120), .B(n2800), .Z(n2802) );
  XOR U4286 ( .A(n3121), .B(n3122), .Z(n2800) );
  ANDN U4287 ( .B(n3123), .A(n3124), .Z(n3121) );
  AND U4288 ( .A(b[19]), .B(a[35]), .Z(n3120) );
  IV U4289 ( .A(n2805), .Z(n2907) );
  XOR U4290 ( .A(n3125), .B(n2805), .Z(n2807) );
  XOR U4291 ( .A(n3126), .B(n3127), .Z(n2805) );
  ANDN U4292 ( .B(n3128), .A(n3129), .Z(n3126) );
  AND U4293 ( .A(b[17]), .B(a[37]), .Z(n3125) );
  XNOR U4294 ( .A(n3130), .B(n2810), .Z(n2812) );
  XOR U4295 ( .A(n3131), .B(n3132), .Z(n2810) );
  ANDN U4296 ( .B(n3133), .A(n3134), .Z(n3131) );
  AND U4297 ( .A(b[16]), .B(a[38]), .Z(n3130) );
  XNOR U4298 ( .A(n3135), .B(n2815), .Z(n2817) );
  XOR U4299 ( .A(n3136), .B(n3137), .Z(n2815) );
  ANDN U4300 ( .B(n3138), .A(n3139), .Z(n3136) );
  AND U4301 ( .A(a[39]), .B(b[15]), .Z(n3135) );
  XNOR U4302 ( .A(n3140), .B(n2820), .Z(n2822) );
  XOR U4303 ( .A(n3141), .B(n3142), .Z(n2820) );
  ANDN U4304 ( .B(n3143), .A(n3144), .Z(n3141) );
  AND U4305 ( .A(b[14]), .B(a[40]), .Z(n3140) );
  XNOR U4306 ( .A(n3145), .B(n2825), .Z(n2827) );
  XOR U4307 ( .A(n3146), .B(n3147), .Z(n2825) );
  ANDN U4308 ( .B(n3148), .A(n3149), .Z(n3146) );
  AND U4309 ( .A(b[13]), .B(a[41]), .Z(n3145) );
  XNOR U4310 ( .A(n3150), .B(n2830), .Z(n2832) );
  XOR U4311 ( .A(n3151), .B(n3152), .Z(n2830) );
  ANDN U4312 ( .B(n3153), .A(n3154), .Z(n3151) );
  AND U4313 ( .A(b[12]), .B(a[42]), .Z(n3150) );
  XNOR U4314 ( .A(n3155), .B(n2835), .Z(n2837) );
  XOR U4315 ( .A(n3156), .B(n3157), .Z(n2835) );
  ANDN U4316 ( .B(n3158), .A(n3159), .Z(n3156) );
  AND U4317 ( .A(b[11]), .B(a[43]), .Z(n3155) );
  XNOR U4318 ( .A(n3160), .B(n2840), .Z(n2842) );
  XOR U4319 ( .A(n3161), .B(n3162), .Z(n2840) );
  ANDN U4320 ( .B(n3163), .A(n3164), .Z(n3161) );
  AND U4321 ( .A(b[10]), .B(a[44]), .Z(n3160) );
  XNOR U4322 ( .A(n3165), .B(n2845), .Z(n2847) );
  XOR U4323 ( .A(n3166), .B(n3167), .Z(n2845) );
  ANDN U4324 ( .B(n3168), .A(n3169), .Z(n3166) );
  AND U4325 ( .A(b[9]), .B(a[45]), .Z(n3165) );
  XNOR U4326 ( .A(n3170), .B(n2850), .Z(n2852) );
  XOR U4327 ( .A(n3171), .B(n3172), .Z(n2850) );
  ANDN U4328 ( .B(n3173), .A(n3174), .Z(n3171) );
  AND U4329 ( .A(b[8]), .B(a[46]), .Z(n3170) );
  XNOR U4330 ( .A(n3175), .B(n2855), .Z(n2857) );
  XOR U4331 ( .A(n3176), .B(n3177), .Z(n2855) );
  ANDN U4332 ( .B(n3178), .A(n3179), .Z(n3176) );
  AND U4333 ( .A(b[7]), .B(a[47]), .Z(n3175) );
  XNOR U4334 ( .A(n3180), .B(n2860), .Z(n2862) );
  XOR U4335 ( .A(n3181), .B(n3182), .Z(n2860) );
  ANDN U4336 ( .B(n3183), .A(n3184), .Z(n3181) );
  AND U4337 ( .A(b[6]), .B(a[48]), .Z(n3180) );
  XNOR U4338 ( .A(n3185), .B(n2865), .Z(n2867) );
  XOR U4339 ( .A(n3186), .B(n3187), .Z(n2865) );
  ANDN U4340 ( .B(n3188), .A(n3189), .Z(n3186) );
  AND U4341 ( .A(b[5]), .B(a[49]), .Z(n3185) );
  XNOR U4342 ( .A(n3190), .B(n2870), .Z(n2872) );
  XOR U4343 ( .A(n3191), .B(n3192), .Z(n2870) );
  ANDN U4344 ( .B(n3193), .A(n3194), .Z(n3191) );
  AND U4345 ( .A(b[4]), .B(a[50]), .Z(n3190) );
  XNOR U4346 ( .A(n3195), .B(n3196), .Z(n2884) );
  NANDN U4347 ( .A(n3197), .B(n3198), .Z(n3196) );
  XNOR U4348 ( .A(n3199), .B(n2875), .Z(n2877) );
  XNOR U4349 ( .A(n3200), .B(n3201), .Z(n2875) );
  AND U4350 ( .A(n3202), .B(n3203), .Z(n3200) );
  AND U4351 ( .A(b[3]), .B(a[51]), .Z(n3199) );
  NAND U4352 ( .A(a[54]), .B(b[0]), .Z(n2566) );
  XNOR U4353 ( .A(n2891), .B(n2890), .Z(c[53]) );
  XNOR U4354 ( .A(n3197), .B(n3198), .Z(n2890) );
  XOR U4355 ( .A(n3195), .B(n3204), .Z(n3198) );
  NAND U4356 ( .A(b[1]), .B(a[52]), .Z(n3204) );
  XOR U4357 ( .A(n3203), .B(n3205), .Z(n3197) );
  XOR U4358 ( .A(n3195), .B(n3202), .Z(n3205) );
  XNOR U4359 ( .A(n3206), .B(n3201), .Z(n3202) );
  AND U4360 ( .A(b[2]), .B(a[51]), .Z(n3206) );
  NANDN U4361 ( .A(n3207), .B(n3208), .Z(n3195) );
  XOR U4362 ( .A(n3201), .B(n3193), .Z(n3209) );
  XNOR U4363 ( .A(n3192), .B(n3188), .Z(n3210) );
  XNOR U4364 ( .A(n3187), .B(n3183), .Z(n3211) );
  XNOR U4365 ( .A(n3182), .B(n3178), .Z(n3212) );
  XNOR U4366 ( .A(n3177), .B(n3173), .Z(n3213) );
  XNOR U4367 ( .A(n3172), .B(n3168), .Z(n3214) );
  XNOR U4368 ( .A(n3167), .B(n3163), .Z(n3215) );
  XNOR U4369 ( .A(n3162), .B(n3158), .Z(n3216) );
  XNOR U4370 ( .A(n3157), .B(n3153), .Z(n3217) );
  XNOR U4371 ( .A(n3152), .B(n3148), .Z(n3218) );
  XNOR U4372 ( .A(n3147), .B(n3143), .Z(n3219) );
  XNOR U4373 ( .A(n3142), .B(n3138), .Z(n3220) );
  XNOR U4374 ( .A(n3137), .B(n3133), .Z(n3221) );
  XNOR U4375 ( .A(n3132), .B(n3128), .Z(n3222) );
  XNOR U4376 ( .A(n3119), .B(n3118), .Z(n3223) );
  XOR U4377 ( .A(n3224), .B(n3117), .Z(n3118) );
  AND U4378 ( .A(b[17]), .B(a[36]), .Z(n3224) );
  XNOR U4379 ( .A(n3117), .B(n3123), .Z(n3225) );
  XNOR U4380 ( .A(n3122), .B(n3114), .Z(n3226) );
  XNOR U4381 ( .A(n3113), .B(n3109), .Z(n3227) );
  XNOR U4382 ( .A(n3108), .B(n3104), .Z(n3228) );
  XNOR U4383 ( .A(n3103), .B(n3099), .Z(n3229) );
  XNOR U4384 ( .A(n3090), .B(n3089), .Z(n3230) );
  XOR U4385 ( .A(n3231), .B(n3088), .Z(n3089) );
  AND U4386 ( .A(b[23]), .B(a[30]), .Z(n3231) );
  XNOR U4387 ( .A(n3088), .B(n3094), .Z(n3232) );
  XNOR U4388 ( .A(n3093), .B(n3085), .Z(n3233) );
  XNOR U4389 ( .A(n3084), .B(n3080), .Z(n3234) );
  XNOR U4390 ( .A(n3079), .B(n3075), .Z(n3235) );
  XNOR U4391 ( .A(n3074), .B(n3070), .Z(n3236) );
  XNOR U4392 ( .A(n3061), .B(n3060), .Z(n3237) );
  XOR U4393 ( .A(n3238), .B(n3059), .Z(n3060) );
  AND U4394 ( .A(b[29]), .B(a[24]), .Z(n3238) );
  XNOR U4395 ( .A(n3059), .B(n3065), .Z(n3239) );
  XNOR U4396 ( .A(n3064), .B(n3056), .Z(n3240) );
  XNOR U4397 ( .A(n3055), .B(n3051), .Z(n3241) );
  XNOR U4398 ( .A(n3050), .B(n3046), .Z(n3242) );
  XNOR U4399 ( .A(n3045), .B(n3041), .Z(n3243) );
  XNOR U4400 ( .A(n3032), .B(n3031), .Z(n3244) );
  XOR U4401 ( .A(n3245), .B(n3030), .Z(n3031) );
  AND U4402 ( .A(b[35]), .B(a[18]), .Z(n3245) );
  XNOR U4403 ( .A(n3030), .B(n3036), .Z(n3246) );
  XNOR U4404 ( .A(n3035), .B(n3027), .Z(n3247) );
  XNOR U4405 ( .A(n3026), .B(n3022), .Z(n3248) );
  XNOR U4406 ( .A(n3021), .B(n3017), .Z(n3249) );
  XNOR U4407 ( .A(n3016), .B(n3012), .Z(n3250) );
  XNOR U4408 ( .A(n3003), .B(n3002), .Z(n3251) );
  XOR U4409 ( .A(n3252), .B(n3001), .Z(n3002) );
  AND U4410 ( .A(b[41]), .B(a[12]), .Z(n3252) );
  XNOR U4411 ( .A(n3001), .B(n3007), .Z(n3253) );
  XNOR U4412 ( .A(n3006), .B(n2998), .Z(n3254) );
  XNOR U4413 ( .A(n2997), .B(n2993), .Z(n3255) );
  XNOR U4414 ( .A(n2992), .B(n2988), .Z(n3256) );
  XNOR U4415 ( .A(n2987), .B(n2983), .Z(n3257) );
  XNOR U4416 ( .A(n2974), .B(n2973), .Z(n3258) );
  XOR U4417 ( .A(n3259), .B(n2972), .Z(n2973) );
  AND U4418 ( .A(a[6]), .B(b[47]), .Z(n3259) );
  XNOR U4419 ( .A(n2972), .B(n2978), .Z(n3260) );
  XNOR U4420 ( .A(n2977), .B(n2969), .Z(n3261) );
  XNOR U4421 ( .A(n2968), .B(n2964), .Z(n3262) );
  XNOR U4422 ( .A(n2963), .B(n2959), .Z(n3263) );
  XNOR U4423 ( .A(n2958), .B(n2954), .Z(n3264) );
  XNOR U4424 ( .A(n3265), .B(n2953), .Z(n2954) );
  AND U4425 ( .A(a[0]), .B(b[53]), .Z(n3265) );
  XOR U4426 ( .A(n3266), .B(n2953), .Z(n2955) );
  XNOR U4427 ( .A(n3267), .B(n3268), .Z(n2953) );
  ANDN U4428 ( .B(n3269), .A(n3270), .Z(n3267) );
  AND U4429 ( .A(a[1]), .B(b[52]), .Z(n3266) );
  XNOR U4430 ( .A(n3271), .B(n2958), .Z(n2960) );
  XOR U4431 ( .A(n3272), .B(n3273), .Z(n2958) );
  ANDN U4432 ( .B(n3274), .A(n3275), .Z(n3272) );
  AND U4433 ( .A(a[2]), .B(b[51]), .Z(n3271) );
  XNOR U4434 ( .A(n3276), .B(n2963), .Z(n2965) );
  XOR U4435 ( .A(n3277), .B(n3278), .Z(n2963) );
  ANDN U4436 ( .B(n3279), .A(n3280), .Z(n3277) );
  AND U4437 ( .A(a[3]), .B(b[50]), .Z(n3276) );
  XNOR U4438 ( .A(n3281), .B(n2968), .Z(n2970) );
  XOR U4439 ( .A(n3282), .B(n3283), .Z(n2968) );
  ANDN U4440 ( .B(n3284), .A(n3285), .Z(n3282) );
  AND U4441 ( .A(a[4]), .B(b[49]), .Z(n3281) );
  XOR U4442 ( .A(n3286), .B(n3287), .Z(n2972) );
  AND U4443 ( .A(n3288), .B(n3289), .Z(n3286) );
  XNOR U4444 ( .A(n3290), .B(n2977), .Z(n2979) );
  XOR U4445 ( .A(n3291), .B(n3292), .Z(n2977) );
  ANDN U4446 ( .B(n3293), .A(n3294), .Z(n3291) );
  AND U4447 ( .A(a[5]), .B(b[48]), .Z(n3290) );
  XOR U4448 ( .A(n3295), .B(n2982), .Z(n2984) );
  XOR U4449 ( .A(n3296), .B(n3297), .Z(n2982) );
  ANDN U4450 ( .B(n3298), .A(n3299), .Z(n3296) );
  AND U4451 ( .A(a[7]), .B(b[46]), .Z(n3295) );
  XNOR U4452 ( .A(n3300), .B(n2987), .Z(n2989) );
  XOR U4453 ( .A(n3301), .B(n3302), .Z(n2987) );
  ANDN U4454 ( .B(n3303), .A(n3304), .Z(n3301) );
  AND U4455 ( .A(a[8]), .B(b[45]), .Z(n3300) );
  XNOR U4456 ( .A(n3305), .B(n2992), .Z(n2994) );
  XOR U4457 ( .A(n3306), .B(n3307), .Z(n2992) );
  ANDN U4458 ( .B(n3308), .A(n3309), .Z(n3306) );
  AND U4459 ( .A(a[9]), .B(b[44]), .Z(n3305) );
  XNOR U4460 ( .A(n3310), .B(n2997), .Z(n2999) );
  XOR U4461 ( .A(n3311), .B(n3312), .Z(n2997) );
  ANDN U4462 ( .B(n3313), .A(n3314), .Z(n3311) );
  AND U4463 ( .A(b[43]), .B(a[10]), .Z(n3310) );
  XOR U4464 ( .A(n3315), .B(n3316), .Z(n3001) );
  AND U4465 ( .A(n3317), .B(n3318), .Z(n3315) );
  XNOR U4466 ( .A(n3319), .B(n3006), .Z(n3008) );
  XOR U4467 ( .A(n3320), .B(n3321), .Z(n3006) );
  ANDN U4468 ( .B(n3322), .A(n3323), .Z(n3320) );
  AND U4469 ( .A(b[42]), .B(a[11]), .Z(n3319) );
  XOR U4470 ( .A(n3324), .B(n3011), .Z(n3013) );
  XOR U4471 ( .A(n3325), .B(n3326), .Z(n3011) );
  ANDN U4472 ( .B(n3327), .A(n3328), .Z(n3325) );
  AND U4473 ( .A(b[40]), .B(a[13]), .Z(n3324) );
  XNOR U4474 ( .A(n3329), .B(n3016), .Z(n3018) );
  XOR U4475 ( .A(n3330), .B(n3331), .Z(n3016) );
  ANDN U4476 ( .B(n3332), .A(n3333), .Z(n3330) );
  AND U4477 ( .A(a[14]), .B(b[39]), .Z(n3329) );
  XNOR U4478 ( .A(n3334), .B(n3021), .Z(n3023) );
  XOR U4479 ( .A(n3335), .B(n3336), .Z(n3021) );
  ANDN U4480 ( .B(n3337), .A(n3338), .Z(n3335) );
  AND U4481 ( .A(b[38]), .B(a[15]), .Z(n3334) );
  XNOR U4482 ( .A(n3339), .B(n3026), .Z(n3028) );
  XOR U4483 ( .A(n3340), .B(n3341), .Z(n3026) );
  ANDN U4484 ( .B(n3342), .A(n3343), .Z(n3340) );
  AND U4485 ( .A(b[37]), .B(a[16]), .Z(n3339) );
  XOR U4486 ( .A(n3344), .B(n3345), .Z(n3030) );
  AND U4487 ( .A(n3346), .B(n3347), .Z(n3344) );
  XNOR U4488 ( .A(n3348), .B(n3035), .Z(n3037) );
  XOR U4489 ( .A(n3349), .B(n3350), .Z(n3035) );
  ANDN U4490 ( .B(n3351), .A(n3352), .Z(n3349) );
  AND U4491 ( .A(b[36]), .B(a[17]), .Z(n3348) );
  XOR U4492 ( .A(n3353), .B(n3040), .Z(n3042) );
  XOR U4493 ( .A(n3354), .B(n3355), .Z(n3040) );
  ANDN U4494 ( .B(n3356), .A(n3357), .Z(n3354) );
  AND U4495 ( .A(b[34]), .B(a[19]), .Z(n3353) );
  XNOR U4496 ( .A(n3358), .B(n3045), .Z(n3047) );
  XOR U4497 ( .A(n3359), .B(n3360), .Z(n3045) );
  ANDN U4498 ( .B(n3361), .A(n3362), .Z(n3359) );
  AND U4499 ( .A(a[20]), .B(b[33]), .Z(n3358) );
  XNOR U4500 ( .A(n3363), .B(n3050), .Z(n3052) );
  XOR U4501 ( .A(n3364), .B(n3365), .Z(n3050) );
  ANDN U4502 ( .B(n3366), .A(n3367), .Z(n3364) );
  AND U4503 ( .A(b[32]), .B(a[21]), .Z(n3363) );
  XNOR U4504 ( .A(n3368), .B(n3055), .Z(n3057) );
  XOR U4505 ( .A(n3369), .B(n3370), .Z(n3055) );
  ANDN U4506 ( .B(n3371), .A(n3372), .Z(n3369) );
  AND U4507 ( .A(b[31]), .B(a[22]), .Z(n3368) );
  XOR U4508 ( .A(n3373), .B(n3374), .Z(n3059) );
  AND U4509 ( .A(n3375), .B(n3376), .Z(n3373) );
  XNOR U4510 ( .A(n3377), .B(n3064), .Z(n3066) );
  XOR U4511 ( .A(n3378), .B(n3379), .Z(n3064) );
  ANDN U4512 ( .B(n3380), .A(n3381), .Z(n3378) );
  AND U4513 ( .A(b[30]), .B(a[23]), .Z(n3377) );
  XOR U4514 ( .A(n3382), .B(n3069), .Z(n3071) );
  XOR U4515 ( .A(n3383), .B(n3384), .Z(n3069) );
  ANDN U4516 ( .B(n3385), .A(n3386), .Z(n3383) );
  AND U4517 ( .A(b[28]), .B(a[25]), .Z(n3382) );
  XNOR U4518 ( .A(n3387), .B(n3074), .Z(n3076) );
  XOR U4519 ( .A(n3388), .B(n3389), .Z(n3074) );
  ANDN U4520 ( .B(n3390), .A(n3391), .Z(n3388) );
  AND U4521 ( .A(a[26]), .B(b[27]), .Z(n3387) );
  XNOR U4522 ( .A(n3392), .B(n3079), .Z(n3081) );
  XOR U4523 ( .A(n3393), .B(n3394), .Z(n3079) );
  ANDN U4524 ( .B(n3395), .A(n3396), .Z(n3393) );
  AND U4525 ( .A(b[26]), .B(a[27]), .Z(n3392) );
  XNOR U4526 ( .A(n3397), .B(n3084), .Z(n3086) );
  XOR U4527 ( .A(n3398), .B(n3399), .Z(n3084) );
  ANDN U4528 ( .B(n3400), .A(n3401), .Z(n3398) );
  AND U4529 ( .A(b[25]), .B(a[28]), .Z(n3397) );
  XOR U4530 ( .A(n3402), .B(n3403), .Z(n3088) );
  AND U4531 ( .A(n3404), .B(n3405), .Z(n3402) );
  XNOR U4532 ( .A(n3406), .B(n3093), .Z(n3095) );
  XOR U4533 ( .A(n3407), .B(n3408), .Z(n3093) );
  ANDN U4534 ( .B(n3409), .A(n3410), .Z(n3407) );
  AND U4535 ( .A(b[24]), .B(a[29]), .Z(n3406) );
  XOR U4536 ( .A(n3411), .B(n3098), .Z(n3100) );
  XOR U4537 ( .A(n3412), .B(n3413), .Z(n3098) );
  ANDN U4538 ( .B(n3414), .A(n3415), .Z(n3412) );
  AND U4539 ( .A(b[22]), .B(a[31]), .Z(n3411) );
  XNOR U4540 ( .A(n3416), .B(n3103), .Z(n3105) );
  XOR U4541 ( .A(n3417), .B(n3418), .Z(n3103) );
  ANDN U4542 ( .B(n3419), .A(n3420), .Z(n3417) );
  AND U4543 ( .A(a[32]), .B(b[21]), .Z(n3416) );
  XNOR U4544 ( .A(n3421), .B(n3108), .Z(n3110) );
  XOR U4545 ( .A(n3422), .B(n3423), .Z(n3108) );
  ANDN U4546 ( .B(n3424), .A(n3425), .Z(n3422) );
  AND U4547 ( .A(b[20]), .B(a[33]), .Z(n3421) );
  XNOR U4548 ( .A(n3426), .B(n3113), .Z(n3115) );
  XOR U4549 ( .A(n3427), .B(n3428), .Z(n3113) );
  ANDN U4550 ( .B(n3429), .A(n3430), .Z(n3427) );
  AND U4551 ( .A(b[19]), .B(a[34]), .Z(n3426) );
  XOR U4552 ( .A(n3431), .B(n3432), .Z(n3117) );
  AND U4553 ( .A(n3433), .B(n3434), .Z(n3431) );
  XNOR U4554 ( .A(n3435), .B(n3122), .Z(n3124) );
  XOR U4555 ( .A(n3436), .B(n3437), .Z(n3122) );
  ANDN U4556 ( .B(n3438), .A(n3439), .Z(n3436) );
  AND U4557 ( .A(b[18]), .B(a[35]), .Z(n3435) );
  XOR U4558 ( .A(n3440), .B(n3127), .Z(n3129) );
  XOR U4559 ( .A(n3441), .B(n3442), .Z(n3127) );
  ANDN U4560 ( .B(n3443), .A(n3444), .Z(n3441) );
  AND U4561 ( .A(b[16]), .B(a[37]), .Z(n3440) );
  XNOR U4562 ( .A(n3445), .B(n3132), .Z(n3134) );
  XOR U4563 ( .A(n3446), .B(n3447), .Z(n3132) );
  ANDN U4564 ( .B(n3448), .A(n3449), .Z(n3446) );
  AND U4565 ( .A(a[38]), .B(b[15]), .Z(n3445) );
  XNOR U4566 ( .A(n3450), .B(n3137), .Z(n3139) );
  XOR U4567 ( .A(n3451), .B(n3452), .Z(n3137) );
  ANDN U4568 ( .B(n3453), .A(n3454), .Z(n3451) );
  AND U4569 ( .A(b[14]), .B(a[39]), .Z(n3450) );
  XNOR U4570 ( .A(n3455), .B(n3142), .Z(n3144) );
  XOR U4571 ( .A(n3456), .B(n3457), .Z(n3142) );
  ANDN U4572 ( .B(n3458), .A(n3459), .Z(n3456) );
  AND U4573 ( .A(b[13]), .B(a[40]), .Z(n3455) );
  XNOR U4574 ( .A(n3460), .B(n3147), .Z(n3149) );
  XOR U4575 ( .A(n3461), .B(n3462), .Z(n3147) );
  ANDN U4576 ( .B(n3463), .A(n3464), .Z(n3461) );
  AND U4577 ( .A(b[12]), .B(a[41]), .Z(n3460) );
  XNOR U4578 ( .A(n3465), .B(n3152), .Z(n3154) );
  XOR U4579 ( .A(n3466), .B(n3467), .Z(n3152) );
  ANDN U4580 ( .B(n3468), .A(n3469), .Z(n3466) );
  AND U4581 ( .A(b[11]), .B(a[42]), .Z(n3465) );
  XNOR U4582 ( .A(n3470), .B(n3157), .Z(n3159) );
  XOR U4583 ( .A(n3471), .B(n3472), .Z(n3157) );
  ANDN U4584 ( .B(n3473), .A(n3474), .Z(n3471) );
  AND U4585 ( .A(b[10]), .B(a[43]), .Z(n3470) );
  XNOR U4586 ( .A(n3475), .B(n3162), .Z(n3164) );
  XOR U4587 ( .A(n3476), .B(n3477), .Z(n3162) );
  ANDN U4588 ( .B(n3478), .A(n3479), .Z(n3476) );
  AND U4589 ( .A(b[9]), .B(a[44]), .Z(n3475) );
  XNOR U4590 ( .A(n3480), .B(n3167), .Z(n3169) );
  XOR U4591 ( .A(n3481), .B(n3482), .Z(n3167) );
  ANDN U4592 ( .B(n3483), .A(n3484), .Z(n3481) );
  AND U4593 ( .A(b[8]), .B(a[45]), .Z(n3480) );
  XNOR U4594 ( .A(n3485), .B(n3172), .Z(n3174) );
  XOR U4595 ( .A(n3486), .B(n3487), .Z(n3172) );
  ANDN U4596 ( .B(n3488), .A(n3489), .Z(n3486) );
  AND U4597 ( .A(b[7]), .B(a[46]), .Z(n3485) );
  XNOR U4598 ( .A(n3490), .B(n3177), .Z(n3179) );
  XOR U4599 ( .A(n3491), .B(n3492), .Z(n3177) );
  ANDN U4600 ( .B(n3493), .A(n3494), .Z(n3491) );
  AND U4601 ( .A(b[6]), .B(a[47]), .Z(n3490) );
  XNOR U4602 ( .A(n3495), .B(n3182), .Z(n3184) );
  XOR U4603 ( .A(n3496), .B(n3497), .Z(n3182) );
  ANDN U4604 ( .B(n3498), .A(n3499), .Z(n3496) );
  AND U4605 ( .A(b[5]), .B(a[48]), .Z(n3495) );
  XNOR U4606 ( .A(n3500), .B(n3187), .Z(n3189) );
  XOR U4607 ( .A(n3501), .B(n3502), .Z(n3187) );
  ANDN U4608 ( .B(n3503), .A(n3504), .Z(n3501) );
  AND U4609 ( .A(b[4]), .B(a[49]), .Z(n3500) );
  XNOR U4610 ( .A(n3505), .B(n3506), .Z(n3201) );
  NANDN U4611 ( .A(n3507), .B(n3508), .Z(n3506) );
  XNOR U4612 ( .A(n3509), .B(n3192), .Z(n3194) );
  XNOR U4613 ( .A(n3510), .B(n3511), .Z(n3192) );
  AND U4614 ( .A(n3512), .B(n3513), .Z(n3510) );
  AND U4615 ( .A(b[3]), .B(a[50]), .Z(n3509) );
  NAND U4616 ( .A(a[53]), .B(b[0]), .Z(n2891) );
  XNOR U4617 ( .A(n3207), .B(n3208), .Z(c[52]) );
  XNOR U4618 ( .A(n3507), .B(n3508), .Z(n3208) );
  XOR U4619 ( .A(n3505), .B(n3514), .Z(n3508) );
  NAND U4620 ( .A(b[1]), .B(a[51]), .Z(n3514) );
  XOR U4621 ( .A(n3513), .B(n3515), .Z(n3507) );
  XOR U4622 ( .A(n3505), .B(n3512), .Z(n3515) );
  XNOR U4623 ( .A(n3516), .B(n3511), .Z(n3512) );
  AND U4624 ( .A(b[2]), .B(a[50]), .Z(n3516) );
  NANDN U4625 ( .A(n3517), .B(n3518), .Z(n3505) );
  XOR U4626 ( .A(n3511), .B(n3503), .Z(n3519) );
  XNOR U4627 ( .A(n3502), .B(n3498), .Z(n3520) );
  XNOR U4628 ( .A(n3497), .B(n3493), .Z(n3521) );
  XNOR U4629 ( .A(n3492), .B(n3488), .Z(n3522) );
  XNOR U4630 ( .A(n3487), .B(n3483), .Z(n3523) );
  XNOR U4631 ( .A(n3482), .B(n3478), .Z(n3524) );
  XNOR U4632 ( .A(n3477), .B(n3473), .Z(n3525) );
  XNOR U4633 ( .A(n3472), .B(n3468), .Z(n3526) );
  XNOR U4634 ( .A(n3467), .B(n3463), .Z(n3527) );
  XNOR U4635 ( .A(n3462), .B(n3458), .Z(n3528) );
  XNOR U4636 ( .A(n3457), .B(n3453), .Z(n3529) );
  XNOR U4637 ( .A(n3452), .B(n3448), .Z(n3530) );
  XNOR U4638 ( .A(n3447), .B(n3443), .Z(n3531) );
  XNOR U4639 ( .A(n3434), .B(n3433), .Z(n3532) );
  XOR U4640 ( .A(n3533), .B(n3432), .Z(n3433) );
  AND U4641 ( .A(b[16]), .B(a[36]), .Z(n3533) );
  XNOR U4642 ( .A(n3432), .B(n3438), .Z(n3534) );
  XNOR U4643 ( .A(n3437), .B(n3429), .Z(n3535) );
  XNOR U4644 ( .A(n3428), .B(n3424), .Z(n3536) );
  XNOR U4645 ( .A(n3423), .B(n3419), .Z(n3537) );
  XNOR U4646 ( .A(n3418), .B(n3414), .Z(n3538) );
  XNOR U4647 ( .A(n3405), .B(n3404), .Z(n3539) );
  XOR U4648 ( .A(n3540), .B(n3403), .Z(n3404) );
  AND U4649 ( .A(b[22]), .B(a[30]), .Z(n3540) );
  XNOR U4650 ( .A(n3403), .B(n3409), .Z(n3541) );
  XNOR U4651 ( .A(n3408), .B(n3400), .Z(n3542) );
  XNOR U4652 ( .A(n3399), .B(n3395), .Z(n3543) );
  XNOR U4653 ( .A(n3394), .B(n3390), .Z(n3544) );
  XNOR U4654 ( .A(n3389), .B(n3385), .Z(n3545) );
  XNOR U4655 ( .A(n3376), .B(n3375), .Z(n3546) );
  XOR U4656 ( .A(n3547), .B(n3374), .Z(n3375) );
  AND U4657 ( .A(b[28]), .B(a[24]), .Z(n3547) );
  XNOR U4658 ( .A(n3374), .B(n3380), .Z(n3548) );
  XNOR U4659 ( .A(n3379), .B(n3371), .Z(n3549) );
  XNOR U4660 ( .A(n3370), .B(n3366), .Z(n3550) );
  XNOR U4661 ( .A(n3365), .B(n3361), .Z(n3551) );
  XNOR U4662 ( .A(n3360), .B(n3356), .Z(n3552) );
  XNOR U4663 ( .A(n3347), .B(n3346), .Z(n3553) );
  XOR U4664 ( .A(n3554), .B(n3345), .Z(n3346) );
  AND U4665 ( .A(b[34]), .B(a[18]), .Z(n3554) );
  XNOR U4666 ( .A(n3345), .B(n3351), .Z(n3555) );
  XNOR U4667 ( .A(n3350), .B(n3342), .Z(n3556) );
  XNOR U4668 ( .A(n3341), .B(n3337), .Z(n3557) );
  XNOR U4669 ( .A(n3336), .B(n3332), .Z(n3558) );
  XNOR U4670 ( .A(n3331), .B(n3327), .Z(n3559) );
  XNOR U4671 ( .A(n3318), .B(n3317), .Z(n3560) );
  XOR U4672 ( .A(n3561), .B(n3316), .Z(n3317) );
  AND U4673 ( .A(b[40]), .B(a[12]), .Z(n3561) );
  XNOR U4674 ( .A(n3316), .B(n3322), .Z(n3562) );
  XNOR U4675 ( .A(n3321), .B(n3313), .Z(n3563) );
  XNOR U4676 ( .A(n3312), .B(n3308), .Z(n3564) );
  XNOR U4677 ( .A(n3307), .B(n3303), .Z(n3565) );
  XNOR U4678 ( .A(n3302), .B(n3298), .Z(n3566) );
  XNOR U4679 ( .A(n3289), .B(n3288), .Z(n3567) );
  XOR U4680 ( .A(n3568), .B(n3287), .Z(n3288) );
  AND U4681 ( .A(a[6]), .B(b[46]), .Z(n3568) );
  XNOR U4682 ( .A(n3287), .B(n3293), .Z(n3569) );
  XNOR U4683 ( .A(n3292), .B(n3284), .Z(n3570) );
  XNOR U4684 ( .A(n3283), .B(n3279), .Z(n3571) );
  XNOR U4685 ( .A(n3278), .B(n3274), .Z(n3572) );
  XNOR U4686 ( .A(n3273), .B(n3269), .Z(n3573) );
  XOR U4687 ( .A(n3574), .B(n3268), .Z(n3269) );
  AND U4688 ( .A(a[0]), .B(b[52]), .Z(n3574) );
  XNOR U4689 ( .A(n3575), .B(n3268), .Z(n3270) );
  XNOR U4690 ( .A(n3576), .B(n3577), .Z(n3268) );
  ANDN U4691 ( .B(n3578), .A(n3579), .Z(n3576) );
  AND U4692 ( .A(a[1]), .B(b[51]), .Z(n3575) );
  XNOR U4693 ( .A(n3580), .B(n3273), .Z(n3275) );
  XOR U4694 ( .A(n3581), .B(n3582), .Z(n3273) );
  ANDN U4695 ( .B(n3583), .A(n3584), .Z(n3581) );
  AND U4696 ( .A(a[2]), .B(b[50]), .Z(n3580) );
  XNOR U4697 ( .A(n3585), .B(n3278), .Z(n3280) );
  XOR U4698 ( .A(n3586), .B(n3587), .Z(n3278) );
  ANDN U4699 ( .B(n3588), .A(n3589), .Z(n3586) );
  AND U4700 ( .A(a[3]), .B(b[49]), .Z(n3585) );
  XNOR U4701 ( .A(n3590), .B(n3283), .Z(n3285) );
  XOR U4702 ( .A(n3591), .B(n3592), .Z(n3283) );
  ANDN U4703 ( .B(n3593), .A(n3594), .Z(n3591) );
  AND U4704 ( .A(a[4]), .B(b[48]), .Z(n3590) );
  XOR U4705 ( .A(n3595), .B(n3596), .Z(n3287) );
  AND U4706 ( .A(n3597), .B(n3598), .Z(n3595) );
  XNOR U4707 ( .A(n3599), .B(n3292), .Z(n3294) );
  XOR U4708 ( .A(n3600), .B(n3601), .Z(n3292) );
  ANDN U4709 ( .B(n3602), .A(n3603), .Z(n3600) );
  AND U4710 ( .A(a[5]), .B(b[47]), .Z(n3599) );
  XOR U4711 ( .A(n3604), .B(n3297), .Z(n3299) );
  XOR U4712 ( .A(n3605), .B(n3606), .Z(n3297) );
  ANDN U4713 ( .B(n3607), .A(n3608), .Z(n3605) );
  AND U4714 ( .A(a[7]), .B(b[45]), .Z(n3604) );
  XNOR U4715 ( .A(n3609), .B(n3302), .Z(n3304) );
  XOR U4716 ( .A(n3610), .B(n3611), .Z(n3302) );
  ANDN U4717 ( .B(n3612), .A(n3613), .Z(n3610) );
  AND U4718 ( .A(a[8]), .B(b[44]), .Z(n3609) );
  XNOR U4719 ( .A(n3614), .B(n3307), .Z(n3309) );
  XOR U4720 ( .A(n3615), .B(n3616), .Z(n3307) );
  ANDN U4721 ( .B(n3617), .A(n3618), .Z(n3615) );
  AND U4722 ( .A(a[9]), .B(b[43]), .Z(n3614) );
  XNOR U4723 ( .A(n3619), .B(n3312), .Z(n3314) );
  XOR U4724 ( .A(n3620), .B(n3621), .Z(n3312) );
  ANDN U4725 ( .B(n3622), .A(n3623), .Z(n3620) );
  AND U4726 ( .A(b[42]), .B(a[10]), .Z(n3619) );
  XOR U4727 ( .A(n3624), .B(n3625), .Z(n3316) );
  AND U4728 ( .A(n3626), .B(n3627), .Z(n3624) );
  XNOR U4729 ( .A(n3628), .B(n3321), .Z(n3323) );
  XOR U4730 ( .A(n3629), .B(n3630), .Z(n3321) );
  ANDN U4731 ( .B(n3631), .A(n3632), .Z(n3629) );
  AND U4732 ( .A(b[41]), .B(a[11]), .Z(n3628) );
  XOR U4733 ( .A(n3633), .B(n3326), .Z(n3328) );
  XOR U4734 ( .A(n3634), .B(n3635), .Z(n3326) );
  ANDN U4735 ( .B(n3636), .A(n3637), .Z(n3634) );
  AND U4736 ( .A(a[13]), .B(b[39]), .Z(n3633) );
  XNOR U4737 ( .A(n3638), .B(n3331), .Z(n3333) );
  XOR U4738 ( .A(n3639), .B(n3640), .Z(n3331) );
  ANDN U4739 ( .B(n3641), .A(n3642), .Z(n3639) );
  AND U4740 ( .A(b[38]), .B(a[14]), .Z(n3638) );
  XNOR U4741 ( .A(n3643), .B(n3336), .Z(n3338) );
  XOR U4742 ( .A(n3644), .B(n3645), .Z(n3336) );
  ANDN U4743 ( .B(n3646), .A(n3647), .Z(n3644) );
  AND U4744 ( .A(b[37]), .B(a[15]), .Z(n3643) );
  XNOR U4745 ( .A(n3648), .B(n3341), .Z(n3343) );
  XOR U4746 ( .A(n3649), .B(n3650), .Z(n3341) );
  ANDN U4747 ( .B(n3651), .A(n3652), .Z(n3649) );
  AND U4748 ( .A(b[36]), .B(a[16]), .Z(n3648) );
  XOR U4749 ( .A(n3653), .B(n3654), .Z(n3345) );
  AND U4750 ( .A(n3655), .B(n3656), .Z(n3653) );
  XNOR U4751 ( .A(n3657), .B(n3350), .Z(n3352) );
  XOR U4752 ( .A(n3658), .B(n3659), .Z(n3350) );
  ANDN U4753 ( .B(n3660), .A(n3661), .Z(n3658) );
  AND U4754 ( .A(b[35]), .B(a[17]), .Z(n3657) );
  XOR U4755 ( .A(n3662), .B(n3355), .Z(n3357) );
  XOR U4756 ( .A(n3663), .B(n3664), .Z(n3355) );
  ANDN U4757 ( .B(n3665), .A(n3666), .Z(n3663) );
  AND U4758 ( .A(a[19]), .B(b[33]), .Z(n3662) );
  XNOR U4759 ( .A(n3667), .B(n3360), .Z(n3362) );
  XOR U4760 ( .A(n3668), .B(n3669), .Z(n3360) );
  ANDN U4761 ( .B(n3670), .A(n3671), .Z(n3668) );
  AND U4762 ( .A(b[32]), .B(a[20]), .Z(n3667) );
  XNOR U4763 ( .A(n3672), .B(n3365), .Z(n3367) );
  XOR U4764 ( .A(n3673), .B(n3674), .Z(n3365) );
  ANDN U4765 ( .B(n3675), .A(n3676), .Z(n3673) );
  AND U4766 ( .A(b[31]), .B(a[21]), .Z(n3672) );
  XNOR U4767 ( .A(n3677), .B(n3370), .Z(n3372) );
  XOR U4768 ( .A(n3678), .B(n3679), .Z(n3370) );
  ANDN U4769 ( .B(n3680), .A(n3681), .Z(n3678) );
  AND U4770 ( .A(b[30]), .B(a[22]), .Z(n3677) );
  XOR U4771 ( .A(n3682), .B(n3683), .Z(n3374) );
  AND U4772 ( .A(n3684), .B(n3685), .Z(n3682) );
  XNOR U4773 ( .A(n3686), .B(n3379), .Z(n3381) );
  XOR U4774 ( .A(n3687), .B(n3688), .Z(n3379) );
  ANDN U4775 ( .B(n3689), .A(n3690), .Z(n3687) );
  AND U4776 ( .A(b[29]), .B(a[23]), .Z(n3686) );
  XOR U4777 ( .A(n3691), .B(n3384), .Z(n3386) );
  XOR U4778 ( .A(n3692), .B(n3693), .Z(n3384) );
  ANDN U4779 ( .B(n3694), .A(n3695), .Z(n3692) );
  AND U4780 ( .A(a[25]), .B(b[27]), .Z(n3691) );
  XNOR U4781 ( .A(n3696), .B(n3389), .Z(n3391) );
  XOR U4782 ( .A(n3697), .B(n3698), .Z(n3389) );
  ANDN U4783 ( .B(n3699), .A(n3700), .Z(n3697) );
  AND U4784 ( .A(b[26]), .B(a[26]), .Z(n3696) );
  XNOR U4785 ( .A(n3701), .B(n3394), .Z(n3396) );
  XOR U4786 ( .A(n3702), .B(n3703), .Z(n3394) );
  ANDN U4787 ( .B(n3704), .A(n3705), .Z(n3702) );
  AND U4788 ( .A(b[25]), .B(a[27]), .Z(n3701) );
  XNOR U4789 ( .A(n3706), .B(n3399), .Z(n3401) );
  XOR U4790 ( .A(n3707), .B(n3708), .Z(n3399) );
  ANDN U4791 ( .B(n3709), .A(n3710), .Z(n3707) );
  AND U4792 ( .A(b[24]), .B(a[28]), .Z(n3706) );
  XOR U4793 ( .A(n3711), .B(n3712), .Z(n3403) );
  AND U4794 ( .A(n3713), .B(n3714), .Z(n3711) );
  XNOR U4795 ( .A(n3715), .B(n3408), .Z(n3410) );
  XOR U4796 ( .A(n3716), .B(n3717), .Z(n3408) );
  ANDN U4797 ( .B(n3718), .A(n3719), .Z(n3716) );
  AND U4798 ( .A(b[23]), .B(a[29]), .Z(n3715) );
  XOR U4799 ( .A(n3720), .B(n3413), .Z(n3415) );
  XOR U4800 ( .A(n3721), .B(n3722), .Z(n3413) );
  ANDN U4801 ( .B(n3723), .A(n3724), .Z(n3721) );
  AND U4802 ( .A(a[31]), .B(b[21]), .Z(n3720) );
  XNOR U4803 ( .A(n3725), .B(n3418), .Z(n3420) );
  XOR U4804 ( .A(n3726), .B(n3727), .Z(n3418) );
  ANDN U4805 ( .B(n3728), .A(n3729), .Z(n3726) );
  AND U4806 ( .A(b[20]), .B(a[32]), .Z(n3725) );
  XNOR U4807 ( .A(n3730), .B(n3423), .Z(n3425) );
  XOR U4808 ( .A(n3731), .B(n3732), .Z(n3423) );
  ANDN U4809 ( .B(n3733), .A(n3734), .Z(n3731) );
  AND U4810 ( .A(b[19]), .B(a[33]), .Z(n3730) );
  XNOR U4811 ( .A(n3735), .B(n3428), .Z(n3430) );
  XOR U4812 ( .A(n3736), .B(n3737), .Z(n3428) );
  ANDN U4813 ( .B(n3738), .A(n3739), .Z(n3736) );
  AND U4814 ( .A(b[18]), .B(a[34]), .Z(n3735) );
  XOR U4815 ( .A(n3740), .B(n3741), .Z(n3432) );
  AND U4816 ( .A(n3742), .B(n3743), .Z(n3740) );
  XNOR U4817 ( .A(n3744), .B(n3437), .Z(n3439) );
  XOR U4818 ( .A(n3745), .B(n3746), .Z(n3437) );
  ANDN U4819 ( .B(n3747), .A(n3748), .Z(n3745) );
  AND U4820 ( .A(b[17]), .B(a[35]), .Z(n3744) );
  XOR U4821 ( .A(n3749), .B(n3442), .Z(n3444) );
  XOR U4822 ( .A(n3750), .B(n3751), .Z(n3442) );
  ANDN U4823 ( .B(n3752), .A(n3753), .Z(n3750) );
  AND U4824 ( .A(a[37]), .B(b[15]), .Z(n3749) );
  XNOR U4825 ( .A(n3754), .B(n3447), .Z(n3449) );
  XOR U4826 ( .A(n3755), .B(n3756), .Z(n3447) );
  ANDN U4827 ( .B(n3757), .A(n3758), .Z(n3755) );
  AND U4828 ( .A(b[14]), .B(a[38]), .Z(n3754) );
  XNOR U4829 ( .A(n3759), .B(n3452), .Z(n3454) );
  XOR U4830 ( .A(n3760), .B(n3761), .Z(n3452) );
  ANDN U4831 ( .B(n3762), .A(n3763), .Z(n3760) );
  AND U4832 ( .A(b[13]), .B(a[39]), .Z(n3759) );
  XNOR U4833 ( .A(n3764), .B(n3457), .Z(n3459) );
  XOR U4834 ( .A(n3765), .B(n3766), .Z(n3457) );
  ANDN U4835 ( .B(n3767), .A(n3768), .Z(n3765) );
  AND U4836 ( .A(b[12]), .B(a[40]), .Z(n3764) );
  XNOR U4837 ( .A(n3769), .B(n3462), .Z(n3464) );
  XOR U4838 ( .A(n3770), .B(n3771), .Z(n3462) );
  ANDN U4839 ( .B(n3772), .A(n3773), .Z(n3770) );
  AND U4840 ( .A(b[11]), .B(a[41]), .Z(n3769) );
  XNOR U4841 ( .A(n3774), .B(n3467), .Z(n3469) );
  XOR U4842 ( .A(n3775), .B(n3776), .Z(n3467) );
  ANDN U4843 ( .B(n3777), .A(n3778), .Z(n3775) );
  AND U4844 ( .A(b[10]), .B(a[42]), .Z(n3774) );
  XNOR U4845 ( .A(n3779), .B(n3472), .Z(n3474) );
  XOR U4846 ( .A(n3780), .B(n3781), .Z(n3472) );
  ANDN U4847 ( .B(n3782), .A(n3783), .Z(n3780) );
  AND U4848 ( .A(b[9]), .B(a[43]), .Z(n3779) );
  XNOR U4849 ( .A(n3784), .B(n3477), .Z(n3479) );
  XOR U4850 ( .A(n3785), .B(n3786), .Z(n3477) );
  ANDN U4851 ( .B(n3787), .A(n3788), .Z(n3785) );
  AND U4852 ( .A(b[8]), .B(a[44]), .Z(n3784) );
  XNOR U4853 ( .A(n3789), .B(n3482), .Z(n3484) );
  XOR U4854 ( .A(n3790), .B(n3791), .Z(n3482) );
  ANDN U4855 ( .B(n3792), .A(n3793), .Z(n3790) );
  AND U4856 ( .A(b[7]), .B(a[45]), .Z(n3789) );
  XNOR U4857 ( .A(n3794), .B(n3487), .Z(n3489) );
  XOR U4858 ( .A(n3795), .B(n3796), .Z(n3487) );
  ANDN U4859 ( .B(n3797), .A(n3798), .Z(n3795) );
  AND U4860 ( .A(b[6]), .B(a[46]), .Z(n3794) );
  XNOR U4861 ( .A(n3799), .B(n3492), .Z(n3494) );
  XOR U4862 ( .A(n3800), .B(n3801), .Z(n3492) );
  ANDN U4863 ( .B(n3802), .A(n3803), .Z(n3800) );
  AND U4864 ( .A(b[5]), .B(a[47]), .Z(n3799) );
  XNOR U4865 ( .A(n3804), .B(n3497), .Z(n3499) );
  XOR U4866 ( .A(n3805), .B(n3806), .Z(n3497) );
  ANDN U4867 ( .B(n3807), .A(n3808), .Z(n3805) );
  AND U4868 ( .A(b[4]), .B(a[48]), .Z(n3804) );
  XNOR U4869 ( .A(n3809), .B(n3810), .Z(n3511) );
  NANDN U4870 ( .A(n3811), .B(n3812), .Z(n3810) );
  XNOR U4871 ( .A(n3813), .B(n3502), .Z(n3504) );
  XNOR U4872 ( .A(n3814), .B(n3815), .Z(n3502) );
  AND U4873 ( .A(n3816), .B(n3817), .Z(n3814) );
  AND U4874 ( .A(b[3]), .B(a[49]), .Z(n3813) );
  NAND U4875 ( .A(a[52]), .B(b[0]), .Z(n3207) );
  XNOR U4876 ( .A(n3517), .B(n3518), .Z(c[51]) );
  XNOR U4877 ( .A(n3811), .B(n3812), .Z(n3518) );
  XOR U4878 ( .A(n3809), .B(n3818), .Z(n3812) );
  NAND U4879 ( .A(b[1]), .B(a[50]), .Z(n3818) );
  XOR U4880 ( .A(n3817), .B(n3819), .Z(n3811) );
  XOR U4881 ( .A(n3809), .B(n3816), .Z(n3819) );
  XNOR U4882 ( .A(n3820), .B(n3815), .Z(n3816) );
  AND U4883 ( .A(b[2]), .B(a[49]), .Z(n3820) );
  NANDN U4884 ( .A(n3821), .B(n3822), .Z(n3809) );
  XOR U4885 ( .A(n3815), .B(n3807), .Z(n3823) );
  XNOR U4886 ( .A(n3806), .B(n3802), .Z(n3824) );
  XNOR U4887 ( .A(n3801), .B(n3797), .Z(n3825) );
  XNOR U4888 ( .A(n3796), .B(n3792), .Z(n3826) );
  XNOR U4889 ( .A(n3791), .B(n3787), .Z(n3827) );
  XNOR U4890 ( .A(n3786), .B(n3782), .Z(n3828) );
  XNOR U4891 ( .A(n3781), .B(n3777), .Z(n3829) );
  XNOR U4892 ( .A(n3776), .B(n3772), .Z(n3830) );
  XNOR U4893 ( .A(n3771), .B(n3767), .Z(n3831) );
  XNOR U4894 ( .A(n3766), .B(n3762), .Z(n3832) );
  XNOR U4895 ( .A(n3761), .B(n3757), .Z(n3833) );
  XNOR U4896 ( .A(n3756), .B(n3752), .Z(n3834) );
  XNOR U4897 ( .A(n3743), .B(n3742), .Z(n3835) );
  XOR U4898 ( .A(n3836), .B(n3741), .Z(n3742) );
  AND U4899 ( .A(b[15]), .B(a[36]), .Z(n3836) );
  XNOR U4900 ( .A(n3741), .B(n3747), .Z(n3837) );
  XNOR U4901 ( .A(n3746), .B(n3738), .Z(n3838) );
  XNOR U4902 ( .A(n3737), .B(n3733), .Z(n3839) );
  XNOR U4903 ( .A(n3732), .B(n3728), .Z(n3840) );
  XNOR U4904 ( .A(n3727), .B(n3723), .Z(n3841) );
  XNOR U4905 ( .A(n3842), .B(n3843), .Z(n3723) );
  XNOR U4906 ( .A(n3714), .B(n3713), .Z(n3843) );
  XOR U4907 ( .A(n3844), .B(n3712), .Z(n3713) );
  AND U4908 ( .A(b[21]), .B(a[30]), .Z(n3844) );
  XNOR U4909 ( .A(n3712), .B(n3718), .Z(n3845) );
  XNOR U4910 ( .A(n3717), .B(n3709), .Z(n3846) );
  XNOR U4911 ( .A(n3708), .B(n3704), .Z(n3847) );
  XNOR U4912 ( .A(n3703), .B(n3699), .Z(n3848) );
  XNOR U4913 ( .A(n3698), .B(n3694), .Z(n3849) );
  XNOR U4914 ( .A(n3685), .B(n3684), .Z(n3850) );
  XOR U4915 ( .A(n3851), .B(n3683), .Z(n3684) );
  AND U4916 ( .A(b[27]), .B(a[24]), .Z(n3851) );
  XNOR U4917 ( .A(n3683), .B(n3689), .Z(n3852) );
  XNOR U4918 ( .A(n3688), .B(n3680), .Z(n3853) );
  XNOR U4919 ( .A(n3679), .B(n3675), .Z(n3854) );
  XNOR U4920 ( .A(n3674), .B(n3670), .Z(n3855) );
  XNOR U4921 ( .A(n3669), .B(n3665), .Z(n3856) );
  XNOR U4922 ( .A(n3656), .B(n3655), .Z(n3857) );
  XOR U4923 ( .A(n3858), .B(n3654), .Z(n3655) );
  AND U4924 ( .A(b[33]), .B(a[18]), .Z(n3858) );
  XNOR U4925 ( .A(n3654), .B(n3660), .Z(n3859) );
  XNOR U4926 ( .A(n3659), .B(n3651), .Z(n3860) );
  XNOR U4927 ( .A(n3650), .B(n3646), .Z(n3861) );
  XNOR U4928 ( .A(n3645), .B(n3641), .Z(n3862) );
  XNOR U4929 ( .A(n3640), .B(n3636), .Z(n3863) );
  XNOR U4930 ( .A(n3627), .B(n3626), .Z(n3864) );
  XOR U4931 ( .A(n3865), .B(n3625), .Z(n3626) );
  AND U4932 ( .A(b[39]), .B(a[12]), .Z(n3865) );
  XNOR U4933 ( .A(n3625), .B(n3631), .Z(n3866) );
  XNOR U4934 ( .A(n3630), .B(n3622), .Z(n3867) );
  XNOR U4935 ( .A(n3621), .B(n3617), .Z(n3868) );
  XNOR U4936 ( .A(n3616), .B(n3612), .Z(n3869) );
  XNOR U4937 ( .A(n3611), .B(n3607), .Z(n3870) );
  XNOR U4938 ( .A(n3598), .B(n3597), .Z(n3871) );
  XOR U4939 ( .A(n3872), .B(n3596), .Z(n3597) );
  AND U4940 ( .A(a[6]), .B(b[45]), .Z(n3872) );
  XNOR U4941 ( .A(n3596), .B(n3602), .Z(n3873) );
  XNOR U4942 ( .A(n3601), .B(n3593), .Z(n3874) );
  XNOR U4943 ( .A(n3592), .B(n3588), .Z(n3875) );
  XNOR U4944 ( .A(n3587), .B(n3583), .Z(n3876) );
  XNOR U4945 ( .A(n3582), .B(n3578), .Z(n3877) );
  XNOR U4946 ( .A(n3878), .B(n3577), .Z(n3578) );
  AND U4947 ( .A(a[0]), .B(b[51]), .Z(n3878) );
  XOR U4948 ( .A(n3879), .B(n3577), .Z(n3579) );
  XNOR U4949 ( .A(n3880), .B(n3881), .Z(n3577) );
  ANDN U4950 ( .B(n3882), .A(n3883), .Z(n3880) );
  AND U4951 ( .A(a[1]), .B(b[50]), .Z(n3879) );
  XNOR U4952 ( .A(n3884), .B(n3582), .Z(n3584) );
  XOR U4953 ( .A(n3885), .B(n3886), .Z(n3582) );
  ANDN U4954 ( .B(n3887), .A(n3888), .Z(n3885) );
  AND U4955 ( .A(a[2]), .B(b[49]), .Z(n3884) );
  XNOR U4956 ( .A(n3889), .B(n3587), .Z(n3589) );
  XOR U4957 ( .A(n3890), .B(n3891), .Z(n3587) );
  ANDN U4958 ( .B(n3892), .A(n3893), .Z(n3890) );
  AND U4959 ( .A(a[3]), .B(b[48]), .Z(n3889) );
  XNOR U4960 ( .A(n3894), .B(n3592), .Z(n3594) );
  XOR U4961 ( .A(n3895), .B(n3896), .Z(n3592) );
  ANDN U4962 ( .B(n3897), .A(n3898), .Z(n3895) );
  AND U4963 ( .A(a[4]), .B(b[47]), .Z(n3894) );
  XOR U4964 ( .A(n3899), .B(n3900), .Z(n3596) );
  AND U4965 ( .A(n3901), .B(n3902), .Z(n3899) );
  XNOR U4966 ( .A(n3903), .B(n3601), .Z(n3603) );
  XOR U4967 ( .A(n3904), .B(n3905), .Z(n3601) );
  ANDN U4968 ( .B(n3906), .A(n3907), .Z(n3904) );
  AND U4969 ( .A(a[5]), .B(b[46]), .Z(n3903) );
  XOR U4970 ( .A(n3908), .B(n3606), .Z(n3608) );
  XOR U4971 ( .A(n3909), .B(n3910), .Z(n3606) );
  ANDN U4972 ( .B(n3911), .A(n3912), .Z(n3909) );
  AND U4973 ( .A(a[7]), .B(b[44]), .Z(n3908) );
  XNOR U4974 ( .A(n3913), .B(n3611), .Z(n3613) );
  XOR U4975 ( .A(n3914), .B(n3915), .Z(n3611) );
  ANDN U4976 ( .B(n3916), .A(n3917), .Z(n3914) );
  AND U4977 ( .A(a[8]), .B(b[43]), .Z(n3913) );
  XNOR U4978 ( .A(n3918), .B(n3616), .Z(n3618) );
  XOR U4979 ( .A(n3919), .B(n3920), .Z(n3616) );
  ANDN U4980 ( .B(n3921), .A(n3922), .Z(n3919) );
  AND U4981 ( .A(a[9]), .B(b[42]), .Z(n3918) );
  XNOR U4982 ( .A(n3923), .B(n3621), .Z(n3623) );
  XOR U4983 ( .A(n3924), .B(n3925), .Z(n3621) );
  ANDN U4984 ( .B(n3926), .A(n3927), .Z(n3924) );
  AND U4985 ( .A(b[41]), .B(a[10]), .Z(n3923) );
  XOR U4986 ( .A(n3928), .B(n3929), .Z(n3625) );
  AND U4987 ( .A(n3930), .B(n3931), .Z(n3928) );
  XNOR U4988 ( .A(n3932), .B(n3630), .Z(n3632) );
  XOR U4989 ( .A(n3933), .B(n3934), .Z(n3630) );
  ANDN U4990 ( .B(n3935), .A(n3936), .Z(n3933) );
  AND U4991 ( .A(b[40]), .B(a[11]), .Z(n3932) );
  XOR U4992 ( .A(n3937), .B(n3635), .Z(n3637) );
  XOR U4993 ( .A(n3938), .B(n3939), .Z(n3635) );
  ANDN U4994 ( .B(n3940), .A(n3941), .Z(n3938) );
  AND U4995 ( .A(b[38]), .B(a[13]), .Z(n3937) );
  XNOR U4996 ( .A(n3942), .B(n3640), .Z(n3642) );
  XOR U4997 ( .A(n3943), .B(n3944), .Z(n3640) );
  ANDN U4998 ( .B(n3945), .A(n3946), .Z(n3943) );
  AND U4999 ( .A(b[37]), .B(a[14]), .Z(n3942) );
  XNOR U5000 ( .A(n3947), .B(n3645), .Z(n3647) );
  XOR U5001 ( .A(n3948), .B(n3949), .Z(n3645) );
  ANDN U5002 ( .B(n3950), .A(n3951), .Z(n3948) );
  AND U5003 ( .A(b[36]), .B(a[15]), .Z(n3947) );
  XNOR U5004 ( .A(n3952), .B(n3650), .Z(n3652) );
  XOR U5005 ( .A(n3953), .B(n3954), .Z(n3650) );
  ANDN U5006 ( .B(n3955), .A(n3956), .Z(n3953) );
  AND U5007 ( .A(b[35]), .B(a[16]), .Z(n3952) );
  XOR U5008 ( .A(n3957), .B(n3958), .Z(n3654) );
  AND U5009 ( .A(n3959), .B(n3960), .Z(n3957) );
  XNOR U5010 ( .A(n3961), .B(n3659), .Z(n3661) );
  XOR U5011 ( .A(n3962), .B(n3963), .Z(n3659) );
  ANDN U5012 ( .B(n3964), .A(n3965), .Z(n3962) );
  AND U5013 ( .A(b[34]), .B(a[17]), .Z(n3961) );
  XOR U5014 ( .A(n3966), .B(n3664), .Z(n3666) );
  XOR U5015 ( .A(n3967), .B(n3968), .Z(n3664) );
  ANDN U5016 ( .B(n3969), .A(n3970), .Z(n3967) );
  AND U5017 ( .A(b[32]), .B(a[19]), .Z(n3966) );
  XNOR U5018 ( .A(n3971), .B(n3669), .Z(n3671) );
  XOR U5019 ( .A(n3972), .B(n3973), .Z(n3669) );
  ANDN U5020 ( .B(n3974), .A(n3975), .Z(n3972) );
  AND U5021 ( .A(b[31]), .B(a[20]), .Z(n3971) );
  XNOR U5022 ( .A(n3976), .B(n3674), .Z(n3676) );
  XOR U5023 ( .A(n3977), .B(n3978), .Z(n3674) );
  ANDN U5024 ( .B(n3979), .A(n3980), .Z(n3977) );
  AND U5025 ( .A(b[30]), .B(a[21]), .Z(n3976) );
  XNOR U5026 ( .A(n3981), .B(n3679), .Z(n3681) );
  XOR U5027 ( .A(n3982), .B(n3983), .Z(n3679) );
  ANDN U5028 ( .B(n3984), .A(n3985), .Z(n3982) );
  AND U5029 ( .A(b[29]), .B(a[22]), .Z(n3981) );
  XOR U5030 ( .A(n3986), .B(n3987), .Z(n3683) );
  AND U5031 ( .A(n3988), .B(n3989), .Z(n3986) );
  XNOR U5032 ( .A(n3990), .B(n3688), .Z(n3690) );
  XOR U5033 ( .A(n3991), .B(n3992), .Z(n3688) );
  ANDN U5034 ( .B(n3993), .A(n3994), .Z(n3991) );
  AND U5035 ( .A(b[28]), .B(a[23]), .Z(n3990) );
  XOR U5036 ( .A(n3995), .B(n3693), .Z(n3695) );
  XOR U5037 ( .A(n3996), .B(n3997), .Z(n3693) );
  ANDN U5038 ( .B(n3998), .A(n3999), .Z(n3996) );
  AND U5039 ( .A(b[26]), .B(a[25]), .Z(n3995) );
  XNOR U5040 ( .A(n4000), .B(n3698), .Z(n3700) );
  XOR U5041 ( .A(n4001), .B(n4002), .Z(n3698) );
  ANDN U5042 ( .B(n4003), .A(n4004), .Z(n4001) );
  AND U5043 ( .A(b[25]), .B(a[26]), .Z(n4000) );
  XNOR U5044 ( .A(n4005), .B(n3703), .Z(n3705) );
  XOR U5045 ( .A(n4006), .B(n4007), .Z(n3703) );
  ANDN U5046 ( .B(n4008), .A(n4009), .Z(n4006) );
  AND U5047 ( .A(b[24]), .B(a[27]), .Z(n4005) );
  XNOR U5048 ( .A(n4010), .B(n3708), .Z(n3710) );
  XOR U5049 ( .A(n4011), .B(n4012), .Z(n3708) );
  ANDN U5050 ( .B(n4013), .A(n4014), .Z(n4011) );
  AND U5051 ( .A(b[23]), .B(a[28]), .Z(n4010) );
  XOR U5052 ( .A(n4015), .B(n4016), .Z(n3712) );
  AND U5053 ( .A(n4017), .B(n4018), .Z(n4015) );
  XNOR U5054 ( .A(n4019), .B(n3717), .Z(n3719) );
  XOR U5055 ( .A(n4020), .B(n4021), .Z(n3717) );
  ANDN U5056 ( .B(n4022), .A(n4023), .Z(n4020) );
  AND U5057 ( .A(b[22]), .B(a[29]), .Z(n4019) );
  IV U5058 ( .A(n3722), .Z(n3842) );
  XOR U5059 ( .A(n4024), .B(n3722), .Z(n3724) );
  XOR U5060 ( .A(n4025), .B(n4026), .Z(n3722) );
  ANDN U5061 ( .B(n4027), .A(n4028), .Z(n4025) );
  AND U5062 ( .A(b[20]), .B(a[31]), .Z(n4024) );
  XNOR U5063 ( .A(n4029), .B(n3727), .Z(n3729) );
  XOR U5064 ( .A(n4030), .B(n4031), .Z(n3727) );
  ANDN U5065 ( .B(n4032), .A(n4033), .Z(n4030) );
  AND U5066 ( .A(b[19]), .B(a[32]), .Z(n4029) );
  XNOR U5067 ( .A(n4034), .B(n3732), .Z(n3734) );
  XOR U5068 ( .A(n4035), .B(n4036), .Z(n3732) );
  ANDN U5069 ( .B(n4037), .A(n4038), .Z(n4035) );
  AND U5070 ( .A(b[18]), .B(a[33]), .Z(n4034) );
  XNOR U5071 ( .A(n4039), .B(n3737), .Z(n3739) );
  XOR U5072 ( .A(n4040), .B(n4041), .Z(n3737) );
  ANDN U5073 ( .B(n4042), .A(n4043), .Z(n4040) );
  AND U5074 ( .A(b[17]), .B(a[34]), .Z(n4039) );
  XOR U5075 ( .A(n4044), .B(n4045), .Z(n3741) );
  AND U5076 ( .A(n4046), .B(n4047), .Z(n4044) );
  XNOR U5077 ( .A(n4048), .B(n3746), .Z(n3748) );
  XOR U5078 ( .A(n4049), .B(n4050), .Z(n3746) );
  ANDN U5079 ( .B(n4051), .A(n4052), .Z(n4049) );
  AND U5080 ( .A(b[16]), .B(a[35]), .Z(n4048) );
  XOR U5081 ( .A(n4053), .B(n3751), .Z(n3753) );
  XOR U5082 ( .A(n4054), .B(n4055), .Z(n3751) );
  ANDN U5083 ( .B(n4056), .A(n4057), .Z(n4054) );
  AND U5084 ( .A(b[14]), .B(a[37]), .Z(n4053) );
  XNOR U5085 ( .A(n4058), .B(n3756), .Z(n3758) );
  XOR U5086 ( .A(n4059), .B(n4060), .Z(n3756) );
  ANDN U5087 ( .B(n4061), .A(n4062), .Z(n4059) );
  AND U5088 ( .A(b[13]), .B(a[38]), .Z(n4058) );
  XNOR U5089 ( .A(n4063), .B(n3761), .Z(n3763) );
  XOR U5090 ( .A(n4064), .B(n4065), .Z(n3761) );
  ANDN U5091 ( .B(n4066), .A(n4067), .Z(n4064) );
  AND U5092 ( .A(b[12]), .B(a[39]), .Z(n4063) );
  XNOR U5093 ( .A(n4068), .B(n3766), .Z(n3768) );
  XOR U5094 ( .A(n4069), .B(n4070), .Z(n3766) );
  ANDN U5095 ( .B(n4071), .A(n4072), .Z(n4069) );
  AND U5096 ( .A(b[11]), .B(a[40]), .Z(n4068) );
  XNOR U5097 ( .A(n4073), .B(n3771), .Z(n3773) );
  XOR U5098 ( .A(n4074), .B(n4075), .Z(n3771) );
  ANDN U5099 ( .B(n4076), .A(n4077), .Z(n4074) );
  AND U5100 ( .A(b[10]), .B(a[41]), .Z(n4073) );
  XNOR U5101 ( .A(n4078), .B(n3776), .Z(n3778) );
  XOR U5102 ( .A(n4079), .B(n4080), .Z(n3776) );
  ANDN U5103 ( .B(n4081), .A(n4082), .Z(n4079) );
  AND U5104 ( .A(b[9]), .B(a[42]), .Z(n4078) );
  XNOR U5105 ( .A(n4083), .B(n3781), .Z(n3783) );
  XOR U5106 ( .A(n4084), .B(n4085), .Z(n3781) );
  ANDN U5107 ( .B(n4086), .A(n4087), .Z(n4084) );
  AND U5108 ( .A(b[8]), .B(a[43]), .Z(n4083) );
  XNOR U5109 ( .A(n4088), .B(n3786), .Z(n3788) );
  XOR U5110 ( .A(n4089), .B(n4090), .Z(n3786) );
  ANDN U5111 ( .B(n4091), .A(n4092), .Z(n4089) );
  AND U5112 ( .A(b[7]), .B(a[44]), .Z(n4088) );
  XNOR U5113 ( .A(n4093), .B(n3791), .Z(n3793) );
  XOR U5114 ( .A(n4094), .B(n4095), .Z(n3791) );
  ANDN U5115 ( .B(n4096), .A(n4097), .Z(n4094) );
  AND U5116 ( .A(b[6]), .B(a[45]), .Z(n4093) );
  XNOR U5117 ( .A(n4098), .B(n3796), .Z(n3798) );
  XOR U5118 ( .A(n4099), .B(n4100), .Z(n3796) );
  ANDN U5119 ( .B(n4101), .A(n4102), .Z(n4099) );
  AND U5120 ( .A(b[5]), .B(a[46]), .Z(n4098) );
  XNOR U5121 ( .A(n4103), .B(n3801), .Z(n3803) );
  XOR U5122 ( .A(n4104), .B(n4105), .Z(n3801) );
  ANDN U5123 ( .B(n4106), .A(n4107), .Z(n4104) );
  AND U5124 ( .A(b[4]), .B(a[47]), .Z(n4103) );
  XNOR U5125 ( .A(n4108), .B(n4109), .Z(n3815) );
  NANDN U5126 ( .A(n4110), .B(n4111), .Z(n4109) );
  XNOR U5127 ( .A(n4112), .B(n3806), .Z(n3808) );
  XNOR U5128 ( .A(n4113), .B(n4114), .Z(n3806) );
  AND U5129 ( .A(n4115), .B(n4116), .Z(n4113) );
  AND U5130 ( .A(b[3]), .B(a[48]), .Z(n4112) );
  NAND U5131 ( .A(a[51]), .B(b[0]), .Z(n3517) );
  XNOR U5132 ( .A(n3821), .B(n3822), .Z(c[50]) );
  XNOR U5133 ( .A(n4110), .B(n4111), .Z(n3822) );
  XOR U5134 ( .A(n4108), .B(n4117), .Z(n4111) );
  NAND U5135 ( .A(b[1]), .B(a[49]), .Z(n4117) );
  XOR U5136 ( .A(n4115), .B(n4118), .Z(n4110) );
  XOR U5137 ( .A(n4108), .B(n4116), .Z(n4118) );
  XNOR U5138 ( .A(n4119), .B(n4114), .Z(n4116) );
  AND U5139 ( .A(b[2]), .B(a[48]), .Z(n4119) );
  NANDN U5140 ( .A(n4120), .B(n4121), .Z(n4108) );
  XOR U5141 ( .A(n4114), .B(n4106), .Z(n4122) );
  XNOR U5142 ( .A(n4105), .B(n4101), .Z(n4123) );
  XNOR U5143 ( .A(n4100), .B(n4096), .Z(n4124) );
  XNOR U5144 ( .A(n4095), .B(n4091), .Z(n4125) );
  XNOR U5145 ( .A(n4090), .B(n4086), .Z(n4126) );
  XNOR U5146 ( .A(n4085), .B(n4081), .Z(n4127) );
  XNOR U5147 ( .A(n4080), .B(n4076), .Z(n4128) );
  XNOR U5148 ( .A(n4075), .B(n4071), .Z(n4129) );
  XNOR U5149 ( .A(n4070), .B(n4066), .Z(n4130) );
  XNOR U5150 ( .A(n4065), .B(n4061), .Z(n4131) );
  XNOR U5151 ( .A(n4060), .B(n4056), .Z(n4132) );
  XNOR U5152 ( .A(n4047), .B(n4046), .Z(n4133) );
  XOR U5153 ( .A(n4134), .B(n4045), .Z(n4046) );
  AND U5154 ( .A(b[14]), .B(a[36]), .Z(n4134) );
  XNOR U5155 ( .A(n4045), .B(n4051), .Z(n4135) );
  XNOR U5156 ( .A(n4050), .B(n4042), .Z(n4136) );
  XNOR U5157 ( .A(n4041), .B(n4037), .Z(n4137) );
  XNOR U5158 ( .A(n4036), .B(n4032), .Z(n4138) );
  XNOR U5159 ( .A(n4031), .B(n4027), .Z(n4139) );
  XNOR U5160 ( .A(n4018), .B(n4017), .Z(n4140) );
  XOR U5161 ( .A(n4141), .B(n4016), .Z(n4017) );
  AND U5162 ( .A(b[20]), .B(a[30]), .Z(n4141) );
  XNOR U5163 ( .A(n4016), .B(n4022), .Z(n4142) );
  XNOR U5164 ( .A(n4021), .B(n4013), .Z(n4143) );
  XNOR U5165 ( .A(n4012), .B(n4008), .Z(n4144) );
  XNOR U5166 ( .A(n4007), .B(n4003), .Z(n4145) );
  XNOR U5167 ( .A(n4002), .B(n3998), .Z(n4146) );
  XNOR U5168 ( .A(n3989), .B(n3988), .Z(n4147) );
  XOR U5169 ( .A(n4148), .B(n3987), .Z(n3988) );
  AND U5170 ( .A(b[26]), .B(a[24]), .Z(n4148) );
  XNOR U5171 ( .A(n3987), .B(n3993), .Z(n4149) );
  XNOR U5172 ( .A(n3992), .B(n3984), .Z(n4150) );
  XNOR U5173 ( .A(n3983), .B(n3979), .Z(n4151) );
  XNOR U5174 ( .A(n3978), .B(n3974), .Z(n4152) );
  XNOR U5175 ( .A(n3973), .B(n3969), .Z(n4153) );
  XNOR U5176 ( .A(n3960), .B(n3959), .Z(n4154) );
  XOR U5177 ( .A(n4155), .B(n3958), .Z(n3959) );
  AND U5178 ( .A(b[32]), .B(a[18]), .Z(n4155) );
  XNOR U5179 ( .A(n3958), .B(n3964), .Z(n4156) );
  XNOR U5180 ( .A(n3963), .B(n3955), .Z(n4157) );
  XNOR U5181 ( .A(n3954), .B(n3950), .Z(n4158) );
  XNOR U5182 ( .A(n3949), .B(n3945), .Z(n4159) );
  XNOR U5183 ( .A(n3944), .B(n3940), .Z(n4160) );
  XNOR U5184 ( .A(n3931), .B(n3930), .Z(n4161) );
  XOR U5185 ( .A(n4162), .B(n3929), .Z(n3930) );
  AND U5186 ( .A(b[38]), .B(a[12]), .Z(n4162) );
  XNOR U5187 ( .A(n3929), .B(n3935), .Z(n4163) );
  XNOR U5188 ( .A(n3934), .B(n3926), .Z(n4164) );
  XNOR U5189 ( .A(n3925), .B(n3921), .Z(n4165) );
  XNOR U5190 ( .A(n3920), .B(n3916), .Z(n4166) );
  XNOR U5191 ( .A(n3915), .B(n3911), .Z(n4167) );
  XNOR U5192 ( .A(n3902), .B(n3901), .Z(n4168) );
  XOR U5193 ( .A(n4169), .B(n3900), .Z(n3901) );
  AND U5194 ( .A(a[6]), .B(b[44]), .Z(n4169) );
  XNOR U5195 ( .A(n3900), .B(n3906), .Z(n4170) );
  XNOR U5196 ( .A(n3905), .B(n3897), .Z(n4171) );
  XNOR U5197 ( .A(n3896), .B(n3892), .Z(n4172) );
  XNOR U5198 ( .A(n3891), .B(n3887), .Z(n4173) );
  XNOR U5199 ( .A(n3886), .B(n3882), .Z(n4174) );
  XOR U5200 ( .A(n4175), .B(n3881), .Z(n3882) );
  AND U5201 ( .A(a[0]), .B(b[50]), .Z(n4175) );
  XNOR U5202 ( .A(n4176), .B(n3881), .Z(n3883) );
  XNOR U5203 ( .A(n4177), .B(n4178), .Z(n3881) );
  ANDN U5204 ( .B(n4179), .A(n4180), .Z(n4177) );
  AND U5205 ( .A(a[1]), .B(b[49]), .Z(n4176) );
  XNOR U5206 ( .A(n4181), .B(n3886), .Z(n3888) );
  XOR U5207 ( .A(n4182), .B(n4183), .Z(n3886) );
  ANDN U5208 ( .B(n4184), .A(n4185), .Z(n4182) );
  AND U5209 ( .A(a[2]), .B(b[48]), .Z(n4181) );
  XNOR U5210 ( .A(n4186), .B(n3891), .Z(n3893) );
  XOR U5211 ( .A(n4187), .B(n4188), .Z(n3891) );
  ANDN U5212 ( .B(n4189), .A(n4190), .Z(n4187) );
  AND U5213 ( .A(a[3]), .B(b[47]), .Z(n4186) );
  XNOR U5214 ( .A(n4191), .B(n3896), .Z(n3898) );
  XOR U5215 ( .A(n4192), .B(n4193), .Z(n3896) );
  ANDN U5216 ( .B(n4194), .A(n4195), .Z(n4192) );
  AND U5217 ( .A(a[4]), .B(b[46]), .Z(n4191) );
  XOR U5218 ( .A(n4196), .B(n4197), .Z(n3900) );
  AND U5219 ( .A(n4198), .B(n4199), .Z(n4196) );
  XNOR U5220 ( .A(n4200), .B(n3905), .Z(n3907) );
  XOR U5221 ( .A(n4201), .B(n4202), .Z(n3905) );
  ANDN U5222 ( .B(n4203), .A(n4204), .Z(n4201) );
  AND U5223 ( .A(a[5]), .B(b[45]), .Z(n4200) );
  XOR U5224 ( .A(n4205), .B(n3910), .Z(n3912) );
  XOR U5225 ( .A(n4206), .B(n4207), .Z(n3910) );
  ANDN U5226 ( .B(n4208), .A(n4209), .Z(n4206) );
  AND U5227 ( .A(a[7]), .B(b[43]), .Z(n4205) );
  XNOR U5228 ( .A(n4210), .B(n3915), .Z(n3917) );
  XOR U5229 ( .A(n4211), .B(n4212), .Z(n3915) );
  ANDN U5230 ( .B(n4213), .A(n4214), .Z(n4211) );
  AND U5231 ( .A(a[8]), .B(b[42]), .Z(n4210) );
  XNOR U5232 ( .A(n4215), .B(n3920), .Z(n3922) );
  XOR U5233 ( .A(n4216), .B(n4217), .Z(n3920) );
  ANDN U5234 ( .B(n4218), .A(n4219), .Z(n4216) );
  AND U5235 ( .A(a[9]), .B(b[41]), .Z(n4215) );
  XNOR U5236 ( .A(n4220), .B(n3925), .Z(n3927) );
  XOR U5237 ( .A(n4221), .B(n4222), .Z(n3925) );
  ANDN U5238 ( .B(n4223), .A(n4224), .Z(n4221) );
  AND U5239 ( .A(b[40]), .B(a[10]), .Z(n4220) );
  XOR U5240 ( .A(n4225), .B(n4226), .Z(n3929) );
  AND U5241 ( .A(n4227), .B(n4228), .Z(n4225) );
  XNOR U5242 ( .A(n4229), .B(n3934), .Z(n3936) );
  XOR U5243 ( .A(n4230), .B(n4231), .Z(n3934) );
  ANDN U5244 ( .B(n4232), .A(n4233), .Z(n4230) );
  AND U5245 ( .A(a[11]), .B(b[39]), .Z(n4229) );
  XOR U5246 ( .A(n4234), .B(n3939), .Z(n3941) );
  XOR U5247 ( .A(n4235), .B(n4236), .Z(n3939) );
  ANDN U5248 ( .B(n4237), .A(n4238), .Z(n4235) );
  AND U5249 ( .A(b[37]), .B(a[13]), .Z(n4234) );
  XNOR U5250 ( .A(n4239), .B(n3944), .Z(n3946) );
  XOR U5251 ( .A(n4240), .B(n4241), .Z(n3944) );
  ANDN U5252 ( .B(n4242), .A(n4243), .Z(n4240) );
  AND U5253 ( .A(b[36]), .B(a[14]), .Z(n4239) );
  XNOR U5254 ( .A(n4244), .B(n3949), .Z(n3951) );
  XOR U5255 ( .A(n4245), .B(n4246), .Z(n3949) );
  ANDN U5256 ( .B(n4247), .A(n4248), .Z(n4245) );
  AND U5257 ( .A(b[35]), .B(a[15]), .Z(n4244) );
  XNOR U5258 ( .A(n4249), .B(n3954), .Z(n3956) );
  XOR U5259 ( .A(n4250), .B(n4251), .Z(n3954) );
  ANDN U5260 ( .B(n4252), .A(n4253), .Z(n4250) );
  AND U5261 ( .A(b[34]), .B(a[16]), .Z(n4249) );
  XOR U5262 ( .A(n4254), .B(n4255), .Z(n3958) );
  AND U5263 ( .A(n4256), .B(n4257), .Z(n4254) );
  XNOR U5264 ( .A(n4258), .B(n3963), .Z(n3965) );
  XOR U5265 ( .A(n4259), .B(n4260), .Z(n3963) );
  ANDN U5266 ( .B(n4261), .A(n4262), .Z(n4259) );
  AND U5267 ( .A(a[17]), .B(b[33]), .Z(n4258) );
  XOR U5268 ( .A(n4263), .B(n3968), .Z(n3970) );
  XOR U5269 ( .A(n4264), .B(n4265), .Z(n3968) );
  ANDN U5270 ( .B(n4266), .A(n4267), .Z(n4264) );
  AND U5271 ( .A(b[31]), .B(a[19]), .Z(n4263) );
  XNOR U5272 ( .A(n4268), .B(n3973), .Z(n3975) );
  XOR U5273 ( .A(n4269), .B(n4270), .Z(n3973) );
  ANDN U5274 ( .B(n4271), .A(n4272), .Z(n4269) );
  AND U5275 ( .A(b[30]), .B(a[20]), .Z(n4268) );
  XNOR U5276 ( .A(n4273), .B(n3978), .Z(n3980) );
  XOR U5277 ( .A(n4274), .B(n4275), .Z(n3978) );
  ANDN U5278 ( .B(n4276), .A(n4277), .Z(n4274) );
  AND U5279 ( .A(b[29]), .B(a[21]), .Z(n4273) );
  XNOR U5280 ( .A(n4278), .B(n3983), .Z(n3985) );
  XOR U5281 ( .A(n4279), .B(n4280), .Z(n3983) );
  ANDN U5282 ( .B(n4281), .A(n4282), .Z(n4279) );
  AND U5283 ( .A(b[28]), .B(a[22]), .Z(n4278) );
  XOR U5284 ( .A(n4283), .B(n4284), .Z(n3987) );
  AND U5285 ( .A(n4285), .B(n4286), .Z(n4283) );
  XNOR U5286 ( .A(n4287), .B(n3992), .Z(n3994) );
  XOR U5287 ( .A(n4288), .B(n4289), .Z(n3992) );
  ANDN U5288 ( .B(n4290), .A(n4291), .Z(n4288) );
  AND U5289 ( .A(a[23]), .B(b[27]), .Z(n4287) );
  XOR U5290 ( .A(n4292), .B(n3997), .Z(n3999) );
  XOR U5291 ( .A(n4293), .B(n4294), .Z(n3997) );
  ANDN U5292 ( .B(n4295), .A(n4296), .Z(n4293) );
  AND U5293 ( .A(b[25]), .B(a[25]), .Z(n4292) );
  XNOR U5294 ( .A(n4297), .B(n4002), .Z(n4004) );
  XOR U5295 ( .A(n4298), .B(n4299), .Z(n4002) );
  ANDN U5296 ( .B(n4300), .A(n4301), .Z(n4298) );
  AND U5297 ( .A(b[24]), .B(a[26]), .Z(n4297) );
  XNOR U5298 ( .A(n4302), .B(n4007), .Z(n4009) );
  XOR U5299 ( .A(n4303), .B(n4304), .Z(n4007) );
  ANDN U5300 ( .B(n4305), .A(n4306), .Z(n4303) );
  AND U5301 ( .A(b[23]), .B(a[27]), .Z(n4302) );
  XNOR U5302 ( .A(n4307), .B(n4012), .Z(n4014) );
  XOR U5303 ( .A(n4308), .B(n4309), .Z(n4012) );
  ANDN U5304 ( .B(n4310), .A(n4311), .Z(n4308) );
  AND U5305 ( .A(b[22]), .B(a[28]), .Z(n4307) );
  XOR U5306 ( .A(n4312), .B(n4313), .Z(n4016) );
  AND U5307 ( .A(n4314), .B(n4315), .Z(n4312) );
  XNOR U5308 ( .A(n4316), .B(n4021), .Z(n4023) );
  XOR U5309 ( .A(n4317), .B(n4318), .Z(n4021) );
  ANDN U5310 ( .B(n4319), .A(n4320), .Z(n4317) );
  AND U5311 ( .A(a[29]), .B(b[21]), .Z(n4316) );
  XOR U5312 ( .A(n4321), .B(n4026), .Z(n4028) );
  XOR U5313 ( .A(n4322), .B(n4323), .Z(n4026) );
  ANDN U5314 ( .B(n4324), .A(n4325), .Z(n4322) );
  AND U5315 ( .A(b[19]), .B(a[31]), .Z(n4321) );
  XNOR U5316 ( .A(n4326), .B(n4031), .Z(n4033) );
  XOR U5317 ( .A(n4327), .B(n4328), .Z(n4031) );
  ANDN U5318 ( .B(n4329), .A(n4330), .Z(n4327) );
  AND U5319 ( .A(b[18]), .B(a[32]), .Z(n4326) );
  XNOR U5320 ( .A(n4331), .B(n4036), .Z(n4038) );
  XOR U5321 ( .A(n4332), .B(n4333), .Z(n4036) );
  ANDN U5322 ( .B(n4334), .A(n4335), .Z(n4332) );
  AND U5323 ( .A(b[17]), .B(a[33]), .Z(n4331) );
  XNOR U5324 ( .A(n4336), .B(n4041), .Z(n4043) );
  XOR U5325 ( .A(n4337), .B(n4338), .Z(n4041) );
  ANDN U5326 ( .B(n4339), .A(n4340), .Z(n4337) );
  AND U5327 ( .A(b[16]), .B(a[34]), .Z(n4336) );
  XOR U5328 ( .A(n4341), .B(n4342), .Z(n4045) );
  AND U5329 ( .A(n4343), .B(n4344), .Z(n4341) );
  XNOR U5330 ( .A(n4345), .B(n4050), .Z(n4052) );
  XOR U5331 ( .A(n4346), .B(n4347), .Z(n4050) );
  ANDN U5332 ( .B(n4348), .A(n4349), .Z(n4346) );
  AND U5333 ( .A(a[35]), .B(b[15]), .Z(n4345) );
  XOR U5334 ( .A(n4350), .B(n4055), .Z(n4057) );
  XOR U5335 ( .A(n4351), .B(n4352), .Z(n4055) );
  ANDN U5336 ( .B(n4353), .A(n4354), .Z(n4351) );
  AND U5337 ( .A(b[13]), .B(a[37]), .Z(n4350) );
  XNOR U5338 ( .A(n4355), .B(n4060), .Z(n4062) );
  XOR U5339 ( .A(n4356), .B(n4357), .Z(n4060) );
  ANDN U5340 ( .B(n4358), .A(n4359), .Z(n4356) );
  AND U5341 ( .A(b[12]), .B(a[38]), .Z(n4355) );
  XNOR U5342 ( .A(n4360), .B(n4065), .Z(n4067) );
  XOR U5343 ( .A(n4361), .B(n4362), .Z(n4065) );
  ANDN U5344 ( .B(n4363), .A(n4364), .Z(n4361) );
  AND U5345 ( .A(b[11]), .B(a[39]), .Z(n4360) );
  XNOR U5346 ( .A(n4365), .B(n4070), .Z(n4072) );
  XOR U5347 ( .A(n4366), .B(n4367), .Z(n4070) );
  ANDN U5348 ( .B(n4368), .A(n4369), .Z(n4366) );
  AND U5349 ( .A(b[10]), .B(a[40]), .Z(n4365) );
  XNOR U5350 ( .A(n4370), .B(n4075), .Z(n4077) );
  XOR U5351 ( .A(n4371), .B(n4372), .Z(n4075) );
  ANDN U5352 ( .B(n4373), .A(n4374), .Z(n4371) );
  AND U5353 ( .A(b[9]), .B(a[41]), .Z(n4370) );
  XNOR U5354 ( .A(n4375), .B(n4080), .Z(n4082) );
  XOR U5355 ( .A(n4376), .B(n4377), .Z(n4080) );
  ANDN U5356 ( .B(n4378), .A(n4379), .Z(n4376) );
  AND U5357 ( .A(b[8]), .B(a[42]), .Z(n4375) );
  XNOR U5358 ( .A(n4380), .B(n4085), .Z(n4087) );
  XOR U5359 ( .A(n4381), .B(n4382), .Z(n4085) );
  ANDN U5360 ( .B(n4383), .A(n4384), .Z(n4381) );
  AND U5361 ( .A(b[7]), .B(a[43]), .Z(n4380) );
  XNOR U5362 ( .A(n4385), .B(n4090), .Z(n4092) );
  XOR U5363 ( .A(n4386), .B(n4387), .Z(n4090) );
  ANDN U5364 ( .B(n4388), .A(n4389), .Z(n4386) );
  AND U5365 ( .A(b[6]), .B(a[44]), .Z(n4385) );
  XNOR U5366 ( .A(n4390), .B(n4095), .Z(n4097) );
  XOR U5367 ( .A(n4391), .B(n4392), .Z(n4095) );
  ANDN U5368 ( .B(n4393), .A(n4394), .Z(n4391) );
  AND U5369 ( .A(b[5]), .B(a[45]), .Z(n4390) );
  XNOR U5370 ( .A(n4395), .B(n4100), .Z(n4102) );
  XOR U5371 ( .A(n4396), .B(n4397), .Z(n4100) );
  ANDN U5372 ( .B(n4398), .A(n4399), .Z(n4396) );
  AND U5373 ( .A(b[4]), .B(a[46]), .Z(n4395) );
  XNOR U5374 ( .A(n4400), .B(n4401), .Z(n4114) );
  NANDN U5375 ( .A(n4402), .B(n4403), .Z(n4401) );
  XNOR U5376 ( .A(n4404), .B(n4105), .Z(n4107) );
  XNOR U5377 ( .A(n4405), .B(n4406), .Z(n4105) );
  NOR U5378 ( .A(n4407), .B(n4408), .Z(n4405) );
  AND U5379 ( .A(b[3]), .B(a[47]), .Z(n4404) );
  NAND U5380 ( .A(a[50]), .B(b[0]), .Z(n3821) );
  XNOR U5381 ( .A(n4409), .B(n4410), .Z(c[4]) );
  XNOR U5382 ( .A(n4120), .B(n4121), .Z(c[49]) );
  XOR U5383 ( .A(n4411), .B(n4412), .Z(n4402) );
  NAND U5384 ( .A(b[1]), .B(a[48]), .Z(n4412) );
  XOR U5385 ( .A(n4411), .B(n4408), .Z(n4413) );
  XOR U5386 ( .A(n4414), .B(n4406), .Z(n4408) );
  AND U5387 ( .A(b[2]), .B(a[47]), .Z(n4414) );
  IV U5388 ( .A(n4400), .Z(n4411) );
  NANDN U5389 ( .A(n4415), .B(n4416), .Z(n4400) );
  XOR U5390 ( .A(n4406), .B(n4398), .Z(n4417) );
  XNOR U5391 ( .A(n4397), .B(n4393), .Z(n4418) );
  XNOR U5392 ( .A(n4392), .B(n4388), .Z(n4419) );
  XNOR U5393 ( .A(n4387), .B(n4383), .Z(n4420) );
  XNOR U5394 ( .A(n4382), .B(n4378), .Z(n4421) );
  XNOR U5395 ( .A(n4377), .B(n4373), .Z(n4422) );
  XNOR U5396 ( .A(n4372), .B(n4368), .Z(n4423) );
  XNOR U5397 ( .A(n4367), .B(n4363), .Z(n4424) );
  XNOR U5398 ( .A(n4362), .B(n4358), .Z(n4425) );
  XNOR U5399 ( .A(n4357), .B(n4353), .Z(n4426) );
  XNOR U5400 ( .A(n4344), .B(n4343), .Z(n4427) );
  XOR U5401 ( .A(n4428), .B(n4342), .Z(n4343) );
  AND U5402 ( .A(b[13]), .B(a[36]), .Z(n4428) );
  XNOR U5403 ( .A(n4342), .B(n4348), .Z(n4429) );
  XNOR U5404 ( .A(n4347), .B(n4339), .Z(n4430) );
  XNOR U5405 ( .A(n4338), .B(n4334), .Z(n4431) );
  XNOR U5406 ( .A(n4333), .B(n4329), .Z(n4432) );
  XNOR U5407 ( .A(n4328), .B(n4324), .Z(n4433) );
  XNOR U5408 ( .A(n4315), .B(n4314), .Z(n4434) );
  XOR U5409 ( .A(n4435), .B(n4313), .Z(n4314) );
  AND U5410 ( .A(b[19]), .B(a[30]), .Z(n4435) );
  XNOR U5411 ( .A(n4313), .B(n4319), .Z(n4436) );
  XNOR U5412 ( .A(n4318), .B(n4310), .Z(n4437) );
  XNOR U5413 ( .A(n4309), .B(n4305), .Z(n4438) );
  XNOR U5414 ( .A(n4304), .B(n4300), .Z(n4439) );
  XNOR U5415 ( .A(n4299), .B(n4295), .Z(n4440) );
  XNOR U5416 ( .A(n4286), .B(n4285), .Z(n4441) );
  XOR U5417 ( .A(n4442), .B(n4284), .Z(n4285) );
  AND U5418 ( .A(b[25]), .B(a[24]), .Z(n4442) );
  XNOR U5419 ( .A(n4284), .B(n4290), .Z(n4443) );
  XNOR U5420 ( .A(n4289), .B(n4281), .Z(n4444) );
  XNOR U5421 ( .A(n4280), .B(n4276), .Z(n4445) );
  XNOR U5422 ( .A(n4275), .B(n4271), .Z(n4446) );
  XNOR U5423 ( .A(n4270), .B(n4266), .Z(n4447) );
  XNOR U5424 ( .A(n4257), .B(n4256), .Z(n4448) );
  XOR U5425 ( .A(n4449), .B(n4255), .Z(n4256) );
  AND U5426 ( .A(b[31]), .B(a[18]), .Z(n4449) );
  XNOR U5427 ( .A(n4255), .B(n4261), .Z(n4450) );
  XNOR U5428 ( .A(n4260), .B(n4252), .Z(n4451) );
  XNOR U5429 ( .A(n4251), .B(n4247), .Z(n4452) );
  XNOR U5430 ( .A(n4246), .B(n4242), .Z(n4453) );
  XNOR U5431 ( .A(n4241), .B(n4237), .Z(n4454) );
  XNOR U5432 ( .A(n4228), .B(n4227), .Z(n4455) );
  XOR U5433 ( .A(n4456), .B(n4226), .Z(n4227) );
  AND U5434 ( .A(b[37]), .B(a[12]), .Z(n4456) );
  XNOR U5435 ( .A(n4226), .B(n4232), .Z(n4457) );
  XNOR U5436 ( .A(n4231), .B(n4223), .Z(n4458) );
  XNOR U5437 ( .A(n4222), .B(n4218), .Z(n4459) );
  XNOR U5438 ( .A(n4217), .B(n4213), .Z(n4460) );
  XNOR U5439 ( .A(n4212), .B(n4208), .Z(n4461) );
  XNOR U5440 ( .A(n4199), .B(n4198), .Z(n4462) );
  XOR U5441 ( .A(n4463), .B(n4197), .Z(n4198) );
  AND U5442 ( .A(a[6]), .B(b[43]), .Z(n4463) );
  XNOR U5443 ( .A(n4197), .B(n4203), .Z(n4464) );
  XNOR U5444 ( .A(n4202), .B(n4194), .Z(n4465) );
  XNOR U5445 ( .A(n4193), .B(n4189), .Z(n4466) );
  XNOR U5446 ( .A(n4188), .B(n4184), .Z(n4467) );
  XNOR U5447 ( .A(n4183), .B(n4179), .Z(n4468) );
  XNOR U5448 ( .A(n4469), .B(n4178), .Z(n4179) );
  AND U5449 ( .A(a[0]), .B(b[49]), .Z(n4469) );
  XOR U5450 ( .A(n4470), .B(n4178), .Z(n4180) );
  XNOR U5451 ( .A(n4471), .B(n4472), .Z(n4178) );
  ANDN U5452 ( .B(n4473), .A(n4474), .Z(n4471) );
  AND U5453 ( .A(a[1]), .B(b[48]), .Z(n4470) );
  XNOR U5454 ( .A(n4475), .B(n4183), .Z(n4185) );
  XOR U5455 ( .A(n4476), .B(n4477), .Z(n4183) );
  ANDN U5456 ( .B(n4478), .A(n4479), .Z(n4476) );
  AND U5457 ( .A(a[2]), .B(b[47]), .Z(n4475) );
  XNOR U5458 ( .A(n4480), .B(n4188), .Z(n4190) );
  XOR U5459 ( .A(n4481), .B(n4482), .Z(n4188) );
  ANDN U5460 ( .B(n4483), .A(n4484), .Z(n4481) );
  AND U5461 ( .A(a[3]), .B(b[46]), .Z(n4480) );
  XNOR U5462 ( .A(n4485), .B(n4193), .Z(n4195) );
  XOR U5463 ( .A(n4486), .B(n4487), .Z(n4193) );
  ANDN U5464 ( .B(n4488), .A(n4489), .Z(n4486) );
  AND U5465 ( .A(a[4]), .B(b[45]), .Z(n4485) );
  XOR U5466 ( .A(n4490), .B(n4491), .Z(n4197) );
  AND U5467 ( .A(n4492), .B(n4493), .Z(n4490) );
  XNOR U5468 ( .A(n4494), .B(n4202), .Z(n4204) );
  XOR U5469 ( .A(n4495), .B(n4496), .Z(n4202) );
  ANDN U5470 ( .B(n4497), .A(n4498), .Z(n4495) );
  AND U5471 ( .A(a[5]), .B(b[44]), .Z(n4494) );
  XOR U5472 ( .A(n4499), .B(n4207), .Z(n4209) );
  XOR U5473 ( .A(n4500), .B(n4501), .Z(n4207) );
  ANDN U5474 ( .B(n4502), .A(n4503), .Z(n4500) );
  AND U5475 ( .A(a[7]), .B(b[42]), .Z(n4499) );
  XNOR U5476 ( .A(n4504), .B(n4212), .Z(n4214) );
  XOR U5477 ( .A(n4505), .B(n4506), .Z(n4212) );
  ANDN U5478 ( .B(n4507), .A(n4508), .Z(n4505) );
  AND U5479 ( .A(a[8]), .B(b[41]), .Z(n4504) );
  XNOR U5480 ( .A(n4509), .B(n4217), .Z(n4219) );
  XOR U5481 ( .A(n4510), .B(n4511), .Z(n4217) );
  ANDN U5482 ( .B(n4512), .A(n4513), .Z(n4510) );
  AND U5483 ( .A(a[9]), .B(b[40]), .Z(n4509) );
  XNOR U5484 ( .A(n4514), .B(n4222), .Z(n4224) );
  XOR U5485 ( .A(n4515), .B(n4516), .Z(n4222) );
  ANDN U5486 ( .B(n4517), .A(n4518), .Z(n4515) );
  AND U5487 ( .A(a[10]), .B(b[39]), .Z(n4514) );
  XOR U5488 ( .A(n4519), .B(n4520), .Z(n4226) );
  AND U5489 ( .A(n4521), .B(n4522), .Z(n4519) );
  XNOR U5490 ( .A(n4523), .B(n4231), .Z(n4233) );
  XOR U5491 ( .A(n4524), .B(n4525), .Z(n4231) );
  ANDN U5492 ( .B(n4526), .A(n4527), .Z(n4524) );
  AND U5493 ( .A(b[38]), .B(a[11]), .Z(n4523) );
  XOR U5494 ( .A(n4528), .B(n4236), .Z(n4238) );
  XOR U5495 ( .A(n4529), .B(n4530), .Z(n4236) );
  ANDN U5496 ( .B(n4531), .A(n4532), .Z(n4529) );
  AND U5497 ( .A(b[36]), .B(a[13]), .Z(n4528) );
  XNOR U5498 ( .A(n4533), .B(n4241), .Z(n4243) );
  XOR U5499 ( .A(n4534), .B(n4535), .Z(n4241) );
  ANDN U5500 ( .B(n4536), .A(n4537), .Z(n4534) );
  AND U5501 ( .A(b[35]), .B(a[14]), .Z(n4533) );
  XNOR U5502 ( .A(n4538), .B(n4246), .Z(n4248) );
  XOR U5503 ( .A(n4539), .B(n4540), .Z(n4246) );
  ANDN U5504 ( .B(n4541), .A(n4542), .Z(n4539) );
  AND U5505 ( .A(b[34]), .B(a[15]), .Z(n4538) );
  XNOR U5506 ( .A(n4543), .B(n4251), .Z(n4253) );
  XOR U5507 ( .A(n4544), .B(n4545), .Z(n4251) );
  ANDN U5508 ( .B(n4546), .A(n4547), .Z(n4544) );
  AND U5509 ( .A(a[16]), .B(b[33]), .Z(n4543) );
  XOR U5510 ( .A(n4548), .B(n4549), .Z(n4255) );
  AND U5511 ( .A(n4550), .B(n4551), .Z(n4548) );
  XNOR U5512 ( .A(n4552), .B(n4260), .Z(n4262) );
  XOR U5513 ( .A(n4553), .B(n4554), .Z(n4260) );
  ANDN U5514 ( .B(n4555), .A(n4556), .Z(n4553) );
  AND U5515 ( .A(b[32]), .B(a[17]), .Z(n4552) );
  XOR U5516 ( .A(n4557), .B(n4265), .Z(n4267) );
  XOR U5517 ( .A(n4558), .B(n4559), .Z(n4265) );
  ANDN U5518 ( .B(n4560), .A(n4561), .Z(n4558) );
  AND U5519 ( .A(b[30]), .B(a[19]), .Z(n4557) );
  XNOR U5520 ( .A(n4562), .B(n4270), .Z(n4272) );
  XOR U5521 ( .A(n4563), .B(n4564), .Z(n4270) );
  ANDN U5522 ( .B(n4565), .A(n4566), .Z(n4563) );
  AND U5523 ( .A(b[29]), .B(a[20]), .Z(n4562) );
  XNOR U5524 ( .A(n4567), .B(n4275), .Z(n4277) );
  XOR U5525 ( .A(n4568), .B(n4569), .Z(n4275) );
  ANDN U5526 ( .B(n4570), .A(n4571), .Z(n4568) );
  AND U5527 ( .A(b[28]), .B(a[21]), .Z(n4567) );
  XNOR U5528 ( .A(n4572), .B(n4280), .Z(n4282) );
  XOR U5529 ( .A(n4573), .B(n4574), .Z(n4280) );
  ANDN U5530 ( .B(n4575), .A(n4576), .Z(n4573) );
  AND U5531 ( .A(a[22]), .B(b[27]), .Z(n4572) );
  XOR U5532 ( .A(n4577), .B(n4578), .Z(n4284) );
  AND U5533 ( .A(n4579), .B(n4580), .Z(n4577) );
  XNOR U5534 ( .A(n4581), .B(n4289), .Z(n4291) );
  XOR U5535 ( .A(n4582), .B(n4583), .Z(n4289) );
  ANDN U5536 ( .B(n4584), .A(n4585), .Z(n4582) );
  AND U5537 ( .A(b[26]), .B(a[23]), .Z(n4581) );
  XOR U5538 ( .A(n4586), .B(n4294), .Z(n4296) );
  XOR U5539 ( .A(n4587), .B(n4588), .Z(n4294) );
  ANDN U5540 ( .B(n4589), .A(n4590), .Z(n4587) );
  AND U5541 ( .A(b[24]), .B(a[25]), .Z(n4586) );
  XNOR U5542 ( .A(n4591), .B(n4299), .Z(n4301) );
  XOR U5543 ( .A(n4592), .B(n4593), .Z(n4299) );
  ANDN U5544 ( .B(n4594), .A(n4595), .Z(n4592) );
  AND U5545 ( .A(b[23]), .B(a[26]), .Z(n4591) );
  XNOR U5546 ( .A(n4596), .B(n4304), .Z(n4306) );
  XOR U5547 ( .A(n4597), .B(n4598), .Z(n4304) );
  ANDN U5548 ( .B(n4599), .A(n4600), .Z(n4597) );
  AND U5549 ( .A(b[22]), .B(a[27]), .Z(n4596) );
  XNOR U5550 ( .A(n4601), .B(n4309), .Z(n4311) );
  XOR U5551 ( .A(n4602), .B(n4603), .Z(n4309) );
  ANDN U5552 ( .B(n4604), .A(n4605), .Z(n4602) );
  AND U5553 ( .A(a[28]), .B(b[21]), .Z(n4601) );
  XOR U5554 ( .A(n4606), .B(n4607), .Z(n4313) );
  AND U5555 ( .A(n4608), .B(n4609), .Z(n4606) );
  XNOR U5556 ( .A(n4610), .B(n4318), .Z(n4320) );
  XOR U5557 ( .A(n4611), .B(n4612), .Z(n4318) );
  ANDN U5558 ( .B(n4613), .A(n4614), .Z(n4611) );
  AND U5559 ( .A(b[20]), .B(a[29]), .Z(n4610) );
  XOR U5560 ( .A(n4615), .B(n4323), .Z(n4325) );
  XOR U5561 ( .A(n4616), .B(n4617), .Z(n4323) );
  ANDN U5562 ( .B(n4618), .A(n4619), .Z(n4616) );
  AND U5563 ( .A(b[18]), .B(a[31]), .Z(n4615) );
  XNOR U5564 ( .A(n4620), .B(n4328), .Z(n4330) );
  XOR U5565 ( .A(n4621), .B(n4622), .Z(n4328) );
  ANDN U5566 ( .B(n4623), .A(n4624), .Z(n4621) );
  AND U5567 ( .A(b[17]), .B(a[32]), .Z(n4620) );
  XNOR U5568 ( .A(n4625), .B(n4333), .Z(n4335) );
  XOR U5569 ( .A(n4626), .B(n4627), .Z(n4333) );
  ANDN U5570 ( .B(n4628), .A(n4629), .Z(n4626) );
  AND U5571 ( .A(b[16]), .B(a[33]), .Z(n4625) );
  XNOR U5572 ( .A(n4630), .B(n4338), .Z(n4340) );
  XOR U5573 ( .A(n4631), .B(n4632), .Z(n4338) );
  ANDN U5574 ( .B(n4633), .A(n4634), .Z(n4631) );
  AND U5575 ( .A(a[34]), .B(b[15]), .Z(n4630) );
  XOR U5576 ( .A(n4635), .B(n4636), .Z(n4342) );
  AND U5577 ( .A(n4637), .B(n4638), .Z(n4635) );
  XNOR U5578 ( .A(n4639), .B(n4347), .Z(n4349) );
  XOR U5579 ( .A(n4640), .B(n4641), .Z(n4347) );
  ANDN U5580 ( .B(n4642), .A(n4643), .Z(n4640) );
  AND U5581 ( .A(b[14]), .B(a[35]), .Z(n4639) );
  XOR U5582 ( .A(n4644), .B(n4352), .Z(n4354) );
  XOR U5583 ( .A(n4645), .B(n4646), .Z(n4352) );
  ANDN U5584 ( .B(n4647), .A(n4648), .Z(n4645) );
  AND U5585 ( .A(b[12]), .B(a[37]), .Z(n4644) );
  XNOR U5586 ( .A(n4649), .B(n4357), .Z(n4359) );
  XOR U5587 ( .A(n4650), .B(n4651), .Z(n4357) );
  ANDN U5588 ( .B(n4652), .A(n4653), .Z(n4650) );
  AND U5589 ( .A(b[11]), .B(a[38]), .Z(n4649) );
  XNOR U5590 ( .A(n4654), .B(n4362), .Z(n4364) );
  XOR U5591 ( .A(n4655), .B(n4656), .Z(n4362) );
  ANDN U5592 ( .B(n4657), .A(n4658), .Z(n4655) );
  AND U5593 ( .A(b[10]), .B(a[39]), .Z(n4654) );
  XNOR U5594 ( .A(n4659), .B(n4367), .Z(n4369) );
  XOR U5595 ( .A(n4660), .B(n4661), .Z(n4367) );
  ANDN U5596 ( .B(n4662), .A(n4663), .Z(n4660) );
  AND U5597 ( .A(b[9]), .B(a[40]), .Z(n4659) );
  XNOR U5598 ( .A(n4664), .B(n4372), .Z(n4374) );
  XOR U5599 ( .A(n4665), .B(n4666), .Z(n4372) );
  ANDN U5600 ( .B(n4667), .A(n4668), .Z(n4665) );
  AND U5601 ( .A(b[8]), .B(a[41]), .Z(n4664) );
  XNOR U5602 ( .A(n4669), .B(n4377), .Z(n4379) );
  XOR U5603 ( .A(n4670), .B(n4671), .Z(n4377) );
  ANDN U5604 ( .B(n4672), .A(n4673), .Z(n4670) );
  AND U5605 ( .A(b[7]), .B(a[42]), .Z(n4669) );
  XNOR U5606 ( .A(n4674), .B(n4382), .Z(n4384) );
  XOR U5607 ( .A(n4675), .B(n4676), .Z(n4382) );
  ANDN U5608 ( .B(n4677), .A(n4678), .Z(n4675) );
  AND U5609 ( .A(b[6]), .B(a[43]), .Z(n4674) );
  XNOR U5610 ( .A(n4679), .B(n4387), .Z(n4389) );
  XOR U5611 ( .A(n4680), .B(n4681), .Z(n4387) );
  ANDN U5612 ( .B(n4682), .A(n4683), .Z(n4680) );
  AND U5613 ( .A(b[5]), .B(a[44]), .Z(n4679) );
  XNOR U5614 ( .A(n4684), .B(n4392), .Z(n4394) );
  XOR U5615 ( .A(n4685), .B(n4686), .Z(n4392) );
  ANDN U5616 ( .B(n4687), .A(n4688), .Z(n4685) );
  AND U5617 ( .A(b[4]), .B(a[45]), .Z(n4684) );
  XOR U5618 ( .A(n4689), .B(n4690), .Z(n4406) );
  NANDN U5619 ( .A(n4691), .B(n4692), .Z(n4690) );
  XNOR U5620 ( .A(n4693), .B(n4397), .Z(n4399) );
  XNOR U5621 ( .A(n4694), .B(n4695), .Z(n4397) );
  AND U5622 ( .A(n4696), .B(n4697), .Z(n4694) );
  AND U5623 ( .A(b[3]), .B(a[46]), .Z(n4693) );
  NAND U5624 ( .A(a[49]), .B(b[0]), .Z(n4120) );
  XNOR U5625 ( .A(n4415), .B(n4416), .Z(c[48]) );
  XNOR U5626 ( .A(n4692), .B(n4691), .Z(n4416) );
  XOR U5627 ( .A(n4689), .B(n4698), .Z(n4691) );
  NAND U5628 ( .A(b[1]), .B(a[47]), .Z(n4698) );
  XNOR U5629 ( .A(n4697), .B(n4699), .Z(n4692) );
  XNOR U5630 ( .A(n4689), .B(n4696), .Z(n4699) );
  XNOR U5631 ( .A(n4700), .B(n4695), .Z(n4696) );
  AND U5632 ( .A(b[2]), .B(a[46]), .Z(n4700) );
  ANDN U5633 ( .B(n4701), .A(n4702), .Z(n4689) );
  XOR U5634 ( .A(n4695), .B(n4687), .Z(n4703) );
  XNOR U5635 ( .A(n4686), .B(n4682), .Z(n4704) );
  XNOR U5636 ( .A(n4681), .B(n4677), .Z(n4705) );
  XNOR U5637 ( .A(n4676), .B(n4672), .Z(n4706) );
  XNOR U5638 ( .A(n4671), .B(n4667), .Z(n4707) );
  XNOR U5639 ( .A(n4666), .B(n4662), .Z(n4708) );
  XNOR U5640 ( .A(n4661), .B(n4657), .Z(n4709) );
  XNOR U5641 ( .A(n4656), .B(n4652), .Z(n4710) );
  XNOR U5642 ( .A(n4651), .B(n4647), .Z(n4711) );
  XNOR U5643 ( .A(n4638), .B(n4637), .Z(n4712) );
  XOR U5644 ( .A(n4713), .B(n4636), .Z(n4637) );
  AND U5645 ( .A(b[12]), .B(a[36]), .Z(n4713) );
  XNOR U5646 ( .A(n4636), .B(n4642), .Z(n4714) );
  XNOR U5647 ( .A(n4641), .B(n4633), .Z(n4715) );
  XNOR U5648 ( .A(n4632), .B(n4628), .Z(n4716) );
  XNOR U5649 ( .A(n4627), .B(n4623), .Z(n4717) );
  XNOR U5650 ( .A(n4622), .B(n4618), .Z(n4718) );
  XNOR U5651 ( .A(n4609), .B(n4608), .Z(n4719) );
  XOR U5652 ( .A(n4720), .B(n4607), .Z(n4608) );
  AND U5653 ( .A(b[18]), .B(a[30]), .Z(n4720) );
  XNOR U5654 ( .A(n4607), .B(n4613), .Z(n4721) );
  XNOR U5655 ( .A(n4612), .B(n4604), .Z(n4722) );
  XNOR U5656 ( .A(n4603), .B(n4599), .Z(n4723) );
  XNOR U5657 ( .A(n4598), .B(n4594), .Z(n4724) );
  XNOR U5658 ( .A(n4593), .B(n4589), .Z(n4725) );
  XNOR U5659 ( .A(n4580), .B(n4579), .Z(n4726) );
  XOR U5660 ( .A(n4727), .B(n4578), .Z(n4579) );
  AND U5661 ( .A(b[24]), .B(a[24]), .Z(n4727) );
  XNOR U5662 ( .A(n4578), .B(n4584), .Z(n4728) );
  XNOR U5663 ( .A(n4583), .B(n4575), .Z(n4729) );
  XNOR U5664 ( .A(n4574), .B(n4570), .Z(n4730) );
  XNOR U5665 ( .A(n4569), .B(n4565), .Z(n4731) );
  XNOR U5666 ( .A(n4564), .B(n4560), .Z(n4732) );
  XNOR U5667 ( .A(n4551), .B(n4550), .Z(n4733) );
  XOR U5668 ( .A(n4734), .B(n4549), .Z(n4550) );
  AND U5669 ( .A(b[30]), .B(a[18]), .Z(n4734) );
  XNOR U5670 ( .A(n4549), .B(n4555), .Z(n4735) );
  XNOR U5671 ( .A(n4554), .B(n4546), .Z(n4736) );
  XNOR U5672 ( .A(n4545), .B(n4541), .Z(n4737) );
  XNOR U5673 ( .A(n4540), .B(n4536), .Z(n4738) );
  XNOR U5674 ( .A(n4535), .B(n4531), .Z(n4739) );
  XNOR U5675 ( .A(n4522), .B(n4521), .Z(n4740) );
  XOR U5676 ( .A(n4741), .B(n4520), .Z(n4521) );
  AND U5677 ( .A(b[36]), .B(a[12]), .Z(n4741) );
  XNOR U5678 ( .A(n4520), .B(n4526), .Z(n4742) );
  XNOR U5679 ( .A(n4525), .B(n4517), .Z(n4743) );
  XNOR U5680 ( .A(n4516), .B(n4512), .Z(n4744) );
  XNOR U5681 ( .A(n4511), .B(n4507), .Z(n4745) );
  XNOR U5682 ( .A(n4506), .B(n4502), .Z(n4746) );
  XNOR U5683 ( .A(n4493), .B(n4492), .Z(n4747) );
  XOR U5684 ( .A(n4748), .B(n4491), .Z(n4492) );
  AND U5685 ( .A(a[6]), .B(b[42]), .Z(n4748) );
  XNOR U5686 ( .A(n4491), .B(n4497), .Z(n4749) );
  XNOR U5687 ( .A(n4496), .B(n4488), .Z(n4750) );
  XNOR U5688 ( .A(n4487), .B(n4483), .Z(n4751) );
  XNOR U5689 ( .A(n4482), .B(n4478), .Z(n4752) );
  XNOR U5690 ( .A(n4477), .B(n4473), .Z(n4753) );
  XOR U5691 ( .A(n4754), .B(n4472), .Z(n4473) );
  AND U5692 ( .A(a[0]), .B(b[48]), .Z(n4754) );
  XNOR U5693 ( .A(n4755), .B(n4472), .Z(n4474) );
  XNOR U5694 ( .A(n4756), .B(n4757), .Z(n4472) );
  ANDN U5695 ( .B(n4758), .A(n4759), .Z(n4756) );
  AND U5696 ( .A(a[1]), .B(b[47]), .Z(n4755) );
  XNOR U5697 ( .A(n4760), .B(n4477), .Z(n4479) );
  XOR U5698 ( .A(n4761), .B(n4762), .Z(n4477) );
  ANDN U5699 ( .B(n4763), .A(n4764), .Z(n4761) );
  AND U5700 ( .A(a[2]), .B(b[46]), .Z(n4760) );
  XNOR U5701 ( .A(n4765), .B(n4482), .Z(n4484) );
  XOR U5702 ( .A(n4766), .B(n4767), .Z(n4482) );
  ANDN U5703 ( .B(n4768), .A(n4769), .Z(n4766) );
  AND U5704 ( .A(a[3]), .B(b[45]), .Z(n4765) );
  XNOR U5705 ( .A(n4770), .B(n4487), .Z(n4489) );
  XOR U5706 ( .A(n4771), .B(n4772), .Z(n4487) );
  ANDN U5707 ( .B(n4773), .A(n4774), .Z(n4771) );
  AND U5708 ( .A(a[4]), .B(b[44]), .Z(n4770) );
  XOR U5709 ( .A(n4775), .B(n4776), .Z(n4491) );
  AND U5710 ( .A(n4777), .B(n4778), .Z(n4775) );
  XNOR U5711 ( .A(n4779), .B(n4496), .Z(n4498) );
  XOR U5712 ( .A(n4780), .B(n4781), .Z(n4496) );
  ANDN U5713 ( .B(n4782), .A(n4783), .Z(n4780) );
  AND U5714 ( .A(a[5]), .B(b[43]), .Z(n4779) );
  XOR U5715 ( .A(n4784), .B(n4501), .Z(n4503) );
  XOR U5716 ( .A(n4785), .B(n4786), .Z(n4501) );
  ANDN U5717 ( .B(n4787), .A(n4788), .Z(n4785) );
  AND U5718 ( .A(a[7]), .B(b[41]), .Z(n4784) );
  XNOR U5719 ( .A(n4789), .B(n4506), .Z(n4508) );
  XOR U5720 ( .A(n4790), .B(n4791), .Z(n4506) );
  ANDN U5721 ( .B(n4792), .A(n4793), .Z(n4790) );
  AND U5722 ( .A(a[8]), .B(b[40]), .Z(n4789) );
  XNOR U5723 ( .A(n4794), .B(n4511), .Z(n4513) );
  XOR U5724 ( .A(n4795), .B(n4796), .Z(n4511) );
  ANDN U5725 ( .B(n4797), .A(n4798), .Z(n4795) );
  AND U5726 ( .A(a[9]), .B(b[39]), .Z(n4794) );
  XNOR U5727 ( .A(n4799), .B(n4516), .Z(n4518) );
  XOR U5728 ( .A(n4800), .B(n4801), .Z(n4516) );
  ANDN U5729 ( .B(n4802), .A(n4803), .Z(n4800) );
  AND U5730 ( .A(b[38]), .B(a[10]), .Z(n4799) );
  XOR U5731 ( .A(n4804), .B(n4805), .Z(n4520) );
  AND U5732 ( .A(n4806), .B(n4807), .Z(n4804) );
  XNOR U5733 ( .A(n4808), .B(n4525), .Z(n4527) );
  XOR U5734 ( .A(n4809), .B(n4810), .Z(n4525) );
  ANDN U5735 ( .B(n4811), .A(n4812), .Z(n4809) );
  AND U5736 ( .A(b[37]), .B(a[11]), .Z(n4808) );
  XOR U5737 ( .A(n4813), .B(n4530), .Z(n4532) );
  XOR U5738 ( .A(n4814), .B(n4815), .Z(n4530) );
  ANDN U5739 ( .B(n4816), .A(n4817), .Z(n4814) );
  AND U5740 ( .A(b[35]), .B(a[13]), .Z(n4813) );
  XNOR U5741 ( .A(n4818), .B(n4535), .Z(n4537) );
  XOR U5742 ( .A(n4819), .B(n4820), .Z(n4535) );
  ANDN U5743 ( .B(n4821), .A(n4822), .Z(n4819) );
  AND U5744 ( .A(b[34]), .B(a[14]), .Z(n4818) );
  XNOR U5745 ( .A(n4823), .B(n4540), .Z(n4542) );
  XOR U5746 ( .A(n4824), .B(n4825), .Z(n4540) );
  ANDN U5747 ( .B(n4826), .A(n4827), .Z(n4824) );
  AND U5748 ( .A(a[15]), .B(b[33]), .Z(n4823) );
  XNOR U5749 ( .A(n4828), .B(n4545), .Z(n4547) );
  XOR U5750 ( .A(n4829), .B(n4830), .Z(n4545) );
  ANDN U5751 ( .B(n4831), .A(n4832), .Z(n4829) );
  AND U5752 ( .A(b[32]), .B(a[16]), .Z(n4828) );
  XOR U5753 ( .A(n4833), .B(n4834), .Z(n4549) );
  AND U5754 ( .A(n4835), .B(n4836), .Z(n4833) );
  XNOR U5755 ( .A(n4837), .B(n4554), .Z(n4556) );
  XOR U5756 ( .A(n4838), .B(n4839), .Z(n4554) );
  ANDN U5757 ( .B(n4840), .A(n4841), .Z(n4838) );
  AND U5758 ( .A(b[31]), .B(a[17]), .Z(n4837) );
  XOR U5759 ( .A(n4842), .B(n4559), .Z(n4561) );
  XOR U5760 ( .A(n4843), .B(n4844), .Z(n4559) );
  ANDN U5761 ( .B(n4845), .A(n4846), .Z(n4843) );
  AND U5762 ( .A(b[29]), .B(a[19]), .Z(n4842) );
  XNOR U5763 ( .A(n4847), .B(n4564), .Z(n4566) );
  XOR U5764 ( .A(n4848), .B(n4849), .Z(n4564) );
  ANDN U5765 ( .B(n4850), .A(n4851), .Z(n4848) );
  AND U5766 ( .A(b[28]), .B(a[20]), .Z(n4847) );
  XNOR U5767 ( .A(n4852), .B(n4569), .Z(n4571) );
  XOR U5768 ( .A(n4853), .B(n4854), .Z(n4569) );
  ANDN U5769 ( .B(n4855), .A(n4856), .Z(n4853) );
  AND U5770 ( .A(a[21]), .B(b[27]), .Z(n4852) );
  XNOR U5771 ( .A(n4857), .B(n4574), .Z(n4576) );
  XOR U5772 ( .A(n4858), .B(n4859), .Z(n4574) );
  ANDN U5773 ( .B(n4860), .A(n4861), .Z(n4858) );
  AND U5774 ( .A(b[26]), .B(a[22]), .Z(n4857) );
  XOR U5775 ( .A(n4862), .B(n4863), .Z(n4578) );
  AND U5776 ( .A(n4864), .B(n4865), .Z(n4862) );
  XNOR U5777 ( .A(n4866), .B(n4583), .Z(n4585) );
  XOR U5778 ( .A(n4867), .B(n4868), .Z(n4583) );
  ANDN U5779 ( .B(n4869), .A(n4870), .Z(n4867) );
  AND U5780 ( .A(b[25]), .B(a[23]), .Z(n4866) );
  XOR U5781 ( .A(n4871), .B(n4588), .Z(n4590) );
  XOR U5782 ( .A(n4872), .B(n4873), .Z(n4588) );
  ANDN U5783 ( .B(n4874), .A(n4875), .Z(n4872) );
  AND U5784 ( .A(b[23]), .B(a[25]), .Z(n4871) );
  XNOR U5785 ( .A(n4876), .B(n4593), .Z(n4595) );
  XOR U5786 ( .A(n4877), .B(n4878), .Z(n4593) );
  ANDN U5787 ( .B(n4879), .A(n4880), .Z(n4877) );
  AND U5788 ( .A(b[22]), .B(a[26]), .Z(n4876) );
  XNOR U5789 ( .A(n4881), .B(n4598), .Z(n4600) );
  XOR U5790 ( .A(n4882), .B(n4883), .Z(n4598) );
  ANDN U5791 ( .B(n4884), .A(n4885), .Z(n4882) );
  AND U5792 ( .A(a[27]), .B(b[21]), .Z(n4881) );
  XNOR U5793 ( .A(n4886), .B(n4603), .Z(n4605) );
  XOR U5794 ( .A(n4887), .B(n4888), .Z(n4603) );
  ANDN U5795 ( .B(n4889), .A(n4890), .Z(n4887) );
  AND U5796 ( .A(b[20]), .B(a[28]), .Z(n4886) );
  XOR U5797 ( .A(n4891), .B(n4892), .Z(n4607) );
  AND U5798 ( .A(n4893), .B(n4894), .Z(n4891) );
  XNOR U5799 ( .A(n4895), .B(n4612), .Z(n4614) );
  XOR U5800 ( .A(n4896), .B(n4897), .Z(n4612) );
  ANDN U5801 ( .B(n4898), .A(n4899), .Z(n4896) );
  AND U5802 ( .A(b[19]), .B(a[29]), .Z(n4895) );
  XOR U5803 ( .A(n4900), .B(n4617), .Z(n4619) );
  XOR U5804 ( .A(n4901), .B(n4902), .Z(n4617) );
  ANDN U5805 ( .B(n4903), .A(n4904), .Z(n4901) );
  AND U5806 ( .A(b[17]), .B(a[31]), .Z(n4900) );
  XNOR U5807 ( .A(n4905), .B(n4622), .Z(n4624) );
  XOR U5808 ( .A(n4906), .B(n4907), .Z(n4622) );
  ANDN U5809 ( .B(n4908), .A(n4909), .Z(n4906) );
  AND U5810 ( .A(b[16]), .B(a[32]), .Z(n4905) );
  XNOR U5811 ( .A(n4910), .B(n4627), .Z(n4629) );
  XOR U5812 ( .A(n4911), .B(n4912), .Z(n4627) );
  ANDN U5813 ( .B(n4913), .A(n4914), .Z(n4911) );
  AND U5814 ( .A(a[33]), .B(b[15]), .Z(n4910) );
  XNOR U5815 ( .A(n4915), .B(n4632), .Z(n4634) );
  XOR U5816 ( .A(n4916), .B(n4917), .Z(n4632) );
  ANDN U5817 ( .B(n4918), .A(n4919), .Z(n4916) );
  AND U5818 ( .A(b[14]), .B(a[34]), .Z(n4915) );
  XOR U5819 ( .A(n4920), .B(n4921), .Z(n4636) );
  AND U5820 ( .A(n4922), .B(n4923), .Z(n4920) );
  XNOR U5821 ( .A(n4924), .B(n4641), .Z(n4643) );
  XOR U5822 ( .A(n4925), .B(n4926), .Z(n4641) );
  ANDN U5823 ( .B(n4927), .A(n4928), .Z(n4925) );
  AND U5824 ( .A(b[13]), .B(a[35]), .Z(n4924) );
  XOR U5825 ( .A(n4929), .B(n4646), .Z(n4648) );
  XOR U5826 ( .A(n4930), .B(n4931), .Z(n4646) );
  ANDN U5827 ( .B(n4932), .A(n4933), .Z(n4930) );
  AND U5828 ( .A(b[11]), .B(a[37]), .Z(n4929) );
  XNOR U5829 ( .A(n4934), .B(n4651), .Z(n4653) );
  XOR U5830 ( .A(n4935), .B(n4936), .Z(n4651) );
  ANDN U5831 ( .B(n4937), .A(n4938), .Z(n4935) );
  AND U5832 ( .A(b[10]), .B(a[38]), .Z(n4934) );
  XNOR U5833 ( .A(n4939), .B(n4656), .Z(n4658) );
  XOR U5834 ( .A(n4940), .B(n4941), .Z(n4656) );
  ANDN U5835 ( .B(n4942), .A(n4943), .Z(n4940) );
  AND U5836 ( .A(b[9]), .B(a[39]), .Z(n4939) );
  XNOR U5837 ( .A(n4944), .B(n4661), .Z(n4663) );
  XOR U5838 ( .A(n4945), .B(n4946), .Z(n4661) );
  ANDN U5839 ( .B(n4947), .A(n4948), .Z(n4945) );
  AND U5840 ( .A(b[8]), .B(a[40]), .Z(n4944) );
  XNOR U5841 ( .A(n4949), .B(n4666), .Z(n4668) );
  XOR U5842 ( .A(n4950), .B(n4951), .Z(n4666) );
  ANDN U5843 ( .B(n4952), .A(n4953), .Z(n4950) );
  AND U5844 ( .A(b[7]), .B(a[41]), .Z(n4949) );
  XNOR U5845 ( .A(n4954), .B(n4671), .Z(n4673) );
  XOR U5846 ( .A(n4955), .B(n4956), .Z(n4671) );
  ANDN U5847 ( .B(n4957), .A(n4958), .Z(n4955) );
  AND U5848 ( .A(b[6]), .B(a[42]), .Z(n4954) );
  XNOR U5849 ( .A(n4959), .B(n4676), .Z(n4678) );
  XOR U5850 ( .A(n4960), .B(n4961), .Z(n4676) );
  ANDN U5851 ( .B(n4962), .A(n4963), .Z(n4960) );
  AND U5852 ( .A(b[5]), .B(a[43]), .Z(n4959) );
  XNOR U5853 ( .A(n4964), .B(n4681), .Z(n4683) );
  XOR U5854 ( .A(n4965), .B(n4966), .Z(n4681) );
  ANDN U5855 ( .B(n4967), .A(n4968), .Z(n4965) );
  AND U5856 ( .A(b[4]), .B(a[44]), .Z(n4964) );
  XNOR U5857 ( .A(n4969), .B(n4970), .Z(n4695) );
  NANDN U5858 ( .A(n4971), .B(n4972), .Z(n4970) );
  XNOR U5859 ( .A(n4973), .B(n4686), .Z(n4688) );
  XNOR U5860 ( .A(n4974), .B(n4975), .Z(n4686) );
  AND U5861 ( .A(n4976), .B(n4977), .Z(n4974) );
  AND U5862 ( .A(b[3]), .B(a[45]), .Z(n4973) );
  NAND U5863 ( .A(a[48]), .B(b[0]), .Z(n4415) );
  XNOR U5864 ( .A(n4702), .B(n4701), .Z(c[47]) );
  XNOR U5865 ( .A(n4971), .B(n4972), .Z(n4701) );
  XOR U5866 ( .A(n4969), .B(n4978), .Z(n4972) );
  NAND U5867 ( .A(b[1]), .B(a[46]), .Z(n4978) );
  XOR U5868 ( .A(n4977), .B(n4979), .Z(n4971) );
  XOR U5869 ( .A(n4969), .B(n4976), .Z(n4979) );
  XNOR U5870 ( .A(n4980), .B(n4975), .Z(n4976) );
  AND U5871 ( .A(b[2]), .B(a[45]), .Z(n4980) );
  NANDN U5872 ( .A(n4981), .B(n4982), .Z(n4969) );
  XOR U5873 ( .A(n4975), .B(n4967), .Z(n4983) );
  XNOR U5874 ( .A(n4966), .B(n4962), .Z(n4984) );
  XNOR U5875 ( .A(n4961), .B(n4957), .Z(n4985) );
  XNOR U5876 ( .A(n4956), .B(n4952), .Z(n4986) );
  XNOR U5877 ( .A(n4951), .B(n4947), .Z(n4987) );
  XNOR U5878 ( .A(n4946), .B(n4942), .Z(n4988) );
  XNOR U5879 ( .A(n4941), .B(n4937), .Z(n4989) );
  XNOR U5880 ( .A(n4936), .B(n4932), .Z(n4990) );
  XNOR U5881 ( .A(n4923), .B(n4922), .Z(n4991) );
  XOR U5882 ( .A(n4992), .B(n4921), .Z(n4922) );
  AND U5883 ( .A(b[11]), .B(a[36]), .Z(n4992) );
  XNOR U5884 ( .A(n4921), .B(n4927), .Z(n4993) );
  XNOR U5885 ( .A(n4926), .B(n4918), .Z(n4994) );
  XNOR U5886 ( .A(n4917), .B(n4913), .Z(n4995) );
  XNOR U5887 ( .A(n4912), .B(n4908), .Z(n4996) );
  XNOR U5888 ( .A(n4907), .B(n4903), .Z(n4997) );
  XNOR U5889 ( .A(n4894), .B(n4893), .Z(n4998) );
  XOR U5890 ( .A(n4999), .B(n4892), .Z(n4893) );
  AND U5891 ( .A(b[17]), .B(a[30]), .Z(n4999) );
  XNOR U5892 ( .A(n4892), .B(n4898), .Z(n5000) );
  XNOR U5893 ( .A(n4897), .B(n4889), .Z(n5001) );
  XNOR U5894 ( .A(n4888), .B(n4884), .Z(n5002) );
  XNOR U5895 ( .A(n4883), .B(n4879), .Z(n5003) );
  XNOR U5896 ( .A(n4878), .B(n4874), .Z(n5004) );
  XNOR U5897 ( .A(n4865), .B(n4864), .Z(n5005) );
  XOR U5898 ( .A(n5006), .B(n4863), .Z(n4864) );
  AND U5899 ( .A(b[23]), .B(a[24]), .Z(n5006) );
  XNOR U5900 ( .A(n4863), .B(n4869), .Z(n5007) );
  XNOR U5901 ( .A(n4868), .B(n4860), .Z(n5008) );
  XNOR U5902 ( .A(n4859), .B(n4855), .Z(n5009) );
  XNOR U5903 ( .A(n4854), .B(n4850), .Z(n5010) );
  XNOR U5904 ( .A(n4849), .B(n4845), .Z(n5011) );
  XNOR U5905 ( .A(n5012), .B(n5013), .Z(n4845) );
  XNOR U5906 ( .A(n4836), .B(n4835), .Z(n5013) );
  XOR U5907 ( .A(n5014), .B(n4834), .Z(n4835) );
  AND U5908 ( .A(b[29]), .B(a[18]), .Z(n5014) );
  XNOR U5909 ( .A(n4834), .B(n4840), .Z(n5015) );
  XNOR U5910 ( .A(n4839), .B(n4831), .Z(n5016) );
  XNOR U5911 ( .A(n4830), .B(n4826), .Z(n5017) );
  XNOR U5912 ( .A(n4825), .B(n4821), .Z(n5018) );
  XNOR U5913 ( .A(n4820), .B(n4816), .Z(n5019) );
  XNOR U5914 ( .A(n4807), .B(n4806), .Z(n5020) );
  XOR U5915 ( .A(n5021), .B(n4805), .Z(n4806) );
  AND U5916 ( .A(b[35]), .B(a[12]), .Z(n5021) );
  XNOR U5917 ( .A(n4805), .B(n4811), .Z(n5022) );
  XNOR U5918 ( .A(n4810), .B(n4802), .Z(n5023) );
  XNOR U5919 ( .A(n4801), .B(n4797), .Z(n5024) );
  XNOR U5920 ( .A(n4796), .B(n4792), .Z(n5025) );
  XNOR U5921 ( .A(n4791), .B(n4787), .Z(n5026) );
  XNOR U5922 ( .A(n4778), .B(n4777), .Z(n5027) );
  XOR U5923 ( .A(n5028), .B(n4776), .Z(n4777) );
  AND U5924 ( .A(a[6]), .B(b[41]), .Z(n5028) );
  XNOR U5925 ( .A(n4776), .B(n4782), .Z(n5029) );
  XNOR U5926 ( .A(n4781), .B(n4773), .Z(n5030) );
  XNOR U5927 ( .A(n4772), .B(n4768), .Z(n5031) );
  XNOR U5928 ( .A(n4767), .B(n4763), .Z(n5032) );
  XNOR U5929 ( .A(n4762), .B(n4758), .Z(n5033) );
  XNOR U5930 ( .A(n5034), .B(n4757), .Z(n4758) );
  AND U5931 ( .A(a[0]), .B(b[47]), .Z(n5034) );
  XOR U5932 ( .A(n5035), .B(n4757), .Z(n4759) );
  XNOR U5933 ( .A(n5036), .B(n5037), .Z(n4757) );
  ANDN U5934 ( .B(n5038), .A(n5039), .Z(n5036) );
  AND U5935 ( .A(a[1]), .B(b[46]), .Z(n5035) );
  XNOR U5936 ( .A(n5040), .B(n4762), .Z(n4764) );
  XOR U5937 ( .A(n5041), .B(n5042), .Z(n4762) );
  ANDN U5938 ( .B(n5043), .A(n5044), .Z(n5041) );
  AND U5939 ( .A(a[2]), .B(b[45]), .Z(n5040) );
  XNOR U5940 ( .A(n5045), .B(n4767), .Z(n4769) );
  XOR U5941 ( .A(n5046), .B(n5047), .Z(n4767) );
  ANDN U5942 ( .B(n5048), .A(n5049), .Z(n5046) );
  AND U5943 ( .A(a[3]), .B(b[44]), .Z(n5045) );
  XNOR U5944 ( .A(n5050), .B(n4772), .Z(n4774) );
  XOR U5945 ( .A(n5051), .B(n5052), .Z(n4772) );
  ANDN U5946 ( .B(n5053), .A(n5054), .Z(n5051) );
  AND U5947 ( .A(a[4]), .B(b[43]), .Z(n5050) );
  XOR U5948 ( .A(n5055), .B(n5056), .Z(n4776) );
  AND U5949 ( .A(n5057), .B(n5058), .Z(n5055) );
  XNOR U5950 ( .A(n5059), .B(n4781), .Z(n4783) );
  XOR U5951 ( .A(n5060), .B(n5061), .Z(n4781) );
  ANDN U5952 ( .B(n5062), .A(n5063), .Z(n5060) );
  AND U5953 ( .A(a[5]), .B(b[42]), .Z(n5059) );
  XOR U5954 ( .A(n5064), .B(n4786), .Z(n4788) );
  XOR U5955 ( .A(n5065), .B(n5066), .Z(n4786) );
  ANDN U5956 ( .B(n5067), .A(n5068), .Z(n5065) );
  AND U5957 ( .A(a[7]), .B(b[40]), .Z(n5064) );
  XNOR U5958 ( .A(n5069), .B(n4791), .Z(n4793) );
  XOR U5959 ( .A(n5070), .B(n5071), .Z(n4791) );
  ANDN U5960 ( .B(n5072), .A(n5073), .Z(n5070) );
  AND U5961 ( .A(a[8]), .B(b[39]), .Z(n5069) );
  XNOR U5962 ( .A(n5074), .B(n4796), .Z(n4798) );
  XOR U5963 ( .A(n5075), .B(n5076), .Z(n4796) );
  ANDN U5964 ( .B(n5077), .A(n5078), .Z(n5075) );
  AND U5965 ( .A(a[9]), .B(b[38]), .Z(n5074) );
  XNOR U5966 ( .A(n5079), .B(n4801), .Z(n4803) );
  XOR U5967 ( .A(n5080), .B(n5081), .Z(n4801) );
  ANDN U5968 ( .B(n5082), .A(n5083), .Z(n5080) );
  AND U5969 ( .A(b[37]), .B(a[10]), .Z(n5079) );
  XOR U5970 ( .A(n5084), .B(n5085), .Z(n4805) );
  AND U5971 ( .A(n5086), .B(n5087), .Z(n5084) );
  XNOR U5972 ( .A(n5088), .B(n4810), .Z(n4812) );
  XOR U5973 ( .A(n5089), .B(n5090), .Z(n4810) );
  ANDN U5974 ( .B(n5091), .A(n5092), .Z(n5089) );
  AND U5975 ( .A(b[36]), .B(a[11]), .Z(n5088) );
  XOR U5976 ( .A(n5093), .B(n4815), .Z(n4817) );
  XOR U5977 ( .A(n5094), .B(n5095), .Z(n4815) );
  ANDN U5978 ( .B(n5096), .A(n5097), .Z(n5094) );
  AND U5979 ( .A(b[34]), .B(a[13]), .Z(n5093) );
  XNOR U5980 ( .A(n5098), .B(n4820), .Z(n4822) );
  XOR U5981 ( .A(n5099), .B(n5100), .Z(n4820) );
  ANDN U5982 ( .B(n5101), .A(n5102), .Z(n5099) );
  AND U5983 ( .A(a[14]), .B(b[33]), .Z(n5098) );
  XNOR U5984 ( .A(n5103), .B(n4825), .Z(n4827) );
  XOR U5985 ( .A(n5104), .B(n5105), .Z(n4825) );
  ANDN U5986 ( .B(n5106), .A(n5107), .Z(n5104) );
  AND U5987 ( .A(b[32]), .B(a[15]), .Z(n5103) );
  XNOR U5988 ( .A(n5108), .B(n4830), .Z(n4832) );
  XOR U5989 ( .A(n5109), .B(n5110), .Z(n4830) );
  ANDN U5990 ( .B(n5111), .A(n5112), .Z(n5109) );
  AND U5991 ( .A(b[31]), .B(a[16]), .Z(n5108) );
  XOR U5992 ( .A(n5113), .B(n5114), .Z(n4834) );
  AND U5993 ( .A(n5115), .B(n5116), .Z(n5113) );
  XNOR U5994 ( .A(n5117), .B(n4839), .Z(n4841) );
  XOR U5995 ( .A(n5118), .B(n5119), .Z(n4839) );
  ANDN U5996 ( .B(n5120), .A(n5121), .Z(n5118) );
  AND U5997 ( .A(b[30]), .B(a[17]), .Z(n5117) );
  IV U5998 ( .A(n4844), .Z(n5012) );
  XOR U5999 ( .A(n5122), .B(n4844), .Z(n4846) );
  XOR U6000 ( .A(n5123), .B(n5124), .Z(n4844) );
  ANDN U6001 ( .B(n5125), .A(n5126), .Z(n5123) );
  AND U6002 ( .A(b[28]), .B(a[19]), .Z(n5122) );
  XNOR U6003 ( .A(n5127), .B(n4849), .Z(n4851) );
  XOR U6004 ( .A(n5128), .B(n5129), .Z(n4849) );
  ANDN U6005 ( .B(n5130), .A(n5131), .Z(n5128) );
  AND U6006 ( .A(a[20]), .B(b[27]), .Z(n5127) );
  XNOR U6007 ( .A(n5132), .B(n4854), .Z(n4856) );
  XOR U6008 ( .A(n5133), .B(n5134), .Z(n4854) );
  ANDN U6009 ( .B(n5135), .A(n5136), .Z(n5133) );
  AND U6010 ( .A(b[26]), .B(a[21]), .Z(n5132) );
  XNOR U6011 ( .A(n5137), .B(n4859), .Z(n4861) );
  XOR U6012 ( .A(n5138), .B(n5139), .Z(n4859) );
  ANDN U6013 ( .B(n5140), .A(n5141), .Z(n5138) );
  AND U6014 ( .A(b[25]), .B(a[22]), .Z(n5137) );
  XOR U6015 ( .A(n5142), .B(n5143), .Z(n4863) );
  AND U6016 ( .A(n5144), .B(n5145), .Z(n5142) );
  XNOR U6017 ( .A(n5146), .B(n4868), .Z(n4870) );
  XOR U6018 ( .A(n5147), .B(n5148), .Z(n4868) );
  ANDN U6019 ( .B(n5149), .A(n5150), .Z(n5147) );
  AND U6020 ( .A(b[24]), .B(a[23]), .Z(n5146) );
  XOR U6021 ( .A(n5151), .B(n4873), .Z(n4875) );
  XOR U6022 ( .A(n5152), .B(n5153), .Z(n4873) );
  ANDN U6023 ( .B(n5154), .A(n5155), .Z(n5152) );
  AND U6024 ( .A(b[22]), .B(a[25]), .Z(n5151) );
  XNOR U6025 ( .A(n5156), .B(n4878), .Z(n4880) );
  XOR U6026 ( .A(n5157), .B(n5158), .Z(n4878) );
  ANDN U6027 ( .B(n5159), .A(n5160), .Z(n5157) );
  AND U6028 ( .A(a[26]), .B(b[21]), .Z(n5156) );
  XNOR U6029 ( .A(n5161), .B(n4883), .Z(n4885) );
  XOR U6030 ( .A(n5162), .B(n5163), .Z(n4883) );
  ANDN U6031 ( .B(n5164), .A(n5165), .Z(n5162) );
  AND U6032 ( .A(b[20]), .B(a[27]), .Z(n5161) );
  XNOR U6033 ( .A(n5166), .B(n4888), .Z(n4890) );
  XOR U6034 ( .A(n5167), .B(n5168), .Z(n4888) );
  ANDN U6035 ( .B(n5169), .A(n5170), .Z(n5167) );
  AND U6036 ( .A(b[19]), .B(a[28]), .Z(n5166) );
  XOR U6037 ( .A(n5171), .B(n5172), .Z(n4892) );
  AND U6038 ( .A(n5173), .B(n5174), .Z(n5171) );
  XNOR U6039 ( .A(n5175), .B(n4897), .Z(n4899) );
  XOR U6040 ( .A(n5176), .B(n5177), .Z(n4897) );
  ANDN U6041 ( .B(n5178), .A(n5179), .Z(n5176) );
  AND U6042 ( .A(b[18]), .B(a[29]), .Z(n5175) );
  XOR U6043 ( .A(n5180), .B(n4902), .Z(n4904) );
  XOR U6044 ( .A(n5181), .B(n5182), .Z(n4902) );
  ANDN U6045 ( .B(n5183), .A(n5184), .Z(n5181) );
  AND U6046 ( .A(b[16]), .B(a[31]), .Z(n5180) );
  XNOR U6047 ( .A(n5185), .B(n4907), .Z(n4909) );
  XOR U6048 ( .A(n5186), .B(n5187), .Z(n4907) );
  ANDN U6049 ( .B(n5188), .A(n5189), .Z(n5186) );
  AND U6050 ( .A(a[32]), .B(b[15]), .Z(n5185) );
  XNOR U6051 ( .A(n5190), .B(n4912), .Z(n4914) );
  XOR U6052 ( .A(n5191), .B(n5192), .Z(n4912) );
  ANDN U6053 ( .B(n5193), .A(n5194), .Z(n5191) );
  AND U6054 ( .A(b[14]), .B(a[33]), .Z(n5190) );
  XNOR U6055 ( .A(n5195), .B(n4917), .Z(n4919) );
  XOR U6056 ( .A(n5196), .B(n5197), .Z(n4917) );
  ANDN U6057 ( .B(n5198), .A(n5199), .Z(n5196) );
  AND U6058 ( .A(b[13]), .B(a[34]), .Z(n5195) );
  XOR U6059 ( .A(n5200), .B(n5201), .Z(n4921) );
  AND U6060 ( .A(n5202), .B(n5203), .Z(n5200) );
  XNOR U6061 ( .A(n5204), .B(n4926), .Z(n4928) );
  XOR U6062 ( .A(n5205), .B(n5206), .Z(n4926) );
  ANDN U6063 ( .B(n5207), .A(n5208), .Z(n5205) );
  AND U6064 ( .A(b[12]), .B(a[35]), .Z(n5204) );
  XOR U6065 ( .A(n5209), .B(n4931), .Z(n4933) );
  XOR U6066 ( .A(n5210), .B(n5211), .Z(n4931) );
  ANDN U6067 ( .B(n5212), .A(n5213), .Z(n5210) );
  AND U6068 ( .A(b[10]), .B(a[37]), .Z(n5209) );
  XNOR U6069 ( .A(n5214), .B(n4936), .Z(n4938) );
  XOR U6070 ( .A(n5215), .B(n5216), .Z(n4936) );
  ANDN U6071 ( .B(n5217), .A(n5218), .Z(n5215) );
  AND U6072 ( .A(b[9]), .B(a[38]), .Z(n5214) );
  XNOR U6073 ( .A(n5219), .B(n4941), .Z(n4943) );
  XOR U6074 ( .A(n5220), .B(n5221), .Z(n4941) );
  ANDN U6075 ( .B(n5222), .A(n5223), .Z(n5220) );
  AND U6076 ( .A(b[8]), .B(a[39]), .Z(n5219) );
  XNOR U6077 ( .A(n5224), .B(n4946), .Z(n4948) );
  XOR U6078 ( .A(n5225), .B(n5226), .Z(n4946) );
  ANDN U6079 ( .B(n5227), .A(n5228), .Z(n5225) );
  AND U6080 ( .A(b[7]), .B(a[40]), .Z(n5224) );
  XNOR U6081 ( .A(n5229), .B(n4951), .Z(n4953) );
  XOR U6082 ( .A(n5230), .B(n5231), .Z(n4951) );
  ANDN U6083 ( .B(n5232), .A(n5233), .Z(n5230) );
  AND U6084 ( .A(b[6]), .B(a[41]), .Z(n5229) );
  XNOR U6085 ( .A(n5234), .B(n4956), .Z(n4958) );
  XOR U6086 ( .A(n5235), .B(n5236), .Z(n4956) );
  ANDN U6087 ( .B(n5237), .A(n5238), .Z(n5235) );
  AND U6088 ( .A(b[5]), .B(a[42]), .Z(n5234) );
  XNOR U6089 ( .A(n5239), .B(n4961), .Z(n4963) );
  XOR U6090 ( .A(n5240), .B(n5241), .Z(n4961) );
  ANDN U6091 ( .B(n5242), .A(n5243), .Z(n5240) );
  AND U6092 ( .A(b[4]), .B(a[43]), .Z(n5239) );
  XNOR U6093 ( .A(n5244), .B(n5245), .Z(n4975) );
  NANDN U6094 ( .A(n5246), .B(n5247), .Z(n5245) );
  XNOR U6095 ( .A(n5248), .B(n4966), .Z(n4968) );
  XNOR U6096 ( .A(n5249), .B(n5250), .Z(n4966) );
  AND U6097 ( .A(n5251), .B(n5252), .Z(n5249) );
  AND U6098 ( .A(b[3]), .B(a[44]), .Z(n5248) );
  NAND U6099 ( .A(a[47]), .B(b[0]), .Z(n4702) );
  XNOR U6100 ( .A(n4981), .B(n4982), .Z(c[46]) );
  XNOR U6101 ( .A(n5246), .B(n5247), .Z(n4982) );
  XOR U6102 ( .A(n5244), .B(n5253), .Z(n5247) );
  NAND U6103 ( .A(b[1]), .B(a[45]), .Z(n5253) );
  XOR U6104 ( .A(n5252), .B(n5254), .Z(n5246) );
  XOR U6105 ( .A(n5244), .B(n5251), .Z(n5254) );
  XNOR U6106 ( .A(n5255), .B(n5250), .Z(n5251) );
  AND U6107 ( .A(b[2]), .B(a[44]), .Z(n5255) );
  NANDN U6108 ( .A(n5256), .B(n5257), .Z(n5244) );
  XOR U6109 ( .A(n5250), .B(n5242), .Z(n5258) );
  XNOR U6110 ( .A(n5241), .B(n5237), .Z(n5259) );
  XNOR U6111 ( .A(n5236), .B(n5232), .Z(n5260) );
  XNOR U6112 ( .A(n5231), .B(n5227), .Z(n5261) );
  XNOR U6113 ( .A(n5226), .B(n5222), .Z(n5262) );
  XNOR U6114 ( .A(n5221), .B(n5217), .Z(n5263) );
  XNOR U6115 ( .A(n5216), .B(n5212), .Z(n5264) );
  XNOR U6116 ( .A(n5203), .B(n5202), .Z(n5265) );
  XOR U6117 ( .A(n5266), .B(n5201), .Z(n5202) );
  AND U6118 ( .A(b[10]), .B(a[36]), .Z(n5266) );
  XNOR U6119 ( .A(n5201), .B(n5207), .Z(n5267) );
  XNOR U6120 ( .A(n5206), .B(n5198), .Z(n5268) );
  XNOR U6121 ( .A(n5197), .B(n5193), .Z(n5269) );
  XNOR U6122 ( .A(n5192), .B(n5188), .Z(n5270) );
  XNOR U6123 ( .A(n5187), .B(n5183), .Z(n5271) );
  XNOR U6124 ( .A(n5174), .B(n5173), .Z(n5272) );
  XOR U6125 ( .A(n5273), .B(n5172), .Z(n5173) );
  AND U6126 ( .A(b[16]), .B(a[30]), .Z(n5273) );
  XNOR U6127 ( .A(n5172), .B(n5178), .Z(n5274) );
  XNOR U6128 ( .A(n5177), .B(n5169), .Z(n5275) );
  XNOR U6129 ( .A(n5168), .B(n5164), .Z(n5276) );
  XNOR U6130 ( .A(n5163), .B(n5159), .Z(n5277) );
  XNOR U6131 ( .A(n5158), .B(n5154), .Z(n5278) );
  XNOR U6132 ( .A(n5145), .B(n5144), .Z(n5279) );
  XOR U6133 ( .A(n5280), .B(n5143), .Z(n5144) );
  AND U6134 ( .A(b[22]), .B(a[24]), .Z(n5280) );
  XNOR U6135 ( .A(n5143), .B(n5149), .Z(n5281) );
  XNOR U6136 ( .A(n5148), .B(n5140), .Z(n5282) );
  XNOR U6137 ( .A(n5139), .B(n5135), .Z(n5283) );
  XNOR U6138 ( .A(n5134), .B(n5130), .Z(n5284) );
  XNOR U6139 ( .A(n5129), .B(n5125), .Z(n5285) );
  XNOR U6140 ( .A(n5116), .B(n5115), .Z(n5286) );
  XOR U6141 ( .A(n5287), .B(n5114), .Z(n5115) );
  AND U6142 ( .A(b[28]), .B(a[18]), .Z(n5287) );
  XNOR U6143 ( .A(n5114), .B(n5120), .Z(n5288) );
  XNOR U6144 ( .A(n5119), .B(n5111), .Z(n5289) );
  XNOR U6145 ( .A(n5110), .B(n5106), .Z(n5290) );
  XNOR U6146 ( .A(n5105), .B(n5101), .Z(n5291) );
  XNOR U6147 ( .A(n5100), .B(n5096), .Z(n5292) );
  XNOR U6148 ( .A(n5087), .B(n5086), .Z(n5293) );
  XOR U6149 ( .A(n5294), .B(n5085), .Z(n5086) );
  AND U6150 ( .A(b[34]), .B(a[12]), .Z(n5294) );
  XNOR U6151 ( .A(n5085), .B(n5091), .Z(n5295) );
  XNOR U6152 ( .A(n5090), .B(n5082), .Z(n5296) );
  XNOR U6153 ( .A(n5081), .B(n5077), .Z(n5297) );
  XNOR U6154 ( .A(n5076), .B(n5072), .Z(n5298) );
  XNOR U6155 ( .A(n5071), .B(n5067), .Z(n5299) );
  XNOR U6156 ( .A(n5058), .B(n5057), .Z(n5300) );
  XOR U6157 ( .A(n5301), .B(n5056), .Z(n5057) );
  AND U6158 ( .A(a[6]), .B(b[40]), .Z(n5301) );
  XNOR U6159 ( .A(n5056), .B(n5062), .Z(n5302) );
  XNOR U6160 ( .A(n5061), .B(n5053), .Z(n5303) );
  XNOR U6161 ( .A(n5052), .B(n5048), .Z(n5304) );
  XNOR U6162 ( .A(n5047), .B(n5043), .Z(n5305) );
  XNOR U6163 ( .A(n5042), .B(n5038), .Z(n5306) );
  XOR U6164 ( .A(n5307), .B(n5037), .Z(n5038) );
  AND U6165 ( .A(a[0]), .B(b[46]), .Z(n5307) );
  XNOR U6166 ( .A(n5308), .B(n5037), .Z(n5039) );
  XNOR U6167 ( .A(n5309), .B(n5310), .Z(n5037) );
  ANDN U6168 ( .B(n5311), .A(n5312), .Z(n5309) );
  AND U6169 ( .A(a[1]), .B(b[45]), .Z(n5308) );
  XNOR U6170 ( .A(n5313), .B(n5042), .Z(n5044) );
  XOR U6171 ( .A(n5314), .B(n5315), .Z(n5042) );
  ANDN U6172 ( .B(n5316), .A(n5317), .Z(n5314) );
  AND U6173 ( .A(a[2]), .B(b[44]), .Z(n5313) );
  XNOR U6174 ( .A(n5318), .B(n5047), .Z(n5049) );
  XOR U6175 ( .A(n5319), .B(n5320), .Z(n5047) );
  ANDN U6176 ( .B(n5321), .A(n5322), .Z(n5319) );
  AND U6177 ( .A(a[3]), .B(b[43]), .Z(n5318) );
  XNOR U6178 ( .A(n5323), .B(n5052), .Z(n5054) );
  XOR U6179 ( .A(n5324), .B(n5325), .Z(n5052) );
  ANDN U6180 ( .B(n5326), .A(n5327), .Z(n5324) );
  AND U6181 ( .A(a[4]), .B(b[42]), .Z(n5323) );
  XOR U6182 ( .A(n5328), .B(n5329), .Z(n5056) );
  AND U6183 ( .A(n5330), .B(n5331), .Z(n5328) );
  XNOR U6184 ( .A(n5332), .B(n5061), .Z(n5063) );
  XOR U6185 ( .A(n5333), .B(n5334), .Z(n5061) );
  ANDN U6186 ( .B(n5335), .A(n5336), .Z(n5333) );
  AND U6187 ( .A(a[5]), .B(b[41]), .Z(n5332) );
  XOR U6188 ( .A(n5337), .B(n5066), .Z(n5068) );
  XOR U6189 ( .A(n5338), .B(n5339), .Z(n5066) );
  ANDN U6190 ( .B(n5340), .A(n5341), .Z(n5338) );
  AND U6191 ( .A(a[7]), .B(b[39]), .Z(n5337) );
  XNOR U6192 ( .A(n5342), .B(n5071), .Z(n5073) );
  XOR U6193 ( .A(n5343), .B(n5344), .Z(n5071) );
  ANDN U6194 ( .B(n5345), .A(n5346), .Z(n5343) );
  AND U6195 ( .A(a[8]), .B(b[38]), .Z(n5342) );
  XNOR U6196 ( .A(n5347), .B(n5076), .Z(n5078) );
  XOR U6197 ( .A(n5348), .B(n5349), .Z(n5076) );
  ANDN U6198 ( .B(n5350), .A(n5351), .Z(n5348) );
  AND U6199 ( .A(a[9]), .B(b[37]), .Z(n5347) );
  XNOR U6200 ( .A(n5352), .B(n5081), .Z(n5083) );
  XOR U6201 ( .A(n5353), .B(n5354), .Z(n5081) );
  ANDN U6202 ( .B(n5355), .A(n5356), .Z(n5353) );
  AND U6203 ( .A(b[36]), .B(a[10]), .Z(n5352) );
  XOR U6204 ( .A(n5357), .B(n5358), .Z(n5085) );
  AND U6205 ( .A(n5359), .B(n5360), .Z(n5357) );
  XNOR U6206 ( .A(n5361), .B(n5090), .Z(n5092) );
  XOR U6207 ( .A(n5362), .B(n5363), .Z(n5090) );
  ANDN U6208 ( .B(n5364), .A(n5365), .Z(n5362) );
  AND U6209 ( .A(b[35]), .B(a[11]), .Z(n5361) );
  XOR U6210 ( .A(n5366), .B(n5095), .Z(n5097) );
  XOR U6211 ( .A(n5367), .B(n5368), .Z(n5095) );
  ANDN U6212 ( .B(n5369), .A(n5370), .Z(n5367) );
  AND U6213 ( .A(a[13]), .B(b[33]), .Z(n5366) );
  XNOR U6214 ( .A(n5371), .B(n5100), .Z(n5102) );
  XOR U6215 ( .A(n5372), .B(n5373), .Z(n5100) );
  ANDN U6216 ( .B(n5374), .A(n5375), .Z(n5372) );
  AND U6217 ( .A(b[32]), .B(a[14]), .Z(n5371) );
  XNOR U6218 ( .A(n5376), .B(n5105), .Z(n5107) );
  XOR U6219 ( .A(n5377), .B(n5378), .Z(n5105) );
  ANDN U6220 ( .B(n5379), .A(n5380), .Z(n5377) );
  AND U6221 ( .A(b[31]), .B(a[15]), .Z(n5376) );
  XNOR U6222 ( .A(n5381), .B(n5110), .Z(n5112) );
  XOR U6223 ( .A(n5382), .B(n5383), .Z(n5110) );
  ANDN U6224 ( .B(n5384), .A(n5385), .Z(n5382) );
  AND U6225 ( .A(b[30]), .B(a[16]), .Z(n5381) );
  XOR U6226 ( .A(n5386), .B(n5387), .Z(n5114) );
  AND U6227 ( .A(n5388), .B(n5389), .Z(n5386) );
  XNOR U6228 ( .A(n5390), .B(n5119), .Z(n5121) );
  XOR U6229 ( .A(n5391), .B(n5392), .Z(n5119) );
  ANDN U6230 ( .B(n5393), .A(n5394), .Z(n5391) );
  AND U6231 ( .A(b[29]), .B(a[17]), .Z(n5390) );
  XOR U6232 ( .A(n5395), .B(n5124), .Z(n5126) );
  XOR U6233 ( .A(n5396), .B(n5397), .Z(n5124) );
  ANDN U6234 ( .B(n5398), .A(n5399), .Z(n5396) );
  AND U6235 ( .A(a[19]), .B(b[27]), .Z(n5395) );
  XNOR U6236 ( .A(n5400), .B(n5129), .Z(n5131) );
  XOR U6237 ( .A(n5401), .B(n5402), .Z(n5129) );
  ANDN U6238 ( .B(n5403), .A(n5404), .Z(n5401) );
  AND U6239 ( .A(b[26]), .B(a[20]), .Z(n5400) );
  XNOR U6240 ( .A(n5405), .B(n5134), .Z(n5136) );
  XOR U6241 ( .A(n5406), .B(n5407), .Z(n5134) );
  ANDN U6242 ( .B(n5408), .A(n5409), .Z(n5406) );
  AND U6243 ( .A(b[25]), .B(a[21]), .Z(n5405) );
  XNOR U6244 ( .A(n5410), .B(n5139), .Z(n5141) );
  XOR U6245 ( .A(n5411), .B(n5412), .Z(n5139) );
  ANDN U6246 ( .B(n5413), .A(n5414), .Z(n5411) );
  AND U6247 ( .A(b[24]), .B(a[22]), .Z(n5410) );
  XOR U6248 ( .A(n5415), .B(n5416), .Z(n5143) );
  AND U6249 ( .A(n5417), .B(n5418), .Z(n5415) );
  XNOR U6250 ( .A(n5419), .B(n5148), .Z(n5150) );
  XOR U6251 ( .A(n5420), .B(n5421), .Z(n5148) );
  ANDN U6252 ( .B(n5422), .A(n5423), .Z(n5420) );
  AND U6253 ( .A(b[23]), .B(a[23]), .Z(n5419) );
  XOR U6254 ( .A(n5424), .B(n5153), .Z(n5155) );
  XOR U6255 ( .A(n5425), .B(n5426), .Z(n5153) );
  ANDN U6256 ( .B(n5427), .A(n5428), .Z(n5425) );
  AND U6257 ( .A(a[25]), .B(b[21]), .Z(n5424) );
  XNOR U6258 ( .A(n5429), .B(n5158), .Z(n5160) );
  XOR U6259 ( .A(n5430), .B(n5431), .Z(n5158) );
  ANDN U6260 ( .B(n5432), .A(n5433), .Z(n5430) );
  AND U6261 ( .A(b[20]), .B(a[26]), .Z(n5429) );
  XNOR U6262 ( .A(n5434), .B(n5163), .Z(n5165) );
  XOR U6263 ( .A(n5435), .B(n5436), .Z(n5163) );
  ANDN U6264 ( .B(n5437), .A(n5438), .Z(n5435) );
  AND U6265 ( .A(b[19]), .B(a[27]), .Z(n5434) );
  XNOR U6266 ( .A(n5439), .B(n5168), .Z(n5170) );
  XOR U6267 ( .A(n5440), .B(n5441), .Z(n5168) );
  ANDN U6268 ( .B(n5442), .A(n5443), .Z(n5440) );
  AND U6269 ( .A(b[18]), .B(a[28]), .Z(n5439) );
  XOR U6270 ( .A(n5444), .B(n5445), .Z(n5172) );
  AND U6271 ( .A(n5446), .B(n5447), .Z(n5444) );
  XNOR U6272 ( .A(n5448), .B(n5177), .Z(n5179) );
  XOR U6273 ( .A(n5449), .B(n5450), .Z(n5177) );
  ANDN U6274 ( .B(n5451), .A(n5452), .Z(n5449) );
  AND U6275 ( .A(b[17]), .B(a[29]), .Z(n5448) );
  XOR U6276 ( .A(n5453), .B(n5182), .Z(n5184) );
  XOR U6277 ( .A(n5454), .B(n5455), .Z(n5182) );
  ANDN U6278 ( .B(n5456), .A(n5457), .Z(n5454) );
  AND U6279 ( .A(a[31]), .B(b[15]), .Z(n5453) );
  XNOR U6280 ( .A(n5458), .B(n5187), .Z(n5189) );
  XOR U6281 ( .A(n5459), .B(n5460), .Z(n5187) );
  ANDN U6282 ( .B(n5461), .A(n5462), .Z(n5459) );
  AND U6283 ( .A(b[14]), .B(a[32]), .Z(n5458) );
  XNOR U6284 ( .A(n5463), .B(n5192), .Z(n5194) );
  XOR U6285 ( .A(n5464), .B(n5465), .Z(n5192) );
  ANDN U6286 ( .B(n5466), .A(n5467), .Z(n5464) );
  AND U6287 ( .A(b[13]), .B(a[33]), .Z(n5463) );
  XNOR U6288 ( .A(n5468), .B(n5197), .Z(n5199) );
  XOR U6289 ( .A(n5469), .B(n5470), .Z(n5197) );
  ANDN U6290 ( .B(n5471), .A(n5472), .Z(n5469) );
  AND U6291 ( .A(b[12]), .B(a[34]), .Z(n5468) );
  XOR U6292 ( .A(n5473), .B(n5474), .Z(n5201) );
  AND U6293 ( .A(n5475), .B(n5476), .Z(n5473) );
  XNOR U6294 ( .A(n5477), .B(n5206), .Z(n5208) );
  XOR U6295 ( .A(n5478), .B(n5479), .Z(n5206) );
  ANDN U6296 ( .B(n5480), .A(n5481), .Z(n5478) );
  AND U6297 ( .A(b[11]), .B(a[35]), .Z(n5477) );
  XOR U6298 ( .A(n5482), .B(n5211), .Z(n5213) );
  XOR U6299 ( .A(n5483), .B(n5484), .Z(n5211) );
  ANDN U6300 ( .B(n5485), .A(n5486), .Z(n5483) );
  AND U6301 ( .A(b[9]), .B(a[37]), .Z(n5482) );
  XNOR U6302 ( .A(n5487), .B(n5216), .Z(n5218) );
  XOR U6303 ( .A(n5488), .B(n5489), .Z(n5216) );
  ANDN U6304 ( .B(n5490), .A(n5491), .Z(n5488) );
  AND U6305 ( .A(b[8]), .B(a[38]), .Z(n5487) );
  XNOR U6306 ( .A(n5492), .B(n5221), .Z(n5223) );
  XOR U6307 ( .A(n5493), .B(n5494), .Z(n5221) );
  ANDN U6308 ( .B(n5495), .A(n5496), .Z(n5493) );
  AND U6309 ( .A(b[7]), .B(a[39]), .Z(n5492) );
  XNOR U6310 ( .A(n5497), .B(n5226), .Z(n5228) );
  XOR U6311 ( .A(n5498), .B(n5499), .Z(n5226) );
  ANDN U6312 ( .B(n5500), .A(n5501), .Z(n5498) );
  AND U6313 ( .A(b[6]), .B(a[40]), .Z(n5497) );
  XNOR U6314 ( .A(n5502), .B(n5231), .Z(n5233) );
  XOR U6315 ( .A(n5503), .B(n5504), .Z(n5231) );
  ANDN U6316 ( .B(n5505), .A(n5506), .Z(n5503) );
  AND U6317 ( .A(b[5]), .B(a[41]), .Z(n5502) );
  XNOR U6318 ( .A(n5507), .B(n5236), .Z(n5238) );
  XOR U6319 ( .A(n5508), .B(n5509), .Z(n5236) );
  ANDN U6320 ( .B(n5510), .A(n5511), .Z(n5508) );
  AND U6321 ( .A(b[4]), .B(a[42]), .Z(n5507) );
  XNOR U6322 ( .A(n5512), .B(n5513), .Z(n5250) );
  NANDN U6323 ( .A(n5514), .B(n5515), .Z(n5513) );
  XNOR U6324 ( .A(n5516), .B(n5241), .Z(n5243) );
  XNOR U6325 ( .A(n5517), .B(n5518), .Z(n5241) );
  AND U6326 ( .A(n5519), .B(n5520), .Z(n5517) );
  AND U6327 ( .A(b[3]), .B(a[43]), .Z(n5516) );
  NAND U6328 ( .A(a[46]), .B(b[0]), .Z(n4981) );
  XNOR U6329 ( .A(n5256), .B(n5257), .Z(c[45]) );
  XNOR U6330 ( .A(n5514), .B(n5515), .Z(n5257) );
  XOR U6331 ( .A(n5512), .B(n5521), .Z(n5515) );
  NAND U6332 ( .A(b[1]), .B(a[44]), .Z(n5521) );
  XOR U6333 ( .A(n5520), .B(n5522), .Z(n5514) );
  XOR U6334 ( .A(n5512), .B(n5519), .Z(n5522) );
  XNOR U6335 ( .A(n5523), .B(n5518), .Z(n5519) );
  AND U6336 ( .A(b[2]), .B(a[43]), .Z(n5523) );
  NANDN U6337 ( .A(n5524), .B(n5525), .Z(n5512) );
  XOR U6338 ( .A(n5518), .B(n5510), .Z(n5526) );
  XNOR U6339 ( .A(n5509), .B(n5505), .Z(n5527) );
  XNOR U6340 ( .A(n5504), .B(n5500), .Z(n5528) );
  XNOR U6341 ( .A(n5499), .B(n5495), .Z(n5529) );
  XNOR U6342 ( .A(n5494), .B(n5490), .Z(n5530) );
  XNOR U6343 ( .A(n5489), .B(n5485), .Z(n5531) );
  XNOR U6344 ( .A(n5476), .B(n5475), .Z(n5532) );
  XOR U6345 ( .A(n5533), .B(n5474), .Z(n5475) );
  AND U6346 ( .A(b[9]), .B(a[36]), .Z(n5533) );
  XNOR U6347 ( .A(n5474), .B(n5480), .Z(n5534) );
  XNOR U6348 ( .A(n5479), .B(n5471), .Z(n5535) );
  XNOR U6349 ( .A(n5470), .B(n5466), .Z(n5536) );
  XNOR U6350 ( .A(n5465), .B(n5461), .Z(n5537) );
  XNOR U6351 ( .A(n5460), .B(n5456), .Z(n5538) );
  XNOR U6352 ( .A(n5447), .B(n5446), .Z(n5539) );
  XOR U6353 ( .A(n5540), .B(n5445), .Z(n5446) );
  AND U6354 ( .A(b[15]), .B(a[30]), .Z(n5540) );
  XNOR U6355 ( .A(n5445), .B(n5451), .Z(n5541) );
  XNOR U6356 ( .A(n5450), .B(n5442), .Z(n5542) );
  XNOR U6357 ( .A(n5441), .B(n5437), .Z(n5543) );
  XNOR U6358 ( .A(n5436), .B(n5432), .Z(n5544) );
  XNOR U6359 ( .A(n5431), .B(n5427), .Z(n5545) );
  XNOR U6360 ( .A(n5418), .B(n5417), .Z(n5546) );
  XOR U6361 ( .A(n5547), .B(n5416), .Z(n5417) );
  AND U6362 ( .A(b[21]), .B(a[24]), .Z(n5547) );
  XNOR U6363 ( .A(n5416), .B(n5422), .Z(n5548) );
  XNOR U6364 ( .A(n5421), .B(n5413), .Z(n5549) );
  XNOR U6365 ( .A(n5412), .B(n5408), .Z(n5550) );
  XNOR U6366 ( .A(n5407), .B(n5403), .Z(n5551) );
  XNOR U6367 ( .A(n5402), .B(n5398), .Z(n5552) );
  XNOR U6368 ( .A(n5389), .B(n5388), .Z(n5553) );
  XOR U6369 ( .A(n5554), .B(n5387), .Z(n5388) );
  AND U6370 ( .A(b[27]), .B(a[18]), .Z(n5554) );
  XNOR U6371 ( .A(n5387), .B(n5393), .Z(n5555) );
  XNOR U6372 ( .A(n5392), .B(n5384), .Z(n5556) );
  XNOR U6373 ( .A(n5383), .B(n5379), .Z(n5557) );
  XNOR U6374 ( .A(n5378), .B(n5374), .Z(n5558) );
  XNOR U6375 ( .A(n5373), .B(n5369), .Z(n5559) );
  XNOR U6376 ( .A(n5360), .B(n5359), .Z(n5560) );
  XOR U6377 ( .A(n5561), .B(n5358), .Z(n5359) );
  AND U6378 ( .A(b[33]), .B(a[12]), .Z(n5561) );
  XNOR U6379 ( .A(n5358), .B(n5364), .Z(n5562) );
  XNOR U6380 ( .A(n5363), .B(n5355), .Z(n5563) );
  XNOR U6381 ( .A(n5354), .B(n5350), .Z(n5564) );
  XNOR U6382 ( .A(n5349), .B(n5345), .Z(n5565) );
  XNOR U6383 ( .A(n5344), .B(n5340), .Z(n5566) );
  XNOR U6384 ( .A(n5331), .B(n5330), .Z(n5567) );
  XOR U6385 ( .A(n5568), .B(n5329), .Z(n5330) );
  AND U6386 ( .A(a[6]), .B(b[39]), .Z(n5568) );
  XNOR U6387 ( .A(n5329), .B(n5335), .Z(n5569) );
  XNOR U6388 ( .A(n5334), .B(n5326), .Z(n5570) );
  XNOR U6389 ( .A(n5325), .B(n5321), .Z(n5571) );
  XNOR U6390 ( .A(n5320), .B(n5316), .Z(n5572) );
  XNOR U6391 ( .A(n5315), .B(n5311), .Z(n5573) );
  XNOR U6392 ( .A(n5574), .B(n5310), .Z(n5311) );
  AND U6393 ( .A(a[0]), .B(b[45]), .Z(n5574) );
  XOR U6394 ( .A(n5575), .B(n5310), .Z(n5312) );
  XNOR U6395 ( .A(n5576), .B(n5577), .Z(n5310) );
  ANDN U6396 ( .B(n5578), .A(n5579), .Z(n5576) );
  AND U6397 ( .A(a[1]), .B(b[44]), .Z(n5575) );
  XNOR U6398 ( .A(n5580), .B(n5315), .Z(n5317) );
  XOR U6399 ( .A(n5581), .B(n5582), .Z(n5315) );
  ANDN U6400 ( .B(n5583), .A(n5584), .Z(n5581) );
  AND U6401 ( .A(a[2]), .B(b[43]), .Z(n5580) );
  XNOR U6402 ( .A(n5585), .B(n5320), .Z(n5322) );
  XOR U6403 ( .A(n5586), .B(n5587), .Z(n5320) );
  ANDN U6404 ( .B(n5588), .A(n5589), .Z(n5586) );
  AND U6405 ( .A(a[3]), .B(b[42]), .Z(n5585) );
  XNOR U6406 ( .A(n5590), .B(n5325), .Z(n5327) );
  XOR U6407 ( .A(n5591), .B(n5592), .Z(n5325) );
  ANDN U6408 ( .B(n5593), .A(n5594), .Z(n5591) );
  AND U6409 ( .A(a[4]), .B(b[41]), .Z(n5590) );
  XOR U6410 ( .A(n5595), .B(n5596), .Z(n5329) );
  AND U6411 ( .A(n5597), .B(n5598), .Z(n5595) );
  XNOR U6412 ( .A(n5599), .B(n5334), .Z(n5336) );
  XOR U6413 ( .A(n5600), .B(n5601), .Z(n5334) );
  ANDN U6414 ( .B(n5602), .A(n5603), .Z(n5600) );
  AND U6415 ( .A(a[5]), .B(b[40]), .Z(n5599) );
  XOR U6416 ( .A(n5604), .B(n5339), .Z(n5341) );
  XOR U6417 ( .A(n5605), .B(n5606), .Z(n5339) );
  ANDN U6418 ( .B(n5607), .A(n5608), .Z(n5605) );
  AND U6419 ( .A(a[7]), .B(b[38]), .Z(n5604) );
  XNOR U6420 ( .A(n5609), .B(n5344), .Z(n5346) );
  XOR U6421 ( .A(n5610), .B(n5611), .Z(n5344) );
  ANDN U6422 ( .B(n5612), .A(n5613), .Z(n5610) );
  AND U6423 ( .A(a[8]), .B(b[37]), .Z(n5609) );
  XNOR U6424 ( .A(n5614), .B(n5349), .Z(n5351) );
  XOR U6425 ( .A(n5615), .B(n5616), .Z(n5349) );
  ANDN U6426 ( .B(n5617), .A(n5618), .Z(n5615) );
  AND U6427 ( .A(a[9]), .B(b[36]), .Z(n5614) );
  XNOR U6428 ( .A(n5619), .B(n5354), .Z(n5356) );
  XOR U6429 ( .A(n5620), .B(n5621), .Z(n5354) );
  ANDN U6430 ( .B(n5622), .A(n5623), .Z(n5620) );
  AND U6431 ( .A(b[35]), .B(a[10]), .Z(n5619) );
  XOR U6432 ( .A(n5624), .B(n5625), .Z(n5358) );
  AND U6433 ( .A(n5626), .B(n5627), .Z(n5624) );
  XNOR U6434 ( .A(n5628), .B(n5363), .Z(n5365) );
  XOR U6435 ( .A(n5629), .B(n5630), .Z(n5363) );
  ANDN U6436 ( .B(n5631), .A(n5632), .Z(n5629) );
  AND U6437 ( .A(b[34]), .B(a[11]), .Z(n5628) );
  XOR U6438 ( .A(n5633), .B(n5368), .Z(n5370) );
  XOR U6439 ( .A(n5634), .B(n5635), .Z(n5368) );
  ANDN U6440 ( .B(n5636), .A(n5637), .Z(n5634) );
  AND U6441 ( .A(b[32]), .B(a[13]), .Z(n5633) );
  XNOR U6442 ( .A(n5638), .B(n5373), .Z(n5375) );
  XOR U6443 ( .A(n5639), .B(n5640), .Z(n5373) );
  ANDN U6444 ( .B(n5641), .A(n5642), .Z(n5639) );
  AND U6445 ( .A(b[31]), .B(a[14]), .Z(n5638) );
  XNOR U6446 ( .A(n5643), .B(n5378), .Z(n5380) );
  XOR U6447 ( .A(n5644), .B(n5645), .Z(n5378) );
  ANDN U6448 ( .B(n5646), .A(n5647), .Z(n5644) );
  AND U6449 ( .A(b[30]), .B(a[15]), .Z(n5643) );
  XNOR U6450 ( .A(n5648), .B(n5383), .Z(n5385) );
  XOR U6451 ( .A(n5649), .B(n5650), .Z(n5383) );
  ANDN U6452 ( .B(n5651), .A(n5652), .Z(n5649) );
  AND U6453 ( .A(b[29]), .B(a[16]), .Z(n5648) );
  XOR U6454 ( .A(n5653), .B(n5654), .Z(n5387) );
  AND U6455 ( .A(n5655), .B(n5656), .Z(n5653) );
  XNOR U6456 ( .A(n5657), .B(n5392), .Z(n5394) );
  XOR U6457 ( .A(n5658), .B(n5659), .Z(n5392) );
  ANDN U6458 ( .B(n5660), .A(n5661), .Z(n5658) );
  AND U6459 ( .A(b[28]), .B(a[17]), .Z(n5657) );
  XOR U6460 ( .A(n5662), .B(n5397), .Z(n5399) );
  XOR U6461 ( .A(n5663), .B(n5664), .Z(n5397) );
  ANDN U6462 ( .B(n5665), .A(n5666), .Z(n5663) );
  AND U6463 ( .A(b[26]), .B(a[19]), .Z(n5662) );
  XNOR U6464 ( .A(n5667), .B(n5402), .Z(n5404) );
  XOR U6465 ( .A(n5668), .B(n5669), .Z(n5402) );
  ANDN U6466 ( .B(n5670), .A(n5671), .Z(n5668) );
  AND U6467 ( .A(b[25]), .B(a[20]), .Z(n5667) );
  XNOR U6468 ( .A(n5672), .B(n5407), .Z(n5409) );
  XOR U6469 ( .A(n5673), .B(n5674), .Z(n5407) );
  ANDN U6470 ( .B(n5675), .A(n5676), .Z(n5673) );
  AND U6471 ( .A(b[24]), .B(a[21]), .Z(n5672) );
  XNOR U6472 ( .A(n5677), .B(n5412), .Z(n5414) );
  XOR U6473 ( .A(n5678), .B(n5679), .Z(n5412) );
  ANDN U6474 ( .B(n5680), .A(n5681), .Z(n5678) );
  AND U6475 ( .A(b[23]), .B(a[22]), .Z(n5677) );
  XOR U6476 ( .A(n5682), .B(n5683), .Z(n5416) );
  AND U6477 ( .A(n5684), .B(n5685), .Z(n5682) );
  XNOR U6478 ( .A(n5686), .B(n5421), .Z(n5423) );
  XOR U6479 ( .A(n5687), .B(n5688), .Z(n5421) );
  ANDN U6480 ( .B(n5689), .A(n5690), .Z(n5687) );
  AND U6481 ( .A(b[22]), .B(a[23]), .Z(n5686) );
  XOR U6482 ( .A(n5691), .B(n5426), .Z(n5428) );
  XOR U6483 ( .A(n5692), .B(n5693), .Z(n5426) );
  ANDN U6484 ( .B(n5694), .A(n5695), .Z(n5692) );
  AND U6485 ( .A(b[20]), .B(a[25]), .Z(n5691) );
  XNOR U6486 ( .A(n5696), .B(n5431), .Z(n5433) );
  XOR U6487 ( .A(n5697), .B(n5698), .Z(n5431) );
  ANDN U6488 ( .B(n5699), .A(n5700), .Z(n5697) );
  AND U6489 ( .A(b[19]), .B(a[26]), .Z(n5696) );
  XNOR U6490 ( .A(n5701), .B(n5436), .Z(n5438) );
  XOR U6491 ( .A(n5702), .B(n5703), .Z(n5436) );
  ANDN U6492 ( .B(n5704), .A(n5705), .Z(n5702) );
  AND U6493 ( .A(b[18]), .B(a[27]), .Z(n5701) );
  XNOR U6494 ( .A(n5706), .B(n5441), .Z(n5443) );
  XOR U6495 ( .A(n5707), .B(n5708), .Z(n5441) );
  ANDN U6496 ( .B(n5709), .A(n5710), .Z(n5707) );
  AND U6497 ( .A(b[17]), .B(a[28]), .Z(n5706) );
  XOR U6498 ( .A(n5711), .B(n5712), .Z(n5445) );
  AND U6499 ( .A(n5713), .B(n5714), .Z(n5711) );
  XNOR U6500 ( .A(n5715), .B(n5450), .Z(n5452) );
  XOR U6501 ( .A(n5716), .B(n5717), .Z(n5450) );
  ANDN U6502 ( .B(n5718), .A(n5719), .Z(n5716) );
  AND U6503 ( .A(b[16]), .B(a[29]), .Z(n5715) );
  XOR U6504 ( .A(n5720), .B(n5455), .Z(n5457) );
  XOR U6505 ( .A(n5721), .B(n5722), .Z(n5455) );
  ANDN U6506 ( .B(n5723), .A(n5724), .Z(n5721) );
  AND U6507 ( .A(b[14]), .B(a[31]), .Z(n5720) );
  XNOR U6508 ( .A(n5725), .B(n5460), .Z(n5462) );
  XOR U6509 ( .A(n5726), .B(n5727), .Z(n5460) );
  ANDN U6510 ( .B(n5728), .A(n5729), .Z(n5726) );
  AND U6511 ( .A(b[13]), .B(a[32]), .Z(n5725) );
  XNOR U6512 ( .A(n5730), .B(n5465), .Z(n5467) );
  XOR U6513 ( .A(n5731), .B(n5732), .Z(n5465) );
  ANDN U6514 ( .B(n5733), .A(n5734), .Z(n5731) );
  AND U6515 ( .A(b[12]), .B(a[33]), .Z(n5730) );
  XNOR U6516 ( .A(n5735), .B(n5470), .Z(n5472) );
  XOR U6517 ( .A(n5736), .B(n5737), .Z(n5470) );
  ANDN U6518 ( .B(n5738), .A(n5739), .Z(n5736) );
  AND U6519 ( .A(b[11]), .B(a[34]), .Z(n5735) );
  XOR U6520 ( .A(n5740), .B(n5741), .Z(n5474) );
  AND U6521 ( .A(n5742), .B(n5743), .Z(n5740) );
  XNOR U6522 ( .A(n5744), .B(n5479), .Z(n5481) );
  XOR U6523 ( .A(n5745), .B(n5746), .Z(n5479) );
  ANDN U6524 ( .B(n5747), .A(n5748), .Z(n5745) );
  AND U6525 ( .A(b[10]), .B(a[35]), .Z(n5744) );
  XOR U6526 ( .A(n5749), .B(n5484), .Z(n5486) );
  XOR U6527 ( .A(n5750), .B(n5751), .Z(n5484) );
  ANDN U6528 ( .B(n5752), .A(n5753), .Z(n5750) );
  AND U6529 ( .A(b[8]), .B(a[37]), .Z(n5749) );
  XNOR U6530 ( .A(n5754), .B(n5489), .Z(n5491) );
  XOR U6531 ( .A(n5755), .B(n5756), .Z(n5489) );
  ANDN U6532 ( .B(n5757), .A(n5758), .Z(n5755) );
  AND U6533 ( .A(b[7]), .B(a[38]), .Z(n5754) );
  XNOR U6534 ( .A(n5759), .B(n5494), .Z(n5496) );
  XOR U6535 ( .A(n5760), .B(n5761), .Z(n5494) );
  ANDN U6536 ( .B(n5762), .A(n5763), .Z(n5760) );
  AND U6537 ( .A(b[6]), .B(a[39]), .Z(n5759) );
  XNOR U6538 ( .A(n5764), .B(n5499), .Z(n5501) );
  XOR U6539 ( .A(n5765), .B(n5766), .Z(n5499) );
  ANDN U6540 ( .B(n5767), .A(n5768), .Z(n5765) );
  AND U6541 ( .A(b[5]), .B(a[40]), .Z(n5764) );
  XNOR U6542 ( .A(n5769), .B(n5504), .Z(n5506) );
  XOR U6543 ( .A(n5770), .B(n5771), .Z(n5504) );
  ANDN U6544 ( .B(n5772), .A(n5773), .Z(n5770) );
  AND U6545 ( .A(b[4]), .B(a[41]), .Z(n5769) );
  XNOR U6546 ( .A(n5774), .B(n5775), .Z(n5518) );
  NANDN U6547 ( .A(n5776), .B(n5777), .Z(n5775) );
  XNOR U6548 ( .A(n5778), .B(n5509), .Z(n5511) );
  XNOR U6549 ( .A(n5779), .B(n5780), .Z(n5509) );
  AND U6550 ( .A(n5781), .B(n5782), .Z(n5779) );
  AND U6551 ( .A(b[3]), .B(a[42]), .Z(n5778) );
  NAND U6552 ( .A(a[45]), .B(b[0]), .Z(n5256) );
  XNOR U6553 ( .A(n5524), .B(n5525), .Z(c[44]) );
  XNOR U6554 ( .A(n5776), .B(n5777), .Z(n5525) );
  XOR U6555 ( .A(n5774), .B(n5783), .Z(n5777) );
  NAND U6556 ( .A(b[1]), .B(a[43]), .Z(n5783) );
  XOR U6557 ( .A(n5781), .B(n5784), .Z(n5776) );
  XOR U6558 ( .A(n5774), .B(n5782), .Z(n5784) );
  XNOR U6559 ( .A(n5785), .B(n5780), .Z(n5782) );
  AND U6560 ( .A(b[2]), .B(a[42]), .Z(n5785) );
  NANDN U6561 ( .A(n5786), .B(n5787), .Z(n5774) );
  XOR U6562 ( .A(n5780), .B(n5772), .Z(n5788) );
  XNOR U6563 ( .A(n5771), .B(n5767), .Z(n5789) );
  XNOR U6564 ( .A(n5766), .B(n5762), .Z(n5790) );
  XNOR U6565 ( .A(n5761), .B(n5757), .Z(n5791) );
  XNOR U6566 ( .A(n5756), .B(n5752), .Z(n5792) );
  XNOR U6567 ( .A(n5743), .B(n5742), .Z(n5793) );
  XOR U6568 ( .A(n5794), .B(n5741), .Z(n5742) );
  AND U6569 ( .A(b[8]), .B(a[36]), .Z(n5794) );
  XNOR U6570 ( .A(n5741), .B(n5747), .Z(n5795) );
  XNOR U6571 ( .A(n5746), .B(n5738), .Z(n5796) );
  XNOR U6572 ( .A(n5737), .B(n5733), .Z(n5797) );
  XNOR U6573 ( .A(n5732), .B(n5728), .Z(n5798) );
  XNOR U6574 ( .A(n5727), .B(n5723), .Z(n5799) );
  XNOR U6575 ( .A(n5714), .B(n5713), .Z(n5800) );
  XOR U6576 ( .A(n5801), .B(n5712), .Z(n5713) );
  AND U6577 ( .A(b[14]), .B(a[30]), .Z(n5801) );
  XNOR U6578 ( .A(n5712), .B(n5718), .Z(n5802) );
  XNOR U6579 ( .A(n5717), .B(n5709), .Z(n5803) );
  XNOR U6580 ( .A(n5708), .B(n5704), .Z(n5804) );
  XNOR U6581 ( .A(n5703), .B(n5699), .Z(n5805) );
  XNOR U6582 ( .A(n5698), .B(n5694), .Z(n5806) );
  XNOR U6583 ( .A(n5685), .B(n5684), .Z(n5807) );
  XOR U6584 ( .A(n5808), .B(n5683), .Z(n5684) );
  AND U6585 ( .A(b[20]), .B(a[24]), .Z(n5808) );
  XNOR U6586 ( .A(n5683), .B(n5689), .Z(n5809) );
  XNOR U6587 ( .A(n5688), .B(n5680), .Z(n5810) );
  XNOR U6588 ( .A(n5679), .B(n5675), .Z(n5811) );
  XNOR U6589 ( .A(n5674), .B(n5670), .Z(n5812) );
  XNOR U6590 ( .A(n5669), .B(n5665), .Z(n5813) );
  XNOR U6591 ( .A(n5656), .B(n5655), .Z(n5814) );
  XOR U6592 ( .A(n5815), .B(n5654), .Z(n5655) );
  AND U6593 ( .A(b[26]), .B(a[18]), .Z(n5815) );
  XNOR U6594 ( .A(n5654), .B(n5660), .Z(n5816) );
  XNOR U6595 ( .A(n5659), .B(n5651), .Z(n5817) );
  XNOR U6596 ( .A(n5650), .B(n5646), .Z(n5818) );
  XNOR U6597 ( .A(n5645), .B(n5641), .Z(n5819) );
  XNOR U6598 ( .A(n5640), .B(n5636), .Z(n5820) );
  XNOR U6599 ( .A(n5821), .B(n5822), .Z(n5636) );
  XNOR U6600 ( .A(n5627), .B(n5626), .Z(n5822) );
  XOR U6601 ( .A(n5823), .B(n5625), .Z(n5626) );
  AND U6602 ( .A(b[32]), .B(a[12]), .Z(n5823) );
  XNOR U6603 ( .A(n5625), .B(n5631), .Z(n5824) );
  XNOR U6604 ( .A(n5630), .B(n5622), .Z(n5825) );
  XNOR U6605 ( .A(n5621), .B(n5617), .Z(n5826) );
  XNOR U6606 ( .A(n5616), .B(n5612), .Z(n5827) );
  XNOR U6607 ( .A(n5611), .B(n5607), .Z(n5828) );
  XNOR U6608 ( .A(n5598), .B(n5597), .Z(n5829) );
  XOR U6609 ( .A(n5830), .B(n5596), .Z(n5597) );
  AND U6610 ( .A(a[6]), .B(b[38]), .Z(n5830) );
  XNOR U6611 ( .A(n5596), .B(n5602), .Z(n5831) );
  XNOR U6612 ( .A(n5601), .B(n5593), .Z(n5832) );
  XNOR U6613 ( .A(n5592), .B(n5588), .Z(n5833) );
  XNOR U6614 ( .A(n5587), .B(n5583), .Z(n5834) );
  XNOR U6615 ( .A(n5582), .B(n5578), .Z(n5835) );
  XOR U6616 ( .A(n5836), .B(n5577), .Z(n5578) );
  AND U6617 ( .A(a[0]), .B(b[44]), .Z(n5836) );
  XNOR U6618 ( .A(n5837), .B(n5577), .Z(n5579) );
  XNOR U6619 ( .A(n5838), .B(n5839), .Z(n5577) );
  ANDN U6620 ( .B(n5840), .A(n5841), .Z(n5838) );
  AND U6621 ( .A(a[1]), .B(b[43]), .Z(n5837) );
  XNOR U6622 ( .A(n5842), .B(n5582), .Z(n5584) );
  XOR U6623 ( .A(n5843), .B(n5844), .Z(n5582) );
  ANDN U6624 ( .B(n5845), .A(n5846), .Z(n5843) );
  AND U6625 ( .A(a[2]), .B(b[42]), .Z(n5842) );
  XNOR U6626 ( .A(n5847), .B(n5587), .Z(n5589) );
  XOR U6627 ( .A(n5848), .B(n5849), .Z(n5587) );
  ANDN U6628 ( .B(n5850), .A(n5851), .Z(n5848) );
  AND U6629 ( .A(a[3]), .B(b[41]), .Z(n5847) );
  XNOR U6630 ( .A(n5852), .B(n5592), .Z(n5594) );
  XOR U6631 ( .A(n5853), .B(n5854), .Z(n5592) );
  ANDN U6632 ( .B(n5855), .A(n5856), .Z(n5853) );
  AND U6633 ( .A(a[4]), .B(b[40]), .Z(n5852) );
  XOR U6634 ( .A(n5857), .B(n5858), .Z(n5596) );
  AND U6635 ( .A(n5859), .B(n5860), .Z(n5857) );
  XNOR U6636 ( .A(n5861), .B(n5601), .Z(n5603) );
  XOR U6637 ( .A(n5862), .B(n5863), .Z(n5601) );
  ANDN U6638 ( .B(n5864), .A(n5865), .Z(n5862) );
  AND U6639 ( .A(a[5]), .B(b[39]), .Z(n5861) );
  XOR U6640 ( .A(n5866), .B(n5606), .Z(n5608) );
  XOR U6641 ( .A(n5867), .B(n5868), .Z(n5606) );
  ANDN U6642 ( .B(n5869), .A(n5870), .Z(n5867) );
  AND U6643 ( .A(a[7]), .B(b[37]), .Z(n5866) );
  XNOR U6644 ( .A(n5871), .B(n5611), .Z(n5613) );
  XOR U6645 ( .A(n5872), .B(n5873), .Z(n5611) );
  ANDN U6646 ( .B(n5874), .A(n5875), .Z(n5872) );
  AND U6647 ( .A(a[8]), .B(b[36]), .Z(n5871) );
  XNOR U6648 ( .A(n5876), .B(n5616), .Z(n5618) );
  XOR U6649 ( .A(n5877), .B(n5878), .Z(n5616) );
  ANDN U6650 ( .B(n5879), .A(n5880), .Z(n5877) );
  AND U6651 ( .A(a[9]), .B(b[35]), .Z(n5876) );
  XNOR U6652 ( .A(n5881), .B(n5621), .Z(n5623) );
  XOR U6653 ( .A(n5882), .B(n5883), .Z(n5621) );
  ANDN U6654 ( .B(n5884), .A(n5885), .Z(n5882) );
  AND U6655 ( .A(b[34]), .B(a[10]), .Z(n5881) );
  XOR U6656 ( .A(n5886), .B(n5887), .Z(n5625) );
  AND U6657 ( .A(n5888), .B(n5889), .Z(n5886) );
  XNOR U6658 ( .A(n5890), .B(n5630), .Z(n5632) );
  XOR U6659 ( .A(n5891), .B(n5892), .Z(n5630) );
  ANDN U6660 ( .B(n5893), .A(n5894), .Z(n5891) );
  AND U6661 ( .A(a[11]), .B(b[33]), .Z(n5890) );
  IV U6662 ( .A(n5635), .Z(n5821) );
  XOR U6663 ( .A(n5895), .B(n5635), .Z(n5637) );
  XOR U6664 ( .A(n5896), .B(n5897), .Z(n5635) );
  ANDN U6665 ( .B(n5898), .A(n5899), .Z(n5896) );
  AND U6666 ( .A(b[31]), .B(a[13]), .Z(n5895) );
  XNOR U6667 ( .A(n5900), .B(n5640), .Z(n5642) );
  XOR U6668 ( .A(n5901), .B(n5902), .Z(n5640) );
  ANDN U6669 ( .B(n5903), .A(n5904), .Z(n5901) );
  AND U6670 ( .A(b[30]), .B(a[14]), .Z(n5900) );
  XNOR U6671 ( .A(n5905), .B(n5645), .Z(n5647) );
  XOR U6672 ( .A(n5906), .B(n5907), .Z(n5645) );
  ANDN U6673 ( .B(n5908), .A(n5909), .Z(n5906) );
  AND U6674 ( .A(b[29]), .B(a[15]), .Z(n5905) );
  XNOR U6675 ( .A(n5910), .B(n5650), .Z(n5652) );
  XOR U6676 ( .A(n5911), .B(n5912), .Z(n5650) );
  ANDN U6677 ( .B(n5913), .A(n5914), .Z(n5911) );
  AND U6678 ( .A(b[28]), .B(a[16]), .Z(n5910) );
  XOR U6679 ( .A(n5915), .B(n5916), .Z(n5654) );
  AND U6680 ( .A(n5917), .B(n5918), .Z(n5915) );
  XNOR U6681 ( .A(n5919), .B(n5659), .Z(n5661) );
  XOR U6682 ( .A(n5920), .B(n5921), .Z(n5659) );
  ANDN U6683 ( .B(n5922), .A(n5923), .Z(n5920) );
  AND U6684 ( .A(a[17]), .B(b[27]), .Z(n5919) );
  XOR U6685 ( .A(n5924), .B(n5664), .Z(n5666) );
  XOR U6686 ( .A(n5925), .B(n5926), .Z(n5664) );
  ANDN U6687 ( .B(n5927), .A(n5928), .Z(n5925) );
  AND U6688 ( .A(b[25]), .B(a[19]), .Z(n5924) );
  XNOR U6689 ( .A(n5929), .B(n5669), .Z(n5671) );
  XOR U6690 ( .A(n5930), .B(n5931), .Z(n5669) );
  ANDN U6691 ( .B(n5932), .A(n5933), .Z(n5930) );
  AND U6692 ( .A(b[24]), .B(a[20]), .Z(n5929) );
  XNOR U6693 ( .A(n5934), .B(n5674), .Z(n5676) );
  XOR U6694 ( .A(n5935), .B(n5936), .Z(n5674) );
  ANDN U6695 ( .B(n5937), .A(n5938), .Z(n5935) );
  AND U6696 ( .A(b[23]), .B(a[21]), .Z(n5934) );
  XNOR U6697 ( .A(n5939), .B(n5679), .Z(n5681) );
  XOR U6698 ( .A(n5940), .B(n5941), .Z(n5679) );
  ANDN U6699 ( .B(n5942), .A(n5943), .Z(n5940) );
  AND U6700 ( .A(b[22]), .B(a[22]), .Z(n5939) );
  XOR U6701 ( .A(n5944), .B(n5945), .Z(n5683) );
  AND U6702 ( .A(n5946), .B(n5947), .Z(n5944) );
  XNOR U6703 ( .A(n5948), .B(n5688), .Z(n5690) );
  XOR U6704 ( .A(n5949), .B(n5950), .Z(n5688) );
  ANDN U6705 ( .B(n5951), .A(n5952), .Z(n5949) );
  AND U6706 ( .A(a[23]), .B(b[21]), .Z(n5948) );
  XOR U6707 ( .A(n5953), .B(n5693), .Z(n5695) );
  XOR U6708 ( .A(n5954), .B(n5955), .Z(n5693) );
  ANDN U6709 ( .B(n5956), .A(n5957), .Z(n5954) );
  AND U6710 ( .A(b[19]), .B(a[25]), .Z(n5953) );
  XNOR U6711 ( .A(n5958), .B(n5698), .Z(n5700) );
  XOR U6712 ( .A(n5959), .B(n5960), .Z(n5698) );
  ANDN U6713 ( .B(n5961), .A(n5962), .Z(n5959) );
  AND U6714 ( .A(b[18]), .B(a[26]), .Z(n5958) );
  XNOR U6715 ( .A(n5963), .B(n5703), .Z(n5705) );
  XOR U6716 ( .A(n5964), .B(n5965), .Z(n5703) );
  ANDN U6717 ( .B(n5966), .A(n5967), .Z(n5964) );
  AND U6718 ( .A(b[17]), .B(a[27]), .Z(n5963) );
  XNOR U6719 ( .A(n5968), .B(n5708), .Z(n5710) );
  XOR U6720 ( .A(n5969), .B(n5970), .Z(n5708) );
  ANDN U6721 ( .B(n5971), .A(n5972), .Z(n5969) );
  AND U6722 ( .A(b[16]), .B(a[28]), .Z(n5968) );
  XOR U6723 ( .A(n5973), .B(n5974), .Z(n5712) );
  AND U6724 ( .A(n5975), .B(n5976), .Z(n5973) );
  XNOR U6725 ( .A(n5977), .B(n5717), .Z(n5719) );
  XOR U6726 ( .A(n5978), .B(n5979), .Z(n5717) );
  ANDN U6727 ( .B(n5980), .A(n5981), .Z(n5978) );
  AND U6728 ( .A(a[29]), .B(b[15]), .Z(n5977) );
  XOR U6729 ( .A(n5982), .B(n5722), .Z(n5724) );
  XOR U6730 ( .A(n5983), .B(n5984), .Z(n5722) );
  ANDN U6731 ( .B(n5985), .A(n5986), .Z(n5983) );
  AND U6732 ( .A(b[13]), .B(a[31]), .Z(n5982) );
  XNOR U6733 ( .A(n5987), .B(n5727), .Z(n5729) );
  XOR U6734 ( .A(n5988), .B(n5989), .Z(n5727) );
  ANDN U6735 ( .B(n5990), .A(n5991), .Z(n5988) );
  AND U6736 ( .A(b[12]), .B(a[32]), .Z(n5987) );
  XNOR U6737 ( .A(n5992), .B(n5732), .Z(n5734) );
  XOR U6738 ( .A(n5993), .B(n5994), .Z(n5732) );
  ANDN U6739 ( .B(n5995), .A(n5996), .Z(n5993) );
  AND U6740 ( .A(b[11]), .B(a[33]), .Z(n5992) );
  XNOR U6741 ( .A(n5997), .B(n5737), .Z(n5739) );
  XOR U6742 ( .A(n5998), .B(n5999), .Z(n5737) );
  ANDN U6743 ( .B(n6000), .A(n6001), .Z(n5998) );
  AND U6744 ( .A(b[10]), .B(a[34]), .Z(n5997) );
  XOR U6745 ( .A(n6002), .B(n6003), .Z(n5741) );
  AND U6746 ( .A(n6004), .B(n6005), .Z(n6002) );
  XNOR U6747 ( .A(n6006), .B(n5746), .Z(n5748) );
  XOR U6748 ( .A(n6007), .B(n6008), .Z(n5746) );
  ANDN U6749 ( .B(n6009), .A(n6010), .Z(n6007) );
  AND U6750 ( .A(b[9]), .B(a[35]), .Z(n6006) );
  XOR U6751 ( .A(n6011), .B(n5751), .Z(n5753) );
  XOR U6752 ( .A(n6012), .B(n6013), .Z(n5751) );
  ANDN U6753 ( .B(n6014), .A(n6015), .Z(n6012) );
  AND U6754 ( .A(b[7]), .B(a[37]), .Z(n6011) );
  XNOR U6755 ( .A(n6016), .B(n5756), .Z(n5758) );
  XOR U6756 ( .A(n6017), .B(n6018), .Z(n5756) );
  ANDN U6757 ( .B(n6019), .A(n6020), .Z(n6017) );
  AND U6758 ( .A(b[6]), .B(a[38]), .Z(n6016) );
  XNOR U6759 ( .A(n6021), .B(n5761), .Z(n5763) );
  XOR U6760 ( .A(n6022), .B(n6023), .Z(n5761) );
  ANDN U6761 ( .B(n6024), .A(n6025), .Z(n6022) );
  AND U6762 ( .A(b[5]), .B(a[39]), .Z(n6021) );
  XNOR U6763 ( .A(n6026), .B(n5766), .Z(n5768) );
  XOR U6764 ( .A(n6027), .B(n6028), .Z(n5766) );
  ANDN U6765 ( .B(n6029), .A(n6030), .Z(n6027) );
  AND U6766 ( .A(b[4]), .B(a[40]), .Z(n6026) );
  XNOR U6767 ( .A(n6031), .B(n6032), .Z(n5780) );
  NANDN U6768 ( .A(n6033), .B(n6034), .Z(n6032) );
  XNOR U6769 ( .A(n6035), .B(n5771), .Z(n5773) );
  XNOR U6770 ( .A(n6036), .B(n6037), .Z(n5771) );
  NOR U6771 ( .A(n6038), .B(n6039), .Z(n6036) );
  AND U6772 ( .A(b[3]), .B(a[41]), .Z(n6035) );
  NAND U6773 ( .A(a[44]), .B(b[0]), .Z(n5524) );
  XNOR U6774 ( .A(n5786), .B(n5787), .Z(c[43]) );
  XOR U6775 ( .A(n6040), .B(n6041), .Z(n6033) );
  NAND U6776 ( .A(b[1]), .B(a[42]), .Z(n6041) );
  XOR U6777 ( .A(n6040), .B(n6039), .Z(n6042) );
  XOR U6778 ( .A(n6043), .B(n6037), .Z(n6039) );
  AND U6779 ( .A(b[2]), .B(a[41]), .Z(n6043) );
  IV U6780 ( .A(n6031), .Z(n6040) );
  NANDN U6781 ( .A(n6044), .B(n6045), .Z(n6031) );
  XOR U6782 ( .A(n6037), .B(n6029), .Z(n6046) );
  XNOR U6783 ( .A(n6028), .B(n6024), .Z(n6047) );
  XNOR U6784 ( .A(n6023), .B(n6019), .Z(n6048) );
  XNOR U6785 ( .A(n6018), .B(n6014), .Z(n6049) );
  XNOR U6786 ( .A(n6005), .B(n6004), .Z(n6050) );
  XOR U6787 ( .A(n6051), .B(n6003), .Z(n6004) );
  AND U6788 ( .A(b[7]), .B(a[36]), .Z(n6051) );
  XNOR U6789 ( .A(n6003), .B(n6009), .Z(n6052) );
  XNOR U6790 ( .A(n6008), .B(n6000), .Z(n6053) );
  XNOR U6791 ( .A(n5999), .B(n5995), .Z(n6054) );
  XNOR U6792 ( .A(n5994), .B(n5990), .Z(n6055) );
  XNOR U6793 ( .A(n5989), .B(n5985), .Z(n6056) );
  XNOR U6794 ( .A(n5976), .B(n5975), .Z(n6057) );
  XOR U6795 ( .A(n6058), .B(n5974), .Z(n5975) );
  AND U6796 ( .A(b[13]), .B(a[30]), .Z(n6058) );
  XNOR U6797 ( .A(n5974), .B(n5980), .Z(n6059) );
  XNOR U6798 ( .A(n5979), .B(n5971), .Z(n6060) );
  XNOR U6799 ( .A(n5970), .B(n5966), .Z(n6061) );
  XNOR U6800 ( .A(n5965), .B(n5961), .Z(n6062) );
  XNOR U6801 ( .A(n5960), .B(n5956), .Z(n6063) );
  XNOR U6802 ( .A(n5947), .B(n5946), .Z(n6064) );
  XOR U6803 ( .A(n6065), .B(n5945), .Z(n5946) );
  AND U6804 ( .A(b[19]), .B(a[24]), .Z(n6065) );
  XNOR U6805 ( .A(n5945), .B(n5951), .Z(n6066) );
  XNOR U6806 ( .A(n5950), .B(n5942), .Z(n6067) );
  XNOR U6807 ( .A(n5941), .B(n5937), .Z(n6068) );
  XNOR U6808 ( .A(n5936), .B(n5932), .Z(n6069) );
  XNOR U6809 ( .A(n5931), .B(n5927), .Z(n6070) );
  XNOR U6810 ( .A(n5918), .B(n5917), .Z(n6071) );
  XOR U6811 ( .A(n6072), .B(n5916), .Z(n5917) );
  AND U6812 ( .A(b[25]), .B(a[18]), .Z(n6072) );
  XNOR U6813 ( .A(n5916), .B(n5922), .Z(n6073) );
  XNOR U6814 ( .A(n5921), .B(n5913), .Z(n6074) );
  XNOR U6815 ( .A(n5912), .B(n5908), .Z(n6075) );
  XNOR U6816 ( .A(n5907), .B(n5903), .Z(n6076) );
  XNOR U6817 ( .A(n5902), .B(n5898), .Z(n6077) );
  XNOR U6818 ( .A(n5889), .B(n5888), .Z(n6078) );
  XOR U6819 ( .A(n6079), .B(n5887), .Z(n5888) );
  AND U6820 ( .A(b[31]), .B(a[12]), .Z(n6079) );
  XNOR U6821 ( .A(n5887), .B(n5893), .Z(n6080) );
  XNOR U6822 ( .A(n5892), .B(n5884), .Z(n6081) );
  XNOR U6823 ( .A(n5883), .B(n5879), .Z(n6082) );
  XNOR U6824 ( .A(n5878), .B(n5874), .Z(n6083) );
  XNOR U6825 ( .A(n5873), .B(n5869), .Z(n6084) );
  XNOR U6826 ( .A(n6085), .B(n6086), .Z(n5869) );
  XNOR U6827 ( .A(n5860), .B(n5859), .Z(n6086) );
  XOR U6828 ( .A(n6087), .B(n5858), .Z(n5859) );
  AND U6829 ( .A(a[6]), .B(b[37]), .Z(n6087) );
  XNOR U6830 ( .A(n5858), .B(n5864), .Z(n6088) );
  XNOR U6831 ( .A(n5863), .B(n5855), .Z(n6089) );
  XNOR U6832 ( .A(n5854), .B(n5850), .Z(n6090) );
  XNOR U6833 ( .A(n5849), .B(n5845), .Z(n6091) );
  XNOR U6834 ( .A(n5844), .B(n5840), .Z(n6092) );
  XNOR U6835 ( .A(n6093), .B(n5839), .Z(n5840) );
  AND U6836 ( .A(a[0]), .B(b[43]), .Z(n6093) );
  XOR U6837 ( .A(n6094), .B(n5839), .Z(n5841) );
  XNOR U6838 ( .A(n6095), .B(n6096), .Z(n5839) );
  ANDN U6839 ( .B(n6097), .A(n6098), .Z(n6095) );
  AND U6840 ( .A(a[1]), .B(b[42]), .Z(n6094) );
  XNOR U6841 ( .A(n6099), .B(n5844), .Z(n5846) );
  XOR U6842 ( .A(n6100), .B(n6101), .Z(n5844) );
  ANDN U6843 ( .B(n6102), .A(n6103), .Z(n6100) );
  AND U6844 ( .A(a[2]), .B(b[41]), .Z(n6099) );
  XNOR U6845 ( .A(n6104), .B(n5849), .Z(n5851) );
  XOR U6846 ( .A(n6105), .B(n6106), .Z(n5849) );
  ANDN U6847 ( .B(n6107), .A(n6108), .Z(n6105) );
  AND U6848 ( .A(a[3]), .B(b[40]), .Z(n6104) );
  XNOR U6849 ( .A(n6109), .B(n5854), .Z(n5856) );
  XOR U6850 ( .A(n6110), .B(n6111), .Z(n5854) );
  ANDN U6851 ( .B(n6112), .A(n6113), .Z(n6110) );
  AND U6852 ( .A(a[4]), .B(b[39]), .Z(n6109) );
  XOR U6853 ( .A(n6114), .B(n6115), .Z(n5858) );
  AND U6854 ( .A(n6116), .B(n6117), .Z(n6114) );
  XNOR U6855 ( .A(n6118), .B(n5863), .Z(n5865) );
  XOR U6856 ( .A(n6119), .B(n6120), .Z(n5863) );
  ANDN U6857 ( .B(n6121), .A(n6122), .Z(n6119) );
  AND U6858 ( .A(a[5]), .B(b[38]), .Z(n6118) );
  IV U6859 ( .A(n5868), .Z(n6085) );
  XOR U6860 ( .A(n6123), .B(n5868), .Z(n5870) );
  XOR U6861 ( .A(n6124), .B(n6125), .Z(n5868) );
  ANDN U6862 ( .B(n6126), .A(n6127), .Z(n6124) );
  AND U6863 ( .A(a[7]), .B(b[36]), .Z(n6123) );
  XNOR U6864 ( .A(n6128), .B(n5873), .Z(n5875) );
  XOR U6865 ( .A(n6129), .B(n6130), .Z(n5873) );
  ANDN U6866 ( .B(n6131), .A(n6132), .Z(n6129) );
  AND U6867 ( .A(a[8]), .B(b[35]), .Z(n6128) );
  XNOR U6868 ( .A(n6133), .B(n5878), .Z(n5880) );
  XOR U6869 ( .A(n6134), .B(n6135), .Z(n5878) );
  ANDN U6870 ( .B(n6136), .A(n6137), .Z(n6134) );
  AND U6871 ( .A(a[9]), .B(b[34]), .Z(n6133) );
  XNOR U6872 ( .A(n6138), .B(n5883), .Z(n5885) );
  XOR U6873 ( .A(n6139), .B(n6140), .Z(n5883) );
  ANDN U6874 ( .B(n6141), .A(n6142), .Z(n6139) );
  AND U6875 ( .A(a[10]), .B(b[33]), .Z(n6138) );
  XOR U6876 ( .A(n6143), .B(n6144), .Z(n5887) );
  AND U6877 ( .A(n6145), .B(n6146), .Z(n6143) );
  XNOR U6878 ( .A(n6147), .B(n5892), .Z(n5894) );
  XOR U6879 ( .A(n6148), .B(n6149), .Z(n5892) );
  ANDN U6880 ( .B(n6150), .A(n6151), .Z(n6148) );
  AND U6881 ( .A(b[32]), .B(a[11]), .Z(n6147) );
  XOR U6882 ( .A(n6152), .B(n5897), .Z(n5899) );
  XOR U6883 ( .A(n6153), .B(n6154), .Z(n5897) );
  ANDN U6884 ( .B(n6155), .A(n6156), .Z(n6153) );
  AND U6885 ( .A(b[30]), .B(a[13]), .Z(n6152) );
  XNOR U6886 ( .A(n6157), .B(n5902), .Z(n5904) );
  XOR U6887 ( .A(n6158), .B(n6159), .Z(n5902) );
  ANDN U6888 ( .B(n6160), .A(n6161), .Z(n6158) );
  AND U6889 ( .A(b[29]), .B(a[14]), .Z(n6157) );
  XNOR U6890 ( .A(n6162), .B(n5907), .Z(n5909) );
  XOR U6891 ( .A(n6163), .B(n6164), .Z(n5907) );
  ANDN U6892 ( .B(n6165), .A(n6166), .Z(n6163) );
  AND U6893 ( .A(b[28]), .B(a[15]), .Z(n6162) );
  XNOR U6894 ( .A(n6167), .B(n5912), .Z(n5914) );
  XOR U6895 ( .A(n6168), .B(n6169), .Z(n5912) );
  ANDN U6896 ( .B(n6170), .A(n6171), .Z(n6168) );
  AND U6897 ( .A(a[16]), .B(b[27]), .Z(n6167) );
  XOR U6898 ( .A(n6172), .B(n6173), .Z(n5916) );
  AND U6899 ( .A(n6174), .B(n6175), .Z(n6172) );
  XNOR U6900 ( .A(n6176), .B(n5921), .Z(n5923) );
  XOR U6901 ( .A(n6177), .B(n6178), .Z(n5921) );
  ANDN U6902 ( .B(n6179), .A(n6180), .Z(n6177) );
  AND U6903 ( .A(b[26]), .B(a[17]), .Z(n6176) );
  XOR U6904 ( .A(n6181), .B(n5926), .Z(n5928) );
  XOR U6905 ( .A(n6182), .B(n6183), .Z(n5926) );
  ANDN U6906 ( .B(n6184), .A(n6185), .Z(n6182) );
  AND U6907 ( .A(b[24]), .B(a[19]), .Z(n6181) );
  XNOR U6908 ( .A(n6186), .B(n5931), .Z(n5933) );
  XOR U6909 ( .A(n6187), .B(n6188), .Z(n5931) );
  ANDN U6910 ( .B(n6189), .A(n6190), .Z(n6187) );
  AND U6911 ( .A(b[23]), .B(a[20]), .Z(n6186) );
  XNOR U6912 ( .A(n6191), .B(n5936), .Z(n5938) );
  XOR U6913 ( .A(n6192), .B(n6193), .Z(n5936) );
  ANDN U6914 ( .B(n6194), .A(n6195), .Z(n6192) );
  AND U6915 ( .A(b[22]), .B(a[21]), .Z(n6191) );
  XNOR U6916 ( .A(n6196), .B(n5941), .Z(n5943) );
  XOR U6917 ( .A(n6197), .B(n6198), .Z(n5941) );
  ANDN U6918 ( .B(n6199), .A(n6200), .Z(n6197) );
  AND U6919 ( .A(a[22]), .B(b[21]), .Z(n6196) );
  XOR U6920 ( .A(n6201), .B(n6202), .Z(n5945) );
  AND U6921 ( .A(n6203), .B(n6204), .Z(n6201) );
  XNOR U6922 ( .A(n6205), .B(n5950), .Z(n5952) );
  XOR U6923 ( .A(n6206), .B(n6207), .Z(n5950) );
  ANDN U6924 ( .B(n6208), .A(n6209), .Z(n6206) );
  AND U6925 ( .A(b[20]), .B(a[23]), .Z(n6205) );
  XOR U6926 ( .A(n6210), .B(n5955), .Z(n5957) );
  XOR U6927 ( .A(n6211), .B(n6212), .Z(n5955) );
  ANDN U6928 ( .B(n6213), .A(n6214), .Z(n6211) );
  AND U6929 ( .A(b[18]), .B(a[25]), .Z(n6210) );
  XNOR U6930 ( .A(n6215), .B(n5960), .Z(n5962) );
  XOR U6931 ( .A(n6216), .B(n6217), .Z(n5960) );
  ANDN U6932 ( .B(n6218), .A(n6219), .Z(n6216) );
  AND U6933 ( .A(b[17]), .B(a[26]), .Z(n6215) );
  XNOR U6934 ( .A(n6220), .B(n5965), .Z(n5967) );
  XOR U6935 ( .A(n6221), .B(n6222), .Z(n5965) );
  ANDN U6936 ( .B(n6223), .A(n6224), .Z(n6221) );
  AND U6937 ( .A(b[16]), .B(a[27]), .Z(n6220) );
  XNOR U6938 ( .A(n6225), .B(n5970), .Z(n5972) );
  XOR U6939 ( .A(n6226), .B(n6227), .Z(n5970) );
  ANDN U6940 ( .B(n6228), .A(n6229), .Z(n6226) );
  AND U6941 ( .A(a[28]), .B(b[15]), .Z(n6225) );
  XOR U6942 ( .A(n6230), .B(n6231), .Z(n5974) );
  AND U6943 ( .A(n6232), .B(n6233), .Z(n6230) );
  XNOR U6944 ( .A(n6234), .B(n5979), .Z(n5981) );
  XOR U6945 ( .A(n6235), .B(n6236), .Z(n5979) );
  ANDN U6946 ( .B(n6237), .A(n6238), .Z(n6235) );
  AND U6947 ( .A(b[14]), .B(a[29]), .Z(n6234) );
  XOR U6948 ( .A(n6239), .B(n5984), .Z(n5986) );
  XOR U6949 ( .A(n6240), .B(n6241), .Z(n5984) );
  ANDN U6950 ( .B(n6242), .A(n6243), .Z(n6240) );
  AND U6951 ( .A(b[12]), .B(a[31]), .Z(n6239) );
  XNOR U6952 ( .A(n6244), .B(n5989), .Z(n5991) );
  XOR U6953 ( .A(n6245), .B(n6246), .Z(n5989) );
  ANDN U6954 ( .B(n6247), .A(n6248), .Z(n6245) );
  AND U6955 ( .A(b[11]), .B(a[32]), .Z(n6244) );
  XNOR U6956 ( .A(n6249), .B(n5994), .Z(n5996) );
  XOR U6957 ( .A(n6250), .B(n6251), .Z(n5994) );
  ANDN U6958 ( .B(n6252), .A(n6253), .Z(n6250) );
  AND U6959 ( .A(b[10]), .B(a[33]), .Z(n6249) );
  XNOR U6960 ( .A(n6254), .B(n5999), .Z(n6001) );
  XOR U6961 ( .A(n6255), .B(n6256), .Z(n5999) );
  ANDN U6962 ( .B(n6257), .A(n6258), .Z(n6255) );
  AND U6963 ( .A(b[9]), .B(a[34]), .Z(n6254) );
  XOR U6964 ( .A(n6259), .B(n6260), .Z(n6003) );
  AND U6965 ( .A(n6261), .B(n6262), .Z(n6259) );
  XNOR U6966 ( .A(n6263), .B(n6008), .Z(n6010) );
  XOR U6967 ( .A(n6264), .B(n6265), .Z(n6008) );
  ANDN U6968 ( .B(n6266), .A(n6267), .Z(n6264) );
  AND U6969 ( .A(b[8]), .B(a[35]), .Z(n6263) );
  XOR U6970 ( .A(n6268), .B(n6013), .Z(n6015) );
  XOR U6971 ( .A(n6269), .B(n6270), .Z(n6013) );
  ANDN U6972 ( .B(n6271), .A(n6272), .Z(n6269) );
  AND U6973 ( .A(b[6]), .B(a[37]), .Z(n6268) );
  XNOR U6974 ( .A(n6273), .B(n6018), .Z(n6020) );
  XOR U6975 ( .A(n6274), .B(n6275), .Z(n6018) );
  ANDN U6976 ( .B(n6276), .A(n6277), .Z(n6274) );
  AND U6977 ( .A(b[5]), .B(a[38]), .Z(n6273) );
  XNOR U6978 ( .A(n6278), .B(n6023), .Z(n6025) );
  XOR U6979 ( .A(n6279), .B(n6280), .Z(n6023) );
  ANDN U6980 ( .B(n6281), .A(n6282), .Z(n6279) );
  AND U6981 ( .A(b[4]), .B(a[39]), .Z(n6278) );
  XOR U6982 ( .A(n6283), .B(n6284), .Z(n6037) );
  NANDN U6983 ( .A(n6285), .B(n6286), .Z(n6284) );
  XNOR U6984 ( .A(n6287), .B(n6028), .Z(n6030) );
  XNOR U6985 ( .A(n6288), .B(n6289), .Z(n6028) );
  AND U6986 ( .A(n6290), .B(n6291), .Z(n6288) );
  AND U6987 ( .A(b[3]), .B(a[40]), .Z(n6287) );
  NAND U6988 ( .A(a[43]), .B(b[0]), .Z(n5786) );
  XNOR U6989 ( .A(n6044), .B(n6045), .Z(c[42]) );
  XNOR U6990 ( .A(n6286), .B(n6285), .Z(n6045) );
  XOR U6991 ( .A(n6283), .B(n6292), .Z(n6285) );
  NAND U6992 ( .A(b[1]), .B(a[41]), .Z(n6292) );
  XNOR U6993 ( .A(n6291), .B(n6293), .Z(n6286) );
  XNOR U6994 ( .A(n6283), .B(n6290), .Z(n6293) );
  XNOR U6995 ( .A(n6294), .B(n6289), .Z(n6290) );
  AND U6996 ( .A(b[2]), .B(a[40]), .Z(n6294) );
  ANDN U6997 ( .B(n6295), .A(n6296), .Z(n6283) );
  XOR U6998 ( .A(n6289), .B(n6281), .Z(n6297) );
  XNOR U6999 ( .A(n6280), .B(n6276), .Z(n6298) );
  XNOR U7000 ( .A(n6275), .B(n6271), .Z(n6299) );
  XNOR U7001 ( .A(n6262), .B(n6261), .Z(n6300) );
  XOR U7002 ( .A(n6301), .B(n6260), .Z(n6261) );
  AND U7003 ( .A(b[6]), .B(a[36]), .Z(n6301) );
  XNOR U7004 ( .A(n6260), .B(n6266), .Z(n6302) );
  XNOR U7005 ( .A(n6265), .B(n6257), .Z(n6303) );
  XNOR U7006 ( .A(n6256), .B(n6252), .Z(n6304) );
  XNOR U7007 ( .A(n6251), .B(n6247), .Z(n6305) );
  XNOR U7008 ( .A(n6246), .B(n6242), .Z(n6306) );
  XNOR U7009 ( .A(n6233), .B(n6232), .Z(n6307) );
  XOR U7010 ( .A(n6308), .B(n6231), .Z(n6232) );
  AND U7011 ( .A(b[12]), .B(a[30]), .Z(n6308) );
  XNOR U7012 ( .A(n6231), .B(n6237), .Z(n6309) );
  XNOR U7013 ( .A(n6236), .B(n6228), .Z(n6310) );
  XNOR U7014 ( .A(n6227), .B(n6223), .Z(n6311) );
  XNOR U7015 ( .A(n6222), .B(n6218), .Z(n6312) );
  XNOR U7016 ( .A(n6217), .B(n6213), .Z(n6313) );
  XNOR U7017 ( .A(n6204), .B(n6203), .Z(n6314) );
  XOR U7018 ( .A(n6315), .B(n6202), .Z(n6203) );
  AND U7019 ( .A(b[18]), .B(a[24]), .Z(n6315) );
  XNOR U7020 ( .A(n6202), .B(n6208), .Z(n6316) );
  XNOR U7021 ( .A(n6207), .B(n6199), .Z(n6317) );
  XNOR U7022 ( .A(n6198), .B(n6194), .Z(n6318) );
  XNOR U7023 ( .A(n6193), .B(n6189), .Z(n6319) );
  XNOR U7024 ( .A(n6188), .B(n6184), .Z(n6320) );
  XNOR U7025 ( .A(n6175), .B(n6174), .Z(n6321) );
  XOR U7026 ( .A(n6322), .B(n6173), .Z(n6174) );
  AND U7027 ( .A(b[24]), .B(a[18]), .Z(n6322) );
  XNOR U7028 ( .A(n6173), .B(n6179), .Z(n6323) );
  XNOR U7029 ( .A(n6178), .B(n6170), .Z(n6324) );
  XNOR U7030 ( .A(n6169), .B(n6165), .Z(n6325) );
  XNOR U7031 ( .A(n6164), .B(n6160), .Z(n6326) );
  XNOR U7032 ( .A(n6159), .B(n6155), .Z(n6327) );
  XNOR U7033 ( .A(n6146), .B(n6145), .Z(n6328) );
  XOR U7034 ( .A(n6329), .B(n6144), .Z(n6145) );
  AND U7035 ( .A(b[30]), .B(a[12]), .Z(n6329) );
  XNOR U7036 ( .A(n6144), .B(n6150), .Z(n6330) );
  XNOR U7037 ( .A(n6149), .B(n6141), .Z(n6331) );
  XNOR U7038 ( .A(n6140), .B(n6136), .Z(n6332) );
  XNOR U7039 ( .A(n6135), .B(n6131), .Z(n6333) );
  XNOR U7040 ( .A(n6130), .B(n6126), .Z(n6334) );
  XNOR U7041 ( .A(n6117), .B(n6116), .Z(n6335) );
  XOR U7042 ( .A(n6336), .B(n6115), .Z(n6116) );
  AND U7043 ( .A(a[6]), .B(b[36]), .Z(n6336) );
  XNOR U7044 ( .A(n6115), .B(n6121), .Z(n6337) );
  XNOR U7045 ( .A(n6120), .B(n6112), .Z(n6338) );
  XNOR U7046 ( .A(n6111), .B(n6107), .Z(n6339) );
  XNOR U7047 ( .A(n6106), .B(n6102), .Z(n6340) );
  XNOR U7048 ( .A(n6101), .B(n6097), .Z(n6341) );
  XOR U7049 ( .A(n6342), .B(n6096), .Z(n6097) );
  AND U7050 ( .A(a[0]), .B(b[42]), .Z(n6342) );
  XNOR U7051 ( .A(n6343), .B(n6096), .Z(n6098) );
  XNOR U7052 ( .A(n6344), .B(n6345), .Z(n6096) );
  ANDN U7053 ( .B(n6346), .A(n6347), .Z(n6344) );
  AND U7054 ( .A(a[1]), .B(b[41]), .Z(n6343) );
  XNOR U7055 ( .A(n6348), .B(n6101), .Z(n6103) );
  XOR U7056 ( .A(n6349), .B(n6350), .Z(n6101) );
  ANDN U7057 ( .B(n6351), .A(n6352), .Z(n6349) );
  AND U7058 ( .A(a[2]), .B(b[40]), .Z(n6348) );
  XNOR U7059 ( .A(n6353), .B(n6106), .Z(n6108) );
  XOR U7060 ( .A(n6354), .B(n6355), .Z(n6106) );
  ANDN U7061 ( .B(n6356), .A(n6357), .Z(n6354) );
  AND U7062 ( .A(a[3]), .B(b[39]), .Z(n6353) );
  XNOR U7063 ( .A(n6358), .B(n6111), .Z(n6113) );
  XOR U7064 ( .A(n6359), .B(n6360), .Z(n6111) );
  ANDN U7065 ( .B(n6361), .A(n6362), .Z(n6359) );
  AND U7066 ( .A(a[4]), .B(b[38]), .Z(n6358) );
  XOR U7067 ( .A(n6363), .B(n6364), .Z(n6115) );
  AND U7068 ( .A(n6365), .B(n6366), .Z(n6363) );
  XNOR U7069 ( .A(n6367), .B(n6120), .Z(n6122) );
  XOR U7070 ( .A(n6368), .B(n6369), .Z(n6120) );
  ANDN U7071 ( .B(n6370), .A(n6371), .Z(n6368) );
  AND U7072 ( .A(a[5]), .B(b[37]), .Z(n6367) );
  XOR U7073 ( .A(n6372), .B(n6125), .Z(n6127) );
  XOR U7074 ( .A(n6373), .B(n6374), .Z(n6125) );
  ANDN U7075 ( .B(n6375), .A(n6376), .Z(n6373) );
  AND U7076 ( .A(a[7]), .B(b[35]), .Z(n6372) );
  XNOR U7077 ( .A(n6377), .B(n6130), .Z(n6132) );
  XOR U7078 ( .A(n6378), .B(n6379), .Z(n6130) );
  ANDN U7079 ( .B(n6380), .A(n6381), .Z(n6378) );
  AND U7080 ( .A(a[8]), .B(b[34]), .Z(n6377) );
  XNOR U7081 ( .A(n6382), .B(n6135), .Z(n6137) );
  XOR U7082 ( .A(n6383), .B(n6384), .Z(n6135) );
  ANDN U7083 ( .B(n6385), .A(n6386), .Z(n6383) );
  AND U7084 ( .A(a[9]), .B(b[33]), .Z(n6382) );
  XNOR U7085 ( .A(n6387), .B(n6140), .Z(n6142) );
  XOR U7086 ( .A(n6388), .B(n6389), .Z(n6140) );
  ANDN U7087 ( .B(n6390), .A(n6391), .Z(n6388) );
  AND U7088 ( .A(b[32]), .B(a[10]), .Z(n6387) );
  XOR U7089 ( .A(n6392), .B(n6393), .Z(n6144) );
  AND U7090 ( .A(n6394), .B(n6395), .Z(n6392) );
  XNOR U7091 ( .A(n6396), .B(n6149), .Z(n6151) );
  XOR U7092 ( .A(n6397), .B(n6398), .Z(n6149) );
  ANDN U7093 ( .B(n6399), .A(n6400), .Z(n6397) );
  AND U7094 ( .A(b[31]), .B(a[11]), .Z(n6396) );
  XOR U7095 ( .A(n6401), .B(n6154), .Z(n6156) );
  XOR U7096 ( .A(n6402), .B(n6403), .Z(n6154) );
  ANDN U7097 ( .B(n6404), .A(n6405), .Z(n6402) );
  AND U7098 ( .A(b[29]), .B(a[13]), .Z(n6401) );
  XNOR U7099 ( .A(n6406), .B(n6159), .Z(n6161) );
  XOR U7100 ( .A(n6407), .B(n6408), .Z(n6159) );
  ANDN U7101 ( .B(n6409), .A(n6410), .Z(n6407) );
  AND U7102 ( .A(b[28]), .B(a[14]), .Z(n6406) );
  XNOR U7103 ( .A(n6411), .B(n6164), .Z(n6166) );
  XOR U7104 ( .A(n6412), .B(n6413), .Z(n6164) );
  ANDN U7105 ( .B(n6414), .A(n6415), .Z(n6412) );
  AND U7106 ( .A(a[15]), .B(b[27]), .Z(n6411) );
  XNOR U7107 ( .A(n6416), .B(n6169), .Z(n6171) );
  XOR U7108 ( .A(n6417), .B(n6418), .Z(n6169) );
  ANDN U7109 ( .B(n6419), .A(n6420), .Z(n6417) );
  AND U7110 ( .A(b[26]), .B(a[16]), .Z(n6416) );
  XOR U7111 ( .A(n6421), .B(n6422), .Z(n6173) );
  AND U7112 ( .A(n6423), .B(n6424), .Z(n6421) );
  XNOR U7113 ( .A(n6425), .B(n6178), .Z(n6180) );
  XOR U7114 ( .A(n6426), .B(n6427), .Z(n6178) );
  ANDN U7115 ( .B(n6428), .A(n6429), .Z(n6426) );
  AND U7116 ( .A(b[25]), .B(a[17]), .Z(n6425) );
  XOR U7117 ( .A(n6430), .B(n6183), .Z(n6185) );
  XOR U7118 ( .A(n6431), .B(n6432), .Z(n6183) );
  ANDN U7119 ( .B(n6433), .A(n6434), .Z(n6431) );
  AND U7120 ( .A(b[23]), .B(a[19]), .Z(n6430) );
  XNOR U7121 ( .A(n6435), .B(n6188), .Z(n6190) );
  XOR U7122 ( .A(n6436), .B(n6437), .Z(n6188) );
  ANDN U7123 ( .B(n6438), .A(n6439), .Z(n6436) );
  AND U7124 ( .A(b[22]), .B(a[20]), .Z(n6435) );
  XNOR U7125 ( .A(n6440), .B(n6193), .Z(n6195) );
  XOR U7126 ( .A(n6441), .B(n6442), .Z(n6193) );
  ANDN U7127 ( .B(n6443), .A(n6444), .Z(n6441) );
  AND U7128 ( .A(a[21]), .B(b[21]), .Z(n6440) );
  XNOR U7129 ( .A(n6445), .B(n6198), .Z(n6200) );
  XOR U7130 ( .A(n6446), .B(n6447), .Z(n6198) );
  ANDN U7131 ( .B(n6448), .A(n6449), .Z(n6446) );
  AND U7132 ( .A(b[20]), .B(a[22]), .Z(n6445) );
  XOR U7133 ( .A(n6450), .B(n6451), .Z(n6202) );
  AND U7134 ( .A(n6452), .B(n6453), .Z(n6450) );
  XNOR U7135 ( .A(n6454), .B(n6207), .Z(n6209) );
  XOR U7136 ( .A(n6455), .B(n6456), .Z(n6207) );
  ANDN U7137 ( .B(n6457), .A(n6458), .Z(n6455) );
  AND U7138 ( .A(b[19]), .B(a[23]), .Z(n6454) );
  XOR U7139 ( .A(n6459), .B(n6212), .Z(n6214) );
  XOR U7140 ( .A(n6460), .B(n6461), .Z(n6212) );
  ANDN U7141 ( .B(n6462), .A(n6463), .Z(n6460) );
  AND U7142 ( .A(b[17]), .B(a[25]), .Z(n6459) );
  XNOR U7143 ( .A(n6464), .B(n6217), .Z(n6219) );
  XOR U7144 ( .A(n6465), .B(n6466), .Z(n6217) );
  ANDN U7145 ( .B(n6467), .A(n6468), .Z(n6465) );
  AND U7146 ( .A(b[16]), .B(a[26]), .Z(n6464) );
  XNOR U7147 ( .A(n6469), .B(n6222), .Z(n6224) );
  XOR U7148 ( .A(n6470), .B(n6471), .Z(n6222) );
  ANDN U7149 ( .B(n6472), .A(n6473), .Z(n6470) );
  AND U7150 ( .A(a[27]), .B(b[15]), .Z(n6469) );
  XNOR U7151 ( .A(n6474), .B(n6227), .Z(n6229) );
  XOR U7152 ( .A(n6475), .B(n6476), .Z(n6227) );
  ANDN U7153 ( .B(n6477), .A(n6478), .Z(n6475) );
  AND U7154 ( .A(b[14]), .B(a[28]), .Z(n6474) );
  XOR U7155 ( .A(n6479), .B(n6480), .Z(n6231) );
  AND U7156 ( .A(n6481), .B(n6482), .Z(n6479) );
  XNOR U7157 ( .A(n6483), .B(n6236), .Z(n6238) );
  XOR U7158 ( .A(n6484), .B(n6485), .Z(n6236) );
  ANDN U7159 ( .B(n6486), .A(n6487), .Z(n6484) );
  AND U7160 ( .A(b[13]), .B(a[29]), .Z(n6483) );
  XOR U7161 ( .A(n6488), .B(n6241), .Z(n6243) );
  XOR U7162 ( .A(n6489), .B(n6490), .Z(n6241) );
  ANDN U7163 ( .B(n6491), .A(n6492), .Z(n6489) );
  AND U7164 ( .A(b[11]), .B(a[31]), .Z(n6488) );
  XNOR U7165 ( .A(n6493), .B(n6246), .Z(n6248) );
  XOR U7166 ( .A(n6494), .B(n6495), .Z(n6246) );
  ANDN U7167 ( .B(n6496), .A(n6497), .Z(n6494) );
  AND U7168 ( .A(b[10]), .B(a[32]), .Z(n6493) );
  XNOR U7169 ( .A(n6498), .B(n6251), .Z(n6253) );
  XOR U7170 ( .A(n6499), .B(n6500), .Z(n6251) );
  ANDN U7171 ( .B(n6501), .A(n6502), .Z(n6499) );
  AND U7172 ( .A(b[9]), .B(a[33]), .Z(n6498) );
  XNOR U7173 ( .A(n6503), .B(n6256), .Z(n6258) );
  XOR U7174 ( .A(n6504), .B(n6505), .Z(n6256) );
  ANDN U7175 ( .B(n6506), .A(n6507), .Z(n6504) );
  AND U7176 ( .A(b[8]), .B(a[34]), .Z(n6503) );
  XOR U7177 ( .A(n6508), .B(n6509), .Z(n6260) );
  AND U7178 ( .A(n6510), .B(n6511), .Z(n6508) );
  XNOR U7179 ( .A(n6512), .B(n6265), .Z(n6267) );
  XOR U7180 ( .A(n6513), .B(n6514), .Z(n6265) );
  ANDN U7181 ( .B(n6515), .A(n6516), .Z(n6513) );
  AND U7182 ( .A(b[7]), .B(a[35]), .Z(n6512) );
  XOR U7183 ( .A(n6517), .B(n6270), .Z(n6272) );
  XOR U7184 ( .A(n6518), .B(n6519), .Z(n6270) );
  ANDN U7185 ( .B(n6520), .A(n6521), .Z(n6518) );
  AND U7186 ( .A(b[5]), .B(a[37]), .Z(n6517) );
  XNOR U7187 ( .A(n6522), .B(n6275), .Z(n6277) );
  XOR U7188 ( .A(n6523), .B(n6524), .Z(n6275) );
  ANDN U7189 ( .B(n6525), .A(n6526), .Z(n6523) );
  AND U7190 ( .A(b[4]), .B(a[38]), .Z(n6522) );
  XNOR U7191 ( .A(n6527), .B(n6528), .Z(n6289) );
  NANDN U7192 ( .A(n6529), .B(n6530), .Z(n6528) );
  XNOR U7193 ( .A(n6531), .B(n6280), .Z(n6282) );
  XNOR U7194 ( .A(n6532), .B(n6533), .Z(n6280) );
  AND U7195 ( .A(n6534), .B(n6535), .Z(n6532) );
  AND U7196 ( .A(b[3]), .B(a[39]), .Z(n6531) );
  NAND U7197 ( .A(a[42]), .B(b[0]), .Z(n6044) );
  XNOR U7198 ( .A(n6296), .B(n6295), .Z(c[41]) );
  XNOR U7199 ( .A(n6529), .B(n6530), .Z(n6295) );
  XOR U7200 ( .A(n6527), .B(n6536), .Z(n6530) );
  NAND U7201 ( .A(b[1]), .B(a[40]), .Z(n6536) );
  XOR U7202 ( .A(n6535), .B(n6537), .Z(n6529) );
  XOR U7203 ( .A(n6527), .B(n6534), .Z(n6537) );
  XNOR U7204 ( .A(n6538), .B(n6533), .Z(n6534) );
  AND U7205 ( .A(b[2]), .B(a[39]), .Z(n6538) );
  NANDN U7206 ( .A(n6539), .B(n6540), .Z(n6527) );
  XOR U7207 ( .A(n6533), .B(n6525), .Z(n6541) );
  XNOR U7208 ( .A(n6524), .B(n6520), .Z(n6542) );
  XNOR U7209 ( .A(n6511), .B(n6510), .Z(n6543) );
  XOR U7210 ( .A(n6544), .B(n6509), .Z(n6510) );
  AND U7211 ( .A(b[5]), .B(a[36]), .Z(n6544) );
  XNOR U7212 ( .A(n6509), .B(n6515), .Z(n6545) );
  XNOR U7213 ( .A(n6514), .B(n6506), .Z(n6546) );
  XNOR U7214 ( .A(n6505), .B(n6501), .Z(n6547) );
  XNOR U7215 ( .A(n6500), .B(n6496), .Z(n6548) );
  XNOR U7216 ( .A(n6495), .B(n6491), .Z(n6549) );
  XNOR U7217 ( .A(n6482), .B(n6481), .Z(n6550) );
  XOR U7218 ( .A(n6551), .B(n6480), .Z(n6481) );
  AND U7219 ( .A(b[11]), .B(a[30]), .Z(n6551) );
  XNOR U7220 ( .A(n6480), .B(n6486), .Z(n6552) );
  XNOR U7221 ( .A(n6485), .B(n6477), .Z(n6553) );
  XNOR U7222 ( .A(n6476), .B(n6472), .Z(n6554) );
  XNOR U7223 ( .A(n6471), .B(n6467), .Z(n6555) );
  XNOR U7224 ( .A(n6466), .B(n6462), .Z(n6556) );
  XNOR U7225 ( .A(n6453), .B(n6452), .Z(n6557) );
  XOR U7226 ( .A(n6558), .B(n6451), .Z(n6452) );
  AND U7227 ( .A(b[17]), .B(a[24]), .Z(n6558) );
  XNOR U7228 ( .A(n6451), .B(n6457), .Z(n6559) );
  XNOR U7229 ( .A(n6456), .B(n6448), .Z(n6560) );
  XNOR U7230 ( .A(n6447), .B(n6443), .Z(n6561) );
  XNOR U7231 ( .A(n6442), .B(n6438), .Z(n6562) );
  XNOR U7232 ( .A(n6437), .B(n6433), .Z(n6563) );
  XNOR U7233 ( .A(n6424), .B(n6423), .Z(n6564) );
  XOR U7234 ( .A(n6565), .B(n6422), .Z(n6423) );
  AND U7235 ( .A(b[23]), .B(a[18]), .Z(n6565) );
  XNOR U7236 ( .A(n6422), .B(n6428), .Z(n6566) );
  XNOR U7237 ( .A(n6427), .B(n6419), .Z(n6567) );
  XNOR U7238 ( .A(n6418), .B(n6414), .Z(n6568) );
  XNOR U7239 ( .A(n6413), .B(n6409), .Z(n6569) );
  XNOR U7240 ( .A(n6408), .B(n6404), .Z(n6570) );
  XNOR U7241 ( .A(n6395), .B(n6394), .Z(n6571) );
  XOR U7242 ( .A(n6572), .B(n6393), .Z(n6394) );
  AND U7243 ( .A(b[29]), .B(a[12]), .Z(n6572) );
  XNOR U7244 ( .A(n6393), .B(n6399), .Z(n6573) );
  XNOR U7245 ( .A(n6398), .B(n6390), .Z(n6574) );
  XNOR U7246 ( .A(n6389), .B(n6385), .Z(n6575) );
  XNOR U7247 ( .A(n6384), .B(n6380), .Z(n6576) );
  XNOR U7248 ( .A(n6379), .B(n6375), .Z(n6577) );
  XNOR U7249 ( .A(n6366), .B(n6365), .Z(n6578) );
  XOR U7250 ( .A(n6579), .B(n6364), .Z(n6365) );
  AND U7251 ( .A(a[6]), .B(b[35]), .Z(n6579) );
  XNOR U7252 ( .A(n6364), .B(n6370), .Z(n6580) );
  XNOR U7253 ( .A(n6369), .B(n6361), .Z(n6581) );
  XNOR U7254 ( .A(n6360), .B(n6356), .Z(n6582) );
  XNOR U7255 ( .A(n6355), .B(n6351), .Z(n6583) );
  XNOR U7256 ( .A(n6350), .B(n6346), .Z(n6584) );
  XNOR U7257 ( .A(n6585), .B(n6345), .Z(n6346) );
  AND U7258 ( .A(a[0]), .B(b[41]), .Z(n6585) );
  XOR U7259 ( .A(n6586), .B(n6345), .Z(n6347) );
  XNOR U7260 ( .A(n6587), .B(n6588), .Z(n6345) );
  ANDN U7261 ( .B(n6589), .A(n6590), .Z(n6587) );
  AND U7262 ( .A(a[1]), .B(b[40]), .Z(n6586) );
  XNOR U7263 ( .A(n6591), .B(n6350), .Z(n6352) );
  XOR U7264 ( .A(n6592), .B(n6593), .Z(n6350) );
  ANDN U7265 ( .B(n6594), .A(n6595), .Z(n6592) );
  AND U7266 ( .A(a[2]), .B(b[39]), .Z(n6591) );
  XNOR U7267 ( .A(n6596), .B(n6355), .Z(n6357) );
  XOR U7268 ( .A(n6597), .B(n6598), .Z(n6355) );
  ANDN U7269 ( .B(n6599), .A(n6600), .Z(n6597) );
  AND U7270 ( .A(a[3]), .B(b[38]), .Z(n6596) );
  XNOR U7271 ( .A(n6601), .B(n6360), .Z(n6362) );
  XOR U7272 ( .A(n6602), .B(n6603), .Z(n6360) );
  ANDN U7273 ( .B(n6604), .A(n6605), .Z(n6602) );
  AND U7274 ( .A(a[4]), .B(b[37]), .Z(n6601) );
  XOR U7275 ( .A(n6606), .B(n6607), .Z(n6364) );
  AND U7276 ( .A(n6608), .B(n6609), .Z(n6606) );
  XNOR U7277 ( .A(n6610), .B(n6369), .Z(n6371) );
  XOR U7278 ( .A(n6611), .B(n6612), .Z(n6369) );
  ANDN U7279 ( .B(n6613), .A(n6614), .Z(n6611) );
  AND U7280 ( .A(a[5]), .B(b[36]), .Z(n6610) );
  XOR U7281 ( .A(n6615), .B(n6374), .Z(n6376) );
  XOR U7282 ( .A(n6616), .B(n6617), .Z(n6374) );
  ANDN U7283 ( .B(n6618), .A(n6619), .Z(n6616) );
  AND U7284 ( .A(a[7]), .B(b[34]), .Z(n6615) );
  XNOR U7285 ( .A(n6620), .B(n6379), .Z(n6381) );
  XOR U7286 ( .A(n6621), .B(n6622), .Z(n6379) );
  ANDN U7287 ( .B(n6623), .A(n6624), .Z(n6621) );
  AND U7288 ( .A(a[8]), .B(b[33]), .Z(n6620) );
  XNOR U7289 ( .A(n6625), .B(n6384), .Z(n6386) );
  XOR U7290 ( .A(n6626), .B(n6627), .Z(n6384) );
  ANDN U7291 ( .B(n6628), .A(n6629), .Z(n6626) );
  AND U7292 ( .A(a[9]), .B(b[32]), .Z(n6625) );
  XNOR U7293 ( .A(n6630), .B(n6389), .Z(n6391) );
  XOR U7294 ( .A(n6631), .B(n6632), .Z(n6389) );
  ANDN U7295 ( .B(n6633), .A(n6634), .Z(n6631) );
  AND U7296 ( .A(b[31]), .B(a[10]), .Z(n6630) );
  XOR U7297 ( .A(n6635), .B(n6636), .Z(n6393) );
  AND U7298 ( .A(n6637), .B(n6638), .Z(n6635) );
  XNOR U7299 ( .A(n6639), .B(n6398), .Z(n6400) );
  XOR U7300 ( .A(n6640), .B(n6641), .Z(n6398) );
  ANDN U7301 ( .B(n6642), .A(n6643), .Z(n6640) );
  AND U7302 ( .A(b[30]), .B(a[11]), .Z(n6639) );
  XOR U7303 ( .A(n6644), .B(n6403), .Z(n6405) );
  XOR U7304 ( .A(n6645), .B(n6646), .Z(n6403) );
  ANDN U7305 ( .B(n6647), .A(n6648), .Z(n6645) );
  AND U7306 ( .A(b[28]), .B(a[13]), .Z(n6644) );
  XNOR U7307 ( .A(n6649), .B(n6408), .Z(n6410) );
  XOR U7308 ( .A(n6650), .B(n6651), .Z(n6408) );
  ANDN U7309 ( .B(n6652), .A(n6653), .Z(n6650) );
  AND U7310 ( .A(a[14]), .B(b[27]), .Z(n6649) );
  XNOR U7311 ( .A(n6654), .B(n6413), .Z(n6415) );
  XOR U7312 ( .A(n6655), .B(n6656), .Z(n6413) );
  ANDN U7313 ( .B(n6657), .A(n6658), .Z(n6655) );
  AND U7314 ( .A(b[26]), .B(a[15]), .Z(n6654) );
  XNOR U7315 ( .A(n6659), .B(n6418), .Z(n6420) );
  XOR U7316 ( .A(n6660), .B(n6661), .Z(n6418) );
  ANDN U7317 ( .B(n6662), .A(n6663), .Z(n6660) );
  AND U7318 ( .A(b[25]), .B(a[16]), .Z(n6659) );
  XOR U7319 ( .A(n6664), .B(n6665), .Z(n6422) );
  AND U7320 ( .A(n6666), .B(n6667), .Z(n6664) );
  XNOR U7321 ( .A(n6668), .B(n6427), .Z(n6429) );
  XOR U7322 ( .A(n6669), .B(n6670), .Z(n6427) );
  ANDN U7323 ( .B(n6671), .A(n6672), .Z(n6669) );
  AND U7324 ( .A(b[24]), .B(a[17]), .Z(n6668) );
  XOR U7325 ( .A(n6673), .B(n6432), .Z(n6434) );
  XOR U7326 ( .A(n6674), .B(n6675), .Z(n6432) );
  ANDN U7327 ( .B(n6676), .A(n6677), .Z(n6674) );
  AND U7328 ( .A(b[22]), .B(a[19]), .Z(n6673) );
  XNOR U7329 ( .A(n6678), .B(n6437), .Z(n6439) );
  XOR U7330 ( .A(n6679), .B(n6680), .Z(n6437) );
  ANDN U7331 ( .B(n6681), .A(n6682), .Z(n6679) );
  AND U7332 ( .A(a[20]), .B(b[21]), .Z(n6678) );
  XNOR U7333 ( .A(n6683), .B(n6442), .Z(n6444) );
  XOR U7334 ( .A(n6684), .B(n6685), .Z(n6442) );
  ANDN U7335 ( .B(n6686), .A(n6687), .Z(n6684) );
  AND U7336 ( .A(b[20]), .B(a[21]), .Z(n6683) );
  XNOR U7337 ( .A(n6688), .B(n6447), .Z(n6449) );
  XOR U7338 ( .A(n6689), .B(n6690), .Z(n6447) );
  ANDN U7339 ( .B(n6691), .A(n6692), .Z(n6689) );
  AND U7340 ( .A(b[19]), .B(a[22]), .Z(n6688) );
  XOR U7341 ( .A(n6693), .B(n6694), .Z(n6451) );
  AND U7342 ( .A(n6695), .B(n6696), .Z(n6693) );
  XNOR U7343 ( .A(n6697), .B(n6456), .Z(n6458) );
  XOR U7344 ( .A(n6698), .B(n6699), .Z(n6456) );
  ANDN U7345 ( .B(n6700), .A(n6701), .Z(n6698) );
  AND U7346 ( .A(b[18]), .B(a[23]), .Z(n6697) );
  XOR U7347 ( .A(n6702), .B(n6461), .Z(n6463) );
  XOR U7348 ( .A(n6703), .B(n6704), .Z(n6461) );
  ANDN U7349 ( .B(n6705), .A(n6706), .Z(n6703) );
  AND U7350 ( .A(b[16]), .B(a[25]), .Z(n6702) );
  XNOR U7351 ( .A(n6707), .B(n6466), .Z(n6468) );
  XOR U7352 ( .A(n6708), .B(n6709), .Z(n6466) );
  ANDN U7353 ( .B(n6710), .A(n6711), .Z(n6708) );
  AND U7354 ( .A(a[26]), .B(b[15]), .Z(n6707) );
  XNOR U7355 ( .A(n6712), .B(n6471), .Z(n6473) );
  XOR U7356 ( .A(n6713), .B(n6714), .Z(n6471) );
  ANDN U7357 ( .B(n6715), .A(n6716), .Z(n6713) );
  AND U7358 ( .A(b[14]), .B(a[27]), .Z(n6712) );
  XNOR U7359 ( .A(n6717), .B(n6476), .Z(n6478) );
  XOR U7360 ( .A(n6718), .B(n6719), .Z(n6476) );
  ANDN U7361 ( .B(n6720), .A(n6721), .Z(n6718) );
  AND U7362 ( .A(b[13]), .B(a[28]), .Z(n6717) );
  XOR U7363 ( .A(n6722), .B(n6723), .Z(n6480) );
  AND U7364 ( .A(n6724), .B(n6725), .Z(n6722) );
  XNOR U7365 ( .A(n6726), .B(n6485), .Z(n6487) );
  XOR U7366 ( .A(n6727), .B(n6728), .Z(n6485) );
  ANDN U7367 ( .B(n6729), .A(n6730), .Z(n6727) );
  AND U7368 ( .A(b[12]), .B(a[29]), .Z(n6726) );
  XOR U7369 ( .A(n6731), .B(n6490), .Z(n6492) );
  XOR U7370 ( .A(n6732), .B(n6733), .Z(n6490) );
  ANDN U7371 ( .B(n6734), .A(n6735), .Z(n6732) );
  AND U7372 ( .A(b[10]), .B(a[31]), .Z(n6731) );
  XNOR U7373 ( .A(n6736), .B(n6495), .Z(n6497) );
  XOR U7374 ( .A(n6737), .B(n6738), .Z(n6495) );
  ANDN U7375 ( .B(n6739), .A(n6740), .Z(n6737) );
  AND U7376 ( .A(b[9]), .B(a[32]), .Z(n6736) );
  XNOR U7377 ( .A(n6741), .B(n6500), .Z(n6502) );
  XOR U7378 ( .A(n6742), .B(n6743), .Z(n6500) );
  ANDN U7379 ( .B(n6744), .A(n6745), .Z(n6742) );
  AND U7380 ( .A(b[8]), .B(a[33]), .Z(n6741) );
  XNOR U7381 ( .A(n6746), .B(n6505), .Z(n6507) );
  XOR U7382 ( .A(n6747), .B(n6748), .Z(n6505) );
  ANDN U7383 ( .B(n6749), .A(n6750), .Z(n6747) );
  AND U7384 ( .A(b[7]), .B(a[34]), .Z(n6746) );
  XOR U7385 ( .A(n6751), .B(n6752), .Z(n6509) );
  AND U7386 ( .A(n6753), .B(n6754), .Z(n6751) );
  XNOR U7387 ( .A(n6755), .B(n6514), .Z(n6516) );
  XOR U7388 ( .A(n6756), .B(n6757), .Z(n6514) );
  ANDN U7389 ( .B(n6758), .A(n6759), .Z(n6756) );
  AND U7390 ( .A(b[6]), .B(a[35]), .Z(n6755) );
  XOR U7391 ( .A(n6760), .B(n6519), .Z(n6521) );
  XOR U7392 ( .A(n6761), .B(n6762), .Z(n6519) );
  ANDN U7393 ( .B(n6763), .A(n6764), .Z(n6761) );
  AND U7394 ( .A(b[4]), .B(a[37]), .Z(n6760) );
  XNOR U7395 ( .A(n6765), .B(n6766), .Z(n6533) );
  NANDN U7396 ( .A(n6767), .B(n6768), .Z(n6766) );
  XNOR U7397 ( .A(n6769), .B(n6524), .Z(n6526) );
  XNOR U7398 ( .A(n6770), .B(n6771), .Z(n6524) );
  AND U7399 ( .A(n6772), .B(n6773), .Z(n6770) );
  AND U7400 ( .A(b[3]), .B(a[38]), .Z(n6769) );
  NAND U7401 ( .A(a[41]), .B(b[0]), .Z(n6296) );
  XNOR U7402 ( .A(n6539), .B(n6540), .Z(c[40]) );
  XNOR U7403 ( .A(n6767), .B(n6768), .Z(n6540) );
  XOR U7404 ( .A(n6765), .B(n6774), .Z(n6768) );
  NAND U7405 ( .A(b[1]), .B(a[39]), .Z(n6774) );
  XOR U7406 ( .A(n6773), .B(n6775), .Z(n6767) );
  XOR U7407 ( .A(n6765), .B(n6772), .Z(n6775) );
  XNOR U7408 ( .A(n6776), .B(n6771), .Z(n6772) );
  AND U7409 ( .A(b[2]), .B(a[38]), .Z(n6776) );
  NANDN U7410 ( .A(n6777), .B(n6778), .Z(n6765) );
  XOR U7411 ( .A(n6771), .B(n6763), .Z(n6779) );
  XNOR U7412 ( .A(n6754), .B(n6753), .Z(n6780) );
  XOR U7413 ( .A(n6781), .B(n6752), .Z(n6753) );
  AND U7414 ( .A(b[4]), .B(a[36]), .Z(n6781) );
  XNOR U7415 ( .A(n6752), .B(n6758), .Z(n6782) );
  XNOR U7416 ( .A(n6757), .B(n6749), .Z(n6783) );
  XNOR U7417 ( .A(n6748), .B(n6744), .Z(n6784) );
  XNOR U7418 ( .A(n6743), .B(n6739), .Z(n6785) );
  XNOR U7419 ( .A(n6738), .B(n6734), .Z(n6786) );
  XNOR U7420 ( .A(n6725), .B(n6724), .Z(n6787) );
  XOR U7421 ( .A(n6788), .B(n6723), .Z(n6724) );
  AND U7422 ( .A(b[10]), .B(a[30]), .Z(n6788) );
  XNOR U7423 ( .A(n6723), .B(n6729), .Z(n6789) );
  XNOR U7424 ( .A(n6728), .B(n6720), .Z(n6790) );
  XNOR U7425 ( .A(n6719), .B(n6715), .Z(n6791) );
  XNOR U7426 ( .A(n6714), .B(n6710), .Z(n6792) );
  XNOR U7427 ( .A(n6709), .B(n6705), .Z(n6793) );
  XNOR U7428 ( .A(n6696), .B(n6695), .Z(n6794) );
  XOR U7429 ( .A(n6795), .B(n6694), .Z(n6695) );
  AND U7430 ( .A(b[16]), .B(a[24]), .Z(n6795) );
  XNOR U7431 ( .A(n6694), .B(n6700), .Z(n6796) );
  XNOR U7432 ( .A(n6699), .B(n6691), .Z(n6797) );
  XNOR U7433 ( .A(n6690), .B(n6686), .Z(n6798) );
  XNOR U7434 ( .A(n6685), .B(n6681), .Z(n6799) );
  XNOR U7435 ( .A(n6680), .B(n6676), .Z(n6800) );
  XNOR U7436 ( .A(n6667), .B(n6666), .Z(n6801) );
  XOR U7437 ( .A(n6802), .B(n6665), .Z(n6666) );
  AND U7438 ( .A(b[22]), .B(a[18]), .Z(n6802) );
  XNOR U7439 ( .A(n6665), .B(n6671), .Z(n6803) );
  XNOR U7440 ( .A(n6670), .B(n6662), .Z(n6804) );
  XNOR U7441 ( .A(n6661), .B(n6657), .Z(n6805) );
  XNOR U7442 ( .A(n6656), .B(n6652), .Z(n6806) );
  XNOR U7443 ( .A(n6651), .B(n6647), .Z(n6807) );
  XNOR U7444 ( .A(n6638), .B(n6637), .Z(n6808) );
  XOR U7445 ( .A(n6809), .B(n6636), .Z(n6637) );
  AND U7446 ( .A(b[28]), .B(a[12]), .Z(n6809) );
  XNOR U7447 ( .A(n6636), .B(n6642), .Z(n6810) );
  XNOR U7448 ( .A(n6641), .B(n6633), .Z(n6811) );
  XNOR U7449 ( .A(n6632), .B(n6628), .Z(n6812) );
  XNOR U7450 ( .A(n6627), .B(n6623), .Z(n6813) );
  XNOR U7451 ( .A(n6622), .B(n6618), .Z(n6814) );
  XNOR U7452 ( .A(n6609), .B(n6608), .Z(n6815) );
  XOR U7453 ( .A(n6816), .B(n6607), .Z(n6608) );
  AND U7454 ( .A(a[6]), .B(b[34]), .Z(n6816) );
  XNOR U7455 ( .A(n6607), .B(n6613), .Z(n6817) );
  XNOR U7456 ( .A(n6612), .B(n6604), .Z(n6818) );
  XNOR U7457 ( .A(n6603), .B(n6599), .Z(n6819) );
  XNOR U7458 ( .A(n6598), .B(n6594), .Z(n6820) );
  XNOR U7459 ( .A(n6593), .B(n6589), .Z(n6821) );
  XOR U7460 ( .A(n6822), .B(n6588), .Z(n6589) );
  AND U7461 ( .A(a[0]), .B(b[40]), .Z(n6822) );
  XNOR U7462 ( .A(n6823), .B(n6588), .Z(n6590) );
  XNOR U7463 ( .A(n6824), .B(n6825), .Z(n6588) );
  ANDN U7464 ( .B(n6826), .A(n6827), .Z(n6824) );
  AND U7465 ( .A(a[1]), .B(b[39]), .Z(n6823) );
  XNOR U7466 ( .A(n6828), .B(n6593), .Z(n6595) );
  XOR U7467 ( .A(n6829), .B(n6830), .Z(n6593) );
  ANDN U7468 ( .B(n6831), .A(n6832), .Z(n6829) );
  AND U7469 ( .A(a[2]), .B(b[38]), .Z(n6828) );
  XNOR U7470 ( .A(n6833), .B(n6598), .Z(n6600) );
  XOR U7471 ( .A(n6834), .B(n6835), .Z(n6598) );
  ANDN U7472 ( .B(n6836), .A(n6837), .Z(n6834) );
  AND U7473 ( .A(a[3]), .B(b[37]), .Z(n6833) );
  XNOR U7474 ( .A(n6838), .B(n6603), .Z(n6605) );
  XOR U7475 ( .A(n6839), .B(n6840), .Z(n6603) );
  ANDN U7476 ( .B(n6841), .A(n6842), .Z(n6839) );
  AND U7477 ( .A(a[4]), .B(b[36]), .Z(n6838) );
  XOR U7478 ( .A(n6843), .B(n6844), .Z(n6607) );
  AND U7479 ( .A(n6845), .B(n6846), .Z(n6843) );
  XNOR U7480 ( .A(n6847), .B(n6612), .Z(n6614) );
  XOR U7481 ( .A(n6848), .B(n6849), .Z(n6612) );
  ANDN U7482 ( .B(n6850), .A(n6851), .Z(n6848) );
  AND U7483 ( .A(a[5]), .B(b[35]), .Z(n6847) );
  XOR U7484 ( .A(n6852), .B(n6617), .Z(n6619) );
  XOR U7485 ( .A(n6853), .B(n6854), .Z(n6617) );
  ANDN U7486 ( .B(n6855), .A(n6856), .Z(n6853) );
  AND U7487 ( .A(a[7]), .B(b[33]), .Z(n6852) );
  XNOR U7488 ( .A(n6857), .B(n6622), .Z(n6624) );
  XOR U7489 ( .A(n6858), .B(n6859), .Z(n6622) );
  ANDN U7490 ( .B(n6860), .A(n6861), .Z(n6858) );
  AND U7491 ( .A(a[8]), .B(b[32]), .Z(n6857) );
  XNOR U7492 ( .A(n6862), .B(n6627), .Z(n6629) );
  XOR U7493 ( .A(n6863), .B(n6864), .Z(n6627) );
  ANDN U7494 ( .B(n6865), .A(n6866), .Z(n6863) );
  AND U7495 ( .A(a[9]), .B(b[31]), .Z(n6862) );
  XNOR U7496 ( .A(n6867), .B(n6632), .Z(n6634) );
  XOR U7497 ( .A(n6868), .B(n6869), .Z(n6632) );
  ANDN U7498 ( .B(n6870), .A(n6871), .Z(n6868) );
  AND U7499 ( .A(b[30]), .B(a[10]), .Z(n6867) );
  XOR U7500 ( .A(n6872), .B(n6873), .Z(n6636) );
  AND U7501 ( .A(n6874), .B(n6875), .Z(n6872) );
  XNOR U7502 ( .A(n6876), .B(n6641), .Z(n6643) );
  XOR U7503 ( .A(n6877), .B(n6878), .Z(n6641) );
  ANDN U7504 ( .B(n6879), .A(n6880), .Z(n6877) );
  AND U7505 ( .A(b[29]), .B(a[11]), .Z(n6876) );
  XOR U7506 ( .A(n6881), .B(n6646), .Z(n6648) );
  XOR U7507 ( .A(n6882), .B(n6883), .Z(n6646) );
  ANDN U7508 ( .B(n6884), .A(n6885), .Z(n6882) );
  AND U7509 ( .A(a[13]), .B(b[27]), .Z(n6881) );
  XNOR U7510 ( .A(n6886), .B(n6651), .Z(n6653) );
  XOR U7511 ( .A(n6887), .B(n6888), .Z(n6651) );
  ANDN U7512 ( .B(n6889), .A(n6890), .Z(n6887) );
  AND U7513 ( .A(b[26]), .B(a[14]), .Z(n6886) );
  XNOR U7514 ( .A(n6891), .B(n6656), .Z(n6658) );
  XOR U7515 ( .A(n6892), .B(n6893), .Z(n6656) );
  ANDN U7516 ( .B(n6894), .A(n6895), .Z(n6892) );
  AND U7517 ( .A(b[25]), .B(a[15]), .Z(n6891) );
  XNOR U7518 ( .A(n6896), .B(n6661), .Z(n6663) );
  XOR U7519 ( .A(n6897), .B(n6898), .Z(n6661) );
  ANDN U7520 ( .B(n6899), .A(n6900), .Z(n6897) );
  AND U7521 ( .A(b[24]), .B(a[16]), .Z(n6896) );
  XOR U7522 ( .A(n6901), .B(n6902), .Z(n6665) );
  AND U7523 ( .A(n6903), .B(n6904), .Z(n6901) );
  XNOR U7524 ( .A(n6905), .B(n6670), .Z(n6672) );
  XOR U7525 ( .A(n6906), .B(n6907), .Z(n6670) );
  ANDN U7526 ( .B(n6908), .A(n6909), .Z(n6906) );
  AND U7527 ( .A(b[23]), .B(a[17]), .Z(n6905) );
  XOR U7528 ( .A(n6910), .B(n6675), .Z(n6677) );
  XOR U7529 ( .A(n6911), .B(n6912), .Z(n6675) );
  ANDN U7530 ( .B(n6913), .A(n6914), .Z(n6911) );
  AND U7531 ( .A(a[19]), .B(b[21]), .Z(n6910) );
  XNOR U7532 ( .A(n6915), .B(n6680), .Z(n6682) );
  XOR U7533 ( .A(n6916), .B(n6917), .Z(n6680) );
  ANDN U7534 ( .B(n6918), .A(n6919), .Z(n6916) );
  AND U7535 ( .A(b[20]), .B(a[20]), .Z(n6915) );
  XNOR U7536 ( .A(n6920), .B(n6685), .Z(n6687) );
  XOR U7537 ( .A(n6921), .B(n6922), .Z(n6685) );
  ANDN U7538 ( .B(n6923), .A(n6924), .Z(n6921) );
  AND U7539 ( .A(b[19]), .B(a[21]), .Z(n6920) );
  XNOR U7540 ( .A(n6925), .B(n6690), .Z(n6692) );
  XOR U7541 ( .A(n6926), .B(n6927), .Z(n6690) );
  ANDN U7542 ( .B(n6928), .A(n6929), .Z(n6926) );
  AND U7543 ( .A(b[18]), .B(a[22]), .Z(n6925) );
  XOR U7544 ( .A(n6930), .B(n6931), .Z(n6694) );
  AND U7545 ( .A(n6932), .B(n6933), .Z(n6930) );
  XNOR U7546 ( .A(n6934), .B(n6699), .Z(n6701) );
  XOR U7547 ( .A(n6935), .B(n6936), .Z(n6699) );
  ANDN U7548 ( .B(n6937), .A(n6938), .Z(n6935) );
  AND U7549 ( .A(b[17]), .B(a[23]), .Z(n6934) );
  XOR U7550 ( .A(n6939), .B(n6704), .Z(n6706) );
  XOR U7551 ( .A(n6940), .B(n6941), .Z(n6704) );
  ANDN U7552 ( .B(n6942), .A(n6943), .Z(n6940) );
  AND U7553 ( .A(a[25]), .B(b[15]), .Z(n6939) );
  XNOR U7554 ( .A(n6944), .B(n6709), .Z(n6711) );
  XOR U7555 ( .A(n6945), .B(n6946), .Z(n6709) );
  ANDN U7556 ( .B(n6947), .A(n6948), .Z(n6945) );
  AND U7557 ( .A(b[14]), .B(a[26]), .Z(n6944) );
  XNOR U7558 ( .A(n6949), .B(n6714), .Z(n6716) );
  XOR U7559 ( .A(n6950), .B(n6951), .Z(n6714) );
  ANDN U7560 ( .B(n6952), .A(n6953), .Z(n6950) );
  AND U7561 ( .A(b[13]), .B(a[27]), .Z(n6949) );
  XNOR U7562 ( .A(n6954), .B(n6719), .Z(n6721) );
  XOR U7563 ( .A(n6955), .B(n6956), .Z(n6719) );
  ANDN U7564 ( .B(n6957), .A(n6958), .Z(n6955) );
  AND U7565 ( .A(b[12]), .B(a[28]), .Z(n6954) );
  XOR U7566 ( .A(n6959), .B(n6960), .Z(n6723) );
  AND U7567 ( .A(n6961), .B(n6962), .Z(n6959) );
  XNOR U7568 ( .A(n6963), .B(n6728), .Z(n6730) );
  XOR U7569 ( .A(n6964), .B(n6965), .Z(n6728) );
  ANDN U7570 ( .B(n6966), .A(n6967), .Z(n6964) );
  AND U7571 ( .A(b[11]), .B(a[29]), .Z(n6963) );
  XOR U7572 ( .A(n6968), .B(n6733), .Z(n6735) );
  XOR U7573 ( .A(n6969), .B(n6970), .Z(n6733) );
  ANDN U7574 ( .B(n6971), .A(n6972), .Z(n6969) );
  AND U7575 ( .A(b[9]), .B(a[31]), .Z(n6968) );
  XNOR U7576 ( .A(n6973), .B(n6738), .Z(n6740) );
  XOR U7577 ( .A(n6974), .B(n6975), .Z(n6738) );
  ANDN U7578 ( .B(n6976), .A(n6977), .Z(n6974) );
  AND U7579 ( .A(b[8]), .B(a[32]), .Z(n6973) );
  XNOR U7580 ( .A(n6978), .B(n6743), .Z(n6745) );
  XOR U7581 ( .A(n6979), .B(n6980), .Z(n6743) );
  ANDN U7582 ( .B(n6981), .A(n6982), .Z(n6979) );
  AND U7583 ( .A(b[7]), .B(a[33]), .Z(n6978) );
  XNOR U7584 ( .A(n6983), .B(n6748), .Z(n6750) );
  XOR U7585 ( .A(n6984), .B(n6985), .Z(n6748) );
  ANDN U7586 ( .B(n6986), .A(n6987), .Z(n6984) );
  AND U7587 ( .A(b[6]), .B(a[34]), .Z(n6983) );
  XOR U7588 ( .A(n6988), .B(n6989), .Z(n6752) );
  AND U7589 ( .A(n6990), .B(n6991), .Z(n6988) );
  XNOR U7590 ( .A(n6992), .B(n6757), .Z(n6759) );
  XOR U7591 ( .A(n6993), .B(n6994), .Z(n6757) );
  ANDN U7592 ( .B(n6995), .A(n6996), .Z(n6993) );
  AND U7593 ( .A(b[5]), .B(a[35]), .Z(n6992) );
  XNOR U7594 ( .A(n6997), .B(n6998), .Z(n6771) );
  NANDN U7595 ( .A(n6999), .B(n7000), .Z(n6998) );
  XOR U7596 ( .A(n7001), .B(n6762), .Z(n6764) );
  XOR U7597 ( .A(n7002), .B(n7003), .Z(n6762) );
  ANDN U7598 ( .B(n7004), .A(n7005), .Z(n7002) );
  AND U7599 ( .A(b[3]), .B(a[37]), .Z(n7001) );
  NAND U7600 ( .A(a[40]), .B(b[0]), .Z(n6539) );
  XNOR U7601 ( .A(n7006), .B(n7007), .Z(c[3]) );
  XNOR U7602 ( .A(n6777), .B(n6778), .Z(c[39]) );
  XNOR U7603 ( .A(n6999), .B(n7000), .Z(n6778) );
  XOR U7604 ( .A(n6997), .B(n7008), .Z(n7000) );
  NAND U7605 ( .A(b[1]), .B(a[38]), .Z(n7008) );
  XNOR U7606 ( .A(n7005), .B(n7009), .Z(n6999) );
  XOR U7607 ( .A(n6997), .B(n7004), .Z(n7009) );
  XNOR U7608 ( .A(n7010), .B(n7003), .Z(n7004) );
  AND U7609 ( .A(b[2]), .B(a[37]), .Z(n7010) );
  NANDN U7610 ( .A(n7011), .B(n7012), .Z(n6997) );
  XNOR U7611 ( .A(n7003), .B(n7013), .Z(n7005) );
  XNOR U7612 ( .A(n6991), .B(n6990), .Z(n7013) );
  XOR U7613 ( .A(n7014), .B(n6989), .Z(n6990) );
  AND U7614 ( .A(b[3]), .B(a[36]), .Z(n7014) );
  XNOR U7615 ( .A(n6989), .B(n6995), .Z(n7015) );
  XNOR U7616 ( .A(n6994), .B(n6986), .Z(n7016) );
  XNOR U7617 ( .A(n6985), .B(n6981), .Z(n7017) );
  XNOR U7618 ( .A(n6980), .B(n6976), .Z(n7018) );
  XNOR U7619 ( .A(n6975), .B(n6971), .Z(n7019) );
  XNOR U7620 ( .A(n6962), .B(n6961), .Z(n7020) );
  XOR U7621 ( .A(n7021), .B(n6960), .Z(n6961) );
  AND U7622 ( .A(b[9]), .B(a[30]), .Z(n7021) );
  XNOR U7623 ( .A(n6960), .B(n6966), .Z(n7022) );
  XNOR U7624 ( .A(n6965), .B(n6957), .Z(n7023) );
  XNOR U7625 ( .A(n6956), .B(n6952), .Z(n7024) );
  XNOR U7626 ( .A(n6951), .B(n6947), .Z(n7025) );
  XNOR U7627 ( .A(n6946), .B(n6942), .Z(n7026) );
  XNOR U7628 ( .A(n6933), .B(n6932), .Z(n7027) );
  XOR U7629 ( .A(n7028), .B(n6931), .Z(n6932) );
  AND U7630 ( .A(b[15]), .B(a[24]), .Z(n7028) );
  XNOR U7631 ( .A(n6931), .B(n6937), .Z(n7029) );
  XNOR U7632 ( .A(n6936), .B(n6928), .Z(n7030) );
  XNOR U7633 ( .A(n6927), .B(n6923), .Z(n7031) );
  XNOR U7634 ( .A(n6922), .B(n6918), .Z(n7032) );
  XNOR U7635 ( .A(n6917), .B(n6913), .Z(n7033) );
  XNOR U7636 ( .A(n6904), .B(n6903), .Z(n7034) );
  XOR U7637 ( .A(n7035), .B(n6902), .Z(n6903) );
  AND U7638 ( .A(b[21]), .B(a[18]), .Z(n7035) );
  XNOR U7639 ( .A(n6902), .B(n6908), .Z(n7036) );
  XNOR U7640 ( .A(n6907), .B(n6899), .Z(n7037) );
  XNOR U7641 ( .A(n6898), .B(n6894), .Z(n7038) );
  XNOR U7642 ( .A(n6893), .B(n6889), .Z(n7039) );
  XNOR U7643 ( .A(n6888), .B(n6884), .Z(n7040) );
  XNOR U7644 ( .A(n6875), .B(n6874), .Z(n7041) );
  XOR U7645 ( .A(n7042), .B(n6873), .Z(n6874) );
  AND U7646 ( .A(b[27]), .B(a[12]), .Z(n7042) );
  XNOR U7647 ( .A(n6873), .B(n6879), .Z(n7043) );
  XNOR U7648 ( .A(n6878), .B(n6870), .Z(n7044) );
  XNOR U7649 ( .A(n6869), .B(n6865), .Z(n7045) );
  XNOR U7650 ( .A(n6864), .B(n6860), .Z(n7046) );
  XNOR U7651 ( .A(n6859), .B(n6855), .Z(n7047) );
  XNOR U7652 ( .A(n6846), .B(n6845), .Z(n7048) );
  XOR U7653 ( .A(n7049), .B(n6844), .Z(n6845) );
  AND U7654 ( .A(a[6]), .B(b[33]), .Z(n7049) );
  XNOR U7655 ( .A(n6844), .B(n6850), .Z(n7050) );
  XNOR U7656 ( .A(n6849), .B(n6841), .Z(n7051) );
  XNOR U7657 ( .A(n6840), .B(n6836), .Z(n7052) );
  XNOR U7658 ( .A(n6835), .B(n6831), .Z(n7053) );
  XNOR U7659 ( .A(n6830), .B(n6826), .Z(n7054) );
  XNOR U7660 ( .A(n7055), .B(n6825), .Z(n6826) );
  AND U7661 ( .A(a[0]), .B(b[39]), .Z(n7055) );
  XOR U7662 ( .A(n7056), .B(n6825), .Z(n6827) );
  XNOR U7663 ( .A(n7057), .B(n7058), .Z(n6825) );
  ANDN U7664 ( .B(n7059), .A(n7060), .Z(n7057) );
  AND U7665 ( .A(a[1]), .B(b[38]), .Z(n7056) );
  XNOR U7666 ( .A(n7061), .B(n6830), .Z(n6832) );
  XOR U7667 ( .A(n7062), .B(n7063), .Z(n6830) );
  ANDN U7668 ( .B(n7064), .A(n7065), .Z(n7062) );
  AND U7669 ( .A(a[2]), .B(b[37]), .Z(n7061) );
  XNOR U7670 ( .A(n7066), .B(n6835), .Z(n6837) );
  XOR U7671 ( .A(n7067), .B(n7068), .Z(n6835) );
  ANDN U7672 ( .B(n7069), .A(n7070), .Z(n7067) );
  AND U7673 ( .A(a[3]), .B(b[36]), .Z(n7066) );
  XNOR U7674 ( .A(n7071), .B(n6840), .Z(n6842) );
  XOR U7675 ( .A(n7072), .B(n7073), .Z(n6840) );
  ANDN U7676 ( .B(n7074), .A(n7075), .Z(n7072) );
  AND U7677 ( .A(a[4]), .B(b[35]), .Z(n7071) );
  XOR U7678 ( .A(n7076), .B(n7077), .Z(n6844) );
  AND U7679 ( .A(n7078), .B(n7079), .Z(n7076) );
  XNOR U7680 ( .A(n7080), .B(n6849), .Z(n6851) );
  XOR U7681 ( .A(n7081), .B(n7082), .Z(n6849) );
  ANDN U7682 ( .B(n7083), .A(n7084), .Z(n7081) );
  AND U7683 ( .A(a[5]), .B(b[34]), .Z(n7080) );
  XOR U7684 ( .A(n7085), .B(n6854), .Z(n6856) );
  XOR U7685 ( .A(n7086), .B(n7087), .Z(n6854) );
  ANDN U7686 ( .B(n7088), .A(n7089), .Z(n7086) );
  AND U7687 ( .A(a[7]), .B(b[32]), .Z(n7085) );
  XNOR U7688 ( .A(n7090), .B(n6859), .Z(n6861) );
  XOR U7689 ( .A(n7091), .B(n7092), .Z(n6859) );
  ANDN U7690 ( .B(n7093), .A(n7094), .Z(n7091) );
  AND U7691 ( .A(a[8]), .B(b[31]), .Z(n7090) );
  XNOR U7692 ( .A(n7095), .B(n6864), .Z(n6866) );
  XOR U7693 ( .A(n7096), .B(n7097), .Z(n6864) );
  ANDN U7694 ( .B(n7098), .A(n7099), .Z(n7096) );
  AND U7695 ( .A(a[9]), .B(b[30]), .Z(n7095) );
  XNOR U7696 ( .A(n7100), .B(n6869), .Z(n6871) );
  XOR U7697 ( .A(n7101), .B(n7102), .Z(n6869) );
  ANDN U7698 ( .B(n7103), .A(n7104), .Z(n7101) );
  AND U7699 ( .A(b[29]), .B(a[10]), .Z(n7100) );
  XOR U7700 ( .A(n7105), .B(n7106), .Z(n6873) );
  AND U7701 ( .A(n7107), .B(n7108), .Z(n7105) );
  XNOR U7702 ( .A(n7109), .B(n6878), .Z(n6880) );
  XOR U7703 ( .A(n7110), .B(n7111), .Z(n6878) );
  ANDN U7704 ( .B(n7112), .A(n7113), .Z(n7110) );
  AND U7705 ( .A(b[28]), .B(a[11]), .Z(n7109) );
  XOR U7706 ( .A(n7114), .B(n6883), .Z(n6885) );
  XOR U7707 ( .A(n7115), .B(n7116), .Z(n6883) );
  ANDN U7708 ( .B(n7117), .A(n7118), .Z(n7115) );
  AND U7709 ( .A(b[26]), .B(a[13]), .Z(n7114) );
  XNOR U7710 ( .A(n7119), .B(n6888), .Z(n6890) );
  XOR U7711 ( .A(n7120), .B(n7121), .Z(n6888) );
  ANDN U7712 ( .B(n7122), .A(n7123), .Z(n7120) );
  AND U7713 ( .A(b[25]), .B(a[14]), .Z(n7119) );
  XNOR U7714 ( .A(n7124), .B(n6893), .Z(n6895) );
  XOR U7715 ( .A(n7125), .B(n7126), .Z(n6893) );
  ANDN U7716 ( .B(n7127), .A(n7128), .Z(n7125) );
  AND U7717 ( .A(b[24]), .B(a[15]), .Z(n7124) );
  XNOR U7718 ( .A(n7129), .B(n6898), .Z(n6900) );
  XOR U7719 ( .A(n7130), .B(n7131), .Z(n6898) );
  ANDN U7720 ( .B(n7132), .A(n7133), .Z(n7130) );
  AND U7721 ( .A(b[23]), .B(a[16]), .Z(n7129) );
  XOR U7722 ( .A(n7134), .B(n7135), .Z(n6902) );
  AND U7723 ( .A(n7136), .B(n7137), .Z(n7134) );
  XNOR U7724 ( .A(n7138), .B(n6907), .Z(n6909) );
  XOR U7725 ( .A(n7139), .B(n7140), .Z(n6907) );
  ANDN U7726 ( .B(n7141), .A(n7142), .Z(n7139) );
  AND U7727 ( .A(b[22]), .B(a[17]), .Z(n7138) );
  XOR U7728 ( .A(n7143), .B(n6912), .Z(n6914) );
  XOR U7729 ( .A(n7144), .B(n7145), .Z(n6912) );
  ANDN U7730 ( .B(n7146), .A(n7147), .Z(n7144) );
  AND U7731 ( .A(b[20]), .B(a[19]), .Z(n7143) );
  XNOR U7732 ( .A(n7148), .B(n6917), .Z(n6919) );
  XOR U7733 ( .A(n7149), .B(n7150), .Z(n6917) );
  ANDN U7734 ( .B(n7151), .A(n7152), .Z(n7149) );
  AND U7735 ( .A(b[19]), .B(a[20]), .Z(n7148) );
  XNOR U7736 ( .A(n7153), .B(n6922), .Z(n6924) );
  XOR U7737 ( .A(n7154), .B(n7155), .Z(n6922) );
  ANDN U7738 ( .B(n7156), .A(n7157), .Z(n7154) );
  AND U7739 ( .A(b[18]), .B(a[21]), .Z(n7153) );
  XNOR U7740 ( .A(n7158), .B(n6927), .Z(n6929) );
  XOR U7741 ( .A(n7159), .B(n7160), .Z(n6927) );
  ANDN U7742 ( .B(n7161), .A(n7162), .Z(n7159) );
  AND U7743 ( .A(b[17]), .B(a[22]), .Z(n7158) );
  XOR U7744 ( .A(n7163), .B(n7164), .Z(n6931) );
  AND U7745 ( .A(n7165), .B(n7166), .Z(n7163) );
  XNOR U7746 ( .A(n7167), .B(n6936), .Z(n6938) );
  XOR U7747 ( .A(n7168), .B(n7169), .Z(n6936) );
  ANDN U7748 ( .B(n7170), .A(n7171), .Z(n7168) );
  AND U7749 ( .A(b[16]), .B(a[23]), .Z(n7167) );
  XOR U7750 ( .A(n7172), .B(n6941), .Z(n6943) );
  XOR U7751 ( .A(n7173), .B(n7174), .Z(n6941) );
  ANDN U7752 ( .B(n7175), .A(n7176), .Z(n7173) );
  AND U7753 ( .A(b[14]), .B(a[25]), .Z(n7172) );
  XNOR U7754 ( .A(n7177), .B(n6946), .Z(n6948) );
  XOR U7755 ( .A(n7178), .B(n7179), .Z(n6946) );
  ANDN U7756 ( .B(n7180), .A(n7181), .Z(n7178) );
  AND U7757 ( .A(b[13]), .B(a[26]), .Z(n7177) );
  XNOR U7758 ( .A(n7182), .B(n6951), .Z(n6953) );
  XOR U7759 ( .A(n7183), .B(n7184), .Z(n6951) );
  ANDN U7760 ( .B(n7185), .A(n7186), .Z(n7183) );
  AND U7761 ( .A(b[12]), .B(a[27]), .Z(n7182) );
  XNOR U7762 ( .A(n7187), .B(n6956), .Z(n6958) );
  XOR U7763 ( .A(n7188), .B(n7189), .Z(n6956) );
  ANDN U7764 ( .B(n7190), .A(n7191), .Z(n7188) );
  AND U7765 ( .A(b[11]), .B(a[28]), .Z(n7187) );
  XOR U7766 ( .A(n7192), .B(n7193), .Z(n6960) );
  AND U7767 ( .A(n7194), .B(n7195), .Z(n7192) );
  XNOR U7768 ( .A(n7196), .B(n6965), .Z(n6967) );
  XOR U7769 ( .A(n7197), .B(n7198), .Z(n6965) );
  ANDN U7770 ( .B(n7199), .A(n7200), .Z(n7197) );
  AND U7771 ( .A(b[10]), .B(a[29]), .Z(n7196) );
  XOR U7772 ( .A(n7201), .B(n6970), .Z(n6972) );
  XOR U7773 ( .A(n7202), .B(n7203), .Z(n6970) );
  ANDN U7774 ( .B(n7204), .A(n7205), .Z(n7202) );
  AND U7775 ( .A(b[8]), .B(a[31]), .Z(n7201) );
  XNOR U7776 ( .A(n7206), .B(n6975), .Z(n6977) );
  XOR U7777 ( .A(n7207), .B(n7208), .Z(n6975) );
  ANDN U7778 ( .B(n7209), .A(n7210), .Z(n7207) );
  AND U7779 ( .A(b[7]), .B(a[32]), .Z(n7206) );
  XNOR U7780 ( .A(n7211), .B(n6980), .Z(n6982) );
  XOR U7781 ( .A(n7212), .B(n7213), .Z(n6980) );
  ANDN U7782 ( .B(n7214), .A(n7215), .Z(n7212) );
  AND U7783 ( .A(b[6]), .B(a[33]), .Z(n7211) );
  XNOR U7784 ( .A(n7216), .B(n6985), .Z(n6987) );
  XOR U7785 ( .A(n7217), .B(n7218), .Z(n6985) );
  ANDN U7786 ( .B(n7219), .A(n7220), .Z(n7217) );
  AND U7787 ( .A(b[5]), .B(a[34]), .Z(n7216) );
  XOR U7788 ( .A(n7221), .B(n7222), .Z(n6989) );
  ANDN U7789 ( .B(n7223), .A(n7224), .Z(n7221) );
  XNOR U7790 ( .A(n7225), .B(n6994), .Z(n6996) );
  XOR U7791 ( .A(n7226), .B(n7227), .Z(n6994) );
  ANDN U7792 ( .B(n7228), .A(n7229), .Z(n7226) );
  AND U7793 ( .A(b[4]), .B(a[35]), .Z(n7225) );
  XNOR U7794 ( .A(n7230), .B(n7231), .Z(n7003) );
  NAND U7795 ( .A(n7232), .B(n7233), .Z(n7231) );
  NAND U7796 ( .A(a[39]), .B(b[0]), .Z(n6777) );
  XNOR U7797 ( .A(n7011), .B(n7012), .Z(c[38]) );
  XOR U7798 ( .A(n7232), .B(n7233), .Z(n7012) );
  XOR U7799 ( .A(n7230), .B(n7234), .Z(n7233) );
  NAND U7800 ( .A(b[1]), .B(a[37]), .Z(n7234) );
  XOR U7801 ( .A(n7230), .B(n7223), .Z(n7235) );
  XNOR U7802 ( .A(n7222), .B(n7228), .Z(n7236) );
  XNOR U7803 ( .A(n7227), .B(n7219), .Z(n7237) );
  XNOR U7804 ( .A(n7218), .B(n7214), .Z(n7238) );
  XNOR U7805 ( .A(n7213), .B(n7209), .Z(n7239) );
  XNOR U7806 ( .A(n7208), .B(n7204), .Z(n7240) );
  XNOR U7807 ( .A(n7195), .B(n7194), .Z(n7241) );
  XOR U7808 ( .A(n7242), .B(n7193), .Z(n7194) );
  AND U7809 ( .A(b[8]), .B(a[30]), .Z(n7242) );
  XNOR U7810 ( .A(n7193), .B(n7199), .Z(n7243) );
  XNOR U7811 ( .A(n7198), .B(n7190), .Z(n7244) );
  XNOR U7812 ( .A(n7189), .B(n7185), .Z(n7245) );
  XNOR U7813 ( .A(n7184), .B(n7180), .Z(n7246) );
  XNOR U7814 ( .A(n7179), .B(n7175), .Z(n7247) );
  XNOR U7815 ( .A(n7166), .B(n7165), .Z(n7248) );
  XOR U7816 ( .A(n7249), .B(n7164), .Z(n7165) );
  AND U7817 ( .A(b[14]), .B(a[24]), .Z(n7249) );
  XNOR U7818 ( .A(n7164), .B(n7170), .Z(n7250) );
  XNOR U7819 ( .A(n7169), .B(n7161), .Z(n7251) );
  XNOR U7820 ( .A(n7160), .B(n7156), .Z(n7252) );
  XNOR U7821 ( .A(n7155), .B(n7151), .Z(n7253) );
  XNOR U7822 ( .A(n7150), .B(n7146), .Z(n7254) );
  XNOR U7823 ( .A(n7137), .B(n7136), .Z(n7255) );
  XOR U7824 ( .A(n7256), .B(n7135), .Z(n7136) );
  AND U7825 ( .A(b[20]), .B(a[18]), .Z(n7256) );
  XNOR U7826 ( .A(n7135), .B(n7141), .Z(n7257) );
  XNOR U7827 ( .A(n7140), .B(n7132), .Z(n7258) );
  XNOR U7828 ( .A(n7131), .B(n7127), .Z(n7259) );
  XNOR U7829 ( .A(n7126), .B(n7122), .Z(n7260) );
  XNOR U7830 ( .A(n7121), .B(n7117), .Z(n7261) );
  XNOR U7831 ( .A(n7108), .B(n7107), .Z(n7262) );
  XOR U7832 ( .A(n7263), .B(n7106), .Z(n7107) );
  AND U7833 ( .A(b[26]), .B(a[12]), .Z(n7263) );
  XNOR U7834 ( .A(n7106), .B(n7112), .Z(n7264) );
  XNOR U7835 ( .A(n7111), .B(n7103), .Z(n7265) );
  XNOR U7836 ( .A(n7102), .B(n7098), .Z(n7266) );
  XNOR U7837 ( .A(n7097), .B(n7093), .Z(n7267) );
  XNOR U7838 ( .A(n7092), .B(n7088), .Z(n7268) );
  XNOR U7839 ( .A(n7079), .B(n7078), .Z(n7269) );
  XOR U7840 ( .A(n7270), .B(n7077), .Z(n7078) );
  AND U7841 ( .A(a[6]), .B(b[32]), .Z(n7270) );
  XNOR U7842 ( .A(n7077), .B(n7083), .Z(n7271) );
  XNOR U7843 ( .A(n7082), .B(n7074), .Z(n7272) );
  XNOR U7844 ( .A(n7073), .B(n7069), .Z(n7273) );
  XNOR U7845 ( .A(n7068), .B(n7064), .Z(n7274) );
  XNOR U7846 ( .A(n7063), .B(n7059), .Z(n7275) );
  XOR U7847 ( .A(n7276), .B(n7058), .Z(n7059) );
  AND U7848 ( .A(a[0]), .B(b[38]), .Z(n7276) );
  XNOR U7849 ( .A(n7277), .B(n7058), .Z(n7060) );
  XNOR U7850 ( .A(n7278), .B(n7279), .Z(n7058) );
  ANDN U7851 ( .B(n7280), .A(n7281), .Z(n7278) );
  AND U7852 ( .A(a[1]), .B(b[37]), .Z(n7277) );
  XNOR U7853 ( .A(n7282), .B(n7063), .Z(n7065) );
  XOR U7854 ( .A(n7283), .B(n7284), .Z(n7063) );
  ANDN U7855 ( .B(n7285), .A(n7286), .Z(n7283) );
  AND U7856 ( .A(a[2]), .B(b[36]), .Z(n7282) );
  XNOR U7857 ( .A(n7287), .B(n7068), .Z(n7070) );
  XOR U7858 ( .A(n7288), .B(n7289), .Z(n7068) );
  ANDN U7859 ( .B(n7290), .A(n7291), .Z(n7288) );
  AND U7860 ( .A(a[3]), .B(b[35]), .Z(n7287) );
  XNOR U7861 ( .A(n7292), .B(n7073), .Z(n7075) );
  XOR U7862 ( .A(n7293), .B(n7294), .Z(n7073) );
  ANDN U7863 ( .B(n7295), .A(n7296), .Z(n7293) );
  AND U7864 ( .A(a[4]), .B(b[34]), .Z(n7292) );
  XOR U7865 ( .A(n7297), .B(n7298), .Z(n7077) );
  AND U7866 ( .A(n7299), .B(n7300), .Z(n7297) );
  XNOR U7867 ( .A(n7301), .B(n7082), .Z(n7084) );
  XOR U7868 ( .A(n7302), .B(n7303), .Z(n7082) );
  ANDN U7869 ( .B(n7304), .A(n7305), .Z(n7302) );
  AND U7870 ( .A(a[5]), .B(b[33]), .Z(n7301) );
  XOR U7871 ( .A(n7306), .B(n7087), .Z(n7089) );
  XOR U7872 ( .A(n7307), .B(n7308), .Z(n7087) );
  ANDN U7873 ( .B(n7309), .A(n7310), .Z(n7307) );
  AND U7874 ( .A(a[7]), .B(b[31]), .Z(n7306) );
  XNOR U7875 ( .A(n7311), .B(n7092), .Z(n7094) );
  XOR U7876 ( .A(n7312), .B(n7313), .Z(n7092) );
  ANDN U7877 ( .B(n7314), .A(n7315), .Z(n7312) );
  AND U7878 ( .A(a[8]), .B(b[30]), .Z(n7311) );
  XNOR U7879 ( .A(n7316), .B(n7097), .Z(n7099) );
  XOR U7880 ( .A(n7317), .B(n7318), .Z(n7097) );
  ANDN U7881 ( .B(n7319), .A(n7320), .Z(n7317) );
  AND U7882 ( .A(a[9]), .B(b[29]), .Z(n7316) );
  XNOR U7883 ( .A(n7321), .B(n7102), .Z(n7104) );
  XOR U7884 ( .A(n7322), .B(n7323), .Z(n7102) );
  ANDN U7885 ( .B(n7324), .A(n7325), .Z(n7322) );
  AND U7886 ( .A(b[28]), .B(a[10]), .Z(n7321) );
  XOR U7887 ( .A(n7326), .B(n7327), .Z(n7106) );
  AND U7888 ( .A(n7328), .B(n7329), .Z(n7326) );
  XNOR U7889 ( .A(n7330), .B(n7111), .Z(n7113) );
  XOR U7890 ( .A(n7331), .B(n7332), .Z(n7111) );
  ANDN U7891 ( .B(n7333), .A(n7334), .Z(n7331) );
  AND U7892 ( .A(a[11]), .B(b[27]), .Z(n7330) );
  XOR U7893 ( .A(n7335), .B(n7116), .Z(n7118) );
  XOR U7894 ( .A(n7336), .B(n7337), .Z(n7116) );
  ANDN U7895 ( .B(n7338), .A(n7339), .Z(n7336) );
  AND U7896 ( .A(b[25]), .B(a[13]), .Z(n7335) );
  XNOR U7897 ( .A(n7340), .B(n7121), .Z(n7123) );
  XOR U7898 ( .A(n7341), .B(n7342), .Z(n7121) );
  ANDN U7899 ( .B(n7343), .A(n7344), .Z(n7341) );
  AND U7900 ( .A(b[24]), .B(a[14]), .Z(n7340) );
  XNOR U7901 ( .A(n7345), .B(n7126), .Z(n7128) );
  XOR U7902 ( .A(n7346), .B(n7347), .Z(n7126) );
  ANDN U7903 ( .B(n7348), .A(n7349), .Z(n7346) );
  AND U7904 ( .A(b[23]), .B(a[15]), .Z(n7345) );
  XNOR U7905 ( .A(n7350), .B(n7131), .Z(n7133) );
  XOR U7906 ( .A(n7351), .B(n7352), .Z(n7131) );
  ANDN U7907 ( .B(n7353), .A(n7354), .Z(n7351) );
  AND U7908 ( .A(b[22]), .B(a[16]), .Z(n7350) );
  XOR U7909 ( .A(n7355), .B(n7356), .Z(n7135) );
  AND U7910 ( .A(n7357), .B(n7358), .Z(n7355) );
  XNOR U7911 ( .A(n7359), .B(n7140), .Z(n7142) );
  XOR U7912 ( .A(n7360), .B(n7361), .Z(n7140) );
  ANDN U7913 ( .B(n7362), .A(n7363), .Z(n7360) );
  AND U7914 ( .A(a[17]), .B(b[21]), .Z(n7359) );
  XOR U7915 ( .A(n7364), .B(n7145), .Z(n7147) );
  XOR U7916 ( .A(n7365), .B(n7366), .Z(n7145) );
  ANDN U7917 ( .B(n7367), .A(n7368), .Z(n7365) );
  AND U7918 ( .A(b[19]), .B(a[19]), .Z(n7364) );
  XNOR U7919 ( .A(n7369), .B(n7150), .Z(n7152) );
  XOR U7920 ( .A(n7370), .B(n7371), .Z(n7150) );
  ANDN U7921 ( .B(n7372), .A(n7373), .Z(n7370) );
  AND U7922 ( .A(b[18]), .B(a[20]), .Z(n7369) );
  XNOR U7923 ( .A(n7374), .B(n7155), .Z(n7157) );
  XOR U7924 ( .A(n7375), .B(n7376), .Z(n7155) );
  ANDN U7925 ( .B(n7377), .A(n7378), .Z(n7375) );
  AND U7926 ( .A(b[17]), .B(a[21]), .Z(n7374) );
  XNOR U7927 ( .A(n7379), .B(n7160), .Z(n7162) );
  XOR U7928 ( .A(n7380), .B(n7381), .Z(n7160) );
  ANDN U7929 ( .B(n7382), .A(n7383), .Z(n7380) );
  AND U7930 ( .A(b[16]), .B(a[22]), .Z(n7379) );
  XOR U7931 ( .A(n7384), .B(n7385), .Z(n7164) );
  AND U7932 ( .A(n7386), .B(n7387), .Z(n7384) );
  XNOR U7933 ( .A(n7388), .B(n7169), .Z(n7171) );
  XOR U7934 ( .A(n7389), .B(n7390), .Z(n7169) );
  ANDN U7935 ( .B(n7391), .A(n7392), .Z(n7389) );
  AND U7936 ( .A(a[23]), .B(b[15]), .Z(n7388) );
  XOR U7937 ( .A(n7393), .B(n7174), .Z(n7176) );
  XOR U7938 ( .A(n7394), .B(n7395), .Z(n7174) );
  ANDN U7939 ( .B(n7396), .A(n7397), .Z(n7394) );
  AND U7940 ( .A(b[13]), .B(a[25]), .Z(n7393) );
  XNOR U7941 ( .A(n7398), .B(n7179), .Z(n7181) );
  XOR U7942 ( .A(n7399), .B(n7400), .Z(n7179) );
  ANDN U7943 ( .B(n7401), .A(n7402), .Z(n7399) );
  AND U7944 ( .A(b[12]), .B(a[26]), .Z(n7398) );
  XNOR U7945 ( .A(n7403), .B(n7184), .Z(n7186) );
  XOR U7946 ( .A(n7404), .B(n7405), .Z(n7184) );
  ANDN U7947 ( .B(n7406), .A(n7407), .Z(n7404) );
  AND U7948 ( .A(b[11]), .B(a[27]), .Z(n7403) );
  XNOR U7949 ( .A(n7408), .B(n7189), .Z(n7191) );
  XOR U7950 ( .A(n7409), .B(n7410), .Z(n7189) );
  ANDN U7951 ( .B(n7411), .A(n7412), .Z(n7409) );
  AND U7952 ( .A(b[10]), .B(a[28]), .Z(n7408) );
  XOR U7953 ( .A(n7413), .B(n7414), .Z(n7193) );
  AND U7954 ( .A(n7415), .B(n7416), .Z(n7413) );
  XNOR U7955 ( .A(n7417), .B(n7198), .Z(n7200) );
  XOR U7956 ( .A(n7418), .B(n7419), .Z(n7198) );
  ANDN U7957 ( .B(n7420), .A(n7421), .Z(n7418) );
  AND U7958 ( .A(b[9]), .B(a[29]), .Z(n7417) );
  XOR U7959 ( .A(n7422), .B(n7203), .Z(n7205) );
  XOR U7960 ( .A(n7423), .B(n7424), .Z(n7203) );
  ANDN U7961 ( .B(n7425), .A(n7426), .Z(n7423) );
  AND U7962 ( .A(b[7]), .B(a[31]), .Z(n7422) );
  XNOR U7963 ( .A(n7427), .B(n7208), .Z(n7210) );
  XOR U7964 ( .A(n7428), .B(n7429), .Z(n7208) );
  ANDN U7965 ( .B(n7430), .A(n7431), .Z(n7428) );
  AND U7966 ( .A(b[6]), .B(a[32]), .Z(n7427) );
  XNOR U7967 ( .A(n7432), .B(n7213), .Z(n7215) );
  XOR U7968 ( .A(n7433), .B(n7434), .Z(n7213) );
  ANDN U7969 ( .B(n7435), .A(n7436), .Z(n7433) );
  AND U7970 ( .A(b[5]), .B(a[33]), .Z(n7432) );
  XNOR U7971 ( .A(n7437), .B(n7218), .Z(n7220) );
  XOR U7972 ( .A(n7438), .B(n7439), .Z(n7218) );
  ANDN U7973 ( .B(n7440), .A(n7441), .Z(n7438) );
  AND U7974 ( .A(b[4]), .B(a[34]), .Z(n7437) );
  XNOR U7975 ( .A(n7442), .B(n7227), .Z(n7229) );
  XNOR U7976 ( .A(n7443), .B(n7444), .Z(n7227) );
  NOR U7977 ( .A(n7445), .B(n7446), .Z(n7443) );
  AND U7978 ( .A(b[3]), .B(a[35]), .Z(n7442) );
  NANDN U7979 ( .A(n7447), .B(n7448), .Z(n7230) );
  XNOR U7980 ( .A(n7449), .B(n7222), .Z(n7224) );
  XNOR U7981 ( .A(n7450), .B(n7451), .Z(n7222) );
  OR U7982 ( .A(n7452), .B(n7453), .Z(n7451) );
  AND U7983 ( .A(b[2]), .B(a[36]), .Z(n7449) );
  NAND U7984 ( .A(a[38]), .B(b[0]), .Z(n7011) );
  XNOR U7985 ( .A(n7447), .B(n7448), .Z(c[37]) );
  XOR U7986 ( .A(n7453), .B(n7452), .Z(n7448) );
  XOR U7987 ( .A(n7450), .B(n7454), .Z(n7452) );
  NAND U7988 ( .A(b[1]), .B(a[36]), .Z(n7454) );
  XOR U7989 ( .A(n7450), .B(n7446), .Z(n7455) );
  XOR U7990 ( .A(n7456), .B(n7444), .Z(n7446) );
  AND U7991 ( .A(b[2]), .B(a[35]), .Z(n7456) );
  ANDN U7992 ( .B(n7457), .A(n7458), .Z(n7450) );
  XOR U7993 ( .A(n7444), .B(n7440), .Z(n7459) );
  XNOR U7994 ( .A(n7439), .B(n7435), .Z(n7460) );
  XNOR U7995 ( .A(n7434), .B(n7430), .Z(n7461) );
  XNOR U7996 ( .A(n7429), .B(n7425), .Z(n7462) );
  XNOR U7997 ( .A(n7416), .B(n7415), .Z(n7463) );
  XOR U7998 ( .A(n7464), .B(n7414), .Z(n7415) );
  AND U7999 ( .A(b[7]), .B(a[30]), .Z(n7464) );
  XNOR U8000 ( .A(n7414), .B(n7420), .Z(n7465) );
  XNOR U8001 ( .A(n7419), .B(n7411), .Z(n7466) );
  XNOR U8002 ( .A(n7410), .B(n7406), .Z(n7467) );
  XNOR U8003 ( .A(n7405), .B(n7401), .Z(n7468) );
  XNOR U8004 ( .A(n7400), .B(n7396), .Z(n7469) );
  XNOR U8005 ( .A(n7387), .B(n7386), .Z(n7470) );
  XOR U8006 ( .A(n7471), .B(n7385), .Z(n7386) );
  AND U8007 ( .A(b[13]), .B(a[24]), .Z(n7471) );
  XNOR U8008 ( .A(n7385), .B(n7391), .Z(n7472) );
  XNOR U8009 ( .A(n7390), .B(n7382), .Z(n7473) );
  XNOR U8010 ( .A(n7381), .B(n7377), .Z(n7474) );
  XNOR U8011 ( .A(n7376), .B(n7372), .Z(n7475) );
  XNOR U8012 ( .A(n7371), .B(n7367), .Z(n7476) );
  XNOR U8013 ( .A(n7358), .B(n7357), .Z(n7477) );
  XOR U8014 ( .A(n7478), .B(n7356), .Z(n7357) );
  AND U8015 ( .A(b[19]), .B(a[18]), .Z(n7478) );
  XNOR U8016 ( .A(n7356), .B(n7362), .Z(n7479) );
  XNOR U8017 ( .A(n7361), .B(n7353), .Z(n7480) );
  XNOR U8018 ( .A(n7352), .B(n7348), .Z(n7481) );
  XNOR U8019 ( .A(n7347), .B(n7343), .Z(n7482) );
  XNOR U8020 ( .A(n7342), .B(n7338), .Z(n7483) );
  XNOR U8021 ( .A(n7329), .B(n7328), .Z(n7484) );
  XOR U8022 ( .A(n7485), .B(n7327), .Z(n7328) );
  AND U8023 ( .A(b[25]), .B(a[12]), .Z(n7485) );
  XNOR U8024 ( .A(n7327), .B(n7333), .Z(n7486) );
  XNOR U8025 ( .A(n7332), .B(n7324), .Z(n7487) );
  XNOR U8026 ( .A(n7323), .B(n7319), .Z(n7488) );
  XNOR U8027 ( .A(n7318), .B(n7314), .Z(n7489) );
  XNOR U8028 ( .A(n7313), .B(n7309), .Z(n7490) );
  XNOR U8029 ( .A(n7300), .B(n7299), .Z(n7491) );
  XOR U8030 ( .A(n7492), .B(n7298), .Z(n7299) );
  AND U8031 ( .A(a[6]), .B(b[31]), .Z(n7492) );
  XNOR U8032 ( .A(n7298), .B(n7304), .Z(n7493) );
  XNOR U8033 ( .A(n7303), .B(n7295), .Z(n7494) );
  XNOR U8034 ( .A(n7294), .B(n7290), .Z(n7495) );
  XNOR U8035 ( .A(n7289), .B(n7285), .Z(n7496) );
  XNOR U8036 ( .A(n7284), .B(n7280), .Z(n7497) );
  XNOR U8037 ( .A(n7498), .B(n7279), .Z(n7280) );
  AND U8038 ( .A(a[0]), .B(b[37]), .Z(n7498) );
  XOR U8039 ( .A(n7499), .B(n7279), .Z(n7281) );
  XNOR U8040 ( .A(n7500), .B(n7501), .Z(n7279) );
  ANDN U8041 ( .B(n7502), .A(n7503), .Z(n7500) );
  AND U8042 ( .A(a[1]), .B(b[36]), .Z(n7499) );
  XNOR U8043 ( .A(n7504), .B(n7284), .Z(n7286) );
  XOR U8044 ( .A(n7505), .B(n7506), .Z(n7284) );
  ANDN U8045 ( .B(n7507), .A(n7508), .Z(n7505) );
  AND U8046 ( .A(a[2]), .B(b[35]), .Z(n7504) );
  XNOR U8047 ( .A(n7509), .B(n7289), .Z(n7291) );
  XOR U8048 ( .A(n7510), .B(n7511), .Z(n7289) );
  ANDN U8049 ( .B(n7512), .A(n7513), .Z(n7510) );
  AND U8050 ( .A(a[3]), .B(b[34]), .Z(n7509) );
  XNOR U8051 ( .A(n7514), .B(n7294), .Z(n7296) );
  XOR U8052 ( .A(n7515), .B(n7516), .Z(n7294) );
  ANDN U8053 ( .B(n7517), .A(n7518), .Z(n7515) );
  AND U8054 ( .A(a[4]), .B(b[33]), .Z(n7514) );
  XOR U8055 ( .A(n7519), .B(n7520), .Z(n7298) );
  AND U8056 ( .A(n7521), .B(n7522), .Z(n7519) );
  XNOR U8057 ( .A(n7523), .B(n7303), .Z(n7305) );
  XOR U8058 ( .A(n7524), .B(n7525), .Z(n7303) );
  ANDN U8059 ( .B(n7526), .A(n7527), .Z(n7524) );
  AND U8060 ( .A(a[5]), .B(b[32]), .Z(n7523) );
  XOR U8061 ( .A(n7528), .B(n7308), .Z(n7310) );
  XOR U8062 ( .A(n7529), .B(n7530), .Z(n7308) );
  ANDN U8063 ( .B(n7531), .A(n7532), .Z(n7529) );
  AND U8064 ( .A(a[7]), .B(b[30]), .Z(n7528) );
  XNOR U8065 ( .A(n7533), .B(n7313), .Z(n7315) );
  XOR U8066 ( .A(n7534), .B(n7535), .Z(n7313) );
  ANDN U8067 ( .B(n7536), .A(n7537), .Z(n7534) );
  AND U8068 ( .A(a[8]), .B(b[29]), .Z(n7533) );
  XNOR U8069 ( .A(n7538), .B(n7318), .Z(n7320) );
  XOR U8070 ( .A(n7539), .B(n7540), .Z(n7318) );
  ANDN U8071 ( .B(n7541), .A(n7542), .Z(n7539) );
  AND U8072 ( .A(a[9]), .B(b[28]), .Z(n7538) );
  XNOR U8073 ( .A(n7543), .B(n7323), .Z(n7325) );
  XOR U8074 ( .A(n7544), .B(n7545), .Z(n7323) );
  ANDN U8075 ( .B(n7546), .A(n7547), .Z(n7544) );
  AND U8076 ( .A(a[10]), .B(b[27]), .Z(n7543) );
  XOR U8077 ( .A(n7548), .B(n7549), .Z(n7327) );
  AND U8078 ( .A(n7550), .B(n7551), .Z(n7548) );
  XNOR U8079 ( .A(n7552), .B(n7332), .Z(n7334) );
  XOR U8080 ( .A(n7553), .B(n7554), .Z(n7332) );
  ANDN U8081 ( .B(n7555), .A(n7556), .Z(n7553) );
  AND U8082 ( .A(b[26]), .B(a[11]), .Z(n7552) );
  XOR U8083 ( .A(n7557), .B(n7337), .Z(n7339) );
  XOR U8084 ( .A(n7558), .B(n7559), .Z(n7337) );
  ANDN U8085 ( .B(n7560), .A(n7561), .Z(n7558) );
  AND U8086 ( .A(b[24]), .B(a[13]), .Z(n7557) );
  XNOR U8087 ( .A(n7562), .B(n7342), .Z(n7344) );
  XOR U8088 ( .A(n7563), .B(n7564), .Z(n7342) );
  ANDN U8089 ( .B(n7565), .A(n7566), .Z(n7563) );
  AND U8090 ( .A(b[23]), .B(a[14]), .Z(n7562) );
  XNOR U8091 ( .A(n7567), .B(n7347), .Z(n7349) );
  XOR U8092 ( .A(n7568), .B(n7569), .Z(n7347) );
  ANDN U8093 ( .B(n7570), .A(n7571), .Z(n7568) );
  AND U8094 ( .A(b[22]), .B(a[15]), .Z(n7567) );
  XNOR U8095 ( .A(n7572), .B(n7352), .Z(n7354) );
  XOR U8096 ( .A(n7573), .B(n7574), .Z(n7352) );
  ANDN U8097 ( .B(n7575), .A(n7576), .Z(n7573) );
  AND U8098 ( .A(a[16]), .B(b[21]), .Z(n7572) );
  XOR U8099 ( .A(n7577), .B(n7578), .Z(n7356) );
  AND U8100 ( .A(n7579), .B(n7580), .Z(n7577) );
  XNOR U8101 ( .A(n7581), .B(n7361), .Z(n7363) );
  XOR U8102 ( .A(n7582), .B(n7583), .Z(n7361) );
  ANDN U8103 ( .B(n7584), .A(n7585), .Z(n7582) );
  AND U8104 ( .A(b[20]), .B(a[17]), .Z(n7581) );
  XOR U8105 ( .A(n7586), .B(n7366), .Z(n7368) );
  XOR U8106 ( .A(n7587), .B(n7588), .Z(n7366) );
  ANDN U8107 ( .B(n7589), .A(n7590), .Z(n7587) );
  AND U8108 ( .A(b[18]), .B(a[19]), .Z(n7586) );
  XNOR U8109 ( .A(n7591), .B(n7371), .Z(n7373) );
  XOR U8110 ( .A(n7592), .B(n7593), .Z(n7371) );
  ANDN U8111 ( .B(n7594), .A(n7595), .Z(n7592) );
  AND U8112 ( .A(b[17]), .B(a[20]), .Z(n7591) );
  XNOR U8113 ( .A(n7596), .B(n7376), .Z(n7378) );
  XOR U8114 ( .A(n7597), .B(n7598), .Z(n7376) );
  ANDN U8115 ( .B(n7599), .A(n7600), .Z(n7597) );
  AND U8116 ( .A(b[16]), .B(a[21]), .Z(n7596) );
  XNOR U8117 ( .A(n7601), .B(n7381), .Z(n7383) );
  XOR U8118 ( .A(n7602), .B(n7603), .Z(n7381) );
  ANDN U8119 ( .B(n7604), .A(n7605), .Z(n7602) );
  AND U8120 ( .A(a[22]), .B(b[15]), .Z(n7601) );
  XOR U8121 ( .A(n7606), .B(n7607), .Z(n7385) );
  AND U8122 ( .A(n7608), .B(n7609), .Z(n7606) );
  XNOR U8123 ( .A(n7610), .B(n7390), .Z(n7392) );
  XOR U8124 ( .A(n7611), .B(n7612), .Z(n7390) );
  ANDN U8125 ( .B(n7613), .A(n7614), .Z(n7611) );
  AND U8126 ( .A(b[14]), .B(a[23]), .Z(n7610) );
  XOR U8127 ( .A(n7615), .B(n7395), .Z(n7397) );
  XOR U8128 ( .A(n7616), .B(n7617), .Z(n7395) );
  ANDN U8129 ( .B(n7618), .A(n7619), .Z(n7616) );
  AND U8130 ( .A(b[12]), .B(a[25]), .Z(n7615) );
  XNOR U8131 ( .A(n7620), .B(n7400), .Z(n7402) );
  XOR U8132 ( .A(n7621), .B(n7622), .Z(n7400) );
  ANDN U8133 ( .B(n7623), .A(n7624), .Z(n7621) );
  AND U8134 ( .A(b[11]), .B(a[26]), .Z(n7620) );
  XNOR U8135 ( .A(n7625), .B(n7405), .Z(n7407) );
  XOR U8136 ( .A(n7626), .B(n7627), .Z(n7405) );
  ANDN U8137 ( .B(n7628), .A(n7629), .Z(n7626) );
  AND U8138 ( .A(b[10]), .B(a[27]), .Z(n7625) );
  XNOR U8139 ( .A(n7630), .B(n7410), .Z(n7412) );
  XOR U8140 ( .A(n7631), .B(n7632), .Z(n7410) );
  ANDN U8141 ( .B(n7633), .A(n7634), .Z(n7631) );
  AND U8142 ( .A(b[9]), .B(a[28]), .Z(n7630) );
  XOR U8143 ( .A(n7635), .B(n7636), .Z(n7414) );
  AND U8144 ( .A(n7637), .B(n7638), .Z(n7635) );
  XNOR U8145 ( .A(n7639), .B(n7419), .Z(n7421) );
  XOR U8146 ( .A(n7640), .B(n7641), .Z(n7419) );
  ANDN U8147 ( .B(n7642), .A(n7643), .Z(n7640) );
  AND U8148 ( .A(b[8]), .B(a[29]), .Z(n7639) );
  XOR U8149 ( .A(n7644), .B(n7424), .Z(n7426) );
  XOR U8150 ( .A(n7645), .B(n7646), .Z(n7424) );
  ANDN U8151 ( .B(n7647), .A(n7648), .Z(n7645) );
  AND U8152 ( .A(b[6]), .B(a[31]), .Z(n7644) );
  XNOR U8153 ( .A(n7649), .B(n7429), .Z(n7431) );
  XOR U8154 ( .A(n7650), .B(n7651), .Z(n7429) );
  ANDN U8155 ( .B(n7652), .A(n7653), .Z(n7650) );
  AND U8156 ( .A(b[5]), .B(a[32]), .Z(n7649) );
  XNOR U8157 ( .A(n7654), .B(n7434), .Z(n7436) );
  XOR U8158 ( .A(n7655), .B(n7656), .Z(n7434) );
  ANDN U8159 ( .B(n7657), .A(n7658), .Z(n7655) );
  AND U8160 ( .A(b[4]), .B(a[33]), .Z(n7654) );
  XNOR U8161 ( .A(n7659), .B(n7660), .Z(n7444) );
  NANDN U8162 ( .A(n7661), .B(n7662), .Z(n7660) );
  XNOR U8163 ( .A(n7663), .B(n7439), .Z(n7441) );
  XNOR U8164 ( .A(n7664), .B(n7665), .Z(n7439) );
  AND U8165 ( .A(n7666), .B(n7667), .Z(n7664) );
  AND U8166 ( .A(b[3]), .B(a[34]), .Z(n7663) );
  NAND U8167 ( .A(a[37]), .B(b[0]), .Z(n7447) );
  XNOR U8168 ( .A(n7458), .B(n7457), .Z(c[36]) );
  XNOR U8169 ( .A(n7661), .B(n7662), .Z(n7457) );
  XOR U8170 ( .A(n7659), .B(n7668), .Z(n7662) );
  NAND U8171 ( .A(b[1]), .B(a[35]), .Z(n7668) );
  XOR U8172 ( .A(n7667), .B(n7669), .Z(n7661) );
  XOR U8173 ( .A(n7659), .B(n7666), .Z(n7669) );
  XNOR U8174 ( .A(n7670), .B(n7665), .Z(n7666) );
  AND U8175 ( .A(b[2]), .B(a[34]), .Z(n7670) );
  NANDN U8176 ( .A(n7671), .B(n7672), .Z(n7659) );
  XOR U8177 ( .A(n7665), .B(n7657), .Z(n7673) );
  XNOR U8178 ( .A(n7656), .B(n7652), .Z(n7674) );
  XNOR U8179 ( .A(n7651), .B(n7647), .Z(n7675) );
  XNOR U8180 ( .A(n7638), .B(n7637), .Z(n7676) );
  XOR U8181 ( .A(n7677), .B(n7636), .Z(n7637) );
  AND U8182 ( .A(b[6]), .B(a[30]), .Z(n7677) );
  XNOR U8183 ( .A(n7636), .B(n7642), .Z(n7678) );
  XNOR U8184 ( .A(n7641), .B(n7633), .Z(n7679) );
  XNOR U8185 ( .A(n7632), .B(n7628), .Z(n7680) );
  XNOR U8186 ( .A(n7627), .B(n7623), .Z(n7681) );
  XNOR U8187 ( .A(n7622), .B(n7618), .Z(n7682) );
  XNOR U8188 ( .A(n7609), .B(n7608), .Z(n7683) );
  XOR U8189 ( .A(n7684), .B(n7607), .Z(n7608) );
  AND U8190 ( .A(b[12]), .B(a[24]), .Z(n7684) );
  XNOR U8191 ( .A(n7607), .B(n7613), .Z(n7685) );
  XNOR U8192 ( .A(n7612), .B(n7604), .Z(n7686) );
  XNOR U8193 ( .A(n7603), .B(n7599), .Z(n7687) );
  XNOR U8194 ( .A(n7598), .B(n7594), .Z(n7688) );
  XNOR U8195 ( .A(n7593), .B(n7589), .Z(n7689) );
  XNOR U8196 ( .A(n7580), .B(n7579), .Z(n7690) );
  XOR U8197 ( .A(n7691), .B(n7578), .Z(n7579) );
  AND U8198 ( .A(b[18]), .B(a[18]), .Z(n7691) );
  XNOR U8199 ( .A(n7578), .B(n7584), .Z(n7692) );
  XNOR U8200 ( .A(n7583), .B(n7575), .Z(n7693) );
  XNOR U8201 ( .A(n7574), .B(n7570), .Z(n7694) );
  XNOR U8202 ( .A(n7569), .B(n7565), .Z(n7695) );
  XNOR U8203 ( .A(n7564), .B(n7560), .Z(n7696) );
  XNOR U8204 ( .A(n7551), .B(n7550), .Z(n7697) );
  XOR U8205 ( .A(n7698), .B(n7549), .Z(n7550) );
  AND U8206 ( .A(b[24]), .B(a[12]), .Z(n7698) );
  XNOR U8207 ( .A(n7549), .B(n7555), .Z(n7699) );
  XNOR U8208 ( .A(n7554), .B(n7546), .Z(n7700) );
  XNOR U8209 ( .A(n7545), .B(n7541), .Z(n7701) );
  XNOR U8210 ( .A(n7540), .B(n7536), .Z(n7702) );
  XNOR U8211 ( .A(n7535), .B(n7531), .Z(n7703) );
  XNOR U8212 ( .A(n7522), .B(n7521), .Z(n7704) );
  XOR U8213 ( .A(n7705), .B(n7520), .Z(n7521) );
  AND U8214 ( .A(a[6]), .B(b[30]), .Z(n7705) );
  XNOR U8215 ( .A(n7520), .B(n7526), .Z(n7706) );
  XNOR U8216 ( .A(n7525), .B(n7517), .Z(n7707) );
  XNOR U8217 ( .A(n7516), .B(n7512), .Z(n7708) );
  XNOR U8218 ( .A(n7511), .B(n7507), .Z(n7709) );
  XNOR U8219 ( .A(n7506), .B(n7502), .Z(n7710) );
  XOR U8220 ( .A(n7711), .B(n7501), .Z(n7502) );
  AND U8221 ( .A(a[0]), .B(b[36]), .Z(n7711) );
  XNOR U8222 ( .A(n7712), .B(n7501), .Z(n7503) );
  XNOR U8223 ( .A(n7713), .B(n7714), .Z(n7501) );
  ANDN U8224 ( .B(n7715), .A(n7716), .Z(n7713) );
  AND U8225 ( .A(a[1]), .B(b[35]), .Z(n7712) );
  XNOR U8226 ( .A(n7717), .B(n7506), .Z(n7508) );
  XOR U8227 ( .A(n7718), .B(n7719), .Z(n7506) );
  ANDN U8228 ( .B(n7720), .A(n7721), .Z(n7718) );
  AND U8229 ( .A(a[2]), .B(b[34]), .Z(n7717) );
  XNOR U8230 ( .A(n7722), .B(n7511), .Z(n7513) );
  XOR U8231 ( .A(n7723), .B(n7724), .Z(n7511) );
  ANDN U8232 ( .B(n7725), .A(n7726), .Z(n7723) );
  AND U8233 ( .A(a[3]), .B(b[33]), .Z(n7722) );
  XNOR U8234 ( .A(n7727), .B(n7516), .Z(n7518) );
  XOR U8235 ( .A(n7728), .B(n7729), .Z(n7516) );
  ANDN U8236 ( .B(n7730), .A(n7731), .Z(n7728) );
  AND U8237 ( .A(a[4]), .B(b[32]), .Z(n7727) );
  XOR U8238 ( .A(n7732), .B(n7733), .Z(n7520) );
  AND U8239 ( .A(n7734), .B(n7735), .Z(n7732) );
  XNOR U8240 ( .A(n7736), .B(n7525), .Z(n7527) );
  XOR U8241 ( .A(n7737), .B(n7738), .Z(n7525) );
  ANDN U8242 ( .B(n7739), .A(n7740), .Z(n7737) );
  AND U8243 ( .A(a[5]), .B(b[31]), .Z(n7736) );
  XOR U8244 ( .A(n7741), .B(n7530), .Z(n7532) );
  XOR U8245 ( .A(n7742), .B(n7743), .Z(n7530) );
  ANDN U8246 ( .B(n7744), .A(n7745), .Z(n7742) );
  AND U8247 ( .A(a[7]), .B(b[29]), .Z(n7741) );
  XNOR U8248 ( .A(n7746), .B(n7535), .Z(n7537) );
  XOR U8249 ( .A(n7747), .B(n7748), .Z(n7535) );
  ANDN U8250 ( .B(n7749), .A(n7750), .Z(n7747) );
  AND U8251 ( .A(a[8]), .B(b[28]), .Z(n7746) );
  XNOR U8252 ( .A(n7751), .B(n7540), .Z(n7542) );
  XOR U8253 ( .A(n7752), .B(n7753), .Z(n7540) );
  ANDN U8254 ( .B(n7754), .A(n7755), .Z(n7752) );
  AND U8255 ( .A(a[9]), .B(b[27]), .Z(n7751) );
  XNOR U8256 ( .A(n7756), .B(n7545), .Z(n7547) );
  XOR U8257 ( .A(n7757), .B(n7758), .Z(n7545) );
  ANDN U8258 ( .B(n7759), .A(n7760), .Z(n7757) );
  AND U8259 ( .A(b[26]), .B(a[10]), .Z(n7756) );
  XOR U8260 ( .A(n7761), .B(n7762), .Z(n7549) );
  AND U8261 ( .A(n7763), .B(n7764), .Z(n7761) );
  XNOR U8262 ( .A(n7765), .B(n7554), .Z(n7556) );
  XOR U8263 ( .A(n7766), .B(n7767), .Z(n7554) );
  ANDN U8264 ( .B(n7768), .A(n7769), .Z(n7766) );
  AND U8265 ( .A(b[25]), .B(a[11]), .Z(n7765) );
  XOR U8266 ( .A(n7770), .B(n7559), .Z(n7561) );
  XOR U8267 ( .A(n7771), .B(n7772), .Z(n7559) );
  ANDN U8268 ( .B(n7773), .A(n7774), .Z(n7771) );
  AND U8269 ( .A(b[23]), .B(a[13]), .Z(n7770) );
  XNOR U8270 ( .A(n7775), .B(n7564), .Z(n7566) );
  XOR U8271 ( .A(n7776), .B(n7777), .Z(n7564) );
  ANDN U8272 ( .B(n7778), .A(n7779), .Z(n7776) );
  AND U8273 ( .A(b[22]), .B(a[14]), .Z(n7775) );
  XNOR U8274 ( .A(n7780), .B(n7569), .Z(n7571) );
  XOR U8275 ( .A(n7781), .B(n7782), .Z(n7569) );
  ANDN U8276 ( .B(n7783), .A(n7784), .Z(n7781) );
  AND U8277 ( .A(a[15]), .B(b[21]), .Z(n7780) );
  XNOR U8278 ( .A(n7785), .B(n7574), .Z(n7576) );
  XOR U8279 ( .A(n7786), .B(n7787), .Z(n7574) );
  ANDN U8280 ( .B(n7788), .A(n7789), .Z(n7786) );
  AND U8281 ( .A(b[20]), .B(a[16]), .Z(n7785) );
  XOR U8282 ( .A(n7790), .B(n7791), .Z(n7578) );
  AND U8283 ( .A(n7792), .B(n7793), .Z(n7790) );
  XNOR U8284 ( .A(n7794), .B(n7583), .Z(n7585) );
  XOR U8285 ( .A(n7795), .B(n7796), .Z(n7583) );
  ANDN U8286 ( .B(n7797), .A(n7798), .Z(n7795) );
  AND U8287 ( .A(b[19]), .B(a[17]), .Z(n7794) );
  XOR U8288 ( .A(n7799), .B(n7588), .Z(n7590) );
  XOR U8289 ( .A(n7800), .B(n7801), .Z(n7588) );
  ANDN U8290 ( .B(n7802), .A(n7803), .Z(n7800) );
  AND U8291 ( .A(b[17]), .B(a[19]), .Z(n7799) );
  XNOR U8292 ( .A(n7804), .B(n7593), .Z(n7595) );
  XOR U8293 ( .A(n7805), .B(n7806), .Z(n7593) );
  ANDN U8294 ( .B(n7807), .A(n7808), .Z(n7805) );
  AND U8295 ( .A(b[16]), .B(a[20]), .Z(n7804) );
  XNOR U8296 ( .A(n7809), .B(n7598), .Z(n7600) );
  XOR U8297 ( .A(n7810), .B(n7811), .Z(n7598) );
  ANDN U8298 ( .B(n7812), .A(n7813), .Z(n7810) );
  AND U8299 ( .A(a[21]), .B(b[15]), .Z(n7809) );
  XNOR U8300 ( .A(n7814), .B(n7603), .Z(n7605) );
  XOR U8301 ( .A(n7815), .B(n7816), .Z(n7603) );
  ANDN U8302 ( .B(n7817), .A(n7818), .Z(n7815) );
  AND U8303 ( .A(b[14]), .B(a[22]), .Z(n7814) );
  XOR U8304 ( .A(n7819), .B(n7820), .Z(n7607) );
  AND U8305 ( .A(n7821), .B(n7822), .Z(n7819) );
  XNOR U8306 ( .A(n7823), .B(n7612), .Z(n7614) );
  XOR U8307 ( .A(n7824), .B(n7825), .Z(n7612) );
  ANDN U8308 ( .B(n7826), .A(n7827), .Z(n7824) );
  AND U8309 ( .A(b[13]), .B(a[23]), .Z(n7823) );
  XOR U8310 ( .A(n7828), .B(n7617), .Z(n7619) );
  XOR U8311 ( .A(n7829), .B(n7830), .Z(n7617) );
  ANDN U8312 ( .B(n7831), .A(n7832), .Z(n7829) );
  AND U8313 ( .A(b[11]), .B(a[25]), .Z(n7828) );
  XNOR U8314 ( .A(n7833), .B(n7622), .Z(n7624) );
  XOR U8315 ( .A(n7834), .B(n7835), .Z(n7622) );
  ANDN U8316 ( .B(n7836), .A(n7837), .Z(n7834) );
  AND U8317 ( .A(b[10]), .B(a[26]), .Z(n7833) );
  XNOR U8318 ( .A(n7838), .B(n7627), .Z(n7629) );
  XOR U8319 ( .A(n7839), .B(n7840), .Z(n7627) );
  ANDN U8320 ( .B(n7841), .A(n7842), .Z(n7839) );
  AND U8321 ( .A(b[9]), .B(a[27]), .Z(n7838) );
  XNOR U8322 ( .A(n7843), .B(n7632), .Z(n7634) );
  XOR U8323 ( .A(n7844), .B(n7845), .Z(n7632) );
  ANDN U8324 ( .B(n7846), .A(n7847), .Z(n7844) );
  AND U8325 ( .A(b[8]), .B(a[28]), .Z(n7843) );
  XOR U8326 ( .A(n7848), .B(n7849), .Z(n7636) );
  AND U8327 ( .A(n7850), .B(n7851), .Z(n7848) );
  XNOR U8328 ( .A(n7852), .B(n7641), .Z(n7643) );
  XOR U8329 ( .A(n7853), .B(n7854), .Z(n7641) );
  ANDN U8330 ( .B(n7855), .A(n7856), .Z(n7853) );
  AND U8331 ( .A(b[7]), .B(a[29]), .Z(n7852) );
  XOR U8332 ( .A(n7857), .B(n7646), .Z(n7648) );
  XOR U8333 ( .A(n7858), .B(n7859), .Z(n7646) );
  ANDN U8334 ( .B(n7860), .A(n7861), .Z(n7858) );
  AND U8335 ( .A(b[5]), .B(a[31]), .Z(n7857) );
  XNOR U8336 ( .A(n7862), .B(n7651), .Z(n7653) );
  XOR U8337 ( .A(n7863), .B(n7864), .Z(n7651) );
  ANDN U8338 ( .B(n7865), .A(n7866), .Z(n7863) );
  AND U8339 ( .A(b[4]), .B(a[32]), .Z(n7862) );
  XNOR U8340 ( .A(n7867), .B(n7868), .Z(n7665) );
  NANDN U8341 ( .A(n7869), .B(n7870), .Z(n7868) );
  XNOR U8342 ( .A(n7871), .B(n7656), .Z(n7658) );
  XNOR U8343 ( .A(n7872), .B(n7873), .Z(n7656) );
  AND U8344 ( .A(n7874), .B(n7875), .Z(n7872) );
  AND U8345 ( .A(b[3]), .B(a[33]), .Z(n7871) );
  NAND U8346 ( .A(a[36]), .B(b[0]), .Z(n7458) );
  XNOR U8347 ( .A(n7671), .B(n7672), .Z(c[35]) );
  XNOR U8348 ( .A(n7869), .B(n7870), .Z(n7672) );
  XOR U8349 ( .A(n7867), .B(n7876), .Z(n7870) );
  NAND U8350 ( .A(b[1]), .B(a[34]), .Z(n7876) );
  XOR U8351 ( .A(n7875), .B(n7877), .Z(n7869) );
  XOR U8352 ( .A(n7867), .B(n7874), .Z(n7877) );
  XNOR U8353 ( .A(n7878), .B(n7873), .Z(n7874) );
  AND U8354 ( .A(b[2]), .B(a[33]), .Z(n7878) );
  NANDN U8355 ( .A(n7879), .B(n7880), .Z(n7867) );
  XOR U8356 ( .A(n7873), .B(n7865), .Z(n7881) );
  XNOR U8357 ( .A(n7864), .B(n7860), .Z(n7882) );
  XNOR U8358 ( .A(n7851), .B(n7850), .Z(n7883) );
  XOR U8359 ( .A(n7884), .B(n7849), .Z(n7850) );
  AND U8360 ( .A(b[5]), .B(a[30]), .Z(n7884) );
  XNOR U8361 ( .A(n7849), .B(n7855), .Z(n7885) );
  XNOR U8362 ( .A(n7854), .B(n7846), .Z(n7886) );
  XNOR U8363 ( .A(n7845), .B(n7841), .Z(n7887) );
  XNOR U8364 ( .A(n7840), .B(n7836), .Z(n7888) );
  XNOR U8365 ( .A(n7835), .B(n7831), .Z(n7889) );
  XNOR U8366 ( .A(n7822), .B(n7821), .Z(n7890) );
  XOR U8367 ( .A(n7891), .B(n7820), .Z(n7821) );
  AND U8368 ( .A(b[11]), .B(a[24]), .Z(n7891) );
  XNOR U8369 ( .A(n7820), .B(n7826), .Z(n7892) );
  XNOR U8370 ( .A(n7825), .B(n7817), .Z(n7893) );
  XNOR U8371 ( .A(n7816), .B(n7812), .Z(n7894) );
  XNOR U8372 ( .A(n7811), .B(n7807), .Z(n7895) );
  XNOR U8373 ( .A(n7806), .B(n7802), .Z(n7896) );
  XNOR U8374 ( .A(n7793), .B(n7792), .Z(n7897) );
  XOR U8375 ( .A(n7898), .B(n7791), .Z(n7792) );
  AND U8376 ( .A(b[17]), .B(a[18]), .Z(n7898) );
  XNOR U8377 ( .A(n7791), .B(n7797), .Z(n7899) );
  XNOR U8378 ( .A(n7796), .B(n7788), .Z(n7900) );
  XNOR U8379 ( .A(n7787), .B(n7783), .Z(n7901) );
  XNOR U8380 ( .A(n7782), .B(n7778), .Z(n7902) );
  XNOR U8381 ( .A(n7777), .B(n7773), .Z(n7903) );
  XNOR U8382 ( .A(n7764), .B(n7763), .Z(n7904) );
  XOR U8383 ( .A(n7905), .B(n7762), .Z(n7763) );
  AND U8384 ( .A(b[23]), .B(a[12]), .Z(n7905) );
  XNOR U8385 ( .A(n7762), .B(n7768), .Z(n7906) );
  XNOR U8386 ( .A(n7767), .B(n7759), .Z(n7907) );
  XNOR U8387 ( .A(n7758), .B(n7754), .Z(n7908) );
  XNOR U8388 ( .A(n7753), .B(n7749), .Z(n7909) );
  XNOR U8389 ( .A(n7748), .B(n7744), .Z(n7910) );
  XNOR U8390 ( .A(n7735), .B(n7734), .Z(n7911) );
  XOR U8391 ( .A(n7912), .B(n7733), .Z(n7734) );
  AND U8392 ( .A(a[6]), .B(b[29]), .Z(n7912) );
  XNOR U8393 ( .A(n7733), .B(n7739), .Z(n7913) );
  XNOR U8394 ( .A(n7738), .B(n7730), .Z(n7914) );
  XNOR U8395 ( .A(n7729), .B(n7725), .Z(n7915) );
  XNOR U8396 ( .A(n7724), .B(n7720), .Z(n7916) );
  XNOR U8397 ( .A(n7719), .B(n7715), .Z(n7917) );
  XNOR U8398 ( .A(n7918), .B(n7714), .Z(n7715) );
  AND U8399 ( .A(a[0]), .B(b[35]), .Z(n7918) );
  XOR U8400 ( .A(n7919), .B(n7714), .Z(n7716) );
  XNOR U8401 ( .A(n7920), .B(n7921), .Z(n7714) );
  ANDN U8402 ( .B(n7922), .A(n7923), .Z(n7920) );
  AND U8403 ( .A(a[1]), .B(b[34]), .Z(n7919) );
  XNOR U8404 ( .A(n7924), .B(n7719), .Z(n7721) );
  XOR U8405 ( .A(n7925), .B(n7926), .Z(n7719) );
  ANDN U8406 ( .B(n7927), .A(n7928), .Z(n7925) );
  AND U8407 ( .A(a[2]), .B(b[33]), .Z(n7924) );
  XNOR U8408 ( .A(n7929), .B(n7724), .Z(n7726) );
  XOR U8409 ( .A(n7930), .B(n7931), .Z(n7724) );
  ANDN U8410 ( .B(n7932), .A(n7933), .Z(n7930) );
  AND U8411 ( .A(a[3]), .B(b[32]), .Z(n7929) );
  XNOR U8412 ( .A(n7934), .B(n7729), .Z(n7731) );
  XOR U8413 ( .A(n7935), .B(n7936), .Z(n7729) );
  ANDN U8414 ( .B(n7937), .A(n7938), .Z(n7935) );
  AND U8415 ( .A(a[4]), .B(b[31]), .Z(n7934) );
  XOR U8416 ( .A(n7939), .B(n7940), .Z(n7733) );
  AND U8417 ( .A(n7941), .B(n7942), .Z(n7939) );
  XNOR U8418 ( .A(n7943), .B(n7738), .Z(n7740) );
  XOR U8419 ( .A(n7944), .B(n7945), .Z(n7738) );
  ANDN U8420 ( .B(n7946), .A(n7947), .Z(n7944) );
  AND U8421 ( .A(a[5]), .B(b[30]), .Z(n7943) );
  XOR U8422 ( .A(n7948), .B(n7743), .Z(n7745) );
  XOR U8423 ( .A(n7949), .B(n7950), .Z(n7743) );
  ANDN U8424 ( .B(n7951), .A(n7952), .Z(n7949) );
  AND U8425 ( .A(a[7]), .B(b[28]), .Z(n7948) );
  XNOR U8426 ( .A(n7953), .B(n7748), .Z(n7750) );
  XOR U8427 ( .A(n7954), .B(n7955), .Z(n7748) );
  ANDN U8428 ( .B(n7956), .A(n7957), .Z(n7954) );
  AND U8429 ( .A(a[8]), .B(b[27]), .Z(n7953) );
  XNOR U8430 ( .A(n7958), .B(n7753), .Z(n7755) );
  XOR U8431 ( .A(n7959), .B(n7960), .Z(n7753) );
  ANDN U8432 ( .B(n7961), .A(n7962), .Z(n7959) );
  AND U8433 ( .A(a[9]), .B(b[26]), .Z(n7958) );
  XNOR U8434 ( .A(n7963), .B(n7758), .Z(n7760) );
  XOR U8435 ( .A(n7964), .B(n7965), .Z(n7758) );
  ANDN U8436 ( .B(n7966), .A(n7967), .Z(n7964) );
  AND U8437 ( .A(b[25]), .B(a[10]), .Z(n7963) );
  XOR U8438 ( .A(n7968), .B(n7969), .Z(n7762) );
  AND U8439 ( .A(n7970), .B(n7971), .Z(n7968) );
  XNOR U8440 ( .A(n7972), .B(n7767), .Z(n7769) );
  XOR U8441 ( .A(n7973), .B(n7974), .Z(n7767) );
  ANDN U8442 ( .B(n7975), .A(n7976), .Z(n7973) );
  AND U8443 ( .A(b[24]), .B(a[11]), .Z(n7972) );
  XOR U8444 ( .A(n7977), .B(n7772), .Z(n7774) );
  XOR U8445 ( .A(n7978), .B(n7979), .Z(n7772) );
  ANDN U8446 ( .B(n7980), .A(n7981), .Z(n7978) );
  AND U8447 ( .A(b[22]), .B(a[13]), .Z(n7977) );
  XNOR U8448 ( .A(n7982), .B(n7777), .Z(n7779) );
  XOR U8449 ( .A(n7983), .B(n7984), .Z(n7777) );
  ANDN U8450 ( .B(n7985), .A(n7986), .Z(n7983) );
  AND U8451 ( .A(a[14]), .B(b[21]), .Z(n7982) );
  XNOR U8452 ( .A(n7987), .B(n7782), .Z(n7784) );
  XOR U8453 ( .A(n7988), .B(n7989), .Z(n7782) );
  ANDN U8454 ( .B(n7990), .A(n7991), .Z(n7988) );
  AND U8455 ( .A(b[20]), .B(a[15]), .Z(n7987) );
  XNOR U8456 ( .A(n7992), .B(n7787), .Z(n7789) );
  XOR U8457 ( .A(n7993), .B(n7994), .Z(n7787) );
  ANDN U8458 ( .B(n7995), .A(n7996), .Z(n7993) );
  AND U8459 ( .A(b[19]), .B(a[16]), .Z(n7992) );
  XOR U8460 ( .A(n7997), .B(n7998), .Z(n7791) );
  AND U8461 ( .A(n7999), .B(n8000), .Z(n7997) );
  XNOR U8462 ( .A(n8001), .B(n7796), .Z(n7798) );
  XOR U8463 ( .A(n8002), .B(n8003), .Z(n7796) );
  ANDN U8464 ( .B(n8004), .A(n8005), .Z(n8002) );
  AND U8465 ( .A(b[18]), .B(a[17]), .Z(n8001) );
  XOR U8466 ( .A(n8006), .B(n7801), .Z(n7803) );
  XOR U8467 ( .A(n8007), .B(n8008), .Z(n7801) );
  ANDN U8468 ( .B(n8009), .A(n8010), .Z(n8007) );
  AND U8469 ( .A(b[16]), .B(a[19]), .Z(n8006) );
  XNOR U8470 ( .A(n8011), .B(n7806), .Z(n7808) );
  XOR U8471 ( .A(n8012), .B(n8013), .Z(n7806) );
  ANDN U8472 ( .B(n8014), .A(n8015), .Z(n8012) );
  AND U8473 ( .A(a[20]), .B(b[15]), .Z(n8011) );
  XNOR U8474 ( .A(n8016), .B(n7811), .Z(n7813) );
  XOR U8475 ( .A(n8017), .B(n8018), .Z(n7811) );
  ANDN U8476 ( .B(n8019), .A(n8020), .Z(n8017) );
  AND U8477 ( .A(b[14]), .B(a[21]), .Z(n8016) );
  XNOR U8478 ( .A(n8021), .B(n7816), .Z(n7818) );
  XOR U8479 ( .A(n8022), .B(n8023), .Z(n7816) );
  ANDN U8480 ( .B(n8024), .A(n8025), .Z(n8022) );
  AND U8481 ( .A(b[13]), .B(a[22]), .Z(n8021) );
  XOR U8482 ( .A(n8026), .B(n8027), .Z(n7820) );
  AND U8483 ( .A(n8028), .B(n8029), .Z(n8026) );
  XNOR U8484 ( .A(n8030), .B(n7825), .Z(n7827) );
  XOR U8485 ( .A(n8031), .B(n8032), .Z(n7825) );
  ANDN U8486 ( .B(n8033), .A(n8034), .Z(n8031) );
  AND U8487 ( .A(b[12]), .B(a[23]), .Z(n8030) );
  XOR U8488 ( .A(n8035), .B(n7830), .Z(n7832) );
  XOR U8489 ( .A(n8036), .B(n8037), .Z(n7830) );
  ANDN U8490 ( .B(n8038), .A(n8039), .Z(n8036) );
  AND U8491 ( .A(b[10]), .B(a[25]), .Z(n8035) );
  XNOR U8492 ( .A(n8040), .B(n7835), .Z(n7837) );
  XOR U8493 ( .A(n8041), .B(n8042), .Z(n7835) );
  ANDN U8494 ( .B(n8043), .A(n8044), .Z(n8041) );
  AND U8495 ( .A(b[9]), .B(a[26]), .Z(n8040) );
  XNOR U8496 ( .A(n8045), .B(n7840), .Z(n7842) );
  XOR U8497 ( .A(n8046), .B(n8047), .Z(n7840) );
  ANDN U8498 ( .B(n8048), .A(n8049), .Z(n8046) );
  AND U8499 ( .A(b[8]), .B(a[27]), .Z(n8045) );
  XNOR U8500 ( .A(n8050), .B(n7845), .Z(n7847) );
  XOR U8501 ( .A(n8051), .B(n8052), .Z(n7845) );
  ANDN U8502 ( .B(n8053), .A(n8054), .Z(n8051) );
  AND U8503 ( .A(b[7]), .B(a[28]), .Z(n8050) );
  XOR U8504 ( .A(n8055), .B(n8056), .Z(n7849) );
  AND U8505 ( .A(n8057), .B(n8058), .Z(n8055) );
  XNOR U8506 ( .A(n8059), .B(n7854), .Z(n7856) );
  XOR U8507 ( .A(n8060), .B(n8061), .Z(n7854) );
  ANDN U8508 ( .B(n8062), .A(n8063), .Z(n8060) );
  AND U8509 ( .A(b[6]), .B(a[29]), .Z(n8059) );
  XOR U8510 ( .A(n8064), .B(n7859), .Z(n7861) );
  XOR U8511 ( .A(n8065), .B(n8066), .Z(n7859) );
  ANDN U8512 ( .B(n8067), .A(n8068), .Z(n8065) );
  AND U8513 ( .A(b[4]), .B(a[31]), .Z(n8064) );
  XNOR U8514 ( .A(n8069), .B(n8070), .Z(n7873) );
  NANDN U8515 ( .A(n8071), .B(n8072), .Z(n8070) );
  XNOR U8516 ( .A(n8073), .B(n7864), .Z(n7866) );
  XNOR U8517 ( .A(n8074), .B(n8075), .Z(n7864) );
  AND U8518 ( .A(n8076), .B(n8077), .Z(n8074) );
  AND U8519 ( .A(b[3]), .B(a[32]), .Z(n8073) );
  NAND U8520 ( .A(a[35]), .B(b[0]), .Z(n7671) );
  XNOR U8521 ( .A(n7879), .B(n7880), .Z(c[34]) );
  XNOR U8522 ( .A(n8071), .B(n8072), .Z(n7880) );
  XOR U8523 ( .A(n8069), .B(n8078), .Z(n8072) );
  NAND U8524 ( .A(b[1]), .B(a[33]), .Z(n8078) );
  XOR U8525 ( .A(n8077), .B(n8079), .Z(n8071) );
  XOR U8526 ( .A(n8069), .B(n8076), .Z(n8079) );
  XNOR U8527 ( .A(n8080), .B(n8075), .Z(n8076) );
  AND U8528 ( .A(b[2]), .B(a[32]), .Z(n8080) );
  NANDN U8529 ( .A(n8081), .B(n8082), .Z(n8069) );
  XOR U8530 ( .A(n8075), .B(n8067), .Z(n8083) );
  XNOR U8531 ( .A(n8058), .B(n8057), .Z(n8084) );
  XOR U8532 ( .A(n8085), .B(n8056), .Z(n8057) );
  AND U8533 ( .A(b[4]), .B(a[30]), .Z(n8085) );
  XNOR U8534 ( .A(n8056), .B(n8062), .Z(n8086) );
  XNOR U8535 ( .A(n8061), .B(n8053), .Z(n8087) );
  XNOR U8536 ( .A(n8052), .B(n8048), .Z(n8088) );
  XNOR U8537 ( .A(n8047), .B(n8043), .Z(n8089) );
  XNOR U8538 ( .A(n8042), .B(n8038), .Z(n8090) );
  XNOR U8539 ( .A(n8029), .B(n8028), .Z(n8091) );
  XOR U8540 ( .A(n8092), .B(n8027), .Z(n8028) );
  AND U8541 ( .A(b[10]), .B(a[24]), .Z(n8092) );
  XNOR U8542 ( .A(n8027), .B(n8033), .Z(n8093) );
  XNOR U8543 ( .A(n8032), .B(n8024), .Z(n8094) );
  XNOR U8544 ( .A(n8023), .B(n8019), .Z(n8095) );
  XNOR U8545 ( .A(n8018), .B(n8014), .Z(n8096) );
  XNOR U8546 ( .A(n8013), .B(n8009), .Z(n8097) );
  XNOR U8547 ( .A(n8000), .B(n7999), .Z(n8098) );
  XOR U8548 ( .A(n8099), .B(n7998), .Z(n7999) );
  AND U8549 ( .A(b[16]), .B(a[18]), .Z(n8099) );
  XNOR U8550 ( .A(n7998), .B(n8004), .Z(n8100) );
  XNOR U8551 ( .A(n8003), .B(n7995), .Z(n8101) );
  XNOR U8552 ( .A(n7994), .B(n7990), .Z(n8102) );
  XNOR U8553 ( .A(n7989), .B(n7985), .Z(n8103) );
  XNOR U8554 ( .A(n7984), .B(n7980), .Z(n8104) );
  XNOR U8555 ( .A(n7971), .B(n7970), .Z(n8105) );
  XOR U8556 ( .A(n8106), .B(n7969), .Z(n7970) );
  AND U8557 ( .A(b[22]), .B(a[12]), .Z(n8106) );
  XNOR U8558 ( .A(n7969), .B(n7975), .Z(n8107) );
  XNOR U8559 ( .A(n7974), .B(n7966), .Z(n8108) );
  XNOR U8560 ( .A(n7965), .B(n7961), .Z(n8109) );
  XNOR U8561 ( .A(n7960), .B(n7956), .Z(n8110) );
  XNOR U8562 ( .A(n7955), .B(n7951), .Z(n8111) );
  XNOR U8563 ( .A(n7942), .B(n7941), .Z(n8112) );
  XOR U8564 ( .A(n8113), .B(n7940), .Z(n7941) );
  AND U8565 ( .A(a[6]), .B(b[28]), .Z(n8113) );
  XNOR U8566 ( .A(n7940), .B(n7946), .Z(n8114) );
  XNOR U8567 ( .A(n7945), .B(n7937), .Z(n8115) );
  XNOR U8568 ( .A(n7936), .B(n7932), .Z(n8116) );
  XNOR U8569 ( .A(n7931), .B(n7927), .Z(n8117) );
  XNOR U8570 ( .A(n7926), .B(n7922), .Z(n8118) );
  XOR U8571 ( .A(n8119), .B(n7921), .Z(n7922) );
  AND U8572 ( .A(a[0]), .B(b[34]), .Z(n8119) );
  XNOR U8573 ( .A(n8120), .B(n7921), .Z(n7923) );
  XNOR U8574 ( .A(n8121), .B(n8122), .Z(n7921) );
  ANDN U8575 ( .B(n8123), .A(n8124), .Z(n8121) );
  AND U8576 ( .A(a[1]), .B(b[33]), .Z(n8120) );
  XNOR U8577 ( .A(n8125), .B(n7926), .Z(n7928) );
  XOR U8578 ( .A(n8126), .B(n8127), .Z(n7926) );
  ANDN U8579 ( .B(n8128), .A(n8129), .Z(n8126) );
  AND U8580 ( .A(a[2]), .B(b[32]), .Z(n8125) );
  XNOR U8581 ( .A(n8130), .B(n7931), .Z(n7933) );
  XOR U8582 ( .A(n8131), .B(n8132), .Z(n7931) );
  ANDN U8583 ( .B(n8133), .A(n8134), .Z(n8131) );
  AND U8584 ( .A(a[3]), .B(b[31]), .Z(n8130) );
  XNOR U8585 ( .A(n8135), .B(n7936), .Z(n7938) );
  XOR U8586 ( .A(n8136), .B(n8137), .Z(n7936) );
  ANDN U8587 ( .B(n8138), .A(n8139), .Z(n8136) );
  AND U8588 ( .A(a[4]), .B(b[30]), .Z(n8135) );
  XOR U8589 ( .A(n8140), .B(n8141), .Z(n7940) );
  AND U8590 ( .A(n8142), .B(n8143), .Z(n8140) );
  XNOR U8591 ( .A(n8144), .B(n7945), .Z(n7947) );
  XOR U8592 ( .A(n8145), .B(n8146), .Z(n7945) );
  ANDN U8593 ( .B(n8147), .A(n8148), .Z(n8145) );
  AND U8594 ( .A(a[5]), .B(b[29]), .Z(n8144) );
  XOR U8595 ( .A(n8149), .B(n7950), .Z(n7952) );
  XOR U8596 ( .A(n8150), .B(n8151), .Z(n7950) );
  ANDN U8597 ( .B(n8152), .A(n8153), .Z(n8150) );
  AND U8598 ( .A(a[7]), .B(b[27]), .Z(n8149) );
  XNOR U8599 ( .A(n8154), .B(n7955), .Z(n7957) );
  XOR U8600 ( .A(n8155), .B(n8156), .Z(n7955) );
  ANDN U8601 ( .B(n8157), .A(n8158), .Z(n8155) );
  AND U8602 ( .A(a[8]), .B(b[26]), .Z(n8154) );
  XNOR U8603 ( .A(n8159), .B(n7960), .Z(n7962) );
  XOR U8604 ( .A(n8160), .B(n8161), .Z(n7960) );
  ANDN U8605 ( .B(n8162), .A(n8163), .Z(n8160) );
  AND U8606 ( .A(a[9]), .B(b[25]), .Z(n8159) );
  XNOR U8607 ( .A(n8164), .B(n7965), .Z(n7967) );
  XOR U8608 ( .A(n8165), .B(n8166), .Z(n7965) );
  ANDN U8609 ( .B(n8167), .A(n8168), .Z(n8165) );
  AND U8610 ( .A(b[24]), .B(a[10]), .Z(n8164) );
  XOR U8611 ( .A(n8169), .B(n8170), .Z(n7969) );
  AND U8612 ( .A(n8171), .B(n8172), .Z(n8169) );
  XNOR U8613 ( .A(n8173), .B(n7974), .Z(n7976) );
  XOR U8614 ( .A(n8174), .B(n8175), .Z(n7974) );
  ANDN U8615 ( .B(n8176), .A(n8177), .Z(n8174) );
  AND U8616 ( .A(b[23]), .B(a[11]), .Z(n8173) );
  XOR U8617 ( .A(n8178), .B(n7979), .Z(n7981) );
  XOR U8618 ( .A(n8179), .B(n8180), .Z(n7979) );
  ANDN U8619 ( .B(n8181), .A(n8182), .Z(n8179) );
  AND U8620 ( .A(a[13]), .B(b[21]), .Z(n8178) );
  XNOR U8621 ( .A(n8183), .B(n7984), .Z(n7986) );
  XOR U8622 ( .A(n8184), .B(n8185), .Z(n7984) );
  ANDN U8623 ( .B(n8186), .A(n8187), .Z(n8184) );
  AND U8624 ( .A(b[20]), .B(a[14]), .Z(n8183) );
  XNOR U8625 ( .A(n8188), .B(n7989), .Z(n7991) );
  XOR U8626 ( .A(n8189), .B(n8190), .Z(n7989) );
  ANDN U8627 ( .B(n8191), .A(n8192), .Z(n8189) );
  AND U8628 ( .A(b[19]), .B(a[15]), .Z(n8188) );
  XNOR U8629 ( .A(n8193), .B(n7994), .Z(n7996) );
  XOR U8630 ( .A(n8194), .B(n8195), .Z(n7994) );
  ANDN U8631 ( .B(n8196), .A(n8197), .Z(n8194) );
  AND U8632 ( .A(b[18]), .B(a[16]), .Z(n8193) );
  XOR U8633 ( .A(n8198), .B(n8199), .Z(n7998) );
  AND U8634 ( .A(n8200), .B(n8201), .Z(n8198) );
  XNOR U8635 ( .A(n8202), .B(n8003), .Z(n8005) );
  XOR U8636 ( .A(n8203), .B(n8204), .Z(n8003) );
  ANDN U8637 ( .B(n8205), .A(n8206), .Z(n8203) );
  AND U8638 ( .A(b[17]), .B(a[17]), .Z(n8202) );
  XOR U8639 ( .A(n8207), .B(n8008), .Z(n8010) );
  XOR U8640 ( .A(n8208), .B(n8209), .Z(n8008) );
  ANDN U8641 ( .B(n8210), .A(n8211), .Z(n8208) );
  AND U8642 ( .A(a[19]), .B(b[15]), .Z(n8207) );
  XNOR U8643 ( .A(n8212), .B(n8013), .Z(n8015) );
  XOR U8644 ( .A(n8213), .B(n8214), .Z(n8013) );
  ANDN U8645 ( .B(n8215), .A(n8216), .Z(n8213) );
  AND U8646 ( .A(b[14]), .B(a[20]), .Z(n8212) );
  XNOR U8647 ( .A(n8217), .B(n8018), .Z(n8020) );
  XOR U8648 ( .A(n8218), .B(n8219), .Z(n8018) );
  ANDN U8649 ( .B(n8220), .A(n8221), .Z(n8218) );
  AND U8650 ( .A(b[13]), .B(a[21]), .Z(n8217) );
  XNOR U8651 ( .A(n8222), .B(n8023), .Z(n8025) );
  XOR U8652 ( .A(n8223), .B(n8224), .Z(n8023) );
  ANDN U8653 ( .B(n8225), .A(n8226), .Z(n8223) );
  AND U8654 ( .A(b[12]), .B(a[22]), .Z(n8222) );
  XOR U8655 ( .A(n8227), .B(n8228), .Z(n8027) );
  AND U8656 ( .A(n8229), .B(n8230), .Z(n8227) );
  XNOR U8657 ( .A(n8231), .B(n8032), .Z(n8034) );
  XOR U8658 ( .A(n8232), .B(n8233), .Z(n8032) );
  ANDN U8659 ( .B(n8234), .A(n8235), .Z(n8232) );
  AND U8660 ( .A(b[11]), .B(a[23]), .Z(n8231) );
  XOR U8661 ( .A(n8236), .B(n8037), .Z(n8039) );
  XOR U8662 ( .A(n8237), .B(n8238), .Z(n8037) );
  ANDN U8663 ( .B(n8239), .A(n8240), .Z(n8237) );
  AND U8664 ( .A(b[9]), .B(a[25]), .Z(n8236) );
  XNOR U8665 ( .A(n8241), .B(n8042), .Z(n8044) );
  XOR U8666 ( .A(n8242), .B(n8243), .Z(n8042) );
  ANDN U8667 ( .B(n8244), .A(n8245), .Z(n8242) );
  AND U8668 ( .A(b[8]), .B(a[26]), .Z(n8241) );
  XNOR U8669 ( .A(n8246), .B(n8047), .Z(n8049) );
  XOR U8670 ( .A(n8247), .B(n8248), .Z(n8047) );
  ANDN U8671 ( .B(n8249), .A(n8250), .Z(n8247) );
  AND U8672 ( .A(b[7]), .B(a[27]), .Z(n8246) );
  XNOR U8673 ( .A(n8251), .B(n8052), .Z(n8054) );
  XOR U8674 ( .A(n8252), .B(n8253), .Z(n8052) );
  ANDN U8675 ( .B(n8254), .A(n8255), .Z(n8252) );
  AND U8676 ( .A(b[6]), .B(a[28]), .Z(n8251) );
  XOR U8677 ( .A(n8256), .B(n8257), .Z(n8056) );
  AND U8678 ( .A(n8258), .B(n8259), .Z(n8256) );
  XNOR U8679 ( .A(n8260), .B(n8061), .Z(n8063) );
  XOR U8680 ( .A(n8261), .B(n8262), .Z(n8061) );
  ANDN U8681 ( .B(n8263), .A(n8264), .Z(n8261) );
  AND U8682 ( .A(b[5]), .B(a[29]), .Z(n8260) );
  XNOR U8683 ( .A(n8265), .B(n8266), .Z(n8075) );
  NANDN U8684 ( .A(n8267), .B(n8268), .Z(n8266) );
  XOR U8685 ( .A(n8269), .B(n8066), .Z(n8068) );
  XOR U8686 ( .A(n8270), .B(n8271), .Z(n8066) );
  ANDN U8687 ( .B(n8272), .A(n8273), .Z(n8270) );
  AND U8688 ( .A(b[3]), .B(a[31]), .Z(n8269) );
  NAND U8689 ( .A(a[34]), .B(b[0]), .Z(n7879) );
  XNOR U8690 ( .A(n8081), .B(n8082), .Z(c[33]) );
  XNOR U8691 ( .A(n8267), .B(n8268), .Z(n8082) );
  XOR U8692 ( .A(n8265), .B(n8274), .Z(n8268) );
  NAND U8693 ( .A(b[1]), .B(a[32]), .Z(n8274) );
  XNOR U8694 ( .A(n8273), .B(n8275), .Z(n8267) );
  XOR U8695 ( .A(n8265), .B(n8272), .Z(n8275) );
  XNOR U8696 ( .A(n8276), .B(n8271), .Z(n8272) );
  AND U8697 ( .A(b[2]), .B(a[31]), .Z(n8276) );
  NANDN U8698 ( .A(n8277), .B(n8278), .Z(n8265) );
  XNOR U8699 ( .A(n8271), .B(n8279), .Z(n8273) );
  XNOR U8700 ( .A(n8259), .B(n8258), .Z(n8279) );
  XOR U8701 ( .A(n8280), .B(n8257), .Z(n8258) );
  AND U8702 ( .A(b[3]), .B(a[30]), .Z(n8280) );
  XNOR U8703 ( .A(n8257), .B(n8263), .Z(n8281) );
  XNOR U8704 ( .A(n8262), .B(n8254), .Z(n8282) );
  XNOR U8705 ( .A(n8253), .B(n8249), .Z(n8283) );
  XNOR U8706 ( .A(n8248), .B(n8244), .Z(n8284) );
  XNOR U8707 ( .A(n8243), .B(n8239), .Z(n8285) );
  XNOR U8708 ( .A(n8230), .B(n8229), .Z(n8286) );
  XOR U8709 ( .A(n8287), .B(n8228), .Z(n8229) );
  AND U8710 ( .A(b[9]), .B(a[24]), .Z(n8287) );
  XNOR U8711 ( .A(n8228), .B(n8234), .Z(n8288) );
  XNOR U8712 ( .A(n8233), .B(n8225), .Z(n8289) );
  XNOR U8713 ( .A(n8224), .B(n8220), .Z(n8290) );
  XNOR U8714 ( .A(n8219), .B(n8215), .Z(n8291) );
  XNOR U8715 ( .A(n8214), .B(n8210), .Z(n8292) );
  XNOR U8716 ( .A(n8201), .B(n8200), .Z(n8293) );
  XOR U8717 ( .A(n8294), .B(n8199), .Z(n8200) );
  AND U8718 ( .A(b[15]), .B(a[18]), .Z(n8294) );
  XNOR U8719 ( .A(n8199), .B(n8205), .Z(n8295) );
  XNOR U8720 ( .A(n8204), .B(n8196), .Z(n8296) );
  XNOR U8721 ( .A(n8195), .B(n8191), .Z(n8297) );
  XNOR U8722 ( .A(n8190), .B(n8186), .Z(n8298) );
  XNOR U8723 ( .A(n8185), .B(n8181), .Z(n8299) );
  XNOR U8724 ( .A(n8172), .B(n8171), .Z(n8300) );
  XOR U8725 ( .A(n8301), .B(n8170), .Z(n8171) );
  AND U8726 ( .A(b[21]), .B(a[12]), .Z(n8301) );
  XNOR U8727 ( .A(n8170), .B(n8176), .Z(n8302) );
  XNOR U8728 ( .A(n8175), .B(n8167), .Z(n8303) );
  XNOR U8729 ( .A(n8166), .B(n8162), .Z(n8304) );
  XNOR U8730 ( .A(n8161), .B(n8157), .Z(n8305) );
  XNOR U8731 ( .A(n8156), .B(n8152), .Z(n8306) );
  XNOR U8732 ( .A(n8143), .B(n8142), .Z(n8307) );
  XOR U8733 ( .A(n8308), .B(n8141), .Z(n8142) );
  AND U8734 ( .A(a[6]), .B(b[27]), .Z(n8308) );
  XNOR U8735 ( .A(n8141), .B(n8147), .Z(n8309) );
  XNOR U8736 ( .A(n8146), .B(n8138), .Z(n8310) );
  XNOR U8737 ( .A(n8137), .B(n8133), .Z(n8311) );
  XNOR U8738 ( .A(n8132), .B(n8128), .Z(n8312) );
  XNOR U8739 ( .A(n8127), .B(n8123), .Z(n8313) );
  XNOR U8740 ( .A(n8314), .B(n8122), .Z(n8123) );
  AND U8741 ( .A(a[0]), .B(b[33]), .Z(n8314) );
  XOR U8742 ( .A(n8315), .B(n8122), .Z(n8124) );
  XNOR U8743 ( .A(n8316), .B(n8317), .Z(n8122) );
  ANDN U8744 ( .B(n8318), .A(n8319), .Z(n8316) );
  AND U8745 ( .A(a[1]), .B(b[32]), .Z(n8315) );
  XNOR U8746 ( .A(n8320), .B(n8127), .Z(n8129) );
  XOR U8747 ( .A(n8321), .B(n8322), .Z(n8127) );
  ANDN U8748 ( .B(n8323), .A(n8324), .Z(n8321) );
  AND U8749 ( .A(a[2]), .B(b[31]), .Z(n8320) );
  XNOR U8750 ( .A(n8325), .B(n8132), .Z(n8134) );
  XOR U8751 ( .A(n8326), .B(n8327), .Z(n8132) );
  ANDN U8752 ( .B(n8328), .A(n8329), .Z(n8326) );
  AND U8753 ( .A(a[3]), .B(b[30]), .Z(n8325) );
  XNOR U8754 ( .A(n8330), .B(n8137), .Z(n8139) );
  XOR U8755 ( .A(n8331), .B(n8332), .Z(n8137) );
  ANDN U8756 ( .B(n8333), .A(n8334), .Z(n8331) );
  AND U8757 ( .A(a[4]), .B(b[29]), .Z(n8330) );
  XOR U8758 ( .A(n8335), .B(n8336), .Z(n8141) );
  AND U8759 ( .A(n8337), .B(n8338), .Z(n8335) );
  XNOR U8760 ( .A(n8339), .B(n8146), .Z(n8148) );
  XOR U8761 ( .A(n8340), .B(n8341), .Z(n8146) );
  ANDN U8762 ( .B(n8342), .A(n8343), .Z(n8340) );
  AND U8763 ( .A(a[5]), .B(b[28]), .Z(n8339) );
  XOR U8764 ( .A(n8344), .B(n8151), .Z(n8153) );
  XOR U8765 ( .A(n8345), .B(n8346), .Z(n8151) );
  ANDN U8766 ( .B(n8347), .A(n8348), .Z(n8345) );
  AND U8767 ( .A(a[7]), .B(b[26]), .Z(n8344) );
  XNOR U8768 ( .A(n8349), .B(n8156), .Z(n8158) );
  XOR U8769 ( .A(n8350), .B(n8351), .Z(n8156) );
  ANDN U8770 ( .B(n8352), .A(n8353), .Z(n8350) );
  AND U8771 ( .A(a[8]), .B(b[25]), .Z(n8349) );
  XNOR U8772 ( .A(n8354), .B(n8161), .Z(n8163) );
  XOR U8773 ( .A(n8355), .B(n8356), .Z(n8161) );
  ANDN U8774 ( .B(n8357), .A(n8358), .Z(n8355) );
  AND U8775 ( .A(a[9]), .B(b[24]), .Z(n8354) );
  XNOR U8776 ( .A(n8359), .B(n8166), .Z(n8168) );
  XOR U8777 ( .A(n8360), .B(n8361), .Z(n8166) );
  ANDN U8778 ( .B(n8362), .A(n8363), .Z(n8360) );
  AND U8779 ( .A(b[23]), .B(a[10]), .Z(n8359) );
  XOR U8780 ( .A(n8364), .B(n8365), .Z(n8170) );
  AND U8781 ( .A(n8366), .B(n8367), .Z(n8364) );
  XNOR U8782 ( .A(n8368), .B(n8175), .Z(n8177) );
  XOR U8783 ( .A(n8369), .B(n8370), .Z(n8175) );
  ANDN U8784 ( .B(n8371), .A(n8372), .Z(n8369) );
  AND U8785 ( .A(b[22]), .B(a[11]), .Z(n8368) );
  XOR U8786 ( .A(n8373), .B(n8180), .Z(n8182) );
  XOR U8787 ( .A(n8374), .B(n8375), .Z(n8180) );
  ANDN U8788 ( .B(n8376), .A(n8377), .Z(n8374) );
  AND U8789 ( .A(b[20]), .B(a[13]), .Z(n8373) );
  XNOR U8790 ( .A(n8378), .B(n8185), .Z(n8187) );
  XOR U8791 ( .A(n8379), .B(n8380), .Z(n8185) );
  ANDN U8792 ( .B(n8381), .A(n8382), .Z(n8379) );
  AND U8793 ( .A(b[19]), .B(a[14]), .Z(n8378) );
  XNOR U8794 ( .A(n8383), .B(n8190), .Z(n8192) );
  XOR U8795 ( .A(n8384), .B(n8385), .Z(n8190) );
  ANDN U8796 ( .B(n8386), .A(n8387), .Z(n8384) );
  AND U8797 ( .A(b[18]), .B(a[15]), .Z(n8383) );
  XNOR U8798 ( .A(n8388), .B(n8195), .Z(n8197) );
  XOR U8799 ( .A(n8389), .B(n8390), .Z(n8195) );
  ANDN U8800 ( .B(n8391), .A(n8392), .Z(n8389) );
  AND U8801 ( .A(b[17]), .B(a[16]), .Z(n8388) );
  XOR U8802 ( .A(n8393), .B(n8394), .Z(n8199) );
  AND U8803 ( .A(n8395), .B(n8396), .Z(n8393) );
  XNOR U8804 ( .A(n8397), .B(n8204), .Z(n8206) );
  XOR U8805 ( .A(n8398), .B(n8399), .Z(n8204) );
  ANDN U8806 ( .B(n8400), .A(n8401), .Z(n8398) );
  AND U8807 ( .A(b[16]), .B(a[17]), .Z(n8397) );
  XOR U8808 ( .A(n8402), .B(n8209), .Z(n8211) );
  XOR U8809 ( .A(n8403), .B(n8404), .Z(n8209) );
  ANDN U8810 ( .B(n8405), .A(n8406), .Z(n8403) );
  AND U8811 ( .A(b[14]), .B(a[19]), .Z(n8402) );
  XNOR U8812 ( .A(n8407), .B(n8214), .Z(n8216) );
  XOR U8813 ( .A(n8408), .B(n8409), .Z(n8214) );
  ANDN U8814 ( .B(n8410), .A(n8411), .Z(n8408) );
  AND U8815 ( .A(b[13]), .B(a[20]), .Z(n8407) );
  XNOR U8816 ( .A(n8412), .B(n8219), .Z(n8221) );
  XOR U8817 ( .A(n8413), .B(n8414), .Z(n8219) );
  ANDN U8818 ( .B(n8415), .A(n8416), .Z(n8413) );
  AND U8819 ( .A(b[12]), .B(a[21]), .Z(n8412) );
  XNOR U8820 ( .A(n8417), .B(n8224), .Z(n8226) );
  XOR U8821 ( .A(n8418), .B(n8419), .Z(n8224) );
  ANDN U8822 ( .B(n8420), .A(n8421), .Z(n8418) );
  AND U8823 ( .A(b[11]), .B(a[22]), .Z(n8417) );
  XOR U8824 ( .A(n8422), .B(n8423), .Z(n8228) );
  AND U8825 ( .A(n8424), .B(n8425), .Z(n8422) );
  XNOR U8826 ( .A(n8426), .B(n8233), .Z(n8235) );
  XOR U8827 ( .A(n8427), .B(n8428), .Z(n8233) );
  ANDN U8828 ( .B(n8429), .A(n8430), .Z(n8427) );
  AND U8829 ( .A(b[10]), .B(a[23]), .Z(n8426) );
  XOR U8830 ( .A(n8431), .B(n8238), .Z(n8240) );
  XOR U8831 ( .A(n8432), .B(n8433), .Z(n8238) );
  ANDN U8832 ( .B(n8434), .A(n8435), .Z(n8432) );
  AND U8833 ( .A(b[8]), .B(a[25]), .Z(n8431) );
  XNOR U8834 ( .A(n8436), .B(n8243), .Z(n8245) );
  XOR U8835 ( .A(n8437), .B(n8438), .Z(n8243) );
  ANDN U8836 ( .B(n8439), .A(n8440), .Z(n8437) );
  AND U8837 ( .A(b[7]), .B(a[26]), .Z(n8436) );
  XNOR U8838 ( .A(n8441), .B(n8248), .Z(n8250) );
  XOR U8839 ( .A(n8442), .B(n8443), .Z(n8248) );
  ANDN U8840 ( .B(n8444), .A(n8445), .Z(n8442) );
  AND U8841 ( .A(b[6]), .B(a[27]), .Z(n8441) );
  XNOR U8842 ( .A(n8446), .B(n8253), .Z(n8255) );
  XOR U8843 ( .A(n8447), .B(n8448), .Z(n8253) );
  ANDN U8844 ( .B(n8449), .A(n8450), .Z(n8447) );
  AND U8845 ( .A(b[5]), .B(a[28]), .Z(n8446) );
  XOR U8846 ( .A(n8451), .B(n8452), .Z(n8257) );
  ANDN U8847 ( .B(n8453), .A(n8454), .Z(n8451) );
  XNOR U8848 ( .A(n8455), .B(n8262), .Z(n8264) );
  XOR U8849 ( .A(n8456), .B(n8457), .Z(n8262) );
  ANDN U8850 ( .B(n8458), .A(n8459), .Z(n8456) );
  AND U8851 ( .A(b[4]), .B(a[29]), .Z(n8455) );
  XNOR U8852 ( .A(n8460), .B(n8461), .Z(n8271) );
  NAND U8853 ( .A(n8462), .B(n8463), .Z(n8461) );
  NAND U8854 ( .A(a[33]), .B(b[0]), .Z(n8081) );
  XNOR U8855 ( .A(n8277), .B(n8278), .Z(c[32]) );
  XOR U8856 ( .A(n8462), .B(n8463), .Z(n8278) );
  XOR U8857 ( .A(n8460), .B(n8464), .Z(n8463) );
  NAND U8858 ( .A(b[1]), .B(a[31]), .Z(n8464) );
  XOR U8859 ( .A(n8460), .B(n8453), .Z(n8465) );
  XNOR U8860 ( .A(n8452), .B(n8458), .Z(n8466) );
  XNOR U8861 ( .A(n8457), .B(n8449), .Z(n8467) );
  XNOR U8862 ( .A(n8448), .B(n8444), .Z(n8468) );
  XNOR U8863 ( .A(n8443), .B(n8439), .Z(n8469) );
  XNOR U8864 ( .A(n8438), .B(n8434), .Z(n8470) );
  XNOR U8865 ( .A(n8425), .B(n8424), .Z(n8471) );
  XOR U8866 ( .A(n8472), .B(n8423), .Z(n8424) );
  AND U8867 ( .A(b[8]), .B(a[24]), .Z(n8472) );
  XNOR U8868 ( .A(n8423), .B(n8429), .Z(n8473) );
  XNOR U8869 ( .A(n8428), .B(n8420), .Z(n8474) );
  XNOR U8870 ( .A(n8419), .B(n8415), .Z(n8475) );
  XNOR U8871 ( .A(n8414), .B(n8410), .Z(n8476) );
  XNOR U8872 ( .A(n8409), .B(n8405), .Z(n8477) );
  XNOR U8873 ( .A(n8396), .B(n8395), .Z(n8478) );
  XOR U8874 ( .A(n8479), .B(n8394), .Z(n8395) );
  AND U8875 ( .A(b[14]), .B(a[18]), .Z(n8479) );
  XNOR U8876 ( .A(n8394), .B(n8400), .Z(n8480) );
  XNOR U8877 ( .A(n8399), .B(n8391), .Z(n8481) );
  XNOR U8878 ( .A(n8390), .B(n8386), .Z(n8482) );
  XNOR U8879 ( .A(n8385), .B(n8381), .Z(n8483) );
  XNOR U8880 ( .A(n8380), .B(n8376), .Z(n8484) );
  XNOR U8881 ( .A(n8367), .B(n8366), .Z(n8485) );
  XOR U8882 ( .A(n8486), .B(n8365), .Z(n8366) );
  AND U8883 ( .A(b[20]), .B(a[12]), .Z(n8486) );
  XNOR U8884 ( .A(n8365), .B(n8371), .Z(n8487) );
  XNOR U8885 ( .A(n8370), .B(n8362), .Z(n8488) );
  XNOR U8886 ( .A(n8361), .B(n8357), .Z(n8489) );
  XNOR U8887 ( .A(n8356), .B(n8352), .Z(n8490) );
  XNOR U8888 ( .A(n8351), .B(n8347), .Z(n8491) );
  XNOR U8889 ( .A(n8338), .B(n8337), .Z(n8492) );
  XOR U8890 ( .A(n8493), .B(n8336), .Z(n8337) );
  AND U8891 ( .A(a[6]), .B(b[26]), .Z(n8493) );
  XNOR U8892 ( .A(n8336), .B(n8342), .Z(n8494) );
  XNOR U8893 ( .A(n8341), .B(n8333), .Z(n8495) );
  XNOR U8894 ( .A(n8332), .B(n8328), .Z(n8496) );
  XNOR U8895 ( .A(n8327), .B(n8323), .Z(n8497) );
  XNOR U8896 ( .A(n8322), .B(n8318), .Z(n8498) );
  XOR U8897 ( .A(n8499), .B(n8317), .Z(n8318) );
  AND U8898 ( .A(a[0]), .B(b[32]), .Z(n8499) );
  XNOR U8899 ( .A(n8500), .B(n8317), .Z(n8319) );
  XNOR U8900 ( .A(n8501), .B(n8502), .Z(n8317) );
  ANDN U8901 ( .B(n8503), .A(n8504), .Z(n8501) );
  AND U8902 ( .A(a[1]), .B(b[31]), .Z(n8500) );
  XNOR U8903 ( .A(n8505), .B(n8322), .Z(n8324) );
  XOR U8904 ( .A(n8506), .B(n8507), .Z(n8322) );
  ANDN U8905 ( .B(n8508), .A(n8509), .Z(n8506) );
  AND U8906 ( .A(a[2]), .B(b[30]), .Z(n8505) );
  XNOR U8907 ( .A(n8510), .B(n8327), .Z(n8329) );
  XOR U8908 ( .A(n8511), .B(n8512), .Z(n8327) );
  ANDN U8909 ( .B(n8513), .A(n8514), .Z(n8511) );
  AND U8910 ( .A(a[3]), .B(b[29]), .Z(n8510) );
  XNOR U8911 ( .A(n8515), .B(n8332), .Z(n8334) );
  XOR U8912 ( .A(n8516), .B(n8517), .Z(n8332) );
  ANDN U8913 ( .B(n8518), .A(n8519), .Z(n8516) );
  AND U8914 ( .A(a[4]), .B(b[28]), .Z(n8515) );
  XOR U8915 ( .A(n8520), .B(n8521), .Z(n8336) );
  AND U8916 ( .A(n8522), .B(n8523), .Z(n8520) );
  XNOR U8917 ( .A(n8524), .B(n8341), .Z(n8343) );
  XOR U8918 ( .A(n8525), .B(n8526), .Z(n8341) );
  ANDN U8919 ( .B(n8527), .A(n8528), .Z(n8525) );
  AND U8920 ( .A(a[5]), .B(b[27]), .Z(n8524) );
  XOR U8921 ( .A(n8529), .B(n8346), .Z(n8348) );
  XOR U8922 ( .A(n8530), .B(n8531), .Z(n8346) );
  ANDN U8923 ( .B(n8532), .A(n8533), .Z(n8530) );
  AND U8924 ( .A(a[7]), .B(b[25]), .Z(n8529) );
  XNOR U8925 ( .A(n8534), .B(n8351), .Z(n8353) );
  XOR U8926 ( .A(n8535), .B(n8536), .Z(n8351) );
  ANDN U8927 ( .B(n8537), .A(n8538), .Z(n8535) );
  AND U8928 ( .A(a[8]), .B(b[24]), .Z(n8534) );
  XNOR U8929 ( .A(n8539), .B(n8356), .Z(n8358) );
  XOR U8930 ( .A(n8540), .B(n8541), .Z(n8356) );
  ANDN U8931 ( .B(n8542), .A(n8543), .Z(n8540) );
  AND U8932 ( .A(a[9]), .B(b[23]), .Z(n8539) );
  XNOR U8933 ( .A(n8544), .B(n8361), .Z(n8363) );
  XOR U8934 ( .A(n8545), .B(n8546), .Z(n8361) );
  ANDN U8935 ( .B(n8547), .A(n8548), .Z(n8545) );
  AND U8936 ( .A(b[22]), .B(a[10]), .Z(n8544) );
  XOR U8937 ( .A(n8549), .B(n8550), .Z(n8365) );
  AND U8938 ( .A(n8551), .B(n8552), .Z(n8549) );
  XNOR U8939 ( .A(n8553), .B(n8370), .Z(n8372) );
  XOR U8940 ( .A(n8554), .B(n8555), .Z(n8370) );
  ANDN U8941 ( .B(n8556), .A(n8557), .Z(n8554) );
  AND U8942 ( .A(a[11]), .B(b[21]), .Z(n8553) );
  XOR U8943 ( .A(n8558), .B(n8375), .Z(n8377) );
  XOR U8944 ( .A(n8559), .B(n8560), .Z(n8375) );
  ANDN U8945 ( .B(n8561), .A(n8562), .Z(n8559) );
  AND U8946 ( .A(b[19]), .B(a[13]), .Z(n8558) );
  XNOR U8947 ( .A(n8563), .B(n8380), .Z(n8382) );
  XOR U8948 ( .A(n8564), .B(n8565), .Z(n8380) );
  ANDN U8949 ( .B(n8566), .A(n8567), .Z(n8564) );
  AND U8950 ( .A(b[18]), .B(a[14]), .Z(n8563) );
  XNOR U8951 ( .A(n8568), .B(n8385), .Z(n8387) );
  XOR U8952 ( .A(n8569), .B(n8570), .Z(n8385) );
  ANDN U8953 ( .B(n8571), .A(n8572), .Z(n8569) );
  AND U8954 ( .A(b[17]), .B(a[15]), .Z(n8568) );
  XNOR U8955 ( .A(n8573), .B(n8390), .Z(n8392) );
  XOR U8956 ( .A(n8574), .B(n8575), .Z(n8390) );
  ANDN U8957 ( .B(n8576), .A(n8577), .Z(n8574) );
  AND U8958 ( .A(b[16]), .B(a[16]), .Z(n8573) );
  XOR U8959 ( .A(n8578), .B(n8579), .Z(n8394) );
  AND U8960 ( .A(n8580), .B(n8581), .Z(n8578) );
  XNOR U8961 ( .A(n8582), .B(n8399), .Z(n8401) );
  XOR U8962 ( .A(n8583), .B(n8584), .Z(n8399) );
  ANDN U8963 ( .B(n8585), .A(n8586), .Z(n8583) );
  AND U8964 ( .A(a[17]), .B(b[15]), .Z(n8582) );
  XOR U8965 ( .A(n8587), .B(n8404), .Z(n8406) );
  XOR U8966 ( .A(n8588), .B(n8589), .Z(n8404) );
  ANDN U8967 ( .B(n8590), .A(n8591), .Z(n8588) );
  AND U8968 ( .A(b[13]), .B(a[19]), .Z(n8587) );
  XNOR U8969 ( .A(n8592), .B(n8409), .Z(n8411) );
  XOR U8970 ( .A(n8593), .B(n8594), .Z(n8409) );
  ANDN U8971 ( .B(n8595), .A(n8596), .Z(n8593) );
  AND U8972 ( .A(b[12]), .B(a[20]), .Z(n8592) );
  XNOR U8973 ( .A(n8597), .B(n8414), .Z(n8416) );
  XOR U8974 ( .A(n8598), .B(n8599), .Z(n8414) );
  ANDN U8975 ( .B(n8600), .A(n8601), .Z(n8598) );
  AND U8976 ( .A(b[11]), .B(a[21]), .Z(n8597) );
  XNOR U8977 ( .A(n8602), .B(n8419), .Z(n8421) );
  XOR U8978 ( .A(n8603), .B(n8604), .Z(n8419) );
  ANDN U8979 ( .B(n8605), .A(n8606), .Z(n8603) );
  AND U8980 ( .A(b[10]), .B(a[22]), .Z(n8602) );
  XOR U8981 ( .A(n8607), .B(n8608), .Z(n8423) );
  AND U8982 ( .A(n8609), .B(n8610), .Z(n8607) );
  XNOR U8983 ( .A(n8611), .B(n8428), .Z(n8430) );
  XOR U8984 ( .A(n8612), .B(n8613), .Z(n8428) );
  ANDN U8985 ( .B(n8614), .A(n8615), .Z(n8612) );
  AND U8986 ( .A(b[9]), .B(a[23]), .Z(n8611) );
  XOR U8987 ( .A(n8616), .B(n8433), .Z(n8435) );
  XOR U8988 ( .A(n8617), .B(n8618), .Z(n8433) );
  ANDN U8989 ( .B(n8619), .A(n8620), .Z(n8617) );
  AND U8990 ( .A(b[7]), .B(a[25]), .Z(n8616) );
  XNOR U8991 ( .A(n8621), .B(n8438), .Z(n8440) );
  XOR U8992 ( .A(n8622), .B(n8623), .Z(n8438) );
  ANDN U8993 ( .B(n8624), .A(n8625), .Z(n8622) );
  AND U8994 ( .A(b[6]), .B(a[26]), .Z(n8621) );
  XNOR U8995 ( .A(n8626), .B(n8443), .Z(n8445) );
  XOR U8996 ( .A(n8627), .B(n8628), .Z(n8443) );
  ANDN U8997 ( .B(n8629), .A(n8630), .Z(n8627) );
  AND U8998 ( .A(b[5]), .B(a[27]), .Z(n8626) );
  XNOR U8999 ( .A(n8631), .B(n8448), .Z(n8450) );
  XOR U9000 ( .A(n8632), .B(n8633), .Z(n8448) );
  ANDN U9001 ( .B(n8634), .A(n8635), .Z(n8632) );
  AND U9002 ( .A(b[4]), .B(a[28]), .Z(n8631) );
  XNOR U9003 ( .A(n8636), .B(n8457), .Z(n8459) );
  XNOR U9004 ( .A(n8637), .B(n8638), .Z(n8457) );
  NOR U9005 ( .A(n8639), .B(n8640), .Z(n8637) );
  AND U9006 ( .A(b[3]), .B(a[29]), .Z(n8636) );
  NANDN U9007 ( .A(n8641), .B(n8642), .Z(n8460) );
  XNOR U9008 ( .A(n8643), .B(n8452), .Z(n8454) );
  XNOR U9009 ( .A(n8644), .B(n8645), .Z(n8452) );
  OR U9010 ( .A(n8646), .B(n8647), .Z(n8645) );
  AND U9011 ( .A(b[2]), .B(a[30]), .Z(n8643) );
  NAND U9012 ( .A(a[32]), .B(b[0]), .Z(n8277) );
  XNOR U9013 ( .A(n8641), .B(n8642), .Z(c[31]) );
  XOR U9014 ( .A(n8647), .B(n8646), .Z(n8642) );
  XOR U9015 ( .A(n8644), .B(n8648), .Z(n8646) );
  NAND U9016 ( .A(b[1]), .B(a[30]), .Z(n8648) );
  XOR U9017 ( .A(n8644), .B(n8640), .Z(n8649) );
  XOR U9018 ( .A(n8650), .B(n8638), .Z(n8640) );
  AND U9019 ( .A(b[2]), .B(a[29]), .Z(n8650) );
  ANDN U9020 ( .B(n8651), .A(n8652), .Z(n8644) );
  XOR U9021 ( .A(n8638), .B(n8634), .Z(n8653) );
  XNOR U9022 ( .A(n8633), .B(n8629), .Z(n8654) );
  XNOR U9023 ( .A(n8628), .B(n8624), .Z(n8655) );
  XNOR U9024 ( .A(n8623), .B(n8619), .Z(n8656) );
  XNOR U9025 ( .A(n8610), .B(n8609), .Z(n8657) );
  XOR U9026 ( .A(n8658), .B(n8608), .Z(n8609) );
  AND U9027 ( .A(b[7]), .B(a[24]), .Z(n8658) );
  XNOR U9028 ( .A(n8608), .B(n8614), .Z(n8659) );
  XNOR U9029 ( .A(n8613), .B(n8605), .Z(n8660) );
  XNOR U9030 ( .A(n8604), .B(n8600), .Z(n8661) );
  XNOR U9031 ( .A(n8599), .B(n8595), .Z(n8662) );
  XNOR U9032 ( .A(n8594), .B(n8590), .Z(n8663) );
  XNOR U9033 ( .A(n8581), .B(n8580), .Z(n8664) );
  XOR U9034 ( .A(n8665), .B(n8579), .Z(n8580) );
  AND U9035 ( .A(b[13]), .B(a[18]), .Z(n8665) );
  XNOR U9036 ( .A(n8579), .B(n8585), .Z(n8666) );
  XNOR U9037 ( .A(n8584), .B(n8576), .Z(n8667) );
  XNOR U9038 ( .A(n8575), .B(n8571), .Z(n8668) );
  XNOR U9039 ( .A(n8570), .B(n8566), .Z(n8669) );
  XNOR U9040 ( .A(n8565), .B(n8561), .Z(n8670) );
  XNOR U9041 ( .A(n8552), .B(n8551), .Z(n8671) );
  XOR U9042 ( .A(n8672), .B(n8550), .Z(n8551) );
  AND U9043 ( .A(b[19]), .B(a[12]), .Z(n8672) );
  XNOR U9044 ( .A(n8550), .B(n8556), .Z(n8673) );
  XNOR U9045 ( .A(n8555), .B(n8547), .Z(n8674) );
  XNOR U9046 ( .A(n8546), .B(n8542), .Z(n8675) );
  XNOR U9047 ( .A(n8541), .B(n8537), .Z(n8676) );
  XNOR U9048 ( .A(n8536), .B(n8532), .Z(n8677) );
  XNOR U9049 ( .A(n8523), .B(n8522), .Z(n8678) );
  XOR U9050 ( .A(n8679), .B(n8521), .Z(n8522) );
  AND U9051 ( .A(a[6]), .B(b[25]), .Z(n8679) );
  XNOR U9052 ( .A(n8521), .B(n8527), .Z(n8680) );
  XNOR U9053 ( .A(n8526), .B(n8518), .Z(n8681) );
  XNOR U9054 ( .A(n8517), .B(n8513), .Z(n8682) );
  XNOR U9055 ( .A(n8512), .B(n8508), .Z(n8683) );
  XNOR U9056 ( .A(n8507), .B(n8503), .Z(n8684) );
  XNOR U9057 ( .A(n8685), .B(n8502), .Z(n8503) );
  AND U9058 ( .A(a[0]), .B(b[31]), .Z(n8685) );
  XOR U9059 ( .A(n8686), .B(n8502), .Z(n8504) );
  XNOR U9060 ( .A(n8687), .B(n8688), .Z(n8502) );
  ANDN U9061 ( .B(n8689), .A(n8690), .Z(n8687) );
  AND U9062 ( .A(a[1]), .B(b[30]), .Z(n8686) );
  XNOR U9063 ( .A(n8691), .B(n8507), .Z(n8509) );
  XOR U9064 ( .A(n8692), .B(n8693), .Z(n8507) );
  ANDN U9065 ( .B(n8694), .A(n8695), .Z(n8692) );
  AND U9066 ( .A(a[2]), .B(b[29]), .Z(n8691) );
  XNOR U9067 ( .A(n8696), .B(n8512), .Z(n8514) );
  XOR U9068 ( .A(n8697), .B(n8698), .Z(n8512) );
  ANDN U9069 ( .B(n8699), .A(n8700), .Z(n8697) );
  AND U9070 ( .A(a[3]), .B(b[28]), .Z(n8696) );
  XNOR U9071 ( .A(n8701), .B(n8517), .Z(n8519) );
  XOR U9072 ( .A(n8702), .B(n8703), .Z(n8517) );
  ANDN U9073 ( .B(n8704), .A(n8705), .Z(n8702) );
  AND U9074 ( .A(a[4]), .B(b[27]), .Z(n8701) );
  XOR U9075 ( .A(n8706), .B(n8707), .Z(n8521) );
  AND U9076 ( .A(n8708), .B(n8709), .Z(n8706) );
  XNOR U9077 ( .A(n8710), .B(n8526), .Z(n8528) );
  XOR U9078 ( .A(n8711), .B(n8712), .Z(n8526) );
  ANDN U9079 ( .B(n8713), .A(n8714), .Z(n8711) );
  AND U9080 ( .A(a[5]), .B(b[26]), .Z(n8710) );
  XOR U9081 ( .A(n8715), .B(n8531), .Z(n8533) );
  XOR U9082 ( .A(n8716), .B(n8717), .Z(n8531) );
  ANDN U9083 ( .B(n8718), .A(n8719), .Z(n8716) );
  AND U9084 ( .A(a[7]), .B(b[24]), .Z(n8715) );
  XNOR U9085 ( .A(n8720), .B(n8536), .Z(n8538) );
  XOR U9086 ( .A(n8721), .B(n8722), .Z(n8536) );
  ANDN U9087 ( .B(n8723), .A(n8724), .Z(n8721) );
  AND U9088 ( .A(a[8]), .B(b[23]), .Z(n8720) );
  XNOR U9089 ( .A(n8725), .B(n8541), .Z(n8543) );
  XOR U9090 ( .A(n8726), .B(n8727), .Z(n8541) );
  ANDN U9091 ( .B(n8728), .A(n8729), .Z(n8726) );
  AND U9092 ( .A(a[9]), .B(b[22]), .Z(n8725) );
  XNOR U9093 ( .A(n8730), .B(n8546), .Z(n8548) );
  XOR U9094 ( .A(n8731), .B(n8732), .Z(n8546) );
  ANDN U9095 ( .B(n8733), .A(n8734), .Z(n8731) );
  AND U9096 ( .A(a[10]), .B(b[21]), .Z(n8730) );
  XOR U9097 ( .A(n8735), .B(n8736), .Z(n8550) );
  AND U9098 ( .A(n8737), .B(n8738), .Z(n8735) );
  XNOR U9099 ( .A(n8739), .B(n8555), .Z(n8557) );
  XOR U9100 ( .A(n8740), .B(n8741), .Z(n8555) );
  ANDN U9101 ( .B(n8742), .A(n8743), .Z(n8740) );
  AND U9102 ( .A(b[20]), .B(a[11]), .Z(n8739) );
  XOR U9103 ( .A(n8744), .B(n8560), .Z(n8562) );
  XOR U9104 ( .A(n8745), .B(n8746), .Z(n8560) );
  ANDN U9105 ( .B(n8747), .A(n8748), .Z(n8745) );
  AND U9106 ( .A(b[18]), .B(a[13]), .Z(n8744) );
  XNOR U9107 ( .A(n8749), .B(n8565), .Z(n8567) );
  XOR U9108 ( .A(n8750), .B(n8751), .Z(n8565) );
  ANDN U9109 ( .B(n8752), .A(n8753), .Z(n8750) );
  AND U9110 ( .A(b[17]), .B(a[14]), .Z(n8749) );
  XNOR U9111 ( .A(n8754), .B(n8570), .Z(n8572) );
  XOR U9112 ( .A(n8755), .B(n8756), .Z(n8570) );
  ANDN U9113 ( .B(n8757), .A(n8758), .Z(n8755) );
  AND U9114 ( .A(b[16]), .B(a[15]), .Z(n8754) );
  XNOR U9115 ( .A(n8759), .B(n8575), .Z(n8577) );
  XOR U9116 ( .A(n8760), .B(n8761), .Z(n8575) );
  ANDN U9117 ( .B(n8762), .A(n8763), .Z(n8760) );
  AND U9118 ( .A(a[16]), .B(b[15]), .Z(n8759) );
  XOR U9119 ( .A(n8764), .B(n8765), .Z(n8579) );
  AND U9120 ( .A(n8766), .B(n8767), .Z(n8764) );
  XNOR U9121 ( .A(n8768), .B(n8584), .Z(n8586) );
  XOR U9122 ( .A(n8769), .B(n8770), .Z(n8584) );
  ANDN U9123 ( .B(n8771), .A(n8772), .Z(n8769) );
  AND U9124 ( .A(b[14]), .B(a[17]), .Z(n8768) );
  XOR U9125 ( .A(n8773), .B(n8589), .Z(n8591) );
  XOR U9126 ( .A(n8774), .B(n8775), .Z(n8589) );
  ANDN U9127 ( .B(n8776), .A(n8777), .Z(n8774) );
  AND U9128 ( .A(b[12]), .B(a[19]), .Z(n8773) );
  XNOR U9129 ( .A(n8778), .B(n8594), .Z(n8596) );
  XOR U9130 ( .A(n8779), .B(n8780), .Z(n8594) );
  ANDN U9131 ( .B(n8781), .A(n8782), .Z(n8779) );
  AND U9132 ( .A(b[11]), .B(a[20]), .Z(n8778) );
  XNOR U9133 ( .A(n8783), .B(n8599), .Z(n8601) );
  XOR U9134 ( .A(n8784), .B(n8785), .Z(n8599) );
  ANDN U9135 ( .B(n8786), .A(n8787), .Z(n8784) );
  AND U9136 ( .A(b[10]), .B(a[21]), .Z(n8783) );
  XNOR U9137 ( .A(n8788), .B(n8604), .Z(n8606) );
  XOR U9138 ( .A(n8789), .B(n8790), .Z(n8604) );
  ANDN U9139 ( .B(n8791), .A(n8792), .Z(n8789) );
  AND U9140 ( .A(b[9]), .B(a[22]), .Z(n8788) );
  XOR U9141 ( .A(n8793), .B(n8794), .Z(n8608) );
  AND U9142 ( .A(n8795), .B(n8796), .Z(n8793) );
  XNOR U9143 ( .A(n8797), .B(n8613), .Z(n8615) );
  XOR U9144 ( .A(n8798), .B(n8799), .Z(n8613) );
  ANDN U9145 ( .B(n8800), .A(n8801), .Z(n8798) );
  AND U9146 ( .A(b[8]), .B(a[23]), .Z(n8797) );
  XOR U9147 ( .A(n8802), .B(n8618), .Z(n8620) );
  XOR U9148 ( .A(n8803), .B(n8804), .Z(n8618) );
  ANDN U9149 ( .B(n8805), .A(n8806), .Z(n8803) );
  AND U9150 ( .A(b[6]), .B(a[25]), .Z(n8802) );
  XNOR U9151 ( .A(n8807), .B(n8623), .Z(n8625) );
  XOR U9152 ( .A(n8808), .B(n8809), .Z(n8623) );
  ANDN U9153 ( .B(n8810), .A(n8811), .Z(n8808) );
  AND U9154 ( .A(b[5]), .B(a[26]), .Z(n8807) );
  XNOR U9155 ( .A(n8812), .B(n8628), .Z(n8630) );
  XOR U9156 ( .A(n8813), .B(n8814), .Z(n8628) );
  ANDN U9157 ( .B(n8815), .A(n8816), .Z(n8813) );
  AND U9158 ( .A(b[4]), .B(a[27]), .Z(n8812) );
  XNOR U9159 ( .A(n8817), .B(n8818), .Z(n8638) );
  NANDN U9160 ( .A(n8819), .B(n8820), .Z(n8818) );
  XNOR U9161 ( .A(n8821), .B(n8633), .Z(n8635) );
  XNOR U9162 ( .A(n8822), .B(n8823), .Z(n8633) );
  AND U9163 ( .A(n8824), .B(n8825), .Z(n8822) );
  AND U9164 ( .A(b[3]), .B(a[28]), .Z(n8821) );
  NAND U9165 ( .A(a[31]), .B(b[0]), .Z(n8641) );
  XNOR U9166 ( .A(n8652), .B(n8651), .Z(c[30]) );
  XNOR U9167 ( .A(n8819), .B(n8820), .Z(n8651) );
  XOR U9168 ( .A(n8817), .B(n8826), .Z(n8820) );
  NAND U9169 ( .A(b[1]), .B(a[29]), .Z(n8826) );
  XOR U9170 ( .A(n8825), .B(n8827), .Z(n8819) );
  XOR U9171 ( .A(n8817), .B(n8824), .Z(n8827) );
  XNOR U9172 ( .A(n8828), .B(n8823), .Z(n8824) );
  AND U9173 ( .A(b[2]), .B(a[28]), .Z(n8828) );
  NANDN U9174 ( .A(n8829), .B(n8830), .Z(n8817) );
  XOR U9175 ( .A(n8823), .B(n8815), .Z(n8831) );
  XNOR U9176 ( .A(n8814), .B(n8810), .Z(n8832) );
  XNOR U9177 ( .A(n8809), .B(n8805), .Z(n8833) );
  XNOR U9178 ( .A(n8796), .B(n8795), .Z(n8834) );
  XOR U9179 ( .A(n8835), .B(n8794), .Z(n8795) );
  AND U9180 ( .A(b[6]), .B(a[24]), .Z(n8835) );
  XNOR U9181 ( .A(n8794), .B(n8800), .Z(n8836) );
  XNOR U9182 ( .A(n8799), .B(n8791), .Z(n8837) );
  XNOR U9183 ( .A(n8790), .B(n8786), .Z(n8838) );
  XNOR U9184 ( .A(n8785), .B(n8781), .Z(n8839) );
  XNOR U9185 ( .A(n8780), .B(n8776), .Z(n8840) );
  XNOR U9186 ( .A(n8767), .B(n8766), .Z(n8841) );
  XOR U9187 ( .A(n8842), .B(n8765), .Z(n8766) );
  AND U9188 ( .A(b[12]), .B(a[18]), .Z(n8842) );
  XNOR U9189 ( .A(n8765), .B(n8771), .Z(n8843) );
  XNOR U9190 ( .A(n8770), .B(n8762), .Z(n8844) );
  XNOR U9191 ( .A(n8761), .B(n8757), .Z(n8845) );
  XNOR U9192 ( .A(n8756), .B(n8752), .Z(n8846) );
  XNOR U9193 ( .A(n8751), .B(n8747), .Z(n8847) );
  XNOR U9194 ( .A(n8738), .B(n8737), .Z(n8848) );
  XOR U9195 ( .A(n8849), .B(n8736), .Z(n8737) );
  AND U9196 ( .A(b[18]), .B(a[12]), .Z(n8849) );
  XNOR U9197 ( .A(n8736), .B(n8742), .Z(n8850) );
  XNOR U9198 ( .A(n8741), .B(n8733), .Z(n8851) );
  XNOR U9199 ( .A(n8732), .B(n8728), .Z(n8852) );
  XNOR U9200 ( .A(n8727), .B(n8723), .Z(n8853) );
  XNOR U9201 ( .A(n8722), .B(n8718), .Z(n8854) );
  XNOR U9202 ( .A(n8709), .B(n8708), .Z(n8855) );
  XOR U9203 ( .A(n8856), .B(n8707), .Z(n8708) );
  AND U9204 ( .A(a[6]), .B(b[24]), .Z(n8856) );
  XNOR U9205 ( .A(n8707), .B(n8713), .Z(n8857) );
  XNOR U9206 ( .A(n8712), .B(n8704), .Z(n8858) );
  XNOR U9207 ( .A(n8703), .B(n8699), .Z(n8859) );
  XNOR U9208 ( .A(n8698), .B(n8694), .Z(n8860) );
  XNOR U9209 ( .A(n8693), .B(n8689), .Z(n8861) );
  XOR U9210 ( .A(n8862), .B(n8688), .Z(n8689) );
  AND U9211 ( .A(a[0]), .B(b[30]), .Z(n8862) );
  XNOR U9212 ( .A(n8863), .B(n8688), .Z(n8690) );
  XNOR U9213 ( .A(n8864), .B(n8865), .Z(n8688) );
  ANDN U9214 ( .B(n8866), .A(n8867), .Z(n8864) );
  AND U9215 ( .A(a[1]), .B(b[29]), .Z(n8863) );
  XNOR U9216 ( .A(n8868), .B(n8693), .Z(n8695) );
  XOR U9217 ( .A(n8869), .B(n8870), .Z(n8693) );
  ANDN U9218 ( .B(n8871), .A(n8872), .Z(n8869) );
  AND U9219 ( .A(a[2]), .B(b[28]), .Z(n8868) );
  XNOR U9220 ( .A(n8873), .B(n8698), .Z(n8700) );
  XOR U9221 ( .A(n8874), .B(n8875), .Z(n8698) );
  ANDN U9222 ( .B(n8876), .A(n8877), .Z(n8874) );
  AND U9223 ( .A(a[3]), .B(b[27]), .Z(n8873) );
  XNOR U9224 ( .A(n8878), .B(n8703), .Z(n8705) );
  XOR U9225 ( .A(n8879), .B(n8880), .Z(n8703) );
  ANDN U9226 ( .B(n8881), .A(n8882), .Z(n8879) );
  AND U9227 ( .A(a[4]), .B(b[26]), .Z(n8878) );
  XOR U9228 ( .A(n8883), .B(n8884), .Z(n8707) );
  AND U9229 ( .A(n8885), .B(n8886), .Z(n8883) );
  XNOR U9230 ( .A(n8887), .B(n8712), .Z(n8714) );
  XOR U9231 ( .A(n8888), .B(n8889), .Z(n8712) );
  ANDN U9232 ( .B(n8890), .A(n8891), .Z(n8888) );
  AND U9233 ( .A(a[5]), .B(b[25]), .Z(n8887) );
  XOR U9234 ( .A(n8892), .B(n8717), .Z(n8719) );
  XOR U9235 ( .A(n8893), .B(n8894), .Z(n8717) );
  ANDN U9236 ( .B(n8895), .A(n8896), .Z(n8893) );
  AND U9237 ( .A(a[7]), .B(b[23]), .Z(n8892) );
  XNOR U9238 ( .A(n8897), .B(n8722), .Z(n8724) );
  XOR U9239 ( .A(n8898), .B(n8899), .Z(n8722) );
  ANDN U9240 ( .B(n8900), .A(n8901), .Z(n8898) );
  AND U9241 ( .A(a[8]), .B(b[22]), .Z(n8897) );
  XNOR U9242 ( .A(n8902), .B(n8727), .Z(n8729) );
  XOR U9243 ( .A(n8903), .B(n8904), .Z(n8727) );
  ANDN U9244 ( .B(n8905), .A(n8906), .Z(n8903) );
  AND U9245 ( .A(a[9]), .B(b[21]), .Z(n8902) );
  XNOR U9246 ( .A(n8907), .B(n8732), .Z(n8734) );
  XOR U9247 ( .A(n8908), .B(n8909), .Z(n8732) );
  ANDN U9248 ( .B(n8910), .A(n8911), .Z(n8908) );
  AND U9249 ( .A(b[20]), .B(a[10]), .Z(n8907) );
  XOR U9250 ( .A(n8912), .B(n8913), .Z(n8736) );
  AND U9251 ( .A(n8914), .B(n8915), .Z(n8912) );
  XNOR U9252 ( .A(n8916), .B(n8741), .Z(n8743) );
  XOR U9253 ( .A(n8917), .B(n8918), .Z(n8741) );
  ANDN U9254 ( .B(n8919), .A(n8920), .Z(n8917) );
  AND U9255 ( .A(b[19]), .B(a[11]), .Z(n8916) );
  XOR U9256 ( .A(n8921), .B(n8746), .Z(n8748) );
  XOR U9257 ( .A(n8922), .B(n8923), .Z(n8746) );
  ANDN U9258 ( .B(n8924), .A(n8925), .Z(n8922) );
  AND U9259 ( .A(b[17]), .B(a[13]), .Z(n8921) );
  XNOR U9260 ( .A(n8926), .B(n8751), .Z(n8753) );
  XOR U9261 ( .A(n8927), .B(n8928), .Z(n8751) );
  ANDN U9262 ( .B(n8929), .A(n8930), .Z(n8927) );
  AND U9263 ( .A(b[16]), .B(a[14]), .Z(n8926) );
  XNOR U9264 ( .A(n8931), .B(n8756), .Z(n8758) );
  XOR U9265 ( .A(n8932), .B(n8933), .Z(n8756) );
  ANDN U9266 ( .B(n8934), .A(n8935), .Z(n8932) );
  AND U9267 ( .A(a[15]), .B(b[15]), .Z(n8931) );
  XNOR U9268 ( .A(n8936), .B(n8761), .Z(n8763) );
  XOR U9269 ( .A(n8937), .B(n8938), .Z(n8761) );
  ANDN U9270 ( .B(n8939), .A(n8940), .Z(n8937) );
  AND U9271 ( .A(b[14]), .B(a[16]), .Z(n8936) );
  XOR U9272 ( .A(n8941), .B(n8942), .Z(n8765) );
  AND U9273 ( .A(n8943), .B(n8944), .Z(n8941) );
  XNOR U9274 ( .A(n8945), .B(n8770), .Z(n8772) );
  XOR U9275 ( .A(n8946), .B(n8947), .Z(n8770) );
  ANDN U9276 ( .B(n8948), .A(n8949), .Z(n8946) );
  AND U9277 ( .A(b[13]), .B(a[17]), .Z(n8945) );
  XOR U9278 ( .A(n8950), .B(n8775), .Z(n8777) );
  XOR U9279 ( .A(n8951), .B(n8952), .Z(n8775) );
  ANDN U9280 ( .B(n8953), .A(n8954), .Z(n8951) );
  AND U9281 ( .A(b[11]), .B(a[19]), .Z(n8950) );
  XNOR U9282 ( .A(n8955), .B(n8780), .Z(n8782) );
  XOR U9283 ( .A(n8956), .B(n8957), .Z(n8780) );
  ANDN U9284 ( .B(n8958), .A(n8959), .Z(n8956) );
  AND U9285 ( .A(b[10]), .B(a[20]), .Z(n8955) );
  XNOR U9286 ( .A(n8960), .B(n8785), .Z(n8787) );
  XOR U9287 ( .A(n8961), .B(n8962), .Z(n8785) );
  ANDN U9288 ( .B(n8963), .A(n8964), .Z(n8961) );
  AND U9289 ( .A(b[9]), .B(a[21]), .Z(n8960) );
  XNOR U9290 ( .A(n8965), .B(n8790), .Z(n8792) );
  XOR U9291 ( .A(n8966), .B(n8967), .Z(n8790) );
  ANDN U9292 ( .B(n8968), .A(n8969), .Z(n8966) );
  AND U9293 ( .A(b[8]), .B(a[22]), .Z(n8965) );
  XOR U9294 ( .A(n8970), .B(n8971), .Z(n8794) );
  AND U9295 ( .A(n8972), .B(n8973), .Z(n8970) );
  XNOR U9296 ( .A(n8974), .B(n8799), .Z(n8801) );
  XOR U9297 ( .A(n8975), .B(n8976), .Z(n8799) );
  ANDN U9298 ( .B(n8977), .A(n8978), .Z(n8975) );
  AND U9299 ( .A(b[7]), .B(a[23]), .Z(n8974) );
  XOR U9300 ( .A(n8979), .B(n8804), .Z(n8806) );
  XOR U9301 ( .A(n8980), .B(n8981), .Z(n8804) );
  ANDN U9302 ( .B(n8982), .A(n8983), .Z(n8980) );
  AND U9303 ( .A(b[5]), .B(a[25]), .Z(n8979) );
  XNOR U9304 ( .A(n8984), .B(n8809), .Z(n8811) );
  XOR U9305 ( .A(n8985), .B(n8986), .Z(n8809) );
  ANDN U9306 ( .B(n8987), .A(n8988), .Z(n8985) );
  AND U9307 ( .A(b[4]), .B(a[26]), .Z(n8984) );
  XNOR U9308 ( .A(n8989), .B(n8990), .Z(n8823) );
  NANDN U9309 ( .A(n8991), .B(n8992), .Z(n8990) );
  XNOR U9310 ( .A(n8993), .B(n8814), .Z(n8816) );
  XNOR U9311 ( .A(n8994), .B(n8995), .Z(n8814) );
  AND U9312 ( .A(n8996), .B(n8997), .Z(n8994) );
  AND U9313 ( .A(b[3]), .B(a[27]), .Z(n8993) );
  NAND U9314 ( .A(a[30]), .B(b[0]), .Z(n8652) );
  XNOR U9315 ( .A(n8998), .B(n8999), .Z(c[2]) );
  XNOR U9316 ( .A(n8829), .B(n8830), .Z(c[29]) );
  XNOR U9317 ( .A(n8991), .B(n8992), .Z(n8830) );
  XOR U9318 ( .A(n8989), .B(n9000), .Z(n8992) );
  NAND U9319 ( .A(b[1]), .B(a[28]), .Z(n9000) );
  XOR U9320 ( .A(n8997), .B(n9001), .Z(n8991) );
  XOR U9321 ( .A(n8989), .B(n8996), .Z(n9001) );
  XNOR U9322 ( .A(n9002), .B(n8995), .Z(n8996) );
  AND U9323 ( .A(b[2]), .B(a[27]), .Z(n9002) );
  NANDN U9324 ( .A(n9003), .B(n9004), .Z(n8989) );
  XOR U9325 ( .A(n8995), .B(n8987), .Z(n9005) );
  XNOR U9326 ( .A(n8986), .B(n8982), .Z(n9006) );
  XNOR U9327 ( .A(n8973), .B(n8972), .Z(n9007) );
  XOR U9328 ( .A(n9008), .B(n8971), .Z(n8972) );
  AND U9329 ( .A(b[5]), .B(a[24]), .Z(n9008) );
  XNOR U9330 ( .A(n8971), .B(n8977), .Z(n9009) );
  XNOR U9331 ( .A(n8976), .B(n8968), .Z(n9010) );
  XNOR U9332 ( .A(n8967), .B(n8963), .Z(n9011) );
  XNOR U9333 ( .A(n8962), .B(n8958), .Z(n9012) );
  XNOR U9334 ( .A(n8957), .B(n8953), .Z(n9013) );
  XNOR U9335 ( .A(n8944), .B(n8943), .Z(n9014) );
  XOR U9336 ( .A(n9015), .B(n8942), .Z(n8943) );
  AND U9337 ( .A(b[11]), .B(a[18]), .Z(n9015) );
  XNOR U9338 ( .A(n8942), .B(n8948), .Z(n9016) );
  XNOR U9339 ( .A(n8947), .B(n8939), .Z(n9017) );
  XNOR U9340 ( .A(n8938), .B(n8934), .Z(n9018) );
  XNOR U9341 ( .A(n8933), .B(n8929), .Z(n9019) );
  XNOR U9342 ( .A(n8928), .B(n8924), .Z(n9020) );
  XNOR U9343 ( .A(n8915), .B(n8914), .Z(n9021) );
  XOR U9344 ( .A(n9022), .B(n8913), .Z(n8914) );
  AND U9345 ( .A(b[17]), .B(a[12]), .Z(n9022) );
  XNOR U9346 ( .A(n8913), .B(n8919), .Z(n9023) );
  XNOR U9347 ( .A(n8918), .B(n8910), .Z(n9024) );
  XNOR U9348 ( .A(n8909), .B(n8905), .Z(n9025) );
  XNOR U9349 ( .A(n8904), .B(n8900), .Z(n9026) );
  XNOR U9350 ( .A(n8899), .B(n8895), .Z(n9027) );
  XNOR U9351 ( .A(n8886), .B(n8885), .Z(n9028) );
  XOR U9352 ( .A(n9029), .B(n8884), .Z(n8885) );
  AND U9353 ( .A(a[6]), .B(b[23]), .Z(n9029) );
  XNOR U9354 ( .A(n8884), .B(n8890), .Z(n9030) );
  XNOR U9355 ( .A(n8889), .B(n8881), .Z(n9031) );
  XNOR U9356 ( .A(n8880), .B(n8876), .Z(n9032) );
  XNOR U9357 ( .A(n8875), .B(n8871), .Z(n9033) );
  XNOR U9358 ( .A(n8870), .B(n8866), .Z(n9034) );
  XNOR U9359 ( .A(n9035), .B(n8865), .Z(n8866) );
  AND U9360 ( .A(a[0]), .B(b[29]), .Z(n9035) );
  XOR U9361 ( .A(n9036), .B(n8865), .Z(n8867) );
  XNOR U9362 ( .A(n9037), .B(n9038), .Z(n8865) );
  ANDN U9363 ( .B(n9039), .A(n9040), .Z(n9037) );
  AND U9364 ( .A(a[1]), .B(b[28]), .Z(n9036) );
  XNOR U9365 ( .A(n9041), .B(n8870), .Z(n8872) );
  XOR U9366 ( .A(n9042), .B(n9043), .Z(n8870) );
  ANDN U9367 ( .B(n9044), .A(n9045), .Z(n9042) );
  AND U9368 ( .A(a[2]), .B(b[27]), .Z(n9041) );
  XNOR U9369 ( .A(n9046), .B(n8875), .Z(n8877) );
  XOR U9370 ( .A(n9047), .B(n9048), .Z(n8875) );
  ANDN U9371 ( .B(n9049), .A(n9050), .Z(n9047) );
  AND U9372 ( .A(a[3]), .B(b[26]), .Z(n9046) );
  XNOR U9373 ( .A(n9051), .B(n8880), .Z(n8882) );
  XOR U9374 ( .A(n9052), .B(n9053), .Z(n8880) );
  ANDN U9375 ( .B(n9054), .A(n9055), .Z(n9052) );
  AND U9376 ( .A(a[4]), .B(b[25]), .Z(n9051) );
  XOR U9377 ( .A(n9056), .B(n9057), .Z(n8884) );
  AND U9378 ( .A(n9058), .B(n9059), .Z(n9056) );
  XNOR U9379 ( .A(n9060), .B(n8889), .Z(n8891) );
  XOR U9380 ( .A(n9061), .B(n9062), .Z(n8889) );
  ANDN U9381 ( .B(n9063), .A(n9064), .Z(n9061) );
  AND U9382 ( .A(a[5]), .B(b[24]), .Z(n9060) );
  XOR U9383 ( .A(n9065), .B(n8894), .Z(n8896) );
  XOR U9384 ( .A(n9066), .B(n9067), .Z(n8894) );
  ANDN U9385 ( .B(n9068), .A(n9069), .Z(n9066) );
  AND U9386 ( .A(a[7]), .B(b[22]), .Z(n9065) );
  XNOR U9387 ( .A(n9070), .B(n8899), .Z(n8901) );
  XOR U9388 ( .A(n9071), .B(n9072), .Z(n8899) );
  ANDN U9389 ( .B(n9073), .A(n9074), .Z(n9071) );
  AND U9390 ( .A(a[8]), .B(b[21]), .Z(n9070) );
  XNOR U9391 ( .A(n9075), .B(n8904), .Z(n8906) );
  XOR U9392 ( .A(n9076), .B(n9077), .Z(n8904) );
  ANDN U9393 ( .B(n9078), .A(n9079), .Z(n9076) );
  AND U9394 ( .A(a[9]), .B(b[20]), .Z(n9075) );
  XNOR U9395 ( .A(n9080), .B(n8909), .Z(n8911) );
  XOR U9396 ( .A(n9081), .B(n9082), .Z(n8909) );
  ANDN U9397 ( .B(n9083), .A(n9084), .Z(n9081) );
  AND U9398 ( .A(b[19]), .B(a[10]), .Z(n9080) );
  XOR U9399 ( .A(n9085), .B(n9086), .Z(n8913) );
  AND U9400 ( .A(n9087), .B(n9088), .Z(n9085) );
  XNOR U9401 ( .A(n9089), .B(n8918), .Z(n8920) );
  XOR U9402 ( .A(n9090), .B(n9091), .Z(n8918) );
  ANDN U9403 ( .B(n9092), .A(n9093), .Z(n9090) );
  AND U9404 ( .A(b[18]), .B(a[11]), .Z(n9089) );
  XOR U9405 ( .A(n9094), .B(n8923), .Z(n8925) );
  XOR U9406 ( .A(n9095), .B(n9096), .Z(n8923) );
  ANDN U9407 ( .B(n9097), .A(n9098), .Z(n9095) );
  AND U9408 ( .A(b[16]), .B(a[13]), .Z(n9094) );
  XNOR U9409 ( .A(n9099), .B(n8928), .Z(n8930) );
  XOR U9410 ( .A(n9100), .B(n9101), .Z(n8928) );
  ANDN U9411 ( .B(n9102), .A(n9103), .Z(n9100) );
  AND U9412 ( .A(a[14]), .B(b[15]), .Z(n9099) );
  XNOR U9413 ( .A(n9104), .B(n8933), .Z(n8935) );
  XOR U9414 ( .A(n9105), .B(n9106), .Z(n8933) );
  ANDN U9415 ( .B(n9107), .A(n9108), .Z(n9105) );
  AND U9416 ( .A(b[14]), .B(a[15]), .Z(n9104) );
  XNOR U9417 ( .A(n9109), .B(n8938), .Z(n8940) );
  XOR U9418 ( .A(n9110), .B(n9111), .Z(n8938) );
  ANDN U9419 ( .B(n9112), .A(n9113), .Z(n9110) );
  AND U9420 ( .A(b[13]), .B(a[16]), .Z(n9109) );
  XOR U9421 ( .A(n9114), .B(n9115), .Z(n8942) );
  AND U9422 ( .A(n9116), .B(n9117), .Z(n9114) );
  XNOR U9423 ( .A(n9118), .B(n8947), .Z(n8949) );
  XOR U9424 ( .A(n9119), .B(n9120), .Z(n8947) );
  ANDN U9425 ( .B(n9121), .A(n9122), .Z(n9119) );
  AND U9426 ( .A(b[12]), .B(a[17]), .Z(n9118) );
  XOR U9427 ( .A(n9123), .B(n8952), .Z(n8954) );
  XOR U9428 ( .A(n9124), .B(n9125), .Z(n8952) );
  ANDN U9429 ( .B(n9126), .A(n9127), .Z(n9124) );
  AND U9430 ( .A(b[10]), .B(a[19]), .Z(n9123) );
  XNOR U9431 ( .A(n9128), .B(n8957), .Z(n8959) );
  XOR U9432 ( .A(n9129), .B(n9130), .Z(n8957) );
  ANDN U9433 ( .B(n9131), .A(n9132), .Z(n9129) );
  AND U9434 ( .A(b[9]), .B(a[20]), .Z(n9128) );
  XNOR U9435 ( .A(n9133), .B(n8962), .Z(n8964) );
  XOR U9436 ( .A(n9134), .B(n9135), .Z(n8962) );
  ANDN U9437 ( .B(n9136), .A(n9137), .Z(n9134) );
  AND U9438 ( .A(b[8]), .B(a[21]), .Z(n9133) );
  XNOR U9439 ( .A(n9138), .B(n8967), .Z(n8969) );
  XOR U9440 ( .A(n9139), .B(n9140), .Z(n8967) );
  ANDN U9441 ( .B(n9141), .A(n9142), .Z(n9139) );
  AND U9442 ( .A(b[7]), .B(a[22]), .Z(n9138) );
  XOR U9443 ( .A(n9143), .B(n9144), .Z(n8971) );
  AND U9444 ( .A(n9145), .B(n9146), .Z(n9143) );
  XNOR U9445 ( .A(n9147), .B(n8976), .Z(n8978) );
  XOR U9446 ( .A(n9148), .B(n9149), .Z(n8976) );
  ANDN U9447 ( .B(n9150), .A(n9151), .Z(n9148) );
  AND U9448 ( .A(b[6]), .B(a[23]), .Z(n9147) );
  XOR U9449 ( .A(n9152), .B(n8981), .Z(n8983) );
  XOR U9450 ( .A(n9153), .B(n9154), .Z(n8981) );
  ANDN U9451 ( .B(n9155), .A(n9156), .Z(n9153) );
  AND U9452 ( .A(b[4]), .B(a[25]), .Z(n9152) );
  XNOR U9453 ( .A(n9157), .B(n9158), .Z(n8995) );
  NANDN U9454 ( .A(n9159), .B(n9160), .Z(n9158) );
  XNOR U9455 ( .A(n9161), .B(n8986), .Z(n8988) );
  XNOR U9456 ( .A(n9162), .B(n9163), .Z(n8986) );
  AND U9457 ( .A(n9164), .B(n9165), .Z(n9162) );
  AND U9458 ( .A(b[3]), .B(a[26]), .Z(n9161) );
  NAND U9459 ( .A(a[29]), .B(b[0]), .Z(n8829) );
  XNOR U9460 ( .A(n9003), .B(n9004), .Z(c[28]) );
  XNOR U9461 ( .A(n9159), .B(n9160), .Z(n9004) );
  XOR U9462 ( .A(n9157), .B(n9166), .Z(n9160) );
  NAND U9463 ( .A(b[1]), .B(a[27]), .Z(n9166) );
  XOR U9464 ( .A(n9165), .B(n9167), .Z(n9159) );
  XOR U9465 ( .A(n9157), .B(n9164), .Z(n9167) );
  XNOR U9466 ( .A(n9168), .B(n9163), .Z(n9164) );
  AND U9467 ( .A(b[2]), .B(a[26]), .Z(n9168) );
  NANDN U9468 ( .A(n9169), .B(n9170), .Z(n9157) );
  XOR U9469 ( .A(n9163), .B(n9155), .Z(n9171) );
  XNOR U9470 ( .A(n9146), .B(n9145), .Z(n9172) );
  XOR U9471 ( .A(n9173), .B(n9144), .Z(n9145) );
  AND U9472 ( .A(b[4]), .B(a[24]), .Z(n9173) );
  XNOR U9473 ( .A(n9144), .B(n9150), .Z(n9174) );
  XNOR U9474 ( .A(n9149), .B(n9141), .Z(n9175) );
  XNOR U9475 ( .A(n9140), .B(n9136), .Z(n9176) );
  XNOR U9476 ( .A(n9135), .B(n9131), .Z(n9177) );
  XNOR U9477 ( .A(n9130), .B(n9126), .Z(n9178) );
  XNOR U9478 ( .A(n9117), .B(n9116), .Z(n9179) );
  XOR U9479 ( .A(n9180), .B(n9115), .Z(n9116) );
  AND U9480 ( .A(b[10]), .B(a[18]), .Z(n9180) );
  XNOR U9481 ( .A(n9115), .B(n9121), .Z(n9181) );
  XNOR U9482 ( .A(n9120), .B(n9112), .Z(n9182) );
  XNOR U9483 ( .A(n9111), .B(n9107), .Z(n9183) );
  XNOR U9484 ( .A(n9106), .B(n9102), .Z(n9184) );
  XNOR U9485 ( .A(n9101), .B(n9097), .Z(n9185) );
  XNOR U9486 ( .A(n9088), .B(n9087), .Z(n9186) );
  XOR U9487 ( .A(n9187), .B(n9086), .Z(n9087) );
  AND U9488 ( .A(b[16]), .B(a[12]), .Z(n9187) );
  XNOR U9489 ( .A(n9086), .B(n9092), .Z(n9188) );
  XNOR U9490 ( .A(n9091), .B(n9083), .Z(n9189) );
  XNOR U9491 ( .A(n9082), .B(n9078), .Z(n9190) );
  XNOR U9492 ( .A(n9077), .B(n9073), .Z(n9191) );
  XNOR U9493 ( .A(n9072), .B(n9068), .Z(n9192) );
  XNOR U9494 ( .A(n9059), .B(n9058), .Z(n9193) );
  XOR U9495 ( .A(n9194), .B(n9057), .Z(n9058) );
  AND U9496 ( .A(a[6]), .B(b[22]), .Z(n9194) );
  XNOR U9497 ( .A(n9057), .B(n9063), .Z(n9195) );
  XNOR U9498 ( .A(n9062), .B(n9054), .Z(n9196) );
  XNOR U9499 ( .A(n9053), .B(n9049), .Z(n9197) );
  XNOR U9500 ( .A(n9048), .B(n9044), .Z(n9198) );
  XNOR U9501 ( .A(n9043), .B(n9039), .Z(n9199) );
  XOR U9502 ( .A(n9200), .B(n9038), .Z(n9039) );
  AND U9503 ( .A(a[0]), .B(b[28]), .Z(n9200) );
  XNOR U9504 ( .A(n9201), .B(n9038), .Z(n9040) );
  XNOR U9505 ( .A(n9202), .B(n9203), .Z(n9038) );
  ANDN U9506 ( .B(n9204), .A(n9205), .Z(n9202) );
  AND U9507 ( .A(a[1]), .B(b[27]), .Z(n9201) );
  XNOR U9508 ( .A(n9206), .B(n9043), .Z(n9045) );
  XOR U9509 ( .A(n9207), .B(n9208), .Z(n9043) );
  ANDN U9510 ( .B(n9209), .A(n9210), .Z(n9207) );
  AND U9511 ( .A(a[2]), .B(b[26]), .Z(n9206) );
  XNOR U9512 ( .A(n9211), .B(n9048), .Z(n9050) );
  XOR U9513 ( .A(n9212), .B(n9213), .Z(n9048) );
  ANDN U9514 ( .B(n9214), .A(n9215), .Z(n9212) );
  AND U9515 ( .A(a[3]), .B(b[25]), .Z(n9211) );
  XNOR U9516 ( .A(n9216), .B(n9053), .Z(n9055) );
  XOR U9517 ( .A(n9217), .B(n9218), .Z(n9053) );
  ANDN U9518 ( .B(n9219), .A(n9220), .Z(n9217) );
  AND U9519 ( .A(a[4]), .B(b[24]), .Z(n9216) );
  XOR U9520 ( .A(n9221), .B(n9222), .Z(n9057) );
  AND U9521 ( .A(n9223), .B(n9224), .Z(n9221) );
  XNOR U9522 ( .A(n9225), .B(n9062), .Z(n9064) );
  XOR U9523 ( .A(n9226), .B(n9227), .Z(n9062) );
  ANDN U9524 ( .B(n9228), .A(n9229), .Z(n9226) );
  AND U9525 ( .A(a[5]), .B(b[23]), .Z(n9225) );
  XOR U9526 ( .A(n9230), .B(n9067), .Z(n9069) );
  XOR U9527 ( .A(n9231), .B(n9232), .Z(n9067) );
  ANDN U9528 ( .B(n9233), .A(n9234), .Z(n9231) );
  AND U9529 ( .A(a[7]), .B(b[21]), .Z(n9230) );
  XNOR U9530 ( .A(n9235), .B(n9072), .Z(n9074) );
  XOR U9531 ( .A(n9236), .B(n9237), .Z(n9072) );
  ANDN U9532 ( .B(n9238), .A(n9239), .Z(n9236) );
  AND U9533 ( .A(a[8]), .B(b[20]), .Z(n9235) );
  XNOR U9534 ( .A(n9240), .B(n9077), .Z(n9079) );
  XOR U9535 ( .A(n9241), .B(n9242), .Z(n9077) );
  ANDN U9536 ( .B(n9243), .A(n9244), .Z(n9241) );
  AND U9537 ( .A(a[9]), .B(b[19]), .Z(n9240) );
  XNOR U9538 ( .A(n9245), .B(n9082), .Z(n9084) );
  XOR U9539 ( .A(n9246), .B(n9247), .Z(n9082) );
  ANDN U9540 ( .B(n9248), .A(n9249), .Z(n9246) );
  AND U9541 ( .A(b[18]), .B(a[10]), .Z(n9245) );
  XOR U9542 ( .A(n9250), .B(n9251), .Z(n9086) );
  AND U9543 ( .A(n9252), .B(n9253), .Z(n9250) );
  XNOR U9544 ( .A(n9254), .B(n9091), .Z(n9093) );
  XOR U9545 ( .A(n9255), .B(n9256), .Z(n9091) );
  ANDN U9546 ( .B(n9257), .A(n9258), .Z(n9255) );
  AND U9547 ( .A(b[17]), .B(a[11]), .Z(n9254) );
  XOR U9548 ( .A(n9259), .B(n9096), .Z(n9098) );
  XOR U9549 ( .A(n9260), .B(n9261), .Z(n9096) );
  ANDN U9550 ( .B(n9262), .A(n9263), .Z(n9260) );
  AND U9551 ( .A(a[13]), .B(b[15]), .Z(n9259) );
  XNOR U9552 ( .A(n9264), .B(n9101), .Z(n9103) );
  XOR U9553 ( .A(n9265), .B(n9266), .Z(n9101) );
  ANDN U9554 ( .B(n9267), .A(n9268), .Z(n9265) );
  AND U9555 ( .A(b[14]), .B(a[14]), .Z(n9264) );
  XNOR U9556 ( .A(n9269), .B(n9106), .Z(n9108) );
  XOR U9557 ( .A(n9270), .B(n9271), .Z(n9106) );
  ANDN U9558 ( .B(n9272), .A(n9273), .Z(n9270) );
  AND U9559 ( .A(b[13]), .B(a[15]), .Z(n9269) );
  XNOR U9560 ( .A(n9274), .B(n9111), .Z(n9113) );
  XOR U9561 ( .A(n9275), .B(n9276), .Z(n9111) );
  ANDN U9562 ( .B(n9277), .A(n9278), .Z(n9275) );
  AND U9563 ( .A(b[12]), .B(a[16]), .Z(n9274) );
  XOR U9564 ( .A(n9279), .B(n9280), .Z(n9115) );
  AND U9565 ( .A(n9281), .B(n9282), .Z(n9279) );
  XNOR U9566 ( .A(n9283), .B(n9120), .Z(n9122) );
  XOR U9567 ( .A(n9284), .B(n9285), .Z(n9120) );
  ANDN U9568 ( .B(n9286), .A(n9287), .Z(n9284) );
  AND U9569 ( .A(b[11]), .B(a[17]), .Z(n9283) );
  XOR U9570 ( .A(n9288), .B(n9125), .Z(n9127) );
  XOR U9571 ( .A(n9289), .B(n9290), .Z(n9125) );
  ANDN U9572 ( .B(n9291), .A(n9292), .Z(n9289) );
  AND U9573 ( .A(b[9]), .B(a[19]), .Z(n9288) );
  XNOR U9574 ( .A(n9293), .B(n9130), .Z(n9132) );
  XOR U9575 ( .A(n9294), .B(n9295), .Z(n9130) );
  ANDN U9576 ( .B(n9296), .A(n9297), .Z(n9294) );
  AND U9577 ( .A(b[8]), .B(a[20]), .Z(n9293) );
  XNOR U9578 ( .A(n9298), .B(n9135), .Z(n9137) );
  XOR U9579 ( .A(n9299), .B(n9300), .Z(n9135) );
  ANDN U9580 ( .B(n9301), .A(n9302), .Z(n9299) );
  AND U9581 ( .A(b[7]), .B(a[21]), .Z(n9298) );
  XNOR U9582 ( .A(n9303), .B(n9140), .Z(n9142) );
  XOR U9583 ( .A(n9304), .B(n9305), .Z(n9140) );
  ANDN U9584 ( .B(n9306), .A(n9307), .Z(n9304) );
  AND U9585 ( .A(b[6]), .B(a[22]), .Z(n9303) );
  XOR U9586 ( .A(n9308), .B(n9309), .Z(n9144) );
  AND U9587 ( .A(n9310), .B(n9311), .Z(n9308) );
  XNOR U9588 ( .A(n9312), .B(n9149), .Z(n9151) );
  XOR U9589 ( .A(n9313), .B(n9314), .Z(n9149) );
  ANDN U9590 ( .B(n9315), .A(n9316), .Z(n9313) );
  AND U9591 ( .A(b[5]), .B(a[23]), .Z(n9312) );
  XNOR U9592 ( .A(n9317), .B(n9318), .Z(n9163) );
  NANDN U9593 ( .A(n9319), .B(n9320), .Z(n9318) );
  XOR U9594 ( .A(n9321), .B(n9154), .Z(n9156) );
  XOR U9595 ( .A(n9322), .B(n9323), .Z(n9154) );
  ANDN U9596 ( .B(n9324), .A(n9325), .Z(n9322) );
  AND U9597 ( .A(b[3]), .B(a[25]), .Z(n9321) );
  NAND U9598 ( .A(a[28]), .B(b[0]), .Z(n9003) );
  XNOR U9599 ( .A(n9169), .B(n9170), .Z(c[27]) );
  XNOR U9600 ( .A(n9319), .B(n9320), .Z(n9170) );
  XOR U9601 ( .A(n9317), .B(n9326), .Z(n9320) );
  NAND U9602 ( .A(b[1]), .B(a[26]), .Z(n9326) );
  XNOR U9603 ( .A(n9325), .B(n9327), .Z(n9319) );
  XOR U9604 ( .A(n9317), .B(n9324), .Z(n9327) );
  XNOR U9605 ( .A(n9328), .B(n9323), .Z(n9324) );
  AND U9606 ( .A(b[2]), .B(a[25]), .Z(n9328) );
  NANDN U9607 ( .A(n9329), .B(n9330), .Z(n9317) );
  XNOR U9608 ( .A(n9323), .B(n9331), .Z(n9325) );
  XNOR U9609 ( .A(n9311), .B(n9310), .Z(n9331) );
  XOR U9610 ( .A(n9332), .B(n9309), .Z(n9310) );
  AND U9611 ( .A(b[3]), .B(a[24]), .Z(n9332) );
  XNOR U9612 ( .A(n9309), .B(n9315), .Z(n9333) );
  XNOR U9613 ( .A(n9314), .B(n9306), .Z(n9334) );
  XNOR U9614 ( .A(n9305), .B(n9301), .Z(n9335) );
  XNOR U9615 ( .A(n9300), .B(n9296), .Z(n9336) );
  XNOR U9616 ( .A(n9295), .B(n9291), .Z(n9337) );
  XNOR U9617 ( .A(n9282), .B(n9281), .Z(n9338) );
  XOR U9618 ( .A(n9339), .B(n9280), .Z(n9281) );
  AND U9619 ( .A(b[9]), .B(a[18]), .Z(n9339) );
  XNOR U9620 ( .A(n9280), .B(n9286), .Z(n9340) );
  XNOR U9621 ( .A(n9285), .B(n9277), .Z(n9341) );
  XNOR U9622 ( .A(n9276), .B(n9272), .Z(n9342) );
  XNOR U9623 ( .A(n9271), .B(n9267), .Z(n9343) );
  XNOR U9624 ( .A(n9266), .B(n9262), .Z(n9344) );
  XNOR U9625 ( .A(n9253), .B(n9252), .Z(n9345) );
  XOR U9626 ( .A(n9346), .B(n9251), .Z(n9252) );
  AND U9627 ( .A(b[15]), .B(a[12]), .Z(n9346) );
  XNOR U9628 ( .A(n9251), .B(n9257), .Z(n9347) );
  XNOR U9629 ( .A(n9256), .B(n9248), .Z(n9348) );
  XNOR U9630 ( .A(n9247), .B(n9243), .Z(n9349) );
  XNOR U9631 ( .A(n9242), .B(n9238), .Z(n9350) );
  XNOR U9632 ( .A(n9237), .B(n9233), .Z(n9351) );
  XNOR U9633 ( .A(n9224), .B(n9223), .Z(n9352) );
  XOR U9634 ( .A(n9353), .B(n9222), .Z(n9223) );
  AND U9635 ( .A(a[6]), .B(b[21]), .Z(n9353) );
  XNOR U9636 ( .A(n9222), .B(n9228), .Z(n9354) );
  XNOR U9637 ( .A(n9227), .B(n9219), .Z(n9355) );
  XNOR U9638 ( .A(n9218), .B(n9214), .Z(n9356) );
  XNOR U9639 ( .A(n9213), .B(n9209), .Z(n9357) );
  XNOR U9640 ( .A(n9208), .B(n9204), .Z(n9358) );
  XNOR U9641 ( .A(n9359), .B(n9203), .Z(n9204) );
  AND U9642 ( .A(a[0]), .B(b[27]), .Z(n9359) );
  XOR U9643 ( .A(n9360), .B(n9203), .Z(n9205) );
  XNOR U9644 ( .A(n9361), .B(n9362), .Z(n9203) );
  ANDN U9645 ( .B(n9363), .A(n9364), .Z(n9361) );
  AND U9646 ( .A(a[1]), .B(b[26]), .Z(n9360) );
  XNOR U9647 ( .A(n9365), .B(n9208), .Z(n9210) );
  XOR U9648 ( .A(n9366), .B(n9367), .Z(n9208) );
  ANDN U9649 ( .B(n9368), .A(n9369), .Z(n9366) );
  AND U9650 ( .A(a[2]), .B(b[25]), .Z(n9365) );
  XNOR U9651 ( .A(n9370), .B(n9213), .Z(n9215) );
  XOR U9652 ( .A(n9371), .B(n9372), .Z(n9213) );
  ANDN U9653 ( .B(n9373), .A(n9374), .Z(n9371) );
  AND U9654 ( .A(a[3]), .B(b[24]), .Z(n9370) );
  XNOR U9655 ( .A(n9375), .B(n9218), .Z(n9220) );
  XOR U9656 ( .A(n9376), .B(n9377), .Z(n9218) );
  ANDN U9657 ( .B(n9378), .A(n9379), .Z(n9376) );
  AND U9658 ( .A(a[4]), .B(b[23]), .Z(n9375) );
  XOR U9659 ( .A(n9380), .B(n9381), .Z(n9222) );
  AND U9660 ( .A(n9382), .B(n9383), .Z(n9380) );
  XNOR U9661 ( .A(n9384), .B(n9227), .Z(n9229) );
  XOR U9662 ( .A(n9385), .B(n9386), .Z(n9227) );
  ANDN U9663 ( .B(n9387), .A(n9388), .Z(n9385) );
  AND U9664 ( .A(a[5]), .B(b[22]), .Z(n9384) );
  XOR U9665 ( .A(n9389), .B(n9232), .Z(n9234) );
  XOR U9666 ( .A(n9390), .B(n9391), .Z(n9232) );
  ANDN U9667 ( .B(n9392), .A(n9393), .Z(n9390) );
  AND U9668 ( .A(a[7]), .B(b[20]), .Z(n9389) );
  XNOR U9669 ( .A(n9394), .B(n9237), .Z(n9239) );
  XOR U9670 ( .A(n9395), .B(n9396), .Z(n9237) );
  ANDN U9671 ( .B(n9397), .A(n9398), .Z(n9395) );
  AND U9672 ( .A(a[8]), .B(b[19]), .Z(n9394) );
  XNOR U9673 ( .A(n9399), .B(n9242), .Z(n9244) );
  XOR U9674 ( .A(n9400), .B(n9401), .Z(n9242) );
  ANDN U9675 ( .B(n9402), .A(n9403), .Z(n9400) );
  AND U9676 ( .A(a[9]), .B(b[18]), .Z(n9399) );
  XNOR U9677 ( .A(n9404), .B(n9247), .Z(n9249) );
  XOR U9678 ( .A(n9405), .B(n9406), .Z(n9247) );
  ANDN U9679 ( .B(n9407), .A(n9408), .Z(n9405) );
  AND U9680 ( .A(b[17]), .B(a[10]), .Z(n9404) );
  XOR U9681 ( .A(n9409), .B(n9410), .Z(n9251) );
  AND U9682 ( .A(n9411), .B(n9412), .Z(n9409) );
  XNOR U9683 ( .A(n9413), .B(n9256), .Z(n9258) );
  XOR U9684 ( .A(n9414), .B(n9415), .Z(n9256) );
  ANDN U9685 ( .B(n9416), .A(n9417), .Z(n9414) );
  AND U9686 ( .A(b[16]), .B(a[11]), .Z(n9413) );
  XOR U9687 ( .A(n9418), .B(n9261), .Z(n9263) );
  XOR U9688 ( .A(n9419), .B(n9420), .Z(n9261) );
  ANDN U9689 ( .B(n9421), .A(n9422), .Z(n9419) );
  AND U9690 ( .A(b[14]), .B(a[13]), .Z(n9418) );
  XNOR U9691 ( .A(n9423), .B(n9266), .Z(n9268) );
  XOR U9692 ( .A(n9424), .B(n9425), .Z(n9266) );
  ANDN U9693 ( .B(n9426), .A(n9427), .Z(n9424) );
  AND U9694 ( .A(b[13]), .B(a[14]), .Z(n9423) );
  XNOR U9695 ( .A(n9428), .B(n9271), .Z(n9273) );
  XOR U9696 ( .A(n9429), .B(n9430), .Z(n9271) );
  ANDN U9697 ( .B(n9431), .A(n9432), .Z(n9429) );
  AND U9698 ( .A(b[12]), .B(a[15]), .Z(n9428) );
  XNOR U9699 ( .A(n9433), .B(n9276), .Z(n9278) );
  XOR U9700 ( .A(n9434), .B(n9435), .Z(n9276) );
  ANDN U9701 ( .B(n9436), .A(n9437), .Z(n9434) );
  AND U9702 ( .A(b[11]), .B(a[16]), .Z(n9433) );
  XOR U9703 ( .A(n9438), .B(n9439), .Z(n9280) );
  AND U9704 ( .A(n9440), .B(n9441), .Z(n9438) );
  XNOR U9705 ( .A(n9442), .B(n9285), .Z(n9287) );
  XOR U9706 ( .A(n9443), .B(n9444), .Z(n9285) );
  ANDN U9707 ( .B(n9445), .A(n9446), .Z(n9443) );
  AND U9708 ( .A(b[10]), .B(a[17]), .Z(n9442) );
  XOR U9709 ( .A(n9447), .B(n9290), .Z(n9292) );
  XOR U9710 ( .A(n9448), .B(n9449), .Z(n9290) );
  ANDN U9711 ( .B(n9450), .A(n9451), .Z(n9448) );
  AND U9712 ( .A(b[8]), .B(a[19]), .Z(n9447) );
  XNOR U9713 ( .A(n9452), .B(n9295), .Z(n9297) );
  XOR U9714 ( .A(n9453), .B(n9454), .Z(n9295) );
  ANDN U9715 ( .B(n9455), .A(n9456), .Z(n9453) );
  AND U9716 ( .A(b[7]), .B(a[20]), .Z(n9452) );
  XNOR U9717 ( .A(n9457), .B(n9300), .Z(n9302) );
  XOR U9718 ( .A(n9458), .B(n9459), .Z(n9300) );
  ANDN U9719 ( .B(n9460), .A(n9461), .Z(n9458) );
  AND U9720 ( .A(b[6]), .B(a[21]), .Z(n9457) );
  XNOR U9721 ( .A(n9462), .B(n9305), .Z(n9307) );
  XOR U9722 ( .A(n9463), .B(n9464), .Z(n9305) );
  ANDN U9723 ( .B(n9465), .A(n9466), .Z(n9463) );
  AND U9724 ( .A(b[5]), .B(a[22]), .Z(n9462) );
  XOR U9725 ( .A(n9467), .B(n9468), .Z(n9309) );
  ANDN U9726 ( .B(n9469), .A(n9470), .Z(n9467) );
  XNOR U9727 ( .A(n9471), .B(n9314), .Z(n9316) );
  XOR U9728 ( .A(n9472), .B(n9473), .Z(n9314) );
  ANDN U9729 ( .B(n9474), .A(n9475), .Z(n9472) );
  AND U9730 ( .A(b[4]), .B(a[23]), .Z(n9471) );
  XNOR U9731 ( .A(n9476), .B(n9477), .Z(n9323) );
  NAND U9732 ( .A(n9478), .B(n9479), .Z(n9477) );
  NAND U9733 ( .A(a[27]), .B(b[0]), .Z(n9169) );
  XNOR U9734 ( .A(n9329), .B(n9330), .Z(c[26]) );
  XOR U9735 ( .A(n9478), .B(n9479), .Z(n9330) );
  XOR U9736 ( .A(n9476), .B(n9480), .Z(n9479) );
  NAND U9737 ( .A(b[1]), .B(a[25]), .Z(n9480) );
  XOR U9738 ( .A(n9476), .B(n9469), .Z(n9481) );
  XNOR U9739 ( .A(n9468), .B(n9474), .Z(n9482) );
  XNOR U9740 ( .A(n9473), .B(n9465), .Z(n9483) );
  XNOR U9741 ( .A(n9464), .B(n9460), .Z(n9484) );
  XNOR U9742 ( .A(n9459), .B(n9455), .Z(n9485) );
  XNOR U9743 ( .A(n9454), .B(n9450), .Z(n9486) );
  XNOR U9744 ( .A(n9441), .B(n9440), .Z(n9487) );
  XOR U9745 ( .A(n9488), .B(n9439), .Z(n9440) );
  AND U9746 ( .A(b[8]), .B(a[18]), .Z(n9488) );
  XNOR U9747 ( .A(n9439), .B(n9445), .Z(n9489) );
  XNOR U9748 ( .A(n9444), .B(n9436), .Z(n9490) );
  XNOR U9749 ( .A(n9435), .B(n9431), .Z(n9491) );
  XNOR U9750 ( .A(n9430), .B(n9426), .Z(n9492) );
  XNOR U9751 ( .A(n9425), .B(n9421), .Z(n9493) );
  XNOR U9752 ( .A(n9412), .B(n9411), .Z(n9494) );
  XOR U9753 ( .A(n9495), .B(n9410), .Z(n9411) );
  AND U9754 ( .A(b[14]), .B(a[12]), .Z(n9495) );
  XNOR U9755 ( .A(n9410), .B(n9416), .Z(n9496) );
  XNOR U9756 ( .A(n9415), .B(n9407), .Z(n9497) );
  XNOR U9757 ( .A(n9406), .B(n9402), .Z(n9498) );
  XNOR U9758 ( .A(n9401), .B(n9397), .Z(n9499) );
  XNOR U9759 ( .A(n9396), .B(n9392), .Z(n9500) );
  XNOR U9760 ( .A(n9383), .B(n9382), .Z(n9501) );
  XOR U9761 ( .A(n9502), .B(n9381), .Z(n9382) );
  AND U9762 ( .A(a[6]), .B(b[20]), .Z(n9502) );
  XNOR U9763 ( .A(n9381), .B(n9387), .Z(n9503) );
  XNOR U9764 ( .A(n9386), .B(n9378), .Z(n9504) );
  XNOR U9765 ( .A(n9377), .B(n9373), .Z(n9505) );
  XNOR U9766 ( .A(n9372), .B(n9368), .Z(n9506) );
  XNOR U9767 ( .A(n9367), .B(n9363), .Z(n9507) );
  XOR U9768 ( .A(n9508), .B(n9362), .Z(n9363) );
  AND U9769 ( .A(a[0]), .B(b[26]), .Z(n9508) );
  XNOR U9770 ( .A(n9509), .B(n9362), .Z(n9364) );
  XNOR U9771 ( .A(n9510), .B(n9511), .Z(n9362) );
  ANDN U9772 ( .B(n9512), .A(n9513), .Z(n9510) );
  AND U9773 ( .A(a[1]), .B(b[25]), .Z(n9509) );
  XNOR U9774 ( .A(n9514), .B(n9367), .Z(n9369) );
  XOR U9775 ( .A(n9515), .B(n9516), .Z(n9367) );
  ANDN U9776 ( .B(n9517), .A(n9518), .Z(n9515) );
  AND U9777 ( .A(a[2]), .B(b[24]), .Z(n9514) );
  XNOR U9778 ( .A(n9519), .B(n9372), .Z(n9374) );
  XOR U9779 ( .A(n9520), .B(n9521), .Z(n9372) );
  ANDN U9780 ( .B(n9522), .A(n9523), .Z(n9520) );
  AND U9781 ( .A(a[3]), .B(b[23]), .Z(n9519) );
  XNOR U9782 ( .A(n9524), .B(n9377), .Z(n9379) );
  XOR U9783 ( .A(n9525), .B(n9526), .Z(n9377) );
  ANDN U9784 ( .B(n9527), .A(n9528), .Z(n9525) );
  AND U9785 ( .A(a[4]), .B(b[22]), .Z(n9524) );
  XOR U9786 ( .A(n9529), .B(n9530), .Z(n9381) );
  AND U9787 ( .A(n9531), .B(n9532), .Z(n9529) );
  XNOR U9788 ( .A(n9533), .B(n9386), .Z(n9388) );
  XOR U9789 ( .A(n9534), .B(n9535), .Z(n9386) );
  ANDN U9790 ( .B(n9536), .A(n9537), .Z(n9534) );
  AND U9791 ( .A(a[5]), .B(b[21]), .Z(n9533) );
  XOR U9792 ( .A(n9538), .B(n9391), .Z(n9393) );
  XOR U9793 ( .A(n9539), .B(n9540), .Z(n9391) );
  ANDN U9794 ( .B(n9541), .A(n9542), .Z(n9539) );
  AND U9795 ( .A(a[7]), .B(b[19]), .Z(n9538) );
  XNOR U9796 ( .A(n9543), .B(n9396), .Z(n9398) );
  XOR U9797 ( .A(n9544), .B(n9545), .Z(n9396) );
  ANDN U9798 ( .B(n9546), .A(n9547), .Z(n9544) );
  AND U9799 ( .A(a[8]), .B(b[18]), .Z(n9543) );
  XNOR U9800 ( .A(n9548), .B(n9401), .Z(n9403) );
  XOR U9801 ( .A(n9549), .B(n9550), .Z(n9401) );
  ANDN U9802 ( .B(n9551), .A(n9552), .Z(n9549) );
  AND U9803 ( .A(a[9]), .B(b[17]), .Z(n9548) );
  XNOR U9804 ( .A(n9553), .B(n9406), .Z(n9408) );
  XOR U9805 ( .A(n9554), .B(n9555), .Z(n9406) );
  ANDN U9806 ( .B(n9556), .A(n9557), .Z(n9554) );
  AND U9807 ( .A(b[16]), .B(a[10]), .Z(n9553) );
  XOR U9808 ( .A(n9558), .B(n9559), .Z(n9410) );
  AND U9809 ( .A(n9560), .B(n9561), .Z(n9558) );
  XNOR U9810 ( .A(n9562), .B(n9415), .Z(n9417) );
  XOR U9811 ( .A(n9563), .B(n9564), .Z(n9415) );
  ANDN U9812 ( .B(n9565), .A(n9566), .Z(n9563) );
  AND U9813 ( .A(a[11]), .B(b[15]), .Z(n9562) );
  XOR U9814 ( .A(n9567), .B(n9420), .Z(n9422) );
  XOR U9815 ( .A(n9568), .B(n9569), .Z(n9420) );
  ANDN U9816 ( .B(n9570), .A(n9571), .Z(n9568) );
  AND U9817 ( .A(b[13]), .B(a[13]), .Z(n9567) );
  XNOR U9818 ( .A(n9572), .B(n9425), .Z(n9427) );
  XOR U9819 ( .A(n9573), .B(n9574), .Z(n9425) );
  ANDN U9820 ( .B(n9575), .A(n9576), .Z(n9573) );
  AND U9821 ( .A(b[12]), .B(a[14]), .Z(n9572) );
  XNOR U9822 ( .A(n9577), .B(n9430), .Z(n9432) );
  XOR U9823 ( .A(n9578), .B(n9579), .Z(n9430) );
  ANDN U9824 ( .B(n9580), .A(n9581), .Z(n9578) );
  AND U9825 ( .A(b[11]), .B(a[15]), .Z(n9577) );
  XNOR U9826 ( .A(n9582), .B(n9435), .Z(n9437) );
  XOR U9827 ( .A(n9583), .B(n9584), .Z(n9435) );
  ANDN U9828 ( .B(n9585), .A(n9586), .Z(n9583) );
  AND U9829 ( .A(b[10]), .B(a[16]), .Z(n9582) );
  XOR U9830 ( .A(n9587), .B(n9588), .Z(n9439) );
  AND U9831 ( .A(n9589), .B(n9590), .Z(n9587) );
  XNOR U9832 ( .A(n9591), .B(n9444), .Z(n9446) );
  XOR U9833 ( .A(n9592), .B(n9593), .Z(n9444) );
  ANDN U9834 ( .B(n9594), .A(n9595), .Z(n9592) );
  AND U9835 ( .A(b[9]), .B(a[17]), .Z(n9591) );
  XOR U9836 ( .A(n9596), .B(n9449), .Z(n9451) );
  XOR U9837 ( .A(n9597), .B(n9598), .Z(n9449) );
  ANDN U9838 ( .B(n9599), .A(n9600), .Z(n9597) );
  AND U9839 ( .A(b[7]), .B(a[19]), .Z(n9596) );
  XNOR U9840 ( .A(n9601), .B(n9454), .Z(n9456) );
  XOR U9841 ( .A(n9602), .B(n9603), .Z(n9454) );
  ANDN U9842 ( .B(n9604), .A(n9605), .Z(n9602) );
  AND U9843 ( .A(b[6]), .B(a[20]), .Z(n9601) );
  XNOR U9844 ( .A(n9606), .B(n9459), .Z(n9461) );
  XOR U9845 ( .A(n9607), .B(n9608), .Z(n9459) );
  ANDN U9846 ( .B(n9609), .A(n9610), .Z(n9607) );
  AND U9847 ( .A(b[5]), .B(a[21]), .Z(n9606) );
  XNOR U9848 ( .A(n9611), .B(n9464), .Z(n9466) );
  XOR U9849 ( .A(n9612), .B(n9613), .Z(n9464) );
  ANDN U9850 ( .B(n9614), .A(n9615), .Z(n9612) );
  AND U9851 ( .A(b[4]), .B(a[22]), .Z(n9611) );
  XNOR U9852 ( .A(n9616), .B(n9473), .Z(n9475) );
  XNOR U9853 ( .A(n9617), .B(n9618), .Z(n9473) );
  NOR U9854 ( .A(n9619), .B(n9620), .Z(n9617) );
  AND U9855 ( .A(b[3]), .B(a[23]), .Z(n9616) );
  NANDN U9856 ( .A(n9621), .B(n9622), .Z(n9476) );
  XNOR U9857 ( .A(n9623), .B(n9468), .Z(n9470) );
  XNOR U9858 ( .A(n9624), .B(n9625), .Z(n9468) );
  OR U9859 ( .A(n9626), .B(n9627), .Z(n9625) );
  AND U9860 ( .A(b[2]), .B(a[24]), .Z(n9623) );
  NAND U9861 ( .A(a[26]), .B(b[0]), .Z(n9329) );
  XNOR U9862 ( .A(n9621), .B(n9622), .Z(c[25]) );
  XOR U9863 ( .A(n9627), .B(n9626), .Z(n9622) );
  XOR U9864 ( .A(n9624), .B(n9628), .Z(n9626) );
  NAND U9865 ( .A(b[1]), .B(a[24]), .Z(n9628) );
  XOR U9866 ( .A(n9624), .B(n9620), .Z(n9629) );
  XOR U9867 ( .A(n9630), .B(n9618), .Z(n9620) );
  AND U9868 ( .A(b[2]), .B(a[23]), .Z(n9630) );
  ANDN U9869 ( .B(n9631), .A(n9632), .Z(n9624) );
  XOR U9870 ( .A(n9618), .B(n9614), .Z(n9633) );
  XNOR U9871 ( .A(n9613), .B(n9609), .Z(n9634) );
  XNOR U9872 ( .A(n9608), .B(n9604), .Z(n9635) );
  XNOR U9873 ( .A(n9603), .B(n9599), .Z(n9636) );
  XNOR U9874 ( .A(n9590), .B(n9589), .Z(n9637) );
  XOR U9875 ( .A(n9638), .B(n9588), .Z(n9589) );
  AND U9876 ( .A(b[7]), .B(a[18]), .Z(n9638) );
  XNOR U9877 ( .A(n9588), .B(n9594), .Z(n9639) );
  XNOR U9878 ( .A(n9593), .B(n9585), .Z(n9640) );
  XNOR U9879 ( .A(n9584), .B(n9580), .Z(n9641) );
  XNOR U9880 ( .A(n9579), .B(n9575), .Z(n9642) );
  XNOR U9881 ( .A(n9574), .B(n9570), .Z(n9643) );
  XNOR U9882 ( .A(n9561), .B(n9560), .Z(n9644) );
  XOR U9883 ( .A(n9645), .B(n9559), .Z(n9560) );
  AND U9884 ( .A(b[13]), .B(a[12]), .Z(n9645) );
  XNOR U9885 ( .A(n9559), .B(n9565), .Z(n9646) );
  XNOR U9886 ( .A(n9564), .B(n9556), .Z(n9647) );
  XNOR U9887 ( .A(n9555), .B(n9551), .Z(n9648) );
  XNOR U9888 ( .A(n9550), .B(n9546), .Z(n9649) );
  XNOR U9889 ( .A(n9545), .B(n9541), .Z(n9650) );
  XNOR U9890 ( .A(n9532), .B(n9531), .Z(n9651) );
  XOR U9891 ( .A(n9652), .B(n9530), .Z(n9531) );
  AND U9892 ( .A(a[6]), .B(b[19]), .Z(n9652) );
  XNOR U9893 ( .A(n9530), .B(n9536), .Z(n9653) );
  XNOR U9894 ( .A(n9535), .B(n9527), .Z(n9654) );
  XNOR U9895 ( .A(n9526), .B(n9522), .Z(n9655) );
  XNOR U9896 ( .A(n9521), .B(n9517), .Z(n9656) );
  XNOR U9897 ( .A(n9516), .B(n9512), .Z(n9657) );
  XNOR U9898 ( .A(n9658), .B(n9511), .Z(n9512) );
  AND U9899 ( .A(a[0]), .B(b[25]), .Z(n9658) );
  XOR U9900 ( .A(n9659), .B(n9511), .Z(n9513) );
  XNOR U9901 ( .A(n9660), .B(n9661), .Z(n9511) );
  ANDN U9902 ( .B(n9662), .A(n9663), .Z(n9660) );
  AND U9903 ( .A(a[1]), .B(b[24]), .Z(n9659) );
  XNOR U9904 ( .A(n9664), .B(n9516), .Z(n9518) );
  XOR U9905 ( .A(n9665), .B(n9666), .Z(n9516) );
  ANDN U9906 ( .B(n9667), .A(n9668), .Z(n9665) );
  AND U9907 ( .A(a[2]), .B(b[23]), .Z(n9664) );
  XNOR U9908 ( .A(n9669), .B(n9521), .Z(n9523) );
  XOR U9909 ( .A(n9670), .B(n9671), .Z(n9521) );
  ANDN U9910 ( .B(n9672), .A(n9673), .Z(n9670) );
  AND U9911 ( .A(a[3]), .B(b[22]), .Z(n9669) );
  XNOR U9912 ( .A(n9674), .B(n9526), .Z(n9528) );
  XOR U9913 ( .A(n9675), .B(n9676), .Z(n9526) );
  ANDN U9914 ( .B(n9677), .A(n9678), .Z(n9675) );
  AND U9915 ( .A(a[4]), .B(b[21]), .Z(n9674) );
  XOR U9916 ( .A(n9679), .B(n9680), .Z(n9530) );
  AND U9917 ( .A(n9681), .B(n9682), .Z(n9679) );
  XNOR U9918 ( .A(n9683), .B(n9535), .Z(n9537) );
  XOR U9919 ( .A(n9684), .B(n9685), .Z(n9535) );
  ANDN U9920 ( .B(n9686), .A(n9687), .Z(n9684) );
  AND U9921 ( .A(a[5]), .B(b[20]), .Z(n9683) );
  XOR U9922 ( .A(n9688), .B(n9540), .Z(n9542) );
  XOR U9923 ( .A(n9689), .B(n9690), .Z(n9540) );
  ANDN U9924 ( .B(n9691), .A(n9692), .Z(n9689) );
  AND U9925 ( .A(a[7]), .B(b[18]), .Z(n9688) );
  XNOR U9926 ( .A(n9693), .B(n9545), .Z(n9547) );
  XOR U9927 ( .A(n9694), .B(n9695), .Z(n9545) );
  ANDN U9928 ( .B(n9696), .A(n9697), .Z(n9694) );
  AND U9929 ( .A(a[8]), .B(b[17]), .Z(n9693) );
  XNOR U9930 ( .A(n9698), .B(n9550), .Z(n9552) );
  XOR U9931 ( .A(n9699), .B(n9700), .Z(n9550) );
  ANDN U9932 ( .B(n9701), .A(n9702), .Z(n9699) );
  AND U9933 ( .A(a[9]), .B(b[16]), .Z(n9698) );
  XNOR U9934 ( .A(n9703), .B(n9555), .Z(n9557) );
  XOR U9935 ( .A(n9704), .B(n9705), .Z(n9555) );
  ANDN U9936 ( .B(n9706), .A(n9707), .Z(n9704) );
  AND U9937 ( .A(a[10]), .B(b[15]), .Z(n9703) );
  XOR U9938 ( .A(n9708), .B(n9709), .Z(n9559) );
  AND U9939 ( .A(n9710), .B(n9711), .Z(n9708) );
  XNOR U9940 ( .A(n9712), .B(n9564), .Z(n9566) );
  XOR U9941 ( .A(n9713), .B(n9714), .Z(n9564) );
  ANDN U9942 ( .B(n9715), .A(n9716), .Z(n9713) );
  AND U9943 ( .A(b[14]), .B(a[11]), .Z(n9712) );
  XOR U9944 ( .A(n9717), .B(n9569), .Z(n9571) );
  XOR U9945 ( .A(n9718), .B(n9719), .Z(n9569) );
  ANDN U9946 ( .B(n9720), .A(n9721), .Z(n9718) );
  AND U9947 ( .A(b[12]), .B(a[13]), .Z(n9717) );
  XNOR U9948 ( .A(n9722), .B(n9574), .Z(n9576) );
  XOR U9949 ( .A(n9723), .B(n9724), .Z(n9574) );
  ANDN U9950 ( .B(n9725), .A(n9726), .Z(n9723) );
  AND U9951 ( .A(b[11]), .B(a[14]), .Z(n9722) );
  XNOR U9952 ( .A(n9727), .B(n9579), .Z(n9581) );
  XOR U9953 ( .A(n9728), .B(n9729), .Z(n9579) );
  ANDN U9954 ( .B(n9730), .A(n9731), .Z(n9728) );
  AND U9955 ( .A(b[10]), .B(a[15]), .Z(n9727) );
  XNOR U9956 ( .A(n9732), .B(n9584), .Z(n9586) );
  XOR U9957 ( .A(n9733), .B(n9734), .Z(n9584) );
  ANDN U9958 ( .B(n9735), .A(n9736), .Z(n9733) );
  AND U9959 ( .A(b[9]), .B(a[16]), .Z(n9732) );
  XOR U9960 ( .A(n9737), .B(n9738), .Z(n9588) );
  AND U9961 ( .A(n9739), .B(n9740), .Z(n9737) );
  XNOR U9962 ( .A(n9741), .B(n9593), .Z(n9595) );
  XOR U9963 ( .A(n9742), .B(n9743), .Z(n9593) );
  ANDN U9964 ( .B(n9744), .A(n9745), .Z(n9742) );
  AND U9965 ( .A(b[8]), .B(a[17]), .Z(n9741) );
  XOR U9966 ( .A(n9746), .B(n9598), .Z(n9600) );
  XOR U9967 ( .A(n9747), .B(n9748), .Z(n9598) );
  ANDN U9968 ( .B(n9749), .A(n9750), .Z(n9747) );
  AND U9969 ( .A(b[6]), .B(a[19]), .Z(n9746) );
  XNOR U9970 ( .A(n9751), .B(n9603), .Z(n9605) );
  XOR U9971 ( .A(n9752), .B(n9753), .Z(n9603) );
  ANDN U9972 ( .B(n9754), .A(n9755), .Z(n9752) );
  AND U9973 ( .A(b[5]), .B(a[20]), .Z(n9751) );
  XNOR U9974 ( .A(n9756), .B(n9608), .Z(n9610) );
  XOR U9975 ( .A(n9757), .B(n9758), .Z(n9608) );
  ANDN U9976 ( .B(n9759), .A(n9760), .Z(n9757) );
  AND U9977 ( .A(b[4]), .B(a[21]), .Z(n9756) );
  XNOR U9978 ( .A(n9761), .B(n9762), .Z(n9618) );
  NANDN U9979 ( .A(n9763), .B(n9764), .Z(n9762) );
  XNOR U9980 ( .A(n9765), .B(n9613), .Z(n9615) );
  XNOR U9981 ( .A(n9766), .B(n9767), .Z(n9613) );
  AND U9982 ( .A(n9768), .B(n9769), .Z(n9766) );
  AND U9983 ( .A(b[3]), .B(a[22]), .Z(n9765) );
  NAND U9984 ( .A(a[25]), .B(b[0]), .Z(n9621) );
  XNOR U9985 ( .A(n9632), .B(n9631), .Z(c[24]) );
  XNOR U9986 ( .A(n9763), .B(n9764), .Z(n9631) );
  XOR U9987 ( .A(n9761), .B(n9770), .Z(n9764) );
  NAND U9988 ( .A(b[1]), .B(a[23]), .Z(n9770) );
  XOR U9989 ( .A(n9769), .B(n9771), .Z(n9763) );
  XOR U9990 ( .A(n9761), .B(n9768), .Z(n9771) );
  XNOR U9991 ( .A(n9772), .B(n9767), .Z(n9768) );
  AND U9992 ( .A(b[2]), .B(a[22]), .Z(n9772) );
  NANDN U9993 ( .A(n9773), .B(n9774), .Z(n9761) );
  XOR U9994 ( .A(n9767), .B(n9759), .Z(n9775) );
  XNOR U9995 ( .A(n9758), .B(n9754), .Z(n9776) );
  XNOR U9996 ( .A(n9753), .B(n9749), .Z(n9777) );
  XNOR U9997 ( .A(n9740), .B(n9739), .Z(n9778) );
  XOR U9998 ( .A(n9779), .B(n9738), .Z(n9739) );
  AND U9999 ( .A(b[6]), .B(a[18]), .Z(n9779) );
  XNOR U10000 ( .A(n9738), .B(n9744), .Z(n9780) );
  XNOR U10001 ( .A(n9743), .B(n9735), .Z(n9781) );
  XNOR U10002 ( .A(n9734), .B(n9730), .Z(n9782) );
  XNOR U10003 ( .A(n9729), .B(n9725), .Z(n9783) );
  XNOR U10004 ( .A(n9724), .B(n9720), .Z(n9784) );
  XNOR U10005 ( .A(n9711), .B(n9710), .Z(n9785) );
  XOR U10006 ( .A(n9786), .B(n9709), .Z(n9710) );
  AND U10007 ( .A(b[12]), .B(a[12]), .Z(n9786) );
  XNOR U10008 ( .A(n9709), .B(n9715), .Z(n9787) );
  XNOR U10009 ( .A(n9714), .B(n9706), .Z(n9788) );
  XNOR U10010 ( .A(n9705), .B(n9701), .Z(n9789) );
  XNOR U10011 ( .A(n9700), .B(n9696), .Z(n9790) );
  XNOR U10012 ( .A(n9695), .B(n9691), .Z(n9791) );
  XNOR U10013 ( .A(n9682), .B(n9681), .Z(n9792) );
  XOR U10014 ( .A(n9793), .B(n9680), .Z(n9681) );
  AND U10015 ( .A(a[6]), .B(b[18]), .Z(n9793) );
  XNOR U10016 ( .A(n9680), .B(n9686), .Z(n9794) );
  XNOR U10017 ( .A(n9685), .B(n9677), .Z(n9795) );
  XNOR U10018 ( .A(n9676), .B(n9672), .Z(n9796) );
  XNOR U10019 ( .A(n9671), .B(n9667), .Z(n9797) );
  XNOR U10020 ( .A(n9666), .B(n9662), .Z(n9798) );
  XOR U10021 ( .A(n9799), .B(n9661), .Z(n9662) );
  AND U10022 ( .A(a[0]), .B(b[24]), .Z(n9799) );
  XNOR U10023 ( .A(n9800), .B(n9661), .Z(n9663) );
  XNOR U10024 ( .A(n9801), .B(n9802), .Z(n9661) );
  ANDN U10025 ( .B(n9803), .A(n9804), .Z(n9801) );
  AND U10026 ( .A(a[1]), .B(b[23]), .Z(n9800) );
  XNOR U10027 ( .A(n9805), .B(n9666), .Z(n9668) );
  XOR U10028 ( .A(n9806), .B(n9807), .Z(n9666) );
  ANDN U10029 ( .B(n9808), .A(n9809), .Z(n9806) );
  AND U10030 ( .A(a[2]), .B(b[22]), .Z(n9805) );
  XNOR U10031 ( .A(n9810), .B(n9671), .Z(n9673) );
  XOR U10032 ( .A(n9811), .B(n9812), .Z(n9671) );
  ANDN U10033 ( .B(n9813), .A(n9814), .Z(n9811) );
  AND U10034 ( .A(a[3]), .B(b[21]), .Z(n9810) );
  XNOR U10035 ( .A(n9815), .B(n9676), .Z(n9678) );
  XOR U10036 ( .A(n9816), .B(n9817), .Z(n9676) );
  ANDN U10037 ( .B(n9818), .A(n9819), .Z(n9816) );
  AND U10038 ( .A(a[4]), .B(b[20]), .Z(n9815) );
  XOR U10039 ( .A(n9820), .B(n9821), .Z(n9680) );
  AND U10040 ( .A(n9822), .B(n9823), .Z(n9820) );
  XNOR U10041 ( .A(n9824), .B(n9685), .Z(n9687) );
  XOR U10042 ( .A(n9825), .B(n9826), .Z(n9685) );
  ANDN U10043 ( .B(n9827), .A(n9828), .Z(n9825) );
  AND U10044 ( .A(a[5]), .B(b[19]), .Z(n9824) );
  XOR U10045 ( .A(n9829), .B(n9690), .Z(n9692) );
  XOR U10046 ( .A(n9830), .B(n9831), .Z(n9690) );
  ANDN U10047 ( .B(n9832), .A(n9833), .Z(n9830) );
  AND U10048 ( .A(a[7]), .B(b[17]), .Z(n9829) );
  XNOR U10049 ( .A(n9834), .B(n9695), .Z(n9697) );
  XOR U10050 ( .A(n9835), .B(n9836), .Z(n9695) );
  ANDN U10051 ( .B(n9837), .A(n9838), .Z(n9835) );
  AND U10052 ( .A(a[8]), .B(b[16]), .Z(n9834) );
  XNOR U10053 ( .A(n9839), .B(n9700), .Z(n9702) );
  XOR U10054 ( .A(n9840), .B(n9841), .Z(n9700) );
  ANDN U10055 ( .B(n9842), .A(n9843), .Z(n9840) );
  AND U10056 ( .A(a[9]), .B(b[15]), .Z(n9839) );
  XNOR U10057 ( .A(n9844), .B(n9705), .Z(n9707) );
  XOR U10058 ( .A(n9845), .B(n9846), .Z(n9705) );
  ANDN U10059 ( .B(n9847), .A(n9848), .Z(n9845) );
  AND U10060 ( .A(b[14]), .B(a[10]), .Z(n9844) );
  XOR U10061 ( .A(n9849), .B(n9850), .Z(n9709) );
  AND U10062 ( .A(n9851), .B(n9852), .Z(n9849) );
  XNOR U10063 ( .A(n9853), .B(n9714), .Z(n9716) );
  XOR U10064 ( .A(n9854), .B(n9855), .Z(n9714) );
  ANDN U10065 ( .B(n9856), .A(n9857), .Z(n9854) );
  AND U10066 ( .A(b[13]), .B(a[11]), .Z(n9853) );
  XOR U10067 ( .A(n9858), .B(n9719), .Z(n9721) );
  XOR U10068 ( .A(n9859), .B(n9860), .Z(n9719) );
  ANDN U10069 ( .B(n9861), .A(n9862), .Z(n9859) );
  AND U10070 ( .A(b[11]), .B(a[13]), .Z(n9858) );
  XNOR U10071 ( .A(n9863), .B(n9724), .Z(n9726) );
  XOR U10072 ( .A(n9864), .B(n9865), .Z(n9724) );
  ANDN U10073 ( .B(n9866), .A(n9867), .Z(n9864) );
  AND U10074 ( .A(b[10]), .B(a[14]), .Z(n9863) );
  XNOR U10075 ( .A(n9868), .B(n9729), .Z(n9731) );
  XOR U10076 ( .A(n9869), .B(n9870), .Z(n9729) );
  ANDN U10077 ( .B(n9871), .A(n9872), .Z(n9869) );
  AND U10078 ( .A(b[9]), .B(a[15]), .Z(n9868) );
  XNOR U10079 ( .A(n9873), .B(n9734), .Z(n9736) );
  XOR U10080 ( .A(n9874), .B(n9875), .Z(n9734) );
  ANDN U10081 ( .B(n9876), .A(n9877), .Z(n9874) );
  AND U10082 ( .A(b[8]), .B(a[16]), .Z(n9873) );
  XOR U10083 ( .A(n9878), .B(n9879), .Z(n9738) );
  AND U10084 ( .A(n9880), .B(n9881), .Z(n9878) );
  XNOR U10085 ( .A(n9882), .B(n9743), .Z(n9745) );
  XOR U10086 ( .A(n9883), .B(n9884), .Z(n9743) );
  ANDN U10087 ( .B(n9885), .A(n9886), .Z(n9883) );
  AND U10088 ( .A(b[7]), .B(a[17]), .Z(n9882) );
  XOR U10089 ( .A(n9887), .B(n9748), .Z(n9750) );
  XOR U10090 ( .A(n9888), .B(n9889), .Z(n9748) );
  ANDN U10091 ( .B(n9890), .A(n9891), .Z(n9888) );
  AND U10092 ( .A(b[5]), .B(a[19]), .Z(n9887) );
  XNOR U10093 ( .A(n9892), .B(n9753), .Z(n9755) );
  XOR U10094 ( .A(n9893), .B(n9894), .Z(n9753) );
  ANDN U10095 ( .B(n9895), .A(n9896), .Z(n9893) );
  AND U10096 ( .A(b[4]), .B(a[20]), .Z(n9892) );
  XNOR U10097 ( .A(n9897), .B(n9898), .Z(n9767) );
  NANDN U10098 ( .A(n9899), .B(n9900), .Z(n9898) );
  XNOR U10099 ( .A(n9901), .B(n9758), .Z(n9760) );
  XNOR U10100 ( .A(n9902), .B(n9903), .Z(n9758) );
  AND U10101 ( .A(n9904), .B(n9905), .Z(n9902) );
  AND U10102 ( .A(b[3]), .B(a[21]), .Z(n9901) );
  NAND U10103 ( .A(a[24]), .B(b[0]), .Z(n9632) );
  XNOR U10104 ( .A(n9773), .B(n9774), .Z(c[23]) );
  XNOR U10105 ( .A(n9899), .B(n9900), .Z(n9774) );
  XOR U10106 ( .A(n9897), .B(n9906), .Z(n9900) );
  NAND U10107 ( .A(b[1]), .B(a[22]), .Z(n9906) );
  XOR U10108 ( .A(n9905), .B(n9907), .Z(n9899) );
  XOR U10109 ( .A(n9897), .B(n9904), .Z(n9907) );
  XNOR U10110 ( .A(n9908), .B(n9903), .Z(n9904) );
  AND U10111 ( .A(b[2]), .B(a[21]), .Z(n9908) );
  NANDN U10112 ( .A(n9909), .B(n9910), .Z(n9897) );
  XOR U10113 ( .A(n9903), .B(n9895), .Z(n9911) );
  XNOR U10114 ( .A(n9894), .B(n9890), .Z(n9912) );
  XNOR U10115 ( .A(n9881), .B(n9880), .Z(n9913) );
  XOR U10116 ( .A(n9914), .B(n9879), .Z(n9880) );
  AND U10117 ( .A(b[5]), .B(a[18]), .Z(n9914) );
  XNOR U10118 ( .A(n9879), .B(n9885), .Z(n9915) );
  XNOR U10119 ( .A(n9884), .B(n9876), .Z(n9916) );
  XNOR U10120 ( .A(n9875), .B(n9871), .Z(n9917) );
  XNOR U10121 ( .A(n9870), .B(n9866), .Z(n9918) );
  XNOR U10122 ( .A(n9865), .B(n9861), .Z(n9919) );
  XNOR U10123 ( .A(n9852), .B(n9851), .Z(n9920) );
  XOR U10124 ( .A(n9921), .B(n9850), .Z(n9851) );
  AND U10125 ( .A(b[11]), .B(a[12]), .Z(n9921) );
  XNOR U10126 ( .A(n9850), .B(n9856), .Z(n9922) );
  XNOR U10127 ( .A(n9855), .B(n9847), .Z(n9923) );
  XNOR U10128 ( .A(n9846), .B(n9842), .Z(n9924) );
  XNOR U10129 ( .A(n9841), .B(n9837), .Z(n9925) );
  XNOR U10130 ( .A(n9836), .B(n9832), .Z(n9926) );
  XNOR U10131 ( .A(n9823), .B(n9822), .Z(n9927) );
  XOR U10132 ( .A(n9928), .B(n9821), .Z(n9822) );
  AND U10133 ( .A(a[6]), .B(b[17]), .Z(n9928) );
  XNOR U10134 ( .A(n9821), .B(n9827), .Z(n9929) );
  XNOR U10135 ( .A(n9826), .B(n9818), .Z(n9930) );
  XNOR U10136 ( .A(n9817), .B(n9813), .Z(n9931) );
  XNOR U10137 ( .A(n9812), .B(n9808), .Z(n9932) );
  XNOR U10138 ( .A(n9807), .B(n9803), .Z(n9933) );
  XNOR U10139 ( .A(n9934), .B(n9802), .Z(n9803) );
  AND U10140 ( .A(a[0]), .B(b[23]), .Z(n9934) );
  XOR U10141 ( .A(n9935), .B(n9802), .Z(n9804) );
  XNOR U10142 ( .A(n9936), .B(n9937), .Z(n9802) );
  ANDN U10143 ( .B(n9938), .A(n9939), .Z(n9936) );
  AND U10144 ( .A(a[1]), .B(b[22]), .Z(n9935) );
  XNOR U10145 ( .A(n9940), .B(n9807), .Z(n9809) );
  XOR U10146 ( .A(n9941), .B(n9942), .Z(n9807) );
  ANDN U10147 ( .B(n9943), .A(n9944), .Z(n9941) );
  AND U10148 ( .A(a[2]), .B(b[21]), .Z(n9940) );
  XNOR U10149 ( .A(n9945), .B(n9812), .Z(n9814) );
  XOR U10150 ( .A(n9946), .B(n9947), .Z(n9812) );
  ANDN U10151 ( .B(n9948), .A(n9949), .Z(n9946) );
  AND U10152 ( .A(a[3]), .B(b[20]), .Z(n9945) );
  XNOR U10153 ( .A(n9950), .B(n9817), .Z(n9819) );
  XOR U10154 ( .A(n9951), .B(n9952), .Z(n9817) );
  ANDN U10155 ( .B(n9953), .A(n9954), .Z(n9951) );
  AND U10156 ( .A(a[4]), .B(b[19]), .Z(n9950) );
  XOR U10157 ( .A(n9955), .B(n9956), .Z(n9821) );
  AND U10158 ( .A(n9957), .B(n9958), .Z(n9955) );
  XNOR U10159 ( .A(n9959), .B(n9826), .Z(n9828) );
  XOR U10160 ( .A(n9960), .B(n9961), .Z(n9826) );
  ANDN U10161 ( .B(n9962), .A(n9963), .Z(n9960) );
  AND U10162 ( .A(a[5]), .B(b[18]), .Z(n9959) );
  XOR U10163 ( .A(n9964), .B(n9831), .Z(n9833) );
  XOR U10164 ( .A(n9965), .B(n9966), .Z(n9831) );
  ANDN U10165 ( .B(n9967), .A(n9968), .Z(n9965) );
  AND U10166 ( .A(a[7]), .B(b[16]), .Z(n9964) );
  XNOR U10167 ( .A(n9969), .B(n9836), .Z(n9838) );
  XOR U10168 ( .A(n9970), .B(n9971), .Z(n9836) );
  ANDN U10169 ( .B(n9972), .A(n9973), .Z(n9970) );
  AND U10170 ( .A(a[8]), .B(b[15]), .Z(n9969) );
  XNOR U10171 ( .A(n9974), .B(n9841), .Z(n9843) );
  XOR U10172 ( .A(n9975), .B(n9976), .Z(n9841) );
  ANDN U10173 ( .B(n9977), .A(n9978), .Z(n9975) );
  AND U10174 ( .A(a[9]), .B(b[14]), .Z(n9974) );
  XNOR U10175 ( .A(n9979), .B(n9846), .Z(n9848) );
  XOR U10176 ( .A(n9980), .B(n9981), .Z(n9846) );
  ANDN U10177 ( .B(n9982), .A(n9983), .Z(n9980) );
  AND U10178 ( .A(b[13]), .B(a[10]), .Z(n9979) );
  XOR U10179 ( .A(n9984), .B(n9985), .Z(n9850) );
  AND U10180 ( .A(n9986), .B(n9987), .Z(n9984) );
  XNOR U10181 ( .A(n9988), .B(n9855), .Z(n9857) );
  XOR U10182 ( .A(n9989), .B(n9990), .Z(n9855) );
  ANDN U10183 ( .B(n9991), .A(n9992), .Z(n9989) );
  AND U10184 ( .A(b[12]), .B(a[11]), .Z(n9988) );
  XOR U10185 ( .A(n9993), .B(n9860), .Z(n9862) );
  XOR U10186 ( .A(n9994), .B(n9995), .Z(n9860) );
  ANDN U10187 ( .B(n9996), .A(n9997), .Z(n9994) );
  AND U10188 ( .A(b[10]), .B(a[13]), .Z(n9993) );
  XNOR U10189 ( .A(n9998), .B(n9865), .Z(n9867) );
  XOR U10190 ( .A(n9999), .B(n10000), .Z(n9865) );
  ANDN U10191 ( .B(n10001), .A(n10002), .Z(n9999) );
  AND U10192 ( .A(b[9]), .B(a[14]), .Z(n9998) );
  XNOR U10193 ( .A(n10003), .B(n9870), .Z(n9872) );
  XOR U10194 ( .A(n10004), .B(n10005), .Z(n9870) );
  ANDN U10195 ( .B(n10006), .A(n10007), .Z(n10004) );
  AND U10196 ( .A(b[8]), .B(a[15]), .Z(n10003) );
  XNOR U10197 ( .A(n10008), .B(n9875), .Z(n9877) );
  XOR U10198 ( .A(n10009), .B(n10010), .Z(n9875) );
  ANDN U10199 ( .B(n10011), .A(n10012), .Z(n10009) );
  AND U10200 ( .A(b[7]), .B(a[16]), .Z(n10008) );
  XOR U10201 ( .A(n10013), .B(n10014), .Z(n9879) );
  AND U10202 ( .A(n10015), .B(n10016), .Z(n10013) );
  XNOR U10203 ( .A(n10017), .B(n9884), .Z(n9886) );
  XOR U10204 ( .A(n10018), .B(n10019), .Z(n9884) );
  ANDN U10205 ( .B(n10020), .A(n10021), .Z(n10018) );
  AND U10206 ( .A(b[6]), .B(a[17]), .Z(n10017) );
  XOR U10207 ( .A(n10022), .B(n9889), .Z(n9891) );
  XOR U10208 ( .A(n10023), .B(n10024), .Z(n9889) );
  ANDN U10209 ( .B(n10025), .A(n10026), .Z(n10023) );
  AND U10210 ( .A(b[4]), .B(a[19]), .Z(n10022) );
  XNOR U10211 ( .A(n10027), .B(n10028), .Z(n9903) );
  NANDN U10212 ( .A(n10029), .B(n10030), .Z(n10028) );
  XNOR U10213 ( .A(n10031), .B(n9894), .Z(n9896) );
  XNOR U10214 ( .A(n10032), .B(n10033), .Z(n9894) );
  AND U10215 ( .A(n10034), .B(n10035), .Z(n10032) );
  AND U10216 ( .A(b[3]), .B(a[20]), .Z(n10031) );
  NAND U10217 ( .A(a[23]), .B(b[0]), .Z(n9773) );
  XNOR U10218 ( .A(n9909), .B(n9910), .Z(c[22]) );
  XNOR U10219 ( .A(n10029), .B(n10030), .Z(n9910) );
  XOR U10220 ( .A(n10027), .B(n10036), .Z(n10030) );
  NAND U10221 ( .A(b[1]), .B(a[21]), .Z(n10036) );
  XOR U10222 ( .A(n10035), .B(n10037), .Z(n10029) );
  XOR U10223 ( .A(n10027), .B(n10034), .Z(n10037) );
  XNOR U10224 ( .A(n10038), .B(n10033), .Z(n10034) );
  AND U10225 ( .A(b[2]), .B(a[20]), .Z(n10038) );
  NANDN U10226 ( .A(n10039), .B(n10040), .Z(n10027) );
  XOR U10227 ( .A(n10033), .B(n10025), .Z(n10041) );
  XNOR U10228 ( .A(n10016), .B(n10015), .Z(n10042) );
  XOR U10229 ( .A(n10043), .B(n10014), .Z(n10015) );
  AND U10230 ( .A(b[4]), .B(a[18]), .Z(n10043) );
  XNOR U10231 ( .A(n10014), .B(n10020), .Z(n10044) );
  XNOR U10232 ( .A(n10019), .B(n10011), .Z(n10045) );
  XNOR U10233 ( .A(n10010), .B(n10006), .Z(n10046) );
  XNOR U10234 ( .A(n10005), .B(n10001), .Z(n10047) );
  XNOR U10235 ( .A(n10000), .B(n9996), .Z(n10048) );
  XNOR U10236 ( .A(n9987), .B(n9986), .Z(n10049) );
  XOR U10237 ( .A(n10050), .B(n9985), .Z(n9986) );
  AND U10238 ( .A(b[10]), .B(a[12]), .Z(n10050) );
  XNOR U10239 ( .A(n9985), .B(n9991), .Z(n10051) );
  XNOR U10240 ( .A(n9990), .B(n9982), .Z(n10052) );
  XNOR U10241 ( .A(n9981), .B(n9977), .Z(n10053) );
  XNOR U10242 ( .A(n9976), .B(n9972), .Z(n10054) );
  XNOR U10243 ( .A(n9971), .B(n9967), .Z(n10055) );
  XNOR U10244 ( .A(n9958), .B(n9957), .Z(n10056) );
  XOR U10245 ( .A(n10057), .B(n9956), .Z(n9957) );
  AND U10246 ( .A(a[6]), .B(b[16]), .Z(n10057) );
  XNOR U10247 ( .A(n9956), .B(n9962), .Z(n10058) );
  XNOR U10248 ( .A(n9961), .B(n9953), .Z(n10059) );
  XNOR U10249 ( .A(n9952), .B(n9948), .Z(n10060) );
  XNOR U10250 ( .A(n9947), .B(n9943), .Z(n10061) );
  XNOR U10251 ( .A(n9942), .B(n9938), .Z(n10062) );
  XOR U10252 ( .A(n10063), .B(n9937), .Z(n9938) );
  AND U10253 ( .A(a[0]), .B(b[22]), .Z(n10063) );
  XNOR U10254 ( .A(n10064), .B(n9937), .Z(n9939) );
  XNOR U10255 ( .A(n10065), .B(n10066), .Z(n9937) );
  ANDN U10256 ( .B(n10067), .A(n10068), .Z(n10065) );
  AND U10257 ( .A(a[1]), .B(b[21]), .Z(n10064) );
  XNOR U10258 ( .A(n10069), .B(n9942), .Z(n9944) );
  XOR U10259 ( .A(n10070), .B(n10071), .Z(n9942) );
  ANDN U10260 ( .B(n10072), .A(n10073), .Z(n10070) );
  AND U10261 ( .A(a[2]), .B(b[20]), .Z(n10069) );
  XNOR U10262 ( .A(n10074), .B(n9947), .Z(n9949) );
  XOR U10263 ( .A(n10075), .B(n10076), .Z(n9947) );
  ANDN U10264 ( .B(n10077), .A(n10078), .Z(n10075) );
  AND U10265 ( .A(a[3]), .B(b[19]), .Z(n10074) );
  XNOR U10266 ( .A(n10079), .B(n9952), .Z(n9954) );
  XOR U10267 ( .A(n10080), .B(n10081), .Z(n9952) );
  ANDN U10268 ( .B(n10082), .A(n10083), .Z(n10080) );
  AND U10269 ( .A(a[4]), .B(b[18]), .Z(n10079) );
  XOR U10270 ( .A(n10084), .B(n10085), .Z(n9956) );
  AND U10271 ( .A(n10086), .B(n10087), .Z(n10084) );
  XNOR U10272 ( .A(n10088), .B(n9961), .Z(n9963) );
  XOR U10273 ( .A(n10089), .B(n10090), .Z(n9961) );
  ANDN U10274 ( .B(n10091), .A(n10092), .Z(n10089) );
  AND U10275 ( .A(a[5]), .B(b[17]), .Z(n10088) );
  XOR U10276 ( .A(n10093), .B(n9966), .Z(n9968) );
  XOR U10277 ( .A(n10094), .B(n10095), .Z(n9966) );
  ANDN U10278 ( .B(n10096), .A(n10097), .Z(n10094) );
  AND U10279 ( .A(a[7]), .B(b[15]), .Z(n10093) );
  XNOR U10280 ( .A(n10098), .B(n9971), .Z(n9973) );
  XOR U10281 ( .A(n10099), .B(n10100), .Z(n9971) );
  ANDN U10282 ( .B(n10101), .A(n10102), .Z(n10099) );
  AND U10283 ( .A(a[8]), .B(b[14]), .Z(n10098) );
  XNOR U10284 ( .A(n10103), .B(n9976), .Z(n9978) );
  XOR U10285 ( .A(n10104), .B(n10105), .Z(n9976) );
  ANDN U10286 ( .B(n10106), .A(n10107), .Z(n10104) );
  AND U10287 ( .A(a[9]), .B(b[13]), .Z(n10103) );
  XNOR U10288 ( .A(n10108), .B(n9981), .Z(n9983) );
  XOR U10289 ( .A(n10109), .B(n10110), .Z(n9981) );
  ANDN U10290 ( .B(n10111), .A(n10112), .Z(n10109) );
  AND U10291 ( .A(b[12]), .B(a[10]), .Z(n10108) );
  XOR U10292 ( .A(n10113), .B(n10114), .Z(n9985) );
  AND U10293 ( .A(n10115), .B(n10116), .Z(n10113) );
  XNOR U10294 ( .A(n10117), .B(n9990), .Z(n9992) );
  XOR U10295 ( .A(n10118), .B(n10119), .Z(n9990) );
  ANDN U10296 ( .B(n10120), .A(n10121), .Z(n10118) );
  AND U10297 ( .A(b[11]), .B(a[11]), .Z(n10117) );
  XOR U10298 ( .A(n10122), .B(n9995), .Z(n9997) );
  XOR U10299 ( .A(n10123), .B(n10124), .Z(n9995) );
  ANDN U10300 ( .B(n10125), .A(n10126), .Z(n10123) );
  AND U10301 ( .A(b[9]), .B(a[13]), .Z(n10122) );
  XNOR U10302 ( .A(n10127), .B(n10000), .Z(n10002) );
  XOR U10303 ( .A(n10128), .B(n10129), .Z(n10000) );
  ANDN U10304 ( .B(n10130), .A(n10131), .Z(n10128) );
  AND U10305 ( .A(b[8]), .B(a[14]), .Z(n10127) );
  XNOR U10306 ( .A(n10132), .B(n10005), .Z(n10007) );
  XOR U10307 ( .A(n10133), .B(n10134), .Z(n10005) );
  ANDN U10308 ( .B(n10135), .A(n10136), .Z(n10133) );
  AND U10309 ( .A(b[7]), .B(a[15]), .Z(n10132) );
  XNOR U10310 ( .A(n10137), .B(n10010), .Z(n10012) );
  XOR U10311 ( .A(n10138), .B(n10139), .Z(n10010) );
  ANDN U10312 ( .B(n10140), .A(n10141), .Z(n10138) );
  AND U10313 ( .A(b[6]), .B(a[16]), .Z(n10137) );
  XOR U10314 ( .A(n10142), .B(n10143), .Z(n10014) );
  AND U10315 ( .A(n10144), .B(n10145), .Z(n10142) );
  XNOR U10316 ( .A(n10146), .B(n10019), .Z(n10021) );
  XOR U10317 ( .A(n10147), .B(n10148), .Z(n10019) );
  ANDN U10318 ( .B(n10149), .A(n10150), .Z(n10147) );
  AND U10319 ( .A(b[5]), .B(a[17]), .Z(n10146) );
  XNOR U10320 ( .A(n10151), .B(n10152), .Z(n10033) );
  NANDN U10321 ( .A(n10153), .B(n10154), .Z(n10152) );
  XOR U10322 ( .A(n10155), .B(n10024), .Z(n10026) );
  XOR U10323 ( .A(n10156), .B(n10157), .Z(n10024) );
  ANDN U10324 ( .B(n10158), .A(n10159), .Z(n10156) );
  AND U10325 ( .A(b[3]), .B(a[19]), .Z(n10155) );
  NAND U10326 ( .A(a[22]), .B(b[0]), .Z(n9909) );
  XNOR U10327 ( .A(n10039), .B(n10040), .Z(c[21]) );
  XNOR U10328 ( .A(n10153), .B(n10154), .Z(n10040) );
  XOR U10329 ( .A(n10151), .B(n10160), .Z(n10154) );
  NAND U10330 ( .A(b[1]), .B(a[20]), .Z(n10160) );
  XNOR U10331 ( .A(n10159), .B(n10161), .Z(n10153) );
  XOR U10332 ( .A(n10151), .B(n10158), .Z(n10161) );
  XNOR U10333 ( .A(n10162), .B(n10157), .Z(n10158) );
  AND U10334 ( .A(b[2]), .B(a[19]), .Z(n10162) );
  NANDN U10335 ( .A(n10163), .B(n10164), .Z(n10151) );
  XNOR U10336 ( .A(n10157), .B(n10165), .Z(n10159) );
  XNOR U10337 ( .A(n10145), .B(n10144), .Z(n10165) );
  XOR U10338 ( .A(n10166), .B(n10143), .Z(n10144) );
  AND U10339 ( .A(b[3]), .B(a[18]), .Z(n10166) );
  XNOR U10340 ( .A(n10143), .B(n10149), .Z(n10167) );
  XNOR U10341 ( .A(n10148), .B(n10140), .Z(n10168) );
  XNOR U10342 ( .A(n10139), .B(n10135), .Z(n10169) );
  XNOR U10343 ( .A(n10134), .B(n10130), .Z(n10170) );
  XNOR U10344 ( .A(n10129), .B(n10125), .Z(n10171) );
  XNOR U10345 ( .A(n10116), .B(n10115), .Z(n10172) );
  XOR U10346 ( .A(n10173), .B(n10114), .Z(n10115) );
  AND U10347 ( .A(b[9]), .B(a[12]), .Z(n10173) );
  XNOR U10348 ( .A(n10114), .B(n10120), .Z(n10174) );
  XNOR U10349 ( .A(n10119), .B(n10111), .Z(n10175) );
  XNOR U10350 ( .A(n10110), .B(n10106), .Z(n10176) );
  XNOR U10351 ( .A(n10105), .B(n10101), .Z(n10177) );
  XNOR U10352 ( .A(n10100), .B(n10096), .Z(n10178) );
  XNOR U10353 ( .A(n10087), .B(n10086), .Z(n10179) );
  XOR U10354 ( .A(n10180), .B(n10085), .Z(n10086) );
  AND U10355 ( .A(a[6]), .B(b[15]), .Z(n10180) );
  XNOR U10356 ( .A(n10085), .B(n10091), .Z(n10181) );
  XNOR U10357 ( .A(n10090), .B(n10082), .Z(n10182) );
  XNOR U10358 ( .A(n10081), .B(n10077), .Z(n10183) );
  XNOR U10359 ( .A(n10076), .B(n10072), .Z(n10184) );
  XNOR U10360 ( .A(n10071), .B(n10067), .Z(n10185) );
  XNOR U10361 ( .A(n10186), .B(n10066), .Z(n10067) );
  AND U10362 ( .A(a[0]), .B(b[21]), .Z(n10186) );
  XOR U10363 ( .A(n10187), .B(n10066), .Z(n10068) );
  XNOR U10364 ( .A(n10188), .B(n10189), .Z(n10066) );
  ANDN U10365 ( .B(n10190), .A(n10191), .Z(n10188) );
  AND U10366 ( .A(a[1]), .B(b[20]), .Z(n10187) );
  XNOR U10367 ( .A(n10192), .B(n10071), .Z(n10073) );
  XOR U10368 ( .A(n10193), .B(n10194), .Z(n10071) );
  ANDN U10369 ( .B(n10195), .A(n10196), .Z(n10193) );
  AND U10370 ( .A(a[2]), .B(b[19]), .Z(n10192) );
  XNOR U10371 ( .A(n10197), .B(n10076), .Z(n10078) );
  XOR U10372 ( .A(n10198), .B(n10199), .Z(n10076) );
  ANDN U10373 ( .B(n10200), .A(n10201), .Z(n10198) );
  AND U10374 ( .A(a[3]), .B(b[18]), .Z(n10197) );
  XNOR U10375 ( .A(n10202), .B(n10081), .Z(n10083) );
  XOR U10376 ( .A(n10203), .B(n10204), .Z(n10081) );
  ANDN U10377 ( .B(n10205), .A(n10206), .Z(n10203) );
  AND U10378 ( .A(a[4]), .B(b[17]), .Z(n10202) );
  XOR U10379 ( .A(n10207), .B(n10208), .Z(n10085) );
  AND U10380 ( .A(n10209), .B(n10210), .Z(n10207) );
  XNOR U10381 ( .A(n10211), .B(n10090), .Z(n10092) );
  XOR U10382 ( .A(n10212), .B(n10213), .Z(n10090) );
  ANDN U10383 ( .B(n10214), .A(n10215), .Z(n10212) );
  AND U10384 ( .A(a[5]), .B(b[16]), .Z(n10211) );
  XOR U10385 ( .A(n10216), .B(n10095), .Z(n10097) );
  XOR U10386 ( .A(n10217), .B(n10218), .Z(n10095) );
  ANDN U10387 ( .B(n10219), .A(n10220), .Z(n10217) );
  AND U10388 ( .A(a[7]), .B(b[14]), .Z(n10216) );
  XNOR U10389 ( .A(n10221), .B(n10100), .Z(n10102) );
  XOR U10390 ( .A(n10222), .B(n10223), .Z(n10100) );
  ANDN U10391 ( .B(n10224), .A(n10225), .Z(n10222) );
  AND U10392 ( .A(a[8]), .B(b[13]), .Z(n10221) );
  XNOR U10393 ( .A(n10226), .B(n10105), .Z(n10107) );
  XOR U10394 ( .A(n10227), .B(n10228), .Z(n10105) );
  ANDN U10395 ( .B(n10229), .A(n10230), .Z(n10227) );
  AND U10396 ( .A(a[9]), .B(b[12]), .Z(n10226) );
  XNOR U10397 ( .A(n10231), .B(n10110), .Z(n10112) );
  XOR U10398 ( .A(n10232), .B(n10233), .Z(n10110) );
  ANDN U10399 ( .B(n10234), .A(n10235), .Z(n10232) );
  AND U10400 ( .A(b[11]), .B(a[10]), .Z(n10231) );
  XOR U10401 ( .A(n10236), .B(n10237), .Z(n10114) );
  AND U10402 ( .A(n10238), .B(n10239), .Z(n10236) );
  XNOR U10403 ( .A(n10240), .B(n10119), .Z(n10121) );
  XOR U10404 ( .A(n10241), .B(n10242), .Z(n10119) );
  ANDN U10405 ( .B(n10243), .A(n10244), .Z(n10241) );
  AND U10406 ( .A(b[10]), .B(a[11]), .Z(n10240) );
  XOR U10407 ( .A(n10245), .B(n10124), .Z(n10126) );
  XOR U10408 ( .A(n10246), .B(n10247), .Z(n10124) );
  ANDN U10409 ( .B(n10248), .A(n10249), .Z(n10246) );
  AND U10410 ( .A(b[8]), .B(a[13]), .Z(n10245) );
  XNOR U10411 ( .A(n10250), .B(n10129), .Z(n10131) );
  XOR U10412 ( .A(n10251), .B(n10252), .Z(n10129) );
  ANDN U10413 ( .B(n10253), .A(n10254), .Z(n10251) );
  AND U10414 ( .A(b[7]), .B(a[14]), .Z(n10250) );
  XNOR U10415 ( .A(n10255), .B(n10134), .Z(n10136) );
  XOR U10416 ( .A(n10256), .B(n10257), .Z(n10134) );
  ANDN U10417 ( .B(n10258), .A(n10259), .Z(n10256) );
  AND U10418 ( .A(b[6]), .B(a[15]), .Z(n10255) );
  XNOR U10419 ( .A(n10260), .B(n10139), .Z(n10141) );
  XOR U10420 ( .A(n10261), .B(n10262), .Z(n10139) );
  ANDN U10421 ( .B(n10263), .A(n10264), .Z(n10261) );
  AND U10422 ( .A(b[5]), .B(a[16]), .Z(n10260) );
  XOR U10423 ( .A(n10265), .B(n10266), .Z(n10143) );
  ANDN U10424 ( .B(n10267), .A(n10268), .Z(n10265) );
  XNOR U10425 ( .A(n10269), .B(n10148), .Z(n10150) );
  XOR U10426 ( .A(n10270), .B(n10271), .Z(n10148) );
  ANDN U10427 ( .B(n10272), .A(n10273), .Z(n10270) );
  AND U10428 ( .A(b[4]), .B(a[17]), .Z(n10269) );
  XNOR U10429 ( .A(n10274), .B(n10275), .Z(n10157) );
  NAND U10430 ( .A(n10276), .B(n10277), .Z(n10275) );
  NAND U10431 ( .A(a[21]), .B(b[0]), .Z(n10039) );
  XNOR U10432 ( .A(n10163), .B(n10164), .Z(c[20]) );
  XOR U10433 ( .A(n10276), .B(n10277), .Z(n10164) );
  XOR U10434 ( .A(n10274), .B(n10278), .Z(n10277) );
  NAND U10435 ( .A(b[1]), .B(a[19]), .Z(n10278) );
  XOR U10436 ( .A(n10274), .B(n10267), .Z(n10279) );
  XNOR U10437 ( .A(n10266), .B(n10272), .Z(n10280) );
  XNOR U10438 ( .A(n10271), .B(n10263), .Z(n10281) );
  XNOR U10439 ( .A(n10262), .B(n10258), .Z(n10282) );
  XNOR U10440 ( .A(n10257), .B(n10253), .Z(n10283) );
  XNOR U10441 ( .A(n10252), .B(n10248), .Z(n10284) );
  XNOR U10442 ( .A(n10239), .B(n10238), .Z(n10285) );
  XOR U10443 ( .A(n10286), .B(n10237), .Z(n10238) );
  AND U10444 ( .A(b[8]), .B(a[12]), .Z(n10286) );
  XNOR U10445 ( .A(n10237), .B(n10243), .Z(n10287) );
  XNOR U10446 ( .A(n10242), .B(n10234), .Z(n10288) );
  XNOR U10447 ( .A(n10233), .B(n10229), .Z(n10289) );
  XNOR U10448 ( .A(n10228), .B(n10224), .Z(n10290) );
  XNOR U10449 ( .A(n10223), .B(n10219), .Z(n10291) );
  XNOR U10450 ( .A(n10210), .B(n10209), .Z(n10292) );
  XOR U10451 ( .A(n10293), .B(n10208), .Z(n10209) );
  AND U10452 ( .A(a[6]), .B(b[14]), .Z(n10293) );
  XNOR U10453 ( .A(n10208), .B(n10214), .Z(n10294) );
  XNOR U10454 ( .A(n10213), .B(n10205), .Z(n10295) );
  XNOR U10455 ( .A(n10204), .B(n10200), .Z(n10296) );
  XNOR U10456 ( .A(n10199), .B(n10195), .Z(n10297) );
  XNOR U10457 ( .A(n10194), .B(n10190), .Z(n10298) );
  XOR U10458 ( .A(n10299), .B(n10189), .Z(n10190) );
  AND U10459 ( .A(a[0]), .B(b[20]), .Z(n10299) );
  XNOR U10460 ( .A(n10300), .B(n10189), .Z(n10191) );
  XNOR U10461 ( .A(n10301), .B(n10302), .Z(n10189) );
  ANDN U10462 ( .B(n10303), .A(n10304), .Z(n10301) );
  AND U10463 ( .A(a[1]), .B(b[19]), .Z(n10300) );
  XNOR U10464 ( .A(n10305), .B(n10194), .Z(n10196) );
  XOR U10465 ( .A(n10306), .B(n10307), .Z(n10194) );
  ANDN U10466 ( .B(n10308), .A(n10309), .Z(n10306) );
  AND U10467 ( .A(a[2]), .B(b[18]), .Z(n10305) );
  XNOR U10468 ( .A(n10310), .B(n10199), .Z(n10201) );
  XOR U10469 ( .A(n10311), .B(n10312), .Z(n10199) );
  ANDN U10470 ( .B(n10313), .A(n10314), .Z(n10311) );
  AND U10471 ( .A(a[3]), .B(b[17]), .Z(n10310) );
  XNOR U10472 ( .A(n10315), .B(n10204), .Z(n10206) );
  XOR U10473 ( .A(n10316), .B(n10317), .Z(n10204) );
  ANDN U10474 ( .B(n10318), .A(n10319), .Z(n10316) );
  AND U10475 ( .A(a[4]), .B(b[16]), .Z(n10315) );
  XOR U10476 ( .A(n10320), .B(n10321), .Z(n10208) );
  AND U10477 ( .A(n10322), .B(n10323), .Z(n10320) );
  XNOR U10478 ( .A(n10324), .B(n10213), .Z(n10215) );
  XOR U10479 ( .A(n10325), .B(n10326), .Z(n10213) );
  ANDN U10480 ( .B(n10327), .A(n10328), .Z(n10325) );
  AND U10481 ( .A(a[5]), .B(b[15]), .Z(n10324) );
  XOR U10482 ( .A(n10329), .B(n10218), .Z(n10220) );
  XOR U10483 ( .A(n10330), .B(n10331), .Z(n10218) );
  ANDN U10484 ( .B(n10332), .A(n10333), .Z(n10330) );
  AND U10485 ( .A(a[7]), .B(b[13]), .Z(n10329) );
  XNOR U10486 ( .A(n10334), .B(n10223), .Z(n10225) );
  XOR U10487 ( .A(n10335), .B(n10336), .Z(n10223) );
  ANDN U10488 ( .B(n10337), .A(n10338), .Z(n10335) );
  AND U10489 ( .A(a[8]), .B(b[12]), .Z(n10334) );
  XNOR U10490 ( .A(n10339), .B(n10228), .Z(n10230) );
  XOR U10491 ( .A(n10340), .B(n10341), .Z(n10228) );
  ANDN U10492 ( .B(n10342), .A(n10343), .Z(n10340) );
  AND U10493 ( .A(a[9]), .B(b[11]), .Z(n10339) );
  XNOR U10494 ( .A(n10344), .B(n10233), .Z(n10235) );
  XOR U10495 ( .A(n10345), .B(n10346), .Z(n10233) );
  ANDN U10496 ( .B(n10347), .A(n10348), .Z(n10345) );
  AND U10497 ( .A(b[10]), .B(a[10]), .Z(n10344) );
  XOR U10498 ( .A(n10349), .B(n10350), .Z(n10237) );
  AND U10499 ( .A(n10351), .B(n10352), .Z(n10349) );
  XNOR U10500 ( .A(n10353), .B(n10242), .Z(n10244) );
  XOR U10501 ( .A(n10354), .B(n10355), .Z(n10242) );
  ANDN U10502 ( .B(n10356), .A(n10357), .Z(n10354) );
  AND U10503 ( .A(b[9]), .B(a[11]), .Z(n10353) );
  XOR U10504 ( .A(n10358), .B(n10247), .Z(n10249) );
  XOR U10505 ( .A(n10359), .B(n10360), .Z(n10247) );
  ANDN U10506 ( .B(n10361), .A(n10362), .Z(n10359) );
  AND U10507 ( .A(b[7]), .B(a[13]), .Z(n10358) );
  XNOR U10508 ( .A(n10363), .B(n10252), .Z(n10254) );
  XOR U10509 ( .A(n10364), .B(n10365), .Z(n10252) );
  ANDN U10510 ( .B(n10366), .A(n10367), .Z(n10364) );
  AND U10511 ( .A(b[6]), .B(a[14]), .Z(n10363) );
  XNOR U10512 ( .A(n10368), .B(n10257), .Z(n10259) );
  XOR U10513 ( .A(n10369), .B(n10370), .Z(n10257) );
  ANDN U10514 ( .B(n10371), .A(n10372), .Z(n10369) );
  AND U10515 ( .A(b[5]), .B(a[15]), .Z(n10368) );
  XNOR U10516 ( .A(n10373), .B(n10262), .Z(n10264) );
  XOR U10517 ( .A(n10374), .B(n10375), .Z(n10262) );
  ANDN U10518 ( .B(n10376), .A(n10377), .Z(n10374) );
  AND U10519 ( .A(b[4]), .B(a[16]), .Z(n10373) );
  XNOR U10520 ( .A(n10378), .B(n10271), .Z(n10273) );
  XNOR U10521 ( .A(n10379), .B(n10380), .Z(n10271) );
  NOR U10522 ( .A(n10381), .B(n10382), .Z(n10379) );
  AND U10523 ( .A(b[3]), .B(a[17]), .Z(n10378) );
  NANDN U10524 ( .A(n10383), .B(n10384), .Z(n10274) );
  XNOR U10525 ( .A(n10385), .B(n10266), .Z(n10268) );
  XNOR U10526 ( .A(n10386), .B(n10387), .Z(n10266) );
  OR U10527 ( .A(n10388), .B(n10389), .Z(n10387) );
  AND U10528 ( .A(b[2]), .B(a[18]), .Z(n10385) );
  NAND U10529 ( .A(a[20]), .B(b[0]), .Z(n10163) );
  XOR U10530 ( .A(n10390), .B(n10391), .Z(c[1]) );
  XNOR U10531 ( .A(n10383), .B(n10384), .Z(c[19]) );
  XOR U10532 ( .A(n10389), .B(n10388), .Z(n10384) );
  XOR U10533 ( .A(n10386), .B(n10392), .Z(n10388) );
  NAND U10534 ( .A(b[1]), .B(a[18]), .Z(n10392) );
  XOR U10535 ( .A(n10386), .B(n10382), .Z(n10393) );
  XOR U10536 ( .A(n10394), .B(n10380), .Z(n10382) );
  AND U10537 ( .A(b[2]), .B(a[17]), .Z(n10394) );
  ANDN U10538 ( .B(n10395), .A(n10396), .Z(n10386) );
  XOR U10539 ( .A(n10380), .B(n10376), .Z(n10397) );
  XNOR U10540 ( .A(n10375), .B(n10371), .Z(n10398) );
  XNOR U10541 ( .A(n10370), .B(n10366), .Z(n10399) );
  XNOR U10542 ( .A(n10365), .B(n10361), .Z(n10400) );
  XNOR U10543 ( .A(n10352), .B(n10351), .Z(n10401) );
  XOR U10544 ( .A(n10402), .B(n10350), .Z(n10351) );
  AND U10545 ( .A(b[7]), .B(a[12]), .Z(n10402) );
  XNOR U10546 ( .A(n10350), .B(n10356), .Z(n10403) );
  XNOR U10547 ( .A(n10355), .B(n10347), .Z(n10404) );
  XNOR U10548 ( .A(n10346), .B(n10342), .Z(n10405) );
  XNOR U10549 ( .A(n10341), .B(n10337), .Z(n10406) );
  XNOR U10550 ( .A(n10336), .B(n10332), .Z(n10407) );
  XNOR U10551 ( .A(n10323), .B(n10322), .Z(n10408) );
  XOR U10552 ( .A(n10409), .B(n10321), .Z(n10322) );
  AND U10553 ( .A(a[6]), .B(b[13]), .Z(n10409) );
  XNOR U10554 ( .A(n10321), .B(n10327), .Z(n10410) );
  XNOR U10555 ( .A(n10326), .B(n10318), .Z(n10411) );
  XNOR U10556 ( .A(n10317), .B(n10313), .Z(n10412) );
  XNOR U10557 ( .A(n10312), .B(n10308), .Z(n10413) );
  XNOR U10558 ( .A(n10307), .B(n10303), .Z(n10414) );
  XNOR U10559 ( .A(n10415), .B(n10302), .Z(n10303) );
  AND U10560 ( .A(a[0]), .B(b[19]), .Z(n10415) );
  XOR U10561 ( .A(n10416), .B(n10302), .Z(n10304) );
  XNOR U10562 ( .A(n10417), .B(n10418), .Z(n10302) );
  ANDN U10563 ( .B(n10419), .A(n10420), .Z(n10417) );
  AND U10564 ( .A(a[1]), .B(b[18]), .Z(n10416) );
  XNOR U10565 ( .A(n10421), .B(n10307), .Z(n10309) );
  XOR U10566 ( .A(n10422), .B(n10423), .Z(n10307) );
  ANDN U10567 ( .B(n10424), .A(n10425), .Z(n10422) );
  AND U10568 ( .A(a[2]), .B(b[17]), .Z(n10421) );
  XNOR U10569 ( .A(n10426), .B(n10312), .Z(n10314) );
  XOR U10570 ( .A(n10427), .B(n10428), .Z(n10312) );
  ANDN U10571 ( .B(n10429), .A(n10430), .Z(n10427) );
  AND U10572 ( .A(a[3]), .B(b[16]), .Z(n10426) );
  XNOR U10573 ( .A(n10431), .B(n10317), .Z(n10319) );
  XOR U10574 ( .A(n10432), .B(n10433), .Z(n10317) );
  ANDN U10575 ( .B(n10434), .A(n10435), .Z(n10432) );
  AND U10576 ( .A(a[4]), .B(b[15]), .Z(n10431) );
  XOR U10577 ( .A(n10436), .B(n10437), .Z(n10321) );
  AND U10578 ( .A(n10438), .B(n10439), .Z(n10436) );
  XNOR U10579 ( .A(n10440), .B(n10326), .Z(n10328) );
  XOR U10580 ( .A(n10441), .B(n10442), .Z(n10326) );
  ANDN U10581 ( .B(n10443), .A(n10444), .Z(n10441) );
  AND U10582 ( .A(a[5]), .B(b[14]), .Z(n10440) );
  XOR U10583 ( .A(n10445), .B(n10331), .Z(n10333) );
  XOR U10584 ( .A(n10446), .B(n10447), .Z(n10331) );
  ANDN U10585 ( .B(n10448), .A(n10449), .Z(n10446) );
  AND U10586 ( .A(a[7]), .B(b[12]), .Z(n10445) );
  XNOR U10587 ( .A(n10450), .B(n10336), .Z(n10338) );
  XOR U10588 ( .A(n10451), .B(n10452), .Z(n10336) );
  ANDN U10589 ( .B(n10453), .A(n10454), .Z(n10451) );
  AND U10590 ( .A(a[8]), .B(b[11]), .Z(n10450) );
  XNOR U10591 ( .A(n10455), .B(n10341), .Z(n10343) );
  XOR U10592 ( .A(n10456), .B(n10457), .Z(n10341) );
  ANDN U10593 ( .B(n10458), .A(n10459), .Z(n10456) );
  AND U10594 ( .A(a[9]), .B(b[10]), .Z(n10455) );
  XNOR U10595 ( .A(n10460), .B(n10346), .Z(n10348) );
  XOR U10596 ( .A(n10461), .B(n10462), .Z(n10346) );
  ANDN U10597 ( .B(n10463), .A(n10464), .Z(n10461) );
  AND U10598 ( .A(b[9]), .B(a[10]), .Z(n10460) );
  XOR U10599 ( .A(n10465), .B(n10466), .Z(n10350) );
  AND U10600 ( .A(n10467), .B(n10468), .Z(n10465) );
  XNOR U10601 ( .A(n10469), .B(n10355), .Z(n10357) );
  XOR U10602 ( .A(n10470), .B(n10471), .Z(n10355) );
  ANDN U10603 ( .B(n10472), .A(n10473), .Z(n10470) );
  AND U10604 ( .A(b[8]), .B(a[11]), .Z(n10469) );
  XOR U10605 ( .A(n10474), .B(n10360), .Z(n10362) );
  XOR U10606 ( .A(n10475), .B(n10476), .Z(n10360) );
  ANDN U10607 ( .B(n10477), .A(n10478), .Z(n10475) );
  AND U10608 ( .A(b[6]), .B(a[13]), .Z(n10474) );
  XNOR U10609 ( .A(n10479), .B(n10365), .Z(n10367) );
  XOR U10610 ( .A(n10480), .B(n10481), .Z(n10365) );
  ANDN U10611 ( .B(n10482), .A(n10483), .Z(n10480) );
  AND U10612 ( .A(b[5]), .B(a[14]), .Z(n10479) );
  XNOR U10613 ( .A(n10484), .B(n10370), .Z(n10372) );
  XOR U10614 ( .A(n10485), .B(n10486), .Z(n10370) );
  ANDN U10615 ( .B(n10487), .A(n10488), .Z(n10485) );
  AND U10616 ( .A(b[4]), .B(a[15]), .Z(n10484) );
  XNOR U10617 ( .A(n10489), .B(n10490), .Z(n10380) );
  NANDN U10618 ( .A(n10491), .B(n10492), .Z(n10490) );
  XNOR U10619 ( .A(n10493), .B(n10375), .Z(n10377) );
  XNOR U10620 ( .A(n10494), .B(n10495), .Z(n10375) );
  AND U10621 ( .A(n10496), .B(n10497), .Z(n10494) );
  AND U10622 ( .A(b[3]), .B(a[16]), .Z(n10493) );
  NAND U10623 ( .A(a[19]), .B(b[0]), .Z(n10383) );
  XNOR U10624 ( .A(n10396), .B(n10395), .Z(c[18]) );
  XNOR U10625 ( .A(n10491), .B(n10492), .Z(n10395) );
  XOR U10626 ( .A(n10489), .B(n10498), .Z(n10492) );
  NAND U10627 ( .A(b[1]), .B(a[17]), .Z(n10498) );
  XOR U10628 ( .A(n10497), .B(n10499), .Z(n10491) );
  XOR U10629 ( .A(n10489), .B(n10496), .Z(n10499) );
  XNOR U10630 ( .A(n10500), .B(n10495), .Z(n10496) );
  AND U10631 ( .A(b[2]), .B(a[16]), .Z(n10500) );
  NANDN U10632 ( .A(n10501), .B(n10502), .Z(n10489) );
  XOR U10633 ( .A(n10495), .B(n10487), .Z(n10503) );
  XNOR U10634 ( .A(n10486), .B(n10482), .Z(n10504) );
  XNOR U10635 ( .A(n10481), .B(n10477), .Z(n10505) );
  XNOR U10636 ( .A(n10468), .B(n10467), .Z(n10506) );
  XOR U10637 ( .A(n10507), .B(n10466), .Z(n10467) );
  AND U10638 ( .A(b[6]), .B(a[12]), .Z(n10507) );
  XNOR U10639 ( .A(n10466), .B(n10472), .Z(n10508) );
  XNOR U10640 ( .A(n10471), .B(n10463), .Z(n10509) );
  XNOR U10641 ( .A(n10462), .B(n10458), .Z(n10510) );
  XNOR U10642 ( .A(n10457), .B(n10453), .Z(n10511) );
  XNOR U10643 ( .A(n10452), .B(n10448), .Z(n10512) );
  XNOR U10644 ( .A(n10439), .B(n10438), .Z(n10513) );
  XOR U10645 ( .A(n10514), .B(n10437), .Z(n10438) );
  AND U10646 ( .A(a[6]), .B(b[12]), .Z(n10514) );
  XNOR U10647 ( .A(n10437), .B(n10443), .Z(n10515) );
  XNOR U10648 ( .A(n10442), .B(n10434), .Z(n10516) );
  XNOR U10649 ( .A(n10433), .B(n10429), .Z(n10517) );
  XNOR U10650 ( .A(n10428), .B(n10424), .Z(n10518) );
  XNOR U10651 ( .A(n10423), .B(n10419), .Z(n10519) );
  XOR U10652 ( .A(n10520), .B(n10418), .Z(n10419) );
  AND U10653 ( .A(a[0]), .B(b[18]), .Z(n10520) );
  XNOR U10654 ( .A(n10521), .B(n10418), .Z(n10420) );
  XNOR U10655 ( .A(n10522), .B(n10523), .Z(n10418) );
  ANDN U10656 ( .B(n10524), .A(n10525), .Z(n10522) );
  AND U10657 ( .A(a[1]), .B(b[17]), .Z(n10521) );
  XNOR U10658 ( .A(n10526), .B(n10423), .Z(n10425) );
  XOR U10659 ( .A(n10527), .B(n10528), .Z(n10423) );
  ANDN U10660 ( .B(n10529), .A(n10530), .Z(n10527) );
  AND U10661 ( .A(a[2]), .B(b[16]), .Z(n10526) );
  XNOR U10662 ( .A(n10531), .B(n10428), .Z(n10430) );
  XOR U10663 ( .A(n10532), .B(n10533), .Z(n10428) );
  ANDN U10664 ( .B(n10534), .A(n10535), .Z(n10532) );
  AND U10665 ( .A(a[3]), .B(b[15]), .Z(n10531) );
  XNOR U10666 ( .A(n10536), .B(n10433), .Z(n10435) );
  XOR U10667 ( .A(n10537), .B(n10538), .Z(n10433) );
  ANDN U10668 ( .B(n10539), .A(n10540), .Z(n10537) );
  AND U10669 ( .A(a[4]), .B(b[14]), .Z(n10536) );
  XOR U10670 ( .A(n10541), .B(n10542), .Z(n10437) );
  AND U10671 ( .A(n10543), .B(n10544), .Z(n10541) );
  XNOR U10672 ( .A(n10545), .B(n10442), .Z(n10444) );
  XOR U10673 ( .A(n10546), .B(n10547), .Z(n10442) );
  ANDN U10674 ( .B(n10548), .A(n10549), .Z(n10546) );
  AND U10675 ( .A(a[5]), .B(b[13]), .Z(n10545) );
  XOR U10676 ( .A(n10550), .B(n10447), .Z(n10449) );
  XOR U10677 ( .A(n10551), .B(n10552), .Z(n10447) );
  ANDN U10678 ( .B(n10553), .A(n10554), .Z(n10551) );
  AND U10679 ( .A(a[7]), .B(b[11]), .Z(n10550) );
  XNOR U10680 ( .A(n10555), .B(n10452), .Z(n10454) );
  XOR U10681 ( .A(n10556), .B(n10557), .Z(n10452) );
  ANDN U10682 ( .B(n10558), .A(n10559), .Z(n10556) );
  AND U10683 ( .A(a[8]), .B(b[10]), .Z(n10555) );
  XNOR U10684 ( .A(n10560), .B(n10457), .Z(n10459) );
  XOR U10685 ( .A(n10561), .B(n10562), .Z(n10457) );
  ANDN U10686 ( .B(n10563), .A(n10564), .Z(n10561) );
  AND U10687 ( .A(a[9]), .B(b[9]), .Z(n10560) );
  XNOR U10688 ( .A(n10565), .B(n10462), .Z(n10464) );
  XOR U10689 ( .A(n10566), .B(n10567), .Z(n10462) );
  ANDN U10690 ( .B(n10568), .A(n10569), .Z(n10566) );
  AND U10691 ( .A(b[8]), .B(a[10]), .Z(n10565) );
  XOR U10692 ( .A(n10570), .B(n10571), .Z(n10466) );
  AND U10693 ( .A(n10572), .B(n10573), .Z(n10570) );
  XNOR U10694 ( .A(n10574), .B(n10471), .Z(n10473) );
  XOR U10695 ( .A(n10575), .B(n10576), .Z(n10471) );
  ANDN U10696 ( .B(n10577), .A(n10578), .Z(n10575) );
  AND U10697 ( .A(b[7]), .B(a[11]), .Z(n10574) );
  XOR U10698 ( .A(n10579), .B(n10476), .Z(n10478) );
  XOR U10699 ( .A(n10580), .B(n10581), .Z(n10476) );
  ANDN U10700 ( .B(n10582), .A(n10583), .Z(n10580) );
  AND U10701 ( .A(b[5]), .B(a[13]), .Z(n10579) );
  XNOR U10702 ( .A(n10584), .B(n10481), .Z(n10483) );
  XOR U10703 ( .A(n10585), .B(n10586), .Z(n10481) );
  ANDN U10704 ( .B(n10587), .A(n10588), .Z(n10585) );
  AND U10705 ( .A(b[4]), .B(a[14]), .Z(n10584) );
  XNOR U10706 ( .A(n10589), .B(n10590), .Z(n10495) );
  NANDN U10707 ( .A(n10591), .B(n10592), .Z(n10590) );
  XNOR U10708 ( .A(n10593), .B(n10486), .Z(n10488) );
  XNOR U10709 ( .A(n10594), .B(n10595), .Z(n10486) );
  AND U10710 ( .A(n10596), .B(n10597), .Z(n10594) );
  AND U10711 ( .A(b[3]), .B(a[15]), .Z(n10593) );
  NAND U10712 ( .A(a[18]), .B(b[0]), .Z(n10396) );
  XNOR U10713 ( .A(n10501), .B(n10502), .Z(c[17]) );
  XNOR U10714 ( .A(n10591), .B(n10592), .Z(n10502) );
  XOR U10715 ( .A(n10589), .B(n10598), .Z(n10592) );
  NAND U10716 ( .A(b[1]), .B(a[16]), .Z(n10598) );
  XOR U10717 ( .A(n10597), .B(n10599), .Z(n10591) );
  XOR U10718 ( .A(n10589), .B(n10596), .Z(n10599) );
  XNOR U10719 ( .A(n10600), .B(n10595), .Z(n10596) );
  AND U10720 ( .A(b[2]), .B(a[15]), .Z(n10600) );
  NANDN U10721 ( .A(n10601), .B(n10602), .Z(n10589) );
  XOR U10722 ( .A(n10595), .B(n10587), .Z(n10603) );
  XNOR U10723 ( .A(n10586), .B(n10582), .Z(n10604) );
  XNOR U10724 ( .A(n10573), .B(n10572), .Z(n10605) );
  XOR U10725 ( .A(n10606), .B(n10571), .Z(n10572) );
  AND U10726 ( .A(b[5]), .B(a[12]), .Z(n10606) );
  XNOR U10727 ( .A(n10571), .B(n10577), .Z(n10607) );
  XNOR U10728 ( .A(n10576), .B(n10568), .Z(n10608) );
  XNOR U10729 ( .A(n10567), .B(n10563), .Z(n10609) );
  XNOR U10730 ( .A(n10562), .B(n10558), .Z(n10610) );
  XNOR U10731 ( .A(n10557), .B(n10553), .Z(n10611) );
  XNOR U10732 ( .A(n10544), .B(n10543), .Z(n10612) );
  XOR U10733 ( .A(n10613), .B(n10542), .Z(n10543) );
  AND U10734 ( .A(a[6]), .B(b[11]), .Z(n10613) );
  XNOR U10735 ( .A(n10542), .B(n10548), .Z(n10614) );
  XNOR U10736 ( .A(n10547), .B(n10539), .Z(n10615) );
  XNOR U10737 ( .A(n10538), .B(n10534), .Z(n10616) );
  XNOR U10738 ( .A(n10533), .B(n10529), .Z(n10617) );
  XNOR U10739 ( .A(n10528), .B(n10524), .Z(n10618) );
  XNOR U10740 ( .A(n10619), .B(n10523), .Z(n10524) );
  AND U10741 ( .A(a[0]), .B(b[17]), .Z(n10619) );
  XOR U10742 ( .A(n10620), .B(n10523), .Z(n10525) );
  XNOR U10743 ( .A(n10621), .B(n10622), .Z(n10523) );
  ANDN U10744 ( .B(n10623), .A(n10624), .Z(n10621) );
  AND U10745 ( .A(a[1]), .B(b[16]), .Z(n10620) );
  XNOR U10746 ( .A(n10625), .B(n10528), .Z(n10530) );
  XOR U10747 ( .A(n10626), .B(n10627), .Z(n10528) );
  ANDN U10748 ( .B(n10628), .A(n10629), .Z(n10626) );
  AND U10749 ( .A(a[2]), .B(b[15]), .Z(n10625) );
  XNOR U10750 ( .A(n10630), .B(n10533), .Z(n10535) );
  XOR U10751 ( .A(n10631), .B(n10632), .Z(n10533) );
  ANDN U10752 ( .B(n10633), .A(n10634), .Z(n10631) );
  AND U10753 ( .A(a[3]), .B(b[14]), .Z(n10630) );
  XNOR U10754 ( .A(n10635), .B(n10538), .Z(n10540) );
  XOR U10755 ( .A(n10636), .B(n10637), .Z(n10538) );
  ANDN U10756 ( .B(n10638), .A(n10639), .Z(n10636) );
  AND U10757 ( .A(a[4]), .B(b[13]), .Z(n10635) );
  XOR U10758 ( .A(n10640), .B(n10641), .Z(n10542) );
  AND U10759 ( .A(n10642), .B(n10643), .Z(n10640) );
  XNOR U10760 ( .A(n10644), .B(n10547), .Z(n10549) );
  XOR U10761 ( .A(n10645), .B(n10646), .Z(n10547) );
  ANDN U10762 ( .B(n10647), .A(n10648), .Z(n10645) );
  AND U10763 ( .A(a[5]), .B(b[12]), .Z(n10644) );
  XOR U10764 ( .A(n10649), .B(n10552), .Z(n10554) );
  XOR U10765 ( .A(n10650), .B(n10651), .Z(n10552) );
  ANDN U10766 ( .B(n10652), .A(n10653), .Z(n10650) );
  AND U10767 ( .A(a[7]), .B(b[10]), .Z(n10649) );
  XNOR U10768 ( .A(n10654), .B(n10557), .Z(n10559) );
  XOR U10769 ( .A(n10655), .B(n10656), .Z(n10557) );
  ANDN U10770 ( .B(n10657), .A(n10658), .Z(n10655) );
  AND U10771 ( .A(a[8]), .B(b[9]), .Z(n10654) );
  XNOR U10772 ( .A(n10659), .B(n10562), .Z(n10564) );
  XOR U10773 ( .A(n10660), .B(n10661), .Z(n10562) );
  ANDN U10774 ( .B(n10662), .A(n10663), .Z(n10660) );
  AND U10775 ( .A(a[9]), .B(b[8]), .Z(n10659) );
  XNOR U10776 ( .A(n10664), .B(n10567), .Z(n10569) );
  XOR U10777 ( .A(n10665), .B(n10666), .Z(n10567) );
  ANDN U10778 ( .B(n10667), .A(n10668), .Z(n10665) );
  AND U10779 ( .A(b[7]), .B(a[10]), .Z(n10664) );
  XOR U10780 ( .A(n10669), .B(n10670), .Z(n10571) );
  AND U10781 ( .A(n10671), .B(n10672), .Z(n10669) );
  XNOR U10782 ( .A(n10673), .B(n10576), .Z(n10578) );
  XOR U10783 ( .A(n10674), .B(n10675), .Z(n10576) );
  ANDN U10784 ( .B(n10676), .A(n10677), .Z(n10674) );
  AND U10785 ( .A(b[6]), .B(a[11]), .Z(n10673) );
  XOR U10786 ( .A(n10678), .B(n10581), .Z(n10583) );
  XOR U10787 ( .A(n10679), .B(n10680), .Z(n10581) );
  ANDN U10788 ( .B(n10681), .A(n10682), .Z(n10679) );
  AND U10789 ( .A(b[4]), .B(a[13]), .Z(n10678) );
  XNOR U10790 ( .A(n10683), .B(n10684), .Z(n10595) );
  NANDN U10791 ( .A(n10685), .B(n10686), .Z(n10684) );
  XNOR U10792 ( .A(n10687), .B(n10586), .Z(n10588) );
  XNOR U10793 ( .A(n10688), .B(n10689), .Z(n10586) );
  AND U10794 ( .A(n10690), .B(n10691), .Z(n10688) );
  AND U10795 ( .A(b[3]), .B(a[14]), .Z(n10687) );
  NAND U10796 ( .A(a[17]), .B(b[0]), .Z(n10501) );
  XNOR U10797 ( .A(n10601), .B(n10602), .Z(c[16]) );
  XNOR U10798 ( .A(n10685), .B(n10686), .Z(n10602) );
  XOR U10799 ( .A(n10683), .B(n10692), .Z(n10686) );
  NAND U10800 ( .A(b[1]), .B(a[15]), .Z(n10692) );
  XOR U10801 ( .A(n10691), .B(n10693), .Z(n10685) );
  XOR U10802 ( .A(n10683), .B(n10690), .Z(n10693) );
  XNOR U10803 ( .A(n10694), .B(n10689), .Z(n10690) );
  AND U10804 ( .A(b[2]), .B(a[14]), .Z(n10694) );
  NANDN U10805 ( .A(n10695), .B(n10696), .Z(n10683) );
  XOR U10806 ( .A(n10689), .B(n10681), .Z(n10697) );
  XNOR U10807 ( .A(n10672), .B(n10671), .Z(n10698) );
  XOR U10808 ( .A(n10699), .B(n10670), .Z(n10671) );
  AND U10809 ( .A(b[4]), .B(a[12]), .Z(n10699) );
  XNOR U10810 ( .A(n10670), .B(n10676), .Z(n10700) );
  XNOR U10811 ( .A(n10675), .B(n10667), .Z(n10701) );
  XNOR U10812 ( .A(n10666), .B(n10662), .Z(n10702) );
  XNOR U10813 ( .A(n10661), .B(n10657), .Z(n10703) );
  XNOR U10814 ( .A(n10656), .B(n10652), .Z(n10704) );
  XNOR U10815 ( .A(n10643), .B(n10642), .Z(n10705) );
  XOR U10816 ( .A(n10706), .B(n10641), .Z(n10642) );
  AND U10817 ( .A(a[6]), .B(b[10]), .Z(n10706) );
  XNOR U10818 ( .A(n10641), .B(n10647), .Z(n10707) );
  XNOR U10819 ( .A(n10646), .B(n10638), .Z(n10708) );
  XNOR U10820 ( .A(n10637), .B(n10633), .Z(n10709) );
  XNOR U10821 ( .A(n10632), .B(n10628), .Z(n10710) );
  XNOR U10822 ( .A(n10627), .B(n10623), .Z(n10711) );
  XOR U10823 ( .A(n10712), .B(n10622), .Z(n10623) );
  AND U10824 ( .A(a[0]), .B(b[16]), .Z(n10712) );
  XNOR U10825 ( .A(n10713), .B(n10622), .Z(n10624) );
  XNOR U10826 ( .A(n10714), .B(n10715), .Z(n10622) );
  ANDN U10827 ( .B(n10716), .A(n10717), .Z(n10714) );
  AND U10828 ( .A(a[1]), .B(b[15]), .Z(n10713) );
  XNOR U10829 ( .A(n10718), .B(n10627), .Z(n10629) );
  XOR U10830 ( .A(n10719), .B(n10720), .Z(n10627) );
  ANDN U10831 ( .B(n10721), .A(n10722), .Z(n10719) );
  AND U10832 ( .A(a[2]), .B(b[14]), .Z(n10718) );
  XNOR U10833 ( .A(n10723), .B(n10632), .Z(n10634) );
  XOR U10834 ( .A(n10724), .B(n10725), .Z(n10632) );
  ANDN U10835 ( .B(n10726), .A(n10727), .Z(n10724) );
  AND U10836 ( .A(a[3]), .B(b[13]), .Z(n10723) );
  XNOR U10837 ( .A(n10728), .B(n10637), .Z(n10639) );
  XOR U10838 ( .A(n10729), .B(n10730), .Z(n10637) );
  ANDN U10839 ( .B(n10731), .A(n10732), .Z(n10729) );
  AND U10840 ( .A(a[4]), .B(b[12]), .Z(n10728) );
  XOR U10841 ( .A(n10733), .B(n10734), .Z(n10641) );
  AND U10842 ( .A(n10735), .B(n10736), .Z(n10733) );
  XNOR U10843 ( .A(n10737), .B(n10646), .Z(n10648) );
  XOR U10844 ( .A(n10738), .B(n10739), .Z(n10646) );
  ANDN U10845 ( .B(n10740), .A(n10741), .Z(n10738) );
  AND U10846 ( .A(a[5]), .B(b[11]), .Z(n10737) );
  XOR U10847 ( .A(n10742), .B(n10651), .Z(n10653) );
  XOR U10848 ( .A(n10743), .B(n10744), .Z(n10651) );
  ANDN U10849 ( .B(n10745), .A(n10746), .Z(n10743) );
  AND U10850 ( .A(a[7]), .B(b[9]), .Z(n10742) );
  XNOR U10851 ( .A(n10747), .B(n10656), .Z(n10658) );
  XOR U10852 ( .A(n10748), .B(n10749), .Z(n10656) );
  ANDN U10853 ( .B(n10750), .A(n10751), .Z(n10748) );
  AND U10854 ( .A(a[8]), .B(b[8]), .Z(n10747) );
  XNOR U10855 ( .A(n10752), .B(n10661), .Z(n10663) );
  XOR U10856 ( .A(n10753), .B(n10754), .Z(n10661) );
  ANDN U10857 ( .B(n10755), .A(n10756), .Z(n10753) );
  AND U10858 ( .A(a[9]), .B(b[7]), .Z(n10752) );
  XNOR U10859 ( .A(n10757), .B(n10666), .Z(n10668) );
  XOR U10860 ( .A(n10758), .B(n10759), .Z(n10666) );
  ANDN U10861 ( .B(n10760), .A(n10761), .Z(n10758) );
  AND U10862 ( .A(b[6]), .B(a[10]), .Z(n10757) );
  XOR U10863 ( .A(n10762), .B(n10763), .Z(n10670) );
  AND U10864 ( .A(n10764), .B(n10765), .Z(n10762) );
  XNOR U10865 ( .A(n10766), .B(n10675), .Z(n10677) );
  XOR U10866 ( .A(n10767), .B(n10768), .Z(n10675) );
  ANDN U10867 ( .B(n10769), .A(n10770), .Z(n10767) );
  AND U10868 ( .A(b[5]), .B(a[11]), .Z(n10766) );
  XNOR U10869 ( .A(n10771), .B(n10772), .Z(n10689) );
  NANDN U10870 ( .A(n10773), .B(n10774), .Z(n10772) );
  XOR U10871 ( .A(n10775), .B(n10680), .Z(n10682) );
  XOR U10872 ( .A(n10776), .B(n10777), .Z(n10680) );
  ANDN U10873 ( .B(n10778), .A(n10779), .Z(n10776) );
  AND U10874 ( .A(b[3]), .B(a[13]), .Z(n10775) );
  NAND U10875 ( .A(a[16]), .B(b[0]), .Z(n10601) );
  XNOR U10876 ( .A(n10695), .B(n10696), .Z(c[15]) );
  XNOR U10877 ( .A(n10773), .B(n10774), .Z(n10696) );
  XOR U10878 ( .A(n10771), .B(n10780), .Z(n10774) );
  NAND U10879 ( .A(b[1]), .B(a[14]), .Z(n10780) );
  XNOR U10880 ( .A(n10779), .B(n10781), .Z(n10773) );
  XOR U10881 ( .A(n10771), .B(n10778), .Z(n10781) );
  XNOR U10882 ( .A(n10782), .B(n10777), .Z(n10778) );
  AND U10883 ( .A(b[2]), .B(a[13]), .Z(n10782) );
  NANDN U10884 ( .A(n10783), .B(n10784), .Z(n10771) );
  XNOR U10885 ( .A(n10777), .B(n10785), .Z(n10779) );
  XNOR U10886 ( .A(n10765), .B(n10764), .Z(n10785) );
  XOR U10887 ( .A(n10786), .B(n10763), .Z(n10764) );
  AND U10888 ( .A(b[3]), .B(a[12]), .Z(n10786) );
  XNOR U10889 ( .A(n10763), .B(n10769), .Z(n10787) );
  XNOR U10890 ( .A(n10768), .B(n10760), .Z(n10788) );
  XNOR U10891 ( .A(n10759), .B(n10755), .Z(n10789) );
  XNOR U10892 ( .A(n10754), .B(n10750), .Z(n10790) );
  XNOR U10893 ( .A(n10749), .B(n10745), .Z(n10791) );
  XNOR U10894 ( .A(n10736), .B(n10735), .Z(n10792) );
  XOR U10895 ( .A(n10793), .B(n10734), .Z(n10735) );
  AND U10896 ( .A(a[6]), .B(b[9]), .Z(n10793) );
  XNOR U10897 ( .A(n10734), .B(n10740), .Z(n10794) );
  XNOR U10898 ( .A(n10739), .B(n10731), .Z(n10795) );
  XNOR U10899 ( .A(n10730), .B(n10726), .Z(n10796) );
  XNOR U10900 ( .A(n10725), .B(n10721), .Z(n10797) );
  XNOR U10901 ( .A(n10720), .B(n10716), .Z(n10798) );
  XNOR U10902 ( .A(n10799), .B(n10715), .Z(n10716) );
  AND U10903 ( .A(a[0]), .B(b[15]), .Z(n10799) );
  XOR U10904 ( .A(n10800), .B(n10715), .Z(n10717) );
  XNOR U10905 ( .A(n10801), .B(n10802), .Z(n10715) );
  ANDN U10906 ( .B(n10803), .A(n10804), .Z(n10801) );
  AND U10907 ( .A(a[1]), .B(b[14]), .Z(n10800) );
  XNOR U10908 ( .A(n10805), .B(n10720), .Z(n10722) );
  XOR U10909 ( .A(n10806), .B(n10807), .Z(n10720) );
  ANDN U10910 ( .B(n10808), .A(n10809), .Z(n10806) );
  AND U10911 ( .A(a[2]), .B(b[13]), .Z(n10805) );
  XNOR U10912 ( .A(n10810), .B(n10725), .Z(n10727) );
  XOR U10913 ( .A(n10811), .B(n10812), .Z(n10725) );
  ANDN U10914 ( .B(n10813), .A(n10814), .Z(n10811) );
  AND U10915 ( .A(a[3]), .B(b[12]), .Z(n10810) );
  XNOR U10916 ( .A(n10815), .B(n10730), .Z(n10732) );
  XOR U10917 ( .A(n10816), .B(n10817), .Z(n10730) );
  ANDN U10918 ( .B(n10818), .A(n10819), .Z(n10816) );
  AND U10919 ( .A(a[4]), .B(b[11]), .Z(n10815) );
  XOR U10920 ( .A(n10820), .B(n10821), .Z(n10734) );
  AND U10921 ( .A(n10822), .B(n10823), .Z(n10820) );
  XNOR U10922 ( .A(n10824), .B(n10739), .Z(n10741) );
  XOR U10923 ( .A(n10825), .B(n10826), .Z(n10739) );
  ANDN U10924 ( .B(n10827), .A(n10828), .Z(n10825) );
  AND U10925 ( .A(a[5]), .B(b[10]), .Z(n10824) );
  XOR U10926 ( .A(n10829), .B(n10744), .Z(n10746) );
  XOR U10927 ( .A(n10830), .B(n10831), .Z(n10744) );
  ANDN U10928 ( .B(n10832), .A(n10833), .Z(n10830) );
  AND U10929 ( .A(a[7]), .B(b[8]), .Z(n10829) );
  XNOR U10930 ( .A(n10834), .B(n10749), .Z(n10751) );
  XOR U10931 ( .A(n10835), .B(n10836), .Z(n10749) );
  ANDN U10932 ( .B(n10837), .A(n10838), .Z(n10835) );
  AND U10933 ( .A(a[8]), .B(b[7]), .Z(n10834) );
  XNOR U10934 ( .A(n10839), .B(n10754), .Z(n10756) );
  XOR U10935 ( .A(n10840), .B(n10841), .Z(n10754) );
  ANDN U10936 ( .B(n10842), .A(n10843), .Z(n10840) );
  AND U10937 ( .A(a[9]), .B(b[6]), .Z(n10839) );
  XNOR U10938 ( .A(n10844), .B(n10759), .Z(n10761) );
  XOR U10939 ( .A(n10845), .B(n10846), .Z(n10759) );
  ANDN U10940 ( .B(n10847), .A(n10848), .Z(n10845) );
  AND U10941 ( .A(b[5]), .B(a[10]), .Z(n10844) );
  XOR U10942 ( .A(n10849), .B(n10850), .Z(n10763) );
  ANDN U10943 ( .B(n10851), .A(n10852), .Z(n10849) );
  XNOR U10944 ( .A(n10853), .B(n10768), .Z(n10770) );
  XOR U10945 ( .A(n10854), .B(n10855), .Z(n10768) );
  ANDN U10946 ( .B(n10856), .A(n10857), .Z(n10854) );
  AND U10947 ( .A(b[4]), .B(a[11]), .Z(n10853) );
  XNOR U10948 ( .A(n10858), .B(n10859), .Z(n10777) );
  NAND U10949 ( .A(n10860), .B(n10861), .Z(n10859) );
  NAND U10950 ( .A(a[15]), .B(b[0]), .Z(n10695) );
  XNOR U10951 ( .A(n10783), .B(n10784), .Z(c[14]) );
  XOR U10952 ( .A(n10860), .B(n10861), .Z(n10784) );
  XOR U10953 ( .A(n10858), .B(n10862), .Z(n10861) );
  NAND U10954 ( .A(b[1]), .B(a[13]), .Z(n10862) );
  XOR U10955 ( .A(n10858), .B(n10851), .Z(n10863) );
  XNOR U10956 ( .A(n10850), .B(n10856), .Z(n10864) );
  XNOR U10957 ( .A(n10855), .B(n10847), .Z(n10865) );
  XNOR U10958 ( .A(n10846), .B(n10842), .Z(n10866) );
  XNOR U10959 ( .A(n10841), .B(n10837), .Z(n10867) );
  XNOR U10960 ( .A(n10836), .B(n10832), .Z(n10868) );
  XNOR U10961 ( .A(n10823), .B(n10822), .Z(n10869) );
  XOR U10962 ( .A(n10870), .B(n10821), .Z(n10822) );
  AND U10963 ( .A(a[6]), .B(b[8]), .Z(n10870) );
  XNOR U10964 ( .A(n10821), .B(n10827), .Z(n10871) );
  XNOR U10965 ( .A(n10826), .B(n10818), .Z(n10872) );
  XNOR U10966 ( .A(n10817), .B(n10813), .Z(n10873) );
  XNOR U10967 ( .A(n10812), .B(n10808), .Z(n10874) );
  XNOR U10968 ( .A(n10807), .B(n10803), .Z(n10875) );
  XOR U10969 ( .A(n10876), .B(n10802), .Z(n10803) );
  AND U10970 ( .A(a[0]), .B(b[14]), .Z(n10876) );
  XNOR U10971 ( .A(n10877), .B(n10802), .Z(n10804) );
  XNOR U10972 ( .A(n10878), .B(n10879), .Z(n10802) );
  ANDN U10973 ( .B(n10880), .A(n10881), .Z(n10878) );
  AND U10974 ( .A(a[1]), .B(b[13]), .Z(n10877) );
  XNOR U10975 ( .A(n10882), .B(n10807), .Z(n10809) );
  XOR U10976 ( .A(n10883), .B(n10884), .Z(n10807) );
  ANDN U10977 ( .B(n10885), .A(n10886), .Z(n10883) );
  AND U10978 ( .A(a[2]), .B(b[12]), .Z(n10882) );
  XNOR U10979 ( .A(n10887), .B(n10812), .Z(n10814) );
  XOR U10980 ( .A(n10888), .B(n10889), .Z(n10812) );
  ANDN U10981 ( .B(n10890), .A(n10891), .Z(n10888) );
  AND U10982 ( .A(a[3]), .B(b[11]), .Z(n10887) );
  XNOR U10983 ( .A(n10892), .B(n10817), .Z(n10819) );
  XOR U10984 ( .A(n10893), .B(n10894), .Z(n10817) );
  ANDN U10985 ( .B(n10895), .A(n10896), .Z(n10893) );
  AND U10986 ( .A(a[4]), .B(b[10]), .Z(n10892) );
  XOR U10987 ( .A(n10897), .B(n10898), .Z(n10821) );
  AND U10988 ( .A(n10899), .B(n10900), .Z(n10897) );
  XNOR U10989 ( .A(n10901), .B(n10826), .Z(n10828) );
  XOR U10990 ( .A(n10902), .B(n10903), .Z(n10826) );
  ANDN U10991 ( .B(n10904), .A(n10905), .Z(n10902) );
  AND U10992 ( .A(a[5]), .B(b[9]), .Z(n10901) );
  XOR U10993 ( .A(n10906), .B(n10831), .Z(n10833) );
  XOR U10994 ( .A(n10907), .B(n10908), .Z(n10831) );
  ANDN U10995 ( .B(n10909), .A(n10910), .Z(n10907) );
  AND U10996 ( .A(a[7]), .B(b[7]), .Z(n10906) );
  XNOR U10997 ( .A(n10911), .B(n10836), .Z(n10838) );
  XOR U10998 ( .A(n10912), .B(n10913), .Z(n10836) );
  ANDN U10999 ( .B(n10914), .A(n10915), .Z(n10912) );
  AND U11000 ( .A(a[8]), .B(b[6]), .Z(n10911) );
  XNOR U11001 ( .A(n10916), .B(n10841), .Z(n10843) );
  XOR U11002 ( .A(n10917), .B(n10918), .Z(n10841) );
  ANDN U11003 ( .B(n10919), .A(n10920), .Z(n10917) );
  AND U11004 ( .A(a[9]), .B(b[5]), .Z(n10916) );
  XNOR U11005 ( .A(n10921), .B(n10846), .Z(n10848) );
  XOR U11006 ( .A(n10922), .B(n10923), .Z(n10846) );
  ANDN U11007 ( .B(n10924), .A(n10925), .Z(n10922) );
  AND U11008 ( .A(b[4]), .B(a[10]), .Z(n10921) );
  XNOR U11009 ( .A(n10926), .B(n10855), .Z(n10857) );
  XNOR U11010 ( .A(n10927), .B(n10928), .Z(n10855) );
  NOR U11011 ( .A(n10929), .B(n10930), .Z(n10927) );
  AND U11012 ( .A(b[3]), .B(a[11]), .Z(n10926) );
  NANDN U11013 ( .A(n10931), .B(n10932), .Z(n10858) );
  XNOR U11014 ( .A(n10933), .B(n10850), .Z(n10852) );
  XNOR U11015 ( .A(n10934), .B(n10935), .Z(n10850) );
  OR U11016 ( .A(n10936), .B(n10937), .Z(n10935) );
  AND U11017 ( .A(b[2]), .B(a[12]), .Z(n10933) );
  NAND U11018 ( .A(a[14]), .B(b[0]), .Z(n10783) );
  XNOR U11019 ( .A(n10931), .B(n10932), .Z(c[13]) );
  XOR U11020 ( .A(n10937), .B(n10936), .Z(n10932) );
  XOR U11021 ( .A(n10934), .B(n10938), .Z(n10936) );
  NAND U11022 ( .A(b[1]), .B(a[12]), .Z(n10938) );
  XOR U11023 ( .A(n10934), .B(n10930), .Z(n10939) );
  XOR U11024 ( .A(n10940), .B(n10928), .Z(n10930) );
  AND U11025 ( .A(b[2]), .B(a[11]), .Z(n10940) );
  ANDN U11026 ( .B(n10941), .A(n10942), .Z(n10934) );
  XOR U11027 ( .A(n10928), .B(n10924), .Z(n10943) );
  XNOR U11028 ( .A(n10923), .B(n10919), .Z(n10944) );
  XNOR U11029 ( .A(n10918), .B(n10914), .Z(n10945) );
  XNOR U11030 ( .A(n10913), .B(n10909), .Z(n10946) );
  XNOR U11031 ( .A(n10900), .B(n10899), .Z(n10947) );
  XOR U11032 ( .A(n10948), .B(n10898), .Z(n10899) );
  AND U11033 ( .A(a[6]), .B(b[7]), .Z(n10948) );
  XNOR U11034 ( .A(n10898), .B(n10904), .Z(n10949) );
  XNOR U11035 ( .A(n10903), .B(n10895), .Z(n10950) );
  XNOR U11036 ( .A(n10894), .B(n10890), .Z(n10951) );
  XNOR U11037 ( .A(n10889), .B(n10885), .Z(n10952) );
  XNOR U11038 ( .A(n10884), .B(n10880), .Z(n10953) );
  XNOR U11039 ( .A(n10954), .B(n10879), .Z(n10880) );
  AND U11040 ( .A(a[0]), .B(b[13]), .Z(n10954) );
  XOR U11041 ( .A(n10955), .B(n10879), .Z(n10881) );
  XNOR U11042 ( .A(n10956), .B(n10957), .Z(n10879) );
  ANDN U11043 ( .B(n10958), .A(n10959), .Z(n10956) );
  AND U11044 ( .A(a[1]), .B(b[12]), .Z(n10955) );
  XNOR U11045 ( .A(n10960), .B(n10884), .Z(n10886) );
  XOR U11046 ( .A(n10961), .B(n10962), .Z(n10884) );
  ANDN U11047 ( .B(n10963), .A(n10964), .Z(n10961) );
  AND U11048 ( .A(a[2]), .B(b[11]), .Z(n10960) );
  XNOR U11049 ( .A(n10965), .B(n10889), .Z(n10891) );
  XOR U11050 ( .A(n10966), .B(n10967), .Z(n10889) );
  ANDN U11051 ( .B(n10968), .A(n10969), .Z(n10966) );
  AND U11052 ( .A(a[3]), .B(b[10]), .Z(n10965) );
  XNOR U11053 ( .A(n10970), .B(n10894), .Z(n10896) );
  XOR U11054 ( .A(n10971), .B(n10972), .Z(n10894) );
  ANDN U11055 ( .B(n10973), .A(n10974), .Z(n10971) );
  AND U11056 ( .A(a[4]), .B(b[9]), .Z(n10970) );
  XOR U11057 ( .A(n10975), .B(n10976), .Z(n10898) );
  AND U11058 ( .A(n10977), .B(n10978), .Z(n10975) );
  XNOR U11059 ( .A(n10979), .B(n10903), .Z(n10905) );
  XOR U11060 ( .A(n10980), .B(n10981), .Z(n10903) );
  ANDN U11061 ( .B(n10982), .A(n10983), .Z(n10980) );
  AND U11062 ( .A(a[5]), .B(b[8]), .Z(n10979) );
  XOR U11063 ( .A(n10984), .B(n10908), .Z(n10910) );
  XOR U11064 ( .A(n10985), .B(n10986), .Z(n10908) );
  ANDN U11065 ( .B(n10987), .A(n10988), .Z(n10985) );
  AND U11066 ( .A(a[7]), .B(b[6]), .Z(n10984) );
  XNOR U11067 ( .A(n10989), .B(n10913), .Z(n10915) );
  XOR U11068 ( .A(n10990), .B(n10991), .Z(n10913) );
  ANDN U11069 ( .B(n10992), .A(n10993), .Z(n10990) );
  AND U11070 ( .A(a[8]), .B(b[5]), .Z(n10989) );
  XNOR U11071 ( .A(n10994), .B(n10918), .Z(n10920) );
  XOR U11072 ( .A(n10995), .B(n10996), .Z(n10918) );
  ANDN U11073 ( .B(n10997), .A(n10998), .Z(n10995) );
  AND U11074 ( .A(a[9]), .B(b[4]), .Z(n10994) );
  XNOR U11075 ( .A(n10999), .B(n11000), .Z(n10928) );
  NANDN U11076 ( .A(n11001), .B(n11002), .Z(n11000) );
  XNOR U11077 ( .A(n11003), .B(n10923), .Z(n10925) );
  XNOR U11078 ( .A(n11004), .B(n11005), .Z(n10923) );
  AND U11079 ( .A(n11006), .B(n11007), .Z(n11004) );
  AND U11080 ( .A(b[3]), .B(a[10]), .Z(n11003) );
  NAND U11081 ( .A(a[13]), .B(b[0]), .Z(n10931) );
  XNOR U11082 ( .A(n10942), .B(n10941), .Z(c[12]) );
  XNOR U11083 ( .A(n11001), .B(n11002), .Z(n10941) );
  XOR U11084 ( .A(n10999), .B(n11008), .Z(n11002) );
  NAND U11085 ( .A(b[1]), .B(a[11]), .Z(n11008) );
  XOR U11086 ( .A(n11007), .B(n11009), .Z(n11001) );
  XOR U11087 ( .A(n10999), .B(n11006), .Z(n11009) );
  XNOR U11088 ( .A(n11010), .B(n11005), .Z(n11006) );
  AND U11089 ( .A(b[2]), .B(a[10]), .Z(n11010) );
  NANDN U11090 ( .A(n11011), .B(n11012), .Z(n10999) );
  XOR U11091 ( .A(n11005), .B(n10997), .Z(n11013) );
  XNOR U11092 ( .A(n10996), .B(n10992), .Z(n11014) );
  XNOR U11093 ( .A(n10991), .B(n10987), .Z(n11015) );
  XNOR U11094 ( .A(n10978), .B(n10977), .Z(n11016) );
  XOR U11095 ( .A(n11017), .B(n10976), .Z(n10977) );
  AND U11096 ( .A(a[6]), .B(b[6]), .Z(n11017) );
  XNOR U11097 ( .A(n10976), .B(n10982), .Z(n11018) );
  XNOR U11098 ( .A(n10981), .B(n10973), .Z(n11019) );
  XNOR U11099 ( .A(n10972), .B(n10968), .Z(n11020) );
  XNOR U11100 ( .A(n10967), .B(n10963), .Z(n11021) );
  XNOR U11101 ( .A(n10962), .B(n10958), .Z(n11022) );
  XOR U11102 ( .A(n11023), .B(n10957), .Z(n10958) );
  AND U11103 ( .A(a[0]), .B(b[12]), .Z(n11023) );
  XNOR U11104 ( .A(n11024), .B(n10957), .Z(n10959) );
  XNOR U11105 ( .A(n11025), .B(n11026), .Z(n10957) );
  ANDN U11106 ( .B(n11027), .A(n11028), .Z(n11025) );
  AND U11107 ( .A(a[1]), .B(b[11]), .Z(n11024) );
  XNOR U11108 ( .A(n11029), .B(n10962), .Z(n10964) );
  XOR U11109 ( .A(n11030), .B(n11031), .Z(n10962) );
  ANDN U11110 ( .B(n11032), .A(n11033), .Z(n11030) );
  AND U11111 ( .A(a[2]), .B(b[10]), .Z(n11029) );
  XNOR U11112 ( .A(n11034), .B(n10967), .Z(n10969) );
  XOR U11113 ( .A(n11035), .B(n11036), .Z(n10967) );
  ANDN U11114 ( .B(n11037), .A(n11038), .Z(n11035) );
  AND U11115 ( .A(a[3]), .B(b[9]), .Z(n11034) );
  XNOR U11116 ( .A(n11039), .B(n10972), .Z(n10974) );
  XOR U11117 ( .A(n11040), .B(n11041), .Z(n10972) );
  ANDN U11118 ( .B(n11042), .A(n11043), .Z(n11040) );
  AND U11119 ( .A(a[4]), .B(b[8]), .Z(n11039) );
  XOR U11120 ( .A(n11044), .B(n11045), .Z(n10976) );
  AND U11121 ( .A(n11046), .B(n11047), .Z(n11044) );
  XNOR U11122 ( .A(n11048), .B(n10981), .Z(n10983) );
  XOR U11123 ( .A(n11049), .B(n11050), .Z(n10981) );
  ANDN U11124 ( .B(n11051), .A(n11052), .Z(n11049) );
  AND U11125 ( .A(a[5]), .B(b[7]), .Z(n11048) );
  XOR U11126 ( .A(n11053), .B(n10986), .Z(n10988) );
  XOR U11127 ( .A(n11054), .B(n11055), .Z(n10986) );
  ANDN U11128 ( .B(n11056), .A(n11057), .Z(n11054) );
  AND U11129 ( .A(a[7]), .B(b[5]), .Z(n11053) );
  XNOR U11130 ( .A(n11058), .B(n10991), .Z(n10993) );
  XOR U11131 ( .A(n11059), .B(n11060), .Z(n10991) );
  ANDN U11132 ( .B(n11061), .A(n11062), .Z(n11059) );
  AND U11133 ( .A(a[8]), .B(b[4]), .Z(n11058) );
  XNOR U11134 ( .A(n11063), .B(n11064), .Z(n11005) );
  NANDN U11135 ( .A(n11065), .B(n11066), .Z(n11064) );
  XNOR U11136 ( .A(n11067), .B(n10996), .Z(n10998) );
  XNOR U11137 ( .A(n11068), .B(n11069), .Z(n10996) );
  AND U11138 ( .A(n11070), .B(n11071), .Z(n11068) );
  AND U11139 ( .A(a[9]), .B(b[3]), .Z(n11067) );
  NAND U11140 ( .A(a[12]), .B(b[0]), .Z(n10942) );
  XNOR U11141 ( .A(n11011), .B(n11012), .Z(c[11]) );
  XNOR U11142 ( .A(n11065), .B(n11066), .Z(n11012) );
  XOR U11143 ( .A(n11063), .B(n11072), .Z(n11066) );
  NAND U11144 ( .A(b[1]), .B(a[10]), .Z(n11072) );
  XOR U11145 ( .A(n11071), .B(n11073), .Z(n11065) );
  XOR U11146 ( .A(n11063), .B(n11070), .Z(n11073) );
  XNOR U11147 ( .A(n11074), .B(n11069), .Z(n11070) );
  AND U11148 ( .A(a[9]), .B(b[2]), .Z(n11074) );
  NANDN U11149 ( .A(n11075), .B(n11076), .Z(n11063) );
  XOR U11150 ( .A(n11069), .B(n11061), .Z(n11077) );
  XNOR U11151 ( .A(n11060), .B(n11056), .Z(n11078) );
  XNOR U11152 ( .A(n11047), .B(n11046), .Z(n11079) );
  XOR U11153 ( .A(n11080), .B(n11045), .Z(n11046) );
  AND U11154 ( .A(a[6]), .B(b[5]), .Z(n11080) );
  XNOR U11155 ( .A(n11045), .B(n11051), .Z(n11081) );
  XNOR U11156 ( .A(n11050), .B(n11042), .Z(n11082) );
  XNOR U11157 ( .A(n11041), .B(n11037), .Z(n11083) );
  XNOR U11158 ( .A(n11036), .B(n11032), .Z(n11084) );
  XNOR U11159 ( .A(n11031), .B(n11027), .Z(n11085) );
  XNOR U11160 ( .A(n11086), .B(n11026), .Z(n11027) );
  AND U11161 ( .A(a[0]), .B(b[11]), .Z(n11086) );
  XOR U11162 ( .A(n11087), .B(n11026), .Z(n11028) );
  XNOR U11163 ( .A(n11088), .B(n11089), .Z(n11026) );
  ANDN U11164 ( .B(n11090), .A(n11091), .Z(n11088) );
  AND U11165 ( .A(a[1]), .B(b[10]), .Z(n11087) );
  XNOR U11166 ( .A(n11092), .B(n11031), .Z(n11033) );
  XOR U11167 ( .A(n11093), .B(n11094), .Z(n11031) );
  ANDN U11168 ( .B(n11095), .A(n11096), .Z(n11093) );
  AND U11169 ( .A(a[2]), .B(b[9]), .Z(n11092) );
  XNOR U11170 ( .A(n11097), .B(n11036), .Z(n11038) );
  XOR U11171 ( .A(n11098), .B(n11099), .Z(n11036) );
  ANDN U11172 ( .B(n11100), .A(n11101), .Z(n11098) );
  AND U11173 ( .A(a[3]), .B(b[8]), .Z(n11097) );
  XNOR U11174 ( .A(n11102), .B(n11041), .Z(n11043) );
  XOR U11175 ( .A(n11103), .B(n11104), .Z(n11041) );
  ANDN U11176 ( .B(n11105), .A(n11106), .Z(n11103) );
  AND U11177 ( .A(a[4]), .B(b[7]), .Z(n11102) );
  XNOR U11178 ( .A(n11107), .B(n11108), .Z(n11045) );
  ANDN U11179 ( .B(n11109), .A(n11110), .Z(n11107) );
  XNOR U11180 ( .A(n11111), .B(n11050), .Z(n11052) );
  XOR U11181 ( .A(n11112), .B(n11113), .Z(n11050) );
  ANDN U11182 ( .B(n11114), .A(n11115), .Z(n11112) );
  AND U11183 ( .A(a[5]), .B(b[6]), .Z(n11111) );
  XOR U11184 ( .A(n11116), .B(n11055), .Z(n11057) );
  XOR U11185 ( .A(n11117), .B(n11118), .Z(n11055) );
  ANDN U11186 ( .B(n11119), .A(n11120), .Z(n11117) );
  AND U11187 ( .A(a[7]), .B(b[4]), .Z(n11116) );
  XNOR U11188 ( .A(n11121), .B(n11122), .Z(n11069) );
  NANDN U11189 ( .A(n11123), .B(n11124), .Z(n11122) );
  XNOR U11190 ( .A(n11125), .B(n11060), .Z(n11062) );
  XNOR U11191 ( .A(n11126), .B(n11127), .Z(n11060) );
  AND U11192 ( .A(n11128), .B(n11129), .Z(n11126) );
  AND U11193 ( .A(a[8]), .B(b[3]), .Z(n11125) );
  NAND U11194 ( .A(a[11]), .B(b[0]), .Z(n11011) );
  XNOR U11195 ( .A(n11075), .B(n11076), .Z(c[10]) );
  XNOR U11196 ( .A(n11123), .B(n11124), .Z(n11076) );
  XOR U11197 ( .A(n11121), .B(n11130), .Z(n11124) );
  NAND U11198 ( .A(a[9]), .B(b[1]), .Z(n11130) );
  XOR U11199 ( .A(n11129), .B(n11131), .Z(n11123) );
  XOR U11200 ( .A(n11121), .B(n11128), .Z(n11131) );
  XNOR U11201 ( .A(n11132), .B(n11127), .Z(n11128) );
  AND U11202 ( .A(a[8]), .B(b[2]), .Z(n11132) );
  OR U11203 ( .A(n1), .B(n2), .Z(n11121) );
  XOR U11204 ( .A(n11133), .B(n11134), .Z(n2) );
  NAND U11205 ( .A(b[0]), .B(a[9]), .Z(n1) );
  XOR U11206 ( .A(n11127), .B(n11119), .Z(n11135) );
  XNOR U11207 ( .A(n11136), .B(n11137), .Z(n11119) );
  XOR U11208 ( .A(n11109), .B(n11110), .Z(n11137) );
  XOR U11209 ( .A(n11138), .B(n11108), .Z(n11110) );
  AND U11210 ( .A(a[6]), .B(b[4]), .Z(n11138) );
  XOR U11211 ( .A(n11108), .B(n11114), .Z(n11139) );
  XNOR U11212 ( .A(n11113), .B(n11105), .Z(n11140) );
  XNOR U11213 ( .A(n11104), .B(n11100), .Z(n11141) );
  XNOR U11214 ( .A(n11099), .B(n11095), .Z(n11142) );
  XNOR U11215 ( .A(n11094), .B(n11090), .Z(n11143) );
  XOR U11216 ( .A(n11144), .B(n11089), .Z(n11090) );
  AND U11217 ( .A(a[0]), .B(b[10]), .Z(n11144) );
  XNOR U11218 ( .A(n11145), .B(n11089), .Z(n11091) );
  XNOR U11219 ( .A(n11146), .B(n11147), .Z(n11089) );
  ANDN U11220 ( .B(n11148), .A(n11149), .Z(n11146) );
  AND U11221 ( .A(a[1]), .B(b[9]), .Z(n11145) );
  XNOR U11222 ( .A(n11150), .B(n11094), .Z(n11096) );
  XNOR U11223 ( .A(n11151), .B(n11152), .Z(n11094) );
  ANDN U11224 ( .B(n11153), .A(n11154), .Z(n11151) );
  AND U11225 ( .A(a[2]), .B(b[8]), .Z(n11150) );
  XNOR U11226 ( .A(n11155), .B(n11099), .Z(n11101) );
  XNOR U11227 ( .A(n11156), .B(n11157), .Z(n11099) );
  ANDN U11228 ( .B(n11158), .A(n11159), .Z(n11156) );
  AND U11229 ( .A(a[3]), .B(b[7]), .Z(n11155) );
  XNOR U11230 ( .A(n11160), .B(n11104), .Z(n11106) );
  XNOR U11231 ( .A(n11161), .B(n11162), .Z(n11104) );
  ANDN U11232 ( .B(n11163), .A(n11164), .Z(n11161) );
  AND U11233 ( .A(a[4]), .B(b[6]), .Z(n11160) );
  XOR U11234 ( .A(n11165), .B(n11166), .Z(n11108) );
  ANDN U11235 ( .B(n11167), .A(n11168), .Z(n11165) );
  XNOR U11236 ( .A(n11169), .B(n11113), .Z(n11115) );
  XNOR U11237 ( .A(n11170), .B(n11171), .Z(n11113) );
  ANDN U11238 ( .B(n11172), .A(n11173), .Z(n11170) );
  AND U11239 ( .A(a[5]), .B(b[5]), .Z(n11169) );
  XNOR U11240 ( .A(n11174), .B(n11175), .Z(n11127) );
  NANDN U11241 ( .A(n11134), .B(n11133), .Z(n11175) );
  XOR U11242 ( .A(n11174), .B(n11176), .Z(n11133) );
  NAND U11243 ( .A(a[8]), .B(b[1]), .Z(n11176) );
  XOR U11244 ( .A(n11174), .B(n11178), .Z(n11177) );
  NANDN U11245 ( .A(n3), .B(n4), .Z(n11174) );
  XOR U11246 ( .A(n11180), .B(n11181), .Z(n4) );
  NAND U11247 ( .A(a[8]), .B(b[0]), .Z(n3) );
  XOR U11248 ( .A(n11182), .B(n11118), .Z(n11120) );
  IV U11249 ( .A(n11136), .Z(n11118) );
  XOR U11250 ( .A(n11183), .B(n11184), .Z(n11136) );
  ANDN U11251 ( .B(n11178), .A(n11179), .Z(n11183) );
  AND U11252 ( .A(a[7]), .B(b[2]), .Z(n11185) );
  XNOR U11253 ( .A(n11167), .B(n11184), .Z(n11186) );
  XOR U11254 ( .A(n11187), .B(n11188), .Z(n11184) );
  OR U11255 ( .A(n11180), .B(n11181), .Z(n11188) );
  XNOR U11256 ( .A(n11190), .B(n11191), .Z(n11189) );
  XOR U11257 ( .A(n11190), .B(n11193), .Z(n11180) );
  NAND U11258 ( .A(a[7]), .B(b[1]), .Z(n11193) );
  IV U11259 ( .A(n11187), .Z(n11190) );
  NANDN U11260 ( .A(n5), .B(n6), .Z(n11187) );
  XOR U11261 ( .A(n11194), .B(n11195), .Z(n6) );
  NAND U11262 ( .A(a[7]), .B(b[0]), .Z(n5) );
  XNOR U11263 ( .A(n11172), .B(n11197), .Z(n11196) );
  XNOR U11264 ( .A(n11163), .B(n11199), .Z(n11198) );
  XNOR U11265 ( .A(n11158), .B(n11201), .Z(n11200) );
  XNOR U11266 ( .A(n11153), .B(n11203), .Z(n11202) );
  XNOR U11267 ( .A(n11148), .B(n11205), .Z(n11204) );
  XNOR U11268 ( .A(n11206), .B(n11147), .Z(n11148) );
  AND U11269 ( .A(a[0]), .B(b[9]), .Z(n11206) );
  XOR U11270 ( .A(n11207), .B(n11147), .Z(n11149) );
  XNOR U11271 ( .A(n11208), .B(n11209), .Z(n11147) );
  ANDN U11272 ( .B(n11210), .A(n11211), .Z(n11208) );
  AND U11273 ( .A(a[1]), .B(b[8]), .Z(n11207) );
  XOR U11274 ( .A(n11212), .B(n11152), .Z(n11154) );
  IV U11275 ( .A(n11205), .Z(n11152) );
  XOR U11276 ( .A(n11213), .B(n11214), .Z(n11205) );
  ANDN U11277 ( .B(n11215), .A(n11216), .Z(n11213) );
  AND U11278 ( .A(a[2]), .B(b[7]), .Z(n11212) );
  XOR U11279 ( .A(n11217), .B(n11157), .Z(n11159) );
  IV U11280 ( .A(n11203), .Z(n11157) );
  XOR U11281 ( .A(n11218), .B(n11219), .Z(n11203) );
  ANDN U11282 ( .B(n11220), .A(n11221), .Z(n11218) );
  AND U11283 ( .A(a[3]), .B(b[6]), .Z(n11217) );
  XOR U11284 ( .A(n11222), .B(n11162), .Z(n11164) );
  IV U11285 ( .A(n11201), .Z(n11162) );
  XOR U11286 ( .A(n11223), .B(n11224), .Z(n11201) );
  ANDN U11287 ( .B(n11225), .A(n11226), .Z(n11223) );
  AND U11288 ( .A(a[4]), .B(b[5]), .Z(n11222) );
  XOR U11289 ( .A(n11227), .B(n11171), .Z(n11173) );
  IV U11290 ( .A(n11199), .Z(n11171) );
  XOR U11291 ( .A(n11228), .B(n11229), .Z(n11199) );
  ANDN U11292 ( .B(n11230), .A(n11231), .Z(n11228) );
  AND U11293 ( .A(a[5]), .B(b[4]), .Z(n11227) );
  XOR U11294 ( .A(n11232), .B(n11166), .Z(n11168) );
  IV U11295 ( .A(n11197), .Z(n11166) );
  XOR U11296 ( .A(n11233), .B(n11234), .Z(n11197) );
  ANDN U11297 ( .B(n11191), .A(n11192), .Z(n11233) );
  AND U11298 ( .A(a[6]), .B(b[2]), .Z(n11235) );
  XNOR U11299 ( .A(n11230), .B(n11234), .Z(n11236) );
  XOR U11300 ( .A(n11237), .B(n11238), .Z(n11234) );
  OR U11301 ( .A(n11194), .B(n11195), .Z(n11238) );
  XNOR U11302 ( .A(n11240), .B(n11241), .Z(n11239) );
  XOR U11303 ( .A(n11240), .B(n11243), .Z(n11194) );
  NAND U11304 ( .A(a[6]), .B(b[1]), .Z(n11243) );
  IV U11305 ( .A(n11237), .Z(n11240) );
  NANDN U11306 ( .A(n7), .B(n8), .Z(n11237) );
  XOR U11307 ( .A(n11244), .B(n11245), .Z(n8) );
  NAND U11308 ( .A(a[6]), .B(b[0]), .Z(n7) );
  XNOR U11309 ( .A(n11225), .B(n11229), .Z(n11246) );
  XNOR U11310 ( .A(n11220), .B(n11224), .Z(n11247) );
  XNOR U11311 ( .A(n11215), .B(n11219), .Z(n11248) );
  XNOR U11312 ( .A(n11210), .B(n11214), .Z(n11249) );
  XOR U11313 ( .A(n11250), .B(n11209), .Z(n11210) );
  AND U11314 ( .A(a[0]), .B(b[8]), .Z(n11250) );
  XNOR U11315 ( .A(n11251), .B(n11209), .Z(n11211) );
  XNOR U11316 ( .A(n11252), .B(n11253), .Z(n11209) );
  ANDN U11317 ( .B(n11254), .A(n11255), .Z(n11252) );
  AND U11318 ( .A(a[1]), .B(b[7]), .Z(n11251) );
  XOR U11319 ( .A(n11257), .B(n11258), .Z(n11214) );
  ANDN U11320 ( .B(n11259), .A(n11260), .Z(n11257) );
  AND U11321 ( .A(a[2]), .B(b[6]), .Z(n11256) );
  XOR U11322 ( .A(n11262), .B(n11263), .Z(n11219) );
  ANDN U11323 ( .B(n11264), .A(n11265), .Z(n11262) );
  AND U11324 ( .A(a[3]), .B(b[5]), .Z(n11261) );
  XOR U11325 ( .A(n11267), .B(n11268), .Z(n11224) );
  ANDN U11326 ( .B(n11269), .A(n11270), .Z(n11267) );
  AND U11327 ( .A(a[4]), .B(b[4]), .Z(n11266) );
  XOR U11328 ( .A(n11272), .B(n11273), .Z(n11229) );
  ANDN U11329 ( .B(n11241), .A(n11242), .Z(n11272) );
  AND U11330 ( .A(a[5]), .B(b[2]), .Z(n11274) );
  XNOR U11331 ( .A(n11269), .B(n11273), .Z(n11275) );
  XOR U11332 ( .A(n11276), .B(n11277), .Z(n11273) );
  OR U11333 ( .A(n11244), .B(n11245), .Z(n11277) );
  XNOR U11334 ( .A(n11279), .B(n11280), .Z(n11278) );
  XOR U11335 ( .A(n11279), .B(n11282), .Z(n11244) );
  NAND U11336 ( .A(a[5]), .B(b[1]), .Z(n11282) );
  IV U11337 ( .A(n11276), .Z(n11279) );
  NANDN U11338 ( .A(n1211), .B(n1212), .Z(n11276) );
  XOR U11339 ( .A(n11283), .B(n11284), .Z(n1212) );
  NAND U11340 ( .A(a[5]), .B(b[0]), .Z(n1211) );
  XNOR U11341 ( .A(n11264), .B(n11268), .Z(n11285) );
  XNOR U11342 ( .A(n11259), .B(n11263), .Z(n11286) );
  XNOR U11343 ( .A(n11254), .B(n11258), .Z(n11287) );
  XNOR U11344 ( .A(n11288), .B(n11253), .Z(n11254) );
  AND U11345 ( .A(a[0]), .B(b[7]), .Z(n11288) );
  XOR U11346 ( .A(n11289), .B(n11253), .Z(n11255) );
  XNOR U11347 ( .A(n11290), .B(n11291), .Z(n11253) );
  ANDN U11348 ( .B(n11292), .A(n11293), .Z(n11290) );
  AND U11349 ( .A(a[1]), .B(b[6]), .Z(n11289) );
  XOR U11350 ( .A(n11295), .B(n11296), .Z(n11258) );
  ANDN U11351 ( .B(n11297), .A(n11298), .Z(n11295) );
  AND U11352 ( .A(a[2]), .B(b[5]), .Z(n11294) );
  XOR U11353 ( .A(n11300), .B(n11301), .Z(n11263) );
  ANDN U11354 ( .B(n11302), .A(n11303), .Z(n11300) );
  AND U11355 ( .A(a[3]), .B(b[4]), .Z(n11299) );
  XOR U11356 ( .A(n11305), .B(n11306), .Z(n11268) );
  ANDN U11357 ( .B(n11280), .A(n11281), .Z(n11305) );
  AND U11358 ( .A(a[4]), .B(b[2]), .Z(n11307) );
  XNOR U11359 ( .A(n11302), .B(n11306), .Z(n11308) );
  XOR U11360 ( .A(n11309), .B(n11310), .Z(n11306) );
  OR U11361 ( .A(n11283), .B(n11284), .Z(n11310) );
  XNOR U11362 ( .A(n11312), .B(n11313), .Z(n11311) );
  XOR U11363 ( .A(n11312), .B(n11315), .Z(n11283) );
  NAND U11364 ( .A(a[4]), .B(b[1]), .Z(n11315) );
  IV U11365 ( .A(n11309), .Z(n11312) );
  NANDN U11366 ( .A(n4409), .B(n4410), .Z(n11309) );
  XOR U11367 ( .A(n11316), .B(n11317), .Z(n4410) );
  NAND U11368 ( .A(a[4]), .B(b[0]), .Z(n4409) );
  XNOR U11369 ( .A(n11297), .B(n11301), .Z(n11318) );
  XNOR U11370 ( .A(n11292), .B(n11296), .Z(n11319) );
  XOR U11371 ( .A(n11320), .B(n11291), .Z(n11292) );
  AND U11372 ( .A(a[0]), .B(b[6]), .Z(n11320) );
  XNOR U11373 ( .A(n11321), .B(n11291), .Z(n11293) );
  XNOR U11374 ( .A(n11322), .B(n11323), .Z(n11291) );
  ANDN U11375 ( .B(n11324), .A(n11325), .Z(n11322) );
  AND U11376 ( .A(a[1]), .B(b[5]), .Z(n11321) );
  XOR U11377 ( .A(n11327), .B(n11328), .Z(n11296) );
  ANDN U11378 ( .B(n11329), .A(n11330), .Z(n11327) );
  AND U11379 ( .A(a[2]), .B(b[4]), .Z(n11326) );
  XOR U11380 ( .A(n11332), .B(n11333), .Z(n11301) );
  ANDN U11381 ( .B(n11313), .A(n11314), .Z(n11332) );
  AND U11382 ( .A(a[3]), .B(b[2]), .Z(n11334) );
  XNOR U11383 ( .A(n11329), .B(n11333), .Z(n11335) );
  XOR U11384 ( .A(n11336), .B(n11337), .Z(n11333) );
  OR U11385 ( .A(n11316), .B(n11317), .Z(n11337) );
  XNOR U11386 ( .A(n11339), .B(n11340), .Z(n11338) );
  XOR U11387 ( .A(n11339), .B(n11342), .Z(n11316) );
  NAND U11388 ( .A(a[3]), .B(b[1]), .Z(n11342) );
  IV U11389 ( .A(n11336), .Z(n11339) );
  NANDN U11390 ( .A(n7006), .B(n7007), .Z(n11336) );
  XOR U11391 ( .A(n11343), .B(n11344), .Z(n7007) );
  NAND U11392 ( .A(a[3]), .B(b[0]), .Z(n7006) );
  XNOR U11393 ( .A(n11324), .B(n11328), .Z(n11345) );
  XNOR U11394 ( .A(n11346), .B(n11323), .Z(n11324) );
  AND U11395 ( .A(a[0]), .B(b[5]), .Z(n11346) );
  XOR U11396 ( .A(n11347), .B(n11323), .Z(n11325) );
  XNOR U11397 ( .A(n11348), .B(n11349), .Z(n11323) );
  ANDN U11398 ( .B(n11350), .A(n11351), .Z(n11348) );
  AND U11399 ( .A(a[1]), .B(b[4]), .Z(n11347) );
  XOR U11400 ( .A(n11353), .B(n11354), .Z(n11328) );
  ANDN U11401 ( .B(n11340), .A(n11341), .Z(n11353) );
  AND U11402 ( .A(a[2]), .B(b[2]), .Z(n11355) );
  XNOR U11403 ( .A(n11350), .B(n11354), .Z(n11356) );
  XOR U11404 ( .A(n11357), .B(n11358), .Z(n11354) );
  OR U11405 ( .A(n11343), .B(n11344), .Z(n11358) );
  XNOR U11406 ( .A(n11360), .B(n11361), .Z(n11359) );
  XOR U11407 ( .A(n11360), .B(n11363), .Z(n11343) );
  NAND U11408 ( .A(a[2]), .B(b[1]), .Z(n11363) );
  IV U11409 ( .A(n11357), .Z(n11360) );
  NANDN U11410 ( .A(n8998), .B(n8999), .Z(n11357) );
  XOR U11411 ( .A(n11364), .B(n11365), .Z(n8999) );
  NAND U11412 ( .A(a[2]), .B(b[0]), .Z(n8998) );
  XOR U11413 ( .A(n11366), .B(n11349), .Z(n11350) );
  AND U11414 ( .A(a[0]), .B(b[4]), .Z(n11366) );
  XNOR U11415 ( .A(n11367), .B(n11349), .Z(n11351) );
  XNOR U11416 ( .A(n11368), .B(n11369), .Z(n11349) );
  ANDN U11417 ( .B(n11361), .A(n11362), .Z(n11368) );
  XOR U11418 ( .A(n11370), .B(n11369), .Z(n11362) );
  AND U11419 ( .A(a[1]), .B(b[2]), .Z(n11370) );
  XNOR U11420 ( .A(n11371), .B(n11369), .Z(n11361) );
  XNOR U11421 ( .A(n11372), .B(n11373), .Z(n11369) );
  OR U11422 ( .A(n11365), .B(n11364), .Z(n11373) );
  XNOR U11423 ( .A(n11372), .B(n11374), .Z(n11364) );
  NAND U11424 ( .A(a[1]), .B(b[1]), .Z(n11374) );
  XNOR U11425 ( .A(n11372), .B(n11375), .Z(n11365) );
  NAND U11426 ( .A(a[0]), .B(b[2]), .Z(n11375) );
  OR U11427 ( .A(n10390), .B(n10391), .Z(n11372) );
  NAND U11428 ( .A(b[1]), .B(a[0]), .Z(n10391) );
  NAND U11429 ( .A(a[1]), .B(b[0]), .Z(n10390) );
  AND U11430 ( .A(a[0]), .B(b[3]), .Z(n11371) );
  AND U11431 ( .A(a[1]), .B(b[3]), .Z(n11367) );
  AND U11432 ( .A(a[2]), .B(b[3]), .Z(n11352) );
  AND U11433 ( .A(a[3]), .B(b[3]), .Z(n11331) );
  AND U11434 ( .A(a[4]), .B(b[3]), .Z(n11304) );
  AND U11435 ( .A(a[5]), .B(b[3]), .Z(n11271) );
  AND U11436 ( .A(a[6]), .B(b[3]), .Z(n11232) );
  AND U11437 ( .A(a[7]), .B(b[3]), .Z(n11182) );
  NAND U11438 ( .A(a[10]), .B(b[0]), .Z(n11075) );
  AND U11439 ( .A(b[0]), .B(a[0]), .Z(c[0]) );
endmodule

