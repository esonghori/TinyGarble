module SubBytes(
x,
z);

	input [127:0] x;
	output [127:0] z;
	wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439;

	assign {w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127} = x;

	assign z = {w331, w332, w327, w321, w333, w322, w334, w324, w538, w539, w534, w528, w540, w529, w541, w531, w745, w746, w741, w735, w747, w736, w748, w738, w952, w953, w948, w942, w954, w943, w955, w945, w1159, w1160, w1155, w1149, w1161, w1150, w1162, w1152, w1366, w1367, w1362, w1356, w1368, w1357, w1369, w1359, w1573, w1574, w1569, w1563, w1575, w1564, w1576, w1566, w1780, w1781, w1776, w1770, w1782, w1771, w1783, w1773, w1987, w1988, w1983, w1977, w1989, w1978, w1990, w1980, w2194, w2195, w2190, w2184, w2196, w2185, w2197, w2187, w2401, w2402, w2397, w2391, w2403, w2392, w2404, w2394, w2608, w2609, w2604, w2598, w2610, w2599, w2611, w2601, w2815, w2816, w2811, w2805, w2817, w2806, w2818, w2808, w3022, w3023, w3018, w3012, w3024, w3013, w3025, w3015, w3229, w3230, w3225, w3219, w3231, w3220, w3232, w3222, w3436, w3437, w3432, w3426, w3438, w3427, w3439, w3429};

	wire w128;
	assign w128 = 1'b0;
	wire w129;
	assign w129 = 1'b0;
	wire w130;
	assign w130 = 1'b0;
	wire w131;
	assign w131 = 1'b0;
	wire w132;
	assign w132 = 1'b0;
	wire w133;
	assign w133 = 1'b0;
	wire w134;
	assign w134 = 1'b0;
	wire w135;
	assign w135 = 1'b0;
	wire w301;
	assign w301 = 1'b1;
	wire w302;
	assign w302 = 1'b1;
	wire w303;
	assign w303 = 1'b1;
	wire w304;
	assign w304 = 1'b1;
	wire w305;
	assign w305 = 1'b1;
	wire w306;
	assign w306 = 1'b1;
	wire w307;
	assign w307 = 1'b1;
	wire w308;
	assign w308 = 1'b1;
	wire w335;
	assign w335 = 1'b0;
	wire w336;
	assign w336 = 1'b0;
	wire w337;
	assign w337 = 1'b0;
	wire w338;
	assign w338 = 1'b0;
	wire w339;
	assign w339 = 1'b0;
	wire w340;
	assign w340 = 1'b0;
	wire w341;
	assign w341 = 1'b0;
	wire w342;
	assign w342 = 1'b0;
	wire w508;
	assign w508 = 1'b1;
	wire w509;
	assign w509 = 1'b1;
	wire w510;
	assign w510 = 1'b1;
	wire w511;
	assign w511 = 1'b1;
	wire w512;
	assign w512 = 1'b1;
	wire w513;
	assign w513 = 1'b1;
	wire w514;
	assign w514 = 1'b1;
	wire w515;
	assign w515 = 1'b1;
	wire w542;
	assign w542 = 1'b0;
	wire w543;
	assign w543 = 1'b0;
	wire w544;
	assign w544 = 1'b0;
	wire w545;
	assign w545 = 1'b0;
	wire w546;
	assign w546 = 1'b0;
	wire w547;
	assign w547 = 1'b0;
	wire w548;
	assign w548 = 1'b0;
	wire w549;
	assign w549 = 1'b0;
	wire w715;
	assign w715 = 1'b1;
	wire w716;
	assign w716 = 1'b1;
	wire w717;
	assign w717 = 1'b1;
	wire w718;
	assign w718 = 1'b1;
	wire w719;
	assign w719 = 1'b1;
	wire w720;
	assign w720 = 1'b1;
	wire w721;
	assign w721 = 1'b1;
	wire w722;
	assign w722 = 1'b1;
	wire w749;
	assign w749 = 1'b0;
	wire w750;
	assign w750 = 1'b0;
	wire w751;
	assign w751 = 1'b0;
	wire w752;
	assign w752 = 1'b0;
	wire w753;
	assign w753 = 1'b0;
	wire w754;
	assign w754 = 1'b0;
	wire w755;
	assign w755 = 1'b0;
	wire w756;
	assign w756 = 1'b0;
	wire w922;
	assign w922 = 1'b1;
	wire w923;
	assign w923 = 1'b1;
	wire w924;
	assign w924 = 1'b1;
	wire w925;
	assign w925 = 1'b1;
	wire w926;
	assign w926 = 1'b1;
	wire w927;
	assign w927 = 1'b1;
	wire w928;
	assign w928 = 1'b1;
	wire w929;
	assign w929 = 1'b1;
	wire w956;
	assign w956 = 1'b0;
	wire w957;
	assign w957 = 1'b0;
	wire w958;
	assign w958 = 1'b0;
	wire w959;
	assign w959 = 1'b0;
	wire w960;
	assign w960 = 1'b0;
	wire w961;
	assign w961 = 1'b0;
	wire w962;
	assign w962 = 1'b0;
	wire w963;
	assign w963 = 1'b0;
	wire w1129;
	assign w1129 = 1'b1;
	wire w1130;
	assign w1130 = 1'b1;
	wire w1131;
	assign w1131 = 1'b1;
	wire w1132;
	assign w1132 = 1'b1;
	wire w1133;
	assign w1133 = 1'b1;
	wire w1134;
	assign w1134 = 1'b1;
	wire w1135;
	assign w1135 = 1'b1;
	wire w1136;
	assign w1136 = 1'b1;
	wire w1163;
	assign w1163 = 1'b0;
	wire w1164;
	assign w1164 = 1'b0;
	wire w1165;
	assign w1165 = 1'b0;
	wire w1166;
	assign w1166 = 1'b0;
	wire w1167;
	assign w1167 = 1'b0;
	wire w1168;
	assign w1168 = 1'b0;
	wire w1169;
	assign w1169 = 1'b0;
	wire w1170;
	assign w1170 = 1'b0;
	wire w1336;
	assign w1336 = 1'b1;
	wire w1337;
	assign w1337 = 1'b1;
	wire w1338;
	assign w1338 = 1'b1;
	wire w1339;
	assign w1339 = 1'b1;
	wire w1340;
	assign w1340 = 1'b1;
	wire w1341;
	assign w1341 = 1'b1;
	wire w1342;
	assign w1342 = 1'b1;
	wire w1343;
	assign w1343 = 1'b1;
	wire w1370;
	assign w1370 = 1'b0;
	wire w1371;
	assign w1371 = 1'b0;
	wire w1372;
	assign w1372 = 1'b0;
	wire w1373;
	assign w1373 = 1'b0;
	wire w1374;
	assign w1374 = 1'b0;
	wire w1375;
	assign w1375 = 1'b0;
	wire w1376;
	assign w1376 = 1'b0;
	wire w1377;
	assign w1377 = 1'b0;
	wire w1543;
	assign w1543 = 1'b1;
	wire w1544;
	assign w1544 = 1'b1;
	wire w1545;
	assign w1545 = 1'b1;
	wire w1546;
	assign w1546 = 1'b1;
	wire w1547;
	assign w1547 = 1'b1;
	wire w1548;
	assign w1548 = 1'b1;
	wire w1549;
	assign w1549 = 1'b1;
	wire w1550;
	assign w1550 = 1'b1;
	wire w1577;
	assign w1577 = 1'b0;
	wire w1578;
	assign w1578 = 1'b0;
	wire w1579;
	assign w1579 = 1'b0;
	wire w1580;
	assign w1580 = 1'b0;
	wire w1581;
	assign w1581 = 1'b0;
	wire w1582;
	assign w1582 = 1'b0;
	wire w1583;
	assign w1583 = 1'b0;
	wire w1584;
	assign w1584 = 1'b0;
	wire w1750;
	assign w1750 = 1'b1;
	wire w1751;
	assign w1751 = 1'b1;
	wire w1752;
	assign w1752 = 1'b1;
	wire w1753;
	assign w1753 = 1'b1;
	wire w1754;
	assign w1754 = 1'b1;
	wire w1755;
	assign w1755 = 1'b1;
	wire w1756;
	assign w1756 = 1'b1;
	wire w1757;
	assign w1757 = 1'b1;
	wire w1784;
	assign w1784 = 1'b0;
	wire w1785;
	assign w1785 = 1'b0;
	wire w1786;
	assign w1786 = 1'b0;
	wire w1787;
	assign w1787 = 1'b0;
	wire w1788;
	assign w1788 = 1'b0;
	wire w1789;
	assign w1789 = 1'b0;
	wire w1790;
	assign w1790 = 1'b0;
	wire w1791;
	assign w1791 = 1'b0;
	wire w1957;
	assign w1957 = 1'b1;
	wire w1958;
	assign w1958 = 1'b1;
	wire w1959;
	assign w1959 = 1'b1;
	wire w1960;
	assign w1960 = 1'b1;
	wire w1961;
	assign w1961 = 1'b1;
	wire w1962;
	assign w1962 = 1'b1;
	wire w1963;
	assign w1963 = 1'b1;
	wire w1964;
	assign w1964 = 1'b1;
	wire w1991;
	assign w1991 = 1'b0;
	wire w1992;
	assign w1992 = 1'b0;
	wire w1993;
	assign w1993 = 1'b0;
	wire w1994;
	assign w1994 = 1'b0;
	wire w1995;
	assign w1995 = 1'b0;
	wire w1996;
	assign w1996 = 1'b0;
	wire w1997;
	assign w1997 = 1'b0;
	wire w1998;
	assign w1998 = 1'b0;
	wire w2164;
	assign w2164 = 1'b1;
	wire w2165;
	assign w2165 = 1'b1;
	wire w2166;
	assign w2166 = 1'b1;
	wire w2167;
	assign w2167 = 1'b1;
	wire w2168;
	assign w2168 = 1'b1;
	wire w2169;
	assign w2169 = 1'b1;
	wire w2170;
	assign w2170 = 1'b1;
	wire w2171;
	assign w2171 = 1'b1;
	wire w2198;
	assign w2198 = 1'b0;
	wire w2199;
	assign w2199 = 1'b0;
	wire w2200;
	assign w2200 = 1'b0;
	wire w2201;
	assign w2201 = 1'b0;
	wire w2202;
	assign w2202 = 1'b0;
	wire w2203;
	assign w2203 = 1'b0;
	wire w2204;
	assign w2204 = 1'b0;
	wire w2205;
	assign w2205 = 1'b0;
	wire w2371;
	assign w2371 = 1'b1;
	wire w2372;
	assign w2372 = 1'b1;
	wire w2373;
	assign w2373 = 1'b1;
	wire w2374;
	assign w2374 = 1'b1;
	wire w2375;
	assign w2375 = 1'b1;
	wire w2376;
	assign w2376 = 1'b1;
	wire w2377;
	assign w2377 = 1'b1;
	wire w2378;
	assign w2378 = 1'b1;
	wire w2405;
	assign w2405 = 1'b0;
	wire w2406;
	assign w2406 = 1'b0;
	wire w2407;
	assign w2407 = 1'b0;
	wire w2408;
	assign w2408 = 1'b0;
	wire w2409;
	assign w2409 = 1'b0;
	wire w2410;
	assign w2410 = 1'b0;
	wire w2411;
	assign w2411 = 1'b0;
	wire w2412;
	assign w2412 = 1'b0;
	wire w2578;
	assign w2578 = 1'b1;
	wire w2579;
	assign w2579 = 1'b1;
	wire w2580;
	assign w2580 = 1'b1;
	wire w2581;
	assign w2581 = 1'b1;
	wire w2582;
	assign w2582 = 1'b1;
	wire w2583;
	assign w2583 = 1'b1;
	wire w2584;
	assign w2584 = 1'b1;
	wire w2585;
	assign w2585 = 1'b1;
	wire w2612;
	assign w2612 = 1'b0;
	wire w2613;
	assign w2613 = 1'b0;
	wire w2614;
	assign w2614 = 1'b0;
	wire w2615;
	assign w2615 = 1'b0;
	wire w2616;
	assign w2616 = 1'b0;
	wire w2617;
	assign w2617 = 1'b0;
	wire w2618;
	assign w2618 = 1'b0;
	wire w2619;
	assign w2619 = 1'b0;
	wire w2785;
	assign w2785 = 1'b1;
	wire w2786;
	assign w2786 = 1'b1;
	wire w2787;
	assign w2787 = 1'b1;
	wire w2788;
	assign w2788 = 1'b1;
	wire w2789;
	assign w2789 = 1'b1;
	wire w2790;
	assign w2790 = 1'b1;
	wire w2791;
	assign w2791 = 1'b1;
	wire w2792;
	assign w2792 = 1'b1;
	wire w2819;
	assign w2819 = 1'b0;
	wire w2820;
	assign w2820 = 1'b0;
	wire w2821;
	assign w2821 = 1'b0;
	wire w2822;
	assign w2822 = 1'b0;
	wire w2823;
	assign w2823 = 1'b0;
	wire w2824;
	assign w2824 = 1'b0;
	wire w2825;
	assign w2825 = 1'b0;
	wire w2826;
	assign w2826 = 1'b0;
	wire w2992;
	assign w2992 = 1'b1;
	wire w2993;
	assign w2993 = 1'b1;
	wire w2994;
	assign w2994 = 1'b1;
	wire w2995;
	assign w2995 = 1'b1;
	wire w2996;
	assign w2996 = 1'b1;
	wire w2997;
	assign w2997 = 1'b1;
	wire w2998;
	assign w2998 = 1'b1;
	wire w2999;
	assign w2999 = 1'b1;
	wire w3026;
	assign w3026 = 1'b0;
	wire w3027;
	assign w3027 = 1'b0;
	wire w3028;
	assign w3028 = 1'b0;
	wire w3029;
	assign w3029 = 1'b0;
	wire w3030;
	assign w3030 = 1'b0;
	wire w3031;
	assign w3031 = 1'b0;
	wire w3032;
	assign w3032 = 1'b0;
	wire w3033;
	assign w3033 = 1'b0;
	wire w3199;
	assign w3199 = 1'b1;
	wire w3200;
	assign w3200 = 1'b1;
	wire w3201;
	assign w3201 = 1'b1;
	wire w3202;
	assign w3202 = 1'b1;
	wire w3203;
	assign w3203 = 1'b1;
	wire w3204;
	assign w3204 = 1'b1;
	wire w3205;
	assign w3205 = 1'b1;
	wire w3206;
	assign w3206 = 1'b1;
	wire w3233;
	assign w3233 = 1'b0;
	wire w3234;
	assign w3234 = 1'b0;
	wire w3235;
	assign w3235 = 1'b0;
	wire w3236;
	assign w3236 = 1'b0;
	wire w3237;
	assign w3237 = 1'b0;
	wire w3238;
	assign w3238 = 1'b0;
	wire w3239;
	assign w3239 = 1'b0;
	wire w3240;
	assign w3240 = 1'b0;
	wire w3406;
	assign w3406 = 1'b1;
	wire w3407;
	assign w3407 = 1'b1;
	wire w3408;
	assign w3408 = 1'b1;
	wire w3409;
	assign w3409 = 1'b1;
	wire w3410;
	assign w3410 = 1'b1;
	wire w3411;
	assign w3411 = 1'b1;
	wire w3412;
	assign w3412 = 1'b1;
	wire w3413;
	assign w3413 = 1'b1;
	
	XOR U0 ( .A(w131), .B(w0), .Z(w136) );
	XOR U1 ( .A(w132), .B(w0), .Z(w137) );
	XOR U2 ( .A(w135), .B(w0), .Z(w138) );
	XOR U3 ( .A(w128), .B(w1), .Z(w139) );
	XOR U4 ( .A(w129), .B(w1), .Z(w140) );
	XOR U5 ( .A(w137), .B(w1), .Z(w141) );
	XOR U6 ( .A(w133), .B(w1), .Z(w142) );
	XOR U7 ( .A(w134), .B(w1), .Z(w143) );
	XOR U8 ( .A(w138), .B(w1), .Z(w144) );
	XOR U9 ( .A(w140), .B(w2), .Z(w145) );
	XOR U10 ( .A(w141), .B(w2), .Z(w146) );
	XOR U11 ( .A(w142), .B(w2), .Z(w147) );
	XOR U12 ( .A(w143), .B(w2), .Z(w148) );
	XOR U13 ( .A(w144), .B(w2), .Z(w149) );
	XOR U14 ( .A(w136), .B(w3), .Z(w150) );
	XOR U15 ( .A(w148), .B(w3), .Z(w151) );
	XOR U16 ( .A(w139), .B(w4), .Z(w152) );
	XOR U17 ( .A(w150), .B(w4), .Z(w153) );
	XOR U18 ( .A(w152), .B(w5), .Z(w154) );
	XOR U19 ( .A(w149), .B(w5), .Z(w155) );
	XOR U20 ( .A(w154), .B(w6), .Z(w156) );
	XOR U21 ( .A(w153), .B(w6), .Z(w157) );
	XOR U22 ( .A(w147), .B(w6), .Z(w158) );
	XOR U23 ( .A(w155), .B(w6), .Z(w159) );
	XOR U24 ( .A(w156), .B(w7), .Z(w160) );
	XOR U25 ( .A(w145), .B(w7), .Z(w161) );
	XOR U26 ( .A(w130), .B(w7), .Z(w162) );
	XOR U27 ( .A(w157), .B(w7), .Z(w163) );
	XOR U28 ( .A(w146), .B(w7), .Z(w164) );
	XOR U29 ( .A(w158), .B(w7), .Z(w165) );
	XOR U30 ( .A(w151), .B(w7), .Z(w166) );
	XOR U31 ( .A(w159), .B(w7), .Z(w167) );
	XOR U32 ( .A(w160), .B(w164), .Z(w168) );
	XOR U33 ( .A(w161), .B(w165), .Z(w169) );
	XOR U34 ( .A(w162), .B(w166), .Z(w170) );
	XOR U35 ( .A(w163), .B(w167), .Z(w171) );
	XOR U36 ( .A(w170), .B(w168), .Z(w172) );
	XOR U37 ( .A(w171), .B(w169), .Z(w173) );
	XOR U38 ( .A(w169), .B(w168), .Z(w174) );
	XOR U39 ( .A(w162), .B(w160), .Z(w177) );
	XOR U40 ( .A(w163), .B(w161), .Z(w178) );
	XOR U41 ( .A(w166), .B(w164), .Z(w179) );
	XOR U42 ( .A(w167), .B(w165), .Z(w180) );
	XOR U43 ( .A(w178), .B(w177), .Z(w181) );
	XOR U44 ( .A(w180), .B(w179), .Z(w182) );
	AND U45 ( .A(w181), .B(w182), .Z(w183) );
	AND U46 ( .A(w178), .B(w180), .Z(w184) );
	XOR U47 ( .A(w184), .B(w183), .Z(w185) );
	AND U48 ( .A(w177), .B(w179), .Z(w186) );
	XOR U49 ( .A(w186), .B(w183), .Z(w187) );
	XOR U50 ( .A(w187), .B(w185), .Z(w188) );
	XOR U51 ( .A(w163), .B(w162), .Z(w189) );
	XOR U52 ( .A(w167), .B(w166), .Z(w190) );
	AND U53 ( .A(w189), .B(w190), .Z(w191) );
	AND U54 ( .A(w163), .B(w167), .Z(w192) );
	XOR U55 ( .A(w192), .B(w191), .Z(w193) );
	AND U56 ( .A(w162), .B(w166), .Z(w194) );
	XOR U57 ( .A(w194), .B(w191), .Z(w195) );
	XOR U58 ( .A(w161), .B(w160), .Z(w196) );
	XOR U59 ( .A(w165), .B(w164), .Z(w197) );
	AND U60 ( .A(w196), .B(w197), .Z(w198) );
	AND U61 ( .A(w161), .B(w165), .Z(w199) );
	XOR U62 ( .A(w199), .B(w198), .Z(w200) );
	AND U63 ( .A(w160), .B(w164), .Z(w201) );
	XOR U64 ( .A(w201), .B(w198), .Z(w202) );
	XOR U65 ( .A(w195), .B(w188), .Z(w203) );
	XOR U66 ( .A(w193), .B(w187), .Z(w204) );
	XOR U67 ( .A(w202), .B(w188), .Z(w205) );
	XOR U68 ( .A(w200), .B(w187), .Z(w206) );
	XOR U69 ( .A(w168), .B(w205), .Z(w207) );
	XOR U70 ( .A(w174), .B(w206), .Z(w208) );
	XOR U71 ( .A(w173), .B(w203), .Z(w209) );
	XOR U72 ( .A(w172), .B(w204), .Z(w210) );
	XOR U73 ( .A(w209), .B(w207), .Z(w211) );
	XOR U74 ( .A(w210), .B(w208), .Z(w212) );
	XOR U75 ( .A(w212), .B(w211), .Z(w213) );
	XOR U76 ( .A(w210), .B(w209), .Z(w214) );
	XOR U77 ( .A(w208), .B(w207), .Z(w215) );
	AND U78 ( .A(w214), .B(w215), .Z(w216) );
	AND U79 ( .A(w210), .B(w208), .Z(w217) );
	XOR U80 ( .A(w217), .B(w216), .Z(w218) );
	AND U81 ( .A(w209), .B(w207), .Z(w219) );
	XOR U82 ( .A(w219), .B(w216), .Z(w220) );
	XOR U83 ( .A(w213), .B(w220), .Z(w221) );
	XOR U84 ( .A(w212), .B(w218), .Z(w222) );
	XOR U85 ( .A(w221), .B(w222), .Z(w223) );
	XOR U86 ( .A(w208), .B(w207), .Z(w224) );
	AND U87 ( .A(w223), .B(w224), .Z(w225) );
	AND U88 ( .A(w221), .B(w208), .Z(w226) );
	XOR U89 ( .A(w226), .B(w225), .Z(w227) );
	AND U90 ( .A(w222), .B(w207), .Z(w228) );
	XOR U91 ( .A(w228), .B(w225), .Z(w229) );
	XOR U92 ( .A(w221), .B(w222), .Z(w230) );
	XOR U93 ( .A(w210), .B(w209), .Z(w231) );
	AND U94 ( .A(w230), .B(w231), .Z(w232) );
	AND U95 ( .A(w221), .B(w210), .Z(w233) );
	XOR U96 ( .A(w233), .B(w232), .Z(w234) );
	AND U97 ( .A(w222), .B(w209), .Z(w235) );
	XOR U98 ( .A(w235), .B(w232), .Z(w236) );
	XOR U99 ( .A(w229), .B(w236), .Z(w239) );
	XOR U100 ( .A(w227), .B(w234), .Z(w240) );
	XOR U101 ( .A(w166), .B(w164), .Z(w241) );
	XOR U102 ( .A(w167), .B(w165), .Z(w242) );
	XOR U103 ( .A(w240), .B(w239), .Z(w243) );
	XOR U104 ( .A(w242), .B(w241), .Z(w244) );
	AND U105 ( .A(w243), .B(w244), .Z(w245) );
	AND U106 ( .A(w240), .B(w242), .Z(w246) );
	XOR U107 ( .A(w246), .B(w245), .Z(w247) );
	AND U108 ( .A(w239), .B(w241), .Z(w248) );
	XOR U109 ( .A(w248), .B(w245), .Z(w249) );
	XOR U110 ( .A(w249), .B(w247), .Z(w250) );
	XOR U111 ( .A(w227), .B(w229), .Z(w251) );
	XOR U112 ( .A(w167), .B(w166), .Z(w252) );
	AND U113 ( .A(w251), .B(w252), .Z(w253) );
	AND U114 ( .A(w227), .B(w167), .Z(w254) );
	XOR U115 ( .A(w254), .B(w253), .Z(w255) );
	AND U116 ( .A(w229), .B(w166), .Z(w256) );
	XOR U117 ( .A(w256), .B(w253), .Z(w257) );
	XOR U118 ( .A(w234), .B(w236), .Z(w258) );
	XOR U119 ( .A(w165), .B(w164), .Z(w259) );
	AND U120 ( .A(w258), .B(w259), .Z(w260) );
	AND U121 ( .A(w234), .B(w165), .Z(w261) );
	XOR U122 ( .A(w261), .B(w260), .Z(w262) );
	AND U123 ( .A(w236), .B(w164), .Z(w263) );
	XOR U124 ( .A(w263), .B(w260), .Z(w264) );
	XOR U125 ( .A(w257), .B(w250), .Z(w265) );
	XOR U126 ( .A(w255), .B(w249), .Z(w266) );
	XOR U127 ( .A(w264), .B(w250), .Z(w267) );
	XOR U128 ( .A(w262), .B(w249), .Z(w268) );
	XOR U129 ( .A(w229), .B(w236), .Z(w271) );
	XOR U130 ( .A(w227), .B(w234), .Z(w272) );
	XOR U131 ( .A(w162), .B(w160), .Z(w273) );
	XOR U132 ( .A(w163), .B(w161), .Z(w274) );
	XOR U133 ( .A(w272), .B(w271), .Z(w275) );
	XOR U134 ( .A(w274), .B(w273), .Z(w276) );
	AND U135 ( .A(w275), .B(w276), .Z(w277) );
	AND U136 ( .A(w272), .B(w274), .Z(w278) );
	XOR U137 ( .A(w278), .B(w277), .Z(w279) );
	AND U138 ( .A(w271), .B(w273), .Z(w280) );
	XOR U139 ( .A(w280), .B(w277), .Z(w281) );
	XOR U140 ( .A(w281), .B(w279), .Z(w282) );
	XOR U141 ( .A(w227), .B(w229), .Z(w283) );
	XOR U142 ( .A(w163), .B(w162), .Z(w284) );
	AND U143 ( .A(w283), .B(w284), .Z(w285) );
	AND U144 ( .A(w227), .B(w163), .Z(w286) );
	XOR U145 ( .A(w286), .B(w285), .Z(w287) );
	AND U146 ( .A(w229), .B(w162), .Z(w288) );
	XOR U147 ( .A(w288), .B(w285), .Z(w289) );
	XOR U148 ( .A(w234), .B(w236), .Z(w290) );
	XOR U149 ( .A(w161), .B(w160), .Z(w291) );
	AND U150 ( .A(w290), .B(w291), .Z(w292) );
	AND U151 ( .A(w234), .B(w161), .Z(w293) );
	XOR U152 ( .A(w293), .B(w292), .Z(w294) );
	AND U153 ( .A(w236), .B(w160), .Z(w295) );
	XOR U154 ( .A(w295), .B(w292), .Z(w296) );
	XOR U155 ( .A(w289), .B(w282), .Z(w297) );
	XOR U156 ( .A(w287), .B(w281), .Z(w298) );
	XOR U157 ( .A(w296), .B(w282), .Z(w299) );
	XOR U158 ( .A(w294), .B(w281), .Z(w300) );
	XOR U159 ( .A(w303), .B(w299), .Z(w309) );
	XOR U160 ( .A(w304), .B(w299), .Z(w310) );
	XOR U161 ( .A(w308), .B(w299), .Z(w311) );
	XOR U162 ( .A(w301), .B(w300), .Z(w312) );
	XOR U163 ( .A(w310), .B(w300), .Z(w313) );
	XOR U164 ( .A(w305), .B(w300), .Z(w314) );
	XOR U165 ( .A(w306), .B(w300), .Z(w315) );
	XOR U166 ( .A(w307), .B(w300), .Z(w316) );
	XOR U167 ( .A(w312), .B(w297), .Z(w317) );
	XOR U168 ( .A(w309), .B(w297), .Z(w318) );
	XOR U169 ( .A(w317), .B(w298), .Z(w319) );
	XOR U170 ( .A(w302), .B(w298), .Z(w320) );
	XOR U171 ( .A(w313), .B(w298), .Z(w321) );
	XOR U172 ( .A(w315), .B(w298), .Z(w322) );
	XOR U173 ( .A(w316), .B(w298), .Z(w323) );
	XOR U174 ( .A(w311), .B(w298), .Z(w324) );
	XOR U175 ( .A(w320), .B(w267), .Z(w325) );
	XOR U176 ( .A(w314), .B(w267), .Z(w326) );
	XOR U177 ( .A(w318), .B(w268), .Z(w327) );
	XOR U178 ( .A(w319), .B(w265), .Z(w328) );
	XOR U179 ( .A(w326), .B(w265), .Z(w329) );
	XOR U180 ( .A(w323), .B(w265), .Z(w330) );
	XOR U181 ( .A(w328), .B(w266), .Z(w331) );
	XOR U182 ( .A(w325), .B(w266), .Z(w332) );
	XOR U183 ( .A(w329), .B(w266), .Z(w333) );
	XOR U184 ( .A(w330), .B(w266), .Z(w334) );
	XOR U185 ( .A(w338), .B(w8), .Z(w343) );
	XOR U186 ( .A(w339), .B(w8), .Z(w344) );
	XOR U187 ( .A(w342), .B(w8), .Z(w345) );
	XOR U188 ( .A(w335), .B(w9), .Z(w346) );
	XOR U189 ( .A(w336), .B(w9), .Z(w347) );
	XOR U190 ( .A(w344), .B(w9), .Z(w348) );
	XOR U191 ( .A(w340), .B(w9), .Z(w349) );
	XOR U192 ( .A(w341), .B(w9), .Z(w350) );
	XOR U193 ( .A(w345), .B(w9), .Z(w351) );
	XOR U194 ( .A(w347), .B(w10), .Z(w352) );
	XOR U195 ( .A(w348), .B(w10), .Z(w353) );
	XOR U196 ( .A(w349), .B(w10), .Z(w354) );
	XOR U197 ( .A(w350), .B(w10), .Z(w355) );
	XOR U198 ( .A(w351), .B(w10), .Z(w356) );
	XOR U199 ( .A(w343), .B(w11), .Z(w357) );
	XOR U200 ( .A(w355), .B(w11), .Z(w358) );
	XOR U201 ( .A(w346), .B(w12), .Z(w359) );
	XOR U202 ( .A(w357), .B(w12), .Z(w360) );
	XOR U203 ( .A(w359), .B(w13), .Z(w361) );
	XOR U204 ( .A(w356), .B(w13), .Z(w362) );
	XOR U205 ( .A(w361), .B(w14), .Z(w363) );
	XOR U206 ( .A(w360), .B(w14), .Z(w364) );
	XOR U207 ( .A(w354), .B(w14), .Z(w365) );
	XOR U208 ( .A(w362), .B(w14), .Z(w366) );
	XOR U209 ( .A(w363), .B(w15), .Z(w367) );
	XOR U210 ( .A(w352), .B(w15), .Z(w368) );
	XOR U211 ( .A(w337), .B(w15), .Z(w369) );
	XOR U212 ( .A(w364), .B(w15), .Z(w370) );
	XOR U213 ( .A(w353), .B(w15), .Z(w371) );
	XOR U214 ( .A(w365), .B(w15), .Z(w372) );
	XOR U215 ( .A(w358), .B(w15), .Z(w373) );
	XOR U216 ( .A(w366), .B(w15), .Z(w374) );
	XOR U217 ( .A(w367), .B(w371), .Z(w375) );
	XOR U218 ( .A(w368), .B(w372), .Z(w376) );
	XOR U219 ( .A(w369), .B(w373), .Z(w377) );
	XOR U220 ( .A(w370), .B(w374), .Z(w378) );
	XOR U221 ( .A(w377), .B(w375), .Z(w379) );
	XOR U222 ( .A(w378), .B(w376), .Z(w380) );
	XOR U223 ( .A(w376), .B(w375), .Z(w381) );
	XOR U224 ( .A(w369), .B(w367), .Z(w384) );
	XOR U225 ( .A(w370), .B(w368), .Z(w385) );
	XOR U226 ( .A(w373), .B(w371), .Z(w386) );
	XOR U227 ( .A(w374), .B(w372), .Z(w387) );
	XOR U228 ( .A(w385), .B(w384), .Z(w388) );
	XOR U229 ( .A(w387), .B(w386), .Z(w389) );
	AND U230 ( .A(w388), .B(w389), .Z(w390) );
	AND U231 ( .A(w385), .B(w387), .Z(w391) );
	XOR U232 ( .A(w391), .B(w390), .Z(w392) );
	AND U233 ( .A(w384), .B(w386), .Z(w393) );
	XOR U234 ( .A(w393), .B(w390), .Z(w394) );
	XOR U235 ( .A(w394), .B(w392), .Z(w395) );
	XOR U236 ( .A(w370), .B(w369), .Z(w396) );
	XOR U237 ( .A(w374), .B(w373), .Z(w397) );
	AND U238 ( .A(w396), .B(w397), .Z(w398) );
	AND U239 ( .A(w370), .B(w374), .Z(w399) );
	XOR U240 ( .A(w399), .B(w398), .Z(w400) );
	AND U241 ( .A(w369), .B(w373), .Z(w401) );
	XOR U242 ( .A(w401), .B(w398), .Z(w402) );
	XOR U243 ( .A(w368), .B(w367), .Z(w403) );
	XOR U244 ( .A(w372), .B(w371), .Z(w404) );
	AND U245 ( .A(w403), .B(w404), .Z(w405) );
	AND U246 ( .A(w368), .B(w372), .Z(w406) );
	XOR U247 ( .A(w406), .B(w405), .Z(w407) );
	AND U248 ( .A(w367), .B(w371), .Z(w408) );
	XOR U249 ( .A(w408), .B(w405), .Z(w409) );
	XOR U250 ( .A(w402), .B(w395), .Z(w410) );
	XOR U251 ( .A(w400), .B(w394), .Z(w411) );
	XOR U252 ( .A(w409), .B(w395), .Z(w412) );
	XOR U253 ( .A(w407), .B(w394), .Z(w413) );
	XOR U254 ( .A(w375), .B(w412), .Z(w414) );
	XOR U255 ( .A(w381), .B(w413), .Z(w415) );
	XOR U256 ( .A(w380), .B(w410), .Z(w416) );
	XOR U257 ( .A(w379), .B(w411), .Z(w417) );
	XOR U258 ( .A(w416), .B(w414), .Z(w418) );
	XOR U259 ( .A(w417), .B(w415), .Z(w419) );
	XOR U260 ( .A(w419), .B(w418), .Z(w420) );
	XOR U261 ( .A(w417), .B(w416), .Z(w421) );
	XOR U262 ( .A(w415), .B(w414), .Z(w422) );
	AND U263 ( .A(w421), .B(w422), .Z(w423) );
	AND U264 ( .A(w417), .B(w415), .Z(w424) );
	XOR U265 ( .A(w424), .B(w423), .Z(w425) );
	AND U266 ( .A(w416), .B(w414), .Z(w426) );
	XOR U267 ( .A(w426), .B(w423), .Z(w427) );
	XOR U268 ( .A(w420), .B(w427), .Z(w428) );
	XOR U269 ( .A(w419), .B(w425), .Z(w429) );
	XOR U270 ( .A(w428), .B(w429), .Z(w430) );
	XOR U271 ( .A(w415), .B(w414), .Z(w431) );
	AND U272 ( .A(w430), .B(w431), .Z(w432) );
	AND U273 ( .A(w428), .B(w415), .Z(w433) );
	XOR U274 ( .A(w433), .B(w432), .Z(w434) );
	AND U275 ( .A(w429), .B(w414), .Z(w435) );
	XOR U276 ( .A(w435), .B(w432), .Z(w436) );
	XOR U277 ( .A(w428), .B(w429), .Z(w437) );
	XOR U278 ( .A(w417), .B(w416), .Z(w438) );
	AND U279 ( .A(w437), .B(w438), .Z(w439) );
	AND U280 ( .A(w428), .B(w417), .Z(w440) );
	XOR U281 ( .A(w440), .B(w439), .Z(w441) );
	AND U282 ( .A(w429), .B(w416), .Z(w442) );
	XOR U283 ( .A(w442), .B(w439), .Z(w443) );
	XOR U284 ( .A(w436), .B(w443), .Z(w446) );
	XOR U285 ( .A(w434), .B(w441), .Z(w447) );
	XOR U286 ( .A(w373), .B(w371), .Z(w448) );
	XOR U287 ( .A(w374), .B(w372), .Z(w449) );
	XOR U288 ( .A(w447), .B(w446), .Z(w450) );
	XOR U289 ( .A(w449), .B(w448), .Z(w451) );
	AND U290 ( .A(w450), .B(w451), .Z(w452) );
	AND U291 ( .A(w447), .B(w449), .Z(w453) );
	XOR U292 ( .A(w453), .B(w452), .Z(w454) );
	AND U293 ( .A(w446), .B(w448), .Z(w455) );
	XOR U294 ( .A(w455), .B(w452), .Z(w456) );
	XOR U295 ( .A(w456), .B(w454), .Z(w457) );
	XOR U296 ( .A(w434), .B(w436), .Z(w458) );
	XOR U297 ( .A(w374), .B(w373), .Z(w459) );
	AND U298 ( .A(w458), .B(w459), .Z(w460) );
	AND U299 ( .A(w434), .B(w374), .Z(w461) );
	XOR U300 ( .A(w461), .B(w460), .Z(w462) );
	AND U301 ( .A(w436), .B(w373), .Z(w463) );
	XOR U302 ( .A(w463), .B(w460), .Z(w464) );
	XOR U303 ( .A(w441), .B(w443), .Z(w465) );
	XOR U304 ( .A(w372), .B(w371), .Z(w466) );
	AND U305 ( .A(w465), .B(w466), .Z(w467) );
	AND U306 ( .A(w441), .B(w372), .Z(w468) );
	XOR U307 ( .A(w468), .B(w467), .Z(w469) );
	AND U308 ( .A(w443), .B(w371), .Z(w470) );
	XOR U309 ( .A(w470), .B(w467), .Z(w471) );
	XOR U310 ( .A(w464), .B(w457), .Z(w472) );
	XOR U311 ( .A(w462), .B(w456), .Z(w473) );
	XOR U312 ( .A(w471), .B(w457), .Z(w474) );
	XOR U313 ( .A(w469), .B(w456), .Z(w475) );
	XOR U314 ( .A(w436), .B(w443), .Z(w478) );
	XOR U315 ( .A(w434), .B(w441), .Z(w479) );
	XOR U316 ( .A(w369), .B(w367), .Z(w480) );
	XOR U317 ( .A(w370), .B(w368), .Z(w481) );
	XOR U318 ( .A(w479), .B(w478), .Z(w482) );
	XOR U319 ( .A(w481), .B(w480), .Z(w483) );
	AND U320 ( .A(w482), .B(w483), .Z(w484) );
	AND U321 ( .A(w479), .B(w481), .Z(w485) );
	XOR U322 ( .A(w485), .B(w484), .Z(w486) );
	AND U323 ( .A(w478), .B(w480), .Z(w487) );
	XOR U324 ( .A(w487), .B(w484), .Z(w488) );
	XOR U325 ( .A(w488), .B(w486), .Z(w489) );
	XOR U326 ( .A(w434), .B(w436), .Z(w490) );
	XOR U327 ( .A(w370), .B(w369), .Z(w491) );
	AND U328 ( .A(w490), .B(w491), .Z(w492) );
	AND U329 ( .A(w434), .B(w370), .Z(w493) );
	XOR U330 ( .A(w493), .B(w492), .Z(w494) );
	AND U331 ( .A(w436), .B(w369), .Z(w495) );
	XOR U332 ( .A(w495), .B(w492), .Z(w496) );
	XOR U333 ( .A(w441), .B(w443), .Z(w497) );
	XOR U334 ( .A(w368), .B(w367), .Z(w498) );
	AND U335 ( .A(w497), .B(w498), .Z(w499) );
	AND U336 ( .A(w441), .B(w368), .Z(w500) );
	XOR U337 ( .A(w500), .B(w499), .Z(w501) );
	AND U338 ( .A(w443), .B(w367), .Z(w502) );
	XOR U339 ( .A(w502), .B(w499), .Z(w503) );
	XOR U340 ( .A(w496), .B(w489), .Z(w504) );
	XOR U341 ( .A(w494), .B(w488), .Z(w505) );
	XOR U342 ( .A(w503), .B(w489), .Z(w506) );
	XOR U343 ( .A(w501), .B(w488), .Z(w507) );
	XOR U344 ( .A(w510), .B(w506), .Z(w516) );
	XOR U345 ( .A(w511), .B(w506), .Z(w517) );
	XOR U346 ( .A(w515), .B(w506), .Z(w518) );
	XOR U347 ( .A(w508), .B(w507), .Z(w519) );
	XOR U348 ( .A(w517), .B(w507), .Z(w520) );
	XOR U349 ( .A(w512), .B(w507), .Z(w521) );
	XOR U350 ( .A(w513), .B(w507), .Z(w522) );
	XOR U351 ( .A(w514), .B(w507), .Z(w523) );
	XOR U352 ( .A(w519), .B(w504), .Z(w524) );
	XOR U353 ( .A(w516), .B(w504), .Z(w525) );
	XOR U354 ( .A(w524), .B(w505), .Z(w526) );
	XOR U355 ( .A(w509), .B(w505), .Z(w527) );
	XOR U356 ( .A(w520), .B(w505), .Z(w528) );
	XOR U357 ( .A(w522), .B(w505), .Z(w529) );
	XOR U358 ( .A(w523), .B(w505), .Z(w530) );
	XOR U359 ( .A(w518), .B(w505), .Z(w531) );
	XOR U360 ( .A(w527), .B(w474), .Z(w532) );
	XOR U361 ( .A(w521), .B(w474), .Z(w533) );
	XOR U362 ( .A(w525), .B(w475), .Z(w534) );
	XOR U363 ( .A(w526), .B(w472), .Z(w535) );
	XOR U364 ( .A(w533), .B(w472), .Z(w536) );
	XOR U365 ( .A(w530), .B(w472), .Z(w537) );
	XOR U366 ( .A(w535), .B(w473), .Z(w538) );
	XOR U367 ( .A(w532), .B(w473), .Z(w539) );
	XOR U368 ( .A(w536), .B(w473), .Z(w540) );
	XOR U369 ( .A(w537), .B(w473), .Z(w541) );
	XOR U370 ( .A(w545), .B(w16), .Z(w550) );
	XOR U371 ( .A(w546), .B(w16), .Z(w551) );
	XOR U372 ( .A(w549), .B(w16), .Z(w552) );
	XOR U373 ( .A(w542), .B(w17), .Z(w553) );
	XOR U374 ( .A(w543), .B(w17), .Z(w554) );
	XOR U375 ( .A(w551), .B(w17), .Z(w555) );
	XOR U376 ( .A(w547), .B(w17), .Z(w556) );
	XOR U377 ( .A(w548), .B(w17), .Z(w557) );
	XOR U378 ( .A(w552), .B(w17), .Z(w558) );
	XOR U379 ( .A(w554), .B(w18), .Z(w559) );
	XOR U380 ( .A(w555), .B(w18), .Z(w560) );
	XOR U381 ( .A(w556), .B(w18), .Z(w561) );
	XOR U382 ( .A(w557), .B(w18), .Z(w562) );
	XOR U383 ( .A(w558), .B(w18), .Z(w563) );
	XOR U384 ( .A(w550), .B(w19), .Z(w564) );
	XOR U385 ( .A(w562), .B(w19), .Z(w565) );
	XOR U386 ( .A(w553), .B(w20), .Z(w566) );
	XOR U387 ( .A(w564), .B(w20), .Z(w567) );
	XOR U388 ( .A(w566), .B(w21), .Z(w568) );
	XOR U389 ( .A(w563), .B(w21), .Z(w569) );
	XOR U390 ( .A(w568), .B(w22), .Z(w570) );
	XOR U391 ( .A(w567), .B(w22), .Z(w571) );
	XOR U392 ( .A(w561), .B(w22), .Z(w572) );
	XOR U393 ( .A(w569), .B(w22), .Z(w573) );
	XOR U394 ( .A(w570), .B(w23), .Z(w574) );
	XOR U395 ( .A(w559), .B(w23), .Z(w575) );
	XOR U396 ( .A(w544), .B(w23), .Z(w576) );
	XOR U397 ( .A(w571), .B(w23), .Z(w577) );
	XOR U398 ( .A(w560), .B(w23), .Z(w578) );
	XOR U399 ( .A(w572), .B(w23), .Z(w579) );
	XOR U400 ( .A(w565), .B(w23), .Z(w580) );
	XOR U401 ( .A(w573), .B(w23), .Z(w581) );
	XOR U402 ( .A(w574), .B(w578), .Z(w582) );
	XOR U403 ( .A(w575), .B(w579), .Z(w583) );
	XOR U404 ( .A(w576), .B(w580), .Z(w584) );
	XOR U405 ( .A(w577), .B(w581), .Z(w585) );
	XOR U406 ( .A(w584), .B(w582), .Z(w586) );
	XOR U407 ( .A(w585), .B(w583), .Z(w587) );
	XOR U408 ( .A(w583), .B(w582), .Z(w588) );
	XOR U409 ( .A(w576), .B(w574), .Z(w591) );
	XOR U410 ( .A(w577), .B(w575), .Z(w592) );
	XOR U411 ( .A(w580), .B(w578), .Z(w593) );
	XOR U412 ( .A(w581), .B(w579), .Z(w594) );
	XOR U413 ( .A(w592), .B(w591), .Z(w595) );
	XOR U414 ( .A(w594), .B(w593), .Z(w596) );
	AND U415 ( .A(w595), .B(w596), .Z(w597) );
	AND U416 ( .A(w592), .B(w594), .Z(w598) );
	XOR U417 ( .A(w598), .B(w597), .Z(w599) );
	AND U418 ( .A(w591), .B(w593), .Z(w600) );
	XOR U419 ( .A(w600), .B(w597), .Z(w601) );
	XOR U420 ( .A(w601), .B(w599), .Z(w602) );
	XOR U421 ( .A(w577), .B(w576), .Z(w603) );
	XOR U422 ( .A(w581), .B(w580), .Z(w604) );
	AND U423 ( .A(w603), .B(w604), .Z(w605) );
	AND U424 ( .A(w577), .B(w581), .Z(w606) );
	XOR U425 ( .A(w606), .B(w605), .Z(w607) );
	AND U426 ( .A(w576), .B(w580), .Z(w608) );
	XOR U427 ( .A(w608), .B(w605), .Z(w609) );
	XOR U428 ( .A(w575), .B(w574), .Z(w610) );
	XOR U429 ( .A(w579), .B(w578), .Z(w611) );
	AND U430 ( .A(w610), .B(w611), .Z(w612) );
	AND U431 ( .A(w575), .B(w579), .Z(w613) );
	XOR U432 ( .A(w613), .B(w612), .Z(w614) );
	AND U433 ( .A(w574), .B(w578), .Z(w615) );
	XOR U434 ( .A(w615), .B(w612), .Z(w616) );
	XOR U435 ( .A(w609), .B(w602), .Z(w617) );
	XOR U436 ( .A(w607), .B(w601), .Z(w618) );
	XOR U437 ( .A(w616), .B(w602), .Z(w619) );
	XOR U438 ( .A(w614), .B(w601), .Z(w620) );
	XOR U439 ( .A(w582), .B(w619), .Z(w621) );
	XOR U440 ( .A(w588), .B(w620), .Z(w622) );
	XOR U441 ( .A(w587), .B(w617), .Z(w623) );
	XOR U442 ( .A(w586), .B(w618), .Z(w624) );
	XOR U443 ( .A(w623), .B(w621), .Z(w625) );
	XOR U444 ( .A(w624), .B(w622), .Z(w626) );
	XOR U445 ( .A(w626), .B(w625), .Z(w627) );
	XOR U446 ( .A(w624), .B(w623), .Z(w628) );
	XOR U447 ( .A(w622), .B(w621), .Z(w629) );
	AND U448 ( .A(w628), .B(w629), .Z(w630) );
	AND U449 ( .A(w624), .B(w622), .Z(w631) );
	XOR U450 ( .A(w631), .B(w630), .Z(w632) );
	AND U451 ( .A(w623), .B(w621), .Z(w633) );
	XOR U452 ( .A(w633), .B(w630), .Z(w634) );
	XOR U453 ( .A(w627), .B(w634), .Z(w635) );
	XOR U454 ( .A(w626), .B(w632), .Z(w636) );
	XOR U455 ( .A(w635), .B(w636), .Z(w637) );
	XOR U456 ( .A(w622), .B(w621), .Z(w638) );
	AND U457 ( .A(w637), .B(w638), .Z(w639) );
	AND U458 ( .A(w635), .B(w622), .Z(w640) );
	XOR U459 ( .A(w640), .B(w639), .Z(w641) );
	AND U460 ( .A(w636), .B(w621), .Z(w642) );
	XOR U461 ( .A(w642), .B(w639), .Z(w643) );
	XOR U462 ( .A(w635), .B(w636), .Z(w644) );
	XOR U463 ( .A(w624), .B(w623), .Z(w645) );
	AND U464 ( .A(w644), .B(w645), .Z(w646) );
	AND U465 ( .A(w635), .B(w624), .Z(w647) );
	XOR U466 ( .A(w647), .B(w646), .Z(w648) );
	AND U467 ( .A(w636), .B(w623), .Z(w649) );
	XOR U468 ( .A(w649), .B(w646), .Z(w650) );
	XOR U469 ( .A(w643), .B(w650), .Z(w653) );
	XOR U470 ( .A(w641), .B(w648), .Z(w654) );
	XOR U471 ( .A(w580), .B(w578), .Z(w655) );
	XOR U472 ( .A(w581), .B(w579), .Z(w656) );
	XOR U473 ( .A(w654), .B(w653), .Z(w657) );
	XOR U474 ( .A(w656), .B(w655), .Z(w658) );
	AND U475 ( .A(w657), .B(w658), .Z(w659) );
	AND U476 ( .A(w654), .B(w656), .Z(w660) );
	XOR U477 ( .A(w660), .B(w659), .Z(w661) );
	AND U478 ( .A(w653), .B(w655), .Z(w662) );
	XOR U479 ( .A(w662), .B(w659), .Z(w663) );
	XOR U480 ( .A(w663), .B(w661), .Z(w664) );
	XOR U481 ( .A(w641), .B(w643), .Z(w665) );
	XOR U482 ( .A(w581), .B(w580), .Z(w666) );
	AND U483 ( .A(w665), .B(w666), .Z(w667) );
	AND U484 ( .A(w641), .B(w581), .Z(w668) );
	XOR U485 ( .A(w668), .B(w667), .Z(w669) );
	AND U486 ( .A(w643), .B(w580), .Z(w670) );
	XOR U487 ( .A(w670), .B(w667), .Z(w671) );
	XOR U488 ( .A(w648), .B(w650), .Z(w672) );
	XOR U489 ( .A(w579), .B(w578), .Z(w673) );
	AND U490 ( .A(w672), .B(w673), .Z(w674) );
	AND U491 ( .A(w648), .B(w579), .Z(w675) );
	XOR U492 ( .A(w675), .B(w674), .Z(w676) );
	AND U493 ( .A(w650), .B(w578), .Z(w677) );
	XOR U494 ( .A(w677), .B(w674), .Z(w678) );
	XOR U495 ( .A(w671), .B(w664), .Z(w679) );
	XOR U496 ( .A(w669), .B(w663), .Z(w680) );
	XOR U497 ( .A(w678), .B(w664), .Z(w681) );
	XOR U498 ( .A(w676), .B(w663), .Z(w682) );
	XOR U499 ( .A(w643), .B(w650), .Z(w685) );
	XOR U500 ( .A(w641), .B(w648), .Z(w686) );
	XOR U501 ( .A(w576), .B(w574), .Z(w687) );
	XOR U502 ( .A(w577), .B(w575), .Z(w688) );
	XOR U503 ( .A(w686), .B(w685), .Z(w689) );
	XOR U504 ( .A(w688), .B(w687), .Z(w690) );
	AND U505 ( .A(w689), .B(w690), .Z(w691) );
	AND U506 ( .A(w686), .B(w688), .Z(w692) );
	XOR U507 ( .A(w692), .B(w691), .Z(w693) );
	AND U508 ( .A(w685), .B(w687), .Z(w694) );
	XOR U509 ( .A(w694), .B(w691), .Z(w695) );
	XOR U510 ( .A(w695), .B(w693), .Z(w696) );
	XOR U511 ( .A(w641), .B(w643), .Z(w697) );
	XOR U512 ( .A(w577), .B(w576), .Z(w698) );
	AND U513 ( .A(w697), .B(w698), .Z(w699) );
	AND U514 ( .A(w641), .B(w577), .Z(w700) );
	XOR U515 ( .A(w700), .B(w699), .Z(w701) );
	AND U516 ( .A(w643), .B(w576), .Z(w702) );
	XOR U517 ( .A(w702), .B(w699), .Z(w703) );
	XOR U518 ( .A(w648), .B(w650), .Z(w704) );
	XOR U519 ( .A(w575), .B(w574), .Z(w705) );
	AND U520 ( .A(w704), .B(w705), .Z(w706) );
	AND U521 ( .A(w648), .B(w575), .Z(w707) );
	XOR U522 ( .A(w707), .B(w706), .Z(w708) );
	AND U523 ( .A(w650), .B(w574), .Z(w709) );
	XOR U524 ( .A(w709), .B(w706), .Z(w710) );
	XOR U525 ( .A(w703), .B(w696), .Z(w711) );
	XOR U526 ( .A(w701), .B(w695), .Z(w712) );
	XOR U527 ( .A(w710), .B(w696), .Z(w713) );
	XOR U528 ( .A(w708), .B(w695), .Z(w714) );
	XOR U529 ( .A(w717), .B(w713), .Z(w723) );
	XOR U530 ( .A(w718), .B(w713), .Z(w724) );
	XOR U531 ( .A(w722), .B(w713), .Z(w725) );
	XOR U532 ( .A(w715), .B(w714), .Z(w726) );
	XOR U533 ( .A(w724), .B(w714), .Z(w727) );
	XOR U534 ( .A(w719), .B(w714), .Z(w728) );
	XOR U535 ( .A(w720), .B(w714), .Z(w729) );
	XOR U536 ( .A(w721), .B(w714), .Z(w730) );
	XOR U537 ( .A(w726), .B(w711), .Z(w731) );
	XOR U538 ( .A(w723), .B(w711), .Z(w732) );
	XOR U539 ( .A(w731), .B(w712), .Z(w733) );
	XOR U540 ( .A(w716), .B(w712), .Z(w734) );
	XOR U541 ( .A(w727), .B(w712), .Z(w735) );
	XOR U542 ( .A(w729), .B(w712), .Z(w736) );
	XOR U543 ( .A(w730), .B(w712), .Z(w737) );
	XOR U544 ( .A(w725), .B(w712), .Z(w738) );
	XOR U545 ( .A(w734), .B(w681), .Z(w739) );
	XOR U546 ( .A(w728), .B(w681), .Z(w740) );
	XOR U547 ( .A(w732), .B(w682), .Z(w741) );
	XOR U548 ( .A(w733), .B(w679), .Z(w742) );
	XOR U549 ( .A(w740), .B(w679), .Z(w743) );
	XOR U550 ( .A(w737), .B(w679), .Z(w744) );
	XOR U551 ( .A(w742), .B(w680), .Z(w745) );
	XOR U552 ( .A(w739), .B(w680), .Z(w746) );
	XOR U553 ( .A(w743), .B(w680), .Z(w747) );
	XOR U554 ( .A(w744), .B(w680), .Z(w748) );
	XOR U555 ( .A(w752), .B(w24), .Z(w757) );
	XOR U556 ( .A(w753), .B(w24), .Z(w758) );
	XOR U557 ( .A(w756), .B(w24), .Z(w759) );
	XOR U558 ( .A(w749), .B(w25), .Z(w760) );
	XOR U559 ( .A(w750), .B(w25), .Z(w761) );
	XOR U560 ( .A(w758), .B(w25), .Z(w762) );
	XOR U561 ( .A(w754), .B(w25), .Z(w763) );
	XOR U562 ( .A(w755), .B(w25), .Z(w764) );
	XOR U563 ( .A(w759), .B(w25), .Z(w765) );
	XOR U564 ( .A(w761), .B(w26), .Z(w766) );
	XOR U565 ( .A(w762), .B(w26), .Z(w767) );
	XOR U566 ( .A(w763), .B(w26), .Z(w768) );
	XOR U567 ( .A(w764), .B(w26), .Z(w769) );
	XOR U568 ( .A(w765), .B(w26), .Z(w770) );
	XOR U569 ( .A(w757), .B(w27), .Z(w771) );
	XOR U570 ( .A(w769), .B(w27), .Z(w772) );
	XOR U571 ( .A(w760), .B(w28), .Z(w773) );
	XOR U572 ( .A(w771), .B(w28), .Z(w774) );
	XOR U573 ( .A(w773), .B(w29), .Z(w775) );
	XOR U574 ( .A(w770), .B(w29), .Z(w776) );
	XOR U575 ( .A(w775), .B(w30), .Z(w777) );
	XOR U576 ( .A(w774), .B(w30), .Z(w778) );
	XOR U577 ( .A(w768), .B(w30), .Z(w779) );
	XOR U578 ( .A(w776), .B(w30), .Z(w780) );
	XOR U579 ( .A(w777), .B(w31), .Z(w781) );
	XOR U580 ( .A(w766), .B(w31), .Z(w782) );
	XOR U581 ( .A(w751), .B(w31), .Z(w783) );
	XOR U582 ( .A(w778), .B(w31), .Z(w784) );
	XOR U583 ( .A(w767), .B(w31), .Z(w785) );
	XOR U584 ( .A(w779), .B(w31), .Z(w786) );
	XOR U585 ( .A(w772), .B(w31), .Z(w787) );
	XOR U586 ( .A(w780), .B(w31), .Z(w788) );
	XOR U587 ( .A(w781), .B(w785), .Z(w789) );
	XOR U588 ( .A(w782), .B(w786), .Z(w790) );
	XOR U589 ( .A(w783), .B(w787), .Z(w791) );
	XOR U590 ( .A(w784), .B(w788), .Z(w792) );
	XOR U591 ( .A(w791), .B(w789), .Z(w793) );
	XOR U592 ( .A(w792), .B(w790), .Z(w794) );
	XOR U593 ( .A(w790), .B(w789), .Z(w795) );
	XOR U594 ( .A(w783), .B(w781), .Z(w798) );
	XOR U595 ( .A(w784), .B(w782), .Z(w799) );
	XOR U596 ( .A(w787), .B(w785), .Z(w800) );
	XOR U597 ( .A(w788), .B(w786), .Z(w801) );
	XOR U598 ( .A(w799), .B(w798), .Z(w802) );
	XOR U599 ( .A(w801), .B(w800), .Z(w803) );
	AND U600 ( .A(w802), .B(w803), .Z(w804) );
	AND U601 ( .A(w799), .B(w801), .Z(w805) );
	XOR U602 ( .A(w805), .B(w804), .Z(w806) );
	AND U603 ( .A(w798), .B(w800), .Z(w807) );
	XOR U604 ( .A(w807), .B(w804), .Z(w808) );
	XOR U605 ( .A(w808), .B(w806), .Z(w809) );
	XOR U606 ( .A(w784), .B(w783), .Z(w810) );
	XOR U607 ( .A(w788), .B(w787), .Z(w811) );
	AND U608 ( .A(w810), .B(w811), .Z(w812) );
	AND U609 ( .A(w784), .B(w788), .Z(w813) );
	XOR U610 ( .A(w813), .B(w812), .Z(w814) );
	AND U611 ( .A(w783), .B(w787), .Z(w815) );
	XOR U612 ( .A(w815), .B(w812), .Z(w816) );
	XOR U613 ( .A(w782), .B(w781), .Z(w817) );
	XOR U614 ( .A(w786), .B(w785), .Z(w818) );
	AND U615 ( .A(w817), .B(w818), .Z(w819) );
	AND U616 ( .A(w782), .B(w786), .Z(w820) );
	XOR U617 ( .A(w820), .B(w819), .Z(w821) );
	AND U618 ( .A(w781), .B(w785), .Z(w822) );
	XOR U619 ( .A(w822), .B(w819), .Z(w823) );
	XOR U620 ( .A(w816), .B(w809), .Z(w824) );
	XOR U621 ( .A(w814), .B(w808), .Z(w825) );
	XOR U622 ( .A(w823), .B(w809), .Z(w826) );
	XOR U623 ( .A(w821), .B(w808), .Z(w827) );
	XOR U624 ( .A(w789), .B(w826), .Z(w828) );
	XOR U625 ( .A(w795), .B(w827), .Z(w829) );
	XOR U626 ( .A(w794), .B(w824), .Z(w830) );
	XOR U627 ( .A(w793), .B(w825), .Z(w831) );
	XOR U628 ( .A(w830), .B(w828), .Z(w832) );
	XOR U629 ( .A(w831), .B(w829), .Z(w833) );
	XOR U630 ( .A(w833), .B(w832), .Z(w834) );
	XOR U631 ( .A(w831), .B(w830), .Z(w835) );
	XOR U632 ( .A(w829), .B(w828), .Z(w836) );
	AND U633 ( .A(w835), .B(w836), .Z(w837) );
	AND U634 ( .A(w831), .B(w829), .Z(w838) );
	XOR U635 ( .A(w838), .B(w837), .Z(w839) );
	AND U636 ( .A(w830), .B(w828), .Z(w840) );
	XOR U637 ( .A(w840), .B(w837), .Z(w841) );
	XOR U638 ( .A(w834), .B(w841), .Z(w842) );
	XOR U639 ( .A(w833), .B(w839), .Z(w843) );
	XOR U640 ( .A(w842), .B(w843), .Z(w844) );
	XOR U641 ( .A(w829), .B(w828), .Z(w845) );
	AND U642 ( .A(w844), .B(w845), .Z(w846) );
	AND U643 ( .A(w842), .B(w829), .Z(w847) );
	XOR U644 ( .A(w847), .B(w846), .Z(w848) );
	AND U645 ( .A(w843), .B(w828), .Z(w849) );
	XOR U646 ( .A(w849), .B(w846), .Z(w850) );
	XOR U647 ( .A(w842), .B(w843), .Z(w851) );
	XOR U648 ( .A(w831), .B(w830), .Z(w852) );
	AND U649 ( .A(w851), .B(w852), .Z(w853) );
	AND U650 ( .A(w842), .B(w831), .Z(w854) );
	XOR U651 ( .A(w854), .B(w853), .Z(w855) );
	AND U652 ( .A(w843), .B(w830), .Z(w856) );
	XOR U653 ( .A(w856), .B(w853), .Z(w857) );
	XOR U654 ( .A(w850), .B(w857), .Z(w860) );
	XOR U655 ( .A(w848), .B(w855), .Z(w861) );
	XOR U656 ( .A(w787), .B(w785), .Z(w862) );
	XOR U657 ( .A(w788), .B(w786), .Z(w863) );
	XOR U658 ( .A(w861), .B(w860), .Z(w864) );
	XOR U659 ( .A(w863), .B(w862), .Z(w865) );
	AND U660 ( .A(w864), .B(w865), .Z(w866) );
	AND U661 ( .A(w861), .B(w863), .Z(w867) );
	XOR U662 ( .A(w867), .B(w866), .Z(w868) );
	AND U663 ( .A(w860), .B(w862), .Z(w869) );
	XOR U664 ( .A(w869), .B(w866), .Z(w870) );
	XOR U665 ( .A(w870), .B(w868), .Z(w871) );
	XOR U666 ( .A(w848), .B(w850), .Z(w872) );
	XOR U667 ( .A(w788), .B(w787), .Z(w873) );
	AND U668 ( .A(w872), .B(w873), .Z(w874) );
	AND U669 ( .A(w848), .B(w788), .Z(w875) );
	XOR U670 ( .A(w875), .B(w874), .Z(w876) );
	AND U671 ( .A(w850), .B(w787), .Z(w877) );
	XOR U672 ( .A(w877), .B(w874), .Z(w878) );
	XOR U673 ( .A(w855), .B(w857), .Z(w879) );
	XOR U674 ( .A(w786), .B(w785), .Z(w880) );
	AND U675 ( .A(w879), .B(w880), .Z(w881) );
	AND U676 ( .A(w855), .B(w786), .Z(w882) );
	XOR U677 ( .A(w882), .B(w881), .Z(w883) );
	AND U678 ( .A(w857), .B(w785), .Z(w884) );
	XOR U679 ( .A(w884), .B(w881), .Z(w885) );
	XOR U680 ( .A(w878), .B(w871), .Z(w886) );
	XOR U681 ( .A(w876), .B(w870), .Z(w887) );
	XOR U682 ( .A(w885), .B(w871), .Z(w888) );
	XOR U683 ( .A(w883), .B(w870), .Z(w889) );
	XOR U684 ( .A(w850), .B(w857), .Z(w892) );
	XOR U685 ( .A(w848), .B(w855), .Z(w893) );
	XOR U686 ( .A(w783), .B(w781), .Z(w894) );
	XOR U687 ( .A(w784), .B(w782), .Z(w895) );
	XOR U688 ( .A(w893), .B(w892), .Z(w896) );
	XOR U689 ( .A(w895), .B(w894), .Z(w897) );
	AND U690 ( .A(w896), .B(w897), .Z(w898) );
	AND U691 ( .A(w893), .B(w895), .Z(w899) );
	XOR U692 ( .A(w899), .B(w898), .Z(w900) );
	AND U693 ( .A(w892), .B(w894), .Z(w901) );
	XOR U694 ( .A(w901), .B(w898), .Z(w902) );
	XOR U695 ( .A(w902), .B(w900), .Z(w903) );
	XOR U696 ( .A(w848), .B(w850), .Z(w904) );
	XOR U697 ( .A(w784), .B(w783), .Z(w905) );
	AND U698 ( .A(w904), .B(w905), .Z(w906) );
	AND U699 ( .A(w848), .B(w784), .Z(w907) );
	XOR U700 ( .A(w907), .B(w906), .Z(w908) );
	AND U701 ( .A(w850), .B(w783), .Z(w909) );
	XOR U702 ( .A(w909), .B(w906), .Z(w910) );
	XOR U703 ( .A(w855), .B(w857), .Z(w911) );
	XOR U704 ( .A(w782), .B(w781), .Z(w912) );
	AND U705 ( .A(w911), .B(w912), .Z(w913) );
	AND U706 ( .A(w855), .B(w782), .Z(w914) );
	XOR U707 ( .A(w914), .B(w913), .Z(w915) );
	AND U708 ( .A(w857), .B(w781), .Z(w916) );
	XOR U709 ( .A(w916), .B(w913), .Z(w917) );
	XOR U710 ( .A(w910), .B(w903), .Z(w918) );
	XOR U711 ( .A(w908), .B(w902), .Z(w919) );
	XOR U712 ( .A(w917), .B(w903), .Z(w920) );
	XOR U713 ( .A(w915), .B(w902), .Z(w921) );
	XOR U714 ( .A(w924), .B(w920), .Z(w930) );
	XOR U715 ( .A(w925), .B(w920), .Z(w931) );
	XOR U716 ( .A(w929), .B(w920), .Z(w932) );
	XOR U717 ( .A(w922), .B(w921), .Z(w933) );
	XOR U718 ( .A(w931), .B(w921), .Z(w934) );
	XOR U719 ( .A(w926), .B(w921), .Z(w935) );
	XOR U720 ( .A(w927), .B(w921), .Z(w936) );
	XOR U721 ( .A(w928), .B(w921), .Z(w937) );
	XOR U722 ( .A(w933), .B(w918), .Z(w938) );
	XOR U723 ( .A(w930), .B(w918), .Z(w939) );
	XOR U724 ( .A(w938), .B(w919), .Z(w940) );
	XOR U725 ( .A(w923), .B(w919), .Z(w941) );
	XOR U726 ( .A(w934), .B(w919), .Z(w942) );
	XOR U727 ( .A(w936), .B(w919), .Z(w943) );
	XOR U728 ( .A(w937), .B(w919), .Z(w944) );
	XOR U729 ( .A(w932), .B(w919), .Z(w945) );
	XOR U730 ( .A(w941), .B(w888), .Z(w946) );
	XOR U731 ( .A(w935), .B(w888), .Z(w947) );
	XOR U732 ( .A(w939), .B(w889), .Z(w948) );
	XOR U733 ( .A(w940), .B(w886), .Z(w949) );
	XOR U734 ( .A(w947), .B(w886), .Z(w950) );
	XOR U735 ( .A(w944), .B(w886), .Z(w951) );
	XOR U736 ( .A(w949), .B(w887), .Z(w952) );
	XOR U737 ( .A(w946), .B(w887), .Z(w953) );
	XOR U738 ( .A(w950), .B(w887), .Z(w954) );
	XOR U739 ( .A(w951), .B(w887), .Z(w955) );
	XOR U740 ( .A(w959), .B(w32), .Z(w964) );
	XOR U741 ( .A(w960), .B(w32), .Z(w965) );
	XOR U742 ( .A(w963), .B(w32), .Z(w966) );
	XOR U743 ( .A(w956), .B(w33), .Z(w967) );
	XOR U744 ( .A(w957), .B(w33), .Z(w968) );
	XOR U745 ( .A(w965), .B(w33), .Z(w969) );
	XOR U746 ( .A(w961), .B(w33), .Z(w970) );
	XOR U747 ( .A(w962), .B(w33), .Z(w971) );
	XOR U748 ( .A(w966), .B(w33), .Z(w972) );
	XOR U749 ( .A(w968), .B(w34), .Z(w973) );
	XOR U750 ( .A(w969), .B(w34), .Z(w974) );
	XOR U751 ( .A(w970), .B(w34), .Z(w975) );
	XOR U752 ( .A(w971), .B(w34), .Z(w976) );
	XOR U753 ( .A(w972), .B(w34), .Z(w977) );
	XOR U754 ( .A(w964), .B(w35), .Z(w978) );
	XOR U755 ( .A(w976), .B(w35), .Z(w979) );
	XOR U756 ( .A(w967), .B(w36), .Z(w980) );
	XOR U757 ( .A(w978), .B(w36), .Z(w981) );
	XOR U758 ( .A(w980), .B(w37), .Z(w982) );
	XOR U759 ( .A(w977), .B(w37), .Z(w983) );
	XOR U760 ( .A(w982), .B(w38), .Z(w984) );
	XOR U761 ( .A(w981), .B(w38), .Z(w985) );
	XOR U762 ( .A(w975), .B(w38), .Z(w986) );
	XOR U763 ( .A(w983), .B(w38), .Z(w987) );
	XOR U764 ( .A(w984), .B(w39), .Z(w988) );
	XOR U765 ( .A(w973), .B(w39), .Z(w989) );
	XOR U766 ( .A(w958), .B(w39), .Z(w990) );
	XOR U767 ( .A(w985), .B(w39), .Z(w991) );
	XOR U768 ( .A(w974), .B(w39), .Z(w992) );
	XOR U769 ( .A(w986), .B(w39), .Z(w993) );
	XOR U770 ( .A(w979), .B(w39), .Z(w994) );
	XOR U771 ( .A(w987), .B(w39), .Z(w995) );
	XOR U772 ( .A(w988), .B(w992), .Z(w996) );
	XOR U773 ( .A(w989), .B(w993), .Z(w997) );
	XOR U774 ( .A(w990), .B(w994), .Z(w998) );
	XOR U775 ( .A(w991), .B(w995), .Z(w999) );
	XOR U776 ( .A(w998), .B(w996), .Z(w1000) );
	XOR U777 ( .A(w999), .B(w997), .Z(w1001) );
	XOR U778 ( .A(w997), .B(w996), .Z(w1002) );
	XOR U779 ( .A(w990), .B(w988), .Z(w1005) );
	XOR U780 ( .A(w991), .B(w989), .Z(w1006) );
	XOR U781 ( .A(w994), .B(w992), .Z(w1007) );
	XOR U782 ( .A(w995), .B(w993), .Z(w1008) );
	XOR U783 ( .A(w1006), .B(w1005), .Z(w1009) );
	XOR U784 ( .A(w1008), .B(w1007), .Z(w1010) );
	AND U785 ( .A(w1009), .B(w1010), .Z(w1011) );
	AND U786 ( .A(w1006), .B(w1008), .Z(w1012) );
	XOR U787 ( .A(w1012), .B(w1011), .Z(w1013) );
	AND U788 ( .A(w1005), .B(w1007), .Z(w1014) );
	XOR U789 ( .A(w1014), .B(w1011), .Z(w1015) );
	XOR U790 ( .A(w1015), .B(w1013), .Z(w1016) );
	XOR U791 ( .A(w991), .B(w990), .Z(w1017) );
	XOR U792 ( .A(w995), .B(w994), .Z(w1018) );
	AND U793 ( .A(w1017), .B(w1018), .Z(w1019) );
	AND U794 ( .A(w991), .B(w995), .Z(w1020) );
	XOR U795 ( .A(w1020), .B(w1019), .Z(w1021) );
	AND U796 ( .A(w990), .B(w994), .Z(w1022) );
	XOR U797 ( .A(w1022), .B(w1019), .Z(w1023) );
	XOR U798 ( .A(w989), .B(w988), .Z(w1024) );
	XOR U799 ( .A(w993), .B(w992), .Z(w1025) );
	AND U800 ( .A(w1024), .B(w1025), .Z(w1026) );
	AND U801 ( .A(w989), .B(w993), .Z(w1027) );
	XOR U802 ( .A(w1027), .B(w1026), .Z(w1028) );
	AND U803 ( .A(w988), .B(w992), .Z(w1029) );
	XOR U804 ( .A(w1029), .B(w1026), .Z(w1030) );
	XOR U805 ( .A(w1023), .B(w1016), .Z(w1031) );
	XOR U806 ( .A(w1021), .B(w1015), .Z(w1032) );
	XOR U807 ( .A(w1030), .B(w1016), .Z(w1033) );
	XOR U808 ( .A(w1028), .B(w1015), .Z(w1034) );
	XOR U809 ( .A(w996), .B(w1033), .Z(w1035) );
	XOR U810 ( .A(w1002), .B(w1034), .Z(w1036) );
	XOR U811 ( .A(w1001), .B(w1031), .Z(w1037) );
	XOR U812 ( .A(w1000), .B(w1032), .Z(w1038) );
	XOR U813 ( .A(w1037), .B(w1035), .Z(w1039) );
	XOR U814 ( .A(w1038), .B(w1036), .Z(w1040) );
	XOR U815 ( .A(w1040), .B(w1039), .Z(w1041) );
	XOR U816 ( .A(w1038), .B(w1037), .Z(w1042) );
	XOR U817 ( .A(w1036), .B(w1035), .Z(w1043) );
	AND U818 ( .A(w1042), .B(w1043), .Z(w1044) );
	AND U819 ( .A(w1038), .B(w1036), .Z(w1045) );
	XOR U820 ( .A(w1045), .B(w1044), .Z(w1046) );
	AND U821 ( .A(w1037), .B(w1035), .Z(w1047) );
	XOR U822 ( .A(w1047), .B(w1044), .Z(w1048) );
	XOR U823 ( .A(w1041), .B(w1048), .Z(w1049) );
	XOR U824 ( .A(w1040), .B(w1046), .Z(w1050) );
	XOR U825 ( .A(w1049), .B(w1050), .Z(w1051) );
	XOR U826 ( .A(w1036), .B(w1035), .Z(w1052) );
	AND U827 ( .A(w1051), .B(w1052), .Z(w1053) );
	AND U828 ( .A(w1049), .B(w1036), .Z(w1054) );
	XOR U829 ( .A(w1054), .B(w1053), .Z(w1055) );
	AND U830 ( .A(w1050), .B(w1035), .Z(w1056) );
	XOR U831 ( .A(w1056), .B(w1053), .Z(w1057) );
	XOR U832 ( .A(w1049), .B(w1050), .Z(w1058) );
	XOR U833 ( .A(w1038), .B(w1037), .Z(w1059) );
	AND U834 ( .A(w1058), .B(w1059), .Z(w1060) );
	AND U835 ( .A(w1049), .B(w1038), .Z(w1061) );
	XOR U836 ( .A(w1061), .B(w1060), .Z(w1062) );
	AND U837 ( .A(w1050), .B(w1037), .Z(w1063) );
	XOR U838 ( .A(w1063), .B(w1060), .Z(w1064) );
	XOR U839 ( .A(w1057), .B(w1064), .Z(w1067) );
	XOR U840 ( .A(w1055), .B(w1062), .Z(w1068) );
	XOR U841 ( .A(w994), .B(w992), .Z(w1069) );
	XOR U842 ( .A(w995), .B(w993), .Z(w1070) );
	XOR U843 ( .A(w1068), .B(w1067), .Z(w1071) );
	XOR U844 ( .A(w1070), .B(w1069), .Z(w1072) );
	AND U845 ( .A(w1071), .B(w1072), .Z(w1073) );
	AND U846 ( .A(w1068), .B(w1070), .Z(w1074) );
	XOR U847 ( .A(w1074), .B(w1073), .Z(w1075) );
	AND U848 ( .A(w1067), .B(w1069), .Z(w1076) );
	XOR U849 ( .A(w1076), .B(w1073), .Z(w1077) );
	XOR U850 ( .A(w1077), .B(w1075), .Z(w1078) );
	XOR U851 ( .A(w1055), .B(w1057), .Z(w1079) );
	XOR U852 ( .A(w995), .B(w994), .Z(w1080) );
	AND U853 ( .A(w1079), .B(w1080), .Z(w1081) );
	AND U854 ( .A(w1055), .B(w995), .Z(w1082) );
	XOR U855 ( .A(w1082), .B(w1081), .Z(w1083) );
	AND U856 ( .A(w1057), .B(w994), .Z(w1084) );
	XOR U857 ( .A(w1084), .B(w1081), .Z(w1085) );
	XOR U858 ( .A(w1062), .B(w1064), .Z(w1086) );
	XOR U859 ( .A(w993), .B(w992), .Z(w1087) );
	AND U860 ( .A(w1086), .B(w1087), .Z(w1088) );
	AND U861 ( .A(w1062), .B(w993), .Z(w1089) );
	XOR U862 ( .A(w1089), .B(w1088), .Z(w1090) );
	AND U863 ( .A(w1064), .B(w992), .Z(w1091) );
	XOR U864 ( .A(w1091), .B(w1088), .Z(w1092) );
	XOR U865 ( .A(w1085), .B(w1078), .Z(w1093) );
	XOR U866 ( .A(w1083), .B(w1077), .Z(w1094) );
	XOR U867 ( .A(w1092), .B(w1078), .Z(w1095) );
	XOR U868 ( .A(w1090), .B(w1077), .Z(w1096) );
	XOR U869 ( .A(w1057), .B(w1064), .Z(w1099) );
	XOR U870 ( .A(w1055), .B(w1062), .Z(w1100) );
	XOR U871 ( .A(w990), .B(w988), .Z(w1101) );
	XOR U872 ( .A(w991), .B(w989), .Z(w1102) );
	XOR U873 ( .A(w1100), .B(w1099), .Z(w1103) );
	XOR U874 ( .A(w1102), .B(w1101), .Z(w1104) );
	AND U875 ( .A(w1103), .B(w1104), .Z(w1105) );
	AND U876 ( .A(w1100), .B(w1102), .Z(w1106) );
	XOR U877 ( .A(w1106), .B(w1105), .Z(w1107) );
	AND U878 ( .A(w1099), .B(w1101), .Z(w1108) );
	XOR U879 ( .A(w1108), .B(w1105), .Z(w1109) );
	XOR U880 ( .A(w1109), .B(w1107), .Z(w1110) );
	XOR U881 ( .A(w1055), .B(w1057), .Z(w1111) );
	XOR U882 ( .A(w991), .B(w990), .Z(w1112) );
	AND U883 ( .A(w1111), .B(w1112), .Z(w1113) );
	AND U884 ( .A(w1055), .B(w991), .Z(w1114) );
	XOR U885 ( .A(w1114), .B(w1113), .Z(w1115) );
	AND U886 ( .A(w1057), .B(w990), .Z(w1116) );
	XOR U887 ( .A(w1116), .B(w1113), .Z(w1117) );
	XOR U888 ( .A(w1062), .B(w1064), .Z(w1118) );
	XOR U889 ( .A(w989), .B(w988), .Z(w1119) );
	AND U890 ( .A(w1118), .B(w1119), .Z(w1120) );
	AND U891 ( .A(w1062), .B(w989), .Z(w1121) );
	XOR U892 ( .A(w1121), .B(w1120), .Z(w1122) );
	AND U893 ( .A(w1064), .B(w988), .Z(w1123) );
	XOR U894 ( .A(w1123), .B(w1120), .Z(w1124) );
	XOR U895 ( .A(w1117), .B(w1110), .Z(w1125) );
	XOR U896 ( .A(w1115), .B(w1109), .Z(w1126) );
	XOR U897 ( .A(w1124), .B(w1110), .Z(w1127) );
	XOR U898 ( .A(w1122), .B(w1109), .Z(w1128) );
	XOR U899 ( .A(w1131), .B(w1127), .Z(w1137) );
	XOR U900 ( .A(w1132), .B(w1127), .Z(w1138) );
	XOR U901 ( .A(w1136), .B(w1127), .Z(w1139) );
	XOR U902 ( .A(w1129), .B(w1128), .Z(w1140) );
	XOR U903 ( .A(w1138), .B(w1128), .Z(w1141) );
	XOR U904 ( .A(w1133), .B(w1128), .Z(w1142) );
	XOR U905 ( .A(w1134), .B(w1128), .Z(w1143) );
	XOR U906 ( .A(w1135), .B(w1128), .Z(w1144) );
	XOR U907 ( .A(w1140), .B(w1125), .Z(w1145) );
	XOR U908 ( .A(w1137), .B(w1125), .Z(w1146) );
	XOR U909 ( .A(w1145), .B(w1126), .Z(w1147) );
	XOR U910 ( .A(w1130), .B(w1126), .Z(w1148) );
	XOR U911 ( .A(w1141), .B(w1126), .Z(w1149) );
	XOR U912 ( .A(w1143), .B(w1126), .Z(w1150) );
	XOR U913 ( .A(w1144), .B(w1126), .Z(w1151) );
	XOR U914 ( .A(w1139), .B(w1126), .Z(w1152) );
	XOR U915 ( .A(w1148), .B(w1095), .Z(w1153) );
	XOR U916 ( .A(w1142), .B(w1095), .Z(w1154) );
	XOR U917 ( .A(w1146), .B(w1096), .Z(w1155) );
	XOR U918 ( .A(w1147), .B(w1093), .Z(w1156) );
	XOR U919 ( .A(w1154), .B(w1093), .Z(w1157) );
	XOR U920 ( .A(w1151), .B(w1093), .Z(w1158) );
	XOR U921 ( .A(w1156), .B(w1094), .Z(w1159) );
	XOR U922 ( .A(w1153), .B(w1094), .Z(w1160) );
	XOR U923 ( .A(w1157), .B(w1094), .Z(w1161) );
	XOR U924 ( .A(w1158), .B(w1094), .Z(w1162) );
	XOR U925 ( .A(w1166), .B(w40), .Z(w1171) );
	XOR U926 ( .A(w1167), .B(w40), .Z(w1172) );
	XOR U927 ( .A(w1170), .B(w40), .Z(w1173) );
	XOR U928 ( .A(w1163), .B(w41), .Z(w1174) );
	XOR U929 ( .A(w1164), .B(w41), .Z(w1175) );
	XOR U930 ( .A(w1172), .B(w41), .Z(w1176) );
	XOR U931 ( .A(w1168), .B(w41), .Z(w1177) );
	XOR U932 ( .A(w1169), .B(w41), .Z(w1178) );
	XOR U933 ( .A(w1173), .B(w41), .Z(w1179) );
	XOR U934 ( .A(w1175), .B(w42), .Z(w1180) );
	XOR U935 ( .A(w1176), .B(w42), .Z(w1181) );
	XOR U936 ( .A(w1177), .B(w42), .Z(w1182) );
	XOR U937 ( .A(w1178), .B(w42), .Z(w1183) );
	XOR U938 ( .A(w1179), .B(w42), .Z(w1184) );
	XOR U939 ( .A(w1171), .B(w43), .Z(w1185) );
	XOR U940 ( .A(w1183), .B(w43), .Z(w1186) );
	XOR U941 ( .A(w1174), .B(w44), .Z(w1187) );
	XOR U942 ( .A(w1185), .B(w44), .Z(w1188) );
	XOR U943 ( .A(w1187), .B(w45), .Z(w1189) );
	XOR U944 ( .A(w1184), .B(w45), .Z(w1190) );
	XOR U945 ( .A(w1189), .B(w46), .Z(w1191) );
	XOR U946 ( .A(w1188), .B(w46), .Z(w1192) );
	XOR U947 ( .A(w1182), .B(w46), .Z(w1193) );
	XOR U948 ( .A(w1190), .B(w46), .Z(w1194) );
	XOR U949 ( .A(w1191), .B(w47), .Z(w1195) );
	XOR U950 ( .A(w1180), .B(w47), .Z(w1196) );
	XOR U951 ( .A(w1165), .B(w47), .Z(w1197) );
	XOR U952 ( .A(w1192), .B(w47), .Z(w1198) );
	XOR U953 ( .A(w1181), .B(w47), .Z(w1199) );
	XOR U954 ( .A(w1193), .B(w47), .Z(w1200) );
	XOR U955 ( .A(w1186), .B(w47), .Z(w1201) );
	XOR U956 ( .A(w1194), .B(w47), .Z(w1202) );
	XOR U957 ( .A(w1195), .B(w1199), .Z(w1203) );
	XOR U958 ( .A(w1196), .B(w1200), .Z(w1204) );
	XOR U959 ( .A(w1197), .B(w1201), .Z(w1205) );
	XOR U960 ( .A(w1198), .B(w1202), .Z(w1206) );
	XOR U961 ( .A(w1205), .B(w1203), .Z(w1207) );
	XOR U962 ( .A(w1206), .B(w1204), .Z(w1208) );
	XOR U963 ( .A(w1204), .B(w1203), .Z(w1209) );
	XOR U964 ( .A(w1197), .B(w1195), .Z(w1212) );
	XOR U965 ( .A(w1198), .B(w1196), .Z(w1213) );
	XOR U966 ( .A(w1201), .B(w1199), .Z(w1214) );
	XOR U967 ( .A(w1202), .B(w1200), .Z(w1215) );
	XOR U968 ( .A(w1213), .B(w1212), .Z(w1216) );
	XOR U969 ( .A(w1215), .B(w1214), .Z(w1217) );
	AND U970 ( .A(w1216), .B(w1217), .Z(w1218) );
	AND U971 ( .A(w1213), .B(w1215), .Z(w1219) );
	XOR U972 ( .A(w1219), .B(w1218), .Z(w1220) );
	AND U973 ( .A(w1212), .B(w1214), .Z(w1221) );
	XOR U974 ( .A(w1221), .B(w1218), .Z(w1222) );
	XOR U975 ( .A(w1222), .B(w1220), .Z(w1223) );
	XOR U976 ( .A(w1198), .B(w1197), .Z(w1224) );
	XOR U977 ( .A(w1202), .B(w1201), .Z(w1225) );
	AND U978 ( .A(w1224), .B(w1225), .Z(w1226) );
	AND U979 ( .A(w1198), .B(w1202), .Z(w1227) );
	XOR U980 ( .A(w1227), .B(w1226), .Z(w1228) );
	AND U981 ( .A(w1197), .B(w1201), .Z(w1229) );
	XOR U982 ( .A(w1229), .B(w1226), .Z(w1230) );
	XOR U983 ( .A(w1196), .B(w1195), .Z(w1231) );
	XOR U984 ( .A(w1200), .B(w1199), .Z(w1232) );
	AND U985 ( .A(w1231), .B(w1232), .Z(w1233) );
	AND U986 ( .A(w1196), .B(w1200), .Z(w1234) );
	XOR U987 ( .A(w1234), .B(w1233), .Z(w1235) );
	AND U988 ( .A(w1195), .B(w1199), .Z(w1236) );
	XOR U989 ( .A(w1236), .B(w1233), .Z(w1237) );
	XOR U990 ( .A(w1230), .B(w1223), .Z(w1238) );
	XOR U991 ( .A(w1228), .B(w1222), .Z(w1239) );
	XOR U992 ( .A(w1237), .B(w1223), .Z(w1240) );
	XOR U993 ( .A(w1235), .B(w1222), .Z(w1241) );
	XOR U994 ( .A(w1203), .B(w1240), .Z(w1242) );
	XOR U995 ( .A(w1209), .B(w1241), .Z(w1243) );
	XOR U996 ( .A(w1208), .B(w1238), .Z(w1244) );
	XOR U997 ( .A(w1207), .B(w1239), .Z(w1245) );
	XOR U998 ( .A(w1244), .B(w1242), .Z(w1246) );
	XOR U999 ( .A(w1245), .B(w1243), .Z(w1247) );
	XOR U1000 ( .A(w1247), .B(w1246), .Z(w1248) );
	XOR U1001 ( .A(w1245), .B(w1244), .Z(w1249) );
	XOR U1002 ( .A(w1243), .B(w1242), .Z(w1250) );
	AND U1003 ( .A(w1249), .B(w1250), .Z(w1251) );
	AND U1004 ( .A(w1245), .B(w1243), .Z(w1252) );
	XOR U1005 ( .A(w1252), .B(w1251), .Z(w1253) );
	AND U1006 ( .A(w1244), .B(w1242), .Z(w1254) );
	XOR U1007 ( .A(w1254), .B(w1251), .Z(w1255) );
	XOR U1008 ( .A(w1248), .B(w1255), .Z(w1256) );
	XOR U1009 ( .A(w1247), .B(w1253), .Z(w1257) );
	XOR U1010 ( .A(w1256), .B(w1257), .Z(w1258) );
	XOR U1011 ( .A(w1243), .B(w1242), .Z(w1259) );
	AND U1012 ( .A(w1258), .B(w1259), .Z(w1260) );
	AND U1013 ( .A(w1256), .B(w1243), .Z(w1261) );
	XOR U1014 ( .A(w1261), .B(w1260), .Z(w1262) );
	AND U1015 ( .A(w1257), .B(w1242), .Z(w1263) );
	XOR U1016 ( .A(w1263), .B(w1260), .Z(w1264) );
	XOR U1017 ( .A(w1256), .B(w1257), .Z(w1265) );
	XOR U1018 ( .A(w1245), .B(w1244), .Z(w1266) );
	AND U1019 ( .A(w1265), .B(w1266), .Z(w1267) );
	AND U1020 ( .A(w1256), .B(w1245), .Z(w1268) );
	XOR U1021 ( .A(w1268), .B(w1267), .Z(w1269) );
	AND U1022 ( .A(w1257), .B(w1244), .Z(w1270) );
	XOR U1023 ( .A(w1270), .B(w1267), .Z(w1271) );
	XOR U1024 ( .A(w1264), .B(w1271), .Z(w1274) );
	XOR U1025 ( .A(w1262), .B(w1269), .Z(w1275) );
	XOR U1026 ( .A(w1201), .B(w1199), .Z(w1276) );
	XOR U1027 ( .A(w1202), .B(w1200), .Z(w1277) );
	XOR U1028 ( .A(w1275), .B(w1274), .Z(w1278) );
	XOR U1029 ( .A(w1277), .B(w1276), .Z(w1279) );
	AND U1030 ( .A(w1278), .B(w1279), .Z(w1280) );
	AND U1031 ( .A(w1275), .B(w1277), .Z(w1281) );
	XOR U1032 ( .A(w1281), .B(w1280), .Z(w1282) );
	AND U1033 ( .A(w1274), .B(w1276), .Z(w1283) );
	XOR U1034 ( .A(w1283), .B(w1280), .Z(w1284) );
	XOR U1035 ( .A(w1284), .B(w1282), .Z(w1285) );
	XOR U1036 ( .A(w1262), .B(w1264), .Z(w1286) );
	XOR U1037 ( .A(w1202), .B(w1201), .Z(w1287) );
	AND U1038 ( .A(w1286), .B(w1287), .Z(w1288) );
	AND U1039 ( .A(w1262), .B(w1202), .Z(w1289) );
	XOR U1040 ( .A(w1289), .B(w1288), .Z(w1290) );
	AND U1041 ( .A(w1264), .B(w1201), .Z(w1291) );
	XOR U1042 ( .A(w1291), .B(w1288), .Z(w1292) );
	XOR U1043 ( .A(w1269), .B(w1271), .Z(w1293) );
	XOR U1044 ( .A(w1200), .B(w1199), .Z(w1294) );
	AND U1045 ( .A(w1293), .B(w1294), .Z(w1295) );
	AND U1046 ( .A(w1269), .B(w1200), .Z(w1296) );
	XOR U1047 ( .A(w1296), .B(w1295), .Z(w1297) );
	AND U1048 ( .A(w1271), .B(w1199), .Z(w1298) );
	XOR U1049 ( .A(w1298), .B(w1295), .Z(w1299) );
	XOR U1050 ( .A(w1292), .B(w1285), .Z(w1300) );
	XOR U1051 ( .A(w1290), .B(w1284), .Z(w1301) );
	XOR U1052 ( .A(w1299), .B(w1285), .Z(w1302) );
	XOR U1053 ( .A(w1297), .B(w1284), .Z(w1303) );
	XOR U1054 ( .A(w1264), .B(w1271), .Z(w1306) );
	XOR U1055 ( .A(w1262), .B(w1269), .Z(w1307) );
	XOR U1056 ( .A(w1197), .B(w1195), .Z(w1308) );
	XOR U1057 ( .A(w1198), .B(w1196), .Z(w1309) );
	XOR U1058 ( .A(w1307), .B(w1306), .Z(w1310) );
	XOR U1059 ( .A(w1309), .B(w1308), .Z(w1311) );
	AND U1060 ( .A(w1310), .B(w1311), .Z(w1312) );
	AND U1061 ( .A(w1307), .B(w1309), .Z(w1313) );
	XOR U1062 ( .A(w1313), .B(w1312), .Z(w1314) );
	AND U1063 ( .A(w1306), .B(w1308), .Z(w1315) );
	XOR U1064 ( .A(w1315), .B(w1312), .Z(w1316) );
	XOR U1065 ( .A(w1316), .B(w1314), .Z(w1317) );
	XOR U1066 ( .A(w1262), .B(w1264), .Z(w1318) );
	XOR U1067 ( .A(w1198), .B(w1197), .Z(w1319) );
	AND U1068 ( .A(w1318), .B(w1319), .Z(w1320) );
	AND U1069 ( .A(w1262), .B(w1198), .Z(w1321) );
	XOR U1070 ( .A(w1321), .B(w1320), .Z(w1322) );
	AND U1071 ( .A(w1264), .B(w1197), .Z(w1323) );
	XOR U1072 ( .A(w1323), .B(w1320), .Z(w1324) );
	XOR U1073 ( .A(w1269), .B(w1271), .Z(w1325) );
	XOR U1074 ( .A(w1196), .B(w1195), .Z(w1326) );
	AND U1075 ( .A(w1325), .B(w1326), .Z(w1327) );
	AND U1076 ( .A(w1269), .B(w1196), .Z(w1328) );
	XOR U1077 ( .A(w1328), .B(w1327), .Z(w1329) );
	AND U1078 ( .A(w1271), .B(w1195), .Z(w1330) );
	XOR U1079 ( .A(w1330), .B(w1327), .Z(w1331) );
	XOR U1080 ( .A(w1324), .B(w1317), .Z(w1332) );
	XOR U1081 ( .A(w1322), .B(w1316), .Z(w1333) );
	XOR U1082 ( .A(w1331), .B(w1317), .Z(w1334) );
	XOR U1083 ( .A(w1329), .B(w1316), .Z(w1335) );
	XOR U1084 ( .A(w1338), .B(w1334), .Z(w1344) );
	XOR U1085 ( .A(w1339), .B(w1334), .Z(w1345) );
	XOR U1086 ( .A(w1343), .B(w1334), .Z(w1346) );
	XOR U1087 ( .A(w1336), .B(w1335), .Z(w1347) );
	XOR U1088 ( .A(w1345), .B(w1335), .Z(w1348) );
	XOR U1089 ( .A(w1340), .B(w1335), .Z(w1349) );
	XOR U1090 ( .A(w1341), .B(w1335), .Z(w1350) );
	XOR U1091 ( .A(w1342), .B(w1335), .Z(w1351) );
	XOR U1092 ( .A(w1347), .B(w1332), .Z(w1352) );
	XOR U1093 ( .A(w1344), .B(w1332), .Z(w1353) );
	XOR U1094 ( .A(w1352), .B(w1333), .Z(w1354) );
	XOR U1095 ( .A(w1337), .B(w1333), .Z(w1355) );
	XOR U1096 ( .A(w1348), .B(w1333), .Z(w1356) );
	XOR U1097 ( .A(w1350), .B(w1333), .Z(w1357) );
	XOR U1098 ( .A(w1351), .B(w1333), .Z(w1358) );
	XOR U1099 ( .A(w1346), .B(w1333), .Z(w1359) );
	XOR U1100 ( .A(w1355), .B(w1302), .Z(w1360) );
	XOR U1101 ( .A(w1349), .B(w1302), .Z(w1361) );
	XOR U1102 ( .A(w1353), .B(w1303), .Z(w1362) );
	XOR U1103 ( .A(w1354), .B(w1300), .Z(w1363) );
	XOR U1104 ( .A(w1361), .B(w1300), .Z(w1364) );
	XOR U1105 ( .A(w1358), .B(w1300), .Z(w1365) );
	XOR U1106 ( .A(w1363), .B(w1301), .Z(w1366) );
	XOR U1107 ( .A(w1360), .B(w1301), .Z(w1367) );
	XOR U1108 ( .A(w1364), .B(w1301), .Z(w1368) );
	XOR U1109 ( .A(w1365), .B(w1301), .Z(w1369) );
	XOR U1110 ( .A(w1373), .B(w48), .Z(w1378) );
	XOR U1111 ( .A(w1374), .B(w48), .Z(w1379) );
	XOR U1112 ( .A(w1377), .B(w48), .Z(w1380) );
	XOR U1113 ( .A(w1370), .B(w49), .Z(w1381) );
	XOR U1114 ( .A(w1371), .B(w49), .Z(w1382) );
	XOR U1115 ( .A(w1379), .B(w49), .Z(w1383) );
	XOR U1116 ( .A(w1375), .B(w49), .Z(w1384) );
	XOR U1117 ( .A(w1376), .B(w49), .Z(w1385) );
	XOR U1118 ( .A(w1380), .B(w49), .Z(w1386) );
	XOR U1119 ( .A(w1382), .B(w50), .Z(w1387) );
	XOR U1120 ( .A(w1383), .B(w50), .Z(w1388) );
	XOR U1121 ( .A(w1384), .B(w50), .Z(w1389) );
	XOR U1122 ( .A(w1385), .B(w50), .Z(w1390) );
	XOR U1123 ( .A(w1386), .B(w50), .Z(w1391) );
	XOR U1124 ( .A(w1378), .B(w51), .Z(w1392) );
	XOR U1125 ( .A(w1390), .B(w51), .Z(w1393) );
	XOR U1126 ( .A(w1381), .B(w52), .Z(w1394) );
	XOR U1127 ( .A(w1392), .B(w52), .Z(w1395) );
	XOR U1128 ( .A(w1394), .B(w53), .Z(w1396) );
	XOR U1129 ( .A(w1391), .B(w53), .Z(w1397) );
	XOR U1130 ( .A(w1396), .B(w54), .Z(w1398) );
	XOR U1131 ( .A(w1395), .B(w54), .Z(w1399) );
	XOR U1132 ( .A(w1389), .B(w54), .Z(w1400) );
	XOR U1133 ( .A(w1397), .B(w54), .Z(w1401) );
	XOR U1134 ( .A(w1398), .B(w55), .Z(w1402) );
	XOR U1135 ( .A(w1387), .B(w55), .Z(w1403) );
	XOR U1136 ( .A(w1372), .B(w55), .Z(w1404) );
	XOR U1137 ( .A(w1399), .B(w55), .Z(w1405) );
	XOR U1138 ( .A(w1388), .B(w55), .Z(w1406) );
	XOR U1139 ( .A(w1400), .B(w55), .Z(w1407) );
	XOR U1140 ( .A(w1393), .B(w55), .Z(w1408) );
	XOR U1141 ( .A(w1401), .B(w55), .Z(w1409) );
	XOR U1142 ( .A(w1402), .B(w1406), .Z(w1410) );
	XOR U1143 ( .A(w1403), .B(w1407), .Z(w1411) );
	XOR U1144 ( .A(w1404), .B(w1408), .Z(w1412) );
	XOR U1145 ( .A(w1405), .B(w1409), .Z(w1413) );
	XOR U1146 ( .A(w1412), .B(w1410), .Z(w1414) );
	XOR U1147 ( .A(w1413), .B(w1411), .Z(w1415) );
	XOR U1148 ( .A(w1411), .B(w1410), .Z(w1416) );
	XOR U1149 ( .A(w1404), .B(w1402), .Z(w1419) );
	XOR U1150 ( .A(w1405), .B(w1403), .Z(w1420) );
	XOR U1151 ( .A(w1408), .B(w1406), .Z(w1421) );
	XOR U1152 ( .A(w1409), .B(w1407), .Z(w1422) );
	XOR U1153 ( .A(w1420), .B(w1419), .Z(w1423) );
	XOR U1154 ( .A(w1422), .B(w1421), .Z(w1424) );
	AND U1155 ( .A(w1423), .B(w1424), .Z(w1425) );
	AND U1156 ( .A(w1420), .B(w1422), .Z(w1426) );
	XOR U1157 ( .A(w1426), .B(w1425), .Z(w1427) );
	AND U1158 ( .A(w1419), .B(w1421), .Z(w1428) );
	XOR U1159 ( .A(w1428), .B(w1425), .Z(w1429) );
	XOR U1160 ( .A(w1429), .B(w1427), .Z(w1430) );
	XOR U1161 ( .A(w1405), .B(w1404), .Z(w1431) );
	XOR U1162 ( .A(w1409), .B(w1408), .Z(w1432) );
	AND U1163 ( .A(w1431), .B(w1432), .Z(w1433) );
	AND U1164 ( .A(w1405), .B(w1409), .Z(w1434) );
	XOR U1165 ( .A(w1434), .B(w1433), .Z(w1435) );
	AND U1166 ( .A(w1404), .B(w1408), .Z(w1436) );
	XOR U1167 ( .A(w1436), .B(w1433), .Z(w1437) );
	XOR U1168 ( .A(w1403), .B(w1402), .Z(w1438) );
	XOR U1169 ( .A(w1407), .B(w1406), .Z(w1439) );
	AND U1170 ( .A(w1438), .B(w1439), .Z(w1440) );
	AND U1171 ( .A(w1403), .B(w1407), .Z(w1441) );
	XOR U1172 ( .A(w1441), .B(w1440), .Z(w1442) );
	AND U1173 ( .A(w1402), .B(w1406), .Z(w1443) );
	XOR U1174 ( .A(w1443), .B(w1440), .Z(w1444) );
	XOR U1175 ( .A(w1437), .B(w1430), .Z(w1445) );
	XOR U1176 ( .A(w1435), .B(w1429), .Z(w1446) );
	XOR U1177 ( .A(w1444), .B(w1430), .Z(w1447) );
	XOR U1178 ( .A(w1442), .B(w1429), .Z(w1448) );
	XOR U1179 ( .A(w1410), .B(w1447), .Z(w1449) );
	XOR U1180 ( .A(w1416), .B(w1448), .Z(w1450) );
	XOR U1181 ( .A(w1415), .B(w1445), .Z(w1451) );
	XOR U1182 ( .A(w1414), .B(w1446), .Z(w1452) );
	XOR U1183 ( .A(w1451), .B(w1449), .Z(w1453) );
	XOR U1184 ( .A(w1452), .B(w1450), .Z(w1454) );
	XOR U1185 ( .A(w1454), .B(w1453), .Z(w1455) );
	XOR U1186 ( .A(w1452), .B(w1451), .Z(w1456) );
	XOR U1187 ( .A(w1450), .B(w1449), .Z(w1457) );
	AND U1188 ( .A(w1456), .B(w1457), .Z(w1458) );
	AND U1189 ( .A(w1452), .B(w1450), .Z(w1459) );
	XOR U1190 ( .A(w1459), .B(w1458), .Z(w1460) );
	AND U1191 ( .A(w1451), .B(w1449), .Z(w1461) );
	XOR U1192 ( .A(w1461), .B(w1458), .Z(w1462) );
	XOR U1193 ( .A(w1455), .B(w1462), .Z(w1463) );
	XOR U1194 ( .A(w1454), .B(w1460), .Z(w1464) );
	XOR U1195 ( .A(w1463), .B(w1464), .Z(w1465) );
	XOR U1196 ( .A(w1450), .B(w1449), .Z(w1466) );
	AND U1197 ( .A(w1465), .B(w1466), .Z(w1467) );
	AND U1198 ( .A(w1463), .B(w1450), .Z(w1468) );
	XOR U1199 ( .A(w1468), .B(w1467), .Z(w1469) );
	AND U1200 ( .A(w1464), .B(w1449), .Z(w1470) );
	XOR U1201 ( .A(w1470), .B(w1467), .Z(w1471) );
	XOR U1202 ( .A(w1463), .B(w1464), .Z(w1472) );
	XOR U1203 ( .A(w1452), .B(w1451), .Z(w1473) );
	AND U1204 ( .A(w1472), .B(w1473), .Z(w1474) );
	AND U1205 ( .A(w1463), .B(w1452), .Z(w1475) );
	XOR U1206 ( .A(w1475), .B(w1474), .Z(w1476) );
	AND U1207 ( .A(w1464), .B(w1451), .Z(w1477) );
	XOR U1208 ( .A(w1477), .B(w1474), .Z(w1478) );
	XOR U1209 ( .A(w1471), .B(w1478), .Z(w1481) );
	XOR U1210 ( .A(w1469), .B(w1476), .Z(w1482) );
	XOR U1211 ( .A(w1408), .B(w1406), .Z(w1483) );
	XOR U1212 ( .A(w1409), .B(w1407), .Z(w1484) );
	XOR U1213 ( .A(w1482), .B(w1481), .Z(w1485) );
	XOR U1214 ( .A(w1484), .B(w1483), .Z(w1486) );
	AND U1215 ( .A(w1485), .B(w1486), .Z(w1487) );
	AND U1216 ( .A(w1482), .B(w1484), .Z(w1488) );
	XOR U1217 ( .A(w1488), .B(w1487), .Z(w1489) );
	AND U1218 ( .A(w1481), .B(w1483), .Z(w1490) );
	XOR U1219 ( .A(w1490), .B(w1487), .Z(w1491) );
	XOR U1220 ( .A(w1491), .B(w1489), .Z(w1492) );
	XOR U1221 ( .A(w1469), .B(w1471), .Z(w1493) );
	XOR U1222 ( .A(w1409), .B(w1408), .Z(w1494) );
	AND U1223 ( .A(w1493), .B(w1494), .Z(w1495) );
	AND U1224 ( .A(w1469), .B(w1409), .Z(w1496) );
	XOR U1225 ( .A(w1496), .B(w1495), .Z(w1497) );
	AND U1226 ( .A(w1471), .B(w1408), .Z(w1498) );
	XOR U1227 ( .A(w1498), .B(w1495), .Z(w1499) );
	XOR U1228 ( .A(w1476), .B(w1478), .Z(w1500) );
	XOR U1229 ( .A(w1407), .B(w1406), .Z(w1501) );
	AND U1230 ( .A(w1500), .B(w1501), .Z(w1502) );
	AND U1231 ( .A(w1476), .B(w1407), .Z(w1503) );
	XOR U1232 ( .A(w1503), .B(w1502), .Z(w1504) );
	AND U1233 ( .A(w1478), .B(w1406), .Z(w1505) );
	XOR U1234 ( .A(w1505), .B(w1502), .Z(w1506) );
	XOR U1235 ( .A(w1499), .B(w1492), .Z(w1507) );
	XOR U1236 ( .A(w1497), .B(w1491), .Z(w1508) );
	XOR U1237 ( .A(w1506), .B(w1492), .Z(w1509) );
	XOR U1238 ( .A(w1504), .B(w1491), .Z(w1510) );
	XOR U1239 ( .A(w1471), .B(w1478), .Z(w1513) );
	XOR U1240 ( .A(w1469), .B(w1476), .Z(w1514) );
	XOR U1241 ( .A(w1404), .B(w1402), .Z(w1515) );
	XOR U1242 ( .A(w1405), .B(w1403), .Z(w1516) );
	XOR U1243 ( .A(w1514), .B(w1513), .Z(w1517) );
	XOR U1244 ( .A(w1516), .B(w1515), .Z(w1518) );
	AND U1245 ( .A(w1517), .B(w1518), .Z(w1519) );
	AND U1246 ( .A(w1514), .B(w1516), .Z(w1520) );
	XOR U1247 ( .A(w1520), .B(w1519), .Z(w1521) );
	AND U1248 ( .A(w1513), .B(w1515), .Z(w1522) );
	XOR U1249 ( .A(w1522), .B(w1519), .Z(w1523) );
	XOR U1250 ( .A(w1523), .B(w1521), .Z(w1524) );
	XOR U1251 ( .A(w1469), .B(w1471), .Z(w1525) );
	XOR U1252 ( .A(w1405), .B(w1404), .Z(w1526) );
	AND U1253 ( .A(w1525), .B(w1526), .Z(w1527) );
	AND U1254 ( .A(w1469), .B(w1405), .Z(w1528) );
	XOR U1255 ( .A(w1528), .B(w1527), .Z(w1529) );
	AND U1256 ( .A(w1471), .B(w1404), .Z(w1530) );
	XOR U1257 ( .A(w1530), .B(w1527), .Z(w1531) );
	XOR U1258 ( .A(w1476), .B(w1478), .Z(w1532) );
	XOR U1259 ( .A(w1403), .B(w1402), .Z(w1533) );
	AND U1260 ( .A(w1532), .B(w1533), .Z(w1534) );
	AND U1261 ( .A(w1476), .B(w1403), .Z(w1535) );
	XOR U1262 ( .A(w1535), .B(w1534), .Z(w1536) );
	AND U1263 ( .A(w1478), .B(w1402), .Z(w1537) );
	XOR U1264 ( .A(w1537), .B(w1534), .Z(w1538) );
	XOR U1265 ( .A(w1531), .B(w1524), .Z(w1539) );
	XOR U1266 ( .A(w1529), .B(w1523), .Z(w1540) );
	XOR U1267 ( .A(w1538), .B(w1524), .Z(w1541) );
	XOR U1268 ( .A(w1536), .B(w1523), .Z(w1542) );
	XOR U1269 ( .A(w1545), .B(w1541), .Z(w1551) );
	XOR U1270 ( .A(w1546), .B(w1541), .Z(w1552) );
	XOR U1271 ( .A(w1550), .B(w1541), .Z(w1553) );
	XOR U1272 ( .A(w1543), .B(w1542), .Z(w1554) );
	XOR U1273 ( .A(w1552), .B(w1542), .Z(w1555) );
	XOR U1274 ( .A(w1547), .B(w1542), .Z(w1556) );
	XOR U1275 ( .A(w1548), .B(w1542), .Z(w1557) );
	XOR U1276 ( .A(w1549), .B(w1542), .Z(w1558) );
	XOR U1277 ( .A(w1554), .B(w1539), .Z(w1559) );
	XOR U1278 ( .A(w1551), .B(w1539), .Z(w1560) );
	XOR U1279 ( .A(w1559), .B(w1540), .Z(w1561) );
	XOR U1280 ( .A(w1544), .B(w1540), .Z(w1562) );
	XOR U1281 ( .A(w1555), .B(w1540), .Z(w1563) );
	XOR U1282 ( .A(w1557), .B(w1540), .Z(w1564) );
	XOR U1283 ( .A(w1558), .B(w1540), .Z(w1565) );
	XOR U1284 ( .A(w1553), .B(w1540), .Z(w1566) );
	XOR U1285 ( .A(w1562), .B(w1509), .Z(w1567) );
	XOR U1286 ( .A(w1556), .B(w1509), .Z(w1568) );
	XOR U1287 ( .A(w1560), .B(w1510), .Z(w1569) );
	XOR U1288 ( .A(w1561), .B(w1507), .Z(w1570) );
	XOR U1289 ( .A(w1568), .B(w1507), .Z(w1571) );
	XOR U1290 ( .A(w1565), .B(w1507), .Z(w1572) );
	XOR U1291 ( .A(w1570), .B(w1508), .Z(w1573) );
	XOR U1292 ( .A(w1567), .B(w1508), .Z(w1574) );
	XOR U1293 ( .A(w1571), .B(w1508), .Z(w1575) );
	XOR U1294 ( .A(w1572), .B(w1508), .Z(w1576) );
	XOR U1295 ( .A(w1580), .B(w56), .Z(w1585) );
	XOR U1296 ( .A(w1581), .B(w56), .Z(w1586) );
	XOR U1297 ( .A(w1584), .B(w56), .Z(w1587) );
	XOR U1298 ( .A(w1577), .B(w57), .Z(w1588) );
	XOR U1299 ( .A(w1578), .B(w57), .Z(w1589) );
	XOR U1300 ( .A(w1586), .B(w57), .Z(w1590) );
	XOR U1301 ( .A(w1582), .B(w57), .Z(w1591) );
	XOR U1302 ( .A(w1583), .B(w57), .Z(w1592) );
	XOR U1303 ( .A(w1587), .B(w57), .Z(w1593) );
	XOR U1304 ( .A(w1589), .B(w58), .Z(w1594) );
	XOR U1305 ( .A(w1590), .B(w58), .Z(w1595) );
	XOR U1306 ( .A(w1591), .B(w58), .Z(w1596) );
	XOR U1307 ( .A(w1592), .B(w58), .Z(w1597) );
	XOR U1308 ( .A(w1593), .B(w58), .Z(w1598) );
	XOR U1309 ( .A(w1585), .B(w59), .Z(w1599) );
	XOR U1310 ( .A(w1597), .B(w59), .Z(w1600) );
	XOR U1311 ( .A(w1588), .B(w60), .Z(w1601) );
	XOR U1312 ( .A(w1599), .B(w60), .Z(w1602) );
	XOR U1313 ( .A(w1601), .B(w61), .Z(w1603) );
	XOR U1314 ( .A(w1598), .B(w61), .Z(w1604) );
	XOR U1315 ( .A(w1603), .B(w62), .Z(w1605) );
	XOR U1316 ( .A(w1602), .B(w62), .Z(w1606) );
	XOR U1317 ( .A(w1596), .B(w62), .Z(w1607) );
	XOR U1318 ( .A(w1604), .B(w62), .Z(w1608) );
	XOR U1319 ( .A(w1605), .B(w63), .Z(w1609) );
	XOR U1320 ( .A(w1594), .B(w63), .Z(w1610) );
	XOR U1321 ( .A(w1579), .B(w63), .Z(w1611) );
	XOR U1322 ( .A(w1606), .B(w63), .Z(w1612) );
	XOR U1323 ( .A(w1595), .B(w63), .Z(w1613) );
	XOR U1324 ( .A(w1607), .B(w63), .Z(w1614) );
	XOR U1325 ( .A(w1600), .B(w63), .Z(w1615) );
	XOR U1326 ( .A(w1608), .B(w63), .Z(w1616) );
	XOR U1327 ( .A(w1609), .B(w1613), .Z(w1617) );
	XOR U1328 ( .A(w1610), .B(w1614), .Z(w1618) );
	XOR U1329 ( .A(w1611), .B(w1615), .Z(w1619) );
	XOR U1330 ( .A(w1612), .B(w1616), .Z(w1620) );
	XOR U1331 ( .A(w1619), .B(w1617), .Z(w1621) );
	XOR U1332 ( .A(w1620), .B(w1618), .Z(w1622) );
	XOR U1333 ( .A(w1618), .B(w1617), .Z(w1623) );
	XOR U1334 ( .A(w1611), .B(w1609), .Z(w1626) );
	XOR U1335 ( .A(w1612), .B(w1610), .Z(w1627) );
	XOR U1336 ( .A(w1615), .B(w1613), .Z(w1628) );
	XOR U1337 ( .A(w1616), .B(w1614), .Z(w1629) );
	XOR U1338 ( .A(w1627), .B(w1626), .Z(w1630) );
	XOR U1339 ( .A(w1629), .B(w1628), .Z(w1631) );
	AND U1340 ( .A(w1630), .B(w1631), .Z(w1632) );
	AND U1341 ( .A(w1627), .B(w1629), .Z(w1633) );
	XOR U1342 ( .A(w1633), .B(w1632), .Z(w1634) );
	AND U1343 ( .A(w1626), .B(w1628), .Z(w1635) );
	XOR U1344 ( .A(w1635), .B(w1632), .Z(w1636) );
	XOR U1345 ( .A(w1636), .B(w1634), .Z(w1637) );
	XOR U1346 ( .A(w1612), .B(w1611), .Z(w1638) );
	XOR U1347 ( .A(w1616), .B(w1615), .Z(w1639) );
	AND U1348 ( .A(w1638), .B(w1639), .Z(w1640) );
	AND U1349 ( .A(w1612), .B(w1616), .Z(w1641) );
	XOR U1350 ( .A(w1641), .B(w1640), .Z(w1642) );
	AND U1351 ( .A(w1611), .B(w1615), .Z(w1643) );
	XOR U1352 ( .A(w1643), .B(w1640), .Z(w1644) );
	XOR U1353 ( .A(w1610), .B(w1609), .Z(w1645) );
	XOR U1354 ( .A(w1614), .B(w1613), .Z(w1646) );
	AND U1355 ( .A(w1645), .B(w1646), .Z(w1647) );
	AND U1356 ( .A(w1610), .B(w1614), .Z(w1648) );
	XOR U1357 ( .A(w1648), .B(w1647), .Z(w1649) );
	AND U1358 ( .A(w1609), .B(w1613), .Z(w1650) );
	XOR U1359 ( .A(w1650), .B(w1647), .Z(w1651) );
	XOR U1360 ( .A(w1644), .B(w1637), .Z(w1652) );
	XOR U1361 ( .A(w1642), .B(w1636), .Z(w1653) );
	XOR U1362 ( .A(w1651), .B(w1637), .Z(w1654) );
	XOR U1363 ( .A(w1649), .B(w1636), .Z(w1655) );
	XOR U1364 ( .A(w1617), .B(w1654), .Z(w1656) );
	XOR U1365 ( .A(w1623), .B(w1655), .Z(w1657) );
	XOR U1366 ( .A(w1622), .B(w1652), .Z(w1658) );
	XOR U1367 ( .A(w1621), .B(w1653), .Z(w1659) );
	XOR U1368 ( .A(w1658), .B(w1656), .Z(w1660) );
	XOR U1369 ( .A(w1659), .B(w1657), .Z(w1661) );
	XOR U1370 ( .A(w1661), .B(w1660), .Z(w1662) );
	XOR U1371 ( .A(w1659), .B(w1658), .Z(w1663) );
	XOR U1372 ( .A(w1657), .B(w1656), .Z(w1664) );
	AND U1373 ( .A(w1663), .B(w1664), .Z(w1665) );
	AND U1374 ( .A(w1659), .B(w1657), .Z(w1666) );
	XOR U1375 ( .A(w1666), .B(w1665), .Z(w1667) );
	AND U1376 ( .A(w1658), .B(w1656), .Z(w1668) );
	XOR U1377 ( .A(w1668), .B(w1665), .Z(w1669) );
	XOR U1378 ( .A(w1662), .B(w1669), .Z(w1670) );
	XOR U1379 ( .A(w1661), .B(w1667), .Z(w1671) );
	XOR U1380 ( .A(w1670), .B(w1671), .Z(w1672) );
	XOR U1381 ( .A(w1657), .B(w1656), .Z(w1673) );
	AND U1382 ( .A(w1672), .B(w1673), .Z(w1674) );
	AND U1383 ( .A(w1670), .B(w1657), .Z(w1675) );
	XOR U1384 ( .A(w1675), .B(w1674), .Z(w1676) );
	AND U1385 ( .A(w1671), .B(w1656), .Z(w1677) );
	XOR U1386 ( .A(w1677), .B(w1674), .Z(w1678) );
	XOR U1387 ( .A(w1670), .B(w1671), .Z(w1679) );
	XOR U1388 ( .A(w1659), .B(w1658), .Z(w1680) );
	AND U1389 ( .A(w1679), .B(w1680), .Z(w1681) );
	AND U1390 ( .A(w1670), .B(w1659), .Z(w1682) );
	XOR U1391 ( .A(w1682), .B(w1681), .Z(w1683) );
	AND U1392 ( .A(w1671), .B(w1658), .Z(w1684) );
	XOR U1393 ( .A(w1684), .B(w1681), .Z(w1685) );
	XOR U1394 ( .A(w1678), .B(w1685), .Z(w1688) );
	XOR U1395 ( .A(w1676), .B(w1683), .Z(w1689) );
	XOR U1396 ( .A(w1615), .B(w1613), .Z(w1690) );
	XOR U1397 ( .A(w1616), .B(w1614), .Z(w1691) );
	XOR U1398 ( .A(w1689), .B(w1688), .Z(w1692) );
	XOR U1399 ( .A(w1691), .B(w1690), .Z(w1693) );
	AND U1400 ( .A(w1692), .B(w1693), .Z(w1694) );
	AND U1401 ( .A(w1689), .B(w1691), .Z(w1695) );
	XOR U1402 ( .A(w1695), .B(w1694), .Z(w1696) );
	AND U1403 ( .A(w1688), .B(w1690), .Z(w1697) );
	XOR U1404 ( .A(w1697), .B(w1694), .Z(w1698) );
	XOR U1405 ( .A(w1698), .B(w1696), .Z(w1699) );
	XOR U1406 ( .A(w1676), .B(w1678), .Z(w1700) );
	XOR U1407 ( .A(w1616), .B(w1615), .Z(w1701) );
	AND U1408 ( .A(w1700), .B(w1701), .Z(w1702) );
	AND U1409 ( .A(w1676), .B(w1616), .Z(w1703) );
	XOR U1410 ( .A(w1703), .B(w1702), .Z(w1704) );
	AND U1411 ( .A(w1678), .B(w1615), .Z(w1705) );
	XOR U1412 ( .A(w1705), .B(w1702), .Z(w1706) );
	XOR U1413 ( .A(w1683), .B(w1685), .Z(w1707) );
	XOR U1414 ( .A(w1614), .B(w1613), .Z(w1708) );
	AND U1415 ( .A(w1707), .B(w1708), .Z(w1709) );
	AND U1416 ( .A(w1683), .B(w1614), .Z(w1710) );
	XOR U1417 ( .A(w1710), .B(w1709), .Z(w1711) );
	AND U1418 ( .A(w1685), .B(w1613), .Z(w1712) );
	XOR U1419 ( .A(w1712), .B(w1709), .Z(w1713) );
	XOR U1420 ( .A(w1706), .B(w1699), .Z(w1714) );
	XOR U1421 ( .A(w1704), .B(w1698), .Z(w1715) );
	XOR U1422 ( .A(w1713), .B(w1699), .Z(w1716) );
	XOR U1423 ( .A(w1711), .B(w1698), .Z(w1717) );
	XOR U1424 ( .A(w1678), .B(w1685), .Z(w1720) );
	XOR U1425 ( .A(w1676), .B(w1683), .Z(w1721) );
	XOR U1426 ( .A(w1611), .B(w1609), .Z(w1722) );
	XOR U1427 ( .A(w1612), .B(w1610), .Z(w1723) );
	XOR U1428 ( .A(w1721), .B(w1720), .Z(w1724) );
	XOR U1429 ( .A(w1723), .B(w1722), .Z(w1725) );
	AND U1430 ( .A(w1724), .B(w1725), .Z(w1726) );
	AND U1431 ( .A(w1721), .B(w1723), .Z(w1727) );
	XOR U1432 ( .A(w1727), .B(w1726), .Z(w1728) );
	AND U1433 ( .A(w1720), .B(w1722), .Z(w1729) );
	XOR U1434 ( .A(w1729), .B(w1726), .Z(w1730) );
	XOR U1435 ( .A(w1730), .B(w1728), .Z(w1731) );
	XOR U1436 ( .A(w1676), .B(w1678), .Z(w1732) );
	XOR U1437 ( .A(w1612), .B(w1611), .Z(w1733) );
	AND U1438 ( .A(w1732), .B(w1733), .Z(w1734) );
	AND U1439 ( .A(w1676), .B(w1612), .Z(w1735) );
	XOR U1440 ( .A(w1735), .B(w1734), .Z(w1736) );
	AND U1441 ( .A(w1678), .B(w1611), .Z(w1737) );
	XOR U1442 ( .A(w1737), .B(w1734), .Z(w1738) );
	XOR U1443 ( .A(w1683), .B(w1685), .Z(w1739) );
	XOR U1444 ( .A(w1610), .B(w1609), .Z(w1740) );
	AND U1445 ( .A(w1739), .B(w1740), .Z(w1741) );
	AND U1446 ( .A(w1683), .B(w1610), .Z(w1742) );
	XOR U1447 ( .A(w1742), .B(w1741), .Z(w1743) );
	AND U1448 ( .A(w1685), .B(w1609), .Z(w1744) );
	XOR U1449 ( .A(w1744), .B(w1741), .Z(w1745) );
	XOR U1450 ( .A(w1738), .B(w1731), .Z(w1746) );
	XOR U1451 ( .A(w1736), .B(w1730), .Z(w1747) );
	XOR U1452 ( .A(w1745), .B(w1731), .Z(w1748) );
	XOR U1453 ( .A(w1743), .B(w1730), .Z(w1749) );
	XOR U1454 ( .A(w1752), .B(w1748), .Z(w1758) );
	XOR U1455 ( .A(w1753), .B(w1748), .Z(w1759) );
	XOR U1456 ( .A(w1757), .B(w1748), .Z(w1760) );
	XOR U1457 ( .A(w1750), .B(w1749), .Z(w1761) );
	XOR U1458 ( .A(w1759), .B(w1749), .Z(w1762) );
	XOR U1459 ( .A(w1754), .B(w1749), .Z(w1763) );
	XOR U1460 ( .A(w1755), .B(w1749), .Z(w1764) );
	XOR U1461 ( .A(w1756), .B(w1749), .Z(w1765) );
	XOR U1462 ( .A(w1761), .B(w1746), .Z(w1766) );
	XOR U1463 ( .A(w1758), .B(w1746), .Z(w1767) );
	XOR U1464 ( .A(w1766), .B(w1747), .Z(w1768) );
	XOR U1465 ( .A(w1751), .B(w1747), .Z(w1769) );
	XOR U1466 ( .A(w1762), .B(w1747), .Z(w1770) );
	XOR U1467 ( .A(w1764), .B(w1747), .Z(w1771) );
	XOR U1468 ( .A(w1765), .B(w1747), .Z(w1772) );
	XOR U1469 ( .A(w1760), .B(w1747), .Z(w1773) );
	XOR U1470 ( .A(w1769), .B(w1716), .Z(w1774) );
	XOR U1471 ( .A(w1763), .B(w1716), .Z(w1775) );
	XOR U1472 ( .A(w1767), .B(w1717), .Z(w1776) );
	XOR U1473 ( .A(w1768), .B(w1714), .Z(w1777) );
	XOR U1474 ( .A(w1775), .B(w1714), .Z(w1778) );
	XOR U1475 ( .A(w1772), .B(w1714), .Z(w1779) );
	XOR U1476 ( .A(w1777), .B(w1715), .Z(w1780) );
	XOR U1477 ( .A(w1774), .B(w1715), .Z(w1781) );
	XOR U1478 ( .A(w1778), .B(w1715), .Z(w1782) );
	XOR U1479 ( .A(w1779), .B(w1715), .Z(w1783) );
	XOR U1480 ( .A(w1787), .B(w64), .Z(w1792) );
	XOR U1481 ( .A(w1788), .B(w64), .Z(w1793) );
	XOR U1482 ( .A(w1791), .B(w64), .Z(w1794) );
	XOR U1483 ( .A(w1784), .B(w65), .Z(w1795) );
	XOR U1484 ( .A(w1785), .B(w65), .Z(w1796) );
	XOR U1485 ( .A(w1793), .B(w65), .Z(w1797) );
	XOR U1486 ( .A(w1789), .B(w65), .Z(w1798) );
	XOR U1487 ( .A(w1790), .B(w65), .Z(w1799) );
	XOR U1488 ( .A(w1794), .B(w65), .Z(w1800) );
	XOR U1489 ( .A(w1796), .B(w66), .Z(w1801) );
	XOR U1490 ( .A(w1797), .B(w66), .Z(w1802) );
	XOR U1491 ( .A(w1798), .B(w66), .Z(w1803) );
	XOR U1492 ( .A(w1799), .B(w66), .Z(w1804) );
	XOR U1493 ( .A(w1800), .B(w66), .Z(w1805) );
	XOR U1494 ( .A(w1792), .B(w67), .Z(w1806) );
	XOR U1495 ( .A(w1804), .B(w67), .Z(w1807) );
	XOR U1496 ( .A(w1795), .B(w68), .Z(w1808) );
	XOR U1497 ( .A(w1806), .B(w68), .Z(w1809) );
	XOR U1498 ( .A(w1808), .B(w69), .Z(w1810) );
	XOR U1499 ( .A(w1805), .B(w69), .Z(w1811) );
	XOR U1500 ( .A(w1810), .B(w70), .Z(w1812) );
	XOR U1501 ( .A(w1809), .B(w70), .Z(w1813) );
	XOR U1502 ( .A(w1803), .B(w70), .Z(w1814) );
	XOR U1503 ( .A(w1811), .B(w70), .Z(w1815) );
	XOR U1504 ( .A(w1812), .B(w71), .Z(w1816) );
	XOR U1505 ( .A(w1801), .B(w71), .Z(w1817) );
	XOR U1506 ( .A(w1786), .B(w71), .Z(w1818) );
	XOR U1507 ( .A(w1813), .B(w71), .Z(w1819) );
	XOR U1508 ( .A(w1802), .B(w71), .Z(w1820) );
	XOR U1509 ( .A(w1814), .B(w71), .Z(w1821) );
	XOR U1510 ( .A(w1807), .B(w71), .Z(w1822) );
	XOR U1511 ( .A(w1815), .B(w71), .Z(w1823) );
	XOR U1512 ( .A(w1816), .B(w1820), .Z(w1824) );
	XOR U1513 ( .A(w1817), .B(w1821), .Z(w1825) );
	XOR U1514 ( .A(w1818), .B(w1822), .Z(w1826) );
	XOR U1515 ( .A(w1819), .B(w1823), .Z(w1827) );
	XOR U1516 ( .A(w1826), .B(w1824), .Z(w1828) );
	XOR U1517 ( .A(w1827), .B(w1825), .Z(w1829) );
	XOR U1518 ( .A(w1825), .B(w1824), .Z(w1830) );
	XOR U1519 ( .A(w1818), .B(w1816), .Z(w1833) );
	XOR U1520 ( .A(w1819), .B(w1817), .Z(w1834) );
	XOR U1521 ( .A(w1822), .B(w1820), .Z(w1835) );
	XOR U1522 ( .A(w1823), .B(w1821), .Z(w1836) );
	XOR U1523 ( .A(w1834), .B(w1833), .Z(w1837) );
	XOR U1524 ( .A(w1836), .B(w1835), .Z(w1838) );
	AND U1525 ( .A(w1837), .B(w1838), .Z(w1839) );
	AND U1526 ( .A(w1834), .B(w1836), .Z(w1840) );
	XOR U1527 ( .A(w1840), .B(w1839), .Z(w1841) );
	AND U1528 ( .A(w1833), .B(w1835), .Z(w1842) );
	XOR U1529 ( .A(w1842), .B(w1839), .Z(w1843) );
	XOR U1530 ( .A(w1843), .B(w1841), .Z(w1844) );
	XOR U1531 ( .A(w1819), .B(w1818), .Z(w1845) );
	XOR U1532 ( .A(w1823), .B(w1822), .Z(w1846) );
	AND U1533 ( .A(w1845), .B(w1846), .Z(w1847) );
	AND U1534 ( .A(w1819), .B(w1823), .Z(w1848) );
	XOR U1535 ( .A(w1848), .B(w1847), .Z(w1849) );
	AND U1536 ( .A(w1818), .B(w1822), .Z(w1850) );
	XOR U1537 ( .A(w1850), .B(w1847), .Z(w1851) );
	XOR U1538 ( .A(w1817), .B(w1816), .Z(w1852) );
	XOR U1539 ( .A(w1821), .B(w1820), .Z(w1853) );
	AND U1540 ( .A(w1852), .B(w1853), .Z(w1854) );
	AND U1541 ( .A(w1817), .B(w1821), .Z(w1855) );
	XOR U1542 ( .A(w1855), .B(w1854), .Z(w1856) );
	AND U1543 ( .A(w1816), .B(w1820), .Z(w1857) );
	XOR U1544 ( .A(w1857), .B(w1854), .Z(w1858) );
	XOR U1545 ( .A(w1851), .B(w1844), .Z(w1859) );
	XOR U1546 ( .A(w1849), .B(w1843), .Z(w1860) );
	XOR U1547 ( .A(w1858), .B(w1844), .Z(w1861) );
	XOR U1548 ( .A(w1856), .B(w1843), .Z(w1862) );
	XOR U1549 ( .A(w1824), .B(w1861), .Z(w1863) );
	XOR U1550 ( .A(w1830), .B(w1862), .Z(w1864) );
	XOR U1551 ( .A(w1829), .B(w1859), .Z(w1865) );
	XOR U1552 ( .A(w1828), .B(w1860), .Z(w1866) );
	XOR U1553 ( .A(w1865), .B(w1863), .Z(w1867) );
	XOR U1554 ( .A(w1866), .B(w1864), .Z(w1868) );
	XOR U1555 ( .A(w1868), .B(w1867), .Z(w1869) );
	XOR U1556 ( .A(w1866), .B(w1865), .Z(w1870) );
	XOR U1557 ( .A(w1864), .B(w1863), .Z(w1871) );
	AND U1558 ( .A(w1870), .B(w1871), .Z(w1872) );
	AND U1559 ( .A(w1866), .B(w1864), .Z(w1873) );
	XOR U1560 ( .A(w1873), .B(w1872), .Z(w1874) );
	AND U1561 ( .A(w1865), .B(w1863), .Z(w1875) );
	XOR U1562 ( .A(w1875), .B(w1872), .Z(w1876) );
	XOR U1563 ( .A(w1869), .B(w1876), .Z(w1877) );
	XOR U1564 ( .A(w1868), .B(w1874), .Z(w1878) );
	XOR U1565 ( .A(w1877), .B(w1878), .Z(w1879) );
	XOR U1566 ( .A(w1864), .B(w1863), .Z(w1880) );
	AND U1567 ( .A(w1879), .B(w1880), .Z(w1881) );
	AND U1568 ( .A(w1877), .B(w1864), .Z(w1882) );
	XOR U1569 ( .A(w1882), .B(w1881), .Z(w1883) );
	AND U1570 ( .A(w1878), .B(w1863), .Z(w1884) );
	XOR U1571 ( .A(w1884), .B(w1881), .Z(w1885) );
	XOR U1572 ( .A(w1877), .B(w1878), .Z(w1886) );
	XOR U1573 ( .A(w1866), .B(w1865), .Z(w1887) );
	AND U1574 ( .A(w1886), .B(w1887), .Z(w1888) );
	AND U1575 ( .A(w1877), .B(w1866), .Z(w1889) );
	XOR U1576 ( .A(w1889), .B(w1888), .Z(w1890) );
	AND U1577 ( .A(w1878), .B(w1865), .Z(w1891) );
	XOR U1578 ( .A(w1891), .B(w1888), .Z(w1892) );
	XOR U1579 ( .A(w1885), .B(w1892), .Z(w1895) );
	XOR U1580 ( .A(w1883), .B(w1890), .Z(w1896) );
	XOR U1581 ( .A(w1822), .B(w1820), .Z(w1897) );
	XOR U1582 ( .A(w1823), .B(w1821), .Z(w1898) );
	XOR U1583 ( .A(w1896), .B(w1895), .Z(w1899) );
	XOR U1584 ( .A(w1898), .B(w1897), .Z(w1900) );
	AND U1585 ( .A(w1899), .B(w1900), .Z(w1901) );
	AND U1586 ( .A(w1896), .B(w1898), .Z(w1902) );
	XOR U1587 ( .A(w1902), .B(w1901), .Z(w1903) );
	AND U1588 ( .A(w1895), .B(w1897), .Z(w1904) );
	XOR U1589 ( .A(w1904), .B(w1901), .Z(w1905) );
	XOR U1590 ( .A(w1905), .B(w1903), .Z(w1906) );
	XOR U1591 ( .A(w1883), .B(w1885), .Z(w1907) );
	XOR U1592 ( .A(w1823), .B(w1822), .Z(w1908) );
	AND U1593 ( .A(w1907), .B(w1908), .Z(w1909) );
	AND U1594 ( .A(w1883), .B(w1823), .Z(w1910) );
	XOR U1595 ( .A(w1910), .B(w1909), .Z(w1911) );
	AND U1596 ( .A(w1885), .B(w1822), .Z(w1912) );
	XOR U1597 ( .A(w1912), .B(w1909), .Z(w1913) );
	XOR U1598 ( .A(w1890), .B(w1892), .Z(w1914) );
	XOR U1599 ( .A(w1821), .B(w1820), .Z(w1915) );
	AND U1600 ( .A(w1914), .B(w1915), .Z(w1916) );
	AND U1601 ( .A(w1890), .B(w1821), .Z(w1917) );
	XOR U1602 ( .A(w1917), .B(w1916), .Z(w1918) );
	AND U1603 ( .A(w1892), .B(w1820), .Z(w1919) );
	XOR U1604 ( .A(w1919), .B(w1916), .Z(w1920) );
	XOR U1605 ( .A(w1913), .B(w1906), .Z(w1921) );
	XOR U1606 ( .A(w1911), .B(w1905), .Z(w1922) );
	XOR U1607 ( .A(w1920), .B(w1906), .Z(w1923) );
	XOR U1608 ( .A(w1918), .B(w1905), .Z(w1924) );
	XOR U1609 ( .A(w1885), .B(w1892), .Z(w1927) );
	XOR U1610 ( .A(w1883), .B(w1890), .Z(w1928) );
	XOR U1611 ( .A(w1818), .B(w1816), .Z(w1929) );
	XOR U1612 ( .A(w1819), .B(w1817), .Z(w1930) );
	XOR U1613 ( .A(w1928), .B(w1927), .Z(w1931) );
	XOR U1614 ( .A(w1930), .B(w1929), .Z(w1932) );
	AND U1615 ( .A(w1931), .B(w1932), .Z(w1933) );
	AND U1616 ( .A(w1928), .B(w1930), .Z(w1934) );
	XOR U1617 ( .A(w1934), .B(w1933), .Z(w1935) );
	AND U1618 ( .A(w1927), .B(w1929), .Z(w1936) );
	XOR U1619 ( .A(w1936), .B(w1933), .Z(w1937) );
	XOR U1620 ( .A(w1937), .B(w1935), .Z(w1938) );
	XOR U1621 ( .A(w1883), .B(w1885), .Z(w1939) );
	XOR U1622 ( .A(w1819), .B(w1818), .Z(w1940) );
	AND U1623 ( .A(w1939), .B(w1940), .Z(w1941) );
	AND U1624 ( .A(w1883), .B(w1819), .Z(w1942) );
	XOR U1625 ( .A(w1942), .B(w1941), .Z(w1943) );
	AND U1626 ( .A(w1885), .B(w1818), .Z(w1944) );
	XOR U1627 ( .A(w1944), .B(w1941), .Z(w1945) );
	XOR U1628 ( .A(w1890), .B(w1892), .Z(w1946) );
	XOR U1629 ( .A(w1817), .B(w1816), .Z(w1947) );
	AND U1630 ( .A(w1946), .B(w1947), .Z(w1948) );
	AND U1631 ( .A(w1890), .B(w1817), .Z(w1949) );
	XOR U1632 ( .A(w1949), .B(w1948), .Z(w1950) );
	AND U1633 ( .A(w1892), .B(w1816), .Z(w1951) );
	XOR U1634 ( .A(w1951), .B(w1948), .Z(w1952) );
	XOR U1635 ( .A(w1945), .B(w1938), .Z(w1953) );
	XOR U1636 ( .A(w1943), .B(w1937), .Z(w1954) );
	XOR U1637 ( .A(w1952), .B(w1938), .Z(w1955) );
	XOR U1638 ( .A(w1950), .B(w1937), .Z(w1956) );
	XOR U1639 ( .A(w1959), .B(w1955), .Z(w1965) );
	XOR U1640 ( .A(w1960), .B(w1955), .Z(w1966) );
	XOR U1641 ( .A(w1964), .B(w1955), .Z(w1967) );
	XOR U1642 ( .A(w1957), .B(w1956), .Z(w1968) );
	XOR U1643 ( .A(w1966), .B(w1956), .Z(w1969) );
	XOR U1644 ( .A(w1961), .B(w1956), .Z(w1970) );
	XOR U1645 ( .A(w1962), .B(w1956), .Z(w1971) );
	XOR U1646 ( .A(w1963), .B(w1956), .Z(w1972) );
	XOR U1647 ( .A(w1968), .B(w1953), .Z(w1973) );
	XOR U1648 ( .A(w1965), .B(w1953), .Z(w1974) );
	XOR U1649 ( .A(w1973), .B(w1954), .Z(w1975) );
	XOR U1650 ( .A(w1958), .B(w1954), .Z(w1976) );
	XOR U1651 ( .A(w1969), .B(w1954), .Z(w1977) );
	XOR U1652 ( .A(w1971), .B(w1954), .Z(w1978) );
	XOR U1653 ( .A(w1972), .B(w1954), .Z(w1979) );
	XOR U1654 ( .A(w1967), .B(w1954), .Z(w1980) );
	XOR U1655 ( .A(w1976), .B(w1923), .Z(w1981) );
	XOR U1656 ( .A(w1970), .B(w1923), .Z(w1982) );
	XOR U1657 ( .A(w1974), .B(w1924), .Z(w1983) );
	XOR U1658 ( .A(w1975), .B(w1921), .Z(w1984) );
	XOR U1659 ( .A(w1982), .B(w1921), .Z(w1985) );
	XOR U1660 ( .A(w1979), .B(w1921), .Z(w1986) );
	XOR U1661 ( .A(w1984), .B(w1922), .Z(w1987) );
	XOR U1662 ( .A(w1981), .B(w1922), .Z(w1988) );
	XOR U1663 ( .A(w1985), .B(w1922), .Z(w1989) );
	XOR U1664 ( .A(w1986), .B(w1922), .Z(w1990) );
	XOR U1665 ( .A(w1994), .B(w72), .Z(w1999) );
	XOR U1666 ( .A(w1995), .B(w72), .Z(w2000) );
	XOR U1667 ( .A(w1998), .B(w72), .Z(w2001) );
	XOR U1668 ( .A(w1991), .B(w73), .Z(w2002) );
	XOR U1669 ( .A(w1992), .B(w73), .Z(w2003) );
	XOR U1670 ( .A(w2000), .B(w73), .Z(w2004) );
	XOR U1671 ( .A(w1996), .B(w73), .Z(w2005) );
	XOR U1672 ( .A(w1997), .B(w73), .Z(w2006) );
	XOR U1673 ( .A(w2001), .B(w73), .Z(w2007) );
	XOR U1674 ( .A(w2003), .B(w74), .Z(w2008) );
	XOR U1675 ( .A(w2004), .B(w74), .Z(w2009) );
	XOR U1676 ( .A(w2005), .B(w74), .Z(w2010) );
	XOR U1677 ( .A(w2006), .B(w74), .Z(w2011) );
	XOR U1678 ( .A(w2007), .B(w74), .Z(w2012) );
	XOR U1679 ( .A(w1999), .B(w75), .Z(w2013) );
	XOR U1680 ( .A(w2011), .B(w75), .Z(w2014) );
	XOR U1681 ( .A(w2002), .B(w76), .Z(w2015) );
	XOR U1682 ( .A(w2013), .B(w76), .Z(w2016) );
	XOR U1683 ( .A(w2015), .B(w77), .Z(w2017) );
	XOR U1684 ( .A(w2012), .B(w77), .Z(w2018) );
	XOR U1685 ( .A(w2017), .B(w78), .Z(w2019) );
	XOR U1686 ( .A(w2016), .B(w78), .Z(w2020) );
	XOR U1687 ( .A(w2010), .B(w78), .Z(w2021) );
	XOR U1688 ( .A(w2018), .B(w78), .Z(w2022) );
	XOR U1689 ( .A(w2019), .B(w79), .Z(w2023) );
	XOR U1690 ( .A(w2008), .B(w79), .Z(w2024) );
	XOR U1691 ( .A(w1993), .B(w79), .Z(w2025) );
	XOR U1692 ( .A(w2020), .B(w79), .Z(w2026) );
	XOR U1693 ( .A(w2009), .B(w79), .Z(w2027) );
	XOR U1694 ( .A(w2021), .B(w79), .Z(w2028) );
	XOR U1695 ( .A(w2014), .B(w79), .Z(w2029) );
	XOR U1696 ( .A(w2022), .B(w79), .Z(w2030) );
	XOR U1697 ( .A(w2023), .B(w2027), .Z(w2031) );
	XOR U1698 ( .A(w2024), .B(w2028), .Z(w2032) );
	XOR U1699 ( .A(w2025), .B(w2029), .Z(w2033) );
	XOR U1700 ( .A(w2026), .B(w2030), .Z(w2034) );
	XOR U1701 ( .A(w2033), .B(w2031), .Z(w2035) );
	XOR U1702 ( .A(w2034), .B(w2032), .Z(w2036) );
	XOR U1703 ( .A(w2032), .B(w2031), .Z(w2037) );
	XOR U1704 ( .A(w2025), .B(w2023), .Z(w2040) );
	XOR U1705 ( .A(w2026), .B(w2024), .Z(w2041) );
	XOR U1706 ( .A(w2029), .B(w2027), .Z(w2042) );
	XOR U1707 ( .A(w2030), .B(w2028), .Z(w2043) );
	XOR U1708 ( .A(w2041), .B(w2040), .Z(w2044) );
	XOR U1709 ( .A(w2043), .B(w2042), .Z(w2045) );
	AND U1710 ( .A(w2044), .B(w2045), .Z(w2046) );
	AND U1711 ( .A(w2041), .B(w2043), .Z(w2047) );
	XOR U1712 ( .A(w2047), .B(w2046), .Z(w2048) );
	AND U1713 ( .A(w2040), .B(w2042), .Z(w2049) );
	XOR U1714 ( .A(w2049), .B(w2046), .Z(w2050) );
	XOR U1715 ( .A(w2050), .B(w2048), .Z(w2051) );
	XOR U1716 ( .A(w2026), .B(w2025), .Z(w2052) );
	XOR U1717 ( .A(w2030), .B(w2029), .Z(w2053) );
	AND U1718 ( .A(w2052), .B(w2053), .Z(w2054) );
	AND U1719 ( .A(w2026), .B(w2030), .Z(w2055) );
	XOR U1720 ( .A(w2055), .B(w2054), .Z(w2056) );
	AND U1721 ( .A(w2025), .B(w2029), .Z(w2057) );
	XOR U1722 ( .A(w2057), .B(w2054), .Z(w2058) );
	XOR U1723 ( .A(w2024), .B(w2023), .Z(w2059) );
	XOR U1724 ( .A(w2028), .B(w2027), .Z(w2060) );
	AND U1725 ( .A(w2059), .B(w2060), .Z(w2061) );
	AND U1726 ( .A(w2024), .B(w2028), .Z(w2062) );
	XOR U1727 ( .A(w2062), .B(w2061), .Z(w2063) );
	AND U1728 ( .A(w2023), .B(w2027), .Z(w2064) );
	XOR U1729 ( .A(w2064), .B(w2061), .Z(w2065) );
	XOR U1730 ( .A(w2058), .B(w2051), .Z(w2066) );
	XOR U1731 ( .A(w2056), .B(w2050), .Z(w2067) );
	XOR U1732 ( .A(w2065), .B(w2051), .Z(w2068) );
	XOR U1733 ( .A(w2063), .B(w2050), .Z(w2069) );
	XOR U1734 ( .A(w2031), .B(w2068), .Z(w2070) );
	XOR U1735 ( .A(w2037), .B(w2069), .Z(w2071) );
	XOR U1736 ( .A(w2036), .B(w2066), .Z(w2072) );
	XOR U1737 ( .A(w2035), .B(w2067), .Z(w2073) );
	XOR U1738 ( .A(w2072), .B(w2070), .Z(w2074) );
	XOR U1739 ( .A(w2073), .B(w2071), .Z(w2075) );
	XOR U1740 ( .A(w2075), .B(w2074), .Z(w2076) );
	XOR U1741 ( .A(w2073), .B(w2072), .Z(w2077) );
	XOR U1742 ( .A(w2071), .B(w2070), .Z(w2078) );
	AND U1743 ( .A(w2077), .B(w2078), .Z(w2079) );
	AND U1744 ( .A(w2073), .B(w2071), .Z(w2080) );
	XOR U1745 ( .A(w2080), .B(w2079), .Z(w2081) );
	AND U1746 ( .A(w2072), .B(w2070), .Z(w2082) );
	XOR U1747 ( .A(w2082), .B(w2079), .Z(w2083) );
	XOR U1748 ( .A(w2076), .B(w2083), .Z(w2084) );
	XOR U1749 ( .A(w2075), .B(w2081), .Z(w2085) );
	XOR U1750 ( .A(w2084), .B(w2085), .Z(w2086) );
	XOR U1751 ( .A(w2071), .B(w2070), .Z(w2087) );
	AND U1752 ( .A(w2086), .B(w2087), .Z(w2088) );
	AND U1753 ( .A(w2084), .B(w2071), .Z(w2089) );
	XOR U1754 ( .A(w2089), .B(w2088), .Z(w2090) );
	AND U1755 ( .A(w2085), .B(w2070), .Z(w2091) );
	XOR U1756 ( .A(w2091), .B(w2088), .Z(w2092) );
	XOR U1757 ( .A(w2084), .B(w2085), .Z(w2093) );
	XOR U1758 ( .A(w2073), .B(w2072), .Z(w2094) );
	AND U1759 ( .A(w2093), .B(w2094), .Z(w2095) );
	AND U1760 ( .A(w2084), .B(w2073), .Z(w2096) );
	XOR U1761 ( .A(w2096), .B(w2095), .Z(w2097) );
	AND U1762 ( .A(w2085), .B(w2072), .Z(w2098) );
	XOR U1763 ( .A(w2098), .B(w2095), .Z(w2099) );
	XOR U1764 ( .A(w2092), .B(w2099), .Z(w2102) );
	XOR U1765 ( .A(w2090), .B(w2097), .Z(w2103) );
	XOR U1766 ( .A(w2029), .B(w2027), .Z(w2104) );
	XOR U1767 ( .A(w2030), .B(w2028), .Z(w2105) );
	XOR U1768 ( .A(w2103), .B(w2102), .Z(w2106) );
	XOR U1769 ( .A(w2105), .B(w2104), .Z(w2107) );
	AND U1770 ( .A(w2106), .B(w2107), .Z(w2108) );
	AND U1771 ( .A(w2103), .B(w2105), .Z(w2109) );
	XOR U1772 ( .A(w2109), .B(w2108), .Z(w2110) );
	AND U1773 ( .A(w2102), .B(w2104), .Z(w2111) );
	XOR U1774 ( .A(w2111), .B(w2108), .Z(w2112) );
	XOR U1775 ( .A(w2112), .B(w2110), .Z(w2113) );
	XOR U1776 ( .A(w2090), .B(w2092), .Z(w2114) );
	XOR U1777 ( .A(w2030), .B(w2029), .Z(w2115) );
	AND U1778 ( .A(w2114), .B(w2115), .Z(w2116) );
	AND U1779 ( .A(w2090), .B(w2030), .Z(w2117) );
	XOR U1780 ( .A(w2117), .B(w2116), .Z(w2118) );
	AND U1781 ( .A(w2092), .B(w2029), .Z(w2119) );
	XOR U1782 ( .A(w2119), .B(w2116), .Z(w2120) );
	XOR U1783 ( .A(w2097), .B(w2099), .Z(w2121) );
	XOR U1784 ( .A(w2028), .B(w2027), .Z(w2122) );
	AND U1785 ( .A(w2121), .B(w2122), .Z(w2123) );
	AND U1786 ( .A(w2097), .B(w2028), .Z(w2124) );
	XOR U1787 ( .A(w2124), .B(w2123), .Z(w2125) );
	AND U1788 ( .A(w2099), .B(w2027), .Z(w2126) );
	XOR U1789 ( .A(w2126), .B(w2123), .Z(w2127) );
	XOR U1790 ( .A(w2120), .B(w2113), .Z(w2128) );
	XOR U1791 ( .A(w2118), .B(w2112), .Z(w2129) );
	XOR U1792 ( .A(w2127), .B(w2113), .Z(w2130) );
	XOR U1793 ( .A(w2125), .B(w2112), .Z(w2131) );
	XOR U1794 ( .A(w2092), .B(w2099), .Z(w2134) );
	XOR U1795 ( .A(w2090), .B(w2097), .Z(w2135) );
	XOR U1796 ( .A(w2025), .B(w2023), .Z(w2136) );
	XOR U1797 ( .A(w2026), .B(w2024), .Z(w2137) );
	XOR U1798 ( .A(w2135), .B(w2134), .Z(w2138) );
	XOR U1799 ( .A(w2137), .B(w2136), .Z(w2139) );
	AND U1800 ( .A(w2138), .B(w2139), .Z(w2140) );
	AND U1801 ( .A(w2135), .B(w2137), .Z(w2141) );
	XOR U1802 ( .A(w2141), .B(w2140), .Z(w2142) );
	AND U1803 ( .A(w2134), .B(w2136), .Z(w2143) );
	XOR U1804 ( .A(w2143), .B(w2140), .Z(w2144) );
	XOR U1805 ( .A(w2144), .B(w2142), .Z(w2145) );
	XOR U1806 ( .A(w2090), .B(w2092), .Z(w2146) );
	XOR U1807 ( .A(w2026), .B(w2025), .Z(w2147) );
	AND U1808 ( .A(w2146), .B(w2147), .Z(w2148) );
	AND U1809 ( .A(w2090), .B(w2026), .Z(w2149) );
	XOR U1810 ( .A(w2149), .B(w2148), .Z(w2150) );
	AND U1811 ( .A(w2092), .B(w2025), .Z(w2151) );
	XOR U1812 ( .A(w2151), .B(w2148), .Z(w2152) );
	XOR U1813 ( .A(w2097), .B(w2099), .Z(w2153) );
	XOR U1814 ( .A(w2024), .B(w2023), .Z(w2154) );
	AND U1815 ( .A(w2153), .B(w2154), .Z(w2155) );
	AND U1816 ( .A(w2097), .B(w2024), .Z(w2156) );
	XOR U1817 ( .A(w2156), .B(w2155), .Z(w2157) );
	AND U1818 ( .A(w2099), .B(w2023), .Z(w2158) );
	XOR U1819 ( .A(w2158), .B(w2155), .Z(w2159) );
	XOR U1820 ( .A(w2152), .B(w2145), .Z(w2160) );
	XOR U1821 ( .A(w2150), .B(w2144), .Z(w2161) );
	XOR U1822 ( .A(w2159), .B(w2145), .Z(w2162) );
	XOR U1823 ( .A(w2157), .B(w2144), .Z(w2163) );
	XOR U1824 ( .A(w2166), .B(w2162), .Z(w2172) );
	XOR U1825 ( .A(w2167), .B(w2162), .Z(w2173) );
	XOR U1826 ( .A(w2171), .B(w2162), .Z(w2174) );
	XOR U1827 ( .A(w2164), .B(w2163), .Z(w2175) );
	XOR U1828 ( .A(w2173), .B(w2163), .Z(w2176) );
	XOR U1829 ( .A(w2168), .B(w2163), .Z(w2177) );
	XOR U1830 ( .A(w2169), .B(w2163), .Z(w2178) );
	XOR U1831 ( .A(w2170), .B(w2163), .Z(w2179) );
	XOR U1832 ( .A(w2175), .B(w2160), .Z(w2180) );
	XOR U1833 ( .A(w2172), .B(w2160), .Z(w2181) );
	XOR U1834 ( .A(w2180), .B(w2161), .Z(w2182) );
	XOR U1835 ( .A(w2165), .B(w2161), .Z(w2183) );
	XOR U1836 ( .A(w2176), .B(w2161), .Z(w2184) );
	XOR U1837 ( .A(w2178), .B(w2161), .Z(w2185) );
	XOR U1838 ( .A(w2179), .B(w2161), .Z(w2186) );
	XOR U1839 ( .A(w2174), .B(w2161), .Z(w2187) );
	XOR U1840 ( .A(w2183), .B(w2130), .Z(w2188) );
	XOR U1841 ( .A(w2177), .B(w2130), .Z(w2189) );
	XOR U1842 ( .A(w2181), .B(w2131), .Z(w2190) );
	XOR U1843 ( .A(w2182), .B(w2128), .Z(w2191) );
	XOR U1844 ( .A(w2189), .B(w2128), .Z(w2192) );
	XOR U1845 ( .A(w2186), .B(w2128), .Z(w2193) );
	XOR U1846 ( .A(w2191), .B(w2129), .Z(w2194) );
	XOR U1847 ( .A(w2188), .B(w2129), .Z(w2195) );
	XOR U1848 ( .A(w2192), .B(w2129), .Z(w2196) );
	XOR U1849 ( .A(w2193), .B(w2129), .Z(w2197) );
	XOR U1850 ( .A(w2201), .B(w80), .Z(w2206) );
	XOR U1851 ( .A(w2202), .B(w80), .Z(w2207) );
	XOR U1852 ( .A(w2205), .B(w80), .Z(w2208) );
	XOR U1853 ( .A(w2198), .B(w81), .Z(w2209) );
	XOR U1854 ( .A(w2199), .B(w81), .Z(w2210) );
	XOR U1855 ( .A(w2207), .B(w81), .Z(w2211) );
	XOR U1856 ( .A(w2203), .B(w81), .Z(w2212) );
	XOR U1857 ( .A(w2204), .B(w81), .Z(w2213) );
	XOR U1858 ( .A(w2208), .B(w81), .Z(w2214) );
	XOR U1859 ( .A(w2210), .B(w82), .Z(w2215) );
	XOR U1860 ( .A(w2211), .B(w82), .Z(w2216) );
	XOR U1861 ( .A(w2212), .B(w82), .Z(w2217) );
	XOR U1862 ( .A(w2213), .B(w82), .Z(w2218) );
	XOR U1863 ( .A(w2214), .B(w82), .Z(w2219) );
	XOR U1864 ( .A(w2206), .B(w83), .Z(w2220) );
	XOR U1865 ( .A(w2218), .B(w83), .Z(w2221) );
	XOR U1866 ( .A(w2209), .B(w84), .Z(w2222) );
	XOR U1867 ( .A(w2220), .B(w84), .Z(w2223) );
	XOR U1868 ( .A(w2222), .B(w85), .Z(w2224) );
	XOR U1869 ( .A(w2219), .B(w85), .Z(w2225) );
	XOR U1870 ( .A(w2224), .B(w86), .Z(w2226) );
	XOR U1871 ( .A(w2223), .B(w86), .Z(w2227) );
	XOR U1872 ( .A(w2217), .B(w86), .Z(w2228) );
	XOR U1873 ( .A(w2225), .B(w86), .Z(w2229) );
	XOR U1874 ( .A(w2226), .B(w87), .Z(w2230) );
	XOR U1875 ( .A(w2215), .B(w87), .Z(w2231) );
	XOR U1876 ( .A(w2200), .B(w87), .Z(w2232) );
	XOR U1877 ( .A(w2227), .B(w87), .Z(w2233) );
	XOR U1878 ( .A(w2216), .B(w87), .Z(w2234) );
	XOR U1879 ( .A(w2228), .B(w87), .Z(w2235) );
	XOR U1880 ( .A(w2221), .B(w87), .Z(w2236) );
	XOR U1881 ( .A(w2229), .B(w87), .Z(w2237) );
	XOR U1882 ( .A(w2230), .B(w2234), .Z(w2238) );
	XOR U1883 ( .A(w2231), .B(w2235), .Z(w2239) );
	XOR U1884 ( .A(w2232), .B(w2236), .Z(w2240) );
	XOR U1885 ( .A(w2233), .B(w2237), .Z(w2241) );
	XOR U1886 ( .A(w2240), .B(w2238), .Z(w2242) );
	XOR U1887 ( .A(w2241), .B(w2239), .Z(w2243) );
	XOR U1888 ( .A(w2239), .B(w2238), .Z(w2244) );
	XOR U1889 ( .A(w2232), .B(w2230), .Z(w2247) );
	XOR U1890 ( .A(w2233), .B(w2231), .Z(w2248) );
	XOR U1891 ( .A(w2236), .B(w2234), .Z(w2249) );
	XOR U1892 ( .A(w2237), .B(w2235), .Z(w2250) );
	XOR U1893 ( .A(w2248), .B(w2247), .Z(w2251) );
	XOR U1894 ( .A(w2250), .B(w2249), .Z(w2252) );
	AND U1895 ( .A(w2251), .B(w2252), .Z(w2253) );
	AND U1896 ( .A(w2248), .B(w2250), .Z(w2254) );
	XOR U1897 ( .A(w2254), .B(w2253), .Z(w2255) );
	AND U1898 ( .A(w2247), .B(w2249), .Z(w2256) );
	XOR U1899 ( .A(w2256), .B(w2253), .Z(w2257) );
	XOR U1900 ( .A(w2257), .B(w2255), .Z(w2258) );
	XOR U1901 ( .A(w2233), .B(w2232), .Z(w2259) );
	XOR U1902 ( .A(w2237), .B(w2236), .Z(w2260) );
	AND U1903 ( .A(w2259), .B(w2260), .Z(w2261) );
	AND U1904 ( .A(w2233), .B(w2237), .Z(w2262) );
	XOR U1905 ( .A(w2262), .B(w2261), .Z(w2263) );
	AND U1906 ( .A(w2232), .B(w2236), .Z(w2264) );
	XOR U1907 ( .A(w2264), .B(w2261), .Z(w2265) );
	XOR U1908 ( .A(w2231), .B(w2230), .Z(w2266) );
	XOR U1909 ( .A(w2235), .B(w2234), .Z(w2267) );
	AND U1910 ( .A(w2266), .B(w2267), .Z(w2268) );
	AND U1911 ( .A(w2231), .B(w2235), .Z(w2269) );
	XOR U1912 ( .A(w2269), .B(w2268), .Z(w2270) );
	AND U1913 ( .A(w2230), .B(w2234), .Z(w2271) );
	XOR U1914 ( .A(w2271), .B(w2268), .Z(w2272) );
	XOR U1915 ( .A(w2265), .B(w2258), .Z(w2273) );
	XOR U1916 ( .A(w2263), .B(w2257), .Z(w2274) );
	XOR U1917 ( .A(w2272), .B(w2258), .Z(w2275) );
	XOR U1918 ( .A(w2270), .B(w2257), .Z(w2276) );
	XOR U1919 ( .A(w2238), .B(w2275), .Z(w2277) );
	XOR U1920 ( .A(w2244), .B(w2276), .Z(w2278) );
	XOR U1921 ( .A(w2243), .B(w2273), .Z(w2279) );
	XOR U1922 ( .A(w2242), .B(w2274), .Z(w2280) );
	XOR U1923 ( .A(w2279), .B(w2277), .Z(w2281) );
	XOR U1924 ( .A(w2280), .B(w2278), .Z(w2282) );
	XOR U1925 ( .A(w2282), .B(w2281), .Z(w2283) );
	XOR U1926 ( .A(w2280), .B(w2279), .Z(w2284) );
	XOR U1927 ( .A(w2278), .B(w2277), .Z(w2285) );
	AND U1928 ( .A(w2284), .B(w2285), .Z(w2286) );
	AND U1929 ( .A(w2280), .B(w2278), .Z(w2287) );
	XOR U1930 ( .A(w2287), .B(w2286), .Z(w2288) );
	AND U1931 ( .A(w2279), .B(w2277), .Z(w2289) );
	XOR U1932 ( .A(w2289), .B(w2286), .Z(w2290) );
	XOR U1933 ( .A(w2283), .B(w2290), .Z(w2291) );
	XOR U1934 ( .A(w2282), .B(w2288), .Z(w2292) );
	XOR U1935 ( .A(w2291), .B(w2292), .Z(w2293) );
	XOR U1936 ( .A(w2278), .B(w2277), .Z(w2294) );
	AND U1937 ( .A(w2293), .B(w2294), .Z(w2295) );
	AND U1938 ( .A(w2291), .B(w2278), .Z(w2296) );
	XOR U1939 ( .A(w2296), .B(w2295), .Z(w2297) );
	AND U1940 ( .A(w2292), .B(w2277), .Z(w2298) );
	XOR U1941 ( .A(w2298), .B(w2295), .Z(w2299) );
	XOR U1942 ( .A(w2291), .B(w2292), .Z(w2300) );
	XOR U1943 ( .A(w2280), .B(w2279), .Z(w2301) );
	AND U1944 ( .A(w2300), .B(w2301), .Z(w2302) );
	AND U1945 ( .A(w2291), .B(w2280), .Z(w2303) );
	XOR U1946 ( .A(w2303), .B(w2302), .Z(w2304) );
	AND U1947 ( .A(w2292), .B(w2279), .Z(w2305) );
	XOR U1948 ( .A(w2305), .B(w2302), .Z(w2306) );
	XOR U1949 ( .A(w2299), .B(w2306), .Z(w2309) );
	XOR U1950 ( .A(w2297), .B(w2304), .Z(w2310) );
	XOR U1951 ( .A(w2236), .B(w2234), .Z(w2311) );
	XOR U1952 ( .A(w2237), .B(w2235), .Z(w2312) );
	XOR U1953 ( .A(w2310), .B(w2309), .Z(w2313) );
	XOR U1954 ( .A(w2312), .B(w2311), .Z(w2314) );
	AND U1955 ( .A(w2313), .B(w2314), .Z(w2315) );
	AND U1956 ( .A(w2310), .B(w2312), .Z(w2316) );
	XOR U1957 ( .A(w2316), .B(w2315), .Z(w2317) );
	AND U1958 ( .A(w2309), .B(w2311), .Z(w2318) );
	XOR U1959 ( .A(w2318), .B(w2315), .Z(w2319) );
	XOR U1960 ( .A(w2319), .B(w2317), .Z(w2320) );
	XOR U1961 ( .A(w2297), .B(w2299), .Z(w2321) );
	XOR U1962 ( .A(w2237), .B(w2236), .Z(w2322) );
	AND U1963 ( .A(w2321), .B(w2322), .Z(w2323) );
	AND U1964 ( .A(w2297), .B(w2237), .Z(w2324) );
	XOR U1965 ( .A(w2324), .B(w2323), .Z(w2325) );
	AND U1966 ( .A(w2299), .B(w2236), .Z(w2326) );
	XOR U1967 ( .A(w2326), .B(w2323), .Z(w2327) );
	XOR U1968 ( .A(w2304), .B(w2306), .Z(w2328) );
	XOR U1969 ( .A(w2235), .B(w2234), .Z(w2329) );
	AND U1970 ( .A(w2328), .B(w2329), .Z(w2330) );
	AND U1971 ( .A(w2304), .B(w2235), .Z(w2331) );
	XOR U1972 ( .A(w2331), .B(w2330), .Z(w2332) );
	AND U1973 ( .A(w2306), .B(w2234), .Z(w2333) );
	XOR U1974 ( .A(w2333), .B(w2330), .Z(w2334) );
	XOR U1975 ( .A(w2327), .B(w2320), .Z(w2335) );
	XOR U1976 ( .A(w2325), .B(w2319), .Z(w2336) );
	XOR U1977 ( .A(w2334), .B(w2320), .Z(w2337) );
	XOR U1978 ( .A(w2332), .B(w2319), .Z(w2338) );
	XOR U1979 ( .A(w2299), .B(w2306), .Z(w2341) );
	XOR U1980 ( .A(w2297), .B(w2304), .Z(w2342) );
	XOR U1981 ( .A(w2232), .B(w2230), .Z(w2343) );
	XOR U1982 ( .A(w2233), .B(w2231), .Z(w2344) );
	XOR U1983 ( .A(w2342), .B(w2341), .Z(w2345) );
	XOR U1984 ( .A(w2344), .B(w2343), .Z(w2346) );
	AND U1985 ( .A(w2345), .B(w2346), .Z(w2347) );
	AND U1986 ( .A(w2342), .B(w2344), .Z(w2348) );
	XOR U1987 ( .A(w2348), .B(w2347), .Z(w2349) );
	AND U1988 ( .A(w2341), .B(w2343), .Z(w2350) );
	XOR U1989 ( .A(w2350), .B(w2347), .Z(w2351) );
	XOR U1990 ( .A(w2351), .B(w2349), .Z(w2352) );
	XOR U1991 ( .A(w2297), .B(w2299), .Z(w2353) );
	XOR U1992 ( .A(w2233), .B(w2232), .Z(w2354) );
	AND U1993 ( .A(w2353), .B(w2354), .Z(w2355) );
	AND U1994 ( .A(w2297), .B(w2233), .Z(w2356) );
	XOR U1995 ( .A(w2356), .B(w2355), .Z(w2357) );
	AND U1996 ( .A(w2299), .B(w2232), .Z(w2358) );
	XOR U1997 ( .A(w2358), .B(w2355), .Z(w2359) );
	XOR U1998 ( .A(w2304), .B(w2306), .Z(w2360) );
	XOR U1999 ( .A(w2231), .B(w2230), .Z(w2361) );
	AND U2000 ( .A(w2360), .B(w2361), .Z(w2362) );
	AND U2001 ( .A(w2304), .B(w2231), .Z(w2363) );
	XOR U2002 ( .A(w2363), .B(w2362), .Z(w2364) );
	AND U2003 ( .A(w2306), .B(w2230), .Z(w2365) );
	XOR U2004 ( .A(w2365), .B(w2362), .Z(w2366) );
	XOR U2005 ( .A(w2359), .B(w2352), .Z(w2367) );
	XOR U2006 ( .A(w2357), .B(w2351), .Z(w2368) );
	XOR U2007 ( .A(w2366), .B(w2352), .Z(w2369) );
	XOR U2008 ( .A(w2364), .B(w2351), .Z(w2370) );
	XOR U2009 ( .A(w2373), .B(w2369), .Z(w2379) );
	XOR U2010 ( .A(w2374), .B(w2369), .Z(w2380) );
	XOR U2011 ( .A(w2378), .B(w2369), .Z(w2381) );
	XOR U2012 ( .A(w2371), .B(w2370), .Z(w2382) );
	XOR U2013 ( .A(w2380), .B(w2370), .Z(w2383) );
	XOR U2014 ( .A(w2375), .B(w2370), .Z(w2384) );
	XOR U2015 ( .A(w2376), .B(w2370), .Z(w2385) );
	XOR U2016 ( .A(w2377), .B(w2370), .Z(w2386) );
	XOR U2017 ( .A(w2382), .B(w2367), .Z(w2387) );
	XOR U2018 ( .A(w2379), .B(w2367), .Z(w2388) );
	XOR U2019 ( .A(w2387), .B(w2368), .Z(w2389) );
	XOR U2020 ( .A(w2372), .B(w2368), .Z(w2390) );
	XOR U2021 ( .A(w2383), .B(w2368), .Z(w2391) );
	XOR U2022 ( .A(w2385), .B(w2368), .Z(w2392) );
	XOR U2023 ( .A(w2386), .B(w2368), .Z(w2393) );
	XOR U2024 ( .A(w2381), .B(w2368), .Z(w2394) );
	XOR U2025 ( .A(w2390), .B(w2337), .Z(w2395) );
	XOR U2026 ( .A(w2384), .B(w2337), .Z(w2396) );
	XOR U2027 ( .A(w2388), .B(w2338), .Z(w2397) );
	XOR U2028 ( .A(w2389), .B(w2335), .Z(w2398) );
	XOR U2029 ( .A(w2396), .B(w2335), .Z(w2399) );
	XOR U2030 ( .A(w2393), .B(w2335), .Z(w2400) );
	XOR U2031 ( .A(w2398), .B(w2336), .Z(w2401) );
	XOR U2032 ( .A(w2395), .B(w2336), .Z(w2402) );
	XOR U2033 ( .A(w2399), .B(w2336), .Z(w2403) );
	XOR U2034 ( .A(w2400), .B(w2336), .Z(w2404) );
	XOR U2035 ( .A(w2408), .B(w88), .Z(w2413) );
	XOR U2036 ( .A(w2409), .B(w88), .Z(w2414) );
	XOR U2037 ( .A(w2412), .B(w88), .Z(w2415) );
	XOR U2038 ( .A(w2405), .B(w89), .Z(w2416) );
	XOR U2039 ( .A(w2406), .B(w89), .Z(w2417) );
	XOR U2040 ( .A(w2414), .B(w89), .Z(w2418) );
	XOR U2041 ( .A(w2410), .B(w89), .Z(w2419) );
	XOR U2042 ( .A(w2411), .B(w89), .Z(w2420) );
	XOR U2043 ( .A(w2415), .B(w89), .Z(w2421) );
	XOR U2044 ( .A(w2417), .B(w90), .Z(w2422) );
	XOR U2045 ( .A(w2418), .B(w90), .Z(w2423) );
	XOR U2046 ( .A(w2419), .B(w90), .Z(w2424) );
	XOR U2047 ( .A(w2420), .B(w90), .Z(w2425) );
	XOR U2048 ( .A(w2421), .B(w90), .Z(w2426) );
	XOR U2049 ( .A(w2413), .B(w91), .Z(w2427) );
	XOR U2050 ( .A(w2425), .B(w91), .Z(w2428) );
	XOR U2051 ( .A(w2416), .B(w92), .Z(w2429) );
	XOR U2052 ( .A(w2427), .B(w92), .Z(w2430) );
	XOR U2053 ( .A(w2429), .B(w93), .Z(w2431) );
	XOR U2054 ( .A(w2426), .B(w93), .Z(w2432) );
	XOR U2055 ( .A(w2431), .B(w94), .Z(w2433) );
	XOR U2056 ( .A(w2430), .B(w94), .Z(w2434) );
	XOR U2057 ( .A(w2424), .B(w94), .Z(w2435) );
	XOR U2058 ( .A(w2432), .B(w94), .Z(w2436) );
	XOR U2059 ( .A(w2433), .B(w95), .Z(w2437) );
	XOR U2060 ( .A(w2422), .B(w95), .Z(w2438) );
	XOR U2061 ( .A(w2407), .B(w95), .Z(w2439) );
	XOR U2062 ( .A(w2434), .B(w95), .Z(w2440) );
	XOR U2063 ( .A(w2423), .B(w95), .Z(w2441) );
	XOR U2064 ( .A(w2435), .B(w95), .Z(w2442) );
	XOR U2065 ( .A(w2428), .B(w95), .Z(w2443) );
	XOR U2066 ( .A(w2436), .B(w95), .Z(w2444) );
	XOR U2067 ( .A(w2437), .B(w2441), .Z(w2445) );
	XOR U2068 ( .A(w2438), .B(w2442), .Z(w2446) );
	XOR U2069 ( .A(w2439), .B(w2443), .Z(w2447) );
	XOR U2070 ( .A(w2440), .B(w2444), .Z(w2448) );
	XOR U2071 ( .A(w2447), .B(w2445), .Z(w2449) );
	XOR U2072 ( .A(w2448), .B(w2446), .Z(w2450) );
	XOR U2073 ( .A(w2446), .B(w2445), .Z(w2451) );
	XOR U2074 ( .A(w2439), .B(w2437), .Z(w2454) );
	XOR U2075 ( .A(w2440), .B(w2438), .Z(w2455) );
	XOR U2076 ( .A(w2443), .B(w2441), .Z(w2456) );
	XOR U2077 ( .A(w2444), .B(w2442), .Z(w2457) );
	XOR U2078 ( .A(w2455), .B(w2454), .Z(w2458) );
	XOR U2079 ( .A(w2457), .B(w2456), .Z(w2459) );
	AND U2080 ( .A(w2458), .B(w2459), .Z(w2460) );
	AND U2081 ( .A(w2455), .B(w2457), .Z(w2461) );
	XOR U2082 ( .A(w2461), .B(w2460), .Z(w2462) );
	AND U2083 ( .A(w2454), .B(w2456), .Z(w2463) );
	XOR U2084 ( .A(w2463), .B(w2460), .Z(w2464) );
	XOR U2085 ( .A(w2464), .B(w2462), .Z(w2465) );
	XOR U2086 ( .A(w2440), .B(w2439), .Z(w2466) );
	XOR U2087 ( .A(w2444), .B(w2443), .Z(w2467) );
	AND U2088 ( .A(w2466), .B(w2467), .Z(w2468) );
	AND U2089 ( .A(w2440), .B(w2444), .Z(w2469) );
	XOR U2090 ( .A(w2469), .B(w2468), .Z(w2470) );
	AND U2091 ( .A(w2439), .B(w2443), .Z(w2471) );
	XOR U2092 ( .A(w2471), .B(w2468), .Z(w2472) );
	XOR U2093 ( .A(w2438), .B(w2437), .Z(w2473) );
	XOR U2094 ( .A(w2442), .B(w2441), .Z(w2474) );
	AND U2095 ( .A(w2473), .B(w2474), .Z(w2475) );
	AND U2096 ( .A(w2438), .B(w2442), .Z(w2476) );
	XOR U2097 ( .A(w2476), .B(w2475), .Z(w2477) );
	AND U2098 ( .A(w2437), .B(w2441), .Z(w2478) );
	XOR U2099 ( .A(w2478), .B(w2475), .Z(w2479) );
	XOR U2100 ( .A(w2472), .B(w2465), .Z(w2480) );
	XOR U2101 ( .A(w2470), .B(w2464), .Z(w2481) );
	XOR U2102 ( .A(w2479), .B(w2465), .Z(w2482) );
	XOR U2103 ( .A(w2477), .B(w2464), .Z(w2483) );
	XOR U2104 ( .A(w2445), .B(w2482), .Z(w2484) );
	XOR U2105 ( .A(w2451), .B(w2483), .Z(w2485) );
	XOR U2106 ( .A(w2450), .B(w2480), .Z(w2486) );
	XOR U2107 ( .A(w2449), .B(w2481), .Z(w2487) );
	XOR U2108 ( .A(w2486), .B(w2484), .Z(w2488) );
	XOR U2109 ( .A(w2487), .B(w2485), .Z(w2489) );
	XOR U2110 ( .A(w2489), .B(w2488), .Z(w2490) );
	XOR U2111 ( .A(w2487), .B(w2486), .Z(w2491) );
	XOR U2112 ( .A(w2485), .B(w2484), .Z(w2492) );
	AND U2113 ( .A(w2491), .B(w2492), .Z(w2493) );
	AND U2114 ( .A(w2487), .B(w2485), .Z(w2494) );
	XOR U2115 ( .A(w2494), .B(w2493), .Z(w2495) );
	AND U2116 ( .A(w2486), .B(w2484), .Z(w2496) );
	XOR U2117 ( .A(w2496), .B(w2493), .Z(w2497) );
	XOR U2118 ( .A(w2490), .B(w2497), .Z(w2498) );
	XOR U2119 ( .A(w2489), .B(w2495), .Z(w2499) );
	XOR U2120 ( .A(w2498), .B(w2499), .Z(w2500) );
	XOR U2121 ( .A(w2485), .B(w2484), .Z(w2501) );
	AND U2122 ( .A(w2500), .B(w2501), .Z(w2502) );
	AND U2123 ( .A(w2498), .B(w2485), .Z(w2503) );
	XOR U2124 ( .A(w2503), .B(w2502), .Z(w2504) );
	AND U2125 ( .A(w2499), .B(w2484), .Z(w2505) );
	XOR U2126 ( .A(w2505), .B(w2502), .Z(w2506) );
	XOR U2127 ( .A(w2498), .B(w2499), .Z(w2507) );
	XOR U2128 ( .A(w2487), .B(w2486), .Z(w2508) );
	AND U2129 ( .A(w2507), .B(w2508), .Z(w2509) );
	AND U2130 ( .A(w2498), .B(w2487), .Z(w2510) );
	XOR U2131 ( .A(w2510), .B(w2509), .Z(w2511) );
	AND U2132 ( .A(w2499), .B(w2486), .Z(w2512) );
	XOR U2133 ( .A(w2512), .B(w2509), .Z(w2513) );
	XOR U2134 ( .A(w2506), .B(w2513), .Z(w2516) );
	XOR U2135 ( .A(w2504), .B(w2511), .Z(w2517) );
	XOR U2136 ( .A(w2443), .B(w2441), .Z(w2518) );
	XOR U2137 ( .A(w2444), .B(w2442), .Z(w2519) );
	XOR U2138 ( .A(w2517), .B(w2516), .Z(w2520) );
	XOR U2139 ( .A(w2519), .B(w2518), .Z(w2521) );
	AND U2140 ( .A(w2520), .B(w2521), .Z(w2522) );
	AND U2141 ( .A(w2517), .B(w2519), .Z(w2523) );
	XOR U2142 ( .A(w2523), .B(w2522), .Z(w2524) );
	AND U2143 ( .A(w2516), .B(w2518), .Z(w2525) );
	XOR U2144 ( .A(w2525), .B(w2522), .Z(w2526) );
	XOR U2145 ( .A(w2526), .B(w2524), .Z(w2527) );
	XOR U2146 ( .A(w2504), .B(w2506), .Z(w2528) );
	XOR U2147 ( .A(w2444), .B(w2443), .Z(w2529) );
	AND U2148 ( .A(w2528), .B(w2529), .Z(w2530) );
	AND U2149 ( .A(w2504), .B(w2444), .Z(w2531) );
	XOR U2150 ( .A(w2531), .B(w2530), .Z(w2532) );
	AND U2151 ( .A(w2506), .B(w2443), .Z(w2533) );
	XOR U2152 ( .A(w2533), .B(w2530), .Z(w2534) );
	XOR U2153 ( .A(w2511), .B(w2513), .Z(w2535) );
	XOR U2154 ( .A(w2442), .B(w2441), .Z(w2536) );
	AND U2155 ( .A(w2535), .B(w2536), .Z(w2537) );
	AND U2156 ( .A(w2511), .B(w2442), .Z(w2538) );
	XOR U2157 ( .A(w2538), .B(w2537), .Z(w2539) );
	AND U2158 ( .A(w2513), .B(w2441), .Z(w2540) );
	XOR U2159 ( .A(w2540), .B(w2537), .Z(w2541) );
	XOR U2160 ( .A(w2534), .B(w2527), .Z(w2542) );
	XOR U2161 ( .A(w2532), .B(w2526), .Z(w2543) );
	XOR U2162 ( .A(w2541), .B(w2527), .Z(w2544) );
	XOR U2163 ( .A(w2539), .B(w2526), .Z(w2545) );
	XOR U2164 ( .A(w2506), .B(w2513), .Z(w2548) );
	XOR U2165 ( .A(w2504), .B(w2511), .Z(w2549) );
	XOR U2166 ( .A(w2439), .B(w2437), .Z(w2550) );
	XOR U2167 ( .A(w2440), .B(w2438), .Z(w2551) );
	XOR U2168 ( .A(w2549), .B(w2548), .Z(w2552) );
	XOR U2169 ( .A(w2551), .B(w2550), .Z(w2553) );
	AND U2170 ( .A(w2552), .B(w2553), .Z(w2554) );
	AND U2171 ( .A(w2549), .B(w2551), .Z(w2555) );
	XOR U2172 ( .A(w2555), .B(w2554), .Z(w2556) );
	AND U2173 ( .A(w2548), .B(w2550), .Z(w2557) );
	XOR U2174 ( .A(w2557), .B(w2554), .Z(w2558) );
	XOR U2175 ( .A(w2558), .B(w2556), .Z(w2559) );
	XOR U2176 ( .A(w2504), .B(w2506), .Z(w2560) );
	XOR U2177 ( .A(w2440), .B(w2439), .Z(w2561) );
	AND U2178 ( .A(w2560), .B(w2561), .Z(w2562) );
	AND U2179 ( .A(w2504), .B(w2440), .Z(w2563) );
	XOR U2180 ( .A(w2563), .B(w2562), .Z(w2564) );
	AND U2181 ( .A(w2506), .B(w2439), .Z(w2565) );
	XOR U2182 ( .A(w2565), .B(w2562), .Z(w2566) );
	XOR U2183 ( .A(w2511), .B(w2513), .Z(w2567) );
	XOR U2184 ( .A(w2438), .B(w2437), .Z(w2568) );
	AND U2185 ( .A(w2567), .B(w2568), .Z(w2569) );
	AND U2186 ( .A(w2511), .B(w2438), .Z(w2570) );
	XOR U2187 ( .A(w2570), .B(w2569), .Z(w2571) );
	AND U2188 ( .A(w2513), .B(w2437), .Z(w2572) );
	XOR U2189 ( .A(w2572), .B(w2569), .Z(w2573) );
	XOR U2190 ( .A(w2566), .B(w2559), .Z(w2574) );
	XOR U2191 ( .A(w2564), .B(w2558), .Z(w2575) );
	XOR U2192 ( .A(w2573), .B(w2559), .Z(w2576) );
	XOR U2193 ( .A(w2571), .B(w2558), .Z(w2577) );
	XOR U2194 ( .A(w2580), .B(w2576), .Z(w2586) );
	XOR U2195 ( .A(w2581), .B(w2576), .Z(w2587) );
	XOR U2196 ( .A(w2585), .B(w2576), .Z(w2588) );
	XOR U2197 ( .A(w2578), .B(w2577), .Z(w2589) );
	XOR U2198 ( .A(w2587), .B(w2577), .Z(w2590) );
	XOR U2199 ( .A(w2582), .B(w2577), .Z(w2591) );
	XOR U2200 ( .A(w2583), .B(w2577), .Z(w2592) );
	XOR U2201 ( .A(w2584), .B(w2577), .Z(w2593) );
	XOR U2202 ( .A(w2589), .B(w2574), .Z(w2594) );
	XOR U2203 ( .A(w2586), .B(w2574), .Z(w2595) );
	XOR U2204 ( .A(w2594), .B(w2575), .Z(w2596) );
	XOR U2205 ( .A(w2579), .B(w2575), .Z(w2597) );
	XOR U2206 ( .A(w2590), .B(w2575), .Z(w2598) );
	XOR U2207 ( .A(w2592), .B(w2575), .Z(w2599) );
	XOR U2208 ( .A(w2593), .B(w2575), .Z(w2600) );
	XOR U2209 ( .A(w2588), .B(w2575), .Z(w2601) );
	XOR U2210 ( .A(w2597), .B(w2544), .Z(w2602) );
	XOR U2211 ( .A(w2591), .B(w2544), .Z(w2603) );
	XOR U2212 ( .A(w2595), .B(w2545), .Z(w2604) );
	XOR U2213 ( .A(w2596), .B(w2542), .Z(w2605) );
	XOR U2214 ( .A(w2603), .B(w2542), .Z(w2606) );
	XOR U2215 ( .A(w2600), .B(w2542), .Z(w2607) );
	XOR U2216 ( .A(w2605), .B(w2543), .Z(w2608) );
	XOR U2217 ( .A(w2602), .B(w2543), .Z(w2609) );
	XOR U2218 ( .A(w2606), .B(w2543), .Z(w2610) );
	XOR U2219 ( .A(w2607), .B(w2543), .Z(w2611) );
	XOR U2220 ( .A(w2615), .B(w96), .Z(w2620) );
	XOR U2221 ( .A(w2616), .B(w96), .Z(w2621) );
	XOR U2222 ( .A(w2619), .B(w96), .Z(w2622) );
	XOR U2223 ( .A(w2612), .B(w97), .Z(w2623) );
	XOR U2224 ( .A(w2613), .B(w97), .Z(w2624) );
	XOR U2225 ( .A(w2621), .B(w97), .Z(w2625) );
	XOR U2226 ( .A(w2617), .B(w97), .Z(w2626) );
	XOR U2227 ( .A(w2618), .B(w97), .Z(w2627) );
	XOR U2228 ( .A(w2622), .B(w97), .Z(w2628) );
	XOR U2229 ( .A(w2624), .B(w98), .Z(w2629) );
	XOR U2230 ( .A(w2625), .B(w98), .Z(w2630) );
	XOR U2231 ( .A(w2626), .B(w98), .Z(w2631) );
	XOR U2232 ( .A(w2627), .B(w98), .Z(w2632) );
	XOR U2233 ( .A(w2628), .B(w98), .Z(w2633) );
	XOR U2234 ( .A(w2620), .B(w99), .Z(w2634) );
	XOR U2235 ( .A(w2632), .B(w99), .Z(w2635) );
	XOR U2236 ( .A(w2623), .B(w100), .Z(w2636) );
	XOR U2237 ( .A(w2634), .B(w100), .Z(w2637) );
	XOR U2238 ( .A(w2636), .B(w101), .Z(w2638) );
	XOR U2239 ( .A(w2633), .B(w101), .Z(w2639) );
	XOR U2240 ( .A(w2638), .B(w102), .Z(w2640) );
	XOR U2241 ( .A(w2637), .B(w102), .Z(w2641) );
	XOR U2242 ( .A(w2631), .B(w102), .Z(w2642) );
	XOR U2243 ( .A(w2639), .B(w102), .Z(w2643) );
	XOR U2244 ( .A(w2640), .B(w103), .Z(w2644) );
	XOR U2245 ( .A(w2629), .B(w103), .Z(w2645) );
	XOR U2246 ( .A(w2614), .B(w103), .Z(w2646) );
	XOR U2247 ( .A(w2641), .B(w103), .Z(w2647) );
	XOR U2248 ( .A(w2630), .B(w103), .Z(w2648) );
	XOR U2249 ( .A(w2642), .B(w103), .Z(w2649) );
	XOR U2250 ( .A(w2635), .B(w103), .Z(w2650) );
	XOR U2251 ( .A(w2643), .B(w103), .Z(w2651) );
	XOR U2252 ( .A(w2644), .B(w2648), .Z(w2652) );
	XOR U2253 ( .A(w2645), .B(w2649), .Z(w2653) );
	XOR U2254 ( .A(w2646), .B(w2650), .Z(w2654) );
	XOR U2255 ( .A(w2647), .B(w2651), .Z(w2655) );
	XOR U2256 ( .A(w2654), .B(w2652), .Z(w2656) );
	XOR U2257 ( .A(w2655), .B(w2653), .Z(w2657) );
	XOR U2258 ( .A(w2653), .B(w2652), .Z(w2658) );
	XOR U2259 ( .A(w2646), .B(w2644), .Z(w2661) );
	XOR U2260 ( .A(w2647), .B(w2645), .Z(w2662) );
	XOR U2261 ( .A(w2650), .B(w2648), .Z(w2663) );
	XOR U2262 ( .A(w2651), .B(w2649), .Z(w2664) );
	XOR U2263 ( .A(w2662), .B(w2661), .Z(w2665) );
	XOR U2264 ( .A(w2664), .B(w2663), .Z(w2666) );
	AND U2265 ( .A(w2665), .B(w2666), .Z(w2667) );
	AND U2266 ( .A(w2662), .B(w2664), .Z(w2668) );
	XOR U2267 ( .A(w2668), .B(w2667), .Z(w2669) );
	AND U2268 ( .A(w2661), .B(w2663), .Z(w2670) );
	XOR U2269 ( .A(w2670), .B(w2667), .Z(w2671) );
	XOR U2270 ( .A(w2671), .B(w2669), .Z(w2672) );
	XOR U2271 ( .A(w2647), .B(w2646), .Z(w2673) );
	XOR U2272 ( .A(w2651), .B(w2650), .Z(w2674) );
	AND U2273 ( .A(w2673), .B(w2674), .Z(w2675) );
	AND U2274 ( .A(w2647), .B(w2651), .Z(w2676) );
	XOR U2275 ( .A(w2676), .B(w2675), .Z(w2677) );
	AND U2276 ( .A(w2646), .B(w2650), .Z(w2678) );
	XOR U2277 ( .A(w2678), .B(w2675), .Z(w2679) );
	XOR U2278 ( .A(w2645), .B(w2644), .Z(w2680) );
	XOR U2279 ( .A(w2649), .B(w2648), .Z(w2681) );
	AND U2280 ( .A(w2680), .B(w2681), .Z(w2682) );
	AND U2281 ( .A(w2645), .B(w2649), .Z(w2683) );
	XOR U2282 ( .A(w2683), .B(w2682), .Z(w2684) );
	AND U2283 ( .A(w2644), .B(w2648), .Z(w2685) );
	XOR U2284 ( .A(w2685), .B(w2682), .Z(w2686) );
	XOR U2285 ( .A(w2679), .B(w2672), .Z(w2687) );
	XOR U2286 ( .A(w2677), .B(w2671), .Z(w2688) );
	XOR U2287 ( .A(w2686), .B(w2672), .Z(w2689) );
	XOR U2288 ( .A(w2684), .B(w2671), .Z(w2690) );
	XOR U2289 ( .A(w2652), .B(w2689), .Z(w2691) );
	XOR U2290 ( .A(w2658), .B(w2690), .Z(w2692) );
	XOR U2291 ( .A(w2657), .B(w2687), .Z(w2693) );
	XOR U2292 ( .A(w2656), .B(w2688), .Z(w2694) );
	XOR U2293 ( .A(w2693), .B(w2691), .Z(w2695) );
	XOR U2294 ( .A(w2694), .B(w2692), .Z(w2696) );
	XOR U2295 ( .A(w2696), .B(w2695), .Z(w2697) );
	XOR U2296 ( .A(w2694), .B(w2693), .Z(w2698) );
	XOR U2297 ( .A(w2692), .B(w2691), .Z(w2699) );
	AND U2298 ( .A(w2698), .B(w2699), .Z(w2700) );
	AND U2299 ( .A(w2694), .B(w2692), .Z(w2701) );
	XOR U2300 ( .A(w2701), .B(w2700), .Z(w2702) );
	AND U2301 ( .A(w2693), .B(w2691), .Z(w2703) );
	XOR U2302 ( .A(w2703), .B(w2700), .Z(w2704) );
	XOR U2303 ( .A(w2697), .B(w2704), .Z(w2705) );
	XOR U2304 ( .A(w2696), .B(w2702), .Z(w2706) );
	XOR U2305 ( .A(w2705), .B(w2706), .Z(w2707) );
	XOR U2306 ( .A(w2692), .B(w2691), .Z(w2708) );
	AND U2307 ( .A(w2707), .B(w2708), .Z(w2709) );
	AND U2308 ( .A(w2705), .B(w2692), .Z(w2710) );
	XOR U2309 ( .A(w2710), .B(w2709), .Z(w2711) );
	AND U2310 ( .A(w2706), .B(w2691), .Z(w2712) );
	XOR U2311 ( .A(w2712), .B(w2709), .Z(w2713) );
	XOR U2312 ( .A(w2705), .B(w2706), .Z(w2714) );
	XOR U2313 ( .A(w2694), .B(w2693), .Z(w2715) );
	AND U2314 ( .A(w2714), .B(w2715), .Z(w2716) );
	AND U2315 ( .A(w2705), .B(w2694), .Z(w2717) );
	XOR U2316 ( .A(w2717), .B(w2716), .Z(w2718) );
	AND U2317 ( .A(w2706), .B(w2693), .Z(w2719) );
	XOR U2318 ( .A(w2719), .B(w2716), .Z(w2720) );
	XOR U2319 ( .A(w2713), .B(w2720), .Z(w2723) );
	XOR U2320 ( .A(w2711), .B(w2718), .Z(w2724) );
	XOR U2321 ( .A(w2650), .B(w2648), .Z(w2725) );
	XOR U2322 ( .A(w2651), .B(w2649), .Z(w2726) );
	XOR U2323 ( .A(w2724), .B(w2723), .Z(w2727) );
	XOR U2324 ( .A(w2726), .B(w2725), .Z(w2728) );
	AND U2325 ( .A(w2727), .B(w2728), .Z(w2729) );
	AND U2326 ( .A(w2724), .B(w2726), .Z(w2730) );
	XOR U2327 ( .A(w2730), .B(w2729), .Z(w2731) );
	AND U2328 ( .A(w2723), .B(w2725), .Z(w2732) );
	XOR U2329 ( .A(w2732), .B(w2729), .Z(w2733) );
	XOR U2330 ( .A(w2733), .B(w2731), .Z(w2734) );
	XOR U2331 ( .A(w2711), .B(w2713), .Z(w2735) );
	XOR U2332 ( .A(w2651), .B(w2650), .Z(w2736) );
	AND U2333 ( .A(w2735), .B(w2736), .Z(w2737) );
	AND U2334 ( .A(w2711), .B(w2651), .Z(w2738) );
	XOR U2335 ( .A(w2738), .B(w2737), .Z(w2739) );
	AND U2336 ( .A(w2713), .B(w2650), .Z(w2740) );
	XOR U2337 ( .A(w2740), .B(w2737), .Z(w2741) );
	XOR U2338 ( .A(w2718), .B(w2720), .Z(w2742) );
	XOR U2339 ( .A(w2649), .B(w2648), .Z(w2743) );
	AND U2340 ( .A(w2742), .B(w2743), .Z(w2744) );
	AND U2341 ( .A(w2718), .B(w2649), .Z(w2745) );
	XOR U2342 ( .A(w2745), .B(w2744), .Z(w2746) );
	AND U2343 ( .A(w2720), .B(w2648), .Z(w2747) );
	XOR U2344 ( .A(w2747), .B(w2744), .Z(w2748) );
	XOR U2345 ( .A(w2741), .B(w2734), .Z(w2749) );
	XOR U2346 ( .A(w2739), .B(w2733), .Z(w2750) );
	XOR U2347 ( .A(w2748), .B(w2734), .Z(w2751) );
	XOR U2348 ( .A(w2746), .B(w2733), .Z(w2752) );
	XOR U2349 ( .A(w2713), .B(w2720), .Z(w2755) );
	XOR U2350 ( .A(w2711), .B(w2718), .Z(w2756) );
	XOR U2351 ( .A(w2646), .B(w2644), .Z(w2757) );
	XOR U2352 ( .A(w2647), .B(w2645), .Z(w2758) );
	XOR U2353 ( .A(w2756), .B(w2755), .Z(w2759) );
	XOR U2354 ( .A(w2758), .B(w2757), .Z(w2760) );
	AND U2355 ( .A(w2759), .B(w2760), .Z(w2761) );
	AND U2356 ( .A(w2756), .B(w2758), .Z(w2762) );
	XOR U2357 ( .A(w2762), .B(w2761), .Z(w2763) );
	AND U2358 ( .A(w2755), .B(w2757), .Z(w2764) );
	XOR U2359 ( .A(w2764), .B(w2761), .Z(w2765) );
	XOR U2360 ( .A(w2765), .B(w2763), .Z(w2766) );
	XOR U2361 ( .A(w2711), .B(w2713), .Z(w2767) );
	XOR U2362 ( .A(w2647), .B(w2646), .Z(w2768) );
	AND U2363 ( .A(w2767), .B(w2768), .Z(w2769) );
	AND U2364 ( .A(w2711), .B(w2647), .Z(w2770) );
	XOR U2365 ( .A(w2770), .B(w2769), .Z(w2771) );
	AND U2366 ( .A(w2713), .B(w2646), .Z(w2772) );
	XOR U2367 ( .A(w2772), .B(w2769), .Z(w2773) );
	XOR U2368 ( .A(w2718), .B(w2720), .Z(w2774) );
	XOR U2369 ( .A(w2645), .B(w2644), .Z(w2775) );
	AND U2370 ( .A(w2774), .B(w2775), .Z(w2776) );
	AND U2371 ( .A(w2718), .B(w2645), .Z(w2777) );
	XOR U2372 ( .A(w2777), .B(w2776), .Z(w2778) );
	AND U2373 ( .A(w2720), .B(w2644), .Z(w2779) );
	XOR U2374 ( .A(w2779), .B(w2776), .Z(w2780) );
	XOR U2375 ( .A(w2773), .B(w2766), .Z(w2781) );
	XOR U2376 ( .A(w2771), .B(w2765), .Z(w2782) );
	XOR U2377 ( .A(w2780), .B(w2766), .Z(w2783) );
	XOR U2378 ( .A(w2778), .B(w2765), .Z(w2784) );
	XOR U2379 ( .A(w2787), .B(w2783), .Z(w2793) );
	XOR U2380 ( .A(w2788), .B(w2783), .Z(w2794) );
	XOR U2381 ( .A(w2792), .B(w2783), .Z(w2795) );
	XOR U2382 ( .A(w2785), .B(w2784), .Z(w2796) );
	XOR U2383 ( .A(w2794), .B(w2784), .Z(w2797) );
	XOR U2384 ( .A(w2789), .B(w2784), .Z(w2798) );
	XOR U2385 ( .A(w2790), .B(w2784), .Z(w2799) );
	XOR U2386 ( .A(w2791), .B(w2784), .Z(w2800) );
	XOR U2387 ( .A(w2796), .B(w2781), .Z(w2801) );
	XOR U2388 ( .A(w2793), .B(w2781), .Z(w2802) );
	XOR U2389 ( .A(w2801), .B(w2782), .Z(w2803) );
	XOR U2390 ( .A(w2786), .B(w2782), .Z(w2804) );
	XOR U2391 ( .A(w2797), .B(w2782), .Z(w2805) );
	XOR U2392 ( .A(w2799), .B(w2782), .Z(w2806) );
	XOR U2393 ( .A(w2800), .B(w2782), .Z(w2807) );
	XOR U2394 ( .A(w2795), .B(w2782), .Z(w2808) );
	XOR U2395 ( .A(w2804), .B(w2751), .Z(w2809) );
	XOR U2396 ( .A(w2798), .B(w2751), .Z(w2810) );
	XOR U2397 ( .A(w2802), .B(w2752), .Z(w2811) );
	XOR U2398 ( .A(w2803), .B(w2749), .Z(w2812) );
	XOR U2399 ( .A(w2810), .B(w2749), .Z(w2813) );
	XOR U2400 ( .A(w2807), .B(w2749), .Z(w2814) );
	XOR U2401 ( .A(w2812), .B(w2750), .Z(w2815) );
	XOR U2402 ( .A(w2809), .B(w2750), .Z(w2816) );
	XOR U2403 ( .A(w2813), .B(w2750), .Z(w2817) );
	XOR U2404 ( .A(w2814), .B(w2750), .Z(w2818) );
	XOR U2405 ( .A(w2822), .B(w104), .Z(w2827) );
	XOR U2406 ( .A(w2823), .B(w104), .Z(w2828) );
	XOR U2407 ( .A(w2826), .B(w104), .Z(w2829) );
	XOR U2408 ( .A(w2819), .B(w105), .Z(w2830) );
	XOR U2409 ( .A(w2820), .B(w105), .Z(w2831) );
	XOR U2410 ( .A(w2828), .B(w105), .Z(w2832) );
	XOR U2411 ( .A(w2824), .B(w105), .Z(w2833) );
	XOR U2412 ( .A(w2825), .B(w105), .Z(w2834) );
	XOR U2413 ( .A(w2829), .B(w105), .Z(w2835) );
	XOR U2414 ( .A(w2831), .B(w106), .Z(w2836) );
	XOR U2415 ( .A(w2832), .B(w106), .Z(w2837) );
	XOR U2416 ( .A(w2833), .B(w106), .Z(w2838) );
	XOR U2417 ( .A(w2834), .B(w106), .Z(w2839) );
	XOR U2418 ( .A(w2835), .B(w106), .Z(w2840) );
	XOR U2419 ( .A(w2827), .B(w107), .Z(w2841) );
	XOR U2420 ( .A(w2839), .B(w107), .Z(w2842) );
	XOR U2421 ( .A(w2830), .B(w108), .Z(w2843) );
	XOR U2422 ( .A(w2841), .B(w108), .Z(w2844) );
	XOR U2423 ( .A(w2843), .B(w109), .Z(w2845) );
	XOR U2424 ( .A(w2840), .B(w109), .Z(w2846) );
	XOR U2425 ( .A(w2845), .B(w110), .Z(w2847) );
	XOR U2426 ( .A(w2844), .B(w110), .Z(w2848) );
	XOR U2427 ( .A(w2838), .B(w110), .Z(w2849) );
	XOR U2428 ( .A(w2846), .B(w110), .Z(w2850) );
	XOR U2429 ( .A(w2847), .B(w111), .Z(w2851) );
	XOR U2430 ( .A(w2836), .B(w111), .Z(w2852) );
	XOR U2431 ( .A(w2821), .B(w111), .Z(w2853) );
	XOR U2432 ( .A(w2848), .B(w111), .Z(w2854) );
	XOR U2433 ( .A(w2837), .B(w111), .Z(w2855) );
	XOR U2434 ( .A(w2849), .B(w111), .Z(w2856) );
	XOR U2435 ( .A(w2842), .B(w111), .Z(w2857) );
	XOR U2436 ( .A(w2850), .B(w111), .Z(w2858) );
	XOR U2437 ( .A(w2851), .B(w2855), .Z(w2859) );
	XOR U2438 ( .A(w2852), .B(w2856), .Z(w2860) );
	XOR U2439 ( .A(w2853), .B(w2857), .Z(w2861) );
	XOR U2440 ( .A(w2854), .B(w2858), .Z(w2862) );
	XOR U2441 ( .A(w2861), .B(w2859), .Z(w2863) );
	XOR U2442 ( .A(w2862), .B(w2860), .Z(w2864) );
	XOR U2443 ( .A(w2860), .B(w2859), .Z(w2865) );
	XOR U2444 ( .A(w2853), .B(w2851), .Z(w2868) );
	XOR U2445 ( .A(w2854), .B(w2852), .Z(w2869) );
	XOR U2446 ( .A(w2857), .B(w2855), .Z(w2870) );
	XOR U2447 ( .A(w2858), .B(w2856), .Z(w2871) );
	XOR U2448 ( .A(w2869), .B(w2868), .Z(w2872) );
	XOR U2449 ( .A(w2871), .B(w2870), .Z(w2873) );
	AND U2450 ( .A(w2872), .B(w2873), .Z(w2874) );
	AND U2451 ( .A(w2869), .B(w2871), .Z(w2875) );
	XOR U2452 ( .A(w2875), .B(w2874), .Z(w2876) );
	AND U2453 ( .A(w2868), .B(w2870), .Z(w2877) );
	XOR U2454 ( .A(w2877), .B(w2874), .Z(w2878) );
	XOR U2455 ( .A(w2878), .B(w2876), .Z(w2879) );
	XOR U2456 ( .A(w2854), .B(w2853), .Z(w2880) );
	XOR U2457 ( .A(w2858), .B(w2857), .Z(w2881) );
	AND U2458 ( .A(w2880), .B(w2881), .Z(w2882) );
	AND U2459 ( .A(w2854), .B(w2858), .Z(w2883) );
	XOR U2460 ( .A(w2883), .B(w2882), .Z(w2884) );
	AND U2461 ( .A(w2853), .B(w2857), .Z(w2885) );
	XOR U2462 ( .A(w2885), .B(w2882), .Z(w2886) );
	XOR U2463 ( .A(w2852), .B(w2851), .Z(w2887) );
	XOR U2464 ( .A(w2856), .B(w2855), .Z(w2888) );
	AND U2465 ( .A(w2887), .B(w2888), .Z(w2889) );
	AND U2466 ( .A(w2852), .B(w2856), .Z(w2890) );
	XOR U2467 ( .A(w2890), .B(w2889), .Z(w2891) );
	AND U2468 ( .A(w2851), .B(w2855), .Z(w2892) );
	XOR U2469 ( .A(w2892), .B(w2889), .Z(w2893) );
	XOR U2470 ( .A(w2886), .B(w2879), .Z(w2894) );
	XOR U2471 ( .A(w2884), .B(w2878), .Z(w2895) );
	XOR U2472 ( .A(w2893), .B(w2879), .Z(w2896) );
	XOR U2473 ( .A(w2891), .B(w2878), .Z(w2897) );
	XOR U2474 ( .A(w2859), .B(w2896), .Z(w2898) );
	XOR U2475 ( .A(w2865), .B(w2897), .Z(w2899) );
	XOR U2476 ( .A(w2864), .B(w2894), .Z(w2900) );
	XOR U2477 ( .A(w2863), .B(w2895), .Z(w2901) );
	XOR U2478 ( .A(w2900), .B(w2898), .Z(w2902) );
	XOR U2479 ( .A(w2901), .B(w2899), .Z(w2903) );
	XOR U2480 ( .A(w2903), .B(w2902), .Z(w2904) );
	XOR U2481 ( .A(w2901), .B(w2900), .Z(w2905) );
	XOR U2482 ( .A(w2899), .B(w2898), .Z(w2906) );
	AND U2483 ( .A(w2905), .B(w2906), .Z(w2907) );
	AND U2484 ( .A(w2901), .B(w2899), .Z(w2908) );
	XOR U2485 ( .A(w2908), .B(w2907), .Z(w2909) );
	AND U2486 ( .A(w2900), .B(w2898), .Z(w2910) );
	XOR U2487 ( .A(w2910), .B(w2907), .Z(w2911) );
	XOR U2488 ( .A(w2904), .B(w2911), .Z(w2912) );
	XOR U2489 ( .A(w2903), .B(w2909), .Z(w2913) );
	XOR U2490 ( .A(w2912), .B(w2913), .Z(w2914) );
	XOR U2491 ( .A(w2899), .B(w2898), .Z(w2915) );
	AND U2492 ( .A(w2914), .B(w2915), .Z(w2916) );
	AND U2493 ( .A(w2912), .B(w2899), .Z(w2917) );
	XOR U2494 ( .A(w2917), .B(w2916), .Z(w2918) );
	AND U2495 ( .A(w2913), .B(w2898), .Z(w2919) );
	XOR U2496 ( .A(w2919), .B(w2916), .Z(w2920) );
	XOR U2497 ( .A(w2912), .B(w2913), .Z(w2921) );
	XOR U2498 ( .A(w2901), .B(w2900), .Z(w2922) );
	AND U2499 ( .A(w2921), .B(w2922), .Z(w2923) );
	AND U2500 ( .A(w2912), .B(w2901), .Z(w2924) );
	XOR U2501 ( .A(w2924), .B(w2923), .Z(w2925) );
	AND U2502 ( .A(w2913), .B(w2900), .Z(w2926) );
	XOR U2503 ( .A(w2926), .B(w2923), .Z(w2927) );
	XOR U2504 ( .A(w2920), .B(w2927), .Z(w2930) );
	XOR U2505 ( .A(w2918), .B(w2925), .Z(w2931) );
	XOR U2506 ( .A(w2857), .B(w2855), .Z(w2932) );
	XOR U2507 ( .A(w2858), .B(w2856), .Z(w2933) );
	XOR U2508 ( .A(w2931), .B(w2930), .Z(w2934) );
	XOR U2509 ( .A(w2933), .B(w2932), .Z(w2935) );
	AND U2510 ( .A(w2934), .B(w2935), .Z(w2936) );
	AND U2511 ( .A(w2931), .B(w2933), .Z(w2937) );
	XOR U2512 ( .A(w2937), .B(w2936), .Z(w2938) );
	AND U2513 ( .A(w2930), .B(w2932), .Z(w2939) );
	XOR U2514 ( .A(w2939), .B(w2936), .Z(w2940) );
	XOR U2515 ( .A(w2940), .B(w2938), .Z(w2941) );
	XOR U2516 ( .A(w2918), .B(w2920), .Z(w2942) );
	XOR U2517 ( .A(w2858), .B(w2857), .Z(w2943) );
	AND U2518 ( .A(w2942), .B(w2943), .Z(w2944) );
	AND U2519 ( .A(w2918), .B(w2858), .Z(w2945) );
	XOR U2520 ( .A(w2945), .B(w2944), .Z(w2946) );
	AND U2521 ( .A(w2920), .B(w2857), .Z(w2947) );
	XOR U2522 ( .A(w2947), .B(w2944), .Z(w2948) );
	XOR U2523 ( .A(w2925), .B(w2927), .Z(w2949) );
	XOR U2524 ( .A(w2856), .B(w2855), .Z(w2950) );
	AND U2525 ( .A(w2949), .B(w2950), .Z(w2951) );
	AND U2526 ( .A(w2925), .B(w2856), .Z(w2952) );
	XOR U2527 ( .A(w2952), .B(w2951), .Z(w2953) );
	AND U2528 ( .A(w2927), .B(w2855), .Z(w2954) );
	XOR U2529 ( .A(w2954), .B(w2951), .Z(w2955) );
	XOR U2530 ( .A(w2948), .B(w2941), .Z(w2956) );
	XOR U2531 ( .A(w2946), .B(w2940), .Z(w2957) );
	XOR U2532 ( .A(w2955), .B(w2941), .Z(w2958) );
	XOR U2533 ( .A(w2953), .B(w2940), .Z(w2959) );
	XOR U2534 ( .A(w2920), .B(w2927), .Z(w2962) );
	XOR U2535 ( .A(w2918), .B(w2925), .Z(w2963) );
	XOR U2536 ( .A(w2853), .B(w2851), .Z(w2964) );
	XOR U2537 ( .A(w2854), .B(w2852), .Z(w2965) );
	XOR U2538 ( .A(w2963), .B(w2962), .Z(w2966) );
	XOR U2539 ( .A(w2965), .B(w2964), .Z(w2967) );
	AND U2540 ( .A(w2966), .B(w2967), .Z(w2968) );
	AND U2541 ( .A(w2963), .B(w2965), .Z(w2969) );
	XOR U2542 ( .A(w2969), .B(w2968), .Z(w2970) );
	AND U2543 ( .A(w2962), .B(w2964), .Z(w2971) );
	XOR U2544 ( .A(w2971), .B(w2968), .Z(w2972) );
	XOR U2545 ( .A(w2972), .B(w2970), .Z(w2973) );
	XOR U2546 ( .A(w2918), .B(w2920), .Z(w2974) );
	XOR U2547 ( .A(w2854), .B(w2853), .Z(w2975) );
	AND U2548 ( .A(w2974), .B(w2975), .Z(w2976) );
	AND U2549 ( .A(w2918), .B(w2854), .Z(w2977) );
	XOR U2550 ( .A(w2977), .B(w2976), .Z(w2978) );
	AND U2551 ( .A(w2920), .B(w2853), .Z(w2979) );
	XOR U2552 ( .A(w2979), .B(w2976), .Z(w2980) );
	XOR U2553 ( .A(w2925), .B(w2927), .Z(w2981) );
	XOR U2554 ( .A(w2852), .B(w2851), .Z(w2982) );
	AND U2555 ( .A(w2981), .B(w2982), .Z(w2983) );
	AND U2556 ( .A(w2925), .B(w2852), .Z(w2984) );
	XOR U2557 ( .A(w2984), .B(w2983), .Z(w2985) );
	AND U2558 ( .A(w2927), .B(w2851), .Z(w2986) );
	XOR U2559 ( .A(w2986), .B(w2983), .Z(w2987) );
	XOR U2560 ( .A(w2980), .B(w2973), .Z(w2988) );
	XOR U2561 ( .A(w2978), .B(w2972), .Z(w2989) );
	XOR U2562 ( .A(w2987), .B(w2973), .Z(w2990) );
	XOR U2563 ( .A(w2985), .B(w2972), .Z(w2991) );
	XOR U2564 ( .A(w2994), .B(w2990), .Z(w3000) );
	XOR U2565 ( .A(w2995), .B(w2990), .Z(w3001) );
	XOR U2566 ( .A(w2999), .B(w2990), .Z(w3002) );
	XOR U2567 ( .A(w2992), .B(w2991), .Z(w3003) );
	XOR U2568 ( .A(w3001), .B(w2991), .Z(w3004) );
	XOR U2569 ( .A(w2996), .B(w2991), .Z(w3005) );
	XOR U2570 ( .A(w2997), .B(w2991), .Z(w3006) );
	XOR U2571 ( .A(w2998), .B(w2991), .Z(w3007) );
	XOR U2572 ( .A(w3003), .B(w2988), .Z(w3008) );
	XOR U2573 ( .A(w3000), .B(w2988), .Z(w3009) );
	XOR U2574 ( .A(w3008), .B(w2989), .Z(w3010) );
	XOR U2575 ( .A(w2993), .B(w2989), .Z(w3011) );
	XOR U2576 ( .A(w3004), .B(w2989), .Z(w3012) );
	XOR U2577 ( .A(w3006), .B(w2989), .Z(w3013) );
	XOR U2578 ( .A(w3007), .B(w2989), .Z(w3014) );
	XOR U2579 ( .A(w3002), .B(w2989), .Z(w3015) );
	XOR U2580 ( .A(w3011), .B(w2958), .Z(w3016) );
	XOR U2581 ( .A(w3005), .B(w2958), .Z(w3017) );
	XOR U2582 ( .A(w3009), .B(w2959), .Z(w3018) );
	XOR U2583 ( .A(w3010), .B(w2956), .Z(w3019) );
	XOR U2584 ( .A(w3017), .B(w2956), .Z(w3020) );
	XOR U2585 ( .A(w3014), .B(w2956), .Z(w3021) );
	XOR U2586 ( .A(w3019), .B(w2957), .Z(w3022) );
	XOR U2587 ( .A(w3016), .B(w2957), .Z(w3023) );
	XOR U2588 ( .A(w3020), .B(w2957), .Z(w3024) );
	XOR U2589 ( .A(w3021), .B(w2957), .Z(w3025) );
	XOR U2590 ( .A(w3029), .B(w112), .Z(w3034) );
	XOR U2591 ( .A(w3030), .B(w112), .Z(w3035) );
	XOR U2592 ( .A(w3033), .B(w112), .Z(w3036) );
	XOR U2593 ( .A(w3026), .B(w113), .Z(w3037) );
	XOR U2594 ( .A(w3027), .B(w113), .Z(w3038) );
	XOR U2595 ( .A(w3035), .B(w113), .Z(w3039) );
	XOR U2596 ( .A(w3031), .B(w113), .Z(w3040) );
	XOR U2597 ( .A(w3032), .B(w113), .Z(w3041) );
	XOR U2598 ( .A(w3036), .B(w113), .Z(w3042) );
	XOR U2599 ( .A(w3038), .B(w114), .Z(w3043) );
	XOR U2600 ( .A(w3039), .B(w114), .Z(w3044) );
	XOR U2601 ( .A(w3040), .B(w114), .Z(w3045) );
	XOR U2602 ( .A(w3041), .B(w114), .Z(w3046) );
	XOR U2603 ( .A(w3042), .B(w114), .Z(w3047) );
	XOR U2604 ( .A(w3034), .B(w115), .Z(w3048) );
	XOR U2605 ( .A(w3046), .B(w115), .Z(w3049) );
	XOR U2606 ( .A(w3037), .B(w116), .Z(w3050) );
	XOR U2607 ( .A(w3048), .B(w116), .Z(w3051) );
	XOR U2608 ( .A(w3050), .B(w117), .Z(w3052) );
	XOR U2609 ( .A(w3047), .B(w117), .Z(w3053) );
	XOR U2610 ( .A(w3052), .B(w118), .Z(w3054) );
	XOR U2611 ( .A(w3051), .B(w118), .Z(w3055) );
	XOR U2612 ( .A(w3045), .B(w118), .Z(w3056) );
	XOR U2613 ( .A(w3053), .B(w118), .Z(w3057) );
	XOR U2614 ( .A(w3054), .B(w119), .Z(w3058) );
	XOR U2615 ( .A(w3043), .B(w119), .Z(w3059) );
	XOR U2616 ( .A(w3028), .B(w119), .Z(w3060) );
	XOR U2617 ( .A(w3055), .B(w119), .Z(w3061) );
	XOR U2618 ( .A(w3044), .B(w119), .Z(w3062) );
	XOR U2619 ( .A(w3056), .B(w119), .Z(w3063) );
	XOR U2620 ( .A(w3049), .B(w119), .Z(w3064) );
	XOR U2621 ( .A(w3057), .B(w119), .Z(w3065) );
	XOR U2622 ( .A(w3058), .B(w3062), .Z(w3066) );
	XOR U2623 ( .A(w3059), .B(w3063), .Z(w3067) );
	XOR U2624 ( .A(w3060), .B(w3064), .Z(w3068) );
	XOR U2625 ( .A(w3061), .B(w3065), .Z(w3069) );
	XOR U2626 ( .A(w3068), .B(w3066), .Z(w3070) );
	XOR U2627 ( .A(w3069), .B(w3067), .Z(w3071) );
	XOR U2628 ( .A(w3067), .B(w3066), .Z(w3072) );
	XOR U2629 ( .A(w3060), .B(w3058), .Z(w3075) );
	XOR U2630 ( .A(w3061), .B(w3059), .Z(w3076) );
	XOR U2631 ( .A(w3064), .B(w3062), .Z(w3077) );
	XOR U2632 ( .A(w3065), .B(w3063), .Z(w3078) );
	XOR U2633 ( .A(w3076), .B(w3075), .Z(w3079) );
	XOR U2634 ( .A(w3078), .B(w3077), .Z(w3080) );
	AND U2635 ( .A(w3079), .B(w3080), .Z(w3081) );
	AND U2636 ( .A(w3076), .B(w3078), .Z(w3082) );
	XOR U2637 ( .A(w3082), .B(w3081), .Z(w3083) );
	AND U2638 ( .A(w3075), .B(w3077), .Z(w3084) );
	XOR U2639 ( .A(w3084), .B(w3081), .Z(w3085) );
	XOR U2640 ( .A(w3085), .B(w3083), .Z(w3086) );
	XOR U2641 ( .A(w3061), .B(w3060), .Z(w3087) );
	XOR U2642 ( .A(w3065), .B(w3064), .Z(w3088) );
	AND U2643 ( .A(w3087), .B(w3088), .Z(w3089) );
	AND U2644 ( .A(w3061), .B(w3065), .Z(w3090) );
	XOR U2645 ( .A(w3090), .B(w3089), .Z(w3091) );
	AND U2646 ( .A(w3060), .B(w3064), .Z(w3092) );
	XOR U2647 ( .A(w3092), .B(w3089), .Z(w3093) );
	XOR U2648 ( .A(w3059), .B(w3058), .Z(w3094) );
	XOR U2649 ( .A(w3063), .B(w3062), .Z(w3095) );
	AND U2650 ( .A(w3094), .B(w3095), .Z(w3096) );
	AND U2651 ( .A(w3059), .B(w3063), .Z(w3097) );
	XOR U2652 ( .A(w3097), .B(w3096), .Z(w3098) );
	AND U2653 ( .A(w3058), .B(w3062), .Z(w3099) );
	XOR U2654 ( .A(w3099), .B(w3096), .Z(w3100) );
	XOR U2655 ( .A(w3093), .B(w3086), .Z(w3101) );
	XOR U2656 ( .A(w3091), .B(w3085), .Z(w3102) );
	XOR U2657 ( .A(w3100), .B(w3086), .Z(w3103) );
	XOR U2658 ( .A(w3098), .B(w3085), .Z(w3104) );
	XOR U2659 ( .A(w3066), .B(w3103), .Z(w3105) );
	XOR U2660 ( .A(w3072), .B(w3104), .Z(w3106) );
	XOR U2661 ( .A(w3071), .B(w3101), .Z(w3107) );
	XOR U2662 ( .A(w3070), .B(w3102), .Z(w3108) );
	XOR U2663 ( .A(w3107), .B(w3105), .Z(w3109) );
	XOR U2664 ( .A(w3108), .B(w3106), .Z(w3110) );
	XOR U2665 ( .A(w3110), .B(w3109), .Z(w3111) );
	XOR U2666 ( .A(w3108), .B(w3107), .Z(w3112) );
	XOR U2667 ( .A(w3106), .B(w3105), .Z(w3113) );
	AND U2668 ( .A(w3112), .B(w3113), .Z(w3114) );
	AND U2669 ( .A(w3108), .B(w3106), .Z(w3115) );
	XOR U2670 ( .A(w3115), .B(w3114), .Z(w3116) );
	AND U2671 ( .A(w3107), .B(w3105), .Z(w3117) );
	XOR U2672 ( .A(w3117), .B(w3114), .Z(w3118) );
	XOR U2673 ( .A(w3111), .B(w3118), .Z(w3119) );
	XOR U2674 ( .A(w3110), .B(w3116), .Z(w3120) );
	XOR U2675 ( .A(w3119), .B(w3120), .Z(w3121) );
	XOR U2676 ( .A(w3106), .B(w3105), .Z(w3122) );
	AND U2677 ( .A(w3121), .B(w3122), .Z(w3123) );
	AND U2678 ( .A(w3119), .B(w3106), .Z(w3124) );
	XOR U2679 ( .A(w3124), .B(w3123), .Z(w3125) );
	AND U2680 ( .A(w3120), .B(w3105), .Z(w3126) );
	XOR U2681 ( .A(w3126), .B(w3123), .Z(w3127) );
	XOR U2682 ( .A(w3119), .B(w3120), .Z(w3128) );
	XOR U2683 ( .A(w3108), .B(w3107), .Z(w3129) );
	AND U2684 ( .A(w3128), .B(w3129), .Z(w3130) );
	AND U2685 ( .A(w3119), .B(w3108), .Z(w3131) );
	XOR U2686 ( .A(w3131), .B(w3130), .Z(w3132) );
	AND U2687 ( .A(w3120), .B(w3107), .Z(w3133) );
	XOR U2688 ( .A(w3133), .B(w3130), .Z(w3134) );
	XOR U2689 ( .A(w3127), .B(w3134), .Z(w3137) );
	XOR U2690 ( .A(w3125), .B(w3132), .Z(w3138) );
	XOR U2691 ( .A(w3064), .B(w3062), .Z(w3139) );
	XOR U2692 ( .A(w3065), .B(w3063), .Z(w3140) );
	XOR U2693 ( .A(w3138), .B(w3137), .Z(w3141) );
	XOR U2694 ( .A(w3140), .B(w3139), .Z(w3142) );
	AND U2695 ( .A(w3141), .B(w3142), .Z(w3143) );
	AND U2696 ( .A(w3138), .B(w3140), .Z(w3144) );
	XOR U2697 ( .A(w3144), .B(w3143), .Z(w3145) );
	AND U2698 ( .A(w3137), .B(w3139), .Z(w3146) );
	XOR U2699 ( .A(w3146), .B(w3143), .Z(w3147) );
	XOR U2700 ( .A(w3147), .B(w3145), .Z(w3148) );
	XOR U2701 ( .A(w3125), .B(w3127), .Z(w3149) );
	XOR U2702 ( .A(w3065), .B(w3064), .Z(w3150) );
	AND U2703 ( .A(w3149), .B(w3150), .Z(w3151) );
	AND U2704 ( .A(w3125), .B(w3065), .Z(w3152) );
	XOR U2705 ( .A(w3152), .B(w3151), .Z(w3153) );
	AND U2706 ( .A(w3127), .B(w3064), .Z(w3154) );
	XOR U2707 ( .A(w3154), .B(w3151), .Z(w3155) );
	XOR U2708 ( .A(w3132), .B(w3134), .Z(w3156) );
	XOR U2709 ( .A(w3063), .B(w3062), .Z(w3157) );
	AND U2710 ( .A(w3156), .B(w3157), .Z(w3158) );
	AND U2711 ( .A(w3132), .B(w3063), .Z(w3159) );
	XOR U2712 ( .A(w3159), .B(w3158), .Z(w3160) );
	AND U2713 ( .A(w3134), .B(w3062), .Z(w3161) );
	XOR U2714 ( .A(w3161), .B(w3158), .Z(w3162) );
	XOR U2715 ( .A(w3155), .B(w3148), .Z(w3163) );
	XOR U2716 ( .A(w3153), .B(w3147), .Z(w3164) );
	XOR U2717 ( .A(w3162), .B(w3148), .Z(w3165) );
	XOR U2718 ( .A(w3160), .B(w3147), .Z(w3166) );
	XOR U2719 ( .A(w3127), .B(w3134), .Z(w3169) );
	XOR U2720 ( .A(w3125), .B(w3132), .Z(w3170) );
	XOR U2721 ( .A(w3060), .B(w3058), .Z(w3171) );
	XOR U2722 ( .A(w3061), .B(w3059), .Z(w3172) );
	XOR U2723 ( .A(w3170), .B(w3169), .Z(w3173) );
	XOR U2724 ( .A(w3172), .B(w3171), .Z(w3174) );
	AND U2725 ( .A(w3173), .B(w3174), .Z(w3175) );
	AND U2726 ( .A(w3170), .B(w3172), .Z(w3176) );
	XOR U2727 ( .A(w3176), .B(w3175), .Z(w3177) );
	AND U2728 ( .A(w3169), .B(w3171), .Z(w3178) );
	XOR U2729 ( .A(w3178), .B(w3175), .Z(w3179) );
	XOR U2730 ( .A(w3179), .B(w3177), .Z(w3180) );
	XOR U2731 ( .A(w3125), .B(w3127), .Z(w3181) );
	XOR U2732 ( .A(w3061), .B(w3060), .Z(w3182) );
	AND U2733 ( .A(w3181), .B(w3182), .Z(w3183) );
	AND U2734 ( .A(w3125), .B(w3061), .Z(w3184) );
	XOR U2735 ( .A(w3184), .B(w3183), .Z(w3185) );
	AND U2736 ( .A(w3127), .B(w3060), .Z(w3186) );
	XOR U2737 ( .A(w3186), .B(w3183), .Z(w3187) );
	XOR U2738 ( .A(w3132), .B(w3134), .Z(w3188) );
	XOR U2739 ( .A(w3059), .B(w3058), .Z(w3189) );
	AND U2740 ( .A(w3188), .B(w3189), .Z(w3190) );
	AND U2741 ( .A(w3132), .B(w3059), .Z(w3191) );
	XOR U2742 ( .A(w3191), .B(w3190), .Z(w3192) );
	AND U2743 ( .A(w3134), .B(w3058), .Z(w3193) );
	XOR U2744 ( .A(w3193), .B(w3190), .Z(w3194) );
	XOR U2745 ( .A(w3187), .B(w3180), .Z(w3195) );
	XOR U2746 ( .A(w3185), .B(w3179), .Z(w3196) );
	XOR U2747 ( .A(w3194), .B(w3180), .Z(w3197) );
	XOR U2748 ( .A(w3192), .B(w3179), .Z(w3198) );
	XOR U2749 ( .A(w3201), .B(w3197), .Z(w3207) );
	XOR U2750 ( .A(w3202), .B(w3197), .Z(w3208) );
	XOR U2751 ( .A(w3206), .B(w3197), .Z(w3209) );
	XOR U2752 ( .A(w3199), .B(w3198), .Z(w3210) );
	XOR U2753 ( .A(w3208), .B(w3198), .Z(w3211) );
	XOR U2754 ( .A(w3203), .B(w3198), .Z(w3212) );
	XOR U2755 ( .A(w3204), .B(w3198), .Z(w3213) );
	XOR U2756 ( .A(w3205), .B(w3198), .Z(w3214) );
	XOR U2757 ( .A(w3210), .B(w3195), .Z(w3215) );
	XOR U2758 ( .A(w3207), .B(w3195), .Z(w3216) );
	XOR U2759 ( .A(w3215), .B(w3196), .Z(w3217) );
	XOR U2760 ( .A(w3200), .B(w3196), .Z(w3218) );
	XOR U2761 ( .A(w3211), .B(w3196), .Z(w3219) );
	XOR U2762 ( .A(w3213), .B(w3196), .Z(w3220) );
	XOR U2763 ( .A(w3214), .B(w3196), .Z(w3221) );
	XOR U2764 ( .A(w3209), .B(w3196), .Z(w3222) );
	XOR U2765 ( .A(w3218), .B(w3165), .Z(w3223) );
	XOR U2766 ( .A(w3212), .B(w3165), .Z(w3224) );
	XOR U2767 ( .A(w3216), .B(w3166), .Z(w3225) );
	XOR U2768 ( .A(w3217), .B(w3163), .Z(w3226) );
	XOR U2769 ( .A(w3224), .B(w3163), .Z(w3227) );
	XOR U2770 ( .A(w3221), .B(w3163), .Z(w3228) );
	XOR U2771 ( .A(w3226), .B(w3164), .Z(w3229) );
	XOR U2772 ( .A(w3223), .B(w3164), .Z(w3230) );
	XOR U2773 ( .A(w3227), .B(w3164), .Z(w3231) );
	XOR U2774 ( .A(w3228), .B(w3164), .Z(w3232) );
	XOR U2775 ( .A(w3236), .B(w120), .Z(w3241) );
	XOR U2776 ( .A(w3237), .B(w120), .Z(w3242) );
	XOR U2777 ( .A(w3240), .B(w120), .Z(w3243) );
	XOR U2778 ( .A(w3233), .B(w121), .Z(w3244) );
	XOR U2779 ( .A(w3234), .B(w121), .Z(w3245) );
	XOR U2780 ( .A(w3242), .B(w121), .Z(w3246) );
	XOR U2781 ( .A(w3238), .B(w121), .Z(w3247) );
	XOR U2782 ( .A(w3239), .B(w121), .Z(w3248) );
	XOR U2783 ( .A(w3243), .B(w121), .Z(w3249) );
	XOR U2784 ( .A(w3245), .B(w122), .Z(w3250) );
	XOR U2785 ( .A(w3246), .B(w122), .Z(w3251) );
	XOR U2786 ( .A(w3247), .B(w122), .Z(w3252) );
	XOR U2787 ( .A(w3248), .B(w122), .Z(w3253) );
	XOR U2788 ( .A(w3249), .B(w122), .Z(w3254) );
	XOR U2789 ( .A(w3241), .B(w123), .Z(w3255) );
	XOR U2790 ( .A(w3253), .B(w123), .Z(w3256) );
	XOR U2791 ( .A(w3244), .B(w124), .Z(w3257) );
	XOR U2792 ( .A(w3255), .B(w124), .Z(w3258) );
	XOR U2793 ( .A(w3257), .B(w125), .Z(w3259) );
	XOR U2794 ( .A(w3254), .B(w125), .Z(w3260) );
	XOR U2795 ( .A(w3259), .B(w126), .Z(w3261) );
	XOR U2796 ( .A(w3258), .B(w126), .Z(w3262) );
	XOR U2797 ( .A(w3252), .B(w126), .Z(w3263) );
	XOR U2798 ( .A(w3260), .B(w126), .Z(w3264) );
	XOR U2799 ( .A(w3261), .B(w127), .Z(w3265) );
	XOR U2800 ( .A(w3250), .B(w127), .Z(w3266) );
	XOR U2801 ( .A(w3235), .B(w127), .Z(w3267) );
	XOR U2802 ( .A(w3262), .B(w127), .Z(w3268) );
	XOR U2803 ( .A(w3251), .B(w127), .Z(w3269) );
	XOR U2804 ( .A(w3263), .B(w127), .Z(w3270) );
	XOR U2805 ( .A(w3256), .B(w127), .Z(w3271) );
	XOR U2806 ( .A(w3264), .B(w127), .Z(w3272) );
	XOR U2807 ( .A(w3265), .B(w3269), .Z(w3273) );
	XOR U2808 ( .A(w3266), .B(w3270), .Z(w3274) );
	XOR U2809 ( .A(w3267), .B(w3271), .Z(w3275) );
	XOR U2810 ( .A(w3268), .B(w3272), .Z(w3276) );
	XOR U2811 ( .A(w3275), .B(w3273), .Z(w3277) );
	XOR U2812 ( .A(w3276), .B(w3274), .Z(w3278) );
	XOR U2813 ( .A(w3274), .B(w3273), .Z(w3279) );
	XOR U2814 ( .A(w3267), .B(w3265), .Z(w3282) );
	XOR U2815 ( .A(w3268), .B(w3266), .Z(w3283) );
	XOR U2816 ( .A(w3271), .B(w3269), .Z(w3284) );
	XOR U2817 ( .A(w3272), .B(w3270), .Z(w3285) );
	XOR U2818 ( .A(w3283), .B(w3282), .Z(w3286) );
	XOR U2819 ( .A(w3285), .B(w3284), .Z(w3287) );
	AND U2820 ( .A(w3286), .B(w3287), .Z(w3288) );
	AND U2821 ( .A(w3283), .B(w3285), .Z(w3289) );
	XOR U2822 ( .A(w3289), .B(w3288), .Z(w3290) );
	AND U2823 ( .A(w3282), .B(w3284), .Z(w3291) );
	XOR U2824 ( .A(w3291), .B(w3288), .Z(w3292) );
	XOR U2825 ( .A(w3292), .B(w3290), .Z(w3293) );
	XOR U2826 ( .A(w3268), .B(w3267), .Z(w3294) );
	XOR U2827 ( .A(w3272), .B(w3271), .Z(w3295) );
	AND U2828 ( .A(w3294), .B(w3295), .Z(w3296) );
	AND U2829 ( .A(w3268), .B(w3272), .Z(w3297) );
	XOR U2830 ( .A(w3297), .B(w3296), .Z(w3298) );
	AND U2831 ( .A(w3267), .B(w3271), .Z(w3299) );
	XOR U2832 ( .A(w3299), .B(w3296), .Z(w3300) );
	XOR U2833 ( .A(w3266), .B(w3265), .Z(w3301) );
	XOR U2834 ( .A(w3270), .B(w3269), .Z(w3302) );
	AND U2835 ( .A(w3301), .B(w3302), .Z(w3303) );
	AND U2836 ( .A(w3266), .B(w3270), .Z(w3304) );
	XOR U2837 ( .A(w3304), .B(w3303), .Z(w3305) );
	AND U2838 ( .A(w3265), .B(w3269), .Z(w3306) );
	XOR U2839 ( .A(w3306), .B(w3303), .Z(w3307) );
	XOR U2840 ( .A(w3300), .B(w3293), .Z(w3308) );
	XOR U2841 ( .A(w3298), .B(w3292), .Z(w3309) );
	XOR U2842 ( .A(w3307), .B(w3293), .Z(w3310) );
	XOR U2843 ( .A(w3305), .B(w3292), .Z(w3311) );
	XOR U2844 ( .A(w3273), .B(w3310), .Z(w3312) );
	XOR U2845 ( .A(w3279), .B(w3311), .Z(w3313) );
	XOR U2846 ( .A(w3278), .B(w3308), .Z(w3314) );
	XOR U2847 ( .A(w3277), .B(w3309), .Z(w3315) );
	XOR U2848 ( .A(w3314), .B(w3312), .Z(w3316) );
	XOR U2849 ( .A(w3315), .B(w3313), .Z(w3317) );
	XOR U2850 ( .A(w3317), .B(w3316), .Z(w3318) );
	XOR U2851 ( .A(w3315), .B(w3314), .Z(w3319) );
	XOR U2852 ( .A(w3313), .B(w3312), .Z(w3320) );
	AND U2853 ( .A(w3319), .B(w3320), .Z(w3321) );
	AND U2854 ( .A(w3315), .B(w3313), .Z(w3322) );
	XOR U2855 ( .A(w3322), .B(w3321), .Z(w3323) );
	AND U2856 ( .A(w3314), .B(w3312), .Z(w3324) );
	XOR U2857 ( .A(w3324), .B(w3321), .Z(w3325) );
	XOR U2858 ( .A(w3318), .B(w3325), .Z(w3326) );
	XOR U2859 ( .A(w3317), .B(w3323), .Z(w3327) );
	XOR U2860 ( .A(w3326), .B(w3327), .Z(w3328) );
	XOR U2861 ( .A(w3313), .B(w3312), .Z(w3329) );
	AND U2862 ( .A(w3328), .B(w3329), .Z(w3330) );
	AND U2863 ( .A(w3326), .B(w3313), .Z(w3331) );
	XOR U2864 ( .A(w3331), .B(w3330), .Z(w3332) );
	AND U2865 ( .A(w3327), .B(w3312), .Z(w3333) );
	XOR U2866 ( .A(w3333), .B(w3330), .Z(w3334) );
	XOR U2867 ( .A(w3326), .B(w3327), .Z(w3335) );
	XOR U2868 ( .A(w3315), .B(w3314), .Z(w3336) );
	AND U2869 ( .A(w3335), .B(w3336), .Z(w3337) );
	AND U2870 ( .A(w3326), .B(w3315), .Z(w3338) );
	XOR U2871 ( .A(w3338), .B(w3337), .Z(w3339) );
	AND U2872 ( .A(w3327), .B(w3314), .Z(w3340) );
	XOR U2873 ( .A(w3340), .B(w3337), .Z(w3341) );
	XOR U2874 ( .A(w3334), .B(w3341), .Z(w3344) );
	XOR U2875 ( .A(w3332), .B(w3339), .Z(w3345) );
	XOR U2876 ( .A(w3271), .B(w3269), .Z(w3346) );
	XOR U2877 ( .A(w3272), .B(w3270), .Z(w3347) );
	XOR U2878 ( .A(w3345), .B(w3344), .Z(w3348) );
	XOR U2879 ( .A(w3347), .B(w3346), .Z(w3349) );
	AND U2880 ( .A(w3348), .B(w3349), .Z(w3350) );
	AND U2881 ( .A(w3345), .B(w3347), .Z(w3351) );
	XOR U2882 ( .A(w3351), .B(w3350), .Z(w3352) );
	AND U2883 ( .A(w3344), .B(w3346), .Z(w3353) );
	XOR U2884 ( .A(w3353), .B(w3350), .Z(w3354) );
	XOR U2885 ( .A(w3354), .B(w3352), .Z(w3355) );
	XOR U2886 ( .A(w3332), .B(w3334), .Z(w3356) );
	XOR U2887 ( .A(w3272), .B(w3271), .Z(w3357) );
	AND U2888 ( .A(w3356), .B(w3357), .Z(w3358) );
	AND U2889 ( .A(w3332), .B(w3272), .Z(w3359) );
	XOR U2890 ( .A(w3359), .B(w3358), .Z(w3360) );
	AND U2891 ( .A(w3334), .B(w3271), .Z(w3361) );
	XOR U2892 ( .A(w3361), .B(w3358), .Z(w3362) );
	XOR U2893 ( .A(w3339), .B(w3341), .Z(w3363) );
	XOR U2894 ( .A(w3270), .B(w3269), .Z(w3364) );
	AND U2895 ( .A(w3363), .B(w3364), .Z(w3365) );
	AND U2896 ( .A(w3339), .B(w3270), .Z(w3366) );
	XOR U2897 ( .A(w3366), .B(w3365), .Z(w3367) );
	AND U2898 ( .A(w3341), .B(w3269), .Z(w3368) );
	XOR U2899 ( .A(w3368), .B(w3365), .Z(w3369) );
	XOR U2900 ( .A(w3362), .B(w3355), .Z(w3370) );
	XOR U2901 ( .A(w3360), .B(w3354), .Z(w3371) );
	XOR U2902 ( .A(w3369), .B(w3355), .Z(w3372) );
	XOR U2903 ( .A(w3367), .B(w3354), .Z(w3373) );
	XOR U2904 ( .A(w3334), .B(w3341), .Z(w3376) );
	XOR U2905 ( .A(w3332), .B(w3339), .Z(w3377) );
	XOR U2906 ( .A(w3267), .B(w3265), .Z(w3378) );
	XOR U2907 ( .A(w3268), .B(w3266), .Z(w3379) );
	XOR U2908 ( .A(w3377), .B(w3376), .Z(w3380) );
	XOR U2909 ( .A(w3379), .B(w3378), .Z(w3381) );
	AND U2910 ( .A(w3380), .B(w3381), .Z(w3382) );
	AND U2911 ( .A(w3377), .B(w3379), .Z(w3383) );
	XOR U2912 ( .A(w3383), .B(w3382), .Z(w3384) );
	AND U2913 ( .A(w3376), .B(w3378), .Z(w3385) );
	XOR U2914 ( .A(w3385), .B(w3382), .Z(w3386) );
	XOR U2915 ( .A(w3386), .B(w3384), .Z(w3387) );
	XOR U2916 ( .A(w3332), .B(w3334), .Z(w3388) );
	XOR U2917 ( .A(w3268), .B(w3267), .Z(w3389) );
	AND U2918 ( .A(w3388), .B(w3389), .Z(w3390) );
	AND U2919 ( .A(w3332), .B(w3268), .Z(w3391) );
	XOR U2920 ( .A(w3391), .B(w3390), .Z(w3392) );
	AND U2921 ( .A(w3334), .B(w3267), .Z(w3393) );
	XOR U2922 ( .A(w3393), .B(w3390), .Z(w3394) );
	XOR U2923 ( .A(w3339), .B(w3341), .Z(w3395) );
	XOR U2924 ( .A(w3266), .B(w3265), .Z(w3396) );
	AND U2925 ( .A(w3395), .B(w3396), .Z(w3397) );
	AND U2926 ( .A(w3339), .B(w3266), .Z(w3398) );
	XOR U2927 ( .A(w3398), .B(w3397), .Z(w3399) );
	AND U2928 ( .A(w3341), .B(w3265), .Z(w3400) );
	XOR U2929 ( .A(w3400), .B(w3397), .Z(w3401) );
	XOR U2930 ( .A(w3394), .B(w3387), .Z(w3402) );
	XOR U2931 ( .A(w3392), .B(w3386), .Z(w3403) );
	XOR U2932 ( .A(w3401), .B(w3387), .Z(w3404) );
	XOR U2933 ( .A(w3399), .B(w3386), .Z(w3405) );
	XOR U2934 ( .A(w3408), .B(w3404), .Z(w3414) );
	XOR U2935 ( .A(w3409), .B(w3404), .Z(w3415) );
	XOR U2936 ( .A(w3413), .B(w3404), .Z(w3416) );
	XOR U2937 ( .A(w3406), .B(w3405), .Z(w3417) );
	XOR U2938 ( .A(w3415), .B(w3405), .Z(w3418) );
	XOR U2939 ( .A(w3410), .B(w3405), .Z(w3419) );
	XOR U2940 ( .A(w3411), .B(w3405), .Z(w3420) );
	XOR U2941 ( .A(w3412), .B(w3405), .Z(w3421) );
	XOR U2942 ( .A(w3417), .B(w3402), .Z(w3422) );
	XOR U2943 ( .A(w3414), .B(w3402), .Z(w3423) );
	XOR U2944 ( .A(w3422), .B(w3403), .Z(w3424) );
	XOR U2945 ( .A(w3407), .B(w3403), .Z(w3425) );
	XOR U2946 ( .A(w3418), .B(w3403), .Z(w3426) );
	XOR U2947 ( .A(w3420), .B(w3403), .Z(w3427) );
	XOR U2948 ( .A(w3421), .B(w3403), .Z(w3428) );
	XOR U2949 ( .A(w3416), .B(w3403), .Z(w3429) );
	XOR U2950 ( .A(w3425), .B(w3372), .Z(w3430) );
	XOR U2951 ( .A(w3419), .B(w3372), .Z(w3431) );
	XOR U2952 ( .A(w3423), .B(w3373), .Z(w3432) );
	XOR U2953 ( .A(w3424), .B(w3370), .Z(w3433) );
	XOR U2954 ( .A(w3431), .B(w3370), .Z(w3434) );
	XOR U2955 ( .A(w3428), .B(w3370), .Z(w3435) );
	XOR U2956 ( .A(w3433), .B(w3371), .Z(w3436) );
	XOR U2957 ( .A(w3430), .B(w3371), .Z(w3437) );
	XOR U2958 ( .A(w3434), .B(w3371), .Z(w3438) );
	XOR U2959 ( .A(w3435), .B(w3371), .Z(w3439) );
endmodule

