
module compare_N16384_CC32 ( clk, rst, x, y, g );
  input [511:0] x;
  input [511:0] y;
  input clk, rst;
  output g;
  wire   ci, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560;

  DFF ci_reg ( .D(g), .CLK(clk), .RST(rst), .I(1'b1), .Q(ci) );
  XOR U516 ( .A(y[3]), .B(n2547), .Z(n2548) );
  XOR U517 ( .A(y[7]), .B(n2531), .Z(n2532) );
  XOR U518 ( .A(y[11]), .B(n2515), .Z(n2516) );
  XOR U519 ( .A(y[15]), .B(n2499), .Z(n2500) );
  XOR U520 ( .A(y[19]), .B(n2483), .Z(n2484) );
  XOR U521 ( .A(y[23]), .B(n2467), .Z(n2468) );
  XOR U522 ( .A(y[27]), .B(n2451), .Z(n2452) );
  XOR U523 ( .A(y[31]), .B(n2435), .Z(n2436) );
  XOR U524 ( .A(y[35]), .B(n2419), .Z(n2420) );
  XOR U525 ( .A(y[39]), .B(n2403), .Z(n2404) );
  XOR U526 ( .A(y[43]), .B(n2387), .Z(n2388) );
  XOR U527 ( .A(y[47]), .B(n2371), .Z(n2372) );
  XOR U528 ( .A(y[51]), .B(n2355), .Z(n2356) );
  XOR U529 ( .A(y[55]), .B(n2339), .Z(n2340) );
  XOR U530 ( .A(y[59]), .B(n2323), .Z(n2324) );
  XOR U531 ( .A(y[63]), .B(n2307), .Z(n2308) );
  XOR U532 ( .A(y[67]), .B(n2291), .Z(n2292) );
  XOR U533 ( .A(y[71]), .B(n2275), .Z(n2276) );
  XOR U534 ( .A(y[75]), .B(n2259), .Z(n2260) );
  XOR U535 ( .A(y[79]), .B(n2243), .Z(n2244) );
  XOR U536 ( .A(y[83]), .B(n2227), .Z(n2228) );
  XOR U537 ( .A(y[87]), .B(n2211), .Z(n2212) );
  XOR U538 ( .A(y[91]), .B(n2195), .Z(n2196) );
  XOR U539 ( .A(y[95]), .B(n2179), .Z(n2180) );
  XOR U540 ( .A(y[99]), .B(n2163), .Z(n2164) );
  XOR U541 ( .A(y[103]), .B(n2147), .Z(n2148) );
  XOR U542 ( .A(y[107]), .B(n2131), .Z(n2132) );
  XOR U543 ( .A(y[111]), .B(n2115), .Z(n2116) );
  XOR U544 ( .A(y[115]), .B(n2099), .Z(n2100) );
  XOR U545 ( .A(y[119]), .B(n2083), .Z(n2084) );
  XOR U546 ( .A(y[123]), .B(n2067), .Z(n2068) );
  XOR U547 ( .A(y[127]), .B(n2051), .Z(n2052) );
  XOR U548 ( .A(y[131]), .B(n2035), .Z(n2036) );
  XOR U549 ( .A(y[135]), .B(n2019), .Z(n2020) );
  XOR U550 ( .A(y[139]), .B(n2003), .Z(n2004) );
  XOR U551 ( .A(y[143]), .B(n1987), .Z(n1988) );
  XOR U552 ( .A(y[147]), .B(n1971), .Z(n1972) );
  XOR U553 ( .A(y[151]), .B(n1955), .Z(n1956) );
  XOR U554 ( .A(y[155]), .B(n1939), .Z(n1940) );
  XOR U555 ( .A(y[159]), .B(n1923), .Z(n1924) );
  XOR U556 ( .A(y[163]), .B(n1907), .Z(n1908) );
  XOR U557 ( .A(y[167]), .B(n1891), .Z(n1892) );
  XOR U558 ( .A(y[171]), .B(n1875), .Z(n1876) );
  XOR U559 ( .A(y[175]), .B(n1859), .Z(n1860) );
  XOR U560 ( .A(y[179]), .B(n1843), .Z(n1844) );
  XOR U561 ( .A(y[183]), .B(n1827), .Z(n1828) );
  XOR U562 ( .A(y[187]), .B(n1811), .Z(n1812) );
  XOR U563 ( .A(y[191]), .B(n1795), .Z(n1796) );
  XOR U564 ( .A(y[195]), .B(n1779), .Z(n1780) );
  XOR U565 ( .A(y[199]), .B(n1763), .Z(n1764) );
  XOR U566 ( .A(y[203]), .B(n1747), .Z(n1748) );
  XOR U567 ( .A(y[207]), .B(n1731), .Z(n1732) );
  XOR U568 ( .A(y[211]), .B(n1715), .Z(n1716) );
  XOR U569 ( .A(y[215]), .B(n1699), .Z(n1700) );
  XOR U570 ( .A(y[219]), .B(n1683), .Z(n1684) );
  XOR U571 ( .A(y[223]), .B(n1667), .Z(n1668) );
  XOR U572 ( .A(y[227]), .B(n1651), .Z(n1652) );
  XOR U573 ( .A(y[231]), .B(n1635), .Z(n1636) );
  XOR U574 ( .A(y[235]), .B(n1619), .Z(n1620) );
  XOR U575 ( .A(y[239]), .B(n1603), .Z(n1604) );
  XOR U576 ( .A(y[243]), .B(n1587), .Z(n1588) );
  XOR U577 ( .A(y[247]), .B(n1571), .Z(n1572) );
  XOR U578 ( .A(y[251]), .B(n1555), .Z(n1556) );
  XOR U579 ( .A(y[255]), .B(n1539), .Z(n1540) );
  XOR U580 ( .A(y[259]), .B(n1523), .Z(n1524) );
  XOR U581 ( .A(y[263]), .B(n1507), .Z(n1508) );
  XOR U582 ( .A(y[267]), .B(n1491), .Z(n1492) );
  XOR U583 ( .A(y[271]), .B(n1475), .Z(n1476) );
  XOR U584 ( .A(y[275]), .B(n1459), .Z(n1460) );
  XOR U585 ( .A(y[279]), .B(n1443), .Z(n1444) );
  XOR U586 ( .A(y[283]), .B(n1427), .Z(n1428) );
  XOR U587 ( .A(y[287]), .B(n1411), .Z(n1412) );
  XOR U588 ( .A(y[291]), .B(n1395), .Z(n1396) );
  XOR U589 ( .A(y[295]), .B(n1379), .Z(n1380) );
  XOR U590 ( .A(y[299]), .B(n1363), .Z(n1364) );
  XOR U591 ( .A(y[303]), .B(n1347), .Z(n1348) );
  XOR U592 ( .A(y[307]), .B(n1331), .Z(n1332) );
  XOR U593 ( .A(y[311]), .B(n1315), .Z(n1316) );
  XOR U594 ( .A(y[315]), .B(n1299), .Z(n1300) );
  XOR U595 ( .A(y[319]), .B(n1283), .Z(n1284) );
  XOR U596 ( .A(y[323]), .B(n1267), .Z(n1268) );
  XOR U597 ( .A(y[327]), .B(n1251), .Z(n1252) );
  XOR U598 ( .A(y[331]), .B(n1235), .Z(n1236) );
  XOR U599 ( .A(y[335]), .B(n1219), .Z(n1220) );
  XOR U600 ( .A(y[339]), .B(n1203), .Z(n1204) );
  XOR U601 ( .A(y[343]), .B(n1187), .Z(n1188) );
  XOR U602 ( .A(y[347]), .B(n1171), .Z(n1172) );
  XOR U603 ( .A(y[351]), .B(n1155), .Z(n1156) );
  XOR U604 ( .A(y[355]), .B(n1139), .Z(n1140) );
  XOR U605 ( .A(y[359]), .B(n1123), .Z(n1124) );
  XOR U606 ( .A(y[363]), .B(n1107), .Z(n1108) );
  XOR U607 ( .A(y[367]), .B(n1091), .Z(n1092) );
  XOR U608 ( .A(y[371]), .B(n1075), .Z(n1076) );
  XOR U609 ( .A(y[375]), .B(n1059), .Z(n1060) );
  XOR U610 ( .A(y[379]), .B(n1043), .Z(n1044) );
  XOR U611 ( .A(y[383]), .B(n1027), .Z(n1028) );
  XOR U612 ( .A(y[387]), .B(n1011), .Z(n1012) );
  XOR U613 ( .A(y[391]), .B(n995), .Z(n996) );
  XOR U614 ( .A(y[395]), .B(n979), .Z(n980) );
  XOR U615 ( .A(y[399]), .B(n963), .Z(n964) );
  XOR U616 ( .A(y[403]), .B(n947), .Z(n948) );
  XOR U617 ( .A(y[407]), .B(n931), .Z(n932) );
  XOR U618 ( .A(y[411]), .B(n915), .Z(n916) );
  XOR U619 ( .A(y[415]), .B(n899), .Z(n900) );
  XOR U620 ( .A(y[419]), .B(n883), .Z(n884) );
  XOR U621 ( .A(y[423]), .B(n867), .Z(n868) );
  XOR U622 ( .A(y[427]), .B(n851), .Z(n852) );
  XOR U623 ( .A(y[431]), .B(n835), .Z(n836) );
  XOR U624 ( .A(y[435]), .B(n819), .Z(n820) );
  XOR U625 ( .A(y[439]), .B(n803), .Z(n804) );
  XOR U626 ( .A(y[443]), .B(n787), .Z(n788) );
  XOR U627 ( .A(y[447]), .B(n771), .Z(n772) );
  XOR U628 ( .A(y[451]), .B(n755), .Z(n756) );
  XOR U629 ( .A(y[455]), .B(n739), .Z(n740) );
  XOR U630 ( .A(y[459]), .B(n723), .Z(n724) );
  XOR U631 ( .A(y[463]), .B(n707), .Z(n708) );
  XOR U632 ( .A(y[467]), .B(n691), .Z(n692) );
  XOR U633 ( .A(y[471]), .B(n675), .Z(n676) );
  XOR U634 ( .A(y[475]), .B(n659), .Z(n660) );
  XOR U635 ( .A(y[479]), .B(n643), .Z(n644) );
  XOR U636 ( .A(y[483]), .B(n627), .Z(n628) );
  XOR U637 ( .A(y[487]), .B(n611), .Z(n612) );
  XOR U638 ( .A(y[491]), .B(n595), .Z(n596) );
  XOR U639 ( .A(y[495]), .B(n579), .Z(n580) );
  XOR U640 ( .A(y[499]), .B(n563), .Z(n564) );
  XOR U641 ( .A(y[503]), .B(n547), .Z(n548) );
  XOR U642 ( .A(y[507]), .B(n531), .Z(n532) );
  XOR U643 ( .A(y[4]), .B(n2543), .Z(n2544) );
  XOR U644 ( .A(y[8]), .B(n2527), .Z(n2528) );
  XOR U645 ( .A(y[12]), .B(n2511), .Z(n2512) );
  XOR U646 ( .A(y[16]), .B(n2495), .Z(n2496) );
  XOR U647 ( .A(y[20]), .B(n2479), .Z(n2480) );
  XOR U648 ( .A(y[24]), .B(n2463), .Z(n2464) );
  XOR U649 ( .A(y[28]), .B(n2447), .Z(n2448) );
  XOR U650 ( .A(y[32]), .B(n2431), .Z(n2432) );
  XOR U651 ( .A(y[36]), .B(n2415), .Z(n2416) );
  XOR U652 ( .A(y[40]), .B(n2399), .Z(n2400) );
  XOR U653 ( .A(y[44]), .B(n2383), .Z(n2384) );
  XOR U654 ( .A(y[48]), .B(n2367), .Z(n2368) );
  XOR U655 ( .A(y[52]), .B(n2351), .Z(n2352) );
  XOR U656 ( .A(y[56]), .B(n2335), .Z(n2336) );
  XOR U657 ( .A(y[60]), .B(n2319), .Z(n2320) );
  XOR U658 ( .A(y[64]), .B(n2303), .Z(n2304) );
  XOR U659 ( .A(y[68]), .B(n2287), .Z(n2288) );
  XOR U660 ( .A(y[72]), .B(n2271), .Z(n2272) );
  XOR U661 ( .A(y[76]), .B(n2255), .Z(n2256) );
  XOR U662 ( .A(y[80]), .B(n2239), .Z(n2240) );
  XOR U663 ( .A(y[84]), .B(n2223), .Z(n2224) );
  XOR U664 ( .A(y[88]), .B(n2207), .Z(n2208) );
  XOR U665 ( .A(y[92]), .B(n2191), .Z(n2192) );
  XOR U666 ( .A(y[96]), .B(n2175), .Z(n2176) );
  XOR U667 ( .A(y[100]), .B(n2159), .Z(n2160) );
  XOR U668 ( .A(y[104]), .B(n2143), .Z(n2144) );
  XOR U669 ( .A(y[108]), .B(n2127), .Z(n2128) );
  XOR U670 ( .A(y[112]), .B(n2111), .Z(n2112) );
  XOR U671 ( .A(y[116]), .B(n2095), .Z(n2096) );
  XOR U672 ( .A(y[120]), .B(n2079), .Z(n2080) );
  XOR U673 ( .A(y[124]), .B(n2063), .Z(n2064) );
  XOR U674 ( .A(y[128]), .B(n2047), .Z(n2048) );
  XOR U675 ( .A(y[132]), .B(n2031), .Z(n2032) );
  XOR U676 ( .A(y[136]), .B(n2015), .Z(n2016) );
  XOR U677 ( .A(y[140]), .B(n1999), .Z(n2000) );
  XOR U678 ( .A(y[144]), .B(n1983), .Z(n1984) );
  XOR U679 ( .A(y[148]), .B(n1967), .Z(n1968) );
  XOR U680 ( .A(y[152]), .B(n1951), .Z(n1952) );
  XOR U681 ( .A(y[156]), .B(n1935), .Z(n1936) );
  XOR U682 ( .A(y[160]), .B(n1919), .Z(n1920) );
  XOR U683 ( .A(y[164]), .B(n1903), .Z(n1904) );
  XOR U684 ( .A(y[168]), .B(n1887), .Z(n1888) );
  XOR U685 ( .A(y[172]), .B(n1871), .Z(n1872) );
  XOR U686 ( .A(y[176]), .B(n1855), .Z(n1856) );
  XOR U687 ( .A(y[180]), .B(n1839), .Z(n1840) );
  XOR U688 ( .A(y[184]), .B(n1823), .Z(n1824) );
  XOR U689 ( .A(y[188]), .B(n1807), .Z(n1808) );
  XOR U690 ( .A(y[192]), .B(n1791), .Z(n1792) );
  XOR U691 ( .A(y[196]), .B(n1775), .Z(n1776) );
  XOR U692 ( .A(y[200]), .B(n1759), .Z(n1760) );
  XOR U693 ( .A(y[204]), .B(n1743), .Z(n1744) );
  XOR U694 ( .A(y[208]), .B(n1727), .Z(n1728) );
  XOR U695 ( .A(y[212]), .B(n1711), .Z(n1712) );
  XOR U696 ( .A(y[216]), .B(n1695), .Z(n1696) );
  XOR U697 ( .A(y[220]), .B(n1679), .Z(n1680) );
  XOR U698 ( .A(y[224]), .B(n1663), .Z(n1664) );
  XOR U699 ( .A(y[228]), .B(n1647), .Z(n1648) );
  XOR U700 ( .A(y[232]), .B(n1631), .Z(n1632) );
  XOR U701 ( .A(y[236]), .B(n1615), .Z(n1616) );
  XOR U702 ( .A(y[240]), .B(n1599), .Z(n1600) );
  XOR U703 ( .A(y[244]), .B(n1583), .Z(n1584) );
  XOR U704 ( .A(y[248]), .B(n1567), .Z(n1568) );
  XOR U705 ( .A(y[252]), .B(n1551), .Z(n1552) );
  XOR U706 ( .A(y[256]), .B(n1535), .Z(n1536) );
  XOR U707 ( .A(y[260]), .B(n1519), .Z(n1520) );
  XOR U708 ( .A(y[264]), .B(n1503), .Z(n1504) );
  XOR U709 ( .A(y[268]), .B(n1487), .Z(n1488) );
  XOR U710 ( .A(y[272]), .B(n1471), .Z(n1472) );
  XOR U711 ( .A(y[276]), .B(n1455), .Z(n1456) );
  XOR U712 ( .A(y[280]), .B(n1439), .Z(n1440) );
  XOR U713 ( .A(y[284]), .B(n1423), .Z(n1424) );
  XOR U714 ( .A(y[288]), .B(n1407), .Z(n1408) );
  XOR U715 ( .A(y[292]), .B(n1391), .Z(n1392) );
  XOR U716 ( .A(y[296]), .B(n1375), .Z(n1376) );
  XOR U717 ( .A(y[300]), .B(n1359), .Z(n1360) );
  XOR U718 ( .A(y[304]), .B(n1343), .Z(n1344) );
  XOR U719 ( .A(y[308]), .B(n1327), .Z(n1328) );
  XOR U720 ( .A(y[312]), .B(n1311), .Z(n1312) );
  XOR U721 ( .A(y[316]), .B(n1295), .Z(n1296) );
  XOR U722 ( .A(y[320]), .B(n1279), .Z(n1280) );
  XOR U723 ( .A(y[324]), .B(n1263), .Z(n1264) );
  XOR U724 ( .A(y[328]), .B(n1247), .Z(n1248) );
  XOR U725 ( .A(y[332]), .B(n1231), .Z(n1232) );
  XOR U726 ( .A(y[336]), .B(n1215), .Z(n1216) );
  XOR U727 ( .A(y[340]), .B(n1199), .Z(n1200) );
  XOR U728 ( .A(y[344]), .B(n1183), .Z(n1184) );
  XOR U729 ( .A(y[348]), .B(n1167), .Z(n1168) );
  XOR U730 ( .A(y[352]), .B(n1151), .Z(n1152) );
  XOR U731 ( .A(y[356]), .B(n1135), .Z(n1136) );
  XOR U732 ( .A(y[360]), .B(n1119), .Z(n1120) );
  XOR U733 ( .A(y[364]), .B(n1103), .Z(n1104) );
  XOR U734 ( .A(y[368]), .B(n1087), .Z(n1088) );
  XOR U735 ( .A(y[372]), .B(n1071), .Z(n1072) );
  XOR U736 ( .A(y[376]), .B(n1055), .Z(n1056) );
  XOR U737 ( .A(y[380]), .B(n1039), .Z(n1040) );
  XOR U738 ( .A(y[384]), .B(n1023), .Z(n1024) );
  XOR U739 ( .A(y[388]), .B(n1007), .Z(n1008) );
  XOR U740 ( .A(y[392]), .B(n991), .Z(n992) );
  XOR U741 ( .A(y[396]), .B(n975), .Z(n976) );
  XOR U742 ( .A(y[400]), .B(n959), .Z(n960) );
  XOR U743 ( .A(y[404]), .B(n943), .Z(n944) );
  XOR U744 ( .A(y[408]), .B(n927), .Z(n928) );
  XOR U745 ( .A(y[412]), .B(n911), .Z(n912) );
  XOR U746 ( .A(y[416]), .B(n895), .Z(n896) );
  XOR U747 ( .A(y[420]), .B(n879), .Z(n880) );
  XOR U748 ( .A(y[424]), .B(n863), .Z(n864) );
  XOR U749 ( .A(y[428]), .B(n847), .Z(n848) );
  XOR U750 ( .A(y[432]), .B(n831), .Z(n832) );
  XOR U751 ( .A(y[436]), .B(n815), .Z(n816) );
  XOR U752 ( .A(y[440]), .B(n799), .Z(n800) );
  XOR U753 ( .A(y[444]), .B(n783), .Z(n784) );
  XOR U754 ( .A(y[448]), .B(n767), .Z(n768) );
  XOR U755 ( .A(y[452]), .B(n751), .Z(n752) );
  XOR U756 ( .A(y[456]), .B(n735), .Z(n736) );
  XOR U757 ( .A(y[460]), .B(n719), .Z(n720) );
  XOR U758 ( .A(y[464]), .B(n703), .Z(n704) );
  XOR U759 ( .A(y[468]), .B(n687), .Z(n688) );
  XOR U760 ( .A(y[472]), .B(n671), .Z(n672) );
  XOR U761 ( .A(y[476]), .B(n655), .Z(n656) );
  XOR U762 ( .A(y[480]), .B(n639), .Z(n640) );
  XOR U763 ( .A(y[484]), .B(n623), .Z(n624) );
  XOR U764 ( .A(y[488]), .B(n607), .Z(n608) );
  XOR U765 ( .A(y[492]), .B(n591), .Z(n592) );
  XOR U766 ( .A(y[496]), .B(n575), .Z(n576) );
  XOR U767 ( .A(y[500]), .B(n559), .Z(n560) );
  XOR U768 ( .A(y[504]), .B(n543), .Z(n544) );
  XOR U769 ( .A(y[508]), .B(n527), .Z(n528) );
  XOR U770 ( .A(y[5]), .B(n2539), .Z(n2540) );
  XOR U771 ( .A(y[9]), .B(n2523), .Z(n2524) );
  XOR U772 ( .A(y[13]), .B(n2507), .Z(n2508) );
  XOR U773 ( .A(y[17]), .B(n2491), .Z(n2492) );
  XOR U774 ( .A(y[21]), .B(n2475), .Z(n2476) );
  XOR U775 ( .A(y[25]), .B(n2459), .Z(n2460) );
  XOR U776 ( .A(y[29]), .B(n2443), .Z(n2444) );
  XOR U777 ( .A(y[33]), .B(n2427), .Z(n2428) );
  XOR U778 ( .A(y[37]), .B(n2411), .Z(n2412) );
  XOR U779 ( .A(y[41]), .B(n2395), .Z(n2396) );
  XOR U780 ( .A(y[45]), .B(n2379), .Z(n2380) );
  XOR U781 ( .A(y[49]), .B(n2363), .Z(n2364) );
  XOR U782 ( .A(y[53]), .B(n2347), .Z(n2348) );
  XOR U783 ( .A(y[57]), .B(n2331), .Z(n2332) );
  XOR U784 ( .A(y[61]), .B(n2315), .Z(n2316) );
  XOR U785 ( .A(y[65]), .B(n2299), .Z(n2300) );
  XOR U786 ( .A(y[69]), .B(n2283), .Z(n2284) );
  XOR U787 ( .A(y[73]), .B(n2267), .Z(n2268) );
  XOR U788 ( .A(y[77]), .B(n2251), .Z(n2252) );
  XOR U789 ( .A(y[81]), .B(n2235), .Z(n2236) );
  XOR U790 ( .A(y[85]), .B(n2219), .Z(n2220) );
  XOR U791 ( .A(y[89]), .B(n2203), .Z(n2204) );
  XOR U792 ( .A(y[93]), .B(n2187), .Z(n2188) );
  XOR U793 ( .A(y[97]), .B(n2171), .Z(n2172) );
  XOR U794 ( .A(y[101]), .B(n2155), .Z(n2156) );
  XOR U795 ( .A(y[105]), .B(n2139), .Z(n2140) );
  XOR U796 ( .A(y[109]), .B(n2123), .Z(n2124) );
  XOR U797 ( .A(y[113]), .B(n2107), .Z(n2108) );
  XOR U798 ( .A(y[117]), .B(n2091), .Z(n2092) );
  XOR U799 ( .A(y[121]), .B(n2075), .Z(n2076) );
  XOR U800 ( .A(y[125]), .B(n2059), .Z(n2060) );
  XOR U801 ( .A(y[129]), .B(n2043), .Z(n2044) );
  XOR U802 ( .A(y[133]), .B(n2027), .Z(n2028) );
  XOR U803 ( .A(y[137]), .B(n2011), .Z(n2012) );
  XOR U804 ( .A(y[141]), .B(n1995), .Z(n1996) );
  XOR U805 ( .A(y[145]), .B(n1979), .Z(n1980) );
  XOR U806 ( .A(y[149]), .B(n1963), .Z(n1964) );
  XOR U807 ( .A(y[153]), .B(n1947), .Z(n1948) );
  XOR U808 ( .A(y[157]), .B(n1931), .Z(n1932) );
  XOR U809 ( .A(y[161]), .B(n1915), .Z(n1916) );
  XOR U810 ( .A(y[165]), .B(n1899), .Z(n1900) );
  XOR U811 ( .A(y[169]), .B(n1883), .Z(n1884) );
  XOR U812 ( .A(y[173]), .B(n1867), .Z(n1868) );
  XOR U813 ( .A(y[177]), .B(n1851), .Z(n1852) );
  XOR U814 ( .A(y[181]), .B(n1835), .Z(n1836) );
  XOR U815 ( .A(y[185]), .B(n1819), .Z(n1820) );
  XOR U816 ( .A(y[189]), .B(n1803), .Z(n1804) );
  XOR U817 ( .A(y[193]), .B(n1787), .Z(n1788) );
  XOR U818 ( .A(y[197]), .B(n1771), .Z(n1772) );
  XOR U819 ( .A(y[201]), .B(n1755), .Z(n1756) );
  XOR U820 ( .A(y[205]), .B(n1739), .Z(n1740) );
  XOR U821 ( .A(y[209]), .B(n1723), .Z(n1724) );
  XOR U822 ( .A(y[213]), .B(n1707), .Z(n1708) );
  XOR U823 ( .A(y[217]), .B(n1691), .Z(n1692) );
  XOR U824 ( .A(y[221]), .B(n1675), .Z(n1676) );
  XOR U825 ( .A(y[225]), .B(n1659), .Z(n1660) );
  XOR U826 ( .A(y[229]), .B(n1643), .Z(n1644) );
  XOR U827 ( .A(y[233]), .B(n1627), .Z(n1628) );
  XOR U828 ( .A(y[237]), .B(n1611), .Z(n1612) );
  XOR U829 ( .A(y[241]), .B(n1595), .Z(n1596) );
  XOR U830 ( .A(y[245]), .B(n1579), .Z(n1580) );
  XOR U831 ( .A(y[249]), .B(n1563), .Z(n1564) );
  XOR U832 ( .A(y[253]), .B(n1547), .Z(n1548) );
  XOR U833 ( .A(y[257]), .B(n1531), .Z(n1532) );
  XOR U834 ( .A(y[261]), .B(n1515), .Z(n1516) );
  XOR U835 ( .A(y[265]), .B(n1499), .Z(n1500) );
  XOR U836 ( .A(y[269]), .B(n1483), .Z(n1484) );
  XOR U837 ( .A(y[273]), .B(n1467), .Z(n1468) );
  XOR U838 ( .A(y[277]), .B(n1451), .Z(n1452) );
  XOR U839 ( .A(y[281]), .B(n1435), .Z(n1436) );
  XOR U840 ( .A(y[285]), .B(n1419), .Z(n1420) );
  XOR U841 ( .A(y[289]), .B(n1403), .Z(n1404) );
  XOR U842 ( .A(y[293]), .B(n1387), .Z(n1388) );
  XOR U843 ( .A(y[297]), .B(n1371), .Z(n1372) );
  XOR U844 ( .A(y[301]), .B(n1355), .Z(n1356) );
  XOR U845 ( .A(y[305]), .B(n1339), .Z(n1340) );
  XOR U846 ( .A(y[309]), .B(n1323), .Z(n1324) );
  XOR U847 ( .A(y[313]), .B(n1307), .Z(n1308) );
  XOR U848 ( .A(y[317]), .B(n1291), .Z(n1292) );
  XOR U849 ( .A(y[321]), .B(n1275), .Z(n1276) );
  XOR U850 ( .A(y[325]), .B(n1259), .Z(n1260) );
  XOR U851 ( .A(y[329]), .B(n1243), .Z(n1244) );
  XOR U852 ( .A(y[333]), .B(n1227), .Z(n1228) );
  XOR U853 ( .A(y[337]), .B(n1211), .Z(n1212) );
  XOR U854 ( .A(y[341]), .B(n1195), .Z(n1196) );
  XOR U855 ( .A(y[345]), .B(n1179), .Z(n1180) );
  XOR U856 ( .A(y[349]), .B(n1163), .Z(n1164) );
  XOR U857 ( .A(y[353]), .B(n1147), .Z(n1148) );
  XOR U858 ( .A(y[357]), .B(n1131), .Z(n1132) );
  XOR U859 ( .A(y[361]), .B(n1115), .Z(n1116) );
  XOR U860 ( .A(y[365]), .B(n1099), .Z(n1100) );
  XOR U861 ( .A(y[369]), .B(n1083), .Z(n1084) );
  XOR U862 ( .A(y[373]), .B(n1067), .Z(n1068) );
  XOR U863 ( .A(y[377]), .B(n1051), .Z(n1052) );
  XOR U864 ( .A(y[381]), .B(n1035), .Z(n1036) );
  XOR U865 ( .A(y[385]), .B(n1019), .Z(n1020) );
  XOR U866 ( .A(y[389]), .B(n1003), .Z(n1004) );
  XOR U867 ( .A(y[393]), .B(n987), .Z(n988) );
  XOR U868 ( .A(y[397]), .B(n971), .Z(n972) );
  XOR U869 ( .A(y[401]), .B(n955), .Z(n956) );
  XOR U870 ( .A(y[405]), .B(n939), .Z(n940) );
  XOR U871 ( .A(y[409]), .B(n923), .Z(n924) );
  XOR U872 ( .A(y[413]), .B(n907), .Z(n908) );
  XOR U873 ( .A(y[417]), .B(n891), .Z(n892) );
  XOR U874 ( .A(y[421]), .B(n875), .Z(n876) );
  XOR U875 ( .A(y[425]), .B(n859), .Z(n860) );
  XOR U876 ( .A(y[429]), .B(n843), .Z(n844) );
  XOR U877 ( .A(y[433]), .B(n827), .Z(n828) );
  XOR U878 ( .A(y[437]), .B(n811), .Z(n812) );
  XOR U879 ( .A(y[441]), .B(n795), .Z(n796) );
  XOR U880 ( .A(y[445]), .B(n779), .Z(n780) );
  XOR U881 ( .A(y[449]), .B(n763), .Z(n764) );
  XOR U882 ( .A(y[453]), .B(n747), .Z(n748) );
  XOR U883 ( .A(y[457]), .B(n731), .Z(n732) );
  XOR U884 ( .A(y[461]), .B(n715), .Z(n716) );
  XOR U885 ( .A(y[465]), .B(n699), .Z(n700) );
  XOR U886 ( .A(y[469]), .B(n683), .Z(n684) );
  XOR U887 ( .A(y[473]), .B(n667), .Z(n668) );
  XOR U888 ( .A(y[477]), .B(n651), .Z(n652) );
  XOR U889 ( .A(y[481]), .B(n635), .Z(n636) );
  XOR U890 ( .A(y[485]), .B(n619), .Z(n620) );
  XOR U891 ( .A(y[489]), .B(n603), .Z(n604) );
  XOR U892 ( .A(y[493]), .B(n587), .Z(n588) );
  XOR U893 ( .A(y[497]), .B(n571), .Z(n572) );
  XOR U894 ( .A(y[501]), .B(n555), .Z(n556) );
  XOR U895 ( .A(y[505]), .B(n539), .Z(n540) );
  XOR U896 ( .A(y[509]), .B(n523), .Z(n524) );
  XOR U897 ( .A(y[2]), .B(n2551), .Z(n2552) );
  XOR U898 ( .A(y[6]), .B(n2535), .Z(n2536) );
  XOR U899 ( .A(y[10]), .B(n2519), .Z(n2520) );
  XOR U900 ( .A(y[14]), .B(n2503), .Z(n2504) );
  XOR U901 ( .A(y[18]), .B(n2487), .Z(n2488) );
  XOR U902 ( .A(y[22]), .B(n2471), .Z(n2472) );
  XOR U903 ( .A(y[26]), .B(n2455), .Z(n2456) );
  XOR U904 ( .A(y[30]), .B(n2439), .Z(n2440) );
  XOR U905 ( .A(y[34]), .B(n2423), .Z(n2424) );
  XOR U906 ( .A(y[38]), .B(n2407), .Z(n2408) );
  XOR U907 ( .A(y[42]), .B(n2391), .Z(n2392) );
  XOR U908 ( .A(y[46]), .B(n2375), .Z(n2376) );
  XOR U909 ( .A(y[50]), .B(n2359), .Z(n2360) );
  XOR U910 ( .A(y[54]), .B(n2343), .Z(n2344) );
  XOR U911 ( .A(y[58]), .B(n2327), .Z(n2328) );
  XOR U912 ( .A(y[62]), .B(n2311), .Z(n2312) );
  XOR U913 ( .A(y[66]), .B(n2295), .Z(n2296) );
  XOR U914 ( .A(y[70]), .B(n2279), .Z(n2280) );
  XOR U915 ( .A(y[74]), .B(n2263), .Z(n2264) );
  XOR U916 ( .A(y[78]), .B(n2247), .Z(n2248) );
  XOR U917 ( .A(y[82]), .B(n2231), .Z(n2232) );
  XOR U918 ( .A(y[86]), .B(n2215), .Z(n2216) );
  XOR U919 ( .A(y[90]), .B(n2199), .Z(n2200) );
  XOR U920 ( .A(y[94]), .B(n2183), .Z(n2184) );
  XOR U921 ( .A(y[98]), .B(n2167), .Z(n2168) );
  XOR U922 ( .A(y[102]), .B(n2151), .Z(n2152) );
  XOR U923 ( .A(y[106]), .B(n2135), .Z(n2136) );
  XOR U924 ( .A(y[110]), .B(n2119), .Z(n2120) );
  XOR U925 ( .A(y[114]), .B(n2103), .Z(n2104) );
  XOR U926 ( .A(y[118]), .B(n2087), .Z(n2088) );
  XOR U927 ( .A(y[122]), .B(n2071), .Z(n2072) );
  XOR U928 ( .A(y[126]), .B(n2055), .Z(n2056) );
  XOR U929 ( .A(y[130]), .B(n2039), .Z(n2040) );
  XOR U930 ( .A(y[134]), .B(n2023), .Z(n2024) );
  XOR U931 ( .A(y[138]), .B(n2007), .Z(n2008) );
  XOR U932 ( .A(y[142]), .B(n1991), .Z(n1992) );
  XOR U933 ( .A(y[146]), .B(n1975), .Z(n1976) );
  XOR U934 ( .A(y[150]), .B(n1959), .Z(n1960) );
  XOR U935 ( .A(y[154]), .B(n1943), .Z(n1944) );
  XOR U936 ( .A(y[158]), .B(n1927), .Z(n1928) );
  XOR U937 ( .A(y[162]), .B(n1911), .Z(n1912) );
  XOR U938 ( .A(y[166]), .B(n1895), .Z(n1896) );
  XOR U939 ( .A(y[170]), .B(n1879), .Z(n1880) );
  XOR U940 ( .A(y[174]), .B(n1863), .Z(n1864) );
  XOR U941 ( .A(y[178]), .B(n1847), .Z(n1848) );
  XOR U942 ( .A(y[182]), .B(n1831), .Z(n1832) );
  XOR U943 ( .A(y[186]), .B(n1815), .Z(n1816) );
  XOR U944 ( .A(y[190]), .B(n1799), .Z(n1800) );
  XOR U945 ( .A(y[194]), .B(n1783), .Z(n1784) );
  XOR U946 ( .A(y[198]), .B(n1767), .Z(n1768) );
  XOR U947 ( .A(y[202]), .B(n1751), .Z(n1752) );
  XOR U948 ( .A(y[206]), .B(n1735), .Z(n1736) );
  XOR U949 ( .A(y[210]), .B(n1719), .Z(n1720) );
  XOR U950 ( .A(y[214]), .B(n1703), .Z(n1704) );
  XOR U951 ( .A(y[218]), .B(n1687), .Z(n1688) );
  XOR U952 ( .A(y[222]), .B(n1671), .Z(n1672) );
  XOR U953 ( .A(y[226]), .B(n1655), .Z(n1656) );
  XOR U954 ( .A(y[230]), .B(n1639), .Z(n1640) );
  XOR U955 ( .A(y[234]), .B(n1623), .Z(n1624) );
  XOR U956 ( .A(y[238]), .B(n1607), .Z(n1608) );
  XOR U957 ( .A(y[242]), .B(n1591), .Z(n1592) );
  XOR U958 ( .A(y[246]), .B(n1575), .Z(n1576) );
  XOR U959 ( .A(y[250]), .B(n1559), .Z(n1560) );
  XOR U960 ( .A(y[254]), .B(n1543), .Z(n1544) );
  XOR U961 ( .A(y[258]), .B(n1527), .Z(n1528) );
  XOR U962 ( .A(y[262]), .B(n1511), .Z(n1512) );
  XOR U963 ( .A(y[266]), .B(n1495), .Z(n1496) );
  XOR U964 ( .A(y[270]), .B(n1479), .Z(n1480) );
  XOR U965 ( .A(y[274]), .B(n1463), .Z(n1464) );
  XOR U966 ( .A(y[278]), .B(n1447), .Z(n1448) );
  XOR U967 ( .A(y[282]), .B(n1431), .Z(n1432) );
  XOR U968 ( .A(y[286]), .B(n1415), .Z(n1416) );
  XOR U969 ( .A(y[290]), .B(n1399), .Z(n1400) );
  XOR U970 ( .A(y[294]), .B(n1383), .Z(n1384) );
  XOR U971 ( .A(y[298]), .B(n1367), .Z(n1368) );
  XOR U972 ( .A(y[302]), .B(n1351), .Z(n1352) );
  XOR U973 ( .A(y[306]), .B(n1335), .Z(n1336) );
  XOR U974 ( .A(y[310]), .B(n1319), .Z(n1320) );
  XOR U975 ( .A(y[314]), .B(n1303), .Z(n1304) );
  XOR U976 ( .A(y[318]), .B(n1287), .Z(n1288) );
  XOR U977 ( .A(y[322]), .B(n1271), .Z(n1272) );
  XOR U978 ( .A(y[326]), .B(n1255), .Z(n1256) );
  XOR U979 ( .A(y[330]), .B(n1239), .Z(n1240) );
  XOR U980 ( .A(y[334]), .B(n1223), .Z(n1224) );
  XOR U981 ( .A(y[338]), .B(n1207), .Z(n1208) );
  XOR U982 ( .A(y[342]), .B(n1191), .Z(n1192) );
  XOR U983 ( .A(y[346]), .B(n1175), .Z(n1176) );
  XOR U984 ( .A(y[350]), .B(n1159), .Z(n1160) );
  XOR U985 ( .A(y[354]), .B(n1143), .Z(n1144) );
  XOR U986 ( .A(y[358]), .B(n1127), .Z(n1128) );
  XOR U987 ( .A(y[362]), .B(n1111), .Z(n1112) );
  XOR U988 ( .A(y[366]), .B(n1095), .Z(n1096) );
  XOR U989 ( .A(y[370]), .B(n1079), .Z(n1080) );
  XOR U990 ( .A(y[374]), .B(n1063), .Z(n1064) );
  XOR U991 ( .A(y[378]), .B(n1047), .Z(n1048) );
  XOR U992 ( .A(y[382]), .B(n1031), .Z(n1032) );
  XOR U993 ( .A(y[386]), .B(n1015), .Z(n1016) );
  XOR U994 ( .A(y[390]), .B(n999), .Z(n1000) );
  XOR U995 ( .A(y[394]), .B(n983), .Z(n984) );
  XOR U996 ( .A(y[398]), .B(n967), .Z(n968) );
  XOR U997 ( .A(y[402]), .B(n951), .Z(n952) );
  XOR U998 ( .A(y[406]), .B(n935), .Z(n936) );
  XOR U999 ( .A(y[410]), .B(n919), .Z(n920) );
  XOR U1000 ( .A(y[414]), .B(n903), .Z(n904) );
  XOR U1001 ( .A(y[418]), .B(n887), .Z(n888) );
  XOR U1002 ( .A(y[422]), .B(n871), .Z(n872) );
  XOR U1003 ( .A(y[426]), .B(n855), .Z(n856) );
  XOR U1004 ( .A(y[430]), .B(n839), .Z(n840) );
  XOR U1005 ( .A(y[434]), .B(n823), .Z(n824) );
  XOR U1006 ( .A(y[438]), .B(n807), .Z(n808) );
  XOR U1007 ( .A(y[442]), .B(n791), .Z(n792) );
  XOR U1008 ( .A(y[446]), .B(n775), .Z(n776) );
  XOR U1009 ( .A(y[450]), .B(n759), .Z(n760) );
  XOR U1010 ( .A(y[454]), .B(n743), .Z(n744) );
  XOR U1011 ( .A(y[458]), .B(n727), .Z(n728) );
  XOR U1012 ( .A(y[462]), .B(n711), .Z(n712) );
  XOR U1013 ( .A(y[466]), .B(n695), .Z(n696) );
  XOR U1014 ( .A(y[470]), .B(n679), .Z(n680) );
  XOR U1015 ( .A(y[474]), .B(n663), .Z(n664) );
  XOR U1016 ( .A(y[478]), .B(n647), .Z(n648) );
  XOR U1017 ( .A(y[482]), .B(n631), .Z(n632) );
  XOR U1018 ( .A(y[486]), .B(n615), .Z(n616) );
  XOR U1019 ( .A(y[490]), .B(n599), .Z(n600) );
  XOR U1020 ( .A(y[494]), .B(n583), .Z(n584) );
  XOR U1021 ( .A(y[498]), .B(n567), .Z(n568) );
  XOR U1022 ( .A(y[502]), .B(n551), .Z(n552) );
  XOR U1023 ( .A(y[506]), .B(n535), .Z(n536) );
  XOR U1024 ( .A(y[510]), .B(n519), .Z(n520) );
  XOR U1025 ( .A(n514), .B(n515), .Z(g) );
  AND U1026 ( .A(n516), .B(n517), .Z(n514) );
  XOR U1027 ( .A(x[511]), .B(n515), .Z(n517) );
  XNOR U1028 ( .A(y[511]), .B(n515), .Z(n516) );
  XNOR U1029 ( .A(n518), .B(n519), .Z(n515) );
  AND U1030 ( .A(n520), .B(n521), .Z(n518) );
  XNOR U1031 ( .A(x[510]), .B(n519), .Z(n521) );
  XOR U1032 ( .A(n522), .B(n523), .Z(n519) );
  AND U1033 ( .A(n524), .B(n525), .Z(n522) );
  XNOR U1034 ( .A(x[509]), .B(n523), .Z(n525) );
  XOR U1035 ( .A(n526), .B(n527), .Z(n523) );
  AND U1036 ( .A(n528), .B(n529), .Z(n526) );
  XNOR U1037 ( .A(x[508]), .B(n527), .Z(n529) );
  XOR U1038 ( .A(n530), .B(n531), .Z(n527) );
  AND U1039 ( .A(n532), .B(n533), .Z(n530) );
  XNOR U1040 ( .A(x[507]), .B(n531), .Z(n533) );
  XOR U1041 ( .A(n534), .B(n535), .Z(n531) );
  AND U1042 ( .A(n536), .B(n537), .Z(n534) );
  XNOR U1043 ( .A(x[506]), .B(n535), .Z(n537) );
  XOR U1044 ( .A(n538), .B(n539), .Z(n535) );
  AND U1045 ( .A(n540), .B(n541), .Z(n538) );
  XNOR U1046 ( .A(x[505]), .B(n539), .Z(n541) );
  XOR U1047 ( .A(n542), .B(n543), .Z(n539) );
  AND U1048 ( .A(n544), .B(n545), .Z(n542) );
  XNOR U1049 ( .A(x[504]), .B(n543), .Z(n545) );
  XOR U1050 ( .A(n546), .B(n547), .Z(n543) );
  AND U1051 ( .A(n548), .B(n549), .Z(n546) );
  XNOR U1052 ( .A(x[503]), .B(n547), .Z(n549) );
  XOR U1053 ( .A(n550), .B(n551), .Z(n547) );
  AND U1054 ( .A(n552), .B(n553), .Z(n550) );
  XNOR U1055 ( .A(x[502]), .B(n551), .Z(n553) );
  XOR U1056 ( .A(n554), .B(n555), .Z(n551) );
  AND U1057 ( .A(n556), .B(n557), .Z(n554) );
  XNOR U1058 ( .A(x[501]), .B(n555), .Z(n557) );
  XOR U1059 ( .A(n558), .B(n559), .Z(n555) );
  AND U1060 ( .A(n560), .B(n561), .Z(n558) );
  XNOR U1061 ( .A(x[500]), .B(n559), .Z(n561) );
  XOR U1062 ( .A(n562), .B(n563), .Z(n559) );
  AND U1063 ( .A(n564), .B(n565), .Z(n562) );
  XNOR U1064 ( .A(x[499]), .B(n563), .Z(n565) );
  XOR U1065 ( .A(n566), .B(n567), .Z(n563) );
  AND U1066 ( .A(n568), .B(n569), .Z(n566) );
  XNOR U1067 ( .A(x[498]), .B(n567), .Z(n569) );
  XOR U1068 ( .A(n570), .B(n571), .Z(n567) );
  AND U1069 ( .A(n572), .B(n573), .Z(n570) );
  XNOR U1070 ( .A(x[497]), .B(n571), .Z(n573) );
  XOR U1071 ( .A(n574), .B(n575), .Z(n571) );
  AND U1072 ( .A(n576), .B(n577), .Z(n574) );
  XNOR U1073 ( .A(x[496]), .B(n575), .Z(n577) );
  XOR U1074 ( .A(n578), .B(n579), .Z(n575) );
  AND U1075 ( .A(n580), .B(n581), .Z(n578) );
  XNOR U1076 ( .A(x[495]), .B(n579), .Z(n581) );
  XOR U1077 ( .A(n582), .B(n583), .Z(n579) );
  AND U1078 ( .A(n584), .B(n585), .Z(n582) );
  XNOR U1079 ( .A(x[494]), .B(n583), .Z(n585) );
  XOR U1080 ( .A(n586), .B(n587), .Z(n583) );
  AND U1081 ( .A(n588), .B(n589), .Z(n586) );
  XNOR U1082 ( .A(x[493]), .B(n587), .Z(n589) );
  XOR U1083 ( .A(n590), .B(n591), .Z(n587) );
  AND U1084 ( .A(n592), .B(n593), .Z(n590) );
  XNOR U1085 ( .A(x[492]), .B(n591), .Z(n593) );
  XOR U1086 ( .A(n594), .B(n595), .Z(n591) );
  AND U1087 ( .A(n596), .B(n597), .Z(n594) );
  XNOR U1088 ( .A(x[491]), .B(n595), .Z(n597) );
  XOR U1089 ( .A(n598), .B(n599), .Z(n595) );
  AND U1090 ( .A(n600), .B(n601), .Z(n598) );
  XNOR U1091 ( .A(x[490]), .B(n599), .Z(n601) );
  XOR U1092 ( .A(n602), .B(n603), .Z(n599) );
  AND U1093 ( .A(n604), .B(n605), .Z(n602) );
  XNOR U1094 ( .A(x[489]), .B(n603), .Z(n605) );
  XOR U1095 ( .A(n606), .B(n607), .Z(n603) );
  AND U1096 ( .A(n608), .B(n609), .Z(n606) );
  XNOR U1097 ( .A(x[488]), .B(n607), .Z(n609) );
  XOR U1098 ( .A(n610), .B(n611), .Z(n607) );
  AND U1099 ( .A(n612), .B(n613), .Z(n610) );
  XNOR U1100 ( .A(x[487]), .B(n611), .Z(n613) );
  XOR U1101 ( .A(n614), .B(n615), .Z(n611) );
  AND U1102 ( .A(n616), .B(n617), .Z(n614) );
  XNOR U1103 ( .A(x[486]), .B(n615), .Z(n617) );
  XOR U1104 ( .A(n618), .B(n619), .Z(n615) );
  AND U1105 ( .A(n620), .B(n621), .Z(n618) );
  XNOR U1106 ( .A(x[485]), .B(n619), .Z(n621) );
  XOR U1107 ( .A(n622), .B(n623), .Z(n619) );
  AND U1108 ( .A(n624), .B(n625), .Z(n622) );
  XNOR U1109 ( .A(x[484]), .B(n623), .Z(n625) );
  XOR U1110 ( .A(n626), .B(n627), .Z(n623) );
  AND U1111 ( .A(n628), .B(n629), .Z(n626) );
  XNOR U1112 ( .A(x[483]), .B(n627), .Z(n629) );
  XOR U1113 ( .A(n630), .B(n631), .Z(n627) );
  AND U1114 ( .A(n632), .B(n633), .Z(n630) );
  XNOR U1115 ( .A(x[482]), .B(n631), .Z(n633) );
  XOR U1116 ( .A(n634), .B(n635), .Z(n631) );
  AND U1117 ( .A(n636), .B(n637), .Z(n634) );
  XNOR U1118 ( .A(x[481]), .B(n635), .Z(n637) );
  XOR U1119 ( .A(n638), .B(n639), .Z(n635) );
  AND U1120 ( .A(n640), .B(n641), .Z(n638) );
  XNOR U1121 ( .A(x[480]), .B(n639), .Z(n641) );
  XOR U1122 ( .A(n642), .B(n643), .Z(n639) );
  AND U1123 ( .A(n644), .B(n645), .Z(n642) );
  XNOR U1124 ( .A(x[479]), .B(n643), .Z(n645) );
  XOR U1125 ( .A(n646), .B(n647), .Z(n643) );
  AND U1126 ( .A(n648), .B(n649), .Z(n646) );
  XNOR U1127 ( .A(x[478]), .B(n647), .Z(n649) );
  XOR U1128 ( .A(n650), .B(n651), .Z(n647) );
  AND U1129 ( .A(n652), .B(n653), .Z(n650) );
  XNOR U1130 ( .A(x[477]), .B(n651), .Z(n653) );
  XOR U1131 ( .A(n654), .B(n655), .Z(n651) );
  AND U1132 ( .A(n656), .B(n657), .Z(n654) );
  XNOR U1133 ( .A(x[476]), .B(n655), .Z(n657) );
  XOR U1134 ( .A(n658), .B(n659), .Z(n655) );
  AND U1135 ( .A(n660), .B(n661), .Z(n658) );
  XNOR U1136 ( .A(x[475]), .B(n659), .Z(n661) );
  XOR U1137 ( .A(n662), .B(n663), .Z(n659) );
  AND U1138 ( .A(n664), .B(n665), .Z(n662) );
  XNOR U1139 ( .A(x[474]), .B(n663), .Z(n665) );
  XOR U1140 ( .A(n666), .B(n667), .Z(n663) );
  AND U1141 ( .A(n668), .B(n669), .Z(n666) );
  XNOR U1142 ( .A(x[473]), .B(n667), .Z(n669) );
  XOR U1143 ( .A(n670), .B(n671), .Z(n667) );
  AND U1144 ( .A(n672), .B(n673), .Z(n670) );
  XNOR U1145 ( .A(x[472]), .B(n671), .Z(n673) );
  XOR U1146 ( .A(n674), .B(n675), .Z(n671) );
  AND U1147 ( .A(n676), .B(n677), .Z(n674) );
  XNOR U1148 ( .A(x[471]), .B(n675), .Z(n677) );
  XOR U1149 ( .A(n678), .B(n679), .Z(n675) );
  AND U1150 ( .A(n680), .B(n681), .Z(n678) );
  XNOR U1151 ( .A(x[470]), .B(n679), .Z(n681) );
  XOR U1152 ( .A(n682), .B(n683), .Z(n679) );
  AND U1153 ( .A(n684), .B(n685), .Z(n682) );
  XNOR U1154 ( .A(x[469]), .B(n683), .Z(n685) );
  XOR U1155 ( .A(n686), .B(n687), .Z(n683) );
  AND U1156 ( .A(n688), .B(n689), .Z(n686) );
  XNOR U1157 ( .A(x[468]), .B(n687), .Z(n689) );
  XOR U1158 ( .A(n690), .B(n691), .Z(n687) );
  AND U1159 ( .A(n692), .B(n693), .Z(n690) );
  XNOR U1160 ( .A(x[467]), .B(n691), .Z(n693) );
  XOR U1161 ( .A(n694), .B(n695), .Z(n691) );
  AND U1162 ( .A(n696), .B(n697), .Z(n694) );
  XNOR U1163 ( .A(x[466]), .B(n695), .Z(n697) );
  XOR U1164 ( .A(n698), .B(n699), .Z(n695) );
  AND U1165 ( .A(n700), .B(n701), .Z(n698) );
  XNOR U1166 ( .A(x[465]), .B(n699), .Z(n701) );
  XOR U1167 ( .A(n702), .B(n703), .Z(n699) );
  AND U1168 ( .A(n704), .B(n705), .Z(n702) );
  XNOR U1169 ( .A(x[464]), .B(n703), .Z(n705) );
  XOR U1170 ( .A(n706), .B(n707), .Z(n703) );
  AND U1171 ( .A(n708), .B(n709), .Z(n706) );
  XNOR U1172 ( .A(x[463]), .B(n707), .Z(n709) );
  XOR U1173 ( .A(n710), .B(n711), .Z(n707) );
  AND U1174 ( .A(n712), .B(n713), .Z(n710) );
  XNOR U1175 ( .A(x[462]), .B(n711), .Z(n713) );
  XOR U1176 ( .A(n714), .B(n715), .Z(n711) );
  AND U1177 ( .A(n716), .B(n717), .Z(n714) );
  XNOR U1178 ( .A(x[461]), .B(n715), .Z(n717) );
  XOR U1179 ( .A(n718), .B(n719), .Z(n715) );
  AND U1180 ( .A(n720), .B(n721), .Z(n718) );
  XNOR U1181 ( .A(x[460]), .B(n719), .Z(n721) );
  XOR U1182 ( .A(n722), .B(n723), .Z(n719) );
  AND U1183 ( .A(n724), .B(n725), .Z(n722) );
  XNOR U1184 ( .A(x[459]), .B(n723), .Z(n725) );
  XOR U1185 ( .A(n726), .B(n727), .Z(n723) );
  AND U1186 ( .A(n728), .B(n729), .Z(n726) );
  XNOR U1187 ( .A(x[458]), .B(n727), .Z(n729) );
  XOR U1188 ( .A(n730), .B(n731), .Z(n727) );
  AND U1189 ( .A(n732), .B(n733), .Z(n730) );
  XNOR U1190 ( .A(x[457]), .B(n731), .Z(n733) );
  XOR U1191 ( .A(n734), .B(n735), .Z(n731) );
  AND U1192 ( .A(n736), .B(n737), .Z(n734) );
  XNOR U1193 ( .A(x[456]), .B(n735), .Z(n737) );
  XOR U1194 ( .A(n738), .B(n739), .Z(n735) );
  AND U1195 ( .A(n740), .B(n741), .Z(n738) );
  XNOR U1196 ( .A(x[455]), .B(n739), .Z(n741) );
  XOR U1197 ( .A(n742), .B(n743), .Z(n739) );
  AND U1198 ( .A(n744), .B(n745), .Z(n742) );
  XNOR U1199 ( .A(x[454]), .B(n743), .Z(n745) );
  XOR U1200 ( .A(n746), .B(n747), .Z(n743) );
  AND U1201 ( .A(n748), .B(n749), .Z(n746) );
  XNOR U1202 ( .A(x[453]), .B(n747), .Z(n749) );
  XOR U1203 ( .A(n750), .B(n751), .Z(n747) );
  AND U1204 ( .A(n752), .B(n753), .Z(n750) );
  XNOR U1205 ( .A(x[452]), .B(n751), .Z(n753) );
  XOR U1206 ( .A(n754), .B(n755), .Z(n751) );
  AND U1207 ( .A(n756), .B(n757), .Z(n754) );
  XNOR U1208 ( .A(x[451]), .B(n755), .Z(n757) );
  XOR U1209 ( .A(n758), .B(n759), .Z(n755) );
  AND U1210 ( .A(n760), .B(n761), .Z(n758) );
  XNOR U1211 ( .A(x[450]), .B(n759), .Z(n761) );
  XOR U1212 ( .A(n762), .B(n763), .Z(n759) );
  AND U1213 ( .A(n764), .B(n765), .Z(n762) );
  XNOR U1214 ( .A(x[449]), .B(n763), .Z(n765) );
  XOR U1215 ( .A(n766), .B(n767), .Z(n763) );
  AND U1216 ( .A(n768), .B(n769), .Z(n766) );
  XNOR U1217 ( .A(x[448]), .B(n767), .Z(n769) );
  XOR U1218 ( .A(n770), .B(n771), .Z(n767) );
  AND U1219 ( .A(n772), .B(n773), .Z(n770) );
  XNOR U1220 ( .A(x[447]), .B(n771), .Z(n773) );
  XOR U1221 ( .A(n774), .B(n775), .Z(n771) );
  AND U1222 ( .A(n776), .B(n777), .Z(n774) );
  XNOR U1223 ( .A(x[446]), .B(n775), .Z(n777) );
  XOR U1224 ( .A(n778), .B(n779), .Z(n775) );
  AND U1225 ( .A(n780), .B(n781), .Z(n778) );
  XNOR U1226 ( .A(x[445]), .B(n779), .Z(n781) );
  XOR U1227 ( .A(n782), .B(n783), .Z(n779) );
  AND U1228 ( .A(n784), .B(n785), .Z(n782) );
  XNOR U1229 ( .A(x[444]), .B(n783), .Z(n785) );
  XOR U1230 ( .A(n786), .B(n787), .Z(n783) );
  AND U1231 ( .A(n788), .B(n789), .Z(n786) );
  XNOR U1232 ( .A(x[443]), .B(n787), .Z(n789) );
  XOR U1233 ( .A(n790), .B(n791), .Z(n787) );
  AND U1234 ( .A(n792), .B(n793), .Z(n790) );
  XNOR U1235 ( .A(x[442]), .B(n791), .Z(n793) );
  XOR U1236 ( .A(n794), .B(n795), .Z(n791) );
  AND U1237 ( .A(n796), .B(n797), .Z(n794) );
  XNOR U1238 ( .A(x[441]), .B(n795), .Z(n797) );
  XOR U1239 ( .A(n798), .B(n799), .Z(n795) );
  AND U1240 ( .A(n800), .B(n801), .Z(n798) );
  XNOR U1241 ( .A(x[440]), .B(n799), .Z(n801) );
  XOR U1242 ( .A(n802), .B(n803), .Z(n799) );
  AND U1243 ( .A(n804), .B(n805), .Z(n802) );
  XNOR U1244 ( .A(x[439]), .B(n803), .Z(n805) );
  XOR U1245 ( .A(n806), .B(n807), .Z(n803) );
  AND U1246 ( .A(n808), .B(n809), .Z(n806) );
  XNOR U1247 ( .A(x[438]), .B(n807), .Z(n809) );
  XOR U1248 ( .A(n810), .B(n811), .Z(n807) );
  AND U1249 ( .A(n812), .B(n813), .Z(n810) );
  XNOR U1250 ( .A(x[437]), .B(n811), .Z(n813) );
  XOR U1251 ( .A(n814), .B(n815), .Z(n811) );
  AND U1252 ( .A(n816), .B(n817), .Z(n814) );
  XNOR U1253 ( .A(x[436]), .B(n815), .Z(n817) );
  XOR U1254 ( .A(n818), .B(n819), .Z(n815) );
  AND U1255 ( .A(n820), .B(n821), .Z(n818) );
  XNOR U1256 ( .A(x[435]), .B(n819), .Z(n821) );
  XOR U1257 ( .A(n822), .B(n823), .Z(n819) );
  AND U1258 ( .A(n824), .B(n825), .Z(n822) );
  XNOR U1259 ( .A(x[434]), .B(n823), .Z(n825) );
  XOR U1260 ( .A(n826), .B(n827), .Z(n823) );
  AND U1261 ( .A(n828), .B(n829), .Z(n826) );
  XNOR U1262 ( .A(x[433]), .B(n827), .Z(n829) );
  XOR U1263 ( .A(n830), .B(n831), .Z(n827) );
  AND U1264 ( .A(n832), .B(n833), .Z(n830) );
  XNOR U1265 ( .A(x[432]), .B(n831), .Z(n833) );
  XOR U1266 ( .A(n834), .B(n835), .Z(n831) );
  AND U1267 ( .A(n836), .B(n837), .Z(n834) );
  XNOR U1268 ( .A(x[431]), .B(n835), .Z(n837) );
  XOR U1269 ( .A(n838), .B(n839), .Z(n835) );
  AND U1270 ( .A(n840), .B(n841), .Z(n838) );
  XNOR U1271 ( .A(x[430]), .B(n839), .Z(n841) );
  XOR U1272 ( .A(n842), .B(n843), .Z(n839) );
  AND U1273 ( .A(n844), .B(n845), .Z(n842) );
  XNOR U1274 ( .A(x[429]), .B(n843), .Z(n845) );
  XOR U1275 ( .A(n846), .B(n847), .Z(n843) );
  AND U1276 ( .A(n848), .B(n849), .Z(n846) );
  XNOR U1277 ( .A(x[428]), .B(n847), .Z(n849) );
  XOR U1278 ( .A(n850), .B(n851), .Z(n847) );
  AND U1279 ( .A(n852), .B(n853), .Z(n850) );
  XNOR U1280 ( .A(x[427]), .B(n851), .Z(n853) );
  XOR U1281 ( .A(n854), .B(n855), .Z(n851) );
  AND U1282 ( .A(n856), .B(n857), .Z(n854) );
  XNOR U1283 ( .A(x[426]), .B(n855), .Z(n857) );
  XOR U1284 ( .A(n858), .B(n859), .Z(n855) );
  AND U1285 ( .A(n860), .B(n861), .Z(n858) );
  XNOR U1286 ( .A(x[425]), .B(n859), .Z(n861) );
  XOR U1287 ( .A(n862), .B(n863), .Z(n859) );
  AND U1288 ( .A(n864), .B(n865), .Z(n862) );
  XNOR U1289 ( .A(x[424]), .B(n863), .Z(n865) );
  XOR U1290 ( .A(n866), .B(n867), .Z(n863) );
  AND U1291 ( .A(n868), .B(n869), .Z(n866) );
  XNOR U1292 ( .A(x[423]), .B(n867), .Z(n869) );
  XOR U1293 ( .A(n870), .B(n871), .Z(n867) );
  AND U1294 ( .A(n872), .B(n873), .Z(n870) );
  XNOR U1295 ( .A(x[422]), .B(n871), .Z(n873) );
  XOR U1296 ( .A(n874), .B(n875), .Z(n871) );
  AND U1297 ( .A(n876), .B(n877), .Z(n874) );
  XNOR U1298 ( .A(x[421]), .B(n875), .Z(n877) );
  XOR U1299 ( .A(n878), .B(n879), .Z(n875) );
  AND U1300 ( .A(n880), .B(n881), .Z(n878) );
  XNOR U1301 ( .A(x[420]), .B(n879), .Z(n881) );
  XOR U1302 ( .A(n882), .B(n883), .Z(n879) );
  AND U1303 ( .A(n884), .B(n885), .Z(n882) );
  XNOR U1304 ( .A(x[419]), .B(n883), .Z(n885) );
  XOR U1305 ( .A(n886), .B(n887), .Z(n883) );
  AND U1306 ( .A(n888), .B(n889), .Z(n886) );
  XNOR U1307 ( .A(x[418]), .B(n887), .Z(n889) );
  XOR U1308 ( .A(n890), .B(n891), .Z(n887) );
  AND U1309 ( .A(n892), .B(n893), .Z(n890) );
  XNOR U1310 ( .A(x[417]), .B(n891), .Z(n893) );
  XOR U1311 ( .A(n894), .B(n895), .Z(n891) );
  AND U1312 ( .A(n896), .B(n897), .Z(n894) );
  XNOR U1313 ( .A(x[416]), .B(n895), .Z(n897) );
  XOR U1314 ( .A(n898), .B(n899), .Z(n895) );
  AND U1315 ( .A(n900), .B(n901), .Z(n898) );
  XNOR U1316 ( .A(x[415]), .B(n899), .Z(n901) );
  XOR U1317 ( .A(n902), .B(n903), .Z(n899) );
  AND U1318 ( .A(n904), .B(n905), .Z(n902) );
  XNOR U1319 ( .A(x[414]), .B(n903), .Z(n905) );
  XOR U1320 ( .A(n906), .B(n907), .Z(n903) );
  AND U1321 ( .A(n908), .B(n909), .Z(n906) );
  XNOR U1322 ( .A(x[413]), .B(n907), .Z(n909) );
  XOR U1323 ( .A(n910), .B(n911), .Z(n907) );
  AND U1324 ( .A(n912), .B(n913), .Z(n910) );
  XNOR U1325 ( .A(x[412]), .B(n911), .Z(n913) );
  XOR U1326 ( .A(n914), .B(n915), .Z(n911) );
  AND U1327 ( .A(n916), .B(n917), .Z(n914) );
  XNOR U1328 ( .A(x[411]), .B(n915), .Z(n917) );
  XOR U1329 ( .A(n918), .B(n919), .Z(n915) );
  AND U1330 ( .A(n920), .B(n921), .Z(n918) );
  XNOR U1331 ( .A(x[410]), .B(n919), .Z(n921) );
  XOR U1332 ( .A(n922), .B(n923), .Z(n919) );
  AND U1333 ( .A(n924), .B(n925), .Z(n922) );
  XNOR U1334 ( .A(x[409]), .B(n923), .Z(n925) );
  XOR U1335 ( .A(n926), .B(n927), .Z(n923) );
  AND U1336 ( .A(n928), .B(n929), .Z(n926) );
  XNOR U1337 ( .A(x[408]), .B(n927), .Z(n929) );
  XOR U1338 ( .A(n930), .B(n931), .Z(n927) );
  AND U1339 ( .A(n932), .B(n933), .Z(n930) );
  XNOR U1340 ( .A(x[407]), .B(n931), .Z(n933) );
  XOR U1341 ( .A(n934), .B(n935), .Z(n931) );
  AND U1342 ( .A(n936), .B(n937), .Z(n934) );
  XNOR U1343 ( .A(x[406]), .B(n935), .Z(n937) );
  XOR U1344 ( .A(n938), .B(n939), .Z(n935) );
  AND U1345 ( .A(n940), .B(n941), .Z(n938) );
  XNOR U1346 ( .A(x[405]), .B(n939), .Z(n941) );
  XOR U1347 ( .A(n942), .B(n943), .Z(n939) );
  AND U1348 ( .A(n944), .B(n945), .Z(n942) );
  XNOR U1349 ( .A(x[404]), .B(n943), .Z(n945) );
  XOR U1350 ( .A(n946), .B(n947), .Z(n943) );
  AND U1351 ( .A(n948), .B(n949), .Z(n946) );
  XNOR U1352 ( .A(x[403]), .B(n947), .Z(n949) );
  XOR U1353 ( .A(n950), .B(n951), .Z(n947) );
  AND U1354 ( .A(n952), .B(n953), .Z(n950) );
  XNOR U1355 ( .A(x[402]), .B(n951), .Z(n953) );
  XOR U1356 ( .A(n954), .B(n955), .Z(n951) );
  AND U1357 ( .A(n956), .B(n957), .Z(n954) );
  XNOR U1358 ( .A(x[401]), .B(n955), .Z(n957) );
  XOR U1359 ( .A(n958), .B(n959), .Z(n955) );
  AND U1360 ( .A(n960), .B(n961), .Z(n958) );
  XNOR U1361 ( .A(x[400]), .B(n959), .Z(n961) );
  XOR U1362 ( .A(n962), .B(n963), .Z(n959) );
  AND U1363 ( .A(n964), .B(n965), .Z(n962) );
  XNOR U1364 ( .A(x[399]), .B(n963), .Z(n965) );
  XOR U1365 ( .A(n966), .B(n967), .Z(n963) );
  AND U1366 ( .A(n968), .B(n969), .Z(n966) );
  XNOR U1367 ( .A(x[398]), .B(n967), .Z(n969) );
  XOR U1368 ( .A(n970), .B(n971), .Z(n967) );
  AND U1369 ( .A(n972), .B(n973), .Z(n970) );
  XNOR U1370 ( .A(x[397]), .B(n971), .Z(n973) );
  XOR U1371 ( .A(n974), .B(n975), .Z(n971) );
  AND U1372 ( .A(n976), .B(n977), .Z(n974) );
  XNOR U1373 ( .A(x[396]), .B(n975), .Z(n977) );
  XOR U1374 ( .A(n978), .B(n979), .Z(n975) );
  AND U1375 ( .A(n980), .B(n981), .Z(n978) );
  XNOR U1376 ( .A(x[395]), .B(n979), .Z(n981) );
  XOR U1377 ( .A(n982), .B(n983), .Z(n979) );
  AND U1378 ( .A(n984), .B(n985), .Z(n982) );
  XNOR U1379 ( .A(x[394]), .B(n983), .Z(n985) );
  XOR U1380 ( .A(n986), .B(n987), .Z(n983) );
  AND U1381 ( .A(n988), .B(n989), .Z(n986) );
  XNOR U1382 ( .A(x[393]), .B(n987), .Z(n989) );
  XOR U1383 ( .A(n990), .B(n991), .Z(n987) );
  AND U1384 ( .A(n992), .B(n993), .Z(n990) );
  XNOR U1385 ( .A(x[392]), .B(n991), .Z(n993) );
  XOR U1386 ( .A(n994), .B(n995), .Z(n991) );
  AND U1387 ( .A(n996), .B(n997), .Z(n994) );
  XNOR U1388 ( .A(x[391]), .B(n995), .Z(n997) );
  XOR U1389 ( .A(n998), .B(n999), .Z(n995) );
  AND U1390 ( .A(n1000), .B(n1001), .Z(n998) );
  XNOR U1391 ( .A(x[390]), .B(n999), .Z(n1001) );
  XOR U1392 ( .A(n1002), .B(n1003), .Z(n999) );
  AND U1393 ( .A(n1004), .B(n1005), .Z(n1002) );
  XNOR U1394 ( .A(x[389]), .B(n1003), .Z(n1005) );
  XOR U1395 ( .A(n1006), .B(n1007), .Z(n1003) );
  AND U1396 ( .A(n1008), .B(n1009), .Z(n1006) );
  XNOR U1397 ( .A(x[388]), .B(n1007), .Z(n1009) );
  XOR U1398 ( .A(n1010), .B(n1011), .Z(n1007) );
  AND U1399 ( .A(n1012), .B(n1013), .Z(n1010) );
  XNOR U1400 ( .A(x[387]), .B(n1011), .Z(n1013) );
  XOR U1401 ( .A(n1014), .B(n1015), .Z(n1011) );
  AND U1402 ( .A(n1016), .B(n1017), .Z(n1014) );
  XNOR U1403 ( .A(x[386]), .B(n1015), .Z(n1017) );
  XOR U1404 ( .A(n1018), .B(n1019), .Z(n1015) );
  AND U1405 ( .A(n1020), .B(n1021), .Z(n1018) );
  XNOR U1406 ( .A(x[385]), .B(n1019), .Z(n1021) );
  XOR U1407 ( .A(n1022), .B(n1023), .Z(n1019) );
  AND U1408 ( .A(n1024), .B(n1025), .Z(n1022) );
  XNOR U1409 ( .A(x[384]), .B(n1023), .Z(n1025) );
  XOR U1410 ( .A(n1026), .B(n1027), .Z(n1023) );
  AND U1411 ( .A(n1028), .B(n1029), .Z(n1026) );
  XNOR U1412 ( .A(x[383]), .B(n1027), .Z(n1029) );
  XOR U1413 ( .A(n1030), .B(n1031), .Z(n1027) );
  AND U1414 ( .A(n1032), .B(n1033), .Z(n1030) );
  XNOR U1415 ( .A(x[382]), .B(n1031), .Z(n1033) );
  XOR U1416 ( .A(n1034), .B(n1035), .Z(n1031) );
  AND U1417 ( .A(n1036), .B(n1037), .Z(n1034) );
  XNOR U1418 ( .A(x[381]), .B(n1035), .Z(n1037) );
  XOR U1419 ( .A(n1038), .B(n1039), .Z(n1035) );
  AND U1420 ( .A(n1040), .B(n1041), .Z(n1038) );
  XNOR U1421 ( .A(x[380]), .B(n1039), .Z(n1041) );
  XOR U1422 ( .A(n1042), .B(n1043), .Z(n1039) );
  AND U1423 ( .A(n1044), .B(n1045), .Z(n1042) );
  XNOR U1424 ( .A(x[379]), .B(n1043), .Z(n1045) );
  XOR U1425 ( .A(n1046), .B(n1047), .Z(n1043) );
  AND U1426 ( .A(n1048), .B(n1049), .Z(n1046) );
  XNOR U1427 ( .A(x[378]), .B(n1047), .Z(n1049) );
  XOR U1428 ( .A(n1050), .B(n1051), .Z(n1047) );
  AND U1429 ( .A(n1052), .B(n1053), .Z(n1050) );
  XNOR U1430 ( .A(x[377]), .B(n1051), .Z(n1053) );
  XOR U1431 ( .A(n1054), .B(n1055), .Z(n1051) );
  AND U1432 ( .A(n1056), .B(n1057), .Z(n1054) );
  XNOR U1433 ( .A(x[376]), .B(n1055), .Z(n1057) );
  XOR U1434 ( .A(n1058), .B(n1059), .Z(n1055) );
  AND U1435 ( .A(n1060), .B(n1061), .Z(n1058) );
  XNOR U1436 ( .A(x[375]), .B(n1059), .Z(n1061) );
  XOR U1437 ( .A(n1062), .B(n1063), .Z(n1059) );
  AND U1438 ( .A(n1064), .B(n1065), .Z(n1062) );
  XNOR U1439 ( .A(x[374]), .B(n1063), .Z(n1065) );
  XOR U1440 ( .A(n1066), .B(n1067), .Z(n1063) );
  AND U1441 ( .A(n1068), .B(n1069), .Z(n1066) );
  XNOR U1442 ( .A(x[373]), .B(n1067), .Z(n1069) );
  XOR U1443 ( .A(n1070), .B(n1071), .Z(n1067) );
  AND U1444 ( .A(n1072), .B(n1073), .Z(n1070) );
  XNOR U1445 ( .A(x[372]), .B(n1071), .Z(n1073) );
  XOR U1446 ( .A(n1074), .B(n1075), .Z(n1071) );
  AND U1447 ( .A(n1076), .B(n1077), .Z(n1074) );
  XNOR U1448 ( .A(x[371]), .B(n1075), .Z(n1077) );
  XOR U1449 ( .A(n1078), .B(n1079), .Z(n1075) );
  AND U1450 ( .A(n1080), .B(n1081), .Z(n1078) );
  XNOR U1451 ( .A(x[370]), .B(n1079), .Z(n1081) );
  XOR U1452 ( .A(n1082), .B(n1083), .Z(n1079) );
  AND U1453 ( .A(n1084), .B(n1085), .Z(n1082) );
  XNOR U1454 ( .A(x[369]), .B(n1083), .Z(n1085) );
  XOR U1455 ( .A(n1086), .B(n1087), .Z(n1083) );
  AND U1456 ( .A(n1088), .B(n1089), .Z(n1086) );
  XNOR U1457 ( .A(x[368]), .B(n1087), .Z(n1089) );
  XOR U1458 ( .A(n1090), .B(n1091), .Z(n1087) );
  AND U1459 ( .A(n1092), .B(n1093), .Z(n1090) );
  XNOR U1460 ( .A(x[367]), .B(n1091), .Z(n1093) );
  XOR U1461 ( .A(n1094), .B(n1095), .Z(n1091) );
  AND U1462 ( .A(n1096), .B(n1097), .Z(n1094) );
  XNOR U1463 ( .A(x[366]), .B(n1095), .Z(n1097) );
  XOR U1464 ( .A(n1098), .B(n1099), .Z(n1095) );
  AND U1465 ( .A(n1100), .B(n1101), .Z(n1098) );
  XNOR U1466 ( .A(x[365]), .B(n1099), .Z(n1101) );
  XOR U1467 ( .A(n1102), .B(n1103), .Z(n1099) );
  AND U1468 ( .A(n1104), .B(n1105), .Z(n1102) );
  XNOR U1469 ( .A(x[364]), .B(n1103), .Z(n1105) );
  XOR U1470 ( .A(n1106), .B(n1107), .Z(n1103) );
  AND U1471 ( .A(n1108), .B(n1109), .Z(n1106) );
  XNOR U1472 ( .A(x[363]), .B(n1107), .Z(n1109) );
  XOR U1473 ( .A(n1110), .B(n1111), .Z(n1107) );
  AND U1474 ( .A(n1112), .B(n1113), .Z(n1110) );
  XNOR U1475 ( .A(x[362]), .B(n1111), .Z(n1113) );
  XOR U1476 ( .A(n1114), .B(n1115), .Z(n1111) );
  AND U1477 ( .A(n1116), .B(n1117), .Z(n1114) );
  XNOR U1478 ( .A(x[361]), .B(n1115), .Z(n1117) );
  XOR U1479 ( .A(n1118), .B(n1119), .Z(n1115) );
  AND U1480 ( .A(n1120), .B(n1121), .Z(n1118) );
  XNOR U1481 ( .A(x[360]), .B(n1119), .Z(n1121) );
  XOR U1482 ( .A(n1122), .B(n1123), .Z(n1119) );
  AND U1483 ( .A(n1124), .B(n1125), .Z(n1122) );
  XNOR U1484 ( .A(x[359]), .B(n1123), .Z(n1125) );
  XOR U1485 ( .A(n1126), .B(n1127), .Z(n1123) );
  AND U1486 ( .A(n1128), .B(n1129), .Z(n1126) );
  XNOR U1487 ( .A(x[358]), .B(n1127), .Z(n1129) );
  XOR U1488 ( .A(n1130), .B(n1131), .Z(n1127) );
  AND U1489 ( .A(n1132), .B(n1133), .Z(n1130) );
  XNOR U1490 ( .A(x[357]), .B(n1131), .Z(n1133) );
  XOR U1491 ( .A(n1134), .B(n1135), .Z(n1131) );
  AND U1492 ( .A(n1136), .B(n1137), .Z(n1134) );
  XNOR U1493 ( .A(x[356]), .B(n1135), .Z(n1137) );
  XOR U1494 ( .A(n1138), .B(n1139), .Z(n1135) );
  AND U1495 ( .A(n1140), .B(n1141), .Z(n1138) );
  XNOR U1496 ( .A(x[355]), .B(n1139), .Z(n1141) );
  XOR U1497 ( .A(n1142), .B(n1143), .Z(n1139) );
  AND U1498 ( .A(n1144), .B(n1145), .Z(n1142) );
  XNOR U1499 ( .A(x[354]), .B(n1143), .Z(n1145) );
  XOR U1500 ( .A(n1146), .B(n1147), .Z(n1143) );
  AND U1501 ( .A(n1148), .B(n1149), .Z(n1146) );
  XNOR U1502 ( .A(x[353]), .B(n1147), .Z(n1149) );
  XOR U1503 ( .A(n1150), .B(n1151), .Z(n1147) );
  AND U1504 ( .A(n1152), .B(n1153), .Z(n1150) );
  XNOR U1505 ( .A(x[352]), .B(n1151), .Z(n1153) );
  XOR U1506 ( .A(n1154), .B(n1155), .Z(n1151) );
  AND U1507 ( .A(n1156), .B(n1157), .Z(n1154) );
  XNOR U1508 ( .A(x[351]), .B(n1155), .Z(n1157) );
  XOR U1509 ( .A(n1158), .B(n1159), .Z(n1155) );
  AND U1510 ( .A(n1160), .B(n1161), .Z(n1158) );
  XNOR U1511 ( .A(x[350]), .B(n1159), .Z(n1161) );
  XOR U1512 ( .A(n1162), .B(n1163), .Z(n1159) );
  AND U1513 ( .A(n1164), .B(n1165), .Z(n1162) );
  XNOR U1514 ( .A(x[349]), .B(n1163), .Z(n1165) );
  XOR U1515 ( .A(n1166), .B(n1167), .Z(n1163) );
  AND U1516 ( .A(n1168), .B(n1169), .Z(n1166) );
  XNOR U1517 ( .A(x[348]), .B(n1167), .Z(n1169) );
  XOR U1518 ( .A(n1170), .B(n1171), .Z(n1167) );
  AND U1519 ( .A(n1172), .B(n1173), .Z(n1170) );
  XNOR U1520 ( .A(x[347]), .B(n1171), .Z(n1173) );
  XOR U1521 ( .A(n1174), .B(n1175), .Z(n1171) );
  AND U1522 ( .A(n1176), .B(n1177), .Z(n1174) );
  XNOR U1523 ( .A(x[346]), .B(n1175), .Z(n1177) );
  XOR U1524 ( .A(n1178), .B(n1179), .Z(n1175) );
  AND U1525 ( .A(n1180), .B(n1181), .Z(n1178) );
  XNOR U1526 ( .A(x[345]), .B(n1179), .Z(n1181) );
  XOR U1527 ( .A(n1182), .B(n1183), .Z(n1179) );
  AND U1528 ( .A(n1184), .B(n1185), .Z(n1182) );
  XNOR U1529 ( .A(x[344]), .B(n1183), .Z(n1185) );
  XOR U1530 ( .A(n1186), .B(n1187), .Z(n1183) );
  AND U1531 ( .A(n1188), .B(n1189), .Z(n1186) );
  XNOR U1532 ( .A(x[343]), .B(n1187), .Z(n1189) );
  XOR U1533 ( .A(n1190), .B(n1191), .Z(n1187) );
  AND U1534 ( .A(n1192), .B(n1193), .Z(n1190) );
  XNOR U1535 ( .A(x[342]), .B(n1191), .Z(n1193) );
  XOR U1536 ( .A(n1194), .B(n1195), .Z(n1191) );
  AND U1537 ( .A(n1196), .B(n1197), .Z(n1194) );
  XNOR U1538 ( .A(x[341]), .B(n1195), .Z(n1197) );
  XOR U1539 ( .A(n1198), .B(n1199), .Z(n1195) );
  AND U1540 ( .A(n1200), .B(n1201), .Z(n1198) );
  XNOR U1541 ( .A(x[340]), .B(n1199), .Z(n1201) );
  XOR U1542 ( .A(n1202), .B(n1203), .Z(n1199) );
  AND U1543 ( .A(n1204), .B(n1205), .Z(n1202) );
  XNOR U1544 ( .A(x[339]), .B(n1203), .Z(n1205) );
  XOR U1545 ( .A(n1206), .B(n1207), .Z(n1203) );
  AND U1546 ( .A(n1208), .B(n1209), .Z(n1206) );
  XNOR U1547 ( .A(x[338]), .B(n1207), .Z(n1209) );
  XOR U1548 ( .A(n1210), .B(n1211), .Z(n1207) );
  AND U1549 ( .A(n1212), .B(n1213), .Z(n1210) );
  XNOR U1550 ( .A(x[337]), .B(n1211), .Z(n1213) );
  XOR U1551 ( .A(n1214), .B(n1215), .Z(n1211) );
  AND U1552 ( .A(n1216), .B(n1217), .Z(n1214) );
  XNOR U1553 ( .A(x[336]), .B(n1215), .Z(n1217) );
  XOR U1554 ( .A(n1218), .B(n1219), .Z(n1215) );
  AND U1555 ( .A(n1220), .B(n1221), .Z(n1218) );
  XNOR U1556 ( .A(x[335]), .B(n1219), .Z(n1221) );
  XOR U1557 ( .A(n1222), .B(n1223), .Z(n1219) );
  AND U1558 ( .A(n1224), .B(n1225), .Z(n1222) );
  XNOR U1559 ( .A(x[334]), .B(n1223), .Z(n1225) );
  XOR U1560 ( .A(n1226), .B(n1227), .Z(n1223) );
  AND U1561 ( .A(n1228), .B(n1229), .Z(n1226) );
  XNOR U1562 ( .A(x[333]), .B(n1227), .Z(n1229) );
  XOR U1563 ( .A(n1230), .B(n1231), .Z(n1227) );
  AND U1564 ( .A(n1232), .B(n1233), .Z(n1230) );
  XNOR U1565 ( .A(x[332]), .B(n1231), .Z(n1233) );
  XOR U1566 ( .A(n1234), .B(n1235), .Z(n1231) );
  AND U1567 ( .A(n1236), .B(n1237), .Z(n1234) );
  XNOR U1568 ( .A(x[331]), .B(n1235), .Z(n1237) );
  XOR U1569 ( .A(n1238), .B(n1239), .Z(n1235) );
  AND U1570 ( .A(n1240), .B(n1241), .Z(n1238) );
  XNOR U1571 ( .A(x[330]), .B(n1239), .Z(n1241) );
  XOR U1572 ( .A(n1242), .B(n1243), .Z(n1239) );
  AND U1573 ( .A(n1244), .B(n1245), .Z(n1242) );
  XNOR U1574 ( .A(x[329]), .B(n1243), .Z(n1245) );
  XOR U1575 ( .A(n1246), .B(n1247), .Z(n1243) );
  AND U1576 ( .A(n1248), .B(n1249), .Z(n1246) );
  XNOR U1577 ( .A(x[328]), .B(n1247), .Z(n1249) );
  XOR U1578 ( .A(n1250), .B(n1251), .Z(n1247) );
  AND U1579 ( .A(n1252), .B(n1253), .Z(n1250) );
  XNOR U1580 ( .A(x[327]), .B(n1251), .Z(n1253) );
  XOR U1581 ( .A(n1254), .B(n1255), .Z(n1251) );
  AND U1582 ( .A(n1256), .B(n1257), .Z(n1254) );
  XNOR U1583 ( .A(x[326]), .B(n1255), .Z(n1257) );
  XOR U1584 ( .A(n1258), .B(n1259), .Z(n1255) );
  AND U1585 ( .A(n1260), .B(n1261), .Z(n1258) );
  XNOR U1586 ( .A(x[325]), .B(n1259), .Z(n1261) );
  XOR U1587 ( .A(n1262), .B(n1263), .Z(n1259) );
  AND U1588 ( .A(n1264), .B(n1265), .Z(n1262) );
  XNOR U1589 ( .A(x[324]), .B(n1263), .Z(n1265) );
  XOR U1590 ( .A(n1266), .B(n1267), .Z(n1263) );
  AND U1591 ( .A(n1268), .B(n1269), .Z(n1266) );
  XNOR U1592 ( .A(x[323]), .B(n1267), .Z(n1269) );
  XOR U1593 ( .A(n1270), .B(n1271), .Z(n1267) );
  AND U1594 ( .A(n1272), .B(n1273), .Z(n1270) );
  XNOR U1595 ( .A(x[322]), .B(n1271), .Z(n1273) );
  XOR U1596 ( .A(n1274), .B(n1275), .Z(n1271) );
  AND U1597 ( .A(n1276), .B(n1277), .Z(n1274) );
  XNOR U1598 ( .A(x[321]), .B(n1275), .Z(n1277) );
  XOR U1599 ( .A(n1278), .B(n1279), .Z(n1275) );
  AND U1600 ( .A(n1280), .B(n1281), .Z(n1278) );
  XNOR U1601 ( .A(x[320]), .B(n1279), .Z(n1281) );
  XOR U1602 ( .A(n1282), .B(n1283), .Z(n1279) );
  AND U1603 ( .A(n1284), .B(n1285), .Z(n1282) );
  XNOR U1604 ( .A(x[319]), .B(n1283), .Z(n1285) );
  XOR U1605 ( .A(n1286), .B(n1287), .Z(n1283) );
  AND U1606 ( .A(n1288), .B(n1289), .Z(n1286) );
  XNOR U1607 ( .A(x[318]), .B(n1287), .Z(n1289) );
  XOR U1608 ( .A(n1290), .B(n1291), .Z(n1287) );
  AND U1609 ( .A(n1292), .B(n1293), .Z(n1290) );
  XNOR U1610 ( .A(x[317]), .B(n1291), .Z(n1293) );
  XOR U1611 ( .A(n1294), .B(n1295), .Z(n1291) );
  AND U1612 ( .A(n1296), .B(n1297), .Z(n1294) );
  XNOR U1613 ( .A(x[316]), .B(n1295), .Z(n1297) );
  XOR U1614 ( .A(n1298), .B(n1299), .Z(n1295) );
  AND U1615 ( .A(n1300), .B(n1301), .Z(n1298) );
  XNOR U1616 ( .A(x[315]), .B(n1299), .Z(n1301) );
  XOR U1617 ( .A(n1302), .B(n1303), .Z(n1299) );
  AND U1618 ( .A(n1304), .B(n1305), .Z(n1302) );
  XNOR U1619 ( .A(x[314]), .B(n1303), .Z(n1305) );
  XOR U1620 ( .A(n1306), .B(n1307), .Z(n1303) );
  AND U1621 ( .A(n1308), .B(n1309), .Z(n1306) );
  XNOR U1622 ( .A(x[313]), .B(n1307), .Z(n1309) );
  XOR U1623 ( .A(n1310), .B(n1311), .Z(n1307) );
  AND U1624 ( .A(n1312), .B(n1313), .Z(n1310) );
  XNOR U1625 ( .A(x[312]), .B(n1311), .Z(n1313) );
  XOR U1626 ( .A(n1314), .B(n1315), .Z(n1311) );
  AND U1627 ( .A(n1316), .B(n1317), .Z(n1314) );
  XNOR U1628 ( .A(x[311]), .B(n1315), .Z(n1317) );
  XOR U1629 ( .A(n1318), .B(n1319), .Z(n1315) );
  AND U1630 ( .A(n1320), .B(n1321), .Z(n1318) );
  XNOR U1631 ( .A(x[310]), .B(n1319), .Z(n1321) );
  XOR U1632 ( .A(n1322), .B(n1323), .Z(n1319) );
  AND U1633 ( .A(n1324), .B(n1325), .Z(n1322) );
  XNOR U1634 ( .A(x[309]), .B(n1323), .Z(n1325) );
  XOR U1635 ( .A(n1326), .B(n1327), .Z(n1323) );
  AND U1636 ( .A(n1328), .B(n1329), .Z(n1326) );
  XNOR U1637 ( .A(x[308]), .B(n1327), .Z(n1329) );
  XOR U1638 ( .A(n1330), .B(n1331), .Z(n1327) );
  AND U1639 ( .A(n1332), .B(n1333), .Z(n1330) );
  XNOR U1640 ( .A(x[307]), .B(n1331), .Z(n1333) );
  XOR U1641 ( .A(n1334), .B(n1335), .Z(n1331) );
  AND U1642 ( .A(n1336), .B(n1337), .Z(n1334) );
  XNOR U1643 ( .A(x[306]), .B(n1335), .Z(n1337) );
  XOR U1644 ( .A(n1338), .B(n1339), .Z(n1335) );
  AND U1645 ( .A(n1340), .B(n1341), .Z(n1338) );
  XNOR U1646 ( .A(x[305]), .B(n1339), .Z(n1341) );
  XOR U1647 ( .A(n1342), .B(n1343), .Z(n1339) );
  AND U1648 ( .A(n1344), .B(n1345), .Z(n1342) );
  XNOR U1649 ( .A(x[304]), .B(n1343), .Z(n1345) );
  XOR U1650 ( .A(n1346), .B(n1347), .Z(n1343) );
  AND U1651 ( .A(n1348), .B(n1349), .Z(n1346) );
  XNOR U1652 ( .A(x[303]), .B(n1347), .Z(n1349) );
  XOR U1653 ( .A(n1350), .B(n1351), .Z(n1347) );
  AND U1654 ( .A(n1352), .B(n1353), .Z(n1350) );
  XNOR U1655 ( .A(x[302]), .B(n1351), .Z(n1353) );
  XOR U1656 ( .A(n1354), .B(n1355), .Z(n1351) );
  AND U1657 ( .A(n1356), .B(n1357), .Z(n1354) );
  XNOR U1658 ( .A(x[301]), .B(n1355), .Z(n1357) );
  XOR U1659 ( .A(n1358), .B(n1359), .Z(n1355) );
  AND U1660 ( .A(n1360), .B(n1361), .Z(n1358) );
  XNOR U1661 ( .A(x[300]), .B(n1359), .Z(n1361) );
  XOR U1662 ( .A(n1362), .B(n1363), .Z(n1359) );
  AND U1663 ( .A(n1364), .B(n1365), .Z(n1362) );
  XNOR U1664 ( .A(x[299]), .B(n1363), .Z(n1365) );
  XOR U1665 ( .A(n1366), .B(n1367), .Z(n1363) );
  AND U1666 ( .A(n1368), .B(n1369), .Z(n1366) );
  XNOR U1667 ( .A(x[298]), .B(n1367), .Z(n1369) );
  XOR U1668 ( .A(n1370), .B(n1371), .Z(n1367) );
  AND U1669 ( .A(n1372), .B(n1373), .Z(n1370) );
  XNOR U1670 ( .A(x[297]), .B(n1371), .Z(n1373) );
  XOR U1671 ( .A(n1374), .B(n1375), .Z(n1371) );
  AND U1672 ( .A(n1376), .B(n1377), .Z(n1374) );
  XNOR U1673 ( .A(x[296]), .B(n1375), .Z(n1377) );
  XOR U1674 ( .A(n1378), .B(n1379), .Z(n1375) );
  AND U1675 ( .A(n1380), .B(n1381), .Z(n1378) );
  XNOR U1676 ( .A(x[295]), .B(n1379), .Z(n1381) );
  XOR U1677 ( .A(n1382), .B(n1383), .Z(n1379) );
  AND U1678 ( .A(n1384), .B(n1385), .Z(n1382) );
  XNOR U1679 ( .A(x[294]), .B(n1383), .Z(n1385) );
  XOR U1680 ( .A(n1386), .B(n1387), .Z(n1383) );
  AND U1681 ( .A(n1388), .B(n1389), .Z(n1386) );
  XNOR U1682 ( .A(x[293]), .B(n1387), .Z(n1389) );
  XOR U1683 ( .A(n1390), .B(n1391), .Z(n1387) );
  AND U1684 ( .A(n1392), .B(n1393), .Z(n1390) );
  XNOR U1685 ( .A(x[292]), .B(n1391), .Z(n1393) );
  XOR U1686 ( .A(n1394), .B(n1395), .Z(n1391) );
  AND U1687 ( .A(n1396), .B(n1397), .Z(n1394) );
  XNOR U1688 ( .A(x[291]), .B(n1395), .Z(n1397) );
  XOR U1689 ( .A(n1398), .B(n1399), .Z(n1395) );
  AND U1690 ( .A(n1400), .B(n1401), .Z(n1398) );
  XNOR U1691 ( .A(x[290]), .B(n1399), .Z(n1401) );
  XOR U1692 ( .A(n1402), .B(n1403), .Z(n1399) );
  AND U1693 ( .A(n1404), .B(n1405), .Z(n1402) );
  XNOR U1694 ( .A(x[289]), .B(n1403), .Z(n1405) );
  XOR U1695 ( .A(n1406), .B(n1407), .Z(n1403) );
  AND U1696 ( .A(n1408), .B(n1409), .Z(n1406) );
  XNOR U1697 ( .A(x[288]), .B(n1407), .Z(n1409) );
  XOR U1698 ( .A(n1410), .B(n1411), .Z(n1407) );
  AND U1699 ( .A(n1412), .B(n1413), .Z(n1410) );
  XNOR U1700 ( .A(x[287]), .B(n1411), .Z(n1413) );
  XOR U1701 ( .A(n1414), .B(n1415), .Z(n1411) );
  AND U1702 ( .A(n1416), .B(n1417), .Z(n1414) );
  XNOR U1703 ( .A(x[286]), .B(n1415), .Z(n1417) );
  XOR U1704 ( .A(n1418), .B(n1419), .Z(n1415) );
  AND U1705 ( .A(n1420), .B(n1421), .Z(n1418) );
  XNOR U1706 ( .A(x[285]), .B(n1419), .Z(n1421) );
  XOR U1707 ( .A(n1422), .B(n1423), .Z(n1419) );
  AND U1708 ( .A(n1424), .B(n1425), .Z(n1422) );
  XNOR U1709 ( .A(x[284]), .B(n1423), .Z(n1425) );
  XOR U1710 ( .A(n1426), .B(n1427), .Z(n1423) );
  AND U1711 ( .A(n1428), .B(n1429), .Z(n1426) );
  XNOR U1712 ( .A(x[283]), .B(n1427), .Z(n1429) );
  XOR U1713 ( .A(n1430), .B(n1431), .Z(n1427) );
  AND U1714 ( .A(n1432), .B(n1433), .Z(n1430) );
  XNOR U1715 ( .A(x[282]), .B(n1431), .Z(n1433) );
  XOR U1716 ( .A(n1434), .B(n1435), .Z(n1431) );
  AND U1717 ( .A(n1436), .B(n1437), .Z(n1434) );
  XNOR U1718 ( .A(x[281]), .B(n1435), .Z(n1437) );
  XOR U1719 ( .A(n1438), .B(n1439), .Z(n1435) );
  AND U1720 ( .A(n1440), .B(n1441), .Z(n1438) );
  XNOR U1721 ( .A(x[280]), .B(n1439), .Z(n1441) );
  XOR U1722 ( .A(n1442), .B(n1443), .Z(n1439) );
  AND U1723 ( .A(n1444), .B(n1445), .Z(n1442) );
  XNOR U1724 ( .A(x[279]), .B(n1443), .Z(n1445) );
  XOR U1725 ( .A(n1446), .B(n1447), .Z(n1443) );
  AND U1726 ( .A(n1448), .B(n1449), .Z(n1446) );
  XNOR U1727 ( .A(x[278]), .B(n1447), .Z(n1449) );
  XOR U1728 ( .A(n1450), .B(n1451), .Z(n1447) );
  AND U1729 ( .A(n1452), .B(n1453), .Z(n1450) );
  XNOR U1730 ( .A(x[277]), .B(n1451), .Z(n1453) );
  XOR U1731 ( .A(n1454), .B(n1455), .Z(n1451) );
  AND U1732 ( .A(n1456), .B(n1457), .Z(n1454) );
  XNOR U1733 ( .A(x[276]), .B(n1455), .Z(n1457) );
  XOR U1734 ( .A(n1458), .B(n1459), .Z(n1455) );
  AND U1735 ( .A(n1460), .B(n1461), .Z(n1458) );
  XNOR U1736 ( .A(x[275]), .B(n1459), .Z(n1461) );
  XOR U1737 ( .A(n1462), .B(n1463), .Z(n1459) );
  AND U1738 ( .A(n1464), .B(n1465), .Z(n1462) );
  XNOR U1739 ( .A(x[274]), .B(n1463), .Z(n1465) );
  XOR U1740 ( .A(n1466), .B(n1467), .Z(n1463) );
  AND U1741 ( .A(n1468), .B(n1469), .Z(n1466) );
  XNOR U1742 ( .A(x[273]), .B(n1467), .Z(n1469) );
  XOR U1743 ( .A(n1470), .B(n1471), .Z(n1467) );
  AND U1744 ( .A(n1472), .B(n1473), .Z(n1470) );
  XNOR U1745 ( .A(x[272]), .B(n1471), .Z(n1473) );
  XOR U1746 ( .A(n1474), .B(n1475), .Z(n1471) );
  AND U1747 ( .A(n1476), .B(n1477), .Z(n1474) );
  XNOR U1748 ( .A(x[271]), .B(n1475), .Z(n1477) );
  XOR U1749 ( .A(n1478), .B(n1479), .Z(n1475) );
  AND U1750 ( .A(n1480), .B(n1481), .Z(n1478) );
  XNOR U1751 ( .A(x[270]), .B(n1479), .Z(n1481) );
  XOR U1752 ( .A(n1482), .B(n1483), .Z(n1479) );
  AND U1753 ( .A(n1484), .B(n1485), .Z(n1482) );
  XNOR U1754 ( .A(x[269]), .B(n1483), .Z(n1485) );
  XOR U1755 ( .A(n1486), .B(n1487), .Z(n1483) );
  AND U1756 ( .A(n1488), .B(n1489), .Z(n1486) );
  XNOR U1757 ( .A(x[268]), .B(n1487), .Z(n1489) );
  XOR U1758 ( .A(n1490), .B(n1491), .Z(n1487) );
  AND U1759 ( .A(n1492), .B(n1493), .Z(n1490) );
  XNOR U1760 ( .A(x[267]), .B(n1491), .Z(n1493) );
  XOR U1761 ( .A(n1494), .B(n1495), .Z(n1491) );
  AND U1762 ( .A(n1496), .B(n1497), .Z(n1494) );
  XNOR U1763 ( .A(x[266]), .B(n1495), .Z(n1497) );
  XOR U1764 ( .A(n1498), .B(n1499), .Z(n1495) );
  AND U1765 ( .A(n1500), .B(n1501), .Z(n1498) );
  XNOR U1766 ( .A(x[265]), .B(n1499), .Z(n1501) );
  XOR U1767 ( .A(n1502), .B(n1503), .Z(n1499) );
  AND U1768 ( .A(n1504), .B(n1505), .Z(n1502) );
  XNOR U1769 ( .A(x[264]), .B(n1503), .Z(n1505) );
  XOR U1770 ( .A(n1506), .B(n1507), .Z(n1503) );
  AND U1771 ( .A(n1508), .B(n1509), .Z(n1506) );
  XNOR U1772 ( .A(x[263]), .B(n1507), .Z(n1509) );
  XOR U1773 ( .A(n1510), .B(n1511), .Z(n1507) );
  AND U1774 ( .A(n1512), .B(n1513), .Z(n1510) );
  XNOR U1775 ( .A(x[262]), .B(n1511), .Z(n1513) );
  XOR U1776 ( .A(n1514), .B(n1515), .Z(n1511) );
  AND U1777 ( .A(n1516), .B(n1517), .Z(n1514) );
  XNOR U1778 ( .A(x[261]), .B(n1515), .Z(n1517) );
  XOR U1779 ( .A(n1518), .B(n1519), .Z(n1515) );
  AND U1780 ( .A(n1520), .B(n1521), .Z(n1518) );
  XNOR U1781 ( .A(x[260]), .B(n1519), .Z(n1521) );
  XOR U1782 ( .A(n1522), .B(n1523), .Z(n1519) );
  AND U1783 ( .A(n1524), .B(n1525), .Z(n1522) );
  XNOR U1784 ( .A(x[259]), .B(n1523), .Z(n1525) );
  XOR U1785 ( .A(n1526), .B(n1527), .Z(n1523) );
  AND U1786 ( .A(n1528), .B(n1529), .Z(n1526) );
  XNOR U1787 ( .A(x[258]), .B(n1527), .Z(n1529) );
  XOR U1788 ( .A(n1530), .B(n1531), .Z(n1527) );
  AND U1789 ( .A(n1532), .B(n1533), .Z(n1530) );
  XNOR U1790 ( .A(x[257]), .B(n1531), .Z(n1533) );
  XOR U1791 ( .A(n1534), .B(n1535), .Z(n1531) );
  AND U1792 ( .A(n1536), .B(n1537), .Z(n1534) );
  XNOR U1793 ( .A(x[256]), .B(n1535), .Z(n1537) );
  XOR U1794 ( .A(n1538), .B(n1539), .Z(n1535) );
  AND U1795 ( .A(n1540), .B(n1541), .Z(n1538) );
  XNOR U1796 ( .A(x[255]), .B(n1539), .Z(n1541) );
  XOR U1797 ( .A(n1542), .B(n1543), .Z(n1539) );
  AND U1798 ( .A(n1544), .B(n1545), .Z(n1542) );
  XNOR U1799 ( .A(x[254]), .B(n1543), .Z(n1545) );
  XOR U1800 ( .A(n1546), .B(n1547), .Z(n1543) );
  AND U1801 ( .A(n1548), .B(n1549), .Z(n1546) );
  XNOR U1802 ( .A(x[253]), .B(n1547), .Z(n1549) );
  XOR U1803 ( .A(n1550), .B(n1551), .Z(n1547) );
  AND U1804 ( .A(n1552), .B(n1553), .Z(n1550) );
  XNOR U1805 ( .A(x[252]), .B(n1551), .Z(n1553) );
  XOR U1806 ( .A(n1554), .B(n1555), .Z(n1551) );
  AND U1807 ( .A(n1556), .B(n1557), .Z(n1554) );
  XNOR U1808 ( .A(x[251]), .B(n1555), .Z(n1557) );
  XOR U1809 ( .A(n1558), .B(n1559), .Z(n1555) );
  AND U1810 ( .A(n1560), .B(n1561), .Z(n1558) );
  XNOR U1811 ( .A(x[250]), .B(n1559), .Z(n1561) );
  XOR U1812 ( .A(n1562), .B(n1563), .Z(n1559) );
  AND U1813 ( .A(n1564), .B(n1565), .Z(n1562) );
  XNOR U1814 ( .A(x[249]), .B(n1563), .Z(n1565) );
  XOR U1815 ( .A(n1566), .B(n1567), .Z(n1563) );
  AND U1816 ( .A(n1568), .B(n1569), .Z(n1566) );
  XNOR U1817 ( .A(x[248]), .B(n1567), .Z(n1569) );
  XOR U1818 ( .A(n1570), .B(n1571), .Z(n1567) );
  AND U1819 ( .A(n1572), .B(n1573), .Z(n1570) );
  XNOR U1820 ( .A(x[247]), .B(n1571), .Z(n1573) );
  XOR U1821 ( .A(n1574), .B(n1575), .Z(n1571) );
  AND U1822 ( .A(n1576), .B(n1577), .Z(n1574) );
  XNOR U1823 ( .A(x[246]), .B(n1575), .Z(n1577) );
  XOR U1824 ( .A(n1578), .B(n1579), .Z(n1575) );
  AND U1825 ( .A(n1580), .B(n1581), .Z(n1578) );
  XNOR U1826 ( .A(x[245]), .B(n1579), .Z(n1581) );
  XOR U1827 ( .A(n1582), .B(n1583), .Z(n1579) );
  AND U1828 ( .A(n1584), .B(n1585), .Z(n1582) );
  XNOR U1829 ( .A(x[244]), .B(n1583), .Z(n1585) );
  XOR U1830 ( .A(n1586), .B(n1587), .Z(n1583) );
  AND U1831 ( .A(n1588), .B(n1589), .Z(n1586) );
  XNOR U1832 ( .A(x[243]), .B(n1587), .Z(n1589) );
  XOR U1833 ( .A(n1590), .B(n1591), .Z(n1587) );
  AND U1834 ( .A(n1592), .B(n1593), .Z(n1590) );
  XNOR U1835 ( .A(x[242]), .B(n1591), .Z(n1593) );
  XOR U1836 ( .A(n1594), .B(n1595), .Z(n1591) );
  AND U1837 ( .A(n1596), .B(n1597), .Z(n1594) );
  XNOR U1838 ( .A(x[241]), .B(n1595), .Z(n1597) );
  XOR U1839 ( .A(n1598), .B(n1599), .Z(n1595) );
  AND U1840 ( .A(n1600), .B(n1601), .Z(n1598) );
  XNOR U1841 ( .A(x[240]), .B(n1599), .Z(n1601) );
  XOR U1842 ( .A(n1602), .B(n1603), .Z(n1599) );
  AND U1843 ( .A(n1604), .B(n1605), .Z(n1602) );
  XNOR U1844 ( .A(x[239]), .B(n1603), .Z(n1605) );
  XOR U1845 ( .A(n1606), .B(n1607), .Z(n1603) );
  AND U1846 ( .A(n1608), .B(n1609), .Z(n1606) );
  XNOR U1847 ( .A(x[238]), .B(n1607), .Z(n1609) );
  XOR U1848 ( .A(n1610), .B(n1611), .Z(n1607) );
  AND U1849 ( .A(n1612), .B(n1613), .Z(n1610) );
  XNOR U1850 ( .A(x[237]), .B(n1611), .Z(n1613) );
  XOR U1851 ( .A(n1614), .B(n1615), .Z(n1611) );
  AND U1852 ( .A(n1616), .B(n1617), .Z(n1614) );
  XNOR U1853 ( .A(x[236]), .B(n1615), .Z(n1617) );
  XOR U1854 ( .A(n1618), .B(n1619), .Z(n1615) );
  AND U1855 ( .A(n1620), .B(n1621), .Z(n1618) );
  XNOR U1856 ( .A(x[235]), .B(n1619), .Z(n1621) );
  XOR U1857 ( .A(n1622), .B(n1623), .Z(n1619) );
  AND U1858 ( .A(n1624), .B(n1625), .Z(n1622) );
  XNOR U1859 ( .A(x[234]), .B(n1623), .Z(n1625) );
  XOR U1860 ( .A(n1626), .B(n1627), .Z(n1623) );
  AND U1861 ( .A(n1628), .B(n1629), .Z(n1626) );
  XNOR U1862 ( .A(x[233]), .B(n1627), .Z(n1629) );
  XOR U1863 ( .A(n1630), .B(n1631), .Z(n1627) );
  AND U1864 ( .A(n1632), .B(n1633), .Z(n1630) );
  XNOR U1865 ( .A(x[232]), .B(n1631), .Z(n1633) );
  XOR U1866 ( .A(n1634), .B(n1635), .Z(n1631) );
  AND U1867 ( .A(n1636), .B(n1637), .Z(n1634) );
  XNOR U1868 ( .A(x[231]), .B(n1635), .Z(n1637) );
  XOR U1869 ( .A(n1638), .B(n1639), .Z(n1635) );
  AND U1870 ( .A(n1640), .B(n1641), .Z(n1638) );
  XNOR U1871 ( .A(x[230]), .B(n1639), .Z(n1641) );
  XOR U1872 ( .A(n1642), .B(n1643), .Z(n1639) );
  AND U1873 ( .A(n1644), .B(n1645), .Z(n1642) );
  XNOR U1874 ( .A(x[229]), .B(n1643), .Z(n1645) );
  XOR U1875 ( .A(n1646), .B(n1647), .Z(n1643) );
  AND U1876 ( .A(n1648), .B(n1649), .Z(n1646) );
  XNOR U1877 ( .A(x[228]), .B(n1647), .Z(n1649) );
  XOR U1878 ( .A(n1650), .B(n1651), .Z(n1647) );
  AND U1879 ( .A(n1652), .B(n1653), .Z(n1650) );
  XNOR U1880 ( .A(x[227]), .B(n1651), .Z(n1653) );
  XOR U1881 ( .A(n1654), .B(n1655), .Z(n1651) );
  AND U1882 ( .A(n1656), .B(n1657), .Z(n1654) );
  XNOR U1883 ( .A(x[226]), .B(n1655), .Z(n1657) );
  XOR U1884 ( .A(n1658), .B(n1659), .Z(n1655) );
  AND U1885 ( .A(n1660), .B(n1661), .Z(n1658) );
  XNOR U1886 ( .A(x[225]), .B(n1659), .Z(n1661) );
  XOR U1887 ( .A(n1662), .B(n1663), .Z(n1659) );
  AND U1888 ( .A(n1664), .B(n1665), .Z(n1662) );
  XNOR U1889 ( .A(x[224]), .B(n1663), .Z(n1665) );
  XOR U1890 ( .A(n1666), .B(n1667), .Z(n1663) );
  AND U1891 ( .A(n1668), .B(n1669), .Z(n1666) );
  XNOR U1892 ( .A(x[223]), .B(n1667), .Z(n1669) );
  XOR U1893 ( .A(n1670), .B(n1671), .Z(n1667) );
  AND U1894 ( .A(n1672), .B(n1673), .Z(n1670) );
  XNOR U1895 ( .A(x[222]), .B(n1671), .Z(n1673) );
  XOR U1896 ( .A(n1674), .B(n1675), .Z(n1671) );
  AND U1897 ( .A(n1676), .B(n1677), .Z(n1674) );
  XNOR U1898 ( .A(x[221]), .B(n1675), .Z(n1677) );
  XOR U1899 ( .A(n1678), .B(n1679), .Z(n1675) );
  AND U1900 ( .A(n1680), .B(n1681), .Z(n1678) );
  XNOR U1901 ( .A(x[220]), .B(n1679), .Z(n1681) );
  XOR U1902 ( .A(n1682), .B(n1683), .Z(n1679) );
  AND U1903 ( .A(n1684), .B(n1685), .Z(n1682) );
  XNOR U1904 ( .A(x[219]), .B(n1683), .Z(n1685) );
  XOR U1905 ( .A(n1686), .B(n1687), .Z(n1683) );
  AND U1906 ( .A(n1688), .B(n1689), .Z(n1686) );
  XNOR U1907 ( .A(x[218]), .B(n1687), .Z(n1689) );
  XOR U1908 ( .A(n1690), .B(n1691), .Z(n1687) );
  AND U1909 ( .A(n1692), .B(n1693), .Z(n1690) );
  XNOR U1910 ( .A(x[217]), .B(n1691), .Z(n1693) );
  XOR U1911 ( .A(n1694), .B(n1695), .Z(n1691) );
  AND U1912 ( .A(n1696), .B(n1697), .Z(n1694) );
  XNOR U1913 ( .A(x[216]), .B(n1695), .Z(n1697) );
  XOR U1914 ( .A(n1698), .B(n1699), .Z(n1695) );
  AND U1915 ( .A(n1700), .B(n1701), .Z(n1698) );
  XNOR U1916 ( .A(x[215]), .B(n1699), .Z(n1701) );
  XOR U1917 ( .A(n1702), .B(n1703), .Z(n1699) );
  AND U1918 ( .A(n1704), .B(n1705), .Z(n1702) );
  XNOR U1919 ( .A(x[214]), .B(n1703), .Z(n1705) );
  XOR U1920 ( .A(n1706), .B(n1707), .Z(n1703) );
  AND U1921 ( .A(n1708), .B(n1709), .Z(n1706) );
  XNOR U1922 ( .A(x[213]), .B(n1707), .Z(n1709) );
  XOR U1923 ( .A(n1710), .B(n1711), .Z(n1707) );
  AND U1924 ( .A(n1712), .B(n1713), .Z(n1710) );
  XNOR U1925 ( .A(x[212]), .B(n1711), .Z(n1713) );
  XOR U1926 ( .A(n1714), .B(n1715), .Z(n1711) );
  AND U1927 ( .A(n1716), .B(n1717), .Z(n1714) );
  XNOR U1928 ( .A(x[211]), .B(n1715), .Z(n1717) );
  XOR U1929 ( .A(n1718), .B(n1719), .Z(n1715) );
  AND U1930 ( .A(n1720), .B(n1721), .Z(n1718) );
  XNOR U1931 ( .A(x[210]), .B(n1719), .Z(n1721) );
  XOR U1932 ( .A(n1722), .B(n1723), .Z(n1719) );
  AND U1933 ( .A(n1724), .B(n1725), .Z(n1722) );
  XNOR U1934 ( .A(x[209]), .B(n1723), .Z(n1725) );
  XOR U1935 ( .A(n1726), .B(n1727), .Z(n1723) );
  AND U1936 ( .A(n1728), .B(n1729), .Z(n1726) );
  XNOR U1937 ( .A(x[208]), .B(n1727), .Z(n1729) );
  XOR U1938 ( .A(n1730), .B(n1731), .Z(n1727) );
  AND U1939 ( .A(n1732), .B(n1733), .Z(n1730) );
  XNOR U1940 ( .A(x[207]), .B(n1731), .Z(n1733) );
  XOR U1941 ( .A(n1734), .B(n1735), .Z(n1731) );
  AND U1942 ( .A(n1736), .B(n1737), .Z(n1734) );
  XNOR U1943 ( .A(x[206]), .B(n1735), .Z(n1737) );
  XOR U1944 ( .A(n1738), .B(n1739), .Z(n1735) );
  AND U1945 ( .A(n1740), .B(n1741), .Z(n1738) );
  XNOR U1946 ( .A(x[205]), .B(n1739), .Z(n1741) );
  XOR U1947 ( .A(n1742), .B(n1743), .Z(n1739) );
  AND U1948 ( .A(n1744), .B(n1745), .Z(n1742) );
  XNOR U1949 ( .A(x[204]), .B(n1743), .Z(n1745) );
  XOR U1950 ( .A(n1746), .B(n1747), .Z(n1743) );
  AND U1951 ( .A(n1748), .B(n1749), .Z(n1746) );
  XNOR U1952 ( .A(x[203]), .B(n1747), .Z(n1749) );
  XOR U1953 ( .A(n1750), .B(n1751), .Z(n1747) );
  AND U1954 ( .A(n1752), .B(n1753), .Z(n1750) );
  XNOR U1955 ( .A(x[202]), .B(n1751), .Z(n1753) );
  XOR U1956 ( .A(n1754), .B(n1755), .Z(n1751) );
  AND U1957 ( .A(n1756), .B(n1757), .Z(n1754) );
  XNOR U1958 ( .A(x[201]), .B(n1755), .Z(n1757) );
  XOR U1959 ( .A(n1758), .B(n1759), .Z(n1755) );
  AND U1960 ( .A(n1760), .B(n1761), .Z(n1758) );
  XNOR U1961 ( .A(x[200]), .B(n1759), .Z(n1761) );
  XOR U1962 ( .A(n1762), .B(n1763), .Z(n1759) );
  AND U1963 ( .A(n1764), .B(n1765), .Z(n1762) );
  XNOR U1964 ( .A(x[199]), .B(n1763), .Z(n1765) );
  XOR U1965 ( .A(n1766), .B(n1767), .Z(n1763) );
  AND U1966 ( .A(n1768), .B(n1769), .Z(n1766) );
  XNOR U1967 ( .A(x[198]), .B(n1767), .Z(n1769) );
  XOR U1968 ( .A(n1770), .B(n1771), .Z(n1767) );
  AND U1969 ( .A(n1772), .B(n1773), .Z(n1770) );
  XNOR U1970 ( .A(x[197]), .B(n1771), .Z(n1773) );
  XOR U1971 ( .A(n1774), .B(n1775), .Z(n1771) );
  AND U1972 ( .A(n1776), .B(n1777), .Z(n1774) );
  XNOR U1973 ( .A(x[196]), .B(n1775), .Z(n1777) );
  XOR U1974 ( .A(n1778), .B(n1779), .Z(n1775) );
  AND U1975 ( .A(n1780), .B(n1781), .Z(n1778) );
  XNOR U1976 ( .A(x[195]), .B(n1779), .Z(n1781) );
  XOR U1977 ( .A(n1782), .B(n1783), .Z(n1779) );
  AND U1978 ( .A(n1784), .B(n1785), .Z(n1782) );
  XNOR U1979 ( .A(x[194]), .B(n1783), .Z(n1785) );
  XOR U1980 ( .A(n1786), .B(n1787), .Z(n1783) );
  AND U1981 ( .A(n1788), .B(n1789), .Z(n1786) );
  XNOR U1982 ( .A(x[193]), .B(n1787), .Z(n1789) );
  XOR U1983 ( .A(n1790), .B(n1791), .Z(n1787) );
  AND U1984 ( .A(n1792), .B(n1793), .Z(n1790) );
  XNOR U1985 ( .A(x[192]), .B(n1791), .Z(n1793) );
  XOR U1986 ( .A(n1794), .B(n1795), .Z(n1791) );
  AND U1987 ( .A(n1796), .B(n1797), .Z(n1794) );
  XNOR U1988 ( .A(x[191]), .B(n1795), .Z(n1797) );
  XOR U1989 ( .A(n1798), .B(n1799), .Z(n1795) );
  AND U1990 ( .A(n1800), .B(n1801), .Z(n1798) );
  XNOR U1991 ( .A(x[190]), .B(n1799), .Z(n1801) );
  XOR U1992 ( .A(n1802), .B(n1803), .Z(n1799) );
  AND U1993 ( .A(n1804), .B(n1805), .Z(n1802) );
  XNOR U1994 ( .A(x[189]), .B(n1803), .Z(n1805) );
  XOR U1995 ( .A(n1806), .B(n1807), .Z(n1803) );
  AND U1996 ( .A(n1808), .B(n1809), .Z(n1806) );
  XNOR U1997 ( .A(x[188]), .B(n1807), .Z(n1809) );
  XOR U1998 ( .A(n1810), .B(n1811), .Z(n1807) );
  AND U1999 ( .A(n1812), .B(n1813), .Z(n1810) );
  XNOR U2000 ( .A(x[187]), .B(n1811), .Z(n1813) );
  XOR U2001 ( .A(n1814), .B(n1815), .Z(n1811) );
  AND U2002 ( .A(n1816), .B(n1817), .Z(n1814) );
  XNOR U2003 ( .A(x[186]), .B(n1815), .Z(n1817) );
  XOR U2004 ( .A(n1818), .B(n1819), .Z(n1815) );
  AND U2005 ( .A(n1820), .B(n1821), .Z(n1818) );
  XNOR U2006 ( .A(x[185]), .B(n1819), .Z(n1821) );
  XOR U2007 ( .A(n1822), .B(n1823), .Z(n1819) );
  AND U2008 ( .A(n1824), .B(n1825), .Z(n1822) );
  XNOR U2009 ( .A(x[184]), .B(n1823), .Z(n1825) );
  XOR U2010 ( .A(n1826), .B(n1827), .Z(n1823) );
  AND U2011 ( .A(n1828), .B(n1829), .Z(n1826) );
  XNOR U2012 ( .A(x[183]), .B(n1827), .Z(n1829) );
  XOR U2013 ( .A(n1830), .B(n1831), .Z(n1827) );
  AND U2014 ( .A(n1832), .B(n1833), .Z(n1830) );
  XNOR U2015 ( .A(x[182]), .B(n1831), .Z(n1833) );
  XOR U2016 ( .A(n1834), .B(n1835), .Z(n1831) );
  AND U2017 ( .A(n1836), .B(n1837), .Z(n1834) );
  XNOR U2018 ( .A(x[181]), .B(n1835), .Z(n1837) );
  XOR U2019 ( .A(n1838), .B(n1839), .Z(n1835) );
  AND U2020 ( .A(n1840), .B(n1841), .Z(n1838) );
  XNOR U2021 ( .A(x[180]), .B(n1839), .Z(n1841) );
  XOR U2022 ( .A(n1842), .B(n1843), .Z(n1839) );
  AND U2023 ( .A(n1844), .B(n1845), .Z(n1842) );
  XNOR U2024 ( .A(x[179]), .B(n1843), .Z(n1845) );
  XOR U2025 ( .A(n1846), .B(n1847), .Z(n1843) );
  AND U2026 ( .A(n1848), .B(n1849), .Z(n1846) );
  XNOR U2027 ( .A(x[178]), .B(n1847), .Z(n1849) );
  XOR U2028 ( .A(n1850), .B(n1851), .Z(n1847) );
  AND U2029 ( .A(n1852), .B(n1853), .Z(n1850) );
  XNOR U2030 ( .A(x[177]), .B(n1851), .Z(n1853) );
  XOR U2031 ( .A(n1854), .B(n1855), .Z(n1851) );
  AND U2032 ( .A(n1856), .B(n1857), .Z(n1854) );
  XNOR U2033 ( .A(x[176]), .B(n1855), .Z(n1857) );
  XOR U2034 ( .A(n1858), .B(n1859), .Z(n1855) );
  AND U2035 ( .A(n1860), .B(n1861), .Z(n1858) );
  XNOR U2036 ( .A(x[175]), .B(n1859), .Z(n1861) );
  XOR U2037 ( .A(n1862), .B(n1863), .Z(n1859) );
  AND U2038 ( .A(n1864), .B(n1865), .Z(n1862) );
  XNOR U2039 ( .A(x[174]), .B(n1863), .Z(n1865) );
  XOR U2040 ( .A(n1866), .B(n1867), .Z(n1863) );
  AND U2041 ( .A(n1868), .B(n1869), .Z(n1866) );
  XNOR U2042 ( .A(x[173]), .B(n1867), .Z(n1869) );
  XOR U2043 ( .A(n1870), .B(n1871), .Z(n1867) );
  AND U2044 ( .A(n1872), .B(n1873), .Z(n1870) );
  XNOR U2045 ( .A(x[172]), .B(n1871), .Z(n1873) );
  XOR U2046 ( .A(n1874), .B(n1875), .Z(n1871) );
  AND U2047 ( .A(n1876), .B(n1877), .Z(n1874) );
  XNOR U2048 ( .A(x[171]), .B(n1875), .Z(n1877) );
  XOR U2049 ( .A(n1878), .B(n1879), .Z(n1875) );
  AND U2050 ( .A(n1880), .B(n1881), .Z(n1878) );
  XNOR U2051 ( .A(x[170]), .B(n1879), .Z(n1881) );
  XOR U2052 ( .A(n1882), .B(n1883), .Z(n1879) );
  AND U2053 ( .A(n1884), .B(n1885), .Z(n1882) );
  XNOR U2054 ( .A(x[169]), .B(n1883), .Z(n1885) );
  XOR U2055 ( .A(n1886), .B(n1887), .Z(n1883) );
  AND U2056 ( .A(n1888), .B(n1889), .Z(n1886) );
  XNOR U2057 ( .A(x[168]), .B(n1887), .Z(n1889) );
  XOR U2058 ( .A(n1890), .B(n1891), .Z(n1887) );
  AND U2059 ( .A(n1892), .B(n1893), .Z(n1890) );
  XNOR U2060 ( .A(x[167]), .B(n1891), .Z(n1893) );
  XOR U2061 ( .A(n1894), .B(n1895), .Z(n1891) );
  AND U2062 ( .A(n1896), .B(n1897), .Z(n1894) );
  XNOR U2063 ( .A(x[166]), .B(n1895), .Z(n1897) );
  XOR U2064 ( .A(n1898), .B(n1899), .Z(n1895) );
  AND U2065 ( .A(n1900), .B(n1901), .Z(n1898) );
  XNOR U2066 ( .A(x[165]), .B(n1899), .Z(n1901) );
  XOR U2067 ( .A(n1902), .B(n1903), .Z(n1899) );
  AND U2068 ( .A(n1904), .B(n1905), .Z(n1902) );
  XNOR U2069 ( .A(x[164]), .B(n1903), .Z(n1905) );
  XOR U2070 ( .A(n1906), .B(n1907), .Z(n1903) );
  AND U2071 ( .A(n1908), .B(n1909), .Z(n1906) );
  XNOR U2072 ( .A(x[163]), .B(n1907), .Z(n1909) );
  XOR U2073 ( .A(n1910), .B(n1911), .Z(n1907) );
  AND U2074 ( .A(n1912), .B(n1913), .Z(n1910) );
  XNOR U2075 ( .A(x[162]), .B(n1911), .Z(n1913) );
  XOR U2076 ( .A(n1914), .B(n1915), .Z(n1911) );
  AND U2077 ( .A(n1916), .B(n1917), .Z(n1914) );
  XNOR U2078 ( .A(x[161]), .B(n1915), .Z(n1917) );
  XOR U2079 ( .A(n1918), .B(n1919), .Z(n1915) );
  AND U2080 ( .A(n1920), .B(n1921), .Z(n1918) );
  XNOR U2081 ( .A(x[160]), .B(n1919), .Z(n1921) );
  XOR U2082 ( .A(n1922), .B(n1923), .Z(n1919) );
  AND U2083 ( .A(n1924), .B(n1925), .Z(n1922) );
  XNOR U2084 ( .A(x[159]), .B(n1923), .Z(n1925) );
  XOR U2085 ( .A(n1926), .B(n1927), .Z(n1923) );
  AND U2086 ( .A(n1928), .B(n1929), .Z(n1926) );
  XNOR U2087 ( .A(x[158]), .B(n1927), .Z(n1929) );
  XOR U2088 ( .A(n1930), .B(n1931), .Z(n1927) );
  AND U2089 ( .A(n1932), .B(n1933), .Z(n1930) );
  XNOR U2090 ( .A(x[157]), .B(n1931), .Z(n1933) );
  XOR U2091 ( .A(n1934), .B(n1935), .Z(n1931) );
  AND U2092 ( .A(n1936), .B(n1937), .Z(n1934) );
  XNOR U2093 ( .A(x[156]), .B(n1935), .Z(n1937) );
  XOR U2094 ( .A(n1938), .B(n1939), .Z(n1935) );
  AND U2095 ( .A(n1940), .B(n1941), .Z(n1938) );
  XNOR U2096 ( .A(x[155]), .B(n1939), .Z(n1941) );
  XOR U2097 ( .A(n1942), .B(n1943), .Z(n1939) );
  AND U2098 ( .A(n1944), .B(n1945), .Z(n1942) );
  XNOR U2099 ( .A(x[154]), .B(n1943), .Z(n1945) );
  XOR U2100 ( .A(n1946), .B(n1947), .Z(n1943) );
  AND U2101 ( .A(n1948), .B(n1949), .Z(n1946) );
  XNOR U2102 ( .A(x[153]), .B(n1947), .Z(n1949) );
  XOR U2103 ( .A(n1950), .B(n1951), .Z(n1947) );
  AND U2104 ( .A(n1952), .B(n1953), .Z(n1950) );
  XNOR U2105 ( .A(x[152]), .B(n1951), .Z(n1953) );
  XOR U2106 ( .A(n1954), .B(n1955), .Z(n1951) );
  AND U2107 ( .A(n1956), .B(n1957), .Z(n1954) );
  XNOR U2108 ( .A(x[151]), .B(n1955), .Z(n1957) );
  XOR U2109 ( .A(n1958), .B(n1959), .Z(n1955) );
  AND U2110 ( .A(n1960), .B(n1961), .Z(n1958) );
  XNOR U2111 ( .A(x[150]), .B(n1959), .Z(n1961) );
  XOR U2112 ( .A(n1962), .B(n1963), .Z(n1959) );
  AND U2113 ( .A(n1964), .B(n1965), .Z(n1962) );
  XNOR U2114 ( .A(x[149]), .B(n1963), .Z(n1965) );
  XOR U2115 ( .A(n1966), .B(n1967), .Z(n1963) );
  AND U2116 ( .A(n1968), .B(n1969), .Z(n1966) );
  XNOR U2117 ( .A(x[148]), .B(n1967), .Z(n1969) );
  XOR U2118 ( .A(n1970), .B(n1971), .Z(n1967) );
  AND U2119 ( .A(n1972), .B(n1973), .Z(n1970) );
  XNOR U2120 ( .A(x[147]), .B(n1971), .Z(n1973) );
  XOR U2121 ( .A(n1974), .B(n1975), .Z(n1971) );
  AND U2122 ( .A(n1976), .B(n1977), .Z(n1974) );
  XNOR U2123 ( .A(x[146]), .B(n1975), .Z(n1977) );
  XOR U2124 ( .A(n1978), .B(n1979), .Z(n1975) );
  AND U2125 ( .A(n1980), .B(n1981), .Z(n1978) );
  XNOR U2126 ( .A(x[145]), .B(n1979), .Z(n1981) );
  XOR U2127 ( .A(n1982), .B(n1983), .Z(n1979) );
  AND U2128 ( .A(n1984), .B(n1985), .Z(n1982) );
  XNOR U2129 ( .A(x[144]), .B(n1983), .Z(n1985) );
  XOR U2130 ( .A(n1986), .B(n1987), .Z(n1983) );
  AND U2131 ( .A(n1988), .B(n1989), .Z(n1986) );
  XNOR U2132 ( .A(x[143]), .B(n1987), .Z(n1989) );
  XOR U2133 ( .A(n1990), .B(n1991), .Z(n1987) );
  AND U2134 ( .A(n1992), .B(n1993), .Z(n1990) );
  XNOR U2135 ( .A(x[142]), .B(n1991), .Z(n1993) );
  XOR U2136 ( .A(n1994), .B(n1995), .Z(n1991) );
  AND U2137 ( .A(n1996), .B(n1997), .Z(n1994) );
  XNOR U2138 ( .A(x[141]), .B(n1995), .Z(n1997) );
  XOR U2139 ( .A(n1998), .B(n1999), .Z(n1995) );
  AND U2140 ( .A(n2000), .B(n2001), .Z(n1998) );
  XNOR U2141 ( .A(x[140]), .B(n1999), .Z(n2001) );
  XOR U2142 ( .A(n2002), .B(n2003), .Z(n1999) );
  AND U2143 ( .A(n2004), .B(n2005), .Z(n2002) );
  XNOR U2144 ( .A(x[139]), .B(n2003), .Z(n2005) );
  XOR U2145 ( .A(n2006), .B(n2007), .Z(n2003) );
  AND U2146 ( .A(n2008), .B(n2009), .Z(n2006) );
  XNOR U2147 ( .A(x[138]), .B(n2007), .Z(n2009) );
  XOR U2148 ( .A(n2010), .B(n2011), .Z(n2007) );
  AND U2149 ( .A(n2012), .B(n2013), .Z(n2010) );
  XNOR U2150 ( .A(x[137]), .B(n2011), .Z(n2013) );
  XOR U2151 ( .A(n2014), .B(n2015), .Z(n2011) );
  AND U2152 ( .A(n2016), .B(n2017), .Z(n2014) );
  XNOR U2153 ( .A(x[136]), .B(n2015), .Z(n2017) );
  XOR U2154 ( .A(n2018), .B(n2019), .Z(n2015) );
  AND U2155 ( .A(n2020), .B(n2021), .Z(n2018) );
  XNOR U2156 ( .A(x[135]), .B(n2019), .Z(n2021) );
  XOR U2157 ( .A(n2022), .B(n2023), .Z(n2019) );
  AND U2158 ( .A(n2024), .B(n2025), .Z(n2022) );
  XNOR U2159 ( .A(x[134]), .B(n2023), .Z(n2025) );
  XOR U2160 ( .A(n2026), .B(n2027), .Z(n2023) );
  AND U2161 ( .A(n2028), .B(n2029), .Z(n2026) );
  XNOR U2162 ( .A(x[133]), .B(n2027), .Z(n2029) );
  XOR U2163 ( .A(n2030), .B(n2031), .Z(n2027) );
  AND U2164 ( .A(n2032), .B(n2033), .Z(n2030) );
  XNOR U2165 ( .A(x[132]), .B(n2031), .Z(n2033) );
  XOR U2166 ( .A(n2034), .B(n2035), .Z(n2031) );
  AND U2167 ( .A(n2036), .B(n2037), .Z(n2034) );
  XNOR U2168 ( .A(x[131]), .B(n2035), .Z(n2037) );
  XOR U2169 ( .A(n2038), .B(n2039), .Z(n2035) );
  AND U2170 ( .A(n2040), .B(n2041), .Z(n2038) );
  XNOR U2171 ( .A(x[130]), .B(n2039), .Z(n2041) );
  XOR U2172 ( .A(n2042), .B(n2043), .Z(n2039) );
  AND U2173 ( .A(n2044), .B(n2045), .Z(n2042) );
  XNOR U2174 ( .A(x[129]), .B(n2043), .Z(n2045) );
  XOR U2175 ( .A(n2046), .B(n2047), .Z(n2043) );
  AND U2176 ( .A(n2048), .B(n2049), .Z(n2046) );
  XNOR U2177 ( .A(x[128]), .B(n2047), .Z(n2049) );
  XOR U2178 ( .A(n2050), .B(n2051), .Z(n2047) );
  AND U2179 ( .A(n2052), .B(n2053), .Z(n2050) );
  XNOR U2180 ( .A(x[127]), .B(n2051), .Z(n2053) );
  XOR U2181 ( .A(n2054), .B(n2055), .Z(n2051) );
  AND U2182 ( .A(n2056), .B(n2057), .Z(n2054) );
  XNOR U2183 ( .A(x[126]), .B(n2055), .Z(n2057) );
  XOR U2184 ( .A(n2058), .B(n2059), .Z(n2055) );
  AND U2185 ( .A(n2060), .B(n2061), .Z(n2058) );
  XNOR U2186 ( .A(x[125]), .B(n2059), .Z(n2061) );
  XOR U2187 ( .A(n2062), .B(n2063), .Z(n2059) );
  AND U2188 ( .A(n2064), .B(n2065), .Z(n2062) );
  XNOR U2189 ( .A(x[124]), .B(n2063), .Z(n2065) );
  XOR U2190 ( .A(n2066), .B(n2067), .Z(n2063) );
  AND U2191 ( .A(n2068), .B(n2069), .Z(n2066) );
  XNOR U2192 ( .A(x[123]), .B(n2067), .Z(n2069) );
  XOR U2193 ( .A(n2070), .B(n2071), .Z(n2067) );
  AND U2194 ( .A(n2072), .B(n2073), .Z(n2070) );
  XNOR U2195 ( .A(x[122]), .B(n2071), .Z(n2073) );
  XOR U2196 ( .A(n2074), .B(n2075), .Z(n2071) );
  AND U2197 ( .A(n2076), .B(n2077), .Z(n2074) );
  XNOR U2198 ( .A(x[121]), .B(n2075), .Z(n2077) );
  XOR U2199 ( .A(n2078), .B(n2079), .Z(n2075) );
  AND U2200 ( .A(n2080), .B(n2081), .Z(n2078) );
  XNOR U2201 ( .A(x[120]), .B(n2079), .Z(n2081) );
  XOR U2202 ( .A(n2082), .B(n2083), .Z(n2079) );
  AND U2203 ( .A(n2084), .B(n2085), .Z(n2082) );
  XNOR U2204 ( .A(x[119]), .B(n2083), .Z(n2085) );
  XOR U2205 ( .A(n2086), .B(n2087), .Z(n2083) );
  AND U2206 ( .A(n2088), .B(n2089), .Z(n2086) );
  XNOR U2207 ( .A(x[118]), .B(n2087), .Z(n2089) );
  XOR U2208 ( .A(n2090), .B(n2091), .Z(n2087) );
  AND U2209 ( .A(n2092), .B(n2093), .Z(n2090) );
  XNOR U2210 ( .A(x[117]), .B(n2091), .Z(n2093) );
  XOR U2211 ( .A(n2094), .B(n2095), .Z(n2091) );
  AND U2212 ( .A(n2096), .B(n2097), .Z(n2094) );
  XNOR U2213 ( .A(x[116]), .B(n2095), .Z(n2097) );
  XOR U2214 ( .A(n2098), .B(n2099), .Z(n2095) );
  AND U2215 ( .A(n2100), .B(n2101), .Z(n2098) );
  XNOR U2216 ( .A(x[115]), .B(n2099), .Z(n2101) );
  XOR U2217 ( .A(n2102), .B(n2103), .Z(n2099) );
  AND U2218 ( .A(n2104), .B(n2105), .Z(n2102) );
  XNOR U2219 ( .A(x[114]), .B(n2103), .Z(n2105) );
  XOR U2220 ( .A(n2106), .B(n2107), .Z(n2103) );
  AND U2221 ( .A(n2108), .B(n2109), .Z(n2106) );
  XNOR U2222 ( .A(x[113]), .B(n2107), .Z(n2109) );
  XOR U2223 ( .A(n2110), .B(n2111), .Z(n2107) );
  AND U2224 ( .A(n2112), .B(n2113), .Z(n2110) );
  XNOR U2225 ( .A(x[112]), .B(n2111), .Z(n2113) );
  XOR U2226 ( .A(n2114), .B(n2115), .Z(n2111) );
  AND U2227 ( .A(n2116), .B(n2117), .Z(n2114) );
  XNOR U2228 ( .A(x[111]), .B(n2115), .Z(n2117) );
  XOR U2229 ( .A(n2118), .B(n2119), .Z(n2115) );
  AND U2230 ( .A(n2120), .B(n2121), .Z(n2118) );
  XNOR U2231 ( .A(x[110]), .B(n2119), .Z(n2121) );
  XOR U2232 ( .A(n2122), .B(n2123), .Z(n2119) );
  AND U2233 ( .A(n2124), .B(n2125), .Z(n2122) );
  XNOR U2234 ( .A(x[109]), .B(n2123), .Z(n2125) );
  XOR U2235 ( .A(n2126), .B(n2127), .Z(n2123) );
  AND U2236 ( .A(n2128), .B(n2129), .Z(n2126) );
  XNOR U2237 ( .A(x[108]), .B(n2127), .Z(n2129) );
  XOR U2238 ( .A(n2130), .B(n2131), .Z(n2127) );
  AND U2239 ( .A(n2132), .B(n2133), .Z(n2130) );
  XNOR U2240 ( .A(x[107]), .B(n2131), .Z(n2133) );
  XOR U2241 ( .A(n2134), .B(n2135), .Z(n2131) );
  AND U2242 ( .A(n2136), .B(n2137), .Z(n2134) );
  XNOR U2243 ( .A(x[106]), .B(n2135), .Z(n2137) );
  XOR U2244 ( .A(n2138), .B(n2139), .Z(n2135) );
  AND U2245 ( .A(n2140), .B(n2141), .Z(n2138) );
  XNOR U2246 ( .A(x[105]), .B(n2139), .Z(n2141) );
  XOR U2247 ( .A(n2142), .B(n2143), .Z(n2139) );
  AND U2248 ( .A(n2144), .B(n2145), .Z(n2142) );
  XNOR U2249 ( .A(x[104]), .B(n2143), .Z(n2145) );
  XOR U2250 ( .A(n2146), .B(n2147), .Z(n2143) );
  AND U2251 ( .A(n2148), .B(n2149), .Z(n2146) );
  XNOR U2252 ( .A(x[103]), .B(n2147), .Z(n2149) );
  XOR U2253 ( .A(n2150), .B(n2151), .Z(n2147) );
  AND U2254 ( .A(n2152), .B(n2153), .Z(n2150) );
  XNOR U2255 ( .A(x[102]), .B(n2151), .Z(n2153) );
  XOR U2256 ( .A(n2154), .B(n2155), .Z(n2151) );
  AND U2257 ( .A(n2156), .B(n2157), .Z(n2154) );
  XNOR U2258 ( .A(x[101]), .B(n2155), .Z(n2157) );
  XOR U2259 ( .A(n2158), .B(n2159), .Z(n2155) );
  AND U2260 ( .A(n2160), .B(n2161), .Z(n2158) );
  XNOR U2261 ( .A(x[100]), .B(n2159), .Z(n2161) );
  XOR U2262 ( .A(n2162), .B(n2163), .Z(n2159) );
  AND U2263 ( .A(n2164), .B(n2165), .Z(n2162) );
  XNOR U2264 ( .A(x[99]), .B(n2163), .Z(n2165) );
  XOR U2265 ( .A(n2166), .B(n2167), .Z(n2163) );
  AND U2266 ( .A(n2168), .B(n2169), .Z(n2166) );
  XNOR U2267 ( .A(x[98]), .B(n2167), .Z(n2169) );
  XOR U2268 ( .A(n2170), .B(n2171), .Z(n2167) );
  AND U2269 ( .A(n2172), .B(n2173), .Z(n2170) );
  XNOR U2270 ( .A(x[97]), .B(n2171), .Z(n2173) );
  XOR U2271 ( .A(n2174), .B(n2175), .Z(n2171) );
  AND U2272 ( .A(n2176), .B(n2177), .Z(n2174) );
  XNOR U2273 ( .A(x[96]), .B(n2175), .Z(n2177) );
  XOR U2274 ( .A(n2178), .B(n2179), .Z(n2175) );
  AND U2275 ( .A(n2180), .B(n2181), .Z(n2178) );
  XNOR U2276 ( .A(x[95]), .B(n2179), .Z(n2181) );
  XOR U2277 ( .A(n2182), .B(n2183), .Z(n2179) );
  AND U2278 ( .A(n2184), .B(n2185), .Z(n2182) );
  XNOR U2279 ( .A(x[94]), .B(n2183), .Z(n2185) );
  XOR U2280 ( .A(n2186), .B(n2187), .Z(n2183) );
  AND U2281 ( .A(n2188), .B(n2189), .Z(n2186) );
  XNOR U2282 ( .A(x[93]), .B(n2187), .Z(n2189) );
  XOR U2283 ( .A(n2190), .B(n2191), .Z(n2187) );
  AND U2284 ( .A(n2192), .B(n2193), .Z(n2190) );
  XNOR U2285 ( .A(x[92]), .B(n2191), .Z(n2193) );
  XOR U2286 ( .A(n2194), .B(n2195), .Z(n2191) );
  AND U2287 ( .A(n2196), .B(n2197), .Z(n2194) );
  XNOR U2288 ( .A(x[91]), .B(n2195), .Z(n2197) );
  XOR U2289 ( .A(n2198), .B(n2199), .Z(n2195) );
  AND U2290 ( .A(n2200), .B(n2201), .Z(n2198) );
  XNOR U2291 ( .A(x[90]), .B(n2199), .Z(n2201) );
  XOR U2292 ( .A(n2202), .B(n2203), .Z(n2199) );
  AND U2293 ( .A(n2204), .B(n2205), .Z(n2202) );
  XNOR U2294 ( .A(x[89]), .B(n2203), .Z(n2205) );
  XOR U2295 ( .A(n2206), .B(n2207), .Z(n2203) );
  AND U2296 ( .A(n2208), .B(n2209), .Z(n2206) );
  XNOR U2297 ( .A(x[88]), .B(n2207), .Z(n2209) );
  XOR U2298 ( .A(n2210), .B(n2211), .Z(n2207) );
  AND U2299 ( .A(n2212), .B(n2213), .Z(n2210) );
  XNOR U2300 ( .A(x[87]), .B(n2211), .Z(n2213) );
  XOR U2301 ( .A(n2214), .B(n2215), .Z(n2211) );
  AND U2302 ( .A(n2216), .B(n2217), .Z(n2214) );
  XNOR U2303 ( .A(x[86]), .B(n2215), .Z(n2217) );
  XOR U2304 ( .A(n2218), .B(n2219), .Z(n2215) );
  AND U2305 ( .A(n2220), .B(n2221), .Z(n2218) );
  XNOR U2306 ( .A(x[85]), .B(n2219), .Z(n2221) );
  XOR U2307 ( .A(n2222), .B(n2223), .Z(n2219) );
  AND U2308 ( .A(n2224), .B(n2225), .Z(n2222) );
  XNOR U2309 ( .A(x[84]), .B(n2223), .Z(n2225) );
  XOR U2310 ( .A(n2226), .B(n2227), .Z(n2223) );
  AND U2311 ( .A(n2228), .B(n2229), .Z(n2226) );
  XNOR U2312 ( .A(x[83]), .B(n2227), .Z(n2229) );
  XOR U2313 ( .A(n2230), .B(n2231), .Z(n2227) );
  AND U2314 ( .A(n2232), .B(n2233), .Z(n2230) );
  XNOR U2315 ( .A(x[82]), .B(n2231), .Z(n2233) );
  XOR U2316 ( .A(n2234), .B(n2235), .Z(n2231) );
  AND U2317 ( .A(n2236), .B(n2237), .Z(n2234) );
  XNOR U2318 ( .A(x[81]), .B(n2235), .Z(n2237) );
  XOR U2319 ( .A(n2238), .B(n2239), .Z(n2235) );
  AND U2320 ( .A(n2240), .B(n2241), .Z(n2238) );
  XNOR U2321 ( .A(x[80]), .B(n2239), .Z(n2241) );
  XOR U2322 ( .A(n2242), .B(n2243), .Z(n2239) );
  AND U2323 ( .A(n2244), .B(n2245), .Z(n2242) );
  XNOR U2324 ( .A(x[79]), .B(n2243), .Z(n2245) );
  XOR U2325 ( .A(n2246), .B(n2247), .Z(n2243) );
  AND U2326 ( .A(n2248), .B(n2249), .Z(n2246) );
  XNOR U2327 ( .A(x[78]), .B(n2247), .Z(n2249) );
  XOR U2328 ( .A(n2250), .B(n2251), .Z(n2247) );
  AND U2329 ( .A(n2252), .B(n2253), .Z(n2250) );
  XNOR U2330 ( .A(x[77]), .B(n2251), .Z(n2253) );
  XOR U2331 ( .A(n2254), .B(n2255), .Z(n2251) );
  AND U2332 ( .A(n2256), .B(n2257), .Z(n2254) );
  XNOR U2333 ( .A(x[76]), .B(n2255), .Z(n2257) );
  XOR U2334 ( .A(n2258), .B(n2259), .Z(n2255) );
  AND U2335 ( .A(n2260), .B(n2261), .Z(n2258) );
  XNOR U2336 ( .A(x[75]), .B(n2259), .Z(n2261) );
  XOR U2337 ( .A(n2262), .B(n2263), .Z(n2259) );
  AND U2338 ( .A(n2264), .B(n2265), .Z(n2262) );
  XNOR U2339 ( .A(x[74]), .B(n2263), .Z(n2265) );
  XOR U2340 ( .A(n2266), .B(n2267), .Z(n2263) );
  AND U2341 ( .A(n2268), .B(n2269), .Z(n2266) );
  XNOR U2342 ( .A(x[73]), .B(n2267), .Z(n2269) );
  XOR U2343 ( .A(n2270), .B(n2271), .Z(n2267) );
  AND U2344 ( .A(n2272), .B(n2273), .Z(n2270) );
  XNOR U2345 ( .A(x[72]), .B(n2271), .Z(n2273) );
  XOR U2346 ( .A(n2274), .B(n2275), .Z(n2271) );
  AND U2347 ( .A(n2276), .B(n2277), .Z(n2274) );
  XNOR U2348 ( .A(x[71]), .B(n2275), .Z(n2277) );
  XOR U2349 ( .A(n2278), .B(n2279), .Z(n2275) );
  AND U2350 ( .A(n2280), .B(n2281), .Z(n2278) );
  XNOR U2351 ( .A(x[70]), .B(n2279), .Z(n2281) );
  XOR U2352 ( .A(n2282), .B(n2283), .Z(n2279) );
  AND U2353 ( .A(n2284), .B(n2285), .Z(n2282) );
  XNOR U2354 ( .A(x[69]), .B(n2283), .Z(n2285) );
  XOR U2355 ( .A(n2286), .B(n2287), .Z(n2283) );
  AND U2356 ( .A(n2288), .B(n2289), .Z(n2286) );
  XNOR U2357 ( .A(x[68]), .B(n2287), .Z(n2289) );
  XOR U2358 ( .A(n2290), .B(n2291), .Z(n2287) );
  AND U2359 ( .A(n2292), .B(n2293), .Z(n2290) );
  XNOR U2360 ( .A(x[67]), .B(n2291), .Z(n2293) );
  XOR U2361 ( .A(n2294), .B(n2295), .Z(n2291) );
  AND U2362 ( .A(n2296), .B(n2297), .Z(n2294) );
  XNOR U2363 ( .A(x[66]), .B(n2295), .Z(n2297) );
  XOR U2364 ( .A(n2298), .B(n2299), .Z(n2295) );
  AND U2365 ( .A(n2300), .B(n2301), .Z(n2298) );
  XNOR U2366 ( .A(x[65]), .B(n2299), .Z(n2301) );
  XOR U2367 ( .A(n2302), .B(n2303), .Z(n2299) );
  AND U2368 ( .A(n2304), .B(n2305), .Z(n2302) );
  XNOR U2369 ( .A(x[64]), .B(n2303), .Z(n2305) );
  XOR U2370 ( .A(n2306), .B(n2307), .Z(n2303) );
  AND U2371 ( .A(n2308), .B(n2309), .Z(n2306) );
  XNOR U2372 ( .A(x[63]), .B(n2307), .Z(n2309) );
  XOR U2373 ( .A(n2310), .B(n2311), .Z(n2307) );
  AND U2374 ( .A(n2312), .B(n2313), .Z(n2310) );
  XNOR U2375 ( .A(x[62]), .B(n2311), .Z(n2313) );
  XOR U2376 ( .A(n2314), .B(n2315), .Z(n2311) );
  AND U2377 ( .A(n2316), .B(n2317), .Z(n2314) );
  XNOR U2378 ( .A(x[61]), .B(n2315), .Z(n2317) );
  XOR U2379 ( .A(n2318), .B(n2319), .Z(n2315) );
  AND U2380 ( .A(n2320), .B(n2321), .Z(n2318) );
  XNOR U2381 ( .A(x[60]), .B(n2319), .Z(n2321) );
  XOR U2382 ( .A(n2322), .B(n2323), .Z(n2319) );
  AND U2383 ( .A(n2324), .B(n2325), .Z(n2322) );
  XNOR U2384 ( .A(x[59]), .B(n2323), .Z(n2325) );
  XOR U2385 ( .A(n2326), .B(n2327), .Z(n2323) );
  AND U2386 ( .A(n2328), .B(n2329), .Z(n2326) );
  XNOR U2387 ( .A(x[58]), .B(n2327), .Z(n2329) );
  XOR U2388 ( .A(n2330), .B(n2331), .Z(n2327) );
  AND U2389 ( .A(n2332), .B(n2333), .Z(n2330) );
  XNOR U2390 ( .A(x[57]), .B(n2331), .Z(n2333) );
  XOR U2391 ( .A(n2334), .B(n2335), .Z(n2331) );
  AND U2392 ( .A(n2336), .B(n2337), .Z(n2334) );
  XNOR U2393 ( .A(x[56]), .B(n2335), .Z(n2337) );
  XOR U2394 ( .A(n2338), .B(n2339), .Z(n2335) );
  AND U2395 ( .A(n2340), .B(n2341), .Z(n2338) );
  XNOR U2396 ( .A(x[55]), .B(n2339), .Z(n2341) );
  XOR U2397 ( .A(n2342), .B(n2343), .Z(n2339) );
  AND U2398 ( .A(n2344), .B(n2345), .Z(n2342) );
  XNOR U2399 ( .A(x[54]), .B(n2343), .Z(n2345) );
  XOR U2400 ( .A(n2346), .B(n2347), .Z(n2343) );
  AND U2401 ( .A(n2348), .B(n2349), .Z(n2346) );
  XNOR U2402 ( .A(x[53]), .B(n2347), .Z(n2349) );
  XOR U2403 ( .A(n2350), .B(n2351), .Z(n2347) );
  AND U2404 ( .A(n2352), .B(n2353), .Z(n2350) );
  XNOR U2405 ( .A(x[52]), .B(n2351), .Z(n2353) );
  XOR U2406 ( .A(n2354), .B(n2355), .Z(n2351) );
  AND U2407 ( .A(n2356), .B(n2357), .Z(n2354) );
  XNOR U2408 ( .A(x[51]), .B(n2355), .Z(n2357) );
  XOR U2409 ( .A(n2358), .B(n2359), .Z(n2355) );
  AND U2410 ( .A(n2360), .B(n2361), .Z(n2358) );
  XNOR U2411 ( .A(x[50]), .B(n2359), .Z(n2361) );
  XOR U2412 ( .A(n2362), .B(n2363), .Z(n2359) );
  AND U2413 ( .A(n2364), .B(n2365), .Z(n2362) );
  XNOR U2414 ( .A(x[49]), .B(n2363), .Z(n2365) );
  XOR U2415 ( .A(n2366), .B(n2367), .Z(n2363) );
  AND U2416 ( .A(n2368), .B(n2369), .Z(n2366) );
  XNOR U2417 ( .A(x[48]), .B(n2367), .Z(n2369) );
  XOR U2418 ( .A(n2370), .B(n2371), .Z(n2367) );
  AND U2419 ( .A(n2372), .B(n2373), .Z(n2370) );
  XNOR U2420 ( .A(x[47]), .B(n2371), .Z(n2373) );
  XOR U2421 ( .A(n2374), .B(n2375), .Z(n2371) );
  AND U2422 ( .A(n2376), .B(n2377), .Z(n2374) );
  XNOR U2423 ( .A(x[46]), .B(n2375), .Z(n2377) );
  XOR U2424 ( .A(n2378), .B(n2379), .Z(n2375) );
  AND U2425 ( .A(n2380), .B(n2381), .Z(n2378) );
  XNOR U2426 ( .A(x[45]), .B(n2379), .Z(n2381) );
  XOR U2427 ( .A(n2382), .B(n2383), .Z(n2379) );
  AND U2428 ( .A(n2384), .B(n2385), .Z(n2382) );
  XNOR U2429 ( .A(x[44]), .B(n2383), .Z(n2385) );
  XOR U2430 ( .A(n2386), .B(n2387), .Z(n2383) );
  AND U2431 ( .A(n2388), .B(n2389), .Z(n2386) );
  XNOR U2432 ( .A(x[43]), .B(n2387), .Z(n2389) );
  XOR U2433 ( .A(n2390), .B(n2391), .Z(n2387) );
  AND U2434 ( .A(n2392), .B(n2393), .Z(n2390) );
  XNOR U2435 ( .A(x[42]), .B(n2391), .Z(n2393) );
  XOR U2436 ( .A(n2394), .B(n2395), .Z(n2391) );
  AND U2437 ( .A(n2396), .B(n2397), .Z(n2394) );
  XNOR U2438 ( .A(x[41]), .B(n2395), .Z(n2397) );
  XOR U2439 ( .A(n2398), .B(n2399), .Z(n2395) );
  AND U2440 ( .A(n2400), .B(n2401), .Z(n2398) );
  XNOR U2441 ( .A(x[40]), .B(n2399), .Z(n2401) );
  XOR U2442 ( .A(n2402), .B(n2403), .Z(n2399) );
  AND U2443 ( .A(n2404), .B(n2405), .Z(n2402) );
  XNOR U2444 ( .A(x[39]), .B(n2403), .Z(n2405) );
  XOR U2445 ( .A(n2406), .B(n2407), .Z(n2403) );
  AND U2446 ( .A(n2408), .B(n2409), .Z(n2406) );
  XNOR U2447 ( .A(x[38]), .B(n2407), .Z(n2409) );
  XOR U2448 ( .A(n2410), .B(n2411), .Z(n2407) );
  AND U2449 ( .A(n2412), .B(n2413), .Z(n2410) );
  XNOR U2450 ( .A(x[37]), .B(n2411), .Z(n2413) );
  XOR U2451 ( .A(n2414), .B(n2415), .Z(n2411) );
  AND U2452 ( .A(n2416), .B(n2417), .Z(n2414) );
  XNOR U2453 ( .A(x[36]), .B(n2415), .Z(n2417) );
  XOR U2454 ( .A(n2418), .B(n2419), .Z(n2415) );
  AND U2455 ( .A(n2420), .B(n2421), .Z(n2418) );
  XNOR U2456 ( .A(x[35]), .B(n2419), .Z(n2421) );
  XOR U2457 ( .A(n2422), .B(n2423), .Z(n2419) );
  AND U2458 ( .A(n2424), .B(n2425), .Z(n2422) );
  XNOR U2459 ( .A(x[34]), .B(n2423), .Z(n2425) );
  XOR U2460 ( .A(n2426), .B(n2427), .Z(n2423) );
  AND U2461 ( .A(n2428), .B(n2429), .Z(n2426) );
  XNOR U2462 ( .A(x[33]), .B(n2427), .Z(n2429) );
  XOR U2463 ( .A(n2430), .B(n2431), .Z(n2427) );
  AND U2464 ( .A(n2432), .B(n2433), .Z(n2430) );
  XNOR U2465 ( .A(x[32]), .B(n2431), .Z(n2433) );
  XOR U2466 ( .A(n2434), .B(n2435), .Z(n2431) );
  AND U2467 ( .A(n2436), .B(n2437), .Z(n2434) );
  XNOR U2468 ( .A(x[31]), .B(n2435), .Z(n2437) );
  XOR U2469 ( .A(n2438), .B(n2439), .Z(n2435) );
  AND U2470 ( .A(n2440), .B(n2441), .Z(n2438) );
  XNOR U2471 ( .A(x[30]), .B(n2439), .Z(n2441) );
  XOR U2472 ( .A(n2442), .B(n2443), .Z(n2439) );
  AND U2473 ( .A(n2444), .B(n2445), .Z(n2442) );
  XNOR U2474 ( .A(x[29]), .B(n2443), .Z(n2445) );
  XOR U2475 ( .A(n2446), .B(n2447), .Z(n2443) );
  AND U2476 ( .A(n2448), .B(n2449), .Z(n2446) );
  XNOR U2477 ( .A(x[28]), .B(n2447), .Z(n2449) );
  XOR U2478 ( .A(n2450), .B(n2451), .Z(n2447) );
  AND U2479 ( .A(n2452), .B(n2453), .Z(n2450) );
  XNOR U2480 ( .A(x[27]), .B(n2451), .Z(n2453) );
  XOR U2481 ( .A(n2454), .B(n2455), .Z(n2451) );
  AND U2482 ( .A(n2456), .B(n2457), .Z(n2454) );
  XNOR U2483 ( .A(x[26]), .B(n2455), .Z(n2457) );
  XOR U2484 ( .A(n2458), .B(n2459), .Z(n2455) );
  AND U2485 ( .A(n2460), .B(n2461), .Z(n2458) );
  XNOR U2486 ( .A(x[25]), .B(n2459), .Z(n2461) );
  XOR U2487 ( .A(n2462), .B(n2463), .Z(n2459) );
  AND U2488 ( .A(n2464), .B(n2465), .Z(n2462) );
  XNOR U2489 ( .A(x[24]), .B(n2463), .Z(n2465) );
  XOR U2490 ( .A(n2466), .B(n2467), .Z(n2463) );
  AND U2491 ( .A(n2468), .B(n2469), .Z(n2466) );
  XNOR U2492 ( .A(x[23]), .B(n2467), .Z(n2469) );
  XOR U2493 ( .A(n2470), .B(n2471), .Z(n2467) );
  AND U2494 ( .A(n2472), .B(n2473), .Z(n2470) );
  XNOR U2495 ( .A(x[22]), .B(n2471), .Z(n2473) );
  XOR U2496 ( .A(n2474), .B(n2475), .Z(n2471) );
  AND U2497 ( .A(n2476), .B(n2477), .Z(n2474) );
  XNOR U2498 ( .A(x[21]), .B(n2475), .Z(n2477) );
  XOR U2499 ( .A(n2478), .B(n2479), .Z(n2475) );
  AND U2500 ( .A(n2480), .B(n2481), .Z(n2478) );
  XNOR U2501 ( .A(x[20]), .B(n2479), .Z(n2481) );
  XOR U2502 ( .A(n2482), .B(n2483), .Z(n2479) );
  AND U2503 ( .A(n2484), .B(n2485), .Z(n2482) );
  XNOR U2504 ( .A(x[19]), .B(n2483), .Z(n2485) );
  XOR U2505 ( .A(n2486), .B(n2487), .Z(n2483) );
  AND U2506 ( .A(n2488), .B(n2489), .Z(n2486) );
  XNOR U2507 ( .A(x[18]), .B(n2487), .Z(n2489) );
  XOR U2508 ( .A(n2490), .B(n2491), .Z(n2487) );
  AND U2509 ( .A(n2492), .B(n2493), .Z(n2490) );
  XNOR U2510 ( .A(x[17]), .B(n2491), .Z(n2493) );
  XOR U2511 ( .A(n2494), .B(n2495), .Z(n2491) );
  AND U2512 ( .A(n2496), .B(n2497), .Z(n2494) );
  XNOR U2513 ( .A(x[16]), .B(n2495), .Z(n2497) );
  XOR U2514 ( .A(n2498), .B(n2499), .Z(n2495) );
  AND U2515 ( .A(n2500), .B(n2501), .Z(n2498) );
  XNOR U2516 ( .A(x[15]), .B(n2499), .Z(n2501) );
  XOR U2517 ( .A(n2502), .B(n2503), .Z(n2499) );
  AND U2518 ( .A(n2504), .B(n2505), .Z(n2502) );
  XNOR U2519 ( .A(x[14]), .B(n2503), .Z(n2505) );
  XOR U2520 ( .A(n2506), .B(n2507), .Z(n2503) );
  AND U2521 ( .A(n2508), .B(n2509), .Z(n2506) );
  XNOR U2522 ( .A(x[13]), .B(n2507), .Z(n2509) );
  XOR U2523 ( .A(n2510), .B(n2511), .Z(n2507) );
  AND U2524 ( .A(n2512), .B(n2513), .Z(n2510) );
  XNOR U2525 ( .A(x[12]), .B(n2511), .Z(n2513) );
  XOR U2526 ( .A(n2514), .B(n2515), .Z(n2511) );
  AND U2527 ( .A(n2516), .B(n2517), .Z(n2514) );
  XNOR U2528 ( .A(x[11]), .B(n2515), .Z(n2517) );
  XOR U2529 ( .A(n2518), .B(n2519), .Z(n2515) );
  AND U2530 ( .A(n2520), .B(n2521), .Z(n2518) );
  XNOR U2531 ( .A(x[10]), .B(n2519), .Z(n2521) );
  XOR U2532 ( .A(n2522), .B(n2523), .Z(n2519) );
  AND U2533 ( .A(n2524), .B(n2525), .Z(n2522) );
  XNOR U2534 ( .A(x[9]), .B(n2523), .Z(n2525) );
  XOR U2535 ( .A(n2526), .B(n2527), .Z(n2523) );
  AND U2536 ( .A(n2528), .B(n2529), .Z(n2526) );
  XNOR U2537 ( .A(x[8]), .B(n2527), .Z(n2529) );
  XOR U2538 ( .A(n2530), .B(n2531), .Z(n2527) );
  AND U2539 ( .A(n2532), .B(n2533), .Z(n2530) );
  XNOR U2540 ( .A(x[7]), .B(n2531), .Z(n2533) );
  XOR U2541 ( .A(n2534), .B(n2535), .Z(n2531) );
  AND U2542 ( .A(n2536), .B(n2537), .Z(n2534) );
  XNOR U2543 ( .A(x[6]), .B(n2535), .Z(n2537) );
  XOR U2544 ( .A(n2538), .B(n2539), .Z(n2535) );
  AND U2545 ( .A(n2540), .B(n2541), .Z(n2538) );
  XNOR U2546 ( .A(x[5]), .B(n2539), .Z(n2541) );
  XOR U2547 ( .A(n2542), .B(n2543), .Z(n2539) );
  AND U2548 ( .A(n2544), .B(n2545), .Z(n2542) );
  XNOR U2549 ( .A(x[4]), .B(n2543), .Z(n2545) );
  XOR U2550 ( .A(n2546), .B(n2547), .Z(n2543) );
  AND U2551 ( .A(n2548), .B(n2549), .Z(n2546) );
  XNOR U2552 ( .A(x[3]), .B(n2547), .Z(n2549) );
  XOR U2553 ( .A(n2550), .B(n2551), .Z(n2547) );
  AND U2554 ( .A(n2552), .B(n2553), .Z(n2550) );
  XNOR U2555 ( .A(x[2]), .B(n2551), .Z(n2553) );
  XOR U2556 ( .A(n2554), .B(n2555), .Z(n2551) );
  AND U2557 ( .A(n2556), .B(n2557), .Z(n2554) );
  XNOR U2558 ( .A(x[1]), .B(n2555), .Z(n2557) );
  XOR U2559 ( .A(y[1]), .B(n2555), .Z(n2556) );
  XOR U2560 ( .A(ci), .B(n2558), .Z(n2555) );
  NANDN U2561 ( .A(n2559), .B(n2560), .Z(n2558) );
  XOR U2562 ( .A(x[0]), .B(ci), .Z(n2560) );
  XOR U2563 ( .A(y[0]), .B(ci), .Z(n2559) );
endmodule

