
module round_0 ( in, round_const, out );
  input [1599:0] in;
  input [63:0] round_const;
  output [1599:0] out;
  wire   round_const_63, round_const_31, round_const_15, round_const_7,
         round_const_3, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614;
  assign round_const_63 = round_const[63];
  assign round_const_31 = round_const[31];
  assign round_const_15 = round_const[15];
  assign round_const_7 = round_const[7];
  assign round_const_3 = round_const[3];

  XOR U1 ( .A(in[1469]), .B(in[509]), .Z(n4809) );
  XNOR U2 ( .A(in[829]), .B(in[189]), .Z(n4808) );
  XNOR U3 ( .A(n4809), .B(n4808), .Z(n4810) );
  XOR U4 ( .A(in[1149]), .B(n4810), .Z(n5679) );
  XOR U5 ( .A(in[1598]), .B(in[638]), .Z(n4812) );
  XNOR U6 ( .A(in[958]), .B(in[318]), .Z(n4811) );
  XNOR U7 ( .A(n4812), .B(n4811), .Z(n4813) );
  XOR U8 ( .A(in[1278]), .B(n4813), .Z(n6280) );
  XNOR U9 ( .A(n5679), .B(n6280), .Z(n8622) );
  XNOR U10 ( .A(in[254]), .B(n8622), .Z(n8384) );
  XOR U11 ( .A(in[1345]), .B(in[65]), .Z(n4815) );
  XNOR U12 ( .A(in[1025]), .B(in[385]), .Z(n4814) );
  XNOR U13 ( .A(n4815), .B(n4814), .Z(n4816) );
  XOR U14 ( .A(in[705]), .B(n4816), .Z(n6288) );
  XOR U15 ( .A(in[1474]), .B(in[514]), .Z(n4818) );
  XNOR U16 ( .A(in[834]), .B(in[194]), .Z(n4817) );
  XNOR U17 ( .A(n4818), .B(n4817), .Z(n4819) );
  XNOR U18 ( .A(in[1154]), .B(n4819), .Z(n5995) );
  XNOR U19 ( .A(n6288), .B(n5995), .Z(n8377) );
  XNOR U20 ( .A(in[1410]), .B(n8377), .Z(n8383) );
  XOR U21 ( .A(in[137]), .B(in[457]), .Z(n4821) );
  XNOR U22 ( .A(in[777]), .B(in[1417]), .Z(n4820) );
  XNOR U23 ( .A(n4821), .B(n4820), .Z(n4822) );
  XOR U24 ( .A(in[1097]), .B(n4822), .Z(n5948) );
  XOR U25 ( .A(in[328]), .B(in[8]), .Z(n4824) );
  XNOR U26 ( .A(in[968]), .B(in[648]), .Z(n4823) );
  XNOR U27 ( .A(n4824), .B(n4823), .Z(n4825) );
  XOR U28 ( .A(in[1288]), .B(n4825), .Z(n6016) );
  XNOR U29 ( .A(n5948), .B(n6016), .Z(n8893) );
  XNOR U30 ( .A(in[1033]), .B(n8893), .Z(n7416) );
  NAND U31 ( .A(n8383), .B(n7416), .Z(n4826) );
  XNOR U32 ( .A(n8384), .B(n4826), .Z(out[0]) );
  XOR U33 ( .A(in[1386]), .B(in[106]), .Z(n4828) );
  XNOR U34 ( .A(in[1066]), .B(in[746]), .Z(n4827) );
  XNOR U35 ( .A(n4828), .B(n4827), .Z(n4829) );
  XOR U36 ( .A(in[426]), .B(n4829), .Z(n5282) );
  XOR U37 ( .A(in[1515]), .B(in[555]), .Z(n4831) );
  XNOR U38 ( .A(in[875]), .B(in[235]), .Z(n4830) );
  XNOR U39 ( .A(n4831), .B(n4830), .Z(n4832) );
  XOR U40 ( .A(in[1195]), .B(n4832), .Z(n6136) );
  XNOR U41 ( .A(n5282), .B(n6136), .Z(n8557) );
  XNOR U42 ( .A(in[171]), .B(n8557), .Z(n6108) );
  XOR U43 ( .A(in[971]), .B(in[1291]), .Z(n4834) );
  XNOR U44 ( .A(in[11]), .B(in[331]), .Z(n4833) );
  XNOR U45 ( .A(n4834), .B(n4833), .Z(n4835) );
  XOR U46 ( .A(in[651]), .B(n4835), .Z(n6027) );
  XOR U47 ( .A(in[140]), .B(in[460]), .Z(n4837) );
  XNOR U48 ( .A(in[1100]), .B(in[1420]), .Z(n4836) );
  XNOR U49 ( .A(n4837), .B(n4836), .Z(n4838) );
  XNOR U50 ( .A(in[780]), .B(n4838), .Z(n5966) );
  XNOR U51 ( .A(n6027), .B(n5966), .Z(n8902) );
  XNOR U52 ( .A(in[1356]), .B(n8902), .Z(n6503) );
  XOR U53 ( .A(in[1364]), .B(in[724]), .Z(n4840) );
  XNOR U54 ( .A(in[84]), .B(in[404]), .Z(n4839) );
  XNOR U55 ( .A(n4840), .B(n4839), .Z(n4841) );
  XOR U56 ( .A(in[1044]), .B(n4841), .Z(n5584) );
  XOR U57 ( .A(in[1555]), .B(in[595]), .Z(n4843) );
  XNOR U58 ( .A(in[915]), .B(in[275]), .Z(n4842) );
  XNOR U59 ( .A(n4843), .B(n4842), .Z(n4844) );
  XOR U60 ( .A(in[1235]), .B(n4844), .Z(n5296) );
  XNOR U61 ( .A(n5584), .B(n5296), .Z(n8689) );
  XNOR U62 ( .A(in[980]), .B(n8689), .Z(n6500) );
  NAND U63 ( .A(n6503), .B(n6500), .Z(n4845) );
  XNOR U64 ( .A(n6108), .B(n4845), .Z(out[1000]) );
  XOR U65 ( .A(in[1387]), .B(in[107]), .Z(n4847) );
  XNOR U66 ( .A(in[1067]), .B(in[747]), .Z(n4846) );
  XNOR U67 ( .A(n4847), .B(n4846), .Z(n4848) );
  XOR U68 ( .A(in[427]), .B(n4848), .Z(n5293) );
  XOR U69 ( .A(in[1516]), .B(in[556]), .Z(n4850) );
  XNOR U70 ( .A(in[876]), .B(in[236]), .Z(n4849) );
  XNOR U71 ( .A(n4850), .B(n4849), .Z(n4851) );
  XOR U72 ( .A(in[1196]), .B(n4851), .Z(n6140) );
  XNOR U73 ( .A(n5293), .B(n6140), .Z(n8565) );
  XNOR U74 ( .A(in[172]), .B(n8565), .Z(n6112) );
  XOR U75 ( .A(in[972]), .B(in[12]), .Z(n4853) );
  XNOR U76 ( .A(in[1292]), .B(in[332]), .Z(n4852) );
  XNOR U77 ( .A(n4853), .B(n4852), .Z(n4854) );
  XOR U78 ( .A(in[652]), .B(n4854), .Z(n6030) );
  XOR U79 ( .A(in[141]), .B(in[461]), .Z(n4856) );
  XNOR U80 ( .A(in[1101]), .B(in[1421]), .Z(n4855) );
  XNOR U81 ( .A(n4856), .B(n4855), .Z(n4857) );
  XNOR U82 ( .A(in[781]), .B(n4857), .Z(n5971) );
  XNOR U83 ( .A(n6030), .B(n5971), .Z(n8905) );
  XNOR U84 ( .A(in[1357]), .B(n8905), .Z(n6507) );
  XOR U85 ( .A(in[1365]), .B(in[725]), .Z(n4859) );
  XNOR U86 ( .A(in[85]), .B(in[405]), .Z(n4858) );
  XNOR U87 ( .A(n4859), .B(n4858), .Z(n4860) );
  XOR U88 ( .A(in[1045]), .B(n4860), .Z(n5597) );
  XOR U89 ( .A(in[1556]), .B(in[596]), .Z(n4862) );
  XNOR U90 ( .A(in[916]), .B(in[276]), .Z(n4861) );
  XNOR U91 ( .A(n4862), .B(n4861), .Z(n4863) );
  XOR U92 ( .A(in[1236]), .B(n4863), .Z(n5311) );
  XNOR U93 ( .A(n5597), .B(n5311), .Z(n8691) );
  XNOR U94 ( .A(in[981]), .B(n8691), .Z(n6504) );
  NAND U95 ( .A(n6507), .B(n6504), .Z(n4864) );
  XNOR U96 ( .A(n6112), .B(n4864), .Z(out[1001]) );
  XOR U97 ( .A(in[1388]), .B(in[108]), .Z(n4866) );
  XNOR U98 ( .A(in[1068]), .B(in[748]), .Z(n4865) );
  XNOR U99 ( .A(n4866), .B(n4865), .Z(n4867) );
  XOR U100 ( .A(in[428]), .B(n4867), .Z(n6202) );
  XOR U101 ( .A(in[1517]), .B(in[557]), .Z(n4869) );
  XNOR U102 ( .A(in[877]), .B(in[237]), .Z(n4868) );
  XNOR U103 ( .A(n4869), .B(n4868), .Z(n4870) );
  XOR U104 ( .A(in[1197]), .B(n4870), .Z(n6144) );
  XNOR U105 ( .A(n6202), .B(n6144), .Z(n8569) );
  XNOR U106 ( .A(in[173]), .B(n8569), .Z(n6117) );
  XOR U107 ( .A(in[973]), .B(in[13]), .Z(n4872) );
  XNOR U108 ( .A(in[1293]), .B(in[333]), .Z(n4871) );
  XNOR U109 ( .A(n4872), .B(n4871), .Z(n4873) );
  XOR U110 ( .A(in[653]), .B(n4873), .Z(n6033) );
  XOR U111 ( .A(in[142]), .B(in[1422]), .Z(n4875) );
  XNOR U112 ( .A(in[1102]), .B(in[782]), .Z(n4874) );
  XNOR U113 ( .A(n4875), .B(n4874), .Z(n4876) );
  XNOR U114 ( .A(in[462]), .B(n4876), .Z(n5976) );
  XNOR U115 ( .A(n6033), .B(n5976), .Z(n8908) );
  XNOR U116 ( .A(in[1358]), .B(n8908), .Z(n6511) );
  XOR U117 ( .A(in[1366]), .B(in[726]), .Z(n4878) );
  XNOR U118 ( .A(in[86]), .B(in[406]), .Z(n4877) );
  XNOR U119 ( .A(n4878), .B(n4877), .Z(n4879) );
  XOR U120 ( .A(in[1046]), .B(n4879), .Z(n5610) );
  XOR U121 ( .A(in[1557]), .B(in[597]), .Z(n4881) );
  XNOR U122 ( .A(in[917]), .B(in[277]), .Z(n4880) );
  XNOR U123 ( .A(n4881), .B(n4880), .Z(n4882) );
  XOR U124 ( .A(in[1237]), .B(n4882), .Z(n5326) );
  XNOR U125 ( .A(n5610), .B(n5326), .Z(n8693) );
  XNOR U126 ( .A(in[982]), .B(n8693), .Z(n6508) );
  NAND U127 ( .A(n6511), .B(n6508), .Z(n4883) );
  XNOR U128 ( .A(n6117), .B(n4883), .Z(out[1002]) );
  XOR U129 ( .A(in[1389]), .B(in[109]), .Z(n4885) );
  XNOR U130 ( .A(in[1069]), .B(in[749]), .Z(n4884) );
  XNOR U131 ( .A(n4885), .B(n4884), .Z(n4886) );
  XOR U132 ( .A(in[429]), .B(n4886), .Z(n6206) );
  XOR U133 ( .A(in[1518]), .B(in[558]), .Z(n4888) );
  XNOR U134 ( .A(in[878]), .B(in[238]), .Z(n4887) );
  XNOR U135 ( .A(n4888), .B(n4887), .Z(n4889) );
  XOR U136 ( .A(in[1198]), .B(n4889), .Z(n6148) );
  XNOR U137 ( .A(n6206), .B(n6148), .Z(n8573) );
  XNOR U138 ( .A(in[174]), .B(n8573), .Z(n6121) );
  XOR U139 ( .A(in[143]), .B(in[1423]), .Z(n4891) );
  XNOR U140 ( .A(in[1103]), .B(in[783]), .Z(n4890) );
  XNOR U141 ( .A(n4891), .B(n4890), .Z(n4892) );
  XOR U142 ( .A(in[463]), .B(n4892), .Z(n5981) );
  XOR U143 ( .A(in[974]), .B(in[14]), .Z(n4894) );
  XNOR U144 ( .A(in[1294]), .B(in[334]), .Z(n4893) );
  XNOR U145 ( .A(n4894), .B(n4893), .Z(n4895) );
  XNOR U146 ( .A(in[654]), .B(n4895), .Z(n6036) );
  XNOR U147 ( .A(n5981), .B(n6036), .Z(n8911) );
  XNOR U148 ( .A(in[1359]), .B(n8911), .Z(n6515) );
  XOR U149 ( .A(in[1367]), .B(in[727]), .Z(n4897) );
  XNOR U150 ( .A(in[87]), .B(in[407]), .Z(n4896) );
  XNOR U151 ( .A(n4897), .B(n4896), .Z(n4898) );
  XOR U152 ( .A(in[1047]), .B(n4898), .Z(n5623) );
  XOR U153 ( .A(in[1558]), .B(in[598]), .Z(n4900) );
  XNOR U154 ( .A(in[918]), .B(in[278]), .Z(n4899) );
  XNOR U155 ( .A(n4900), .B(n4899), .Z(n4901) );
  XOR U156 ( .A(in[1238]), .B(n4901), .Z(n5341) );
  XNOR U157 ( .A(n5623), .B(n5341), .Z(n8695) );
  XNOR U158 ( .A(in[983]), .B(n8695), .Z(n6512) );
  NAND U159 ( .A(n6515), .B(n6512), .Z(n4902) );
  XNOR U160 ( .A(n6121), .B(n4902), .Z(out[1003]) );
  XOR U161 ( .A(in[1390]), .B(in[110]), .Z(n4904) );
  XNOR U162 ( .A(in[1070]), .B(in[750]), .Z(n4903) );
  XNOR U163 ( .A(n4904), .B(n4903), .Z(n4905) );
  XOR U164 ( .A(in[430]), .B(n4905), .Z(n6210) );
  XOR U165 ( .A(in[1519]), .B(in[559]), .Z(n4907) );
  XNOR U166 ( .A(in[879]), .B(in[239]), .Z(n4906) );
  XNOR U167 ( .A(n4907), .B(n4906), .Z(n4908) );
  XOR U168 ( .A(in[1199]), .B(n4908), .Z(n6152) );
  XNOR U169 ( .A(n6210), .B(n6152), .Z(n8577) );
  XNOR U170 ( .A(in[175]), .B(n8577), .Z(n6125) );
  XOR U171 ( .A(in[144]), .B(in[1424]), .Z(n4910) );
  XNOR U172 ( .A(in[1104]), .B(in[784]), .Z(n4909) );
  XNOR U173 ( .A(n4910), .B(n4909), .Z(n4911) );
  XOR U174 ( .A(in[464]), .B(n4911), .Z(n5986) );
  XOR U175 ( .A(in[975]), .B(in[15]), .Z(n4913) );
  XNOR U176 ( .A(in[1295]), .B(in[335]), .Z(n4912) );
  XNOR U177 ( .A(n4913), .B(n4912), .Z(n4914) );
  XNOR U178 ( .A(in[655]), .B(n4914), .Z(n6039) );
  XNOR U179 ( .A(n5986), .B(n6039), .Z(n8914) );
  XNOR U180 ( .A(in[1360]), .B(n8914), .Z(n6520) );
  XOR U181 ( .A(in[1368]), .B(in[728]), .Z(n4916) );
  XNOR U182 ( .A(in[88]), .B(in[408]), .Z(n4915) );
  XNOR U183 ( .A(n4916), .B(n4915), .Z(n4917) );
  XOR U184 ( .A(in[1048]), .B(n4917), .Z(n5636) );
  XOR U185 ( .A(in[1559]), .B(in[599]), .Z(n4919) );
  XNOR U186 ( .A(in[919]), .B(in[279]), .Z(n4918) );
  XNOR U187 ( .A(n4919), .B(n4918), .Z(n4920) );
  XOR U188 ( .A(in[1239]), .B(n4920), .Z(n5356) );
  XNOR U189 ( .A(n5636), .B(n5356), .Z(n8697) );
  XNOR U190 ( .A(in[984]), .B(n8697), .Z(n6517) );
  NAND U191 ( .A(n6520), .B(n6517), .Z(n4921) );
  XNOR U192 ( .A(n6125), .B(n4921), .Z(out[1004]) );
  XOR U193 ( .A(in[1391]), .B(in[111]), .Z(n4923) );
  XNOR U194 ( .A(in[1071]), .B(in[751]), .Z(n4922) );
  XNOR U195 ( .A(n4923), .B(n4922), .Z(n4924) );
  XOR U196 ( .A(in[431]), .B(n4924), .Z(n6214) );
  XOR U197 ( .A(in[1520]), .B(in[560]), .Z(n4926) );
  XNOR U198 ( .A(in[880]), .B(in[240]), .Z(n4925) );
  XNOR U199 ( .A(n4926), .B(n4925), .Z(n4927) );
  XOR U200 ( .A(in[1200]), .B(n4927), .Z(n6157) );
  XNOR U201 ( .A(n6214), .B(n6157), .Z(n8581) );
  XNOR U202 ( .A(in[176]), .B(n8581), .Z(n6129) );
  XOR U203 ( .A(in[145]), .B(in[1425]), .Z(n4929) );
  XNOR U204 ( .A(in[1105]), .B(in[785]), .Z(n4928) );
  XNOR U205 ( .A(n4929), .B(n4928), .Z(n4930) );
  XOR U206 ( .A(in[465]), .B(n4930), .Z(n5991) );
  XOR U207 ( .A(in[976]), .B(in[16]), .Z(n4932) );
  XNOR U208 ( .A(in[1296]), .B(in[336]), .Z(n4931) );
  XNOR U209 ( .A(n4932), .B(n4931), .Z(n4933) );
  XNOR U210 ( .A(in[656]), .B(n4933), .Z(n6042) );
  XNOR U211 ( .A(n5991), .B(n6042), .Z(n8921) );
  XNOR U212 ( .A(in[1361]), .B(n8921), .Z(n6524) );
  XOR U213 ( .A(in[1369]), .B(in[729]), .Z(n4935) );
  XNOR U214 ( .A(in[89]), .B(in[409]), .Z(n4934) );
  XNOR U215 ( .A(n4935), .B(n4934), .Z(n4936) );
  XOR U216 ( .A(in[1049]), .B(n4936), .Z(n5649) );
  XOR U217 ( .A(in[1560]), .B(in[600]), .Z(n4938) );
  XNOR U218 ( .A(in[920]), .B(in[280]), .Z(n4937) );
  XNOR U219 ( .A(n4938), .B(n4937), .Z(n4939) );
  XOR U220 ( .A(in[1240]), .B(n4939), .Z(n5371) );
  XNOR U221 ( .A(n5649), .B(n5371), .Z(n8699) );
  XNOR U222 ( .A(in[985]), .B(n8699), .Z(n6521) );
  NAND U223 ( .A(n6524), .B(n6521), .Z(n4940) );
  XNOR U224 ( .A(n6129), .B(n4940), .Z(out[1005]) );
  XOR U225 ( .A(in[1392]), .B(in[112]), .Z(n4942) );
  XNOR U226 ( .A(in[1072]), .B(in[752]), .Z(n4941) );
  XNOR U227 ( .A(n4942), .B(n4941), .Z(n4943) );
  XOR U228 ( .A(in[432]), .B(n4943), .Z(n6218) );
  XOR U229 ( .A(in[1521]), .B(in[561]), .Z(n4945) );
  XNOR U230 ( .A(in[881]), .B(in[241]), .Z(n4944) );
  XNOR U231 ( .A(n4945), .B(n4944), .Z(n4946) );
  XOR U232 ( .A(in[1201]), .B(n4946), .Z(n6161) );
  XNOR U233 ( .A(n6218), .B(n6161), .Z(n8585) );
  XNOR U234 ( .A(in[177]), .B(n8585), .Z(n6133) );
  XOR U235 ( .A(in[17]), .B(in[657]), .Z(n4948) );
  XNOR U236 ( .A(in[977]), .B(in[337]), .Z(n4947) );
  XNOR U237 ( .A(n4948), .B(n4947), .Z(n4949) );
  XOR U238 ( .A(in[1297]), .B(n4949), .Z(n6045) );
  XOR U239 ( .A(in[1426]), .B(in[466]), .Z(n4951) );
  XNOR U240 ( .A(in[786]), .B(in[146]), .Z(n4950) );
  XNOR U241 ( .A(n4951), .B(n4950), .Z(n4952) );
  XNOR U242 ( .A(in[1106]), .B(n4952), .Z(n5295) );
  XNOR U243 ( .A(n6045), .B(n5295), .Z(n8924) );
  XNOR U244 ( .A(n8924), .B(in[1362]), .Z(n6528) );
  XOR U245 ( .A(in[1370]), .B(in[730]), .Z(n4954) );
  XNOR U246 ( .A(in[90]), .B(in[410]), .Z(n4953) );
  XNOR U247 ( .A(n4954), .B(n4953), .Z(n4955) );
  XOR U248 ( .A(in[1050]), .B(n4955), .Z(n5664) );
  XOR U249 ( .A(in[1561]), .B(in[601]), .Z(n4957) );
  XNOR U250 ( .A(in[921]), .B(in[281]), .Z(n4956) );
  XNOR U251 ( .A(n4957), .B(n4956), .Z(n4958) );
  XOR U252 ( .A(in[1241]), .B(n4958), .Z(n5397) );
  XNOR U253 ( .A(n5664), .B(n5397), .Z(n8701) );
  XNOR U254 ( .A(in[986]), .B(n8701), .Z(n6525) );
  NAND U255 ( .A(n6528), .B(n6525), .Z(n4959) );
  XNOR U256 ( .A(n6133), .B(n4959), .Z(out[1006]) );
  XOR U257 ( .A(in[1393]), .B(in[113]), .Z(n4961) );
  XNOR U258 ( .A(in[1073]), .B(in[753]), .Z(n4960) );
  XNOR U259 ( .A(n4961), .B(n4960), .Z(n4962) );
  XOR U260 ( .A(in[433]), .B(n4962), .Z(n6222) );
  XOR U261 ( .A(in[1522]), .B(in[562]), .Z(n4964) );
  XNOR U262 ( .A(in[882]), .B(in[242]), .Z(n4963) );
  XNOR U263 ( .A(n4964), .B(n4963), .Z(n4965) );
  XOR U264 ( .A(in[1202]), .B(n4965), .Z(n6165) );
  XNOR U265 ( .A(n6222), .B(n6165), .Z(n8589) );
  XNOR U266 ( .A(in[178]), .B(n8589), .Z(n6137) );
  XOR U267 ( .A(in[147]), .B(in[1427]), .Z(n4967) );
  XNOR U268 ( .A(in[1107]), .B(in[787]), .Z(n4966) );
  XNOR U269 ( .A(n4967), .B(n4966), .Z(n4968) );
  XOR U270 ( .A(in[467]), .B(n4968), .Z(n5310) );
  XOR U271 ( .A(in[978]), .B(in[18]), .Z(n4970) );
  XNOR U272 ( .A(in[1298]), .B(in[338]), .Z(n4969) );
  XNOR U273 ( .A(n4970), .B(n4969), .Z(n4971) );
  XNOR U274 ( .A(in[658]), .B(n4971), .Z(n6048) );
  XNOR U275 ( .A(n5310), .B(n6048), .Z(n8927) );
  XNOR U276 ( .A(in[1363]), .B(n8927), .Z(n6532) );
  XOR U277 ( .A(in[1371]), .B(in[731]), .Z(n4973) );
  XNOR U278 ( .A(in[91]), .B(in[411]), .Z(n4972) );
  XNOR U279 ( .A(n4973), .B(n4972), .Z(n4974) );
  XOR U280 ( .A(in[1051]), .B(n4974), .Z(n5677) );
  XOR U281 ( .A(in[1562]), .B(in[602]), .Z(n4976) );
  XNOR U282 ( .A(in[922]), .B(in[282]), .Z(n4975) );
  XNOR U283 ( .A(n4976), .B(n4975), .Z(n4977) );
  XOR U284 ( .A(in[1242]), .B(n4977), .Z(n5412) );
  XNOR U285 ( .A(n5677), .B(n5412), .Z(n8703) );
  XNOR U286 ( .A(in[987]), .B(n8703), .Z(n6529) );
  NAND U287 ( .A(n6532), .B(n6529), .Z(n4978) );
  XNOR U288 ( .A(n6137), .B(n4978), .Z(out[1007]) );
  XOR U289 ( .A(in[1394]), .B(in[114]), .Z(n4980) );
  XNOR U290 ( .A(in[1074]), .B(in[754]), .Z(n4979) );
  XNOR U291 ( .A(n4980), .B(n4979), .Z(n4981) );
  XOR U292 ( .A(in[434]), .B(n4981), .Z(n6226) );
  XOR U293 ( .A(in[1523]), .B(in[563]), .Z(n4983) );
  XNOR U294 ( .A(in[883]), .B(in[243]), .Z(n4982) );
  XNOR U295 ( .A(n4983), .B(n4982), .Z(n4984) );
  XOR U296 ( .A(in[1203]), .B(n4984), .Z(n6169) );
  XNOR U297 ( .A(n6226), .B(n6169), .Z(n8593) );
  XNOR U298 ( .A(in[179]), .B(n8593), .Z(n6141) );
  XOR U299 ( .A(in[148]), .B(in[1428]), .Z(n4986) );
  XNOR U300 ( .A(in[1108]), .B(in[788]), .Z(n4985) );
  XNOR U301 ( .A(n4986), .B(n4985), .Z(n4987) );
  XOR U302 ( .A(in[468]), .B(n4987), .Z(n5325) );
  XOR U303 ( .A(in[979]), .B(in[19]), .Z(n4989) );
  XNOR U304 ( .A(in[1299]), .B(in[339]), .Z(n4988) );
  XNOR U305 ( .A(n4989), .B(n4988), .Z(n4990) );
  XNOR U306 ( .A(in[659]), .B(n4990), .Z(n6052) );
  XNOR U307 ( .A(n5325), .B(n6052), .Z(n8930) );
  XNOR U308 ( .A(in[1364]), .B(n8930), .Z(n6536) );
  XOR U309 ( .A(in[1372]), .B(in[732]), .Z(n4992) );
  XNOR U310 ( .A(in[92]), .B(in[412]), .Z(n4991) );
  XNOR U311 ( .A(n4992), .B(n4991), .Z(n4993) );
  XOR U312 ( .A(in[1052]), .B(n4993), .Z(n5697) );
  XOR U313 ( .A(in[1563]), .B(in[603]), .Z(n4995) );
  XNOR U314 ( .A(in[923]), .B(in[283]), .Z(n4994) );
  XNOR U315 ( .A(n4995), .B(n4994), .Z(n4996) );
  XOR U316 ( .A(in[1243]), .B(n4996), .Z(n5427) );
  XNOR U317 ( .A(n5697), .B(n5427), .Z(n8707) );
  XNOR U318 ( .A(in[988]), .B(n8707), .Z(n6533) );
  NAND U319 ( .A(n6536), .B(n6533), .Z(n4997) );
  XNOR U320 ( .A(n6141), .B(n4997), .Z(out[1008]) );
  XOR U321 ( .A(in[1395]), .B(in[115]), .Z(n4999) );
  XNOR U322 ( .A(in[1075]), .B(in[755]), .Z(n4998) );
  XNOR U323 ( .A(n4999), .B(n4998), .Z(n5000) );
  XOR U324 ( .A(in[435]), .B(n5000), .Z(n6230) );
  XOR U325 ( .A(in[1524]), .B(in[564]), .Z(n5002) );
  XNOR U326 ( .A(in[884]), .B(in[244]), .Z(n5001) );
  XNOR U327 ( .A(n5002), .B(n5001), .Z(n5003) );
  XOR U328 ( .A(in[1204]), .B(n5003), .Z(n6173) );
  XNOR U329 ( .A(n6230), .B(n6173), .Z(n8597) );
  XNOR U330 ( .A(in[180]), .B(n8597), .Z(n6145) );
  XOR U331 ( .A(in[340]), .B(in[660]), .Z(n5005) );
  XNOR U332 ( .A(in[20]), .B(in[1300]), .Z(n5004) );
  XNOR U333 ( .A(n5005), .B(n5004), .Z(n5006) );
  XOR U334 ( .A(in[980]), .B(n5006), .Z(n6055) );
  XOR U335 ( .A(in[149]), .B(in[1429]), .Z(n5008) );
  XNOR U336 ( .A(in[1109]), .B(in[789]), .Z(n5007) );
  XNOR U337 ( .A(n5008), .B(n5007), .Z(n5009) );
  XNOR U338 ( .A(in[469]), .B(n5009), .Z(n5340) );
  XNOR U339 ( .A(n6055), .B(n5340), .Z(n8933) );
  XNOR U340 ( .A(in[1365]), .B(n8933), .Z(n6540) );
  XOR U341 ( .A(in[1373]), .B(in[733]), .Z(n5011) );
  XNOR U342 ( .A(in[93]), .B(in[413]), .Z(n5010) );
  XNOR U343 ( .A(n5011), .B(n5010), .Z(n5012) );
  XOR U344 ( .A(in[1053]), .B(n5012), .Z(n5710) );
  XOR U345 ( .A(in[1564]), .B(in[604]), .Z(n5014) );
  XNOR U346 ( .A(in[924]), .B(in[284]), .Z(n5013) );
  XNOR U347 ( .A(n5014), .B(n5013), .Z(n5015) );
  XOR U348 ( .A(in[1244]), .B(n5015), .Z(n5442) );
  XNOR U349 ( .A(n5710), .B(n5442), .Z(n8709) );
  XNOR U350 ( .A(in[989]), .B(n8709), .Z(n6537) );
  NAND U351 ( .A(n6540), .B(n6537), .Z(n5016) );
  XNOR U352 ( .A(n6145), .B(n5016), .Z(out[1009]) );
  XOR U353 ( .A(in[1339]), .B(in[59]), .Z(n5018) );
  XNOR U354 ( .A(in[699]), .B(in[379]), .Z(n5017) );
  XNOR U355 ( .A(n5018), .B(n5017), .Z(n5019) );
  XOR U356 ( .A(in[1019]), .B(n5019), .Z(n5668) );
  XOR U357 ( .A(in[1530]), .B(in[570]), .Z(n5021) );
  XNOR U358 ( .A(in[1210]), .B(in[250]), .Z(n5020) );
  XNOR U359 ( .A(n5021), .B(n5020), .Z(n5022) );
  XOR U360 ( .A(in[890]), .B(n5022), .Z(n5134) );
  XNOR U361 ( .A(n5668), .B(n5134), .Z(n8399) );
  XNOR U362 ( .A(in[635]), .B(n8399), .Z(n7357) );
  XOR U363 ( .A(in[161]), .B(in[1441]), .Z(n5024) );
  XNOR U364 ( .A(in[801]), .B(in[1121]), .Z(n5023) );
  XNOR U365 ( .A(n5024), .B(n5023), .Z(n5025) );
  XOR U366 ( .A(in[481]), .B(n5025), .Z(n5261) );
  XOR U367 ( .A(in[1570]), .B(in[610]), .Z(n5027) );
  XNOR U368 ( .A(in[930]), .B(in[290]), .Z(n5026) );
  XNOR U369 ( .A(n5027), .B(n5026), .Z(n5028) );
  XNOR U370 ( .A(in[1250]), .B(n5028), .Z(n5144) );
  XNOR U371 ( .A(n5261), .B(n5144), .Z(n8496) );
  XNOR U372 ( .A(in[226]), .B(n8496), .Z(n7638) );
  XOR U373 ( .A(in[1510]), .B(in[550]), .Z(n5030) );
  XNOR U374 ( .A(in[870]), .B(in[230]), .Z(n5029) );
  XNOR U375 ( .A(n5030), .B(n5029), .Z(n5031) );
  XOR U376 ( .A(in[1190]), .B(n5031), .Z(n6116) );
  XOR U377 ( .A(in[1061]), .B(in[421]), .Z(n5033) );
  XNOR U378 ( .A(in[741]), .B(in[1381]), .Z(n5032) );
  XNOR U379 ( .A(n5033), .B(n5032), .Z(n5034) );
  XOR U380 ( .A(in[101]), .B(n5034), .Z(n5180) );
  XNOR U381 ( .A(n6116), .B(n5180), .Z(n8537) );
  XNOR U382 ( .A(in[1446]), .B(n8537), .Z(n7635) );
  NAND U383 ( .A(n7638), .B(n7635), .Z(n5035) );
  XNOR U384 ( .A(n7357), .B(n5035), .Z(out[100]) );
  XOR U385 ( .A(in[1396]), .B(in[116]), .Z(n5037) );
  XNOR U386 ( .A(in[1076]), .B(in[756]), .Z(n5036) );
  XNOR U387 ( .A(n5037), .B(n5036), .Z(n5038) );
  XOR U388 ( .A(in[436]), .B(n5038), .Z(n6235) );
  XOR U389 ( .A(in[1525]), .B(in[565]), .Z(n5040) );
  XNOR U390 ( .A(in[885]), .B(in[245]), .Z(n5039) );
  XNOR U391 ( .A(n5040), .B(n5039), .Z(n5041) );
  XOR U392 ( .A(in[1205]), .B(n5041), .Z(n6177) );
  XNOR U393 ( .A(n6235), .B(n6177), .Z(n8601) );
  XNOR U394 ( .A(in[181]), .B(n8601), .Z(n6149) );
  XOR U395 ( .A(in[341]), .B(in[661]), .Z(n5043) );
  XNOR U396 ( .A(in[21]), .B(in[1301]), .Z(n5042) );
  XNOR U397 ( .A(n5043), .B(n5042), .Z(n5044) );
  XOR U398 ( .A(in[981]), .B(n5044), .Z(n6058) );
  XOR U399 ( .A(in[150]), .B(in[1430]), .Z(n5046) );
  XNOR U400 ( .A(in[1110]), .B(in[790]), .Z(n5045) );
  XNOR U401 ( .A(n5046), .B(n5045), .Z(n5047) );
  XNOR U402 ( .A(in[470]), .B(n5047), .Z(n5355) );
  XNOR U403 ( .A(n6058), .B(n5355), .Z(n8936) );
  XNOR U404 ( .A(in[1366]), .B(n8936), .Z(n6544) );
  XOR U405 ( .A(in[1374]), .B(in[734]), .Z(n5049) );
  XNOR U406 ( .A(in[94]), .B(in[414]), .Z(n5048) );
  XNOR U407 ( .A(n5049), .B(n5048), .Z(n5050) );
  XOR U408 ( .A(in[1054]), .B(n5050), .Z(n5723) );
  XOR U409 ( .A(in[1565]), .B(in[605]), .Z(n5052) );
  XNOR U410 ( .A(in[925]), .B(in[285]), .Z(n5051) );
  XNOR U411 ( .A(n5052), .B(n5051), .Z(n5053) );
  XOR U412 ( .A(in[1245]), .B(n5053), .Z(n5457) );
  XNOR U413 ( .A(n5723), .B(n5457), .Z(n8711) );
  XNOR U414 ( .A(in[990]), .B(n8711), .Z(n6541) );
  NAND U415 ( .A(n6544), .B(n6541), .Z(n5054) );
  XNOR U416 ( .A(n6149), .B(n5054), .Z(out[1010]) );
  XOR U417 ( .A(in[1526]), .B(in[566]), .Z(n5056) );
  XNOR U418 ( .A(in[886]), .B(in[246]), .Z(n5055) );
  XNOR U419 ( .A(n5056), .B(n5055), .Z(n5057) );
  XOR U420 ( .A(in[1206]), .B(n5057), .Z(n6181) );
  XOR U421 ( .A(in[1397]), .B(in[117]), .Z(n5059) );
  XNOR U422 ( .A(in[1077]), .B(in[757]), .Z(n5058) );
  XNOR U423 ( .A(n5059), .B(n5058), .Z(n5060) );
  XOR U424 ( .A(in[437]), .B(n5060), .Z(n6239) );
  XNOR U425 ( .A(n6181), .B(n6239), .Z(n8611) );
  XNOR U426 ( .A(in[182]), .B(n8611), .Z(n6153) );
  XOR U427 ( .A(in[151]), .B(in[1431]), .Z(n5062) );
  XNOR U428 ( .A(in[1111]), .B(in[791]), .Z(n5061) );
  XNOR U429 ( .A(n5062), .B(n5061), .Z(n5063) );
  XOR U430 ( .A(in[471]), .B(n5063), .Z(n5370) );
  XOR U431 ( .A(in[342]), .B(in[662]), .Z(n5065) );
  XNOR U432 ( .A(in[22]), .B(in[1302]), .Z(n5064) );
  XNOR U433 ( .A(n5065), .B(n5064), .Z(n5066) );
  XNOR U434 ( .A(in[982]), .B(n5066), .Z(n6061) );
  XNOR U435 ( .A(n5370), .B(n6061), .Z(n8939) );
  XNOR U436 ( .A(in[1367]), .B(n8939), .Z(n6548) );
  XOR U437 ( .A(in[1375]), .B(in[735]), .Z(n5068) );
  XNOR U438 ( .A(in[95]), .B(in[415]), .Z(n5067) );
  XNOR U439 ( .A(n5068), .B(n5067), .Z(n5069) );
  XOR U440 ( .A(in[1055]), .B(n5069), .Z(n5736) );
  XOR U441 ( .A(in[1566]), .B(in[606]), .Z(n5071) );
  XNOR U442 ( .A(in[926]), .B(in[286]), .Z(n5070) );
  XNOR U443 ( .A(n5071), .B(n5070), .Z(n5072) );
  XOR U444 ( .A(in[1246]), .B(n5072), .Z(n5472) );
  XNOR U445 ( .A(n5736), .B(n5472), .Z(n8713) );
  XNOR U446 ( .A(in[991]), .B(n8713), .Z(n6545) );
  NAND U447 ( .A(n6548), .B(n6545), .Z(n5073) );
  XNOR U448 ( .A(n6153), .B(n5073), .Z(out[1011]) );
  XOR U449 ( .A(in[1527]), .B(in[567]), .Z(n5075) );
  XNOR U450 ( .A(in[887]), .B(in[247]), .Z(n5074) );
  XNOR U451 ( .A(n5075), .B(n5074), .Z(n5076) );
  XOR U452 ( .A(in[1207]), .B(n5076), .Z(n6185) );
  XOR U453 ( .A(in[1398]), .B(in[118]), .Z(n5078) );
  XNOR U454 ( .A(in[1078]), .B(in[758]), .Z(n5077) );
  XNOR U455 ( .A(n5078), .B(n5077), .Z(n5079) );
  XOR U456 ( .A(in[438]), .B(n5079), .Z(n6243) );
  XNOR U457 ( .A(n6185), .B(n6243), .Z(n8615) );
  XNOR U458 ( .A(in[183]), .B(n8615), .Z(n6158) );
  XOR U459 ( .A(in[343]), .B(in[663]), .Z(n5081) );
  XNOR U460 ( .A(in[23]), .B(in[1303]), .Z(n5080) );
  XNOR U461 ( .A(n5081), .B(n5080), .Z(n5082) );
  XOR U462 ( .A(in[983]), .B(n5082), .Z(n6064) );
  XOR U463 ( .A(in[152]), .B(in[1432]), .Z(n5084) );
  XNOR U464 ( .A(in[1112]), .B(in[792]), .Z(n5083) );
  XNOR U465 ( .A(n5084), .B(n5083), .Z(n5085) );
  XNOR U466 ( .A(in[472]), .B(n5085), .Z(n5396) );
  XNOR U467 ( .A(n6064), .B(n5396), .Z(n8942) );
  XNOR U468 ( .A(in[1368]), .B(n8942), .Z(n6552) );
  XOR U469 ( .A(in[1376]), .B(in[736]), .Z(n5087) );
  XNOR U470 ( .A(in[96]), .B(in[416]), .Z(n5086) );
  XNOR U471 ( .A(n5087), .B(n5086), .Z(n5088) );
  XOR U472 ( .A(in[1056]), .B(n5088), .Z(n5751) );
  XOR U473 ( .A(in[1567]), .B(in[607]), .Z(n5090) );
  XNOR U474 ( .A(in[927]), .B(in[287]), .Z(n5089) );
  XNOR U475 ( .A(n5090), .B(n5089), .Z(n5091) );
  XOR U476 ( .A(in[1247]), .B(n5091), .Z(n5487) );
  XNOR U477 ( .A(n5751), .B(n5487), .Z(n8715) );
  XNOR U478 ( .A(in[992]), .B(n8715), .Z(n6549) );
  NAND U479 ( .A(n6552), .B(n6549), .Z(n5092) );
  XNOR U480 ( .A(n6158), .B(n5092), .Z(out[1012]) );
  XOR U481 ( .A(in[1528]), .B(in[568]), .Z(n5094) );
  XNOR U482 ( .A(in[888]), .B(in[248]), .Z(n5093) );
  XNOR U483 ( .A(n5094), .B(n5093), .Z(n5095) );
  XOR U484 ( .A(in[1208]), .B(n5095), .Z(n6189) );
  XOR U485 ( .A(in[1399]), .B(in[119]), .Z(n5097) );
  XNOR U486 ( .A(in[1079]), .B(in[759]), .Z(n5096) );
  XNOR U487 ( .A(n5097), .B(n5096), .Z(n5098) );
  XOR U488 ( .A(in[439]), .B(n5098), .Z(n6247) );
  XNOR U489 ( .A(n6189), .B(n6247), .Z(n8619) );
  XNOR U490 ( .A(in[184]), .B(n8619), .Z(n6162) );
  XOR U491 ( .A(in[344]), .B(in[664]), .Z(n5100) );
  XNOR U492 ( .A(in[24]), .B(in[1304]), .Z(n5099) );
  XNOR U493 ( .A(n5100), .B(n5099), .Z(n5101) );
  XOR U494 ( .A(in[984]), .B(n5101), .Z(n6067) );
  XOR U495 ( .A(in[153]), .B(in[1433]), .Z(n5103) );
  XNOR U496 ( .A(in[1113]), .B(in[793]), .Z(n5102) );
  XNOR U497 ( .A(n5103), .B(n5102), .Z(n5104) );
  XNOR U498 ( .A(in[473]), .B(n5104), .Z(n5411) );
  XNOR U499 ( .A(n6067), .B(n5411), .Z(n8945) );
  XNOR U500 ( .A(in[1369]), .B(n8945), .Z(n6556) );
  XOR U501 ( .A(in[1377]), .B(in[737]), .Z(n5106) );
  XNOR U502 ( .A(in[97]), .B(in[417]), .Z(n5105) );
  XNOR U503 ( .A(n5106), .B(n5105), .Z(n5107) );
  XOR U504 ( .A(in[1057]), .B(n5107), .Z(n5766) );
  XOR U505 ( .A(in[1568]), .B(in[608]), .Z(n5109) );
  XNOR U506 ( .A(in[928]), .B(in[288]), .Z(n5108) );
  XNOR U507 ( .A(n5109), .B(n5108), .Z(n5110) );
  XOR U508 ( .A(in[1248]), .B(n5110), .Z(n5502) );
  XNOR U509 ( .A(n5766), .B(n5502), .Z(n8717) );
  XNOR U510 ( .A(in[993]), .B(n8717), .Z(n6553) );
  NAND U511 ( .A(n6556), .B(n6553), .Z(n5111) );
  XNOR U512 ( .A(n6162), .B(n5111), .Z(out[1013]) );
  XOR U513 ( .A(in[1529]), .B(in[569]), .Z(n5113) );
  XNOR U514 ( .A(in[889]), .B(in[249]), .Z(n5112) );
  XNOR U515 ( .A(n5113), .B(n5112), .Z(n5114) );
  XOR U516 ( .A(in[1209]), .B(n5114), .Z(n6193) );
  XOR U517 ( .A(in[1400]), .B(in[120]), .Z(n5116) );
  XNOR U518 ( .A(in[1080]), .B(in[760]), .Z(n5115) );
  XNOR U519 ( .A(n5116), .B(n5115), .Z(n5117) );
  XOR U520 ( .A(in[440]), .B(n5117), .Z(n6251) );
  XNOR U521 ( .A(n6193), .B(n6251), .Z(n8623) );
  XNOR U522 ( .A(in[185]), .B(n8623), .Z(n6166) );
  XOR U523 ( .A(in[345]), .B(in[665]), .Z(n5119) );
  XNOR U524 ( .A(in[25]), .B(in[1305]), .Z(n5118) );
  XNOR U525 ( .A(n5119), .B(n5118), .Z(n5120) );
  XOR U526 ( .A(in[985]), .B(n5120), .Z(n6070) );
  XOR U527 ( .A(in[154]), .B(in[1434]), .Z(n5122) );
  XNOR U528 ( .A(in[1114]), .B(in[794]), .Z(n5121) );
  XNOR U529 ( .A(n5122), .B(n5121), .Z(n5123) );
  XNOR U530 ( .A(in[474]), .B(n5123), .Z(n5426) );
  XNOR U531 ( .A(n6070), .B(n5426), .Z(n8948) );
  XNOR U532 ( .A(in[1370]), .B(n8948), .Z(n6561) );
  XOR U533 ( .A(in[1569]), .B(in[609]), .Z(n5125) );
  XNOR U534 ( .A(in[929]), .B(in[289]), .Z(n5124) );
  XNOR U535 ( .A(n5125), .B(n5124), .Z(n5126) );
  XOR U536 ( .A(in[1249]), .B(n5126), .Z(n5517) );
  XOR U537 ( .A(in[1378]), .B(in[738]), .Z(n5128) );
  XNOR U538 ( .A(in[98]), .B(in[418]), .Z(n5127) );
  XNOR U539 ( .A(n5128), .B(n5127), .Z(n5129) );
  XOR U540 ( .A(in[1058]), .B(n5129), .Z(n5781) );
  XNOR U541 ( .A(n5517), .B(n5781), .Z(n8719) );
  XNOR U542 ( .A(in[994]), .B(n8719), .Z(n6558) );
  NAND U543 ( .A(n6561), .B(n6558), .Z(n5130) );
  XNOR U544 ( .A(n6166), .B(n5130), .Z(out[1014]) );
  XOR U545 ( .A(in[1401]), .B(in[121]), .Z(n5132) );
  XNOR U546 ( .A(in[1081]), .B(in[761]), .Z(n5131) );
  XNOR U547 ( .A(n5132), .B(n5131), .Z(n5133) );
  XOR U548 ( .A(in[441]), .B(n5133), .Z(n6255) );
  XNOR U549 ( .A(n5134), .B(n6255), .Z(n8345) );
  XNOR U550 ( .A(in[186]), .B(n8345), .Z(n6170) );
  XOR U551 ( .A(in[155]), .B(in[1435]), .Z(n5136) );
  XNOR U552 ( .A(in[1115]), .B(in[795]), .Z(n5135) );
  XNOR U553 ( .A(n5136), .B(n5135), .Z(n5137) );
  XOR U554 ( .A(in[475]), .B(n5137), .Z(n5441) );
  XOR U555 ( .A(in[346]), .B(in[666]), .Z(n5139) );
  XNOR U556 ( .A(in[26]), .B(in[1306]), .Z(n5138) );
  XNOR U557 ( .A(n5139), .B(n5138), .Z(n5140) );
  XNOR U558 ( .A(in[986]), .B(n5140), .Z(n6073) );
  XNOR U559 ( .A(n5441), .B(n6073), .Z(n8955) );
  XNOR U560 ( .A(in[1371]), .B(n8955), .Z(n6565) );
  XOR U561 ( .A(in[1379]), .B(in[739]), .Z(n5142) );
  XNOR U562 ( .A(in[99]), .B(in[419]), .Z(n5141) );
  XNOR U563 ( .A(n5142), .B(n5141), .Z(n5143) );
  XNOR U564 ( .A(in[1059]), .B(n5143), .Z(n5796) );
  XNOR U565 ( .A(n5144), .B(n5796), .Z(n8721) );
  XNOR U566 ( .A(in[995]), .B(n8721), .Z(n6562) );
  NAND U567 ( .A(n6565), .B(n6562), .Z(n5145) );
  XNOR U568 ( .A(n6170), .B(n5145), .Z(out[1015]) );
  XOR U569 ( .A(in[1402]), .B(in[122]), .Z(n5147) );
  XNOR U570 ( .A(in[1082]), .B(in[762]), .Z(n5146) );
  XNOR U571 ( .A(n5147), .B(n5146), .Z(n5148) );
  XOR U572 ( .A(in[442]), .B(n5148), .Z(n6259) );
  XOR U573 ( .A(in[1531]), .B(in[571]), .Z(n5150) );
  XNOR U574 ( .A(in[1211]), .B(in[251]), .Z(n5149) );
  XNOR U575 ( .A(n5150), .B(n5149), .Z(n5151) );
  XOR U576 ( .A(in[891]), .B(n5151), .Z(n5223) );
  XNOR U577 ( .A(n6259), .B(n5223), .Z(n8349) );
  XNOR U578 ( .A(in[187]), .B(n8349), .Z(n6174) );
  XOR U579 ( .A(in[156]), .B(in[1436]), .Z(n5153) );
  XNOR U580 ( .A(in[1116]), .B(in[796]), .Z(n5152) );
  XNOR U581 ( .A(n5153), .B(n5152), .Z(n5154) );
  XOR U582 ( .A(in[476]), .B(n5154), .Z(n5456) );
  XOR U583 ( .A(in[347]), .B(in[667]), .Z(n5156) );
  XNOR U584 ( .A(in[27]), .B(in[1307]), .Z(n5155) );
  XNOR U585 ( .A(n5156), .B(n5155), .Z(n5157) );
  XNOR U586 ( .A(in[987]), .B(n5157), .Z(n6076) );
  XNOR U587 ( .A(n5456), .B(n6076), .Z(n8958) );
  XNOR U588 ( .A(in[1372]), .B(n8958), .Z(n6569) );
  XOR U589 ( .A(in[1060]), .B(in[420]), .Z(n5159) );
  XNOR U590 ( .A(in[740]), .B(in[1380]), .Z(n5158) );
  XNOR U591 ( .A(n5159), .B(n5158), .Z(n5160) );
  XOR U592 ( .A(in[100]), .B(n5160), .Z(n5811) );
  XOR U593 ( .A(in[1571]), .B(in[611]), .Z(n5162) );
  XNOR U594 ( .A(in[931]), .B(in[291]), .Z(n5161) );
  XNOR U595 ( .A(n5162), .B(n5161), .Z(n5163) );
  XOR U596 ( .A(in[1251]), .B(n5163), .Z(n5227) );
  XNOR U597 ( .A(n5811), .B(n5227), .Z(n8723) );
  XNOR U598 ( .A(in[996]), .B(n8723), .Z(n6566) );
  NAND U599 ( .A(n6569), .B(n6566), .Z(n5164) );
  XNOR U600 ( .A(n6174), .B(n5164), .Z(out[1016]) );
  XOR U601 ( .A(in[1403]), .B(in[123]), .Z(n5166) );
  XNOR U602 ( .A(in[1083]), .B(in[763]), .Z(n5165) );
  XNOR U603 ( .A(n5166), .B(n5165), .Z(n5167) );
  XOR U604 ( .A(in[443]), .B(n5167), .Z(n6263) );
  XOR U605 ( .A(in[1532]), .B(in[572]), .Z(n5169) );
  XNOR U606 ( .A(in[1212]), .B(in[252]), .Z(n5168) );
  XNOR U607 ( .A(n5169), .B(n5168), .Z(n5170) );
  XOR U608 ( .A(in[892]), .B(n5170), .Z(n5388) );
  XNOR U609 ( .A(n6263), .B(n5388), .Z(n8353) );
  XNOR U610 ( .A(in[188]), .B(n8353), .Z(n6178) );
  XOR U611 ( .A(in[157]), .B(in[1437]), .Z(n5172) );
  XNOR U612 ( .A(in[1117]), .B(in[797]), .Z(n5171) );
  XNOR U613 ( .A(n5172), .B(n5171), .Z(n5173) );
  XOR U614 ( .A(in[477]), .B(n5173), .Z(n5471) );
  XOR U615 ( .A(in[348]), .B(in[668]), .Z(n5175) );
  XNOR U616 ( .A(in[28]), .B(in[1308]), .Z(n5174) );
  XNOR U617 ( .A(n5175), .B(n5174), .Z(n5176) );
  XNOR U618 ( .A(in[988]), .B(n5176), .Z(n6079) );
  XNOR U619 ( .A(n5471), .B(n6079), .Z(n8961) );
  XNOR U620 ( .A(in[1373]), .B(n8961), .Z(n6573) );
  XOR U621 ( .A(in[1572]), .B(in[612]), .Z(n5178) );
  XNOR U622 ( .A(in[932]), .B(in[292]), .Z(n5177) );
  XNOR U623 ( .A(n5178), .B(n5177), .Z(n5179) );
  XOR U624 ( .A(in[1252]), .B(n5179), .Z(n5390) );
  XNOR U625 ( .A(n5180), .B(n5390), .Z(n8725) );
  XNOR U626 ( .A(in[997]), .B(n8725), .Z(n6570) );
  NAND U627 ( .A(n6573), .B(n6570), .Z(n5181) );
  XNOR U628 ( .A(n6178), .B(n5181), .Z(out[1017]) );
  XOR U629 ( .A(in[1404]), .B(in[124]), .Z(n5183) );
  XNOR U630 ( .A(in[1084]), .B(in[764]), .Z(n5182) );
  XNOR U631 ( .A(n5183), .B(n5182), .Z(n5184) );
  XOR U632 ( .A(in[444]), .B(n5184), .Z(n6267) );
  XOR U633 ( .A(in[1533]), .B(in[573]), .Z(n5186) );
  XNOR U634 ( .A(in[1213]), .B(in[253]), .Z(n5185) );
  XNOR U635 ( .A(n5186), .B(n5185), .Z(n5187) );
  XOR U636 ( .A(in[893]), .B(n5187), .Z(n5547) );
  XNOR U637 ( .A(n6267), .B(n5547), .Z(n8357) );
  XNOR U638 ( .A(in[189]), .B(n8357), .Z(n6182) );
  XOR U639 ( .A(in[158]), .B(in[1438]), .Z(n5189) );
  XNOR U640 ( .A(in[1118]), .B(in[798]), .Z(n5188) );
  XNOR U641 ( .A(n5189), .B(n5188), .Z(n5190) );
  XOR U642 ( .A(in[478]), .B(n5190), .Z(n5486) );
  XOR U643 ( .A(in[349]), .B(in[669]), .Z(n5192) );
  XNOR U644 ( .A(in[29]), .B(in[1309]), .Z(n5191) );
  XNOR U645 ( .A(n5192), .B(n5191), .Z(n5193) );
  XNOR U646 ( .A(in[989]), .B(n5193), .Z(n6083) );
  XNOR U647 ( .A(n5486), .B(n6083), .Z(n8964) );
  XNOR U648 ( .A(in[1374]), .B(n8964), .Z(n6577) );
  XOR U649 ( .A(in[1062]), .B(in[422]), .Z(n5195) );
  XNOR U650 ( .A(in[742]), .B(in[1382]), .Z(n5194) );
  XNOR U651 ( .A(n5195), .B(n5194), .Z(n5196) );
  XOR U652 ( .A(in[102]), .B(n5196), .Z(n5231) );
  XOR U653 ( .A(in[1573]), .B(in[613]), .Z(n5198) );
  XNOR U654 ( .A(in[933]), .B(in[293]), .Z(n5197) );
  XNOR U655 ( .A(n5198), .B(n5197), .Z(n5199) );
  XOR U656 ( .A(in[1253]), .B(n5199), .Z(n5549) );
  XNOR U657 ( .A(n5231), .B(n5549), .Z(n8731) );
  XNOR U658 ( .A(in[998]), .B(n8731), .Z(n6574) );
  NAND U659 ( .A(n6577), .B(n6574), .Z(n5200) );
  XNOR U660 ( .A(n6182), .B(n5200), .Z(out[1018]) );
  XOR U661 ( .A(in[1405]), .B(in[125]), .Z(n5202) );
  XNOR U662 ( .A(in[1085]), .B(in[765]), .Z(n5201) );
  XNOR U663 ( .A(n5202), .B(n5201), .Z(n5203) );
  XOR U664 ( .A(in[445]), .B(n5203), .Z(n6271) );
  XOR U665 ( .A(in[1534]), .B(in[894]), .Z(n5205) );
  XNOR U666 ( .A(in[574]), .B(in[1214]), .Z(n5204) );
  XNOR U667 ( .A(n5205), .B(n5204), .Z(n5206) );
  XOR U668 ( .A(in[254]), .B(n5206), .Z(n5684) );
  XNOR U669 ( .A(n6271), .B(n5684), .Z(n8361) );
  XNOR U670 ( .A(in[190]), .B(n8361), .Z(n6186) );
  XOR U671 ( .A(in[1439]), .B(in[479]), .Z(n5208) );
  XNOR U672 ( .A(in[799]), .B(in[159]), .Z(n5207) );
  XNOR U673 ( .A(n5208), .B(n5207), .Z(n5209) );
  XOR U674 ( .A(in[1119]), .B(n5209), .Z(n5501) );
  XOR U675 ( .A(in[350]), .B(in[670]), .Z(n5211) );
  XNOR U676 ( .A(in[30]), .B(in[1310]), .Z(n5210) );
  XNOR U677 ( .A(n5211), .B(n5210), .Z(n5212) );
  XNOR U678 ( .A(in[990]), .B(n5212), .Z(n6086) );
  XNOR U679 ( .A(n5501), .B(n6086), .Z(n8967) );
  XNOR U680 ( .A(in[1375]), .B(n8967), .Z(n6581) );
  XOR U681 ( .A(in[1063]), .B(in[423]), .Z(n5214) );
  XNOR U682 ( .A(in[743]), .B(in[1383]), .Z(n5213) );
  XNOR U683 ( .A(n5214), .B(n5213), .Z(n5215) );
  XOR U684 ( .A(in[103]), .B(n5215), .Z(n5394) );
  XOR U685 ( .A(in[1574]), .B(in[614]), .Z(n5217) );
  XNOR U686 ( .A(in[934]), .B(in[294]), .Z(n5216) );
  XNOR U687 ( .A(n5217), .B(n5216), .Z(n5218) );
  XOR U688 ( .A(in[1254]), .B(n5218), .Z(n5593) );
  XNOR U689 ( .A(n5394), .B(n5593), .Z(n8733) );
  XNOR U690 ( .A(in[999]), .B(n8733), .Z(n6578) );
  NAND U691 ( .A(n6581), .B(n6578), .Z(n5219) );
  XNOR U692 ( .A(n6186), .B(n5219), .Z(out[1019]) );
  XOR U693 ( .A(in[1340]), .B(in[60]), .Z(n5221) );
  XNOR U694 ( .A(in[700]), .B(in[380]), .Z(n5220) );
  XNOR U695 ( .A(n5221), .B(n5220), .Z(n5222) );
  XOR U696 ( .A(in[1020]), .B(n5222), .Z(n5678) );
  XNOR U697 ( .A(n5223), .B(n5678), .Z(n8403) );
  XNOR U698 ( .A(in[636]), .B(n8403), .Z(n7359) );
  XOR U699 ( .A(in[162]), .B(in[1442]), .Z(n5225) );
  XNOR U700 ( .A(in[802]), .B(in[1122]), .Z(n5224) );
  XNOR U701 ( .A(n5225), .B(n5224), .Z(n5226) );
  XNOR U702 ( .A(in[482]), .B(n5226), .Z(n5278) );
  XNOR U703 ( .A(n5227), .B(n5278), .Z(n8500) );
  XNOR U704 ( .A(in[227]), .B(n8500), .Z(n7652) );
  XOR U705 ( .A(in[1511]), .B(in[551]), .Z(n5229) );
  XNOR U706 ( .A(in[871]), .B(in[231]), .Z(n5228) );
  XNOR U707 ( .A(n5229), .B(n5228), .Z(n5230) );
  XOR U708 ( .A(in[1191]), .B(n5230), .Z(n6120) );
  XNOR U709 ( .A(n5231), .B(n6120), .Z(n8541) );
  XNOR U710 ( .A(in[1447]), .B(n8541), .Z(n7649) );
  NAND U711 ( .A(n7652), .B(n7649), .Z(n5232) );
  XNOR U712 ( .A(n7359), .B(n5232), .Z(out[101]) );
  XOR U713 ( .A(in[1406]), .B(in[126]), .Z(n5234) );
  XNOR U714 ( .A(in[1086]), .B(in[766]), .Z(n5233) );
  XNOR U715 ( .A(n5234), .B(n5233), .Z(n5235) );
  XOR U716 ( .A(in[446]), .B(n5235), .Z(n6276) );
  XOR U717 ( .A(in[1535]), .B(in[575]), .Z(n5237) );
  XNOR U718 ( .A(in[895]), .B(in[255]), .Z(n5236) );
  XNOR U719 ( .A(n5237), .B(n5236), .Z(n5238) );
  XOR U720 ( .A(in[1215]), .B(n5238), .Z(n5831) );
  XNOR U721 ( .A(n6276), .B(n5831), .Z(n8365) );
  XNOR U722 ( .A(in[191]), .B(n8365), .Z(n6190) );
  XOR U723 ( .A(in[1440]), .B(in[480]), .Z(n5240) );
  XNOR U724 ( .A(in[800]), .B(in[160]), .Z(n5239) );
  XNOR U725 ( .A(n5240), .B(n5239), .Z(n5241) );
  XOR U726 ( .A(in[1120]), .B(n5241), .Z(n5516) );
  XOR U727 ( .A(in[351]), .B(in[671]), .Z(n5243) );
  XNOR U728 ( .A(in[31]), .B(in[1311]), .Z(n5242) );
  XNOR U729 ( .A(n5243), .B(n5242), .Z(n5244) );
  XNOR U730 ( .A(in[991]), .B(n5244), .Z(n6089) );
  XNOR U731 ( .A(n5516), .B(n6089), .Z(n8970) );
  XNOR U732 ( .A(in[1376]), .B(n8970), .Z(n6585) );
  XOR U733 ( .A(in[1064]), .B(in[424]), .Z(n5246) );
  XNOR U734 ( .A(in[744]), .B(in[1384]), .Z(n5245) );
  XNOR U735 ( .A(n5246), .B(n5245), .Z(n5247) );
  XOR U736 ( .A(in[104]), .B(n5247), .Z(n5553) );
  XOR U737 ( .A(in[1575]), .B(in[615]), .Z(n5249) );
  XNOR U738 ( .A(in[935]), .B(in[295]), .Z(n5248) );
  XNOR U739 ( .A(n5249), .B(n5248), .Z(n5250) );
  XOR U740 ( .A(in[1255]), .B(n5250), .Z(n5606) );
  XNOR U741 ( .A(n5553), .B(n5606), .Z(n8735) );
  XNOR U742 ( .A(in[1000]), .B(n8735), .Z(n6582) );
  NAND U743 ( .A(n6585), .B(n6582), .Z(n5251) );
  XNOR U744 ( .A(n6190), .B(n5251), .Z(out[1020]) );
  XOR U745 ( .A(in[1407]), .B(in[127]), .Z(n5253) );
  XNOR U746 ( .A(in[1087]), .B(in[767]), .Z(n5252) );
  XNOR U747 ( .A(n5253), .B(n5252), .Z(n5254) );
  XOR U748 ( .A(in[447]), .B(n5254), .Z(n6279) );
  XOR U749 ( .A(in[1472]), .B(in[512]), .Z(n5256) );
  XNOR U750 ( .A(in[832]), .B(in[192]), .Z(n5255) );
  XNOR U751 ( .A(n5256), .B(n5255), .Z(n5257) );
  XOR U752 ( .A(in[1152]), .B(n5257), .Z(n5898) );
  XNOR U753 ( .A(n6279), .B(n5898), .Z(n8369) );
  XNOR U754 ( .A(in[128]), .B(n8369), .Z(n6194) );
  XOR U755 ( .A(in[352]), .B(in[672]), .Z(n5259) );
  XNOR U756 ( .A(in[32]), .B(in[1312]), .Z(n5258) );
  XNOR U757 ( .A(n5259), .B(n5258), .Z(n5260) );
  XNOR U758 ( .A(in[992]), .B(n5260), .Z(n6092) );
  XNOR U759 ( .A(n5261), .B(n6092), .Z(n8973) );
  XNOR U760 ( .A(in[1377]), .B(n8973), .Z(n6589) );
  XOR U761 ( .A(in[1065]), .B(in[425]), .Z(n5263) );
  XNOR U762 ( .A(in[745]), .B(in[1385]), .Z(n5262) );
  XNOR U763 ( .A(n5263), .B(n5262), .Z(n5264) );
  XOR U764 ( .A(in[105]), .B(n5264), .Z(n5688) );
  XOR U765 ( .A(in[1576]), .B(in[616]), .Z(n5266) );
  XNOR U766 ( .A(in[936]), .B(in[296]), .Z(n5265) );
  XNOR U767 ( .A(n5266), .B(n5265), .Z(n5267) );
  XOR U768 ( .A(in[1256]), .B(n5267), .Z(n5619) );
  XNOR U769 ( .A(n5688), .B(n5619), .Z(n8737) );
  XNOR U770 ( .A(in[1001]), .B(n8737), .Z(n6586) );
  NAND U771 ( .A(n6589), .B(n6586), .Z(n5268) );
  XNOR U772 ( .A(n6194), .B(n5268), .Z(out[1021]) );
  XOR U773 ( .A(in[1344]), .B(in[64]), .Z(n5270) );
  XNOR U774 ( .A(in[1024]), .B(in[384]), .Z(n5269) );
  XNOR U775 ( .A(n5270), .B(n5269), .Z(n5271) );
  XOR U776 ( .A(in[704]), .B(n5271), .Z(n6284) );
  XOR U777 ( .A(in[1473]), .B(in[513]), .Z(n5273) );
  XNOR U778 ( .A(in[833]), .B(in[193]), .Z(n5272) );
  XNOR U779 ( .A(n5273), .B(n5272), .Z(n5274) );
  XOR U780 ( .A(in[1153]), .B(n5274), .Z(n5951) );
  XNOR U781 ( .A(n6284), .B(n5951), .Z(n8373) );
  XNOR U782 ( .A(in[129]), .B(n8373), .Z(n6197) );
  XOR U783 ( .A(in[353]), .B(in[673]), .Z(n5276) );
  XNOR U784 ( .A(in[33]), .B(in[1313]), .Z(n5275) );
  XNOR U785 ( .A(n5276), .B(n5275), .Z(n5277) );
  XOR U786 ( .A(in[993]), .B(n5277), .Z(n6095) );
  XNOR U787 ( .A(n6095), .B(n5278), .Z(n8976) );
  XNOR U788 ( .A(in[1378]), .B(n8976), .Z(n6593) );
  XOR U789 ( .A(in[1577]), .B(in[617]), .Z(n5280) );
  XNOR U790 ( .A(in[937]), .B(in[297]), .Z(n5279) );
  XNOR U791 ( .A(n5280), .B(n5279), .Z(n5281) );
  XOR U792 ( .A(in[1257]), .B(n5281), .Z(n5632) );
  XNOR U793 ( .A(n5282), .B(n5632), .Z(n8739) );
  XNOR U794 ( .A(in[1002]), .B(n8739), .Z(n6590) );
  NAND U795 ( .A(n6593), .B(n6590), .Z(n5283) );
  XNOR U796 ( .A(n6197), .B(n5283), .Z(out[1022]) );
  XOR U797 ( .A(n8377), .B(in[130]), .Z(n6199) );
  XOR U798 ( .A(in[354]), .B(in[674]), .Z(n5285) );
  XNOR U799 ( .A(in[34]), .B(in[1314]), .Z(n5284) );
  XNOR U800 ( .A(n5285), .B(n5284), .Z(n5286) );
  XOR U801 ( .A(in[994]), .B(n5286), .Z(n6098) );
  XOR U802 ( .A(in[163]), .B(in[1443]), .Z(n5288) );
  XNOR U803 ( .A(in[803]), .B(in[1123]), .Z(n5287) );
  XNOR U804 ( .A(n5288), .B(n5287), .Z(n5289) );
  XNOR U805 ( .A(in[483]), .B(n5289), .Z(n5389) );
  XNOR U806 ( .A(n6098), .B(n5389), .Z(n8979) );
  XNOR U807 ( .A(in[1379]), .B(n8979), .Z(n6597) );
  XOR U808 ( .A(in[1578]), .B(in[618]), .Z(n5291) );
  XNOR U809 ( .A(in[938]), .B(in[298]), .Z(n5290) );
  XNOR U810 ( .A(n5291), .B(n5290), .Z(n5292) );
  XOR U811 ( .A(in[1258]), .B(n5292), .Z(n5645) );
  XNOR U812 ( .A(n5293), .B(n5645), .Z(n8741) );
  XNOR U813 ( .A(in[1003]), .B(n8741), .Z(n6594) );
  NAND U814 ( .A(n6597), .B(n6594), .Z(n5294) );
  XNOR U815 ( .A(n6199), .B(n5294), .Z(out[1023]) );
  XOR U816 ( .A(n5296), .B(n5295), .Z(n8432) );
  XNOR U817 ( .A(in[531]), .B(n8432), .Z(n6203) );
  XOR U818 ( .A(in[1346]), .B(in[66]), .Z(n5298) );
  XNOR U819 ( .A(in[1026]), .B(in[386]), .Z(n5297) );
  XNOR U820 ( .A(n5298), .B(n5297), .Z(n5299) );
  XOR U821 ( .A(in[706]), .B(n5299), .Z(n6292) );
  XOR U822 ( .A(in[1475]), .B(in[515]), .Z(n5301) );
  XNOR U823 ( .A(in[835]), .B(in[195]), .Z(n5300) );
  XNOR U824 ( .A(n5301), .B(n5300), .Z(n5302) );
  XNOR U825 ( .A(in[1155]), .B(n5302), .Z(n6003) );
  XNOR U826 ( .A(n6292), .B(n6003), .Z(n8381) );
  XNOR U827 ( .A(in[131]), .B(n8381), .Z(n9438) );
  XOR U828 ( .A(in[164]), .B(in[1444]), .Z(n5304) );
  XNOR U829 ( .A(in[804]), .B(in[1124]), .Z(n5303) );
  XNOR U830 ( .A(n5304), .B(n5303), .Z(n5305) );
  XOR U831 ( .A(in[484]), .B(n5305), .Z(n5548) );
  XOR U832 ( .A(in[35]), .B(in[675]), .Z(n5307) );
  XNOR U833 ( .A(in[355]), .B(in[1315]), .Z(n5306) );
  XNOR U834 ( .A(n5307), .B(n5306), .Z(n5308) );
  XOR U835 ( .A(in[995]), .B(n5308), .Z(n6101) );
  XNOR U836 ( .A(n5548), .B(n6101), .Z(n8982) );
  XNOR U837 ( .A(in[1380]), .B(n8982), .Z(n9435) );
  NAND U838 ( .A(n9438), .B(n9435), .Z(n5309) );
  XNOR U839 ( .A(n6203), .B(n5309), .Z(out[1024]) );
  XNOR U840 ( .A(n5311), .B(n5310), .Z(n8436) );
  XNOR U841 ( .A(in[532]), .B(n8436), .Z(n6207) );
  XOR U842 ( .A(in[1347]), .B(in[67]), .Z(n5313) );
  XNOR U843 ( .A(in[1027]), .B(in[387]), .Z(n5312) );
  XNOR U844 ( .A(n5313), .B(n5312), .Z(n5314) );
  XOR U845 ( .A(in[707]), .B(n5314), .Z(n6296) );
  XOR U846 ( .A(in[1476]), .B(in[516]), .Z(n5316) );
  XNOR U847 ( .A(in[836]), .B(in[196]), .Z(n5315) );
  XNOR U848 ( .A(n5316), .B(n5315), .Z(n5317) );
  XNOR U849 ( .A(in[1156]), .B(n5317), .Z(n6006) );
  XNOR U850 ( .A(n6296), .B(n6006), .Z(n8389) );
  XNOR U851 ( .A(in[132]), .B(n8389), .Z(n9442) );
  XOR U852 ( .A(in[36]), .B(in[676]), .Z(n5319) );
  XNOR U853 ( .A(in[356]), .B(in[1316]), .Z(n5318) );
  XNOR U854 ( .A(n5319), .B(n5318), .Z(n5320) );
  XOR U855 ( .A(in[996]), .B(n5320), .Z(n6104) );
  XOR U856 ( .A(in[1445]), .B(in[165]), .Z(n5322) );
  XNOR U857 ( .A(in[805]), .B(in[1125]), .Z(n5321) );
  XNOR U858 ( .A(n5322), .B(n5321), .Z(n5323) );
  XOR U859 ( .A(in[485]), .B(n5323), .Z(n5592) );
  XNOR U860 ( .A(n6104), .B(n5592), .Z(n8989) );
  XNOR U861 ( .A(in[1381]), .B(n8989), .Z(n9439) );
  NAND U862 ( .A(n9442), .B(n9439), .Z(n5324) );
  XNOR U863 ( .A(n6207), .B(n5324), .Z(out[1025]) );
  XNOR U864 ( .A(n5326), .B(n5325), .Z(n8440) );
  XNOR U865 ( .A(in[533]), .B(n8440), .Z(n6211) );
  XOR U866 ( .A(in[1348]), .B(in[68]), .Z(n5328) );
  XNOR U867 ( .A(in[1028]), .B(in[388]), .Z(n5327) );
  XNOR U868 ( .A(n5328), .B(n5327), .Z(n5329) );
  XOR U869 ( .A(in[708]), .B(n5329), .Z(n6300) );
  XOR U870 ( .A(in[1477]), .B(in[517]), .Z(n5331) );
  XNOR U871 ( .A(in[837]), .B(in[197]), .Z(n5330) );
  XNOR U872 ( .A(n5331), .B(n5330), .Z(n5332) );
  XNOR U873 ( .A(in[1157]), .B(n5332), .Z(n6009) );
  XNOR U874 ( .A(n6300), .B(n6009), .Z(n8393) );
  XNOR U875 ( .A(in[133]), .B(n8393), .Z(n9446) );
  XOR U876 ( .A(in[166]), .B(in[806]), .Z(n5334) );
  XNOR U877 ( .A(in[1126]), .B(in[486]), .Z(n5333) );
  XNOR U878 ( .A(n5334), .B(n5333), .Z(n5335) );
  XOR U879 ( .A(in[1446]), .B(n5335), .Z(n5605) );
  XOR U880 ( .A(in[37]), .B(in[677]), .Z(n5337) );
  XNOR U881 ( .A(in[357]), .B(in[1317]), .Z(n5336) );
  XNOR U882 ( .A(n5337), .B(n5336), .Z(n5338) );
  XOR U883 ( .A(in[997]), .B(n5338), .Z(n6107) );
  XNOR U884 ( .A(n5605), .B(n6107), .Z(n8992) );
  XNOR U885 ( .A(in[1382]), .B(n8992), .Z(n9443) );
  NAND U886 ( .A(n9446), .B(n9443), .Z(n5339) );
  XNOR U887 ( .A(n6211), .B(n5339), .Z(out[1026]) );
  XOR U888 ( .A(n5341), .B(n5340), .Z(n8444) );
  XNOR U889 ( .A(in[534]), .B(n8444), .Z(n6215) );
  XOR U890 ( .A(in[1349]), .B(in[69]), .Z(n5343) );
  XNOR U891 ( .A(in[1029]), .B(in[389]), .Z(n5342) );
  XNOR U892 ( .A(n5343), .B(n5342), .Z(n5344) );
  XOR U893 ( .A(in[709]), .B(n5344), .Z(n6304) );
  XOR U894 ( .A(in[1478]), .B(in[518]), .Z(n5346) );
  XNOR U895 ( .A(in[838]), .B(in[198]), .Z(n5345) );
  XNOR U896 ( .A(n5346), .B(n5345), .Z(n5347) );
  XNOR U897 ( .A(in[1158]), .B(n5347), .Z(n6012) );
  XNOR U898 ( .A(n6304), .B(n6012), .Z(n8397) );
  XNOR U899 ( .A(in[134]), .B(n8397), .Z(n9450) );
  XOR U900 ( .A(in[38]), .B(in[678]), .Z(n5349) );
  XNOR U901 ( .A(in[358]), .B(in[1318]), .Z(n5348) );
  XNOR U902 ( .A(n5349), .B(n5348), .Z(n5350) );
  XOR U903 ( .A(in[998]), .B(n5350), .Z(n6111) );
  XOR U904 ( .A(in[167]), .B(in[807]), .Z(n5352) );
  XNOR U905 ( .A(in[1127]), .B(in[487]), .Z(n5351) );
  XNOR U906 ( .A(n5352), .B(n5351), .Z(n5353) );
  XOR U907 ( .A(in[1447]), .B(n5353), .Z(n5618) );
  XNOR U908 ( .A(n6111), .B(n5618), .Z(n8771) );
  XNOR U909 ( .A(in[1383]), .B(n8771), .Z(n9447) );
  NAND U910 ( .A(n9450), .B(n9447), .Z(n5354) );
  XNOR U911 ( .A(n6215), .B(n5354), .Z(out[1027]) );
  XOR U912 ( .A(n5356), .B(n5355), .Z(n8448) );
  XNOR U913 ( .A(in[535]), .B(n8448), .Z(n6219) );
  XOR U914 ( .A(in[1350]), .B(in[70]), .Z(n5358) );
  XNOR U915 ( .A(in[1030]), .B(in[390]), .Z(n5357) );
  XNOR U916 ( .A(n5358), .B(n5357), .Z(n5359) );
  XOR U917 ( .A(in[710]), .B(n5359), .Z(n6308) );
  XOR U918 ( .A(in[199]), .B(in[1479]), .Z(n5361) );
  XNOR U919 ( .A(in[1159]), .B(in[839]), .Z(n5360) );
  XNOR U920 ( .A(n5361), .B(n5360), .Z(n5362) );
  XNOR U921 ( .A(in[519]), .B(n5362), .Z(n6015) );
  XNOR U922 ( .A(n6308), .B(n6015), .Z(n8401) );
  XNOR U923 ( .A(in[135]), .B(n8401), .Z(n9454) );
  XOR U924 ( .A(in[168]), .B(in[1448]), .Z(n5364) );
  XNOR U925 ( .A(in[1128]), .B(in[808]), .Z(n5363) );
  XNOR U926 ( .A(n5364), .B(n5363), .Z(n5365) );
  XOR U927 ( .A(in[488]), .B(n5365), .Z(n5631) );
  XOR U928 ( .A(in[39]), .B(in[679]), .Z(n5367) );
  XNOR U929 ( .A(in[359]), .B(in[1319]), .Z(n5366) );
  XNOR U930 ( .A(n5367), .B(n5366), .Z(n5368) );
  XOR U931 ( .A(in[999]), .B(n5368), .Z(n6115) );
  XNOR U932 ( .A(n5631), .B(n6115), .Z(n8774) );
  XNOR U933 ( .A(in[1384]), .B(n8774), .Z(n9451) );
  NAND U934 ( .A(n9454), .B(n9451), .Z(n5369) );
  XNOR U935 ( .A(n6219), .B(n5369), .Z(out[1028]) );
  XNOR U936 ( .A(n5371), .B(n5370), .Z(n8452) );
  XNOR U937 ( .A(in[536]), .B(n8452), .Z(n6223) );
  XOR U938 ( .A(in[1351]), .B(in[711]), .Z(n5373) );
  XNOR U939 ( .A(in[1031]), .B(in[391]), .Z(n5372) );
  XNOR U940 ( .A(n5373), .B(n5372), .Z(n5374) );
  XOR U941 ( .A(in[71]), .B(n5374), .Z(n6312) );
  XOR U942 ( .A(in[1480]), .B(in[520]), .Z(n5376) );
  XNOR U943 ( .A(in[840]), .B(in[200]), .Z(n5375) );
  XNOR U944 ( .A(n5376), .B(n5375), .Z(n5377) );
  XNOR U945 ( .A(in[1160]), .B(n5377), .Z(n6020) );
  XNOR U946 ( .A(n6312), .B(n6020), .Z(n8405) );
  XNOR U947 ( .A(in[136]), .B(n8405), .Z(n9458) );
  XOR U948 ( .A(in[680]), .B(in[1320]), .Z(n5379) );
  XNOR U949 ( .A(in[40]), .B(in[360]), .Z(n5378) );
  XNOR U950 ( .A(n5379), .B(n5378), .Z(n5380) );
  XOR U951 ( .A(in[1000]), .B(n5380), .Z(n6119) );
  XOR U952 ( .A(in[169]), .B(in[1449]), .Z(n5382) );
  XNOR U953 ( .A(in[1129]), .B(in[809]), .Z(n5381) );
  XNOR U954 ( .A(n5382), .B(n5381), .Z(n5383) );
  XOR U955 ( .A(in[489]), .B(n5383), .Z(n5644) );
  XNOR U956 ( .A(n6119), .B(n5644), .Z(n8781) );
  XNOR U957 ( .A(in[1385]), .B(n8781), .Z(n9455) );
  NAND U958 ( .A(n9458), .B(n9455), .Z(n5384) );
  XNOR U959 ( .A(n6223), .B(n5384), .Z(out[1029]) );
  XOR U960 ( .A(in[1341]), .B(in[61]), .Z(n5386) );
  XNOR U961 ( .A(in[701]), .B(in[381]), .Z(n5385) );
  XNOR U962 ( .A(n5386), .B(n5385), .Z(n5387) );
  XOR U963 ( .A(in[1021]), .B(n5387), .Z(n5701) );
  XNOR U964 ( .A(n5388), .B(n5701), .Z(n8407) );
  XNOR U965 ( .A(in[637]), .B(n8407), .Z(n7362) );
  XNOR U966 ( .A(n5390), .B(n5389), .Z(n8504) );
  XNOR U967 ( .A(in[228]), .B(n8504), .Z(n7666) );
  XOR U968 ( .A(in[1512]), .B(in[552]), .Z(n5392) );
  XNOR U969 ( .A(in[872]), .B(in[232]), .Z(n5391) );
  XNOR U970 ( .A(n5392), .B(n5391), .Z(n5393) );
  XOR U971 ( .A(in[1192]), .B(n5393), .Z(n6124) );
  XNOR U972 ( .A(n5394), .B(n6124), .Z(n8545) );
  XNOR U973 ( .A(in[1448]), .B(n8545), .Z(n7663) );
  NAND U974 ( .A(n7666), .B(n7663), .Z(n5395) );
  XNOR U975 ( .A(n7362), .B(n5395), .Z(out[102]) );
  XOR U976 ( .A(n5397), .B(n5396), .Z(n8456) );
  XNOR U977 ( .A(in[537]), .B(n8456), .Z(n6227) );
  XOR U978 ( .A(in[1352]), .B(in[712]), .Z(n5399) );
  XNOR U979 ( .A(in[1032]), .B(in[392]), .Z(n5398) );
  XNOR U980 ( .A(n5399), .B(n5398), .Z(n5400) );
  XOR U981 ( .A(in[72]), .B(n5400), .Z(n6317) );
  XOR U982 ( .A(in[1481]), .B(in[521]), .Z(n5402) );
  XNOR U983 ( .A(in[841]), .B(in[201]), .Z(n5401) );
  XNOR U984 ( .A(n5402), .B(n5401), .Z(n5403) );
  XNOR U985 ( .A(in[1161]), .B(n5403), .Z(n6023) );
  XNOR U986 ( .A(n6317), .B(n6023), .Z(n8409) );
  XNOR U987 ( .A(in[137]), .B(n8409), .Z(n9462) );
  XOR U988 ( .A(in[681]), .B(in[1321]), .Z(n5405) );
  XNOR U989 ( .A(in[41]), .B(in[361]), .Z(n5404) );
  XNOR U990 ( .A(n5405), .B(n5404), .Z(n5406) );
  XOR U991 ( .A(in[1001]), .B(n5406), .Z(n6123) );
  XOR U992 ( .A(in[170]), .B(in[1450]), .Z(n5408) );
  XNOR U993 ( .A(in[1130]), .B(in[810]), .Z(n5407) );
  XNOR U994 ( .A(n5408), .B(n5407), .Z(n5409) );
  XOR U995 ( .A(in[490]), .B(n5409), .Z(n5660) );
  XNOR U996 ( .A(n6123), .B(n5660), .Z(n8784) );
  XNOR U997 ( .A(in[1386]), .B(n8784), .Z(n9459) );
  NAND U998 ( .A(n9462), .B(n9459), .Z(n5410) );
  XNOR U999 ( .A(n6227), .B(n5410), .Z(out[1030]) );
  XOR U1000 ( .A(n5412), .B(n5411), .Z(n8460) );
  XNOR U1001 ( .A(in[538]), .B(n8460), .Z(n6231) );
  XOR U1002 ( .A(in[1353]), .B(in[393]), .Z(n5414) );
  XNOR U1003 ( .A(in[713]), .B(in[73]), .Z(n5413) );
  XNOR U1004 ( .A(n5414), .B(n5413), .Z(n5415) );
  XOR U1005 ( .A(in[1033]), .B(n5415), .Z(n6321) );
  XOR U1006 ( .A(in[1482]), .B(in[522]), .Z(n5417) );
  XNOR U1007 ( .A(in[842]), .B(in[202]), .Z(n5416) );
  XNOR U1008 ( .A(n5417), .B(n5416), .Z(n5418) );
  XNOR U1009 ( .A(in[1162]), .B(n5418), .Z(n6026) );
  XNOR U1010 ( .A(n6321), .B(n6026), .Z(n8413) );
  XNOR U1011 ( .A(in[138]), .B(n8413), .Z(n9466) );
  XOR U1012 ( .A(in[811]), .B(in[491]), .Z(n5420) );
  XNOR U1013 ( .A(in[1451]), .B(in[1131]), .Z(n5419) );
  XNOR U1014 ( .A(n5420), .B(n5419), .Z(n5421) );
  XOR U1015 ( .A(in[171]), .B(n5421), .Z(n5673) );
  XOR U1016 ( .A(in[682]), .B(in[1322]), .Z(n5423) );
  XNOR U1017 ( .A(in[42]), .B(in[362]), .Z(n5422) );
  XNOR U1018 ( .A(n5423), .B(n5422), .Z(n5424) );
  XOR U1019 ( .A(in[1002]), .B(n5424), .Z(n6128) );
  XNOR U1020 ( .A(n5673), .B(n6128), .Z(n8787) );
  XNOR U1021 ( .A(in[1387]), .B(n8787), .Z(n9463) );
  NAND U1022 ( .A(n9466), .B(n9463), .Z(n5425) );
  XNOR U1023 ( .A(n6231), .B(n5425), .Z(out[1031]) );
  XOR U1024 ( .A(n5427), .B(n5426), .Z(n8464) );
  XNOR U1025 ( .A(in[539]), .B(n8464), .Z(n6236) );
  XOR U1026 ( .A(in[1483]), .B(in[523]), .Z(n5429) );
  XNOR U1027 ( .A(in[843]), .B(in[203]), .Z(n5428) );
  XNOR U1028 ( .A(n5429), .B(n5428), .Z(n5430) );
  XOR U1029 ( .A(in[1163]), .B(n5430), .Z(n6029) );
  XOR U1030 ( .A(in[1354]), .B(in[714]), .Z(n5432) );
  XNOR U1031 ( .A(in[74]), .B(in[394]), .Z(n5431) );
  XNOR U1032 ( .A(n5432), .B(n5431), .Z(n5433) );
  XNOR U1033 ( .A(in[1034]), .B(n5433), .Z(n6325) );
  XNOR U1034 ( .A(n6029), .B(n6325), .Z(n8417) );
  XNOR U1035 ( .A(n8417), .B(in[139]), .Z(n9470) );
  XOR U1036 ( .A(in[812]), .B(in[492]), .Z(n5435) );
  XNOR U1037 ( .A(in[1452]), .B(in[1132]), .Z(n5434) );
  XNOR U1038 ( .A(n5435), .B(n5434), .Z(n5436) );
  XOR U1039 ( .A(in[172]), .B(n5436), .Z(n5693) );
  XOR U1040 ( .A(in[683]), .B(in[1323]), .Z(n5438) );
  XNOR U1041 ( .A(in[43]), .B(in[363]), .Z(n5437) );
  XNOR U1042 ( .A(n5438), .B(n5437), .Z(n5439) );
  XOR U1043 ( .A(in[1003]), .B(n5439), .Z(n6132) );
  XNOR U1044 ( .A(n5693), .B(n6132), .Z(n8790) );
  XNOR U1045 ( .A(in[1388]), .B(n8790), .Z(n9467) );
  NAND U1046 ( .A(n9470), .B(n9467), .Z(n5440) );
  XNOR U1047 ( .A(n6236), .B(n5440), .Z(out[1032]) );
  XNOR U1048 ( .A(n5442), .B(n5441), .Z(n8468) );
  XNOR U1049 ( .A(in[540]), .B(n8468), .Z(n6240) );
  XOR U1050 ( .A(in[1355]), .B(in[715]), .Z(n5444) );
  XNOR U1051 ( .A(in[1035]), .B(in[395]), .Z(n5443) );
  XNOR U1052 ( .A(n5444), .B(n5443), .Z(n5445) );
  XOR U1053 ( .A(in[75]), .B(n5445), .Z(n6329) );
  XOR U1054 ( .A(in[1484]), .B(in[524]), .Z(n5447) );
  XNOR U1055 ( .A(in[844]), .B(in[204]), .Z(n5446) );
  XNOR U1056 ( .A(n5447), .B(n5446), .Z(n5448) );
  XNOR U1057 ( .A(in[1164]), .B(n5448), .Z(n6032) );
  XNOR U1058 ( .A(n6329), .B(n6032), .Z(n8421) );
  XNOR U1059 ( .A(in[140]), .B(n8421), .Z(n9474) );
  XOR U1060 ( .A(in[813]), .B(in[493]), .Z(n5450) );
  XNOR U1061 ( .A(in[1453]), .B(in[1133]), .Z(n5449) );
  XNOR U1062 ( .A(n5450), .B(n5449), .Z(n5451) );
  XOR U1063 ( .A(in[173]), .B(n5451), .Z(n5706) );
  XOR U1064 ( .A(in[1324]), .B(in[44]), .Z(n5453) );
  XNOR U1065 ( .A(in[684]), .B(in[364]), .Z(n5452) );
  XNOR U1066 ( .A(n5453), .B(n5452), .Z(n5454) );
  XOR U1067 ( .A(in[1004]), .B(n5454), .Z(n6135) );
  XNOR U1068 ( .A(n5706), .B(n6135), .Z(n8793) );
  XNOR U1069 ( .A(in[1389]), .B(n8793), .Z(n9471) );
  NAND U1070 ( .A(n9474), .B(n9471), .Z(n5455) );
  XNOR U1071 ( .A(n6240), .B(n5455), .Z(out[1033]) );
  XNOR U1072 ( .A(n5457), .B(n5456), .Z(n8476) );
  XNOR U1073 ( .A(in[541]), .B(n8476), .Z(n6244) );
  XOR U1074 ( .A(in[76]), .B(in[1036]), .Z(n5459) );
  XNOR U1075 ( .A(in[716]), .B(in[396]), .Z(n5458) );
  XNOR U1076 ( .A(n5459), .B(n5458), .Z(n5460) );
  XOR U1077 ( .A(in[1356]), .B(n5460), .Z(n6333) );
  XOR U1078 ( .A(in[1485]), .B(in[525]), .Z(n5462) );
  XNOR U1079 ( .A(in[845]), .B(in[205]), .Z(n5461) );
  XNOR U1080 ( .A(n5462), .B(n5461), .Z(n5463) );
  XNOR U1081 ( .A(in[1165]), .B(n5463), .Z(n6035) );
  XNOR U1082 ( .A(n6333), .B(n6035), .Z(n8425) );
  XNOR U1083 ( .A(in[141]), .B(n8425), .Z(n9482) );
  XOR U1084 ( .A(in[814]), .B(in[494]), .Z(n5465) );
  XNOR U1085 ( .A(in[1454]), .B(in[1134]), .Z(n5464) );
  XNOR U1086 ( .A(n5465), .B(n5464), .Z(n5466) );
  XOR U1087 ( .A(in[174]), .B(n5466), .Z(n5719) );
  XOR U1088 ( .A(in[1325]), .B(in[45]), .Z(n5468) );
  XNOR U1089 ( .A(in[685]), .B(in[365]), .Z(n5467) );
  XNOR U1090 ( .A(n5468), .B(n5467), .Z(n5469) );
  XOR U1091 ( .A(in[1005]), .B(n5469), .Z(n6139) );
  XNOR U1092 ( .A(n5719), .B(n6139), .Z(n8796) );
  XNOR U1093 ( .A(in[1390]), .B(n8796), .Z(n9479) );
  NAND U1094 ( .A(n9482), .B(n9479), .Z(n5470) );
  XNOR U1095 ( .A(n6244), .B(n5470), .Z(out[1034]) );
  XNOR U1096 ( .A(n5472), .B(n5471), .Z(n8480) );
  XNOR U1097 ( .A(in[542]), .B(n8480), .Z(n6248) );
  XOR U1098 ( .A(in[77]), .B(in[1037]), .Z(n5474) );
  XNOR U1099 ( .A(in[717]), .B(in[397]), .Z(n5473) );
  XNOR U1100 ( .A(n5474), .B(n5473), .Z(n5475) );
  XOR U1101 ( .A(in[1357]), .B(n5475), .Z(n6337) );
  XOR U1102 ( .A(in[1486]), .B(in[526]), .Z(n5477) );
  XNOR U1103 ( .A(in[846]), .B(in[206]), .Z(n5476) );
  XNOR U1104 ( .A(n5477), .B(n5476), .Z(n5478) );
  XNOR U1105 ( .A(in[1166]), .B(n5478), .Z(n6038) );
  XNOR U1106 ( .A(n6337), .B(n6038), .Z(n8433) );
  XNOR U1107 ( .A(in[142]), .B(n8433), .Z(n9486) );
  XOR U1108 ( .A(in[1326]), .B(in[46]), .Z(n5480) );
  XNOR U1109 ( .A(in[686]), .B(in[366]), .Z(n5479) );
  XNOR U1110 ( .A(n5480), .B(n5479), .Z(n5481) );
  XOR U1111 ( .A(in[1006]), .B(n5481), .Z(n6143) );
  XOR U1112 ( .A(in[815]), .B(in[495]), .Z(n5483) );
  XNOR U1113 ( .A(in[1455]), .B(in[1135]), .Z(n5482) );
  XNOR U1114 ( .A(n5483), .B(n5482), .Z(n5484) );
  XOR U1115 ( .A(in[175]), .B(n5484), .Z(n5732) );
  XNOR U1116 ( .A(n6143), .B(n5732), .Z(n8799) );
  XNOR U1117 ( .A(in[1391]), .B(n8799), .Z(n9483) );
  NAND U1118 ( .A(n9486), .B(n9483), .Z(n5485) );
  XNOR U1119 ( .A(n6248), .B(n5485), .Z(out[1035]) );
  XNOR U1120 ( .A(n5487), .B(n5486), .Z(n8484) );
  XNOR U1121 ( .A(in[543]), .B(n8484), .Z(n6252) );
  XOR U1122 ( .A(in[78]), .B(in[1038]), .Z(n5489) );
  XNOR U1123 ( .A(in[718]), .B(in[398]), .Z(n5488) );
  XNOR U1124 ( .A(n5489), .B(n5488), .Z(n5490) );
  XOR U1125 ( .A(in[1358]), .B(n5490), .Z(n6341) );
  XOR U1126 ( .A(in[1487]), .B(in[527]), .Z(n5492) );
  XNOR U1127 ( .A(in[847]), .B(in[207]), .Z(n5491) );
  XNOR U1128 ( .A(n5492), .B(n5491), .Z(n5493) );
  XNOR U1129 ( .A(in[1167]), .B(n5493), .Z(n6041) );
  XNOR U1130 ( .A(n6341), .B(n6041), .Z(n8437) );
  XNOR U1131 ( .A(in[143]), .B(n8437), .Z(n9490) );
  XOR U1132 ( .A(in[1327]), .B(in[47]), .Z(n5495) );
  XNOR U1133 ( .A(in[687]), .B(in[367]), .Z(n5494) );
  XNOR U1134 ( .A(n5495), .B(n5494), .Z(n5496) );
  XOR U1135 ( .A(in[1007]), .B(n5496), .Z(n6147) );
  XOR U1136 ( .A(in[816]), .B(in[496]), .Z(n5498) );
  XNOR U1137 ( .A(in[1456]), .B(in[1136]), .Z(n5497) );
  XNOR U1138 ( .A(n5498), .B(n5497), .Z(n5499) );
  XOR U1139 ( .A(in[176]), .B(n5499), .Z(n5747) );
  XNOR U1140 ( .A(n6147), .B(n5747), .Z(n8802) );
  XNOR U1141 ( .A(in[1392]), .B(n8802), .Z(n9487) );
  NAND U1142 ( .A(n9490), .B(n9487), .Z(n5500) );
  XNOR U1143 ( .A(n6252), .B(n5500), .Z(out[1036]) );
  XNOR U1144 ( .A(n5502), .B(n5501), .Z(n8488) );
  XNOR U1145 ( .A(in[544]), .B(n8488), .Z(n6256) );
  XOR U1146 ( .A(in[79]), .B(in[1039]), .Z(n5504) );
  XNOR U1147 ( .A(in[719]), .B(in[399]), .Z(n5503) );
  XNOR U1148 ( .A(n5504), .B(n5503), .Z(n5505) );
  XOR U1149 ( .A(in[1359]), .B(n5505), .Z(n6345) );
  XOR U1150 ( .A(in[1488]), .B(in[528]), .Z(n5507) );
  XNOR U1151 ( .A(in[848]), .B(in[208]), .Z(n5506) );
  XNOR U1152 ( .A(n5507), .B(n5506), .Z(n5508) );
  XNOR U1153 ( .A(in[1168]), .B(n5508), .Z(n6044) );
  XNOR U1154 ( .A(n6345), .B(n6044), .Z(n8441) );
  XNOR U1155 ( .A(in[144]), .B(n8441), .Z(n9494) );
  XOR U1156 ( .A(in[1328]), .B(in[48]), .Z(n5510) );
  XNOR U1157 ( .A(in[688]), .B(in[368]), .Z(n5509) );
  XNOR U1158 ( .A(n5510), .B(n5509), .Z(n5511) );
  XOR U1159 ( .A(in[1008]), .B(n5511), .Z(n6151) );
  XOR U1160 ( .A(in[817]), .B(in[497]), .Z(n5513) );
  XNOR U1161 ( .A(in[1457]), .B(in[1137]), .Z(n5512) );
  XNOR U1162 ( .A(n5513), .B(n5512), .Z(n5514) );
  XOR U1163 ( .A(in[177]), .B(n5514), .Z(n5762) );
  XNOR U1164 ( .A(n6151), .B(n5762), .Z(n8805) );
  XNOR U1165 ( .A(in[1393]), .B(n8805), .Z(n9491) );
  NAND U1166 ( .A(n9494), .B(n9491), .Z(n5515) );
  XNOR U1167 ( .A(n6256), .B(n5515), .Z(out[1037]) );
  XNOR U1168 ( .A(n5517), .B(n5516), .Z(n8492) );
  XNOR U1169 ( .A(in[545]), .B(n8492), .Z(n6260) );
  XOR U1170 ( .A(in[80]), .B(in[1040]), .Z(n5519) );
  XNOR U1171 ( .A(in[720]), .B(in[400]), .Z(n5518) );
  XNOR U1172 ( .A(n5519), .B(n5518), .Z(n5520) );
  XOR U1173 ( .A(in[1360]), .B(n5520), .Z(n6349) );
  XOR U1174 ( .A(in[1489]), .B(in[529]), .Z(n5522) );
  XNOR U1175 ( .A(in[849]), .B(in[209]), .Z(n5521) );
  XNOR U1176 ( .A(n5522), .B(n5521), .Z(n5523) );
  XNOR U1177 ( .A(in[1169]), .B(n5523), .Z(n6047) );
  XNOR U1178 ( .A(n6349), .B(n6047), .Z(n8445) );
  XNOR U1179 ( .A(in[145]), .B(n8445), .Z(n9498) );
  XOR U1180 ( .A(in[818]), .B(in[498]), .Z(n5525) );
  XNOR U1181 ( .A(in[1458]), .B(in[1138]), .Z(n5524) );
  XNOR U1182 ( .A(n5525), .B(n5524), .Z(n5526) );
  XOR U1183 ( .A(in[178]), .B(n5526), .Z(n5777) );
  XOR U1184 ( .A(in[1329]), .B(in[49]), .Z(n5528) );
  XNOR U1185 ( .A(in[689]), .B(in[369]), .Z(n5527) );
  XNOR U1186 ( .A(n5528), .B(n5527), .Z(n5529) );
  XOR U1187 ( .A(in[1009]), .B(n5529), .Z(n6156) );
  XNOR U1188 ( .A(n5777), .B(n6156), .Z(n8808) );
  XNOR U1189 ( .A(in[1394]), .B(n8808), .Z(n9495) );
  NAND U1190 ( .A(n9498), .B(n9495), .Z(n5530) );
  XNOR U1191 ( .A(n6260), .B(n5530), .Z(out[1038]) );
  XOR U1192 ( .A(n8496), .B(in[546]), .Z(n6264) );
  XOR U1193 ( .A(in[81]), .B(in[1041]), .Z(n5532) );
  XNOR U1194 ( .A(in[721]), .B(in[401]), .Z(n5531) );
  XNOR U1195 ( .A(n5532), .B(n5531), .Z(n5533) );
  XOR U1196 ( .A(in[1361]), .B(n5533), .Z(n6353) );
  XOR U1197 ( .A(in[1490]), .B(in[530]), .Z(n5535) );
  XNOR U1198 ( .A(in[850]), .B(in[210]), .Z(n5534) );
  XNOR U1199 ( .A(n5535), .B(n5534), .Z(n5536) );
  XNOR U1200 ( .A(in[1170]), .B(n5536), .Z(n6051) );
  XNOR U1201 ( .A(n6353), .B(n6051), .Z(n8449) );
  XNOR U1202 ( .A(in[146]), .B(n8449), .Z(n9502) );
  XOR U1203 ( .A(in[1330]), .B(in[50]), .Z(n5538) );
  XNOR U1204 ( .A(in[690]), .B(in[370]), .Z(n5537) );
  XNOR U1205 ( .A(n5538), .B(n5537), .Z(n5539) );
  XOR U1206 ( .A(in[1010]), .B(n5539), .Z(n6160) );
  XOR U1207 ( .A(in[819]), .B(in[499]), .Z(n5541) );
  XNOR U1208 ( .A(in[1459]), .B(in[1139]), .Z(n5540) );
  XNOR U1209 ( .A(n5541), .B(n5540), .Z(n5542) );
  XOR U1210 ( .A(in[179]), .B(n5542), .Z(n5792) );
  XNOR U1211 ( .A(n6160), .B(n5792), .Z(n8815) );
  XNOR U1212 ( .A(in[1395]), .B(n8815), .Z(n9499) );
  NAND U1213 ( .A(n9502), .B(n9499), .Z(n5543) );
  XNOR U1214 ( .A(n6264), .B(n5543), .Z(out[1039]) );
  XOR U1215 ( .A(in[1342]), .B(in[62]), .Z(n5545) );
  XNOR U1216 ( .A(in[702]), .B(in[382]), .Z(n5544) );
  XNOR U1217 ( .A(n5545), .B(n5544), .Z(n5546) );
  XOR U1218 ( .A(in[1022]), .B(n5546), .Z(n5714) );
  XNOR U1219 ( .A(n5547), .B(n5714), .Z(n8411) );
  XNOR U1220 ( .A(in[638]), .B(n8411), .Z(n7364) );
  XOR U1221 ( .A(n5549), .B(n5548), .Z(n8508) );
  XNOR U1222 ( .A(in[229]), .B(n8508), .Z(n7680) );
  XOR U1223 ( .A(in[1513]), .B(in[553]), .Z(n5551) );
  XNOR U1224 ( .A(in[873]), .B(in[233]), .Z(n5550) );
  XNOR U1225 ( .A(n5551), .B(n5550), .Z(n5552) );
  XOR U1226 ( .A(in[1193]), .B(n5552), .Z(n6127) );
  XNOR U1227 ( .A(n5553), .B(n6127), .Z(n8549) );
  XNOR U1228 ( .A(in[1449]), .B(n8549), .Z(n7677) );
  NAND U1229 ( .A(n7680), .B(n7677), .Z(n5554) );
  XNOR U1230 ( .A(n7364), .B(n5554), .Z(out[103]) );
  XOR U1231 ( .A(n8500), .B(in[547]), .Z(n6268) );
  XOR U1232 ( .A(in[1042]), .B(in[402]), .Z(n5556) );
  XNOR U1233 ( .A(in[722]), .B(in[82]), .Z(n5555) );
  XNOR U1234 ( .A(n5556), .B(n5555), .Z(n5557) );
  XOR U1235 ( .A(in[1362]), .B(n5557), .Z(n6358) );
  XOR U1236 ( .A(in[851]), .B(in[1171]), .Z(n5559) );
  XNOR U1237 ( .A(in[1491]), .B(in[211]), .Z(n5558) );
  XNOR U1238 ( .A(n5559), .B(n5558), .Z(n5560) );
  XNOR U1239 ( .A(in[531]), .B(n5560), .Z(n6054) );
  XNOR U1240 ( .A(n6358), .B(n6054), .Z(n8453) );
  XNOR U1241 ( .A(in[147]), .B(n8453), .Z(n9506) );
  XOR U1242 ( .A(in[1331]), .B(in[51]), .Z(n5562) );
  XNOR U1243 ( .A(in[691]), .B(in[371]), .Z(n5561) );
  XNOR U1244 ( .A(n5562), .B(n5561), .Z(n5563) );
  XOR U1245 ( .A(in[1011]), .B(n5563), .Z(n6164) );
  XOR U1246 ( .A(in[820]), .B(in[500]), .Z(n5565) );
  XNOR U1247 ( .A(in[1460]), .B(in[1140]), .Z(n5564) );
  XNOR U1248 ( .A(n5565), .B(n5564), .Z(n5566) );
  XOR U1249 ( .A(in[180]), .B(n5566), .Z(n5807) );
  XNOR U1250 ( .A(n6164), .B(n5807), .Z(n8818) );
  XNOR U1251 ( .A(in[1396]), .B(n8818), .Z(n9503) );
  NAND U1252 ( .A(n9506), .B(n9503), .Z(n5567) );
  XNOR U1253 ( .A(n6268), .B(n5567), .Z(out[1040]) );
  XOR U1254 ( .A(n8504), .B(in[548]), .Z(n6272) );
  XOR U1255 ( .A(in[83]), .B(in[1043]), .Z(n5569) );
  XNOR U1256 ( .A(in[723]), .B(in[403]), .Z(n5568) );
  XNOR U1257 ( .A(n5569), .B(n5568), .Z(n5570) );
  XOR U1258 ( .A(in[1363]), .B(n5570), .Z(n6362) );
  XOR U1259 ( .A(in[852]), .B(in[1172]), .Z(n5572) );
  XNOR U1260 ( .A(in[1492]), .B(in[212]), .Z(n5571) );
  XNOR U1261 ( .A(n5572), .B(n5571), .Z(n5573) );
  XNOR U1262 ( .A(in[532]), .B(n5573), .Z(n6057) );
  XNOR U1263 ( .A(n6362), .B(n6057), .Z(n8457) );
  XNOR U1264 ( .A(in[148]), .B(n8457), .Z(n9510) );
  XOR U1265 ( .A(in[821]), .B(in[501]), .Z(n5575) );
  XNOR U1266 ( .A(in[1461]), .B(in[1141]), .Z(n5574) );
  XNOR U1267 ( .A(n5575), .B(n5574), .Z(n5576) );
  XOR U1268 ( .A(in[181]), .B(n5576), .Z(n5822) );
  XOR U1269 ( .A(in[1332]), .B(in[52]), .Z(n5578) );
  XNOR U1270 ( .A(in[692]), .B(in[372]), .Z(n5577) );
  XNOR U1271 ( .A(n5578), .B(n5577), .Z(n5579) );
  XOR U1272 ( .A(in[1012]), .B(n5579), .Z(n6168) );
  XNOR U1273 ( .A(n5822), .B(n6168), .Z(n8821) );
  XNOR U1274 ( .A(in[1397]), .B(n8821), .Z(n9507) );
  NAND U1275 ( .A(n9510), .B(n9507), .Z(n5580) );
  XNOR U1276 ( .A(n6272), .B(n5580), .Z(out[1041]) );
  XOR U1277 ( .A(n8508), .B(in[549]), .Z(n6277) );
  XOR U1278 ( .A(in[853]), .B(in[1173]), .Z(n5582) );
  XNOR U1279 ( .A(in[1493]), .B(in[213]), .Z(n5581) );
  XNOR U1280 ( .A(n5582), .B(n5581), .Z(n5583) );
  XNOR U1281 ( .A(in[533]), .B(n5583), .Z(n6060) );
  XNOR U1282 ( .A(n5584), .B(n6060), .Z(n8461) );
  XNOR U1283 ( .A(in[149]), .B(n8461), .Z(n9514) );
  XOR U1284 ( .A(in[822]), .B(in[502]), .Z(n5586) );
  XNOR U1285 ( .A(in[1462]), .B(in[1142]), .Z(n5585) );
  XNOR U1286 ( .A(n5586), .B(n5585), .Z(n5587) );
  XOR U1287 ( .A(in[182]), .B(n5587), .Z(n5836) );
  XOR U1288 ( .A(in[1333]), .B(in[53]), .Z(n5589) );
  XNOR U1289 ( .A(in[693]), .B(in[373]), .Z(n5588) );
  XNOR U1290 ( .A(n5589), .B(n5588), .Z(n5590) );
  XOR U1291 ( .A(in[1013]), .B(n5590), .Z(n6172) );
  XNOR U1292 ( .A(n5836), .B(n6172), .Z(n8824) );
  XNOR U1293 ( .A(in[1398]), .B(n8824), .Z(n9511) );
  NAND U1294 ( .A(n9514), .B(n9511), .Z(n5591) );
  XNOR U1295 ( .A(n6277), .B(n5591), .Z(out[1042]) );
  XNOR U1296 ( .A(n5593), .B(n5592), .Z(n8512) );
  XNOR U1297 ( .A(in[550]), .B(n8512), .Z(n6281) );
  XOR U1298 ( .A(in[854]), .B(in[1174]), .Z(n5595) );
  XNOR U1299 ( .A(in[1494]), .B(in[214]), .Z(n5594) );
  XNOR U1300 ( .A(n5595), .B(n5594), .Z(n5596) );
  XNOR U1301 ( .A(in[534]), .B(n5596), .Z(n6063) );
  XNOR U1302 ( .A(n5597), .B(n6063), .Z(n8465) );
  XNOR U1303 ( .A(in[150]), .B(n8465), .Z(n9518) );
  XOR U1304 ( .A(in[823]), .B(in[503]), .Z(n5599) );
  XNOR U1305 ( .A(in[1463]), .B(in[1143]), .Z(n5598) );
  XNOR U1306 ( .A(n5599), .B(n5598), .Z(n5600) );
  XOR U1307 ( .A(in[183]), .B(n5600), .Z(n5847) );
  XOR U1308 ( .A(in[1334]), .B(in[54]), .Z(n5602) );
  XNOR U1309 ( .A(in[694]), .B(in[374]), .Z(n5601) );
  XNOR U1310 ( .A(n5602), .B(n5601), .Z(n5603) );
  XOR U1311 ( .A(in[1014]), .B(n5603), .Z(n6176) );
  XNOR U1312 ( .A(n5847), .B(n6176), .Z(n8827) );
  XNOR U1313 ( .A(in[1399]), .B(n8827), .Z(n9515) );
  NAND U1314 ( .A(n9518), .B(n9515), .Z(n5604) );
  XNOR U1315 ( .A(n6281), .B(n5604), .Z(out[1043]) );
  XNOR U1316 ( .A(n5606), .B(n5605), .Z(n8520) );
  XNOR U1317 ( .A(in[551]), .B(n8520), .Z(n6285) );
  XOR U1318 ( .A(in[855]), .B(in[1175]), .Z(n5608) );
  XNOR U1319 ( .A(in[1495]), .B(in[215]), .Z(n5607) );
  XNOR U1320 ( .A(n5608), .B(n5607), .Z(n5609) );
  XNOR U1321 ( .A(in[535]), .B(n5609), .Z(n6066) );
  XNOR U1322 ( .A(n5610), .B(n6066), .Z(n8469) );
  XNOR U1323 ( .A(in[151]), .B(n8469), .Z(n9526) );
  XOR U1324 ( .A(in[1335]), .B(in[55]), .Z(n5612) );
  XNOR U1325 ( .A(in[695]), .B(in[375]), .Z(n5611) );
  XNOR U1326 ( .A(n5612), .B(n5611), .Z(n5613) );
  XOR U1327 ( .A(in[1015]), .B(n5613), .Z(n6180) );
  XOR U1328 ( .A(in[824]), .B(in[504]), .Z(n5615) );
  XNOR U1329 ( .A(in[1464]), .B(in[1144]), .Z(n5614) );
  XNOR U1330 ( .A(n5615), .B(n5614), .Z(n5616) );
  XOR U1331 ( .A(in[184]), .B(n5616), .Z(n5852) );
  XNOR U1332 ( .A(n6180), .B(n5852), .Z(n8830) );
  XNOR U1333 ( .A(in[1400]), .B(n8830), .Z(n9523) );
  NAND U1334 ( .A(n9526), .B(n9523), .Z(n5617) );
  XNOR U1335 ( .A(n6285), .B(n5617), .Z(out[1044]) );
  XNOR U1336 ( .A(n5619), .B(n5618), .Z(n8524) );
  XNOR U1337 ( .A(in[552]), .B(n8524), .Z(n6289) );
  XOR U1338 ( .A(in[856]), .B(in[1176]), .Z(n5621) );
  XNOR U1339 ( .A(in[1496]), .B(in[216]), .Z(n5620) );
  XNOR U1340 ( .A(n5621), .B(n5620), .Z(n5622) );
  XNOR U1341 ( .A(in[536]), .B(n5622), .Z(n6069) );
  XNOR U1342 ( .A(n5623), .B(n6069), .Z(n8477) );
  XNOR U1343 ( .A(in[152]), .B(n8477), .Z(n9530) );
  XOR U1344 ( .A(in[1336]), .B(in[56]), .Z(n5625) );
  XNOR U1345 ( .A(in[696]), .B(in[376]), .Z(n5624) );
  XNOR U1346 ( .A(n5625), .B(n5624), .Z(n5626) );
  XOR U1347 ( .A(in[1016]), .B(n5626), .Z(n6184) );
  XOR U1348 ( .A(in[825]), .B(in[505]), .Z(n5628) );
  XNOR U1349 ( .A(in[1465]), .B(in[1145]), .Z(n5627) );
  XNOR U1350 ( .A(n5628), .B(n5627), .Z(n5629) );
  XOR U1351 ( .A(in[185]), .B(n5629), .Z(n5863) );
  XNOR U1352 ( .A(n6184), .B(n5863), .Z(n8833) );
  XNOR U1353 ( .A(in[1401]), .B(n8833), .Z(n9527) );
  NAND U1354 ( .A(n9530), .B(n9527), .Z(n5630) );
  XNOR U1355 ( .A(n6289), .B(n5630), .Z(out[1045]) );
  XNOR U1356 ( .A(n5632), .B(n5631), .Z(n8528) );
  XNOR U1357 ( .A(in[553]), .B(n8528), .Z(n6293) );
  XOR U1358 ( .A(in[857]), .B(in[1177]), .Z(n5634) );
  XNOR U1359 ( .A(in[1497]), .B(in[217]), .Z(n5633) );
  XNOR U1360 ( .A(n5634), .B(n5633), .Z(n5635) );
  XNOR U1361 ( .A(in[537]), .B(n5635), .Z(n6072) );
  XNOR U1362 ( .A(n5636), .B(n6072), .Z(n8481) );
  XNOR U1363 ( .A(in[153]), .B(n8481), .Z(n9534) );
  XOR U1364 ( .A(in[1337]), .B(in[57]), .Z(n5638) );
  XNOR U1365 ( .A(in[697]), .B(in[377]), .Z(n5637) );
  XNOR U1366 ( .A(n5638), .B(n5637), .Z(n5639) );
  XOR U1367 ( .A(in[1017]), .B(n5639), .Z(n6188) );
  XOR U1368 ( .A(in[826]), .B(in[506]), .Z(n5641) );
  XNOR U1369 ( .A(in[1466]), .B(in[1146]), .Z(n5640) );
  XNOR U1370 ( .A(n5641), .B(n5640), .Z(n5642) );
  XOR U1371 ( .A(in[186]), .B(n5642), .Z(n5874) );
  XNOR U1372 ( .A(n6188), .B(n5874), .Z(n8836) );
  XNOR U1373 ( .A(in[1402]), .B(n8836), .Z(n9531) );
  NAND U1374 ( .A(n9534), .B(n9531), .Z(n5643) );
  XNOR U1375 ( .A(n6293), .B(n5643), .Z(out[1046]) );
  XNOR U1376 ( .A(n5645), .B(n5644), .Z(n8532) );
  XNOR U1377 ( .A(in[554]), .B(n8532), .Z(n6297) );
  XOR U1378 ( .A(in[858]), .B(in[1178]), .Z(n5647) );
  XNOR U1379 ( .A(in[1498]), .B(in[218]), .Z(n5646) );
  XNOR U1380 ( .A(n5647), .B(n5646), .Z(n5648) );
  XNOR U1381 ( .A(in[538]), .B(n5648), .Z(n6075) );
  XNOR U1382 ( .A(n5649), .B(n6075), .Z(n8485) );
  XNOR U1383 ( .A(in[154]), .B(n8485), .Z(n9538) );
  XOR U1384 ( .A(in[1338]), .B(in[58]), .Z(n5651) );
  XNOR U1385 ( .A(in[698]), .B(in[378]), .Z(n5650) );
  XNOR U1386 ( .A(n5651), .B(n5650), .Z(n5652) );
  XOR U1387 ( .A(in[1018]), .B(n5652), .Z(n6192) );
  XOR U1388 ( .A(in[827]), .B(in[507]), .Z(n5654) );
  XNOR U1389 ( .A(in[1467]), .B(in[1147]), .Z(n5653) );
  XNOR U1390 ( .A(n5654), .B(n5653), .Z(n5655) );
  XOR U1391 ( .A(in[187]), .B(n5655), .Z(n5879) );
  XNOR U1392 ( .A(n6192), .B(n5879), .Z(n8839) );
  XNOR U1393 ( .A(in[1403]), .B(n8839), .Z(n9535) );
  NAND U1394 ( .A(n9538), .B(n9535), .Z(n5656) );
  XNOR U1395 ( .A(n6297), .B(n5656), .Z(out[1047]) );
  XOR U1396 ( .A(in[1579]), .B(in[619]), .Z(n5658) );
  XNOR U1397 ( .A(in[939]), .B(in[299]), .Z(n5657) );
  XNOR U1398 ( .A(n5658), .B(n5657), .Z(n5659) );
  XOR U1399 ( .A(in[1259]), .B(n5659), .Z(n6201) );
  XNOR U1400 ( .A(n5660), .B(n6201), .Z(n8536) );
  XNOR U1401 ( .A(in[555]), .B(n8536), .Z(n6301) );
  XOR U1402 ( .A(in[859]), .B(in[1179]), .Z(n5662) );
  XNOR U1403 ( .A(in[1499]), .B(in[219]), .Z(n5661) );
  XNOR U1404 ( .A(n5662), .B(n5661), .Z(n5663) );
  XNOR U1405 ( .A(in[539]), .B(n5663), .Z(n6078) );
  XNOR U1406 ( .A(n5664), .B(n6078), .Z(n8489) );
  XNOR U1407 ( .A(in[155]), .B(n8489), .Z(n9542) );
  XOR U1408 ( .A(in[828]), .B(in[508]), .Z(n5666) );
  XNOR U1409 ( .A(in[1468]), .B(in[1148]), .Z(n5665) );
  XNOR U1410 ( .A(n5666), .B(n5665), .Z(n5667) );
  XOR U1411 ( .A(in[188]), .B(n5667), .Z(n5884) );
  XNOR U1412 ( .A(n5668), .B(n5884), .Z(n8842) );
  XNOR U1413 ( .A(in[1404]), .B(n8842), .Z(n9539) );
  NAND U1414 ( .A(n9542), .B(n9539), .Z(n5669) );
  XNOR U1415 ( .A(n6301), .B(n5669), .Z(out[1048]) );
  XOR U1416 ( .A(in[1580]), .B(in[620]), .Z(n5671) );
  XNOR U1417 ( .A(in[940]), .B(in[300]), .Z(n5670) );
  XNOR U1418 ( .A(n5671), .B(n5670), .Z(n5672) );
  XOR U1419 ( .A(in[1260]), .B(n5672), .Z(n6205) );
  XNOR U1420 ( .A(n5673), .B(n6205), .Z(n8540) );
  XNOR U1421 ( .A(in[556]), .B(n8540), .Z(n6305) );
  XOR U1422 ( .A(in[860]), .B(in[1180]), .Z(n5675) );
  XNOR U1423 ( .A(in[1500]), .B(in[220]), .Z(n5674) );
  XNOR U1424 ( .A(n5675), .B(n5674), .Z(n5676) );
  XNOR U1425 ( .A(in[540]), .B(n5676), .Z(n6082) );
  XNOR U1426 ( .A(n5677), .B(n6082), .Z(n8493) );
  XNOR U1427 ( .A(in[156]), .B(n8493), .Z(n9546) );
  XNOR U1428 ( .A(n5679), .B(n5678), .Z(n8849) );
  XNOR U1429 ( .A(in[1405]), .B(n8849), .Z(n9543) );
  NAND U1430 ( .A(n9546), .B(n9543), .Z(n5680) );
  XNOR U1431 ( .A(n6305), .B(n5680), .Z(out[1049]) );
  XOR U1432 ( .A(in[1343]), .B(in[63]), .Z(n5682) );
  XNOR U1433 ( .A(in[703]), .B(in[383]), .Z(n5681) );
  XNOR U1434 ( .A(n5682), .B(n5681), .Z(n5683) );
  XOR U1435 ( .A(in[1023]), .B(n5683), .Z(n5727) );
  XNOR U1436 ( .A(n5684), .B(n5727), .Z(n8415) );
  XNOR U1437 ( .A(in[639]), .B(n8415), .Z(n7366) );
  XOR U1438 ( .A(in[230]), .B(n8512), .Z(n7696) );
  XOR U1439 ( .A(in[874]), .B(in[1194]), .Z(n5686) );
  XNOR U1440 ( .A(in[1514]), .B(in[234]), .Z(n5685) );
  XNOR U1441 ( .A(n5686), .B(n5685), .Z(n5687) );
  XOR U1442 ( .A(in[554]), .B(n5687), .Z(n6131) );
  XNOR U1443 ( .A(n5688), .B(n6131), .Z(n8553) );
  XNOR U1444 ( .A(in[1450]), .B(n8553), .Z(n7693) );
  NAND U1445 ( .A(n7696), .B(n7693), .Z(n5689) );
  XNOR U1446 ( .A(n7366), .B(n5689), .Z(out[104]) );
  XOR U1447 ( .A(in[1581]), .B(in[621]), .Z(n5691) );
  XNOR U1448 ( .A(in[941]), .B(in[301]), .Z(n5690) );
  XNOR U1449 ( .A(n5691), .B(n5690), .Z(n5692) );
  XOR U1450 ( .A(in[1261]), .B(n5692), .Z(n6209) );
  XNOR U1451 ( .A(n5693), .B(n6209), .Z(n8544) );
  XNOR U1452 ( .A(in[557]), .B(n8544), .Z(n6309) );
  XOR U1453 ( .A(in[861]), .B(in[1181]), .Z(n5695) );
  XNOR U1454 ( .A(in[1501]), .B(in[221]), .Z(n5694) );
  XNOR U1455 ( .A(n5695), .B(n5694), .Z(n5696) );
  XNOR U1456 ( .A(in[541]), .B(n5696), .Z(n6085) );
  XNOR U1457 ( .A(n5697), .B(n6085), .Z(n8497) );
  XNOR U1458 ( .A(in[157]), .B(n8497), .Z(n9550) );
  XOR U1459 ( .A(in[830]), .B(in[510]), .Z(n5699) );
  XNOR U1460 ( .A(in[1470]), .B(in[1150]), .Z(n5698) );
  XNOR U1461 ( .A(n5699), .B(n5698), .Z(n5700) );
  XOR U1462 ( .A(in[190]), .B(n5700), .Z(n5890) );
  XNOR U1463 ( .A(n5701), .B(n5890), .Z(n8852) );
  XNOR U1464 ( .A(in[1406]), .B(n8852), .Z(n9547) );
  NAND U1465 ( .A(n9550), .B(n9547), .Z(n5702) );
  XNOR U1466 ( .A(n6309), .B(n5702), .Z(out[1050]) );
  XOR U1467 ( .A(in[1582]), .B(in[622]), .Z(n5704) );
  XNOR U1468 ( .A(in[942]), .B(in[302]), .Z(n5703) );
  XNOR U1469 ( .A(n5704), .B(n5703), .Z(n5705) );
  XOR U1470 ( .A(in[1262]), .B(n5705), .Z(n6213) );
  XNOR U1471 ( .A(n5706), .B(n6213), .Z(n8548) );
  XNOR U1472 ( .A(in[558]), .B(n8548), .Z(n6313) );
  XOR U1473 ( .A(in[862]), .B(in[1182]), .Z(n5708) );
  XNOR U1474 ( .A(in[1502]), .B(in[222]), .Z(n5707) );
  XNOR U1475 ( .A(n5708), .B(n5707), .Z(n5709) );
  XNOR U1476 ( .A(in[542]), .B(n5709), .Z(n6088) );
  XNOR U1477 ( .A(n5710), .B(n6088), .Z(n8501) );
  XNOR U1478 ( .A(in[158]), .B(n8501), .Z(n9554) );
  XOR U1479 ( .A(in[831]), .B(in[511]), .Z(n5712) );
  XNOR U1480 ( .A(in[1471]), .B(in[1151]), .Z(n5711) );
  XNOR U1481 ( .A(n5712), .B(n5711), .Z(n5713) );
  XOR U1482 ( .A(in[191]), .B(n5713), .Z(n5895) );
  XNOR U1483 ( .A(n5714), .B(n5895), .Z(n8855) );
  XNOR U1484 ( .A(in[1407]), .B(n8855), .Z(n9551) );
  NAND U1485 ( .A(n9554), .B(n9551), .Z(n5715) );
  XNOR U1486 ( .A(n6313), .B(n5715), .Z(out[1051]) );
  XOR U1487 ( .A(in[1583]), .B(in[623]), .Z(n5717) );
  XNOR U1488 ( .A(in[943]), .B(in[303]), .Z(n5716) );
  XNOR U1489 ( .A(n5717), .B(n5716), .Z(n5718) );
  XOR U1490 ( .A(in[1263]), .B(n5718), .Z(n6217) );
  XNOR U1491 ( .A(n5719), .B(n6217), .Z(n8552) );
  XNOR U1492 ( .A(in[559]), .B(n8552), .Z(n6318) );
  XOR U1493 ( .A(in[863]), .B(in[1183]), .Z(n5721) );
  XNOR U1494 ( .A(in[1503]), .B(in[223]), .Z(n5720) );
  XNOR U1495 ( .A(n5721), .B(n5720), .Z(n5722) );
  XNOR U1496 ( .A(in[543]), .B(n5722), .Z(n6091) );
  XNOR U1497 ( .A(n5723), .B(n6091), .Z(n8505) );
  XNOR U1498 ( .A(in[159]), .B(n8505), .Z(n9558) );
  XOR U1499 ( .A(in[768]), .B(in[1088]), .Z(n5725) );
  XNOR U1500 ( .A(in[448]), .B(in[1408]), .Z(n5724) );
  XNOR U1501 ( .A(n5725), .B(n5724), .Z(n5726) );
  XOR U1502 ( .A(in[128]), .B(n5726), .Z(n5903) );
  XNOR U1503 ( .A(n5727), .B(n5903), .Z(n8858) );
  XNOR U1504 ( .A(in[1344]), .B(n8858), .Z(n9555) );
  NAND U1505 ( .A(n9558), .B(n9555), .Z(n5728) );
  XNOR U1506 ( .A(n6318), .B(n5728), .Z(out[1052]) );
  XOR U1507 ( .A(in[1584]), .B(in[624]), .Z(n5730) );
  XNOR U1508 ( .A(in[944]), .B(in[304]), .Z(n5729) );
  XNOR U1509 ( .A(n5730), .B(n5729), .Z(n5731) );
  XOR U1510 ( .A(in[1264]), .B(n5731), .Z(n6221) );
  XNOR U1511 ( .A(n5732), .B(n6221), .Z(n8556) );
  XNOR U1512 ( .A(in[560]), .B(n8556), .Z(n6322) );
  XOR U1513 ( .A(in[224]), .B(in[864]), .Z(n5734) );
  XNOR U1514 ( .A(in[1184]), .B(in[1504]), .Z(n5733) );
  XNOR U1515 ( .A(n5734), .B(n5733), .Z(n5735) );
  XNOR U1516 ( .A(in[544]), .B(n5735), .Z(n6094) );
  XNOR U1517 ( .A(n5736), .B(n6094), .Z(n8509) );
  XNOR U1518 ( .A(in[160]), .B(n8509), .Z(n9562) );
  XOR U1519 ( .A(in[1280]), .B(in[640]), .Z(n5738) );
  XNOR U1520 ( .A(in[960]), .B(in[320]), .Z(n5737) );
  XNOR U1521 ( .A(n5738), .B(n5737), .Z(n5739) );
  XOR U1522 ( .A(in[0]), .B(n5739), .Z(n5830) );
  XOR U1523 ( .A(in[769]), .B(in[1089]), .Z(n5741) );
  XNOR U1524 ( .A(in[449]), .B(in[1409]), .Z(n5740) );
  XNOR U1525 ( .A(n5741), .B(n5740), .Z(n5742) );
  XOR U1526 ( .A(in[129]), .B(n5742), .Z(n5908) );
  XNOR U1527 ( .A(n5830), .B(n5908), .Z(n8861) );
  XNOR U1528 ( .A(in[1345]), .B(n8861), .Z(n9559) );
  NAND U1529 ( .A(n9562), .B(n9559), .Z(n5743) );
  XNOR U1530 ( .A(n6322), .B(n5743), .Z(out[1053]) );
  XOR U1531 ( .A(in[1585]), .B(in[625]), .Z(n5745) );
  XNOR U1532 ( .A(in[945]), .B(in[305]), .Z(n5744) );
  XNOR U1533 ( .A(n5745), .B(n5744), .Z(n5746) );
  XOR U1534 ( .A(in[1265]), .B(n5746), .Z(n6225) );
  XNOR U1535 ( .A(n5747), .B(n6225), .Z(n8564) );
  XNOR U1536 ( .A(in[561]), .B(n8564), .Z(n6326) );
  XOR U1537 ( .A(in[225]), .B(in[865]), .Z(n5749) );
  XNOR U1538 ( .A(in[1185]), .B(in[1505]), .Z(n5748) );
  XNOR U1539 ( .A(n5749), .B(n5748), .Z(n5750) );
  XNOR U1540 ( .A(in[545]), .B(n5750), .Z(n6097) );
  XNOR U1541 ( .A(n5751), .B(n6097), .Z(n8513) );
  XNOR U1542 ( .A(in[161]), .B(n8513), .Z(n9570) );
  XOR U1543 ( .A(in[1]), .B(in[641]), .Z(n5753) );
  XNOR U1544 ( .A(in[961]), .B(in[321]), .Z(n5752) );
  XNOR U1545 ( .A(n5753), .B(n5752), .Z(n5754) );
  XOR U1546 ( .A(in[1281]), .B(n5754), .Z(n5897) );
  XOR U1547 ( .A(in[1090]), .B(in[450]), .Z(n5756) );
  XNOR U1548 ( .A(in[130]), .B(in[770]), .Z(n5755) );
  XNOR U1549 ( .A(n5756), .B(n5755), .Z(n5757) );
  XOR U1550 ( .A(in[1410]), .B(n5757), .Z(n5913) );
  XNOR U1551 ( .A(n5897), .B(n5913), .Z(n8864) );
  XNOR U1552 ( .A(in[1346]), .B(n8864), .Z(n9567) );
  NAND U1553 ( .A(n9570), .B(n9567), .Z(n5758) );
  XNOR U1554 ( .A(n6326), .B(n5758), .Z(out[1054]) );
  XOR U1555 ( .A(in[1586]), .B(in[626]), .Z(n5760) );
  XNOR U1556 ( .A(in[946]), .B(in[306]), .Z(n5759) );
  XNOR U1557 ( .A(n5760), .B(n5759), .Z(n5761) );
  XOR U1558 ( .A(in[1266]), .B(n5761), .Z(n6229) );
  XNOR U1559 ( .A(n5762), .B(n6229), .Z(n8568) );
  XNOR U1560 ( .A(in[562]), .B(n8568), .Z(n6330) );
  XOR U1561 ( .A(in[1186]), .B(in[1506]), .Z(n5764) );
  XNOR U1562 ( .A(in[546]), .B(in[866]), .Z(n5763) );
  XNOR U1563 ( .A(n5764), .B(n5763), .Z(n5765) );
  XNOR U1564 ( .A(in[226]), .B(n5765), .Z(n6100) );
  XNOR U1565 ( .A(n5766), .B(n6100), .Z(n8521) );
  XNOR U1566 ( .A(in[162]), .B(n8521), .Z(n9574) );
  XOR U1567 ( .A(in[771]), .B(in[1091]), .Z(n5768) );
  XNOR U1568 ( .A(in[451]), .B(in[1411]), .Z(n5767) );
  XNOR U1569 ( .A(n5768), .B(n5767), .Z(n5769) );
  XOR U1570 ( .A(in[131]), .B(n5769), .Z(n5918) );
  XOR U1571 ( .A(in[2]), .B(in[642]), .Z(n5771) );
  XNOR U1572 ( .A(in[962]), .B(in[322]), .Z(n5770) );
  XNOR U1573 ( .A(n5771), .B(n5770), .Z(n5772) );
  XOR U1574 ( .A(in[1282]), .B(n5772), .Z(n5950) );
  XNOR U1575 ( .A(n5918), .B(n5950), .Z(n8867) );
  XNOR U1576 ( .A(in[1347]), .B(n8867), .Z(n9571) );
  NAND U1577 ( .A(n9574), .B(n9571), .Z(n5773) );
  XNOR U1578 ( .A(n6330), .B(n5773), .Z(out[1055]) );
  XOR U1579 ( .A(in[1587]), .B(in[627]), .Z(n5775) );
  XNOR U1580 ( .A(in[947]), .B(in[307]), .Z(n5774) );
  XNOR U1581 ( .A(n5775), .B(n5774), .Z(n5776) );
  XOR U1582 ( .A(in[1267]), .B(n5776), .Z(n6234) );
  XNOR U1583 ( .A(n5777), .B(n6234), .Z(n8572) );
  XNOR U1584 ( .A(in[563]), .B(n8572), .Z(n6334) );
  XOR U1585 ( .A(in[1187]), .B(in[1507]), .Z(n5779) );
  XNOR U1586 ( .A(in[547]), .B(in[867]), .Z(n5778) );
  XNOR U1587 ( .A(n5779), .B(n5778), .Z(n5780) );
  XNOR U1588 ( .A(in[227]), .B(n5780), .Z(n6103) );
  XNOR U1589 ( .A(n5781), .B(n6103), .Z(n8525) );
  XNOR U1590 ( .A(in[163]), .B(n8525), .Z(n9578) );
  XOR U1591 ( .A(in[323]), .B(in[643]), .Z(n5783) );
  XNOR U1592 ( .A(in[963]), .B(in[3]), .Z(n5782) );
  XNOR U1593 ( .A(n5783), .B(n5782), .Z(n5784) );
  XOR U1594 ( .A(in[1283]), .B(n5784), .Z(n5996) );
  XOR U1595 ( .A(in[772]), .B(in[1092]), .Z(n5786) );
  XNOR U1596 ( .A(in[452]), .B(in[1412]), .Z(n5785) );
  XNOR U1597 ( .A(n5786), .B(n5785), .Z(n5787) );
  XOR U1598 ( .A(in[132]), .B(n5787), .Z(n5923) );
  XNOR U1599 ( .A(n5996), .B(n5923), .Z(n8870) );
  XNOR U1600 ( .A(in[1348]), .B(n8870), .Z(n9575) );
  NAND U1601 ( .A(n9578), .B(n9575), .Z(n5788) );
  XNOR U1602 ( .A(n6334), .B(n5788), .Z(out[1056]) );
  XOR U1603 ( .A(in[1588]), .B(in[628]), .Z(n5790) );
  XNOR U1604 ( .A(in[948]), .B(in[308]), .Z(n5789) );
  XNOR U1605 ( .A(n5790), .B(n5789), .Z(n5791) );
  XOR U1606 ( .A(in[1268]), .B(n5791), .Z(n6238) );
  XNOR U1607 ( .A(n5792), .B(n6238), .Z(n8576) );
  XNOR U1608 ( .A(in[564]), .B(n8576), .Z(n6338) );
  XOR U1609 ( .A(in[1188]), .B(in[1508]), .Z(n5794) );
  XNOR U1610 ( .A(in[548]), .B(in[868]), .Z(n5793) );
  XNOR U1611 ( .A(n5794), .B(n5793), .Z(n5795) );
  XOR U1612 ( .A(in[228]), .B(n5795), .Z(n6106) );
  XNOR U1613 ( .A(n6106), .B(n5796), .Z(n8529) );
  XNOR U1614 ( .A(in[164]), .B(n8529), .Z(n9582) );
  XOR U1615 ( .A(in[324]), .B(in[644]), .Z(n5798) );
  XNOR U1616 ( .A(in[964]), .B(in[4]), .Z(n5797) );
  XNOR U1617 ( .A(n5798), .B(n5797), .Z(n5799) );
  XOR U1618 ( .A(in[1284]), .B(n5799), .Z(n6004) );
  XOR U1619 ( .A(in[773]), .B(in[1093]), .Z(n5801) );
  XNOR U1620 ( .A(in[453]), .B(in[1413]), .Z(n5800) );
  XNOR U1621 ( .A(n5801), .B(n5800), .Z(n5802) );
  XOR U1622 ( .A(in[133]), .B(n5802), .Z(n5928) );
  XNOR U1623 ( .A(n6004), .B(n5928), .Z(n8873) );
  XNOR U1624 ( .A(in[1349]), .B(n8873), .Z(n9579) );
  NAND U1625 ( .A(n9582), .B(n9579), .Z(n5803) );
  XNOR U1626 ( .A(n6338), .B(n5803), .Z(out[1057]) );
  XOR U1627 ( .A(in[1589]), .B(in[629]), .Z(n5805) );
  XNOR U1628 ( .A(in[949]), .B(in[309]), .Z(n5804) );
  XNOR U1629 ( .A(n5805), .B(n5804), .Z(n5806) );
  XOR U1630 ( .A(in[1269]), .B(n5806), .Z(n6242) );
  XNOR U1631 ( .A(n5807), .B(n6242), .Z(n8580) );
  XNOR U1632 ( .A(in[565]), .B(n8580), .Z(n6342) );
  XOR U1633 ( .A(in[1189]), .B(in[1509]), .Z(n5809) );
  XNOR U1634 ( .A(in[549]), .B(in[869]), .Z(n5808) );
  XNOR U1635 ( .A(n5809), .B(n5808), .Z(n5810) );
  XNOR U1636 ( .A(in[229]), .B(n5810), .Z(n6110) );
  XNOR U1637 ( .A(n5811), .B(n6110), .Z(n8533) );
  XNOR U1638 ( .A(in[165]), .B(n8533), .Z(n9586) );
  XOR U1639 ( .A(in[774]), .B(in[1094]), .Z(n5813) );
  XNOR U1640 ( .A(in[454]), .B(in[1414]), .Z(n5812) );
  XNOR U1641 ( .A(n5813), .B(n5812), .Z(n5814) );
  XOR U1642 ( .A(in[134]), .B(n5814), .Z(n5933) );
  XOR U1643 ( .A(in[325]), .B(in[645]), .Z(n5816) );
  XNOR U1644 ( .A(in[965]), .B(in[5]), .Z(n5815) );
  XNOR U1645 ( .A(n5816), .B(n5815), .Z(n5817) );
  XOR U1646 ( .A(in[1285]), .B(n5817), .Z(n6007) );
  XNOR U1647 ( .A(n5933), .B(n6007), .Z(n8876) );
  XNOR U1648 ( .A(in[1350]), .B(n8876), .Z(n9583) );
  NAND U1649 ( .A(n9586), .B(n9583), .Z(n5818) );
  XNOR U1650 ( .A(n6342), .B(n5818), .Z(out[1058]) );
  XOR U1651 ( .A(in[1590]), .B(in[630]), .Z(n5820) );
  XNOR U1652 ( .A(in[950]), .B(in[310]), .Z(n5819) );
  XNOR U1653 ( .A(n5820), .B(n5819), .Z(n5821) );
  XOR U1654 ( .A(in[1270]), .B(n5821), .Z(n6246) );
  XNOR U1655 ( .A(n5822), .B(n6246), .Z(n8584) );
  XNOR U1656 ( .A(in[566]), .B(n8584), .Z(n6346) );
  XOR U1657 ( .A(in[166]), .B(n8537), .Z(n9590) );
  XOR U1658 ( .A(in[775]), .B(in[1095]), .Z(n5824) );
  XNOR U1659 ( .A(in[455]), .B(in[1415]), .Z(n5823) );
  XNOR U1660 ( .A(n5824), .B(n5823), .Z(n5825) );
  XOR U1661 ( .A(in[135]), .B(n5825), .Z(n5938) );
  XOR U1662 ( .A(in[326]), .B(in[6]), .Z(n5827) );
  XNOR U1663 ( .A(in[966]), .B(in[646]), .Z(n5826) );
  XNOR U1664 ( .A(n5827), .B(n5826), .Z(n5828) );
  XOR U1665 ( .A(in[1286]), .B(n5828), .Z(n6010) );
  XNOR U1666 ( .A(n5938), .B(n6010), .Z(n8887) );
  XNOR U1667 ( .A(in[1351]), .B(n8887), .Z(n9587) );
  NAND U1668 ( .A(n9590), .B(n9587), .Z(n5829) );
  XNOR U1669 ( .A(n6346), .B(n5829), .Z(out[1059]) );
  XNOR U1670 ( .A(n5831), .B(n5830), .Z(n8419) );
  XNOR U1671 ( .A(in[576]), .B(n8419), .Z(n7368) );
  XOR U1672 ( .A(in[231]), .B(n8520), .Z(n7710) );
  XNOR U1673 ( .A(in[1451]), .B(n8557), .Z(n7707) );
  NAND U1674 ( .A(n7710), .B(n7707), .Z(n5832) );
  XNOR U1675 ( .A(n7368), .B(n5832), .Z(out[105]) );
  XOR U1676 ( .A(in[1591]), .B(in[631]), .Z(n5834) );
  XNOR U1677 ( .A(in[951]), .B(in[311]), .Z(n5833) );
  XNOR U1678 ( .A(n5834), .B(n5833), .Z(n5835) );
  XOR U1679 ( .A(in[1271]), .B(n5835), .Z(n6250) );
  XNOR U1680 ( .A(n5836), .B(n6250), .Z(n8588) );
  XNOR U1681 ( .A(in[567]), .B(n8588), .Z(n6350) );
  XOR U1682 ( .A(in[167]), .B(n8541), .Z(n9594) );
  XOR U1683 ( .A(in[327]), .B(in[7]), .Z(n5838) );
  XNOR U1684 ( .A(in[967]), .B(in[647]), .Z(n5837) );
  XNOR U1685 ( .A(n5838), .B(n5837), .Z(n5839) );
  XOR U1686 ( .A(in[1287]), .B(n5839), .Z(n6013) );
  XOR U1687 ( .A(in[776]), .B(in[1096]), .Z(n5841) );
  XNOR U1688 ( .A(in[456]), .B(in[1416]), .Z(n5840) );
  XNOR U1689 ( .A(n5841), .B(n5840), .Z(n5842) );
  XOR U1690 ( .A(in[136]), .B(n5842), .Z(n5943) );
  XNOR U1691 ( .A(n6013), .B(n5943), .Z(n8890) );
  XNOR U1692 ( .A(in[1352]), .B(n8890), .Z(n9591) );
  NAND U1693 ( .A(n9594), .B(n9591), .Z(n5843) );
  XNOR U1694 ( .A(n6350), .B(n5843), .Z(out[1060]) );
  XOR U1695 ( .A(in[632]), .B(in[1592]), .Z(n5845) );
  XNOR U1696 ( .A(in[1272]), .B(in[312]), .Z(n5844) );
  XNOR U1697 ( .A(n5845), .B(n5844), .Z(n5846) );
  XOR U1698 ( .A(in[952]), .B(n5846), .Z(n6254) );
  XNOR U1699 ( .A(n5847), .B(n6254), .Z(n8592) );
  XNOR U1700 ( .A(in[568]), .B(n8592), .Z(n6354) );
  XOR U1701 ( .A(in[168]), .B(n8545), .Z(n9598) );
  XNOR U1702 ( .A(in[1353]), .B(n8893), .Z(n9595) );
  NAND U1703 ( .A(n9598), .B(n9595), .Z(n5848) );
  XNOR U1704 ( .A(n6354), .B(n5848), .Z(out[1061]) );
  XOR U1705 ( .A(in[633]), .B(in[1593]), .Z(n5850) );
  XNOR U1706 ( .A(in[1273]), .B(in[313]), .Z(n5849) );
  XNOR U1707 ( .A(n5850), .B(n5849), .Z(n5851) );
  XOR U1708 ( .A(in[953]), .B(n5851), .Z(n6258) );
  XNOR U1709 ( .A(n5852), .B(n6258), .Z(n8596) );
  XNOR U1710 ( .A(in[569]), .B(n8596), .Z(n6359) );
  XOR U1711 ( .A(in[169]), .B(n8549), .Z(n9602) );
  XOR U1712 ( .A(in[329]), .B(in[969]), .Z(n5854) );
  XNOR U1713 ( .A(in[9]), .B(in[649]), .Z(n5853) );
  XNOR U1714 ( .A(n5854), .B(n5853), .Z(n5855) );
  XOR U1715 ( .A(in[1289]), .B(n5855), .Z(n6021) );
  XOR U1716 ( .A(in[778]), .B(in[1098]), .Z(n5857) );
  XNOR U1717 ( .A(in[458]), .B(in[1418]), .Z(n5856) );
  XNOR U1718 ( .A(n5857), .B(n5856), .Z(n5858) );
  XOR U1719 ( .A(in[138]), .B(n5858), .Z(n5956) );
  XNOR U1720 ( .A(n6021), .B(n5956), .Z(n8896) );
  XNOR U1721 ( .A(in[1354]), .B(n8896), .Z(n9599) );
  NAND U1722 ( .A(n9602), .B(n9599), .Z(n5859) );
  XNOR U1723 ( .A(n6359), .B(n5859), .Z(out[1062]) );
  XOR U1724 ( .A(in[634]), .B(in[1594]), .Z(n5861) );
  XNOR U1725 ( .A(in[1274]), .B(in[314]), .Z(n5860) );
  XNOR U1726 ( .A(n5861), .B(n5860), .Z(n5862) );
  XOR U1727 ( .A(in[954]), .B(n5862), .Z(n6262) );
  XNOR U1728 ( .A(n5863), .B(n6262), .Z(n8600) );
  XNOR U1729 ( .A(in[570]), .B(n8600), .Z(n6363) );
  XOR U1730 ( .A(in[170]), .B(n8553), .Z(n9606) );
  XOR U1731 ( .A(in[1290]), .B(in[650]), .Z(n5865) );
  XNOR U1732 ( .A(in[970]), .B(in[330]), .Z(n5864) );
  XNOR U1733 ( .A(n5865), .B(n5864), .Z(n5866) );
  XOR U1734 ( .A(in[10]), .B(n5866), .Z(n6024) );
  XOR U1735 ( .A(in[1419]), .B(in[779]), .Z(n5868) );
  XNOR U1736 ( .A(in[1099]), .B(in[459]), .Z(n5867) );
  XNOR U1737 ( .A(n5868), .B(n5867), .Z(n5869) );
  XOR U1738 ( .A(in[139]), .B(n5869), .Z(n5961) );
  XNOR U1739 ( .A(n6024), .B(n5961), .Z(n8899) );
  XNOR U1740 ( .A(in[1355]), .B(n8899), .Z(n9603) );
  NAND U1741 ( .A(n9606), .B(n9603), .Z(n5870) );
  XNOR U1742 ( .A(n6363), .B(n5870), .Z(out[1063]) );
  XOR U1743 ( .A(in[955]), .B(in[1275]), .Z(n5872) );
  XNOR U1744 ( .A(in[1595]), .B(in[315]), .Z(n5871) );
  XNOR U1745 ( .A(n5872), .B(n5871), .Z(n5873) );
  XNOR U1746 ( .A(in[635]), .B(n5873), .Z(n6266) );
  XNOR U1747 ( .A(n5874), .B(n6266), .Z(n8610) );
  XNOR U1748 ( .A(in[571]), .B(n8610), .Z(n6365) );
  NOR U1749 ( .A(n6108), .B(n6503), .Z(n5875) );
  XNOR U1750 ( .A(n6365), .B(n5875), .Z(out[1064]) );
  XOR U1751 ( .A(in[956]), .B(in[1276]), .Z(n5877) );
  XNOR U1752 ( .A(in[1596]), .B(in[316]), .Z(n5876) );
  XNOR U1753 ( .A(n5877), .B(n5876), .Z(n5878) );
  XNOR U1754 ( .A(in[636]), .B(n5878), .Z(n6270) );
  XNOR U1755 ( .A(n5879), .B(n6270), .Z(n8614) );
  XNOR U1756 ( .A(in[572]), .B(n8614), .Z(n6367) );
  NOR U1757 ( .A(n6112), .B(n6507), .Z(n5880) );
  XNOR U1758 ( .A(n6367), .B(n5880), .Z(out[1065]) );
  XOR U1759 ( .A(in[957]), .B(in[1277]), .Z(n5882) );
  XNOR U1760 ( .A(in[1597]), .B(in[317]), .Z(n5881) );
  XNOR U1761 ( .A(n5882), .B(n5881), .Z(n5883) );
  XNOR U1762 ( .A(in[637]), .B(n5883), .Z(n6275) );
  XNOR U1763 ( .A(n5884), .B(n6275), .Z(n8618) );
  XNOR U1764 ( .A(in[573]), .B(n8618), .Z(n6369) );
  NOR U1765 ( .A(n6117), .B(n6511), .Z(n5885) );
  XNOR U1766 ( .A(n6369), .B(n5885), .Z(out[1066]) );
  XOR U1767 ( .A(in[574]), .B(n8622), .Z(n6371) );
  NOR U1768 ( .A(n6121), .B(n6515), .Z(n5886) );
  XNOR U1769 ( .A(n6371), .B(n5886), .Z(out[1067]) );
  XOR U1770 ( .A(in[959]), .B(in[1279]), .Z(n5888) );
  XNOR U1771 ( .A(in[1599]), .B(in[319]), .Z(n5887) );
  XNOR U1772 ( .A(n5888), .B(n5887), .Z(n5889) );
  XNOR U1773 ( .A(in[639]), .B(n5889), .Z(n6283) );
  XNOR U1774 ( .A(n5890), .B(n6283), .Z(n8344) );
  XNOR U1775 ( .A(in[575]), .B(n8344), .Z(n6373) );
  NOR U1776 ( .A(n6125), .B(n6520), .Z(n5891) );
  XNOR U1777 ( .A(n6373), .B(n5891), .Z(out[1068]) );
  XOR U1778 ( .A(in[896]), .B(in[1216]), .Z(n5893) );
  XNOR U1779 ( .A(in[1536]), .B(in[256]), .Z(n5892) );
  XNOR U1780 ( .A(n5893), .B(n5892), .Z(n5894) );
  XNOR U1781 ( .A(in[576]), .B(n5894), .Z(n6287) );
  XNOR U1782 ( .A(n5895), .B(n6287), .Z(n8348) );
  XNOR U1783 ( .A(in[512]), .B(n8348), .Z(n6375) );
  NOR U1784 ( .A(n6129), .B(n6524), .Z(n5896) );
  XNOR U1785 ( .A(n6375), .B(n5896), .Z(out[1069]) );
  XNOR U1786 ( .A(n5898), .B(n5897), .Z(n8423) );
  XNOR U1787 ( .A(in[577]), .B(n8423), .Z(n7370) );
  XOR U1788 ( .A(in[232]), .B(n8524), .Z(n7724) );
  XNOR U1789 ( .A(in[1452]), .B(n8565), .Z(n7721) );
  NAND U1790 ( .A(n7724), .B(n7721), .Z(n5899) );
  XNOR U1791 ( .A(n7370), .B(n5899), .Z(out[106]) );
  XOR U1792 ( .A(in[897]), .B(in[1217]), .Z(n5901) );
  XNOR U1793 ( .A(in[1537]), .B(in[257]), .Z(n5900) );
  XNOR U1794 ( .A(n5901), .B(n5900), .Z(n5902) );
  XNOR U1795 ( .A(in[577]), .B(n5902), .Z(n6291) );
  XNOR U1796 ( .A(n5903), .B(n6291), .Z(n8352) );
  XNOR U1797 ( .A(in[513]), .B(n8352), .Z(n6377) );
  NOR U1798 ( .A(n6133), .B(n6528), .Z(n5904) );
  XNOR U1799 ( .A(n6377), .B(n5904), .Z(out[1070]) );
  XOR U1800 ( .A(in[1538]), .B(in[578]), .Z(n5906) );
  XNOR U1801 ( .A(in[898]), .B(in[258]), .Z(n5905) );
  XNOR U1802 ( .A(n5906), .B(n5905), .Z(n5907) );
  XNOR U1803 ( .A(in[1218]), .B(n5907), .Z(n6295) );
  XNOR U1804 ( .A(n5908), .B(n6295), .Z(n8356) );
  XNOR U1805 ( .A(in[514]), .B(n8356), .Z(n6379) );
  NOR U1806 ( .A(n6137), .B(n6532), .Z(n5909) );
  XNOR U1807 ( .A(n6379), .B(n5909), .Z(out[1071]) );
  XOR U1808 ( .A(in[1539]), .B(in[579]), .Z(n5911) );
  XNOR U1809 ( .A(in[899]), .B(in[259]), .Z(n5910) );
  XNOR U1810 ( .A(n5911), .B(n5910), .Z(n5912) );
  XNOR U1811 ( .A(in[1219]), .B(n5912), .Z(n6299) );
  XNOR U1812 ( .A(n5913), .B(n6299), .Z(n8360) );
  XNOR U1813 ( .A(in[515]), .B(n8360), .Z(n6383) );
  NOR U1814 ( .A(n6141), .B(n6536), .Z(n5914) );
  XNOR U1815 ( .A(n6383), .B(n5914), .Z(out[1072]) );
  XOR U1816 ( .A(in[1540]), .B(in[580]), .Z(n5916) );
  XNOR U1817 ( .A(in[900]), .B(in[260]), .Z(n5915) );
  XNOR U1818 ( .A(n5916), .B(n5915), .Z(n5917) );
  XNOR U1819 ( .A(in[1220]), .B(n5917), .Z(n6303) );
  XNOR U1820 ( .A(n5918), .B(n6303), .Z(n8364) );
  XNOR U1821 ( .A(in[516]), .B(n8364), .Z(n6385) );
  NOR U1822 ( .A(n6145), .B(n6540), .Z(n5919) );
  XNOR U1823 ( .A(n6385), .B(n5919), .Z(out[1073]) );
  XOR U1824 ( .A(in[1541]), .B(in[581]), .Z(n5921) );
  XNOR U1825 ( .A(in[901]), .B(in[261]), .Z(n5920) );
  XNOR U1826 ( .A(n5921), .B(n5920), .Z(n5922) );
  XNOR U1827 ( .A(in[1221]), .B(n5922), .Z(n6307) );
  XNOR U1828 ( .A(n5923), .B(n6307), .Z(n8368) );
  XNOR U1829 ( .A(in[517]), .B(n8368), .Z(n6387) );
  NOR U1830 ( .A(n6149), .B(n6544), .Z(n5924) );
  XNOR U1831 ( .A(n6387), .B(n5924), .Z(out[1074]) );
  XOR U1832 ( .A(in[1542]), .B(in[582]), .Z(n5926) );
  XNOR U1833 ( .A(in[902]), .B(in[262]), .Z(n5925) );
  XNOR U1834 ( .A(n5926), .B(n5925), .Z(n5927) );
  XNOR U1835 ( .A(in[1222]), .B(n5927), .Z(n6311) );
  XNOR U1836 ( .A(n5928), .B(n6311), .Z(n8372) );
  XNOR U1837 ( .A(in[518]), .B(n8372), .Z(n6389) );
  NOR U1838 ( .A(n6153), .B(n6548), .Z(n5929) );
  XNOR U1839 ( .A(n6389), .B(n5929), .Z(out[1075]) );
  XOR U1840 ( .A(in[1543]), .B(in[583]), .Z(n5931) );
  XNOR U1841 ( .A(in[903]), .B(in[263]), .Z(n5930) );
  XNOR U1842 ( .A(n5931), .B(n5930), .Z(n5932) );
  XNOR U1843 ( .A(in[1223]), .B(n5932), .Z(n6316) );
  XNOR U1844 ( .A(n5933), .B(n6316), .Z(n8376) );
  XNOR U1845 ( .A(in[519]), .B(n8376), .Z(n6391) );
  NOR U1846 ( .A(n6158), .B(n6552), .Z(n5934) );
  XNOR U1847 ( .A(n6391), .B(n5934), .Z(out[1076]) );
  XOR U1848 ( .A(in[1544]), .B(in[584]), .Z(n5936) );
  XNOR U1849 ( .A(in[904]), .B(in[264]), .Z(n5935) );
  XNOR U1850 ( .A(n5936), .B(n5935), .Z(n5937) );
  XNOR U1851 ( .A(in[1224]), .B(n5937), .Z(n6320) );
  XNOR U1852 ( .A(n5938), .B(n6320), .Z(n8380) );
  XNOR U1853 ( .A(in[520]), .B(n8380), .Z(n6393) );
  NOR U1854 ( .A(n6162), .B(n6556), .Z(n5939) );
  XNOR U1855 ( .A(n6393), .B(n5939), .Z(out[1077]) );
  XOR U1856 ( .A(in[1545]), .B(in[585]), .Z(n5941) );
  XNOR U1857 ( .A(in[905]), .B(in[265]), .Z(n5940) );
  XNOR U1858 ( .A(n5941), .B(n5940), .Z(n5942) );
  XNOR U1859 ( .A(in[1225]), .B(n5942), .Z(n6324) );
  XNOR U1860 ( .A(n5943), .B(n6324), .Z(n8388) );
  XNOR U1861 ( .A(in[521]), .B(n8388), .Z(n6395) );
  NOR U1862 ( .A(n6166), .B(n6561), .Z(n5944) );
  XNOR U1863 ( .A(n6395), .B(n5944), .Z(out[1078]) );
  XOR U1864 ( .A(in[1546]), .B(in[586]), .Z(n5946) );
  XNOR U1865 ( .A(in[906]), .B(in[266]), .Z(n5945) );
  XNOR U1866 ( .A(n5946), .B(n5945), .Z(n5947) );
  XNOR U1867 ( .A(in[1226]), .B(n5947), .Z(n6328) );
  XNOR U1868 ( .A(n5948), .B(n6328), .Z(n8392) );
  XNOR U1869 ( .A(in[522]), .B(n8392), .Z(n6397) );
  NOR U1870 ( .A(n6170), .B(n6565), .Z(n5949) );
  XNOR U1871 ( .A(n6397), .B(n5949), .Z(out[1079]) );
  XNOR U1872 ( .A(n5951), .B(n5950), .Z(n8431) );
  XNOR U1873 ( .A(in[578]), .B(n8431), .Z(n7372) );
  XOR U1874 ( .A(in[233]), .B(n8528), .Z(n7738) );
  XNOR U1875 ( .A(in[1453]), .B(n8569), .Z(n7735) );
  NAND U1876 ( .A(n7738), .B(n7735), .Z(n5952) );
  XNOR U1877 ( .A(n7372), .B(n5952), .Z(out[107]) );
  XOR U1878 ( .A(in[1547]), .B(in[587]), .Z(n5954) );
  XNOR U1879 ( .A(in[907]), .B(in[267]), .Z(n5953) );
  XNOR U1880 ( .A(n5954), .B(n5953), .Z(n5955) );
  XNOR U1881 ( .A(in[1227]), .B(n5955), .Z(n6332) );
  XNOR U1882 ( .A(n5956), .B(n6332), .Z(n8396) );
  XNOR U1883 ( .A(in[523]), .B(n8396), .Z(n6399) );
  NOR U1884 ( .A(n6174), .B(n6569), .Z(n5957) );
  XNOR U1885 ( .A(n6399), .B(n5957), .Z(out[1080]) );
  XOR U1886 ( .A(in[1548]), .B(in[588]), .Z(n5959) );
  XNOR U1887 ( .A(in[908]), .B(in[268]), .Z(n5958) );
  XNOR U1888 ( .A(n5959), .B(n5958), .Z(n5960) );
  XNOR U1889 ( .A(in[1228]), .B(n5960), .Z(n6336) );
  XNOR U1890 ( .A(n5961), .B(n6336), .Z(n8400) );
  XNOR U1891 ( .A(in[524]), .B(n8400), .Z(n6401) );
  NOR U1892 ( .A(n6178), .B(n6573), .Z(n5962) );
  XNOR U1893 ( .A(n6401), .B(n5962), .Z(out[1081]) );
  XOR U1894 ( .A(in[1549]), .B(in[589]), .Z(n5964) );
  XNOR U1895 ( .A(in[909]), .B(in[269]), .Z(n5963) );
  XNOR U1896 ( .A(n5964), .B(n5963), .Z(n5965) );
  XOR U1897 ( .A(in[1229]), .B(n5965), .Z(n6340) );
  XNOR U1898 ( .A(n6340), .B(n5966), .Z(n8404) );
  XNOR U1899 ( .A(in[525]), .B(n8404), .Z(n6404) );
  NOR U1900 ( .A(n6182), .B(n6577), .Z(n5967) );
  XNOR U1901 ( .A(n6404), .B(n5967), .Z(out[1082]) );
  XOR U1902 ( .A(in[1550]), .B(in[590]), .Z(n5969) );
  XNOR U1903 ( .A(in[910]), .B(in[270]), .Z(n5968) );
  XNOR U1904 ( .A(n5969), .B(n5968), .Z(n5970) );
  XOR U1905 ( .A(in[1230]), .B(n5970), .Z(n6344) );
  XNOR U1906 ( .A(n6344), .B(n5971), .Z(n8408) );
  XNOR U1907 ( .A(in[526]), .B(n8408), .Z(n6406) );
  NOR U1908 ( .A(n6186), .B(n6581), .Z(n5972) );
  XNOR U1909 ( .A(n6406), .B(n5972), .Z(out[1083]) );
  XOR U1910 ( .A(in[1551]), .B(in[591]), .Z(n5974) );
  XNOR U1911 ( .A(in[911]), .B(in[271]), .Z(n5973) );
  XNOR U1912 ( .A(n5974), .B(n5973), .Z(n5975) );
  XOR U1913 ( .A(in[1231]), .B(n5975), .Z(n6348) );
  XNOR U1914 ( .A(n6348), .B(n5976), .Z(n8412) );
  XNOR U1915 ( .A(in[527]), .B(n8412), .Z(n6408) );
  NOR U1916 ( .A(n6190), .B(n6585), .Z(n5977) );
  XNOR U1917 ( .A(n6408), .B(n5977), .Z(out[1084]) );
  XOR U1918 ( .A(in[1552]), .B(in[592]), .Z(n5979) );
  XNOR U1919 ( .A(in[912]), .B(in[272]), .Z(n5978) );
  XNOR U1920 ( .A(n5979), .B(n5978), .Z(n5980) );
  XNOR U1921 ( .A(in[1232]), .B(n5980), .Z(n6352) );
  XNOR U1922 ( .A(n5981), .B(n6352), .Z(n8416) );
  XNOR U1923 ( .A(in[528]), .B(n8416), .Z(n6410) );
  NOR U1924 ( .A(n6194), .B(n6589), .Z(n5982) );
  XNOR U1925 ( .A(n6410), .B(n5982), .Z(out[1085]) );
  XOR U1926 ( .A(in[1553]), .B(in[593]), .Z(n5984) );
  XNOR U1927 ( .A(in[913]), .B(in[273]), .Z(n5983) );
  XNOR U1928 ( .A(n5984), .B(n5983), .Z(n5985) );
  XNOR U1929 ( .A(in[1233]), .B(n5985), .Z(n6357) );
  XNOR U1930 ( .A(n5986), .B(n6357), .Z(n8420) );
  XNOR U1931 ( .A(in[529]), .B(n8420), .Z(n6412) );
  NOR U1932 ( .A(n6197), .B(n6593), .Z(n5987) );
  XNOR U1933 ( .A(n6412), .B(n5987), .Z(out[1086]) );
  XOR U1934 ( .A(in[1554]), .B(in[594]), .Z(n5989) );
  XNOR U1935 ( .A(in[914]), .B(in[274]), .Z(n5988) );
  XNOR U1936 ( .A(n5989), .B(n5988), .Z(n5990) );
  XNOR U1937 ( .A(in[1234]), .B(n5990), .Z(n6361) );
  XNOR U1938 ( .A(n5991), .B(n6361), .Z(n8424) );
  XNOR U1939 ( .A(in[530]), .B(n8424), .Z(n6414) );
  NOR U1940 ( .A(n6199), .B(n6597), .Z(n5992) );
  XNOR U1941 ( .A(n6414), .B(n5992), .Z(out[1087]) );
  XOR U1942 ( .A(in[957]), .B(n8407), .Z(n6416) );
  NOR U1943 ( .A(n6203), .B(n9438), .Z(n5993) );
  XNOR U1944 ( .A(n6416), .B(n5993), .Z(out[1088]) );
  XOR U1945 ( .A(in[958]), .B(n8411), .Z(n6418) );
  NOR U1946 ( .A(n6207), .B(n9442), .Z(n5994) );
  XNOR U1947 ( .A(n6418), .B(n5994), .Z(out[1089]) );
  XOR U1948 ( .A(n5996), .B(n5995), .Z(n8435) );
  XNOR U1949 ( .A(in[579]), .B(n8435), .Z(n7374) );
  XOR U1950 ( .A(in[234]), .B(n8532), .Z(n7754) );
  XNOR U1951 ( .A(in[1454]), .B(n8573), .Z(n7751) );
  NAND U1952 ( .A(n7754), .B(n7751), .Z(n5997) );
  XNOR U1953 ( .A(n7374), .B(n5997), .Z(out[108]) );
  XOR U1954 ( .A(in[959]), .B(n8415), .Z(n6420) );
  NOR U1955 ( .A(n6211), .B(n9446), .Z(n5998) );
  XNOR U1956 ( .A(n6420), .B(n5998), .Z(out[1090]) );
  XOR U1957 ( .A(in[896]), .B(n8419), .Z(n6422) );
  NOR U1958 ( .A(n6215), .B(n9450), .Z(n5999) );
  XNOR U1959 ( .A(n6422), .B(n5999), .Z(out[1091]) );
  XOR U1960 ( .A(in[897]), .B(n8423), .Z(n6425) );
  NOR U1961 ( .A(n6219), .B(n9454), .Z(n6000) );
  XNOR U1962 ( .A(n6425), .B(n6000), .Z(out[1092]) );
  XOR U1963 ( .A(in[898]), .B(n8431), .Z(n6427) );
  NOR U1964 ( .A(n6223), .B(n9458), .Z(n6001) );
  XNOR U1965 ( .A(n6427), .B(n6001), .Z(out[1093]) );
  XOR U1966 ( .A(in[899]), .B(n8435), .Z(n6429) );
  NOR U1967 ( .A(n6227), .B(n9462), .Z(n6002) );
  XNOR U1968 ( .A(n6429), .B(n6002), .Z(out[1094]) );
  XNOR U1969 ( .A(n6004), .B(n6003), .Z(n8439) );
  XNOR U1970 ( .A(in[900]), .B(n8439), .Z(n6431) );
  NOR U1971 ( .A(n6231), .B(n9466), .Z(n6005) );
  XNOR U1972 ( .A(n6431), .B(n6005), .Z(out[1095]) );
  XNOR U1973 ( .A(n6007), .B(n6006), .Z(n8443) );
  XNOR U1974 ( .A(in[901]), .B(n8443), .Z(n6433) );
  NOR U1975 ( .A(n6236), .B(n9470), .Z(n6008) );
  XNOR U1976 ( .A(n6433), .B(n6008), .Z(out[1096]) );
  XNOR U1977 ( .A(n6010), .B(n6009), .Z(n8447) );
  XNOR U1978 ( .A(in[902]), .B(n8447), .Z(n6435) );
  NOR U1979 ( .A(n6240), .B(n9474), .Z(n6011) );
  XNOR U1980 ( .A(n6435), .B(n6011), .Z(out[1097]) );
  XNOR U1981 ( .A(n6013), .B(n6012), .Z(n8451) );
  XNOR U1982 ( .A(in[903]), .B(n8451), .Z(n6437) );
  NOR U1983 ( .A(n6244), .B(n9482), .Z(n6014) );
  XNOR U1984 ( .A(n6437), .B(n6014), .Z(out[1098]) );
  XNOR U1985 ( .A(n6016), .B(n6015), .Z(n8455) );
  XNOR U1986 ( .A(in[904]), .B(n8455), .Z(n6439) );
  NOR U1987 ( .A(n6248), .B(n9486), .Z(n6017) );
  XNOR U1988 ( .A(n6439), .B(n6017), .Z(out[1099]) );
  XOR U1989 ( .A(in[580]), .B(n8439), .Z(n7376) );
  XOR U1990 ( .A(in[235]), .B(n8536), .Z(n7778) );
  XNOR U1991 ( .A(in[1455]), .B(n8577), .Z(n7775) );
  NAND U1992 ( .A(n7778), .B(n7775), .Z(n6018) );
  XNOR U1993 ( .A(n7376), .B(n6018), .Z(out[109]) );
  XOR U1994 ( .A(in[200]), .B(n8380), .Z(n8728) );
  XNOR U1995 ( .A(in[1420]), .B(n8421), .Z(n8727) );
  XOR U1996 ( .A(n8927), .B(in[1043]), .Z(n7439) );
  NAND U1997 ( .A(n8727), .B(n7439), .Z(n6019) );
  XNOR U1998 ( .A(n8728), .B(n6019), .Z(out[10]) );
  XNOR U1999 ( .A(n6021), .B(n6020), .Z(n8459) );
  XNOR U2000 ( .A(in[905]), .B(n8459), .Z(n6441) );
  NOR U2001 ( .A(n6252), .B(n9490), .Z(n6022) );
  XNOR U2002 ( .A(n6441), .B(n6022), .Z(out[1100]) );
  XNOR U2003 ( .A(n6024), .B(n6023), .Z(n8463) );
  XNOR U2004 ( .A(in[906]), .B(n8463), .Z(n6443) );
  NOR U2005 ( .A(n6256), .B(n9494), .Z(n6025) );
  XNOR U2006 ( .A(n6443), .B(n6025), .Z(out[1101]) );
  XNOR U2007 ( .A(n6027), .B(n6026), .Z(n8467) );
  XNOR U2008 ( .A(in[907]), .B(n8467), .Z(n6446) );
  NOR U2009 ( .A(n6260), .B(n9498), .Z(n6028) );
  XNOR U2010 ( .A(n6446), .B(n6028), .Z(out[1102]) );
  XOR U2011 ( .A(n6030), .B(n6029), .Z(n8475) );
  XNOR U2012 ( .A(in[908]), .B(n8475), .Z(n6448) );
  NOR U2013 ( .A(n6264), .B(n9502), .Z(n6031) );
  XNOR U2014 ( .A(n6448), .B(n6031), .Z(out[1103]) );
  XNOR U2015 ( .A(n6033), .B(n6032), .Z(n8479) );
  XNOR U2016 ( .A(in[909]), .B(n8479), .Z(n6450) );
  NOR U2017 ( .A(n6268), .B(n9506), .Z(n6034) );
  XNOR U2018 ( .A(n6450), .B(n6034), .Z(out[1104]) );
  XOR U2019 ( .A(n6036), .B(n6035), .Z(n8483) );
  XNOR U2020 ( .A(in[910]), .B(n8483), .Z(n6452) );
  NOR U2021 ( .A(n6272), .B(n9510), .Z(n6037) );
  XNOR U2022 ( .A(n6452), .B(n6037), .Z(out[1105]) );
  XOR U2023 ( .A(n6039), .B(n6038), .Z(n8487) );
  XNOR U2024 ( .A(in[911]), .B(n8487), .Z(n6454) );
  NOR U2025 ( .A(n6277), .B(n9514), .Z(n6040) );
  XNOR U2026 ( .A(n6454), .B(n6040), .Z(out[1106]) );
  XOR U2027 ( .A(n6042), .B(n6041), .Z(n8491) );
  XNOR U2028 ( .A(in[912]), .B(n8491), .Z(n6456) );
  NOR U2029 ( .A(n6281), .B(n9518), .Z(n6043) );
  XNOR U2030 ( .A(n6456), .B(n6043), .Z(out[1107]) );
  XNOR U2031 ( .A(n6045), .B(n6044), .Z(n8495) );
  XNOR U2032 ( .A(in[913]), .B(n8495), .Z(n6458) );
  NOR U2033 ( .A(n6285), .B(n9526), .Z(n6046) );
  XNOR U2034 ( .A(n6458), .B(n6046), .Z(out[1108]) );
  XOR U2035 ( .A(n6048), .B(n6047), .Z(n8499) );
  XNOR U2036 ( .A(in[914]), .B(n8499), .Z(n6460) );
  NOR U2037 ( .A(n6289), .B(n9530), .Z(n6049) );
  XNOR U2038 ( .A(n6460), .B(n6049), .Z(out[1109]) );
  XOR U2039 ( .A(in[581]), .B(n8443), .Z(n7378) );
  XOR U2040 ( .A(in[236]), .B(n8540), .Z(n7802) );
  XNOR U2041 ( .A(in[1456]), .B(n8581), .Z(n7799) );
  NAND U2042 ( .A(n7802), .B(n7799), .Z(n6050) );
  XNOR U2043 ( .A(n7378), .B(n6050), .Z(out[110]) );
  XOR U2044 ( .A(n6052), .B(n6051), .Z(n8503) );
  XNOR U2045 ( .A(in[915]), .B(n8503), .Z(n6462) );
  NOR U2046 ( .A(n6293), .B(n9534), .Z(n6053) );
  XNOR U2047 ( .A(n6462), .B(n6053), .Z(out[1110]) );
  XNOR U2048 ( .A(n6055), .B(n6054), .Z(n8507) );
  XNOR U2049 ( .A(in[916]), .B(n8507), .Z(n6464) );
  NOR U2050 ( .A(n6297), .B(n9538), .Z(n6056) );
  XNOR U2051 ( .A(n6464), .B(n6056), .Z(out[1111]) );
  XNOR U2052 ( .A(n6058), .B(n6057), .Z(n8511) );
  XNOR U2053 ( .A(in[917]), .B(n8511), .Z(n6467) );
  NOR U2054 ( .A(n6301), .B(n9542), .Z(n6059) );
  XNOR U2055 ( .A(n6467), .B(n6059), .Z(out[1112]) );
  XOR U2056 ( .A(n6061), .B(n6060), .Z(n8519) );
  XNOR U2057 ( .A(in[918]), .B(n8519), .Z(n6469) );
  NOR U2058 ( .A(n6305), .B(n9546), .Z(n6062) );
  XNOR U2059 ( .A(n6469), .B(n6062), .Z(out[1113]) );
  XNOR U2060 ( .A(n6064), .B(n6063), .Z(n8523) );
  XNOR U2061 ( .A(in[919]), .B(n8523), .Z(n6471) );
  NOR U2062 ( .A(n6309), .B(n9550), .Z(n6065) );
  XNOR U2063 ( .A(n6471), .B(n6065), .Z(out[1114]) );
  XNOR U2064 ( .A(n6067), .B(n6066), .Z(n8527) );
  XNOR U2065 ( .A(in[920]), .B(n8527), .Z(n6473) );
  NOR U2066 ( .A(n6313), .B(n9554), .Z(n6068) );
  XNOR U2067 ( .A(n6473), .B(n6068), .Z(out[1115]) );
  XNOR U2068 ( .A(n6070), .B(n6069), .Z(n8531) );
  XNOR U2069 ( .A(in[921]), .B(n8531), .Z(n6475) );
  NOR U2070 ( .A(n6318), .B(n9558), .Z(n6071) );
  XNOR U2071 ( .A(n6475), .B(n6071), .Z(out[1116]) );
  XOR U2072 ( .A(n6073), .B(n6072), .Z(n8535) );
  XNOR U2073 ( .A(in[922]), .B(n8535), .Z(n6477) );
  NOR U2074 ( .A(n6322), .B(n9562), .Z(n6074) );
  XNOR U2075 ( .A(n6477), .B(n6074), .Z(out[1117]) );
  XOR U2076 ( .A(n6076), .B(n6075), .Z(n8539) );
  XNOR U2077 ( .A(in[923]), .B(n8539), .Z(n6479) );
  NOR U2078 ( .A(n6326), .B(n9570), .Z(n6077) );
  XNOR U2079 ( .A(n6479), .B(n6077), .Z(out[1118]) );
  XOR U2080 ( .A(n6079), .B(n6078), .Z(n8543) );
  XNOR U2081 ( .A(in[924]), .B(n8543), .Z(n6481) );
  NOR U2082 ( .A(n6330), .B(n9574), .Z(n6080) );
  XNOR U2083 ( .A(n6481), .B(n6080), .Z(out[1119]) );
  XOR U2084 ( .A(in[582]), .B(n8447), .Z(n7380) );
  XOR U2085 ( .A(in[237]), .B(n8544), .Z(n7826) );
  XNOR U2086 ( .A(in[1457]), .B(n8585), .Z(n7823) );
  NAND U2087 ( .A(n7826), .B(n7823), .Z(n6081) );
  XNOR U2088 ( .A(n7380), .B(n6081), .Z(out[111]) );
  XOR U2089 ( .A(n6083), .B(n6082), .Z(n8547) );
  XNOR U2090 ( .A(in[925]), .B(n8547), .Z(n6483) );
  NOR U2091 ( .A(n6334), .B(n9578), .Z(n6084) );
  XNOR U2092 ( .A(n6483), .B(n6084), .Z(out[1120]) );
  XOR U2093 ( .A(n6086), .B(n6085), .Z(n8551) );
  XNOR U2094 ( .A(in[926]), .B(n8551), .Z(n6485) );
  NOR U2095 ( .A(n6338), .B(n9582), .Z(n6087) );
  XNOR U2096 ( .A(n6485), .B(n6087), .Z(out[1121]) );
  XOR U2097 ( .A(n6089), .B(n6088), .Z(n8555) );
  XNOR U2098 ( .A(in[927]), .B(n8555), .Z(n6488) );
  NOR U2099 ( .A(n6342), .B(n9586), .Z(n6090) );
  XNOR U2100 ( .A(n6488), .B(n6090), .Z(out[1122]) );
  XOR U2101 ( .A(n6092), .B(n6091), .Z(n8563) );
  XNOR U2102 ( .A(in[928]), .B(n8563), .Z(n6490) );
  NOR U2103 ( .A(n6346), .B(n9590), .Z(n6093) );
  XNOR U2104 ( .A(n6490), .B(n6093), .Z(out[1123]) );
  XNOR U2105 ( .A(n6095), .B(n6094), .Z(n8567) );
  XNOR U2106 ( .A(in[929]), .B(n8567), .Z(n6492) );
  NOR U2107 ( .A(n6350), .B(n9594), .Z(n6096) );
  XNOR U2108 ( .A(n6492), .B(n6096), .Z(out[1124]) );
  XNOR U2109 ( .A(n6098), .B(n6097), .Z(n8571) );
  XNOR U2110 ( .A(in[930]), .B(n8571), .Z(n6494) );
  NOR U2111 ( .A(n6354), .B(n9598), .Z(n6099) );
  XNOR U2112 ( .A(n6494), .B(n6099), .Z(out[1125]) );
  XNOR U2113 ( .A(n6101), .B(n6100), .Z(n8575) );
  XNOR U2114 ( .A(in[931]), .B(n8575), .Z(n6496) );
  NOR U2115 ( .A(n6359), .B(n9602), .Z(n6102) );
  XNOR U2116 ( .A(n6496), .B(n6102), .Z(out[1126]) );
  XNOR U2117 ( .A(n6104), .B(n6103), .Z(n8579) );
  XNOR U2118 ( .A(in[932]), .B(n8579), .Z(n6498) );
  NOR U2119 ( .A(n6363), .B(n9606), .Z(n6105) );
  XNOR U2120 ( .A(n6498), .B(n6105), .Z(out[1127]) );
  XNOR U2121 ( .A(n6107), .B(n6106), .Z(n8583) );
  XNOR U2122 ( .A(in[933]), .B(n8583), .Z(n6501) );
  NAND U2123 ( .A(n6365), .B(n6108), .Z(n6109) );
  XNOR U2124 ( .A(n6501), .B(n6109), .Z(out[1128]) );
  XOR U2125 ( .A(n6111), .B(n6110), .Z(n8587) );
  XNOR U2126 ( .A(in[934]), .B(n8587), .Z(n6505) );
  NAND U2127 ( .A(n6367), .B(n6112), .Z(n6113) );
  XNOR U2128 ( .A(n6505), .B(n6113), .Z(out[1129]) );
  XOR U2129 ( .A(in[583]), .B(n8451), .Z(n7383) );
  XOR U2130 ( .A(in[238]), .B(n8548), .Z(n7850) );
  XNOR U2131 ( .A(in[1458]), .B(n8589), .Z(n7847) );
  NAND U2132 ( .A(n7850), .B(n7847), .Z(n6114) );
  XNOR U2133 ( .A(n7383), .B(n6114), .Z(out[112]) );
  XNOR U2134 ( .A(n6116), .B(n6115), .Z(n8591) );
  XNOR U2135 ( .A(in[935]), .B(n8591), .Z(n6509) );
  NAND U2136 ( .A(n6369), .B(n6117), .Z(n6118) );
  XNOR U2137 ( .A(n6509), .B(n6118), .Z(out[1130]) );
  XNOR U2138 ( .A(n6120), .B(n6119), .Z(n8595) );
  XNOR U2139 ( .A(in[936]), .B(n8595), .Z(n6513) );
  NAND U2140 ( .A(n6371), .B(n6121), .Z(n6122) );
  XNOR U2141 ( .A(n6513), .B(n6122), .Z(out[1131]) );
  XNOR U2142 ( .A(n6124), .B(n6123), .Z(n8599) );
  XNOR U2143 ( .A(in[937]), .B(n8599), .Z(n6518) );
  NAND U2144 ( .A(n6373), .B(n6125), .Z(n6126) );
  XNOR U2145 ( .A(n6518), .B(n6126), .Z(out[1132]) );
  XNOR U2146 ( .A(n6128), .B(n6127), .Z(n8609) );
  XNOR U2147 ( .A(in[938]), .B(n8609), .Z(n6522) );
  NAND U2148 ( .A(n6375), .B(n6129), .Z(n6130) );
  XNOR U2149 ( .A(n6522), .B(n6130), .Z(out[1133]) );
  XNOR U2150 ( .A(n6132), .B(n6131), .Z(n8613) );
  XNOR U2151 ( .A(in[939]), .B(n8613), .Z(n6526) );
  NAND U2152 ( .A(n6377), .B(n6133), .Z(n6134) );
  XNOR U2153 ( .A(n6526), .B(n6134), .Z(out[1134]) );
  XNOR U2154 ( .A(n6136), .B(n6135), .Z(n8617) );
  XNOR U2155 ( .A(in[940]), .B(n8617), .Z(n6530) );
  NAND U2156 ( .A(n6379), .B(n6137), .Z(n6138) );
  XNOR U2157 ( .A(n6530), .B(n6138), .Z(out[1135]) );
  XNOR U2158 ( .A(n6140), .B(n6139), .Z(n8621) );
  XNOR U2159 ( .A(in[941]), .B(n8621), .Z(n6534) );
  NAND U2160 ( .A(n6383), .B(n6141), .Z(n6142) );
  XNOR U2161 ( .A(n6534), .B(n6142), .Z(out[1136]) );
  XNOR U2162 ( .A(n6144), .B(n6143), .Z(n8343) );
  XNOR U2163 ( .A(in[942]), .B(n8343), .Z(n6538) );
  NAND U2164 ( .A(n6385), .B(n6145), .Z(n6146) );
  XNOR U2165 ( .A(n6538), .B(n6146), .Z(out[1137]) );
  XNOR U2166 ( .A(n6148), .B(n6147), .Z(n8347) );
  XNOR U2167 ( .A(in[943]), .B(n8347), .Z(n6542) );
  NAND U2168 ( .A(n6387), .B(n6149), .Z(n6150) );
  XNOR U2169 ( .A(n6542), .B(n6150), .Z(out[1138]) );
  XNOR U2170 ( .A(n6152), .B(n6151), .Z(n8351) );
  XNOR U2171 ( .A(in[944]), .B(n8351), .Z(n6546) );
  NAND U2172 ( .A(n6389), .B(n6153), .Z(n6154) );
  XNOR U2173 ( .A(n6546), .B(n6154), .Z(out[1139]) );
  XOR U2174 ( .A(in[584]), .B(n8455), .Z(n7385) );
  XOR U2175 ( .A(in[239]), .B(n8552), .Z(n7874) );
  XNOR U2176 ( .A(in[1459]), .B(n8593), .Z(n7871) );
  NAND U2177 ( .A(n7874), .B(n7871), .Z(n6155) );
  XNOR U2178 ( .A(n7385), .B(n6155), .Z(out[113]) );
  XNOR U2179 ( .A(n6157), .B(n6156), .Z(n8355) );
  XNOR U2180 ( .A(in[945]), .B(n8355), .Z(n6550) );
  NAND U2181 ( .A(n6391), .B(n6158), .Z(n6159) );
  XNOR U2182 ( .A(n6550), .B(n6159), .Z(out[1140]) );
  XNOR U2183 ( .A(n6161), .B(n6160), .Z(n8359) );
  XNOR U2184 ( .A(in[946]), .B(n8359), .Z(n6554) );
  NAND U2185 ( .A(n6393), .B(n6162), .Z(n6163) );
  XNOR U2186 ( .A(n6554), .B(n6163), .Z(out[1141]) );
  XNOR U2187 ( .A(n6165), .B(n6164), .Z(n8363) );
  XNOR U2188 ( .A(in[947]), .B(n8363), .Z(n6559) );
  NAND U2189 ( .A(n6395), .B(n6166), .Z(n6167) );
  XNOR U2190 ( .A(n6559), .B(n6167), .Z(out[1142]) );
  XNOR U2191 ( .A(n6169), .B(n6168), .Z(n8367) );
  XNOR U2192 ( .A(in[948]), .B(n8367), .Z(n6563) );
  NAND U2193 ( .A(n6397), .B(n6170), .Z(n6171) );
  XNOR U2194 ( .A(n6563), .B(n6171), .Z(out[1143]) );
  XNOR U2195 ( .A(n6173), .B(n6172), .Z(n8371) );
  XNOR U2196 ( .A(in[949]), .B(n8371), .Z(n6567) );
  NAND U2197 ( .A(n6399), .B(n6174), .Z(n6175) );
  XNOR U2198 ( .A(n6567), .B(n6175), .Z(out[1144]) );
  XNOR U2199 ( .A(n6177), .B(n6176), .Z(n8375) );
  XNOR U2200 ( .A(in[950]), .B(n8375), .Z(n6571) );
  NAND U2201 ( .A(n6401), .B(n6178), .Z(n6179) );
  XNOR U2202 ( .A(n6571), .B(n6179), .Z(out[1145]) );
  XNOR U2203 ( .A(n6181), .B(n6180), .Z(n8379) );
  XNOR U2204 ( .A(in[951]), .B(n8379), .Z(n6575) );
  NAND U2205 ( .A(n6404), .B(n6182), .Z(n6183) );
  XNOR U2206 ( .A(n6575), .B(n6183), .Z(out[1146]) );
  XNOR U2207 ( .A(n6185), .B(n6184), .Z(n8387) );
  XNOR U2208 ( .A(in[952]), .B(n8387), .Z(n6579) );
  NAND U2209 ( .A(n6406), .B(n6186), .Z(n6187) );
  XNOR U2210 ( .A(n6579), .B(n6187), .Z(out[1147]) );
  XNOR U2211 ( .A(n6189), .B(n6188), .Z(n8391) );
  XNOR U2212 ( .A(in[953]), .B(n8391), .Z(n6583) );
  NAND U2213 ( .A(n6408), .B(n6190), .Z(n6191) );
  XNOR U2214 ( .A(n6583), .B(n6191), .Z(out[1148]) );
  XNOR U2215 ( .A(n6193), .B(n6192), .Z(n8395) );
  XNOR U2216 ( .A(in[954]), .B(n8395), .Z(n6587) );
  NAND U2217 ( .A(n6410), .B(n6194), .Z(n6195) );
  XNOR U2218 ( .A(n6587), .B(n6195), .Z(out[1149]) );
  XOR U2219 ( .A(in[585]), .B(n8459), .Z(n7387) );
  XOR U2220 ( .A(in[240]), .B(n8556), .Z(n7900) );
  XNOR U2221 ( .A(in[1460]), .B(n8597), .Z(n7897) );
  NAND U2222 ( .A(n7900), .B(n7897), .Z(n6196) );
  XNOR U2223 ( .A(n7387), .B(n6196), .Z(out[114]) );
  XNOR U2224 ( .A(in[955]), .B(n8399), .Z(n6591) );
  NAND U2225 ( .A(n6412), .B(n6197), .Z(n6198) );
  XNOR U2226 ( .A(n6591), .B(n6198), .Z(out[1150]) );
  XNOR U2227 ( .A(in[956]), .B(n8403), .Z(n6595) );
  NAND U2228 ( .A(n6414), .B(n6199), .Z(n6200) );
  XNOR U2229 ( .A(n6595), .B(n6200), .Z(out[1151]) );
  XNOR U2230 ( .A(n6202), .B(n6201), .Z(n8743) );
  XNOR U2231 ( .A(in[1004]), .B(n8743), .Z(n9436) );
  NAND U2232 ( .A(n6416), .B(n6203), .Z(n6204) );
  XNOR U2233 ( .A(n9436), .B(n6204), .Z(out[1152]) );
  XNOR U2234 ( .A(n6206), .B(n6205), .Z(n8745) );
  XNOR U2235 ( .A(in[1005]), .B(n8745), .Z(n9440) );
  NAND U2236 ( .A(n6418), .B(n6207), .Z(n6208) );
  XNOR U2237 ( .A(n9440), .B(n6208), .Z(out[1153]) );
  XNOR U2238 ( .A(n6210), .B(n6209), .Z(n8747) );
  XNOR U2239 ( .A(in[1006]), .B(n8747), .Z(n9444) );
  NAND U2240 ( .A(n6420), .B(n6211), .Z(n6212) );
  XNOR U2241 ( .A(n9444), .B(n6212), .Z(out[1154]) );
  XNOR U2242 ( .A(n6214), .B(n6213), .Z(n8749) );
  XNOR U2243 ( .A(in[1007]), .B(n8749), .Z(n9448) );
  NAND U2244 ( .A(n6422), .B(n6215), .Z(n6216) );
  XNOR U2245 ( .A(n9448), .B(n6216), .Z(out[1155]) );
  XNOR U2246 ( .A(n6218), .B(n6217), .Z(n8755) );
  XNOR U2247 ( .A(in[1008]), .B(n8755), .Z(n9452) );
  NAND U2248 ( .A(n6425), .B(n6219), .Z(n6220) );
  XNOR U2249 ( .A(n9452), .B(n6220), .Z(out[1156]) );
  XNOR U2250 ( .A(n6222), .B(n6221), .Z(n8757) );
  XNOR U2251 ( .A(in[1009]), .B(n8757), .Z(n9456) );
  NAND U2252 ( .A(n6427), .B(n6223), .Z(n6224) );
  XNOR U2253 ( .A(n9456), .B(n6224), .Z(out[1157]) );
  XNOR U2254 ( .A(n6226), .B(n6225), .Z(n8759) );
  XNOR U2255 ( .A(in[1010]), .B(n8759), .Z(n9460) );
  NAND U2256 ( .A(n6429), .B(n6227), .Z(n6228) );
  XNOR U2257 ( .A(n9460), .B(n6228), .Z(out[1158]) );
  XNOR U2258 ( .A(n6230), .B(n6229), .Z(n8761) );
  XNOR U2259 ( .A(in[1011]), .B(n8761), .Z(n9464) );
  NAND U2260 ( .A(n6431), .B(n6231), .Z(n6232) );
  XNOR U2261 ( .A(n9464), .B(n6232), .Z(out[1159]) );
  XOR U2262 ( .A(in[586]), .B(n8463), .Z(n7389) );
  XOR U2263 ( .A(in[241]), .B(n8564), .Z(n7924) );
  XNOR U2264 ( .A(in[1461]), .B(n8601), .Z(n7921) );
  NAND U2265 ( .A(n7924), .B(n7921), .Z(n6233) );
  XNOR U2266 ( .A(n7389), .B(n6233), .Z(out[115]) );
  XNOR U2267 ( .A(n6235), .B(n6234), .Z(n8763) );
  XNOR U2268 ( .A(in[1012]), .B(n8763), .Z(n9468) );
  NAND U2269 ( .A(n6433), .B(n6236), .Z(n6237) );
  XNOR U2270 ( .A(n9468), .B(n6237), .Z(out[1160]) );
  XNOR U2271 ( .A(n6239), .B(n6238), .Z(n8765) );
  XNOR U2272 ( .A(in[1013]), .B(n8765), .Z(n9472) );
  NAND U2273 ( .A(n6435), .B(n6240), .Z(n6241) );
  XNOR U2274 ( .A(n9472), .B(n6241), .Z(out[1161]) );
  XNOR U2275 ( .A(n6243), .B(n6242), .Z(n8767) );
  XNOR U2276 ( .A(in[1014]), .B(n8767), .Z(n9480) );
  NAND U2277 ( .A(n6437), .B(n6244), .Z(n6245) );
  XNOR U2278 ( .A(n9480), .B(n6245), .Z(out[1162]) );
  XNOR U2279 ( .A(n6247), .B(n6246), .Z(n8769) );
  XNOR U2280 ( .A(in[1015]), .B(n8769), .Z(n9484) );
  NAND U2281 ( .A(n6439), .B(n6248), .Z(n6249) );
  XNOR U2282 ( .A(n9484), .B(n6249), .Z(out[1163]) );
  XNOR U2283 ( .A(n6251), .B(n6250), .Z(n8625) );
  XNOR U2284 ( .A(in[1016]), .B(n8625), .Z(n9488) );
  NAND U2285 ( .A(n6441), .B(n6252), .Z(n6253) );
  XNOR U2286 ( .A(n9488), .B(n6253), .Z(out[1164]) );
  XNOR U2287 ( .A(n6255), .B(n6254), .Z(n8627) );
  XNOR U2288 ( .A(in[1017]), .B(n8627), .Z(n9492) );
  NAND U2289 ( .A(n6443), .B(n6256), .Z(n6257) );
  XNOR U2290 ( .A(n9492), .B(n6257), .Z(out[1165]) );
  XNOR U2291 ( .A(n6259), .B(n6258), .Z(n8629) );
  XNOR U2292 ( .A(in[1018]), .B(n8629), .Z(n9496) );
  NAND U2293 ( .A(n6446), .B(n6260), .Z(n6261) );
  XNOR U2294 ( .A(n9496), .B(n6261), .Z(out[1166]) );
  XNOR U2295 ( .A(n6263), .B(n6262), .Z(n8631) );
  XNOR U2296 ( .A(in[1019]), .B(n8631), .Z(n9500) );
  NAND U2297 ( .A(n6448), .B(n6264), .Z(n6265) );
  XNOR U2298 ( .A(n9500), .B(n6265), .Z(out[1167]) );
  XOR U2299 ( .A(n6267), .B(n6266), .Z(n8633) );
  XNOR U2300 ( .A(in[1020]), .B(n8633), .Z(n9504) );
  NAND U2301 ( .A(n6450), .B(n6268), .Z(n6269) );
  XNOR U2302 ( .A(n9504), .B(n6269), .Z(out[1168]) );
  XOR U2303 ( .A(n6271), .B(n6270), .Z(n8635) );
  XNOR U2304 ( .A(in[1021]), .B(n8635), .Z(n9508) );
  NAND U2305 ( .A(n6452), .B(n6272), .Z(n6273) );
  XNOR U2306 ( .A(n9508), .B(n6273), .Z(out[1169]) );
  XOR U2307 ( .A(in[587]), .B(n8467), .Z(n7391) );
  XOR U2308 ( .A(in[242]), .B(n8568), .Z(n7948) );
  XNOR U2309 ( .A(in[1462]), .B(n8611), .Z(n7945) );
  NAND U2310 ( .A(n7948), .B(n7945), .Z(n6274) );
  XNOR U2311 ( .A(n7391), .B(n6274), .Z(out[116]) );
  XOR U2312 ( .A(n6276), .B(n6275), .Z(n8641) );
  XNOR U2313 ( .A(in[1022]), .B(n8641), .Z(n9512) );
  NAND U2314 ( .A(n6454), .B(n6277), .Z(n6278) );
  XNOR U2315 ( .A(n9512), .B(n6278), .Z(out[1170]) );
  XNOR U2316 ( .A(n6280), .B(n6279), .Z(n8643) );
  XNOR U2317 ( .A(in[1023]), .B(n8643), .Z(n9516) );
  NAND U2318 ( .A(n6456), .B(n6281), .Z(n6282) );
  XNOR U2319 ( .A(n9516), .B(n6282), .Z(out[1171]) );
  XOR U2320 ( .A(n6284), .B(n6283), .Z(n8645) );
  XNOR U2321 ( .A(in[960]), .B(n8645), .Z(n9524) );
  NAND U2322 ( .A(n6458), .B(n6285), .Z(n6286) );
  XNOR U2323 ( .A(n9524), .B(n6286), .Z(out[1172]) );
  XOR U2324 ( .A(n6288), .B(n6287), .Z(n8647) );
  XNOR U2325 ( .A(in[961]), .B(n8647), .Z(n9528) );
  NAND U2326 ( .A(n6460), .B(n6289), .Z(n6290) );
  XNOR U2327 ( .A(n9528), .B(n6290), .Z(out[1173]) );
  XOR U2328 ( .A(n6292), .B(n6291), .Z(n8649) );
  XNOR U2329 ( .A(in[962]), .B(n8649), .Z(n9532) );
  NAND U2330 ( .A(n6462), .B(n6293), .Z(n6294) );
  XNOR U2331 ( .A(n9532), .B(n6294), .Z(out[1174]) );
  XOR U2332 ( .A(n6296), .B(n6295), .Z(n8651) );
  XNOR U2333 ( .A(in[963]), .B(n8651), .Z(n9536) );
  NAND U2334 ( .A(n6464), .B(n6297), .Z(n6298) );
  XNOR U2335 ( .A(n9536), .B(n6298), .Z(out[1175]) );
  XOR U2336 ( .A(n6300), .B(n6299), .Z(n8653) );
  XNOR U2337 ( .A(in[964]), .B(n8653), .Z(n9540) );
  NAND U2338 ( .A(n6467), .B(n6301), .Z(n6302) );
  XNOR U2339 ( .A(n9540), .B(n6302), .Z(out[1176]) );
  XOR U2340 ( .A(n6304), .B(n6303), .Z(n8655) );
  XNOR U2341 ( .A(in[965]), .B(n8655), .Z(n9544) );
  NAND U2342 ( .A(n6469), .B(n6305), .Z(n6306) );
  XNOR U2343 ( .A(n9544), .B(n6306), .Z(out[1177]) );
  XOR U2344 ( .A(n6308), .B(n6307), .Z(n8657) );
  XNOR U2345 ( .A(in[966]), .B(n8657), .Z(n9548) );
  NAND U2346 ( .A(n6471), .B(n6309), .Z(n6310) );
  XNOR U2347 ( .A(n9548), .B(n6310), .Z(out[1178]) );
  XOR U2348 ( .A(n6312), .B(n6311), .Z(n8659) );
  XNOR U2349 ( .A(in[967]), .B(n8659), .Z(n9552) );
  NAND U2350 ( .A(n6473), .B(n6313), .Z(n6314) );
  XNOR U2351 ( .A(n9552), .B(n6314), .Z(out[1179]) );
  XOR U2352 ( .A(in[588]), .B(n8475), .Z(n7393) );
  XOR U2353 ( .A(in[243]), .B(n8572), .Z(n7972) );
  XNOR U2354 ( .A(in[1463]), .B(n8615), .Z(n7969) );
  NAND U2355 ( .A(n7972), .B(n7969), .Z(n6315) );
  XNOR U2356 ( .A(n7393), .B(n6315), .Z(out[117]) );
  XOR U2357 ( .A(n6317), .B(n6316), .Z(n8663) );
  XNOR U2358 ( .A(in[968]), .B(n8663), .Z(n9556) );
  NAND U2359 ( .A(n6475), .B(n6318), .Z(n6319) );
  XNOR U2360 ( .A(n9556), .B(n6319), .Z(out[1180]) );
  XOR U2361 ( .A(n6321), .B(n6320), .Z(n8665) );
  XNOR U2362 ( .A(in[969]), .B(n8665), .Z(n9560) );
  NAND U2363 ( .A(n6477), .B(n6322), .Z(n6323) );
  XNOR U2364 ( .A(n9560), .B(n6323), .Z(out[1181]) );
  XNOR U2365 ( .A(n6325), .B(n6324), .Z(n8667) );
  XNOR U2366 ( .A(in[970]), .B(n8667), .Z(n9568) );
  NAND U2367 ( .A(n6479), .B(n6326), .Z(n6327) );
  XNOR U2368 ( .A(n9568), .B(n6327), .Z(out[1182]) );
  XOR U2369 ( .A(n6329), .B(n6328), .Z(n8669) );
  XNOR U2370 ( .A(in[971]), .B(n8669), .Z(n9572) );
  NAND U2371 ( .A(n6481), .B(n6330), .Z(n6331) );
  XNOR U2372 ( .A(n9572), .B(n6331), .Z(out[1183]) );
  XOR U2373 ( .A(n6333), .B(n6332), .Z(n8671) );
  XNOR U2374 ( .A(in[972]), .B(n8671), .Z(n9576) );
  NAND U2375 ( .A(n6483), .B(n6334), .Z(n6335) );
  XNOR U2376 ( .A(n9576), .B(n6335), .Z(out[1184]) );
  XOR U2377 ( .A(n6337), .B(n6336), .Z(n8673) );
  XNOR U2378 ( .A(in[973]), .B(n8673), .Z(n9580) );
  NAND U2379 ( .A(n6485), .B(n6338), .Z(n6339) );
  XNOR U2380 ( .A(n9580), .B(n6339), .Z(out[1185]) );
  XNOR U2381 ( .A(n6341), .B(n6340), .Z(n8675) );
  XNOR U2382 ( .A(in[974]), .B(n8675), .Z(n9584) );
  NAND U2383 ( .A(n6488), .B(n6342), .Z(n6343) );
  XNOR U2384 ( .A(n9584), .B(n6343), .Z(out[1186]) );
  XNOR U2385 ( .A(n6345), .B(n6344), .Z(n8677) );
  XNOR U2386 ( .A(in[975]), .B(n8677), .Z(n9588) );
  NAND U2387 ( .A(n6490), .B(n6346), .Z(n6347) );
  XNOR U2388 ( .A(n9588), .B(n6347), .Z(out[1187]) );
  XNOR U2389 ( .A(n6349), .B(n6348), .Z(n8679) );
  XNOR U2390 ( .A(in[976]), .B(n8679), .Z(n9592) );
  NAND U2391 ( .A(n6492), .B(n6350), .Z(n6351) );
  XNOR U2392 ( .A(n9592), .B(n6351), .Z(out[1188]) );
  XOR U2393 ( .A(n6353), .B(n6352), .Z(n8681) );
  XNOR U2394 ( .A(in[977]), .B(n8681), .Z(n9596) );
  NAND U2395 ( .A(n6494), .B(n6354), .Z(n6355) );
  XNOR U2396 ( .A(n9596), .B(n6355), .Z(out[1189]) );
  XOR U2397 ( .A(in[589]), .B(n8479), .Z(n7395) );
  XOR U2398 ( .A(in[244]), .B(n8576), .Z(n7996) );
  XNOR U2399 ( .A(in[1464]), .B(n8619), .Z(n7993) );
  NAND U2400 ( .A(n7996), .B(n7993), .Z(n6356) );
  XNOR U2401 ( .A(n7395), .B(n6356), .Z(out[118]) );
  XOR U2402 ( .A(n6358), .B(n6357), .Z(n8685) );
  XNOR U2403 ( .A(in[978]), .B(n8685), .Z(n9600) );
  NAND U2404 ( .A(n6496), .B(n6359), .Z(n6360) );
  XNOR U2405 ( .A(n9600), .B(n6360), .Z(out[1190]) );
  XOR U2406 ( .A(n6362), .B(n6361), .Z(n8687) );
  XNOR U2407 ( .A(in[979]), .B(n8687), .Z(n9604) );
  NAND U2408 ( .A(n6498), .B(n6363), .Z(n6364) );
  XNOR U2409 ( .A(n9604), .B(n6364), .Z(out[1191]) );
  OR U2410 ( .A(n6501), .B(n6365), .Z(n6366) );
  XNOR U2411 ( .A(n6500), .B(n6366), .Z(out[1192]) );
  OR U2412 ( .A(n6505), .B(n6367), .Z(n6368) );
  XNOR U2413 ( .A(n6504), .B(n6368), .Z(out[1193]) );
  OR U2414 ( .A(n6509), .B(n6369), .Z(n6370) );
  XNOR U2415 ( .A(n6508), .B(n6370), .Z(out[1194]) );
  OR U2416 ( .A(n6513), .B(n6371), .Z(n6372) );
  XNOR U2417 ( .A(n6512), .B(n6372), .Z(out[1195]) );
  OR U2418 ( .A(n6518), .B(n6373), .Z(n6374) );
  XNOR U2419 ( .A(n6517), .B(n6374), .Z(out[1196]) );
  OR U2420 ( .A(n6522), .B(n6375), .Z(n6376) );
  XNOR U2421 ( .A(n6521), .B(n6376), .Z(out[1197]) );
  OR U2422 ( .A(n6526), .B(n6377), .Z(n6378) );
  XNOR U2423 ( .A(n6525), .B(n6378), .Z(out[1198]) );
  OR U2424 ( .A(n6530), .B(n6379), .Z(n6380) );
  XNOR U2425 ( .A(n6529), .B(n6380), .Z(out[1199]) );
  XOR U2426 ( .A(in[590]), .B(n8483), .Z(n7397) );
  XOR U2427 ( .A(in[245]), .B(n8580), .Z(n8020) );
  XNOR U2428 ( .A(in[1465]), .B(n8623), .Z(n8017) );
  NAND U2429 ( .A(n8020), .B(n8017), .Z(n6381) );
  XNOR U2430 ( .A(n7397), .B(n6381), .Z(out[119]) );
  XOR U2431 ( .A(in[201]), .B(n8388), .Z(n8752) );
  XNOR U2432 ( .A(in[1421]), .B(n8425), .Z(n8751) );
  XOR U2433 ( .A(in[1044]), .B(n8930), .Z(n7442) );
  NAND U2434 ( .A(n8751), .B(n7442), .Z(n6382) );
  XNOR U2435 ( .A(n8752), .B(n6382), .Z(out[11]) );
  OR U2436 ( .A(n6534), .B(n6383), .Z(n6384) );
  XNOR U2437 ( .A(n6533), .B(n6384), .Z(out[1200]) );
  OR U2438 ( .A(n6538), .B(n6385), .Z(n6386) );
  XNOR U2439 ( .A(n6537), .B(n6386), .Z(out[1201]) );
  OR U2440 ( .A(n6542), .B(n6387), .Z(n6388) );
  XNOR U2441 ( .A(n6541), .B(n6388), .Z(out[1202]) );
  OR U2442 ( .A(n6546), .B(n6389), .Z(n6390) );
  XNOR U2443 ( .A(n6545), .B(n6390), .Z(out[1203]) );
  OR U2444 ( .A(n6550), .B(n6391), .Z(n6392) );
  XNOR U2445 ( .A(n6549), .B(n6392), .Z(out[1204]) );
  OR U2446 ( .A(n6554), .B(n6393), .Z(n6394) );
  XNOR U2447 ( .A(n6553), .B(n6394), .Z(out[1205]) );
  OR U2448 ( .A(n6559), .B(n6395), .Z(n6396) );
  XNOR U2449 ( .A(n6558), .B(n6396), .Z(out[1206]) );
  OR U2450 ( .A(n6563), .B(n6397), .Z(n6398) );
  XNOR U2451 ( .A(n6562), .B(n6398), .Z(out[1207]) );
  OR U2452 ( .A(n6567), .B(n6399), .Z(n6400) );
  XNOR U2453 ( .A(n6566), .B(n6400), .Z(out[1208]) );
  OR U2454 ( .A(n6571), .B(n6401), .Z(n6402) );
  XNOR U2455 ( .A(n6570), .B(n6402), .Z(out[1209]) );
  XOR U2456 ( .A(in[591]), .B(n8487), .Z(n7399) );
  XOR U2457 ( .A(in[246]), .B(n8584), .Z(n8044) );
  XNOR U2458 ( .A(in[1466]), .B(n8345), .Z(n8041) );
  NAND U2459 ( .A(n8044), .B(n8041), .Z(n6403) );
  XNOR U2460 ( .A(n7399), .B(n6403), .Z(out[120]) );
  OR U2461 ( .A(n6575), .B(n6404), .Z(n6405) );
  XNOR U2462 ( .A(n6574), .B(n6405), .Z(out[1210]) );
  OR U2463 ( .A(n6579), .B(n6406), .Z(n6407) );
  XNOR U2464 ( .A(n6578), .B(n6407), .Z(out[1211]) );
  OR U2465 ( .A(n6583), .B(n6408), .Z(n6409) );
  XNOR U2466 ( .A(n6582), .B(n6409), .Z(out[1212]) );
  OR U2467 ( .A(n6587), .B(n6410), .Z(n6411) );
  XNOR U2468 ( .A(n6586), .B(n6411), .Z(out[1213]) );
  OR U2469 ( .A(n6591), .B(n6412), .Z(n6413) );
  XNOR U2470 ( .A(n6590), .B(n6413), .Z(out[1214]) );
  OR U2471 ( .A(n6595), .B(n6414), .Z(n6415) );
  XNOR U2472 ( .A(n6594), .B(n6415), .Z(out[1215]) );
  OR U2473 ( .A(n9436), .B(n6416), .Z(n6417) );
  XNOR U2474 ( .A(n9435), .B(n6417), .Z(out[1216]) );
  OR U2475 ( .A(n9440), .B(n6418), .Z(n6419) );
  XNOR U2476 ( .A(n9439), .B(n6419), .Z(out[1217]) );
  OR U2477 ( .A(n9444), .B(n6420), .Z(n6421) );
  XNOR U2478 ( .A(n9443), .B(n6421), .Z(out[1218]) );
  OR U2479 ( .A(n9448), .B(n6422), .Z(n6423) );
  XNOR U2480 ( .A(n9447), .B(n6423), .Z(out[1219]) );
  XOR U2481 ( .A(in[592]), .B(n8491), .Z(n7401) );
  XOR U2482 ( .A(in[247]), .B(n8588), .Z(n8076) );
  XNOR U2483 ( .A(in[1467]), .B(n8349), .Z(n8073) );
  NAND U2484 ( .A(n8076), .B(n8073), .Z(n6424) );
  XNOR U2485 ( .A(n7401), .B(n6424), .Z(out[121]) );
  OR U2486 ( .A(n9452), .B(n6425), .Z(n6426) );
  XNOR U2487 ( .A(n9451), .B(n6426), .Z(out[1220]) );
  OR U2488 ( .A(n9456), .B(n6427), .Z(n6428) );
  XNOR U2489 ( .A(n9455), .B(n6428), .Z(out[1221]) );
  OR U2490 ( .A(n9460), .B(n6429), .Z(n6430) );
  XNOR U2491 ( .A(n9459), .B(n6430), .Z(out[1222]) );
  OR U2492 ( .A(n9464), .B(n6431), .Z(n6432) );
  XNOR U2493 ( .A(n9463), .B(n6432), .Z(out[1223]) );
  OR U2494 ( .A(n9468), .B(n6433), .Z(n6434) );
  XNOR U2495 ( .A(n9467), .B(n6434), .Z(out[1224]) );
  OR U2496 ( .A(n9472), .B(n6435), .Z(n6436) );
  XNOR U2497 ( .A(n9471), .B(n6436), .Z(out[1225]) );
  OR U2498 ( .A(n9480), .B(n6437), .Z(n6438) );
  XNOR U2499 ( .A(n9479), .B(n6438), .Z(out[1226]) );
  OR U2500 ( .A(n9484), .B(n6439), .Z(n6440) );
  XNOR U2501 ( .A(n9483), .B(n6440), .Z(out[1227]) );
  OR U2502 ( .A(n9488), .B(n6441), .Z(n6442) );
  XNOR U2503 ( .A(n9487), .B(n6442), .Z(out[1228]) );
  OR U2504 ( .A(n9492), .B(n6443), .Z(n6444) );
  XNOR U2505 ( .A(n9491), .B(n6444), .Z(out[1229]) );
  XOR U2506 ( .A(in[593]), .B(n8495), .Z(n7404) );
  XOR U2507 ( .A(in[248]), .B(n8592), .Z(n8120) );
  XNOR U2508 ( .A(in[1468]), .B(n8353), .Z(n8117) );
  NAND U2509 ( .A(n8120), .B(n8117), .Z(n6445) );
  XNOR U2510 ( .A(n7404), .B(n6445), .Z(out[122]) );
  OR U2511 ( .A(n9496), .B(n6446), .Z(n6447) );
  XNOR U2512 ( .A(n9495), .B(n6447), .Z(out[1230]) );
  OR U2513 ( .A(n9500), .B(n6448), .Z(n6449) );
  XNOR U2514 ( .A(n9499), .B(n6449), .Z(out[1231]) );
  OR U2515 ( .A(n9504), .B(n6450), .Z(n6451) );
  XNOR U2516 ( .A(n9503), .B(n6451), .Z(out[1232]) );
  OR U2517 ( .A(n9508), .B(n6452), .Z(n6453) );
  XNOR U2518 ( .A(n9507), .B(n6453), .Z(out[1233]) );
  OR U2519 ( .A(n9512), .B(n6454), .Z(n6455) );
  XNOR U2520 ( .A(n9511), .B(n6455), .Z(out[1234]) );
  OR U2521 ( .A(n9516), .B(n6456), .Z(n6457) );
  XNOR U2522 ( .A(n9515), .B(n6457), .Z(out[1235]) );
  OR U2523 ( .A(n9524), .B(n6458), .Z(n6459) );
  XNOR U2524 ( .A(n9523), .B(n6459), .Z(out[1236]) );
  OR U2525 ( .A(n9528), .B(n6460), .Z(n6461) );
  XNOR U2526 ( .A(n9527), .B(n6461), .Z(out[1237]) );
  OR U2527 ( .A(n9532), .B(n6462), .Z(n6463) );
  XNOR U2528 ( .A(n9531), .B(n6463), .Z(out[1238]) );
  OR U2529 ( .A(n9536), .B(n6464), .Z(n6465) );
  XNOR U2530 ( .A(n9535), .B(n6465), .Z(out[1239]) );
  XOR U2531 ( .A(in[594]), .B(n8499), .Z(n7406) );
  XOR U2532 ( .A(in[249]), .B(n8596), .Z(n8164) );
  XNOR U2533 ( .A(in[1469]), .B(n8357), .Z(n8161) );
  NAND U2534 ( .A(n8164), .B(n8161), .Z(n6466) );
  XNOR U2535 ( .A(n7406), .B(n6466), .Z(out[123]) );
  OR U2536 ( .A(n9540), .B(n6467), .Z(n6468) );
  XNOR U2537 ( .A(n9539), .B(n6468), .Z(out[1240]) );
  OR U2538 ( .A(n9544), .B(n6469), .Z(n6470) );
  XNOR U2539 ( .A(n9543), .B(n6470), .Z(out[1241]) );
  OR U2540 ( .A(n9548), .B(n6471), .Z(n6472) );
  XNOR U2541 ( .A(n9547), .B(n6472), .Z(out[1242]) );
  OR U2542 ( .A(n9552), .B(n6473), .Z(n6474) );
  XNOR U2543 ( .A(n9551), .B(n6474), .Z(out[1243]) );
  OR U2544 ( .A(n9556), .B(n6475), .Z(n6476) );
  XNOR U2545 ( .A(n9555), .B(n6476), .Z(out[1244]) );
  OR U2546 ( .A(n9560), .B(n6477), .Z(n6478) );
  XNOR U2547 ( .A(n9559), .B(n6478), .Z(out[1245]) );
  OR U2548 ( .A(n9568), .B(n6479), .Z(n6480) );
  XNOR U2549 ( .A(n9567), .B(n6480), .Z(out[1246]) );
  OR U2550 ( .A(n9572), .B(n6481), .Z(n6482) );
  XNOR U2551 ( .A(n9571), .B(n6482), .Z(out[1247]) );
  OR U2552 ( .A(n9576), .B(n6483), .Z(n6484) );
  XNOR U2553 ( .A(n9575), .B(n6484), .Z(out[1248]) );
  OR U2554 ( .A(n9580), .B(n6485), .Z(n6486) );
  XNOR U2555 ( .A(n9579), .B(n6486), .Z(out[1249]) );
  XOR U2556 ( .A(in[595]), .B(n8503), .Z(n7408) );
  XOR U2557 ( .A(in[250]), .B(n8600), .Z(n8210) );
  XNOR U2558 ( .A(in[1470]), .B(n8361), .Z(n8207) );
  NAND U2559 ( .A(n8210), .B(n8207), .Z(n6487) );
  XNOR U2560 ( .A(n7408), .B(n6487), .Z(out[124]) );
  OR U2561 ( .A(n9584), .B(n6488), .Z(n6489) );
  XNOR U2562 ( .A(n9583), .B(n6489), .Z(out[1250]) );
  OR U2563 ( .A(n9588), .B(n6490), .Z(n6491) );
  XNOR U2564 ( .A(n9587), .B(n6491), .Z(out[1251]) );
  OR U2565 ( .A(n9592), .B(n6492), .Z(n6493) );
  XNOR U2566 ( .A(n9591), .B(n6493), .Z(out[1252]) );
  OR U2567 ( .A(n9596), .B(n6494), .Z(n6495) );
  XNOR U2568 ( .A(n9595), .B(n6495), .Z(out[1253]) );
  OR U2569 ( .A(n9600), .B(n6496), .Z(n6497) );
  XNOR U2570 ( .A(n9599), .B(n6497), .Z(out[1254]) );
  OR U2571 ( .A(n9604), .B(n6498), .Z(n6499) );
  XNOR U2572 ( .A(n9603), .B(n6499), .Z(out[1255]) );
  ANDN U2573 ( .B(n6501), .A(n6500), .Z(n6502) );
  XNOR U2574 ( .A(n6503), .B(n6502), .Z(out[1256]) );
  ANDN U2575 ( .B(n6505), .A(n6504), .Z(n6506) );
  XNOR U2576 ( .A(n6507), .B(n6506), .Z(out[1257]) );
  ANDN U2577 ( .B(n6509), .A(n6508), .Z(n6510) );
  XNOR U2578 ( .A(n6511), .B(n6510), .Z(out[1258]) );
  ANDN U2579 ( .B(n6513), .A(n6512), .Z(n6514) );
  XNOR U2580 ( .A(n6515), .B(n6514), .Z(out[1259]) );
  XOR U2581 ( .A(in[596]), .B(n8507), .Z(n7410) );
  XNOR U2582 ( .A(in[251]), .B(n8610), .Z(n8254) );
  XNOR U2583 ( .A(in[1471]), .B(n8365), .Z(n8251) );
  NAND U2584 ( .A(n8254), .B(n8251), .Z(n6516) );
  XNOR U2585 ( .A(n7410), .B(n6516), .Z(out[125]) );
  ANDN U2586 ( .B(n6518), .A(n6517), .Z(n6519) );
  XNOR U2587 ( .A(n6520), .B(n6519), .Z(out[1260]) );
  ANDN U2588 ( .B(n6522), .A(n6521), .Z(n6523) );
  XNOR U2589 ( .A(n6524), .B(n6523), .Z(out[1261]) );
  ANDN U2590 ( .B(n6526), .A(n6525), .Z(n6527) );
  XNOR U2591 ( .A(n6528), .B(n6527), .Z(out[1262]) );
  ANDN U2592 ( .B(n6530), .A(n6529), .Z(n6531) );
  XNOR U2593 ( .A(n6532), .B(n6531), .Z(out[1263]) );
  ANDN U2594 ( .B(n6534), .A(n6533), .Z(n6535) );
  XNOR U2595 ( .A(n6536), .B(n6535), .Z(out[1264]) );
  ANDN U2596 ( .B(n6538), .A(n6537), .Z(n6539) );
  XNOR U2597 ( .A(n6540), .B(n6539), .Z(out[1265]) );
  ANDN U2598 ( .B(n6542), .A(n6541), .Z(n6543) );
  XNOR U2599 ( .A(n6544), .B(n6543), .Z(out[1266]) );
  ANDN U2600 ( .B(n6546), .A(n6545), .Z(n6547) );
  XNOR U2601 ( .A(n6548), .B(n6547), .Z(out[1267]) );
  ANDN U2602 ( .B(n6550), .A(n6549), .Z(n6551) );
  XNOR U2603 ( .A(n6552), .B(n6551), .Z(out[1268]) );
  ANDN U2604 ( .B(n6554), .A(n6553), .Z(n6555) );
  XNOR U2605 ( .A(n6556), .B(n6555), .Z(out[1269]) );
  XOR U2606 ( .A(in[597]), .B(n8511), .Z(n7412) );
  XNOR U2607 ( .A(in[252]), .B(n8614), .Z(n8298) );
  XNOR U2608 ( .A(in[1408]), .B(n8369), .Z(n8295) );
  NAND U2609 ( .A(n8298), .B(n8295), .Z(n6557) );
  XNOR U2610 ( .A(n7412), .B(n6557), .Z(out[126]) );
  ANDN U2611 ( .B(n6559), .A(n6558), .Z(n6560) );
  XNOR U2612 ( .A(n6561), .B(n6560), .Z(out[1270]) );
  ANDN U2613 ( .B(n6563), .A(n6562), .Z(n6564) );
  XNOR U2614 ( .A(n6565), .B(n6564), .Z(out[1271]) );
  ANDN U2615 ( .B(n6567), .A(n6566), .Z(n6568) );
  XNOR U2616 ( .A(n6569), .B(n6568), .Z(out[1272]) );
  ANDN U2617 ( .B(n6571), .A(n6570), .Z(n6572) );
  XNOR U2618 ( .A(n6573), .B(n6572), .Z(out[1273]) );
  ANDN U2619 ( .B(n6575), .A(n6574), .Z(n6576) );
  XNOR U2620 ( .A(n6577), .B(n6576), .Z(out[1274]) );
  ANDN U2621 ( .B(n6579), .A(n6578), .Z(n6580) );
  XNOR U2622 ( .A(n6581), .B(n6580), .Z(out[1275]) );
  ANDN U2623 ( .B(n6583), .A(n6582), .Z(n6584) );
  XNOR U2624 ( .A(n6585), .B(n6584), .Z(out[1276]) );
  ANDN U2625 ( .B(n6587), .A(n6586), .Z(n6588) );
  XNOR U2626 ( .A(n6589), .B(n6588), .Z(out[1277]) );
  ANDN U2627 ( .B(n6591), .A(n6590), .Z(n6592) );
  XNOR U2628 ( .A(n6593), .B(n6592), .Z(out[1278]) );
  ANDN U2629 ( .B(n6595), .A(n6594), .Z(n6596) );
  XNOR U2630 ( .A(n6597), .B(n6596), .Z(out[1279]) );
  XOR U2631 ( .A(in[598]), .B(n8519), .Z(n7414) );
  XNOR U2632 ( .A(in[253]), .B(n8618), .Z(n8342) );
  XNOR U2633 ( .A(in[1409]), .B(n8373), .Z(n8339) );
  NAND U2634 ( .A(n8342), .B(n8339), .Z(n6598) );
  XNOR U2635 ( .A(n7414), .B(n6598), .Z(out[127]) );
  XNOR U2636 ( .A(in[50]), .B(n8759), .Z(n6741) );
  XOR U2637 ( .A(in[1536]), .B(n8419), .Z(n7013) );
  XNOR U2638 ( .A(in[1172]), .B(n8436), .Z(n7011) );
  NAND U2639 ( .A(n7013), .B(n7011), .Z(n6599) );
  XNOR U2640 ( .A(n6741), .B(n6599), .Z(out[1280]) );
  XNOR U2641 ( .A(in[51]), .B(n8761), .Z(n6743) );
  XOR U2642 ( .A(in[1537]), .B(n8423), .Z(n7018) );
  XNOR U2643 ( .A(in[1173]), .B(n8440), .Z(n7016) );
  NAND U2644 ( .A(n7018), .B(n7016), .Z(n6600) );
  XNOR U2645 ( .A(n6743), .B(n6600), .Z(out[1281]) );
  XNOR U2646 ( .A(in[52]), .B(n8763), .Z(n6746) );
  XOR U2647 ( .A(in[1538]), .B(n8431), .Z(n7024) );
  XNOR U2648 ( .A(in[1174]), .B(n8444), .Z(n7021) );
  NAND U2649 ( .A(n7024), .B(n7021), .Z(n6601) );
  XNOR U2650 ( .A(n6746), .B(n6601), .Z(out[1282]) );
  XNOR U2651 ( .A(in[53]), .B(n8765), .Z(n6748) );
  XOR U2652 ( .A(in[1539]), .B(n8435), .Z(n7027) );
  XNOR U2653 ( .A(in[1175]), .B(n8448), .Z(n7025) );
  NAND U2654 ( .A(n7027), .B(n7025), .Z(n6602) );
  XNOR U2655 ( .A(n6748), .B(n6602), .Z(out[1283]) );
  XNOR U2656 ( .A(in[54]), .B(n8767), .Z(n6750) );
  XNOR U2657 ( .A(in[1540]), .B(n8439), .Z(n7034) );
  XNOR U2658 ( .A(in[1176]), .B(n8452), .Z(n7031) );
  NAND U2659 ( .A(n7034), .B(n7031), .Z(n6603) );
  XNOR U2660 ( .A(n6750), .B(n6603), .Z(out[1284]) );
  XNOR U2661 ( .A(in[55]), .B(n8769), .Z(n6752) );
  XNOR U2662 ( .A(in[1541]), .B(n8443), .Z(n7038) );
  XNOR U2663 ( .A(in[1177]), .B(n8456), .Z(n7035) );
  NAND U2664 ( .A(n7038), .B(n7035), .Z(n6604) );
  XNOR U2665 ( .A(n6752), .B(n6604), .Z(out[1285]) );
  XNOR U2666 ( .A(in[56]), .B(n8625), .Z(n6754) );
  XNOR U2667 ( .A(in[1542]), .B(n8447), .Z(n7042) );
  XNOR U2668 ( .A(in[1178]), .B(n8460), .Z(n7039) );
  NAND U2669 ( .A(n7042), .B(n7039), .Z(n6605) );
  XNOR U2670 ( .A(n6754), .B(n6605), .Z(out[1286]) );
  XNOR U2671 ( .A(in[57]), .B(n8627), .Z(n6756) );
  XNOR U2672 ( .A(in[1543]), .B(n8451), .Z(n7045) );
  XNOR U2673 ( .A(in[1179]), .B(n8464), .Z(n7043) );
  NAND U2674 ( .A(n7045), .B(n7043), .Z(n6606) );
  XNOR U2675 ( .A(n6756), .B(n6606), .Z(out[1287]) );
  XNOR U2676 ( .A(in[58]), .B(n8629), .Z(n6758) );
  XNOR U2677 ( .A(in[1544]), .B(n8455), .Z(n7051) );
  XNOR U2678 ( .A(in[1180]), .B(n8468), .Z(n7048) );
  NAND U2679 ( .A(n7051), .B(n7048), .Z(n6607) );
  XNOR U2680 ( .A(n6758), .B(n6607), .Z(out[1288]) );
  XNOR U2681 ( .A(in[59]), .B(n8631), .Z(n6760) );
  XNOR U2682 ( .A(in[1545]), .B(n8459), .Z(n7055) );
  XNOR U2683 ( .A(in[1181]), .B(n8476), .Z(n7052) );
  NAND U2684 ( .A(n7055), .B(n7052), .Z(n6608) );
  XNOR U2685 ( .A(n6760), .B(n6608), .Z(out[1289]) );
  XNOR U2686 ( .A(in[665]), .B(n8699), .Z(n7417) );
  XNOR U2687 ( .A(in[599]), .B(n8523), .Z(n8386) );
  NAND U2688 ( .A(n8386), .B(n8384), .Z(n6609) );
  XNOR U2689 ( .A(n7417), .B(n6609), .Z(out[128]) );
  XNOR U2690 ( .A(in[60]), .B(n8633), .Z(n6762) );
  XNOR U2691 ( .A(in[1546]), .B(n8463), .Z(n7059) );
  XNOR U2692 ( .A(in[1182]), .B(n8480), .Z(n7056) );
  NAND U2693 ( .A(n7059), .B(n7056), .Z(n6610) );
  XNOR U2694 ( .A(n6762), .B(n6610), .Z(out[1290]) );
  XNOR U2695 ( .A(in[61]), .B(n8635), .Z(n6764) );
  XNOR U2696 ( .A(in[1547]), .B(n8467), .Z(n7063) );
  XNOR U2697 ( .A(in[1183]), .B(n8484), .Z(n7060) );
  NAND U2698 ( .A(n7063), .B(n7060), .Z(n6611) );
  XNOR U2699 ( .A(n6764), .B(n6611), .Z(out[1291]) );
  XNOR U2700 ( .A(in[62]), .B(n8641), .Z(n6767) );
  XNOR U2701 ( .A(in[1548]), .B(n8475), .Z(n7067) );
  XNOR U2702 ( .A(in[1184]), .B(n8488), .Z(n7064) );
  NAND U2703 ( .A(n7067), .B(n7064), .Z(n6612) );
  XNOR U2704 ( .A(n6767), .B(n6612), .Z(out[1292]) );
  XNOR U2705 ( .A(in[63]), .B(n8643), .Z(n6769) );
  XNOR U2706 ( .A(in[1549]), .B(n8479), .Z(n7071) );
  XNOR U2707 ( .A(in[1185]), .B(n8492), .Z(n7068) );
  NAND U2708 ( .A(n7071), .B(n7068), .Z(n6613) );
  XNOR U2709 ( .A(n6769), .B(n6613), .Z(out[1293]) );
  XNOR U2710 ( .A(in[0]), .B(n8645), .Z(n6771) );
  XNOR U2711 ( .A(in[1550]), .B(n8483), .Z(n7076) );
  XOR U2712 ( .A(n8496), .B(in[1186]), .Z(n7073) );
  NAND U2713 ( .A(n7076), .B(n7073), .Z(n6614) );
  XNOR U2714 ( .A(n6771), .B(n6614), .Z(out[1294]) );
  XNOR U2715 ( .A(in[1]), .B(n8647), .Z(n6773) );
  XNOR U2716 ( .A(in[1551]), .B(n8487), .Z(n7079) );
  XOR U2717 ( .A(n8500), .B(in[1187]), .Z(n7077) );
  NAND U2718 ( .A(n7079), .B(n7077), .Z(n6615) );
  XNOR U2719 ( .A(n6773), .B(n6615), .Z(out[1295]) );
  XNOR U2720 ( .A(in[2]), .B(n8649), .Z(n6775) );
  XNOR U2721 ( .A(in[1552]), .B(n8491), .Z(n7085) );
  XOR U2722 ( .A(n8504), .B(in[1188]), .Z(n7082) );
  NAND U2723 ( .A(n7085), .B(n7082), .Z(n6616) );
  XNOR U2724 ( .A(n6775), .B(n6616), .Z(out[1296]) );
  XNOR U2725 ( .A(in[3]), .B(n8651), .Z(n6777) );
  XNOR U2726 ( .A(in[1553]), .B(n8495), .Z(n7089) );
  XOR U2727 ( .A(n8508), .B(in[1189]), .Z(n7086) );
  NAND U2728 ( .A(n7089), .B(n7086), .Z(n6617) );
  XNOR U2729 ( .A(n6777), .B(n6617), .Z(out[1297]) );
  XNOR U2730 ( .A(in[4]), .B(n8653), .Z(n6779) );
  XNOR U2731 ( .A(in[1554]), .B(n8499), .Z(n7093) );
  XNOR U2732 ( .A(in[1190]), .B(n8512), .Z(n7090) );
  NAND U2733 ( .A(n7093), .B(n7090), .Z(n6618) );
  XNOR U2734 ( .A(n6779), .B(n6618), .Z(out[1298]) );
  XNOR U2735 ( .A(in[5]), .B(n8655), .Z(n6781) );
  XNOR U2736 ( .A(in[1555]), .B(n8503), .Z(n7097) );
  XNOR U2737 ( .A(in[1191]), .B(n8520), .Z(n7094) );
  NAND U2738 ( .A(n7097), .B(n7094), .Z(n6619) );
  XNOR U2739 ( .A(n6781), .B(n6619), .Z(out[1299]) );
  XNOR U2740 ( .A(in[666]), .B(n8701), .Z(n7419) );
  XNOR U2741 ( .A(in[600]), .B(n8527), .Z(n8430) );
  XOR U2742 ( .A(in[255]), .B(n8344), .Z(n8428) );
  NAND U2743 ( .A(n8430), .B(n8428), .Z(n6620) );
  XNOR U2744 ( .A(n7419), .B(n6620), .Z(out[129]) );
  XOR U2745 ( .A(in[202]), .B(n8392), .Z(n8778) );
  XNOR U2746 ( .A(in[1422]), .B(n8433), .Z(n8777) );
  XOR U2747 ( .A(in[1045]), .B(n8933), .Z(n7445) );
  NAND U2748 ( .A(n8777), .B(n7445), .Z(n6621) );
  XNOR U2749 ( .A(n8778), .B(n6621), .Z(out[12]) );
  XNOR U2750 ( .A(in[6]), .B(n8657), .Z(n6783) );
  XNOR U2751 ( .A(in[1556]), .B(n8507), .Z(n7101) );
  XNOR U2752 ( .A(in[1192]), .B(n8524), .Z(n7098) );
  NAND U2753 ( .A(n7101), .B(n7098), .Z(n6622) );
  XNOR U2754 ( .A(n6783), .B(n6622), .Z(out[1300]) );
  XNOR U2755 ( .A(in[7]), .B(n8659), .Z(n6785) );
  XNOR U2756 ( .A(in[1557]), .B(n8511), .Z(n7105) );
  XNOR U2757 ( .A(in[1193]), .B(n8528), .Z(n7102) );
  NAND U2758 ( .A(n7105), .B(n7102), .Z(n6623) );
  XNOR U2759 ( .A(n6785), .B(n6623), .Z(out[1301]) );
  XNOR U2760 ( .A(in[8]), .B(n8663), .Z(n6788) );
  XNOR U2761 ( .A(in[1558]), .B(n8519), .Z(n7109) );
  XNOR U2762 ( .A(in[1194]), .B(n8532), .Z(n7106) );
  NAND U2763 ( .A(n7109), .B(n7106), .Z(n6624) );
  XNOR U2764 ( .A(n6788), .B(n6624), .Z(out[1302]) );
  XNOR U2765 ( .A(in[9]), .B(n8665), .Z(n6790) );
  XNOR U2766 ( .A(in[1559]), .B(n8523), .Z(n7113) );
  XNOR U2767 ( .A(in[1195]), .B(n8536), .Z(n7110) );
  NAND U2768 ( .A(n7113), .B(n7110), .Z(n6625) );
  XNOR U2769 ( .A(n6790), .B(n6625), .Z(out[1303]) );
  XNOR U2770 ( .A(in[10]), .B(n8667), .Z(n6792) );
  XNOR U2771 ( .A(in[1560]), .B(n8527), .Z(n7118) );
  XNOR U2772 ( .A(in[1196]), .B(n8540), .Z(n7115) );
  NAND U2773 ( .A(n7118), .B(n7115), .Z(n6626) );
  XNOR U2774 ( .A(n6792), .B(n6626), .Z(out[1304]) );
  XNOR U2775 ( .A(in[11]), .B(n8669), .Z(n6794) );
  XNOR U2776 ( .A(in[1561]), .B(n8531), .Z(n7122) );
  XNOR U2777 ( .A(in[1197]), .B(n8544), .Z(n7119) );
  NAND U2778 ( .A(n7122), .B(n7119), .Z(n6627) );
  XNOR U2779 ( .A(n6794), .B(n6627), .Z(out[1305]) );
  XNOR U2780 ( .A(in[12]), .B(n8671), .Z(n6796) );
  XNOR U2781 ( .A(in[1562]), .B(n8535), .Z(n7126) );
  XNOR U2782 ( .A(in[1198]), .B(n8548), .Z(n7123) );
  NAND U2783 ( .A(n7126), .B(n7123), .Z(n6628) );
  XNOR U2784 ( .A(n6796), .B(n6628), .Z(out[1306]) );
  XNOR U2785 ( .A(in[13]), .B(n8673), .Z(n6798) );
  XNOR U2786 ( .A(in[1563]), .B(n8539), .Z(n7130) );
  XNOR U2787 ( .A(in[1199]), .B(n8552), .Z(n7127) );
  NAND U2788 ( .A(n7130), .B(n7127), .Z(n6629) );
  XNOR U2789 ( .A(n6798), .B(n6629), .Z(out[1307]) );
  XNOR U2790 ( .A(in[14]), .B(n8675), .Z(n6800) );
  XNOR U2791 ( .A(in[1564]), .B(n8543), .Z(n7134) );
  XNOR U2792 ( .A(in[1200]), .B(n8556), .Z(n7131) );
  NAND U2793 ( .A(n7134), .B(n7131), .Z(n6630) );
  XNOR U2794 ( .A(n6800), .B(n6630), .Z(out[1308]) );
  XNOR U2795 ( .A(in[15]), .B(n8677), .Z(n6802) );
  XNOR U2796 ( .A(in[1565]), .B(n8547), .Z(n7138) );
  XNOR U2797 ( .A(in[1201]), .B(n8564), .Z(n7135) );
  NAND U2798 ( .A(n7138), .B(n7135), .Z(n6631) );
  XNOR U2799 ( .A(n6802), .B(n6631), .Z(out[1309]) );
  XNOR U2800 ( .A(in[667]), .B(n8703), .Z(n7422) );
  XNOR U2801 ( .A(in[601]), .B(n8531), .Z(n8474) );
  XOR U2802 ( .A(in[192]), .B(n8348), .Z(n8471) );
  NAND U2803 ( .A(n8474), .B(n8471), .Z(n6632) );
  XNOR U2804 ( .A(n7422), .B(n6632), .Z(out[130]) );
  XNOR U2805 ( .A(in[16]), .B(n8679), .Z(n6804) );
  XNOR U2806 ( .A(in[1566]), .B(n8551), .Z(n7142) );
  XNOR U2807 ( .A(in[1202]), .B(n8568), .Z(n7139) );
  NAND U2808 ( .A(n7142), .B(n7139), .Z(n6633) );
  XNOR U2809 ( .A(n6804), .B(n6633), .Z(out[1310]) );
  XNOR U2810 ( .A(in[17]), .B(n8681), .Z(n6806) );
  XNOR U2811 ( .A(in[1567]), .B(n8555), .Z(n7145) );
  XNOR U2812 ( .A(in[1203]), .B(n8572), .Z(n7143) );
  NAND U2813 ( .A(n7145), .B(n7143), .Z(n6634) );
  XNOR U2814 ( .A(n6806), .B(n6634), .Z(out[1311]) );
  XNOR U2815 ( .A(in[18]), .B(n8685), .Z(n6809) );
  XNOR U2816 ( .A(in[1568]), .B(n8563), .Z(n7151) );
  XNOR U2817 ( .A(in[1204]), .B(n8576), .Z(n7148) );
  NAND U2818 ( .A(n7151), .B(n7148), .Z(n6635) );
  XNOR U2819 ( .A(n6809), .B(n6635), .Z(out[1312]) );
  XNOR U2820 ( .A(in[19]), .B(n8687), .Z(n6811) );
  XNOR U2821 ( .A(in[1569]), .B(n8567), .Z(n7155) );
  XNOR U2822 ( .A(in[1205]), .B(n8580), .Z(n7152) );
  NAND U2823 ( .A(n7155), .B(n7152), .Z(n6636) );
  XNOR U2824 ( .A(n6811), .B(n6636), .Z(out[1313]) );
  XNOR U2825 ( .A(in[20]), .B(n8689), .Z(n6813) );
  XNOR U2826 ( .A(in[1570]), .B(n8571), .Z(n7160) );
  XNOR U2827 ( .A(in[1206]), .B(n8584), .Z(n7157) );
  NAND U2828 ( .A(n7160), .B(n7157), .Z(n6637) );
  XNOR U2829 ( .A(n6813), .B(n6637), .Z(out[1314]) );
  XNOR U2830 ( .A(in[21]), .B(n8691), .Z(n6815) );
  XNOR U2831 ( .A(in[1571]), .B(n8575), .Z(n7164) );
  XNOR U2832 ( .A(in[1207]), .B(n8588), .Z(n7161) );
  NAND U2833 ( .A(n7164), .B(n7161), .Z(n6638) );
  XNOR U2834 ( .A(n6815), .B(n6638), .Z(out[1315]) );
  XNOR U2835 ( .A(in[22]), .B(n8693), .Z(n6817) );
  XNOR U2836 ( .A(in[1572]), .B(n8579), .Z(n7168) );
  XNOR U2837 ( .A(in[1208]), .B(n8592), .Z(n7165) );
  NAND U2838 ( .A(n7168), .B(n7165), .Z(n6639) );
  XNOR U2839 ( .A(n6817), .B(n6639), .Z(out[1316]) );
  XNOR U2840 ( .A(in[23]), .B(n8695), .Z(n6819) );
  XOR U2841 ( .A(in[1573]), .B(n8583), .Z(n7172) );
  XNOR U2842 ( .A(in[1209]), .B(n8596), .Z(n7169) );
  NAND U2843 ( .A(n7172), .B(n7169), .Z(n6640) );
  XNOR U2844 ( .A(n6819), .B(n6640), .Z(out[1317]) );
  XNOR U2845 ( .A(in[24]), .B(n8697), .Z(n6821) );
  XOR U2846 ( .A(in[1574]), .B(n8587), .Z(n7176) );
  XNOR U2847 ( .A(in[1210]), .B(n8600), .Z(n7173) );
  NAND U2848 ( .A(n7176), .B(n7173), .Z(n6641) );
  XNOR U2849 ( .A(n6821), .B(n6641), .Z(out[1318]) );
  XNOR U2850 ( .A(in[25]), .B(n8699), .Z(n6823) );
  XOR U2851 ( .A(in[1575]), .B(n8591), .Z(n7180) );
  XOR U2852 ( .A(in[1211]), .B(n8610), .Z(n7177) );
  NAND U2853 ( .A(n7180), .B(n7177), .Z(n6642) );
  XNOR U2854 ( .A(n6823), .B(n6642), .Z(out[1319]) );
  XNOR U2855 ( .A(in[668]), .B(n8707), .Z(n7424) );
  XNOR U2856 ( .A(in[602]), .B(n8535), .Z(n8518) );
  XOR U2857 ( .A(in[193]), .B(n8352), .Z(n8515) );
  NAND U2858 ( .A(n8518), .B(n8515), .Z(n6643) );
  XNOR U2859 ( .A(n7424), .B(n6643), .Z(out[131]) );
  XNOR U2860 ( .A(in[26]), .B(n8701), .Z(n6825) );
  XOR U2861 ( .A(in[1576]), .B(n8595), .Z(n7184) );
  XOR U2862 ( .A(in[1212]), .B(n8614), .Z(n7181) );
  NAND U2863 ( .A(n7184), .B(n7181), .Z(n6644) );
  XNOR U2864 ( .A(n6825), .B(n6644), .Z(out[1320]) );
  XNOR U2865 ( .A(in[27]), .B(n8703), .Z(n6827) );
  XOR U2866 ( .A(in[1577]), .B(n8599), .Z(n7188) );
  XOR U2867 ( .A(in[1213]), .B(n8618), .Z(n7185) );
  NAND U2868 ( .A(n7188), .B(n7185), .Z(n6645) );
  XNOR U2869 ( .A(n6827), .B(n6645), .Z(out[1321]) );
  XNOR U2870 ( .A(in[28]), .B(n8707), .Z(n6830) );
  XOR U2871 ( .A(in[1578]), .B(n8609), .Z(n7192) );
  XNOR U2872 ( .A(in[1214]), .B(n8622), .Z(n7189) );
  NAND U2873 ( .A(n7192), .B(n7189), .Z(n6646) );
  XNOR U2874 ( .A(n6830), .B(n6646), .Z(out[1322]) );
  XNOR U2875 ( .A(in[29]), .B(n8709), .Z(n6832) );
  XOR U2876 ( .A(in[1579]), .B(n8613), .Z(n7196) );
  XOR U2877 ( .A(in[1215]), .B(n8344), .Z(n7193) );
  NAND U2878 ( .A(n7196), .B(n7193), .Z(n6647) );
  XNOR U2879 ( .A(n6832), .B(n6647), .Z(out[1323]) );
  XNOR U2880 ( .A(in[30]), .B(n8711), .Z(n6834) );
  XOR U2881 ( .A(in[1580]), .B(n8617), .Z(n7201) );
  XOR U2882 ( .A(in[1152]), .B(n8348), .Z(n7198) );
  NAND U2883 ( .A(n7201), .B(n7198), .Z(n6648) );
  XNOR U2884 ( .A(n6834), .B(n6648), .Z(out[1324]) );
  XNOR U2885 ( .A(in[31]), .B(n8713), .Z(n6836) );
  XOR U2886 ( .A(in[1581]), .B(n8621), .Z(n7205) );
  XOR U2887 ( .A(in[1153]), .B(n8352), .Z(n7202) );
  NAND U2888 ( .A(n7205), .B(n7202), .Z(n6649) );
  XNOR U2889 ( .A(n6836), .B(n6649), .Z(out[1325]) );
  XNOR U2890 ( .A(in[32]), .B(n8715), .Z(n6838) );
  XOR U2891 ( .A(in[1582]), .B(n8343), .Z(n7209) );
  XOR U2892 ( .A(in[1154]), .B(n8356), .Z(n7206) );
  NAND U2893 ( .A(n7209), .B(n7206), .Z(n6650) );
  XNOR U2894 ( .A(n6838), .B(n6650), .Z(out[1326]) );
  XNOR U2895 ( .A(in[33]), .B(n8717), .Z(n6840) );
  XOR U2896 ( .A(in[1583]), .B(n8347), .Z(n7213) );
  XOR U2897 ( .A(in[1155]), .B(n8360), .Z(n7210) );
  NAND U2898 ( .A(n7213), .B(n7210), .Z(n6651) );
  XNOR U2899 ( .A(n6840), .B(n6651), .Z(out[1327]) );
  XNOR U2900 ( .A(in[34]), .B(n8719), .Z(n6842) );
  XOR U2901 ( .A(in[1584]), .B(n8351), .Z(n7217) );
  XOR U2902 ( .A(in[1156]), .B(n8364), .Z(n7214) );
  NAND U2903 ( .A(n7217), .B(n7214), .Z(n6652) );
  XNOR U2904 ( .A(n6842), .B(n6652), .Z(out[1328]) );
  XNOR U2905 ( .A(in[35]), .B(n8721), .Z(n6844) );
  XOR U2906 ( .A(in[1585]), .B(n8355), .Z(n7221) );
  XOR U2907 ( .A(in[1157]), .B(n8368), .Z(n7218) );
  NAND U2908 ( .A(n7221), .B(n7218), .Z(n6653) );
  XNOR U2909 ( .A(n6844), .B(n6653), .Z(out[1329]) );
  XNOR U2910 ( .A(in[669]), .B(n8709), .Z(n7427) );
  XNOR U2911 ( .A(in[603]), .B(n8539), .Z(n8562) );
  XOR U2912 ( .A(in[194]), .B(n8356), .Z(n8559) );
  NAND U2913 ( .A(n8562), .B(n8559), .Z(n6654) );
  XNOR U2914 ( .A(n7427), .B(n6654), .Z(out[132]) );
  XNOR U2915 ( .A(in[36]), .B(n8723), .Z(n6846) );
  XOR U2916 ( .A(in[1586]), .B(n8359), .Z(n7225) );
  XOR U2917 ( .A(in[1158]), .B(n8372), .Z(n7222) );
  NAND U2918 ( .A(n7225), .B(n7222), .Z(n6655) );
  XNOR U2919 ( .A(n6846), .B(n6655), .Z(out[1330]) );
  XNOR U2920 ( .A(in[37]), .B(n8725), .Z(n6848) );
  XOR U2921 ( .A(in[1587]), .B(n8363), .Z(n7229) );
  XOR U2922 ( .A(in[1159]), .B(n8376), .Z(n7226) );
  NAND U2923 ( .A(n7229), .B(n7226), .Z(n6656) );
  XNOR U2924 ( .A(n6848), .B(n6656), .Z(out[1331]) );
  XNOR U2925 ( .A(in[38]), .B(n8731), .Z(n6851) );
  XOR U2926 ( .A(in[1588]), .B(n8367), .Z(n7233) );
  XOR U2927 ( .A(in[1160]), .B(n8380), .Z(n7230) );
  NAND U2928 ( .A(n7233), .B(n7230), .Z(n6657) );
  XNOR U2929 ( .A(n6851), .B(n6657), .Z(out[1332]) );
  XNOR U2930 ( .A(in[39]), .B(n8733), .Z(n6853) );
  XOR U2931 ( .A(in[1589]), .B(n8371), .Z(n7237) );
  XOR U2932 ( .A(in[1161]), .B(n8388), .Z(n7234) );
  NAND U2933 ( .A(n7237), .B(n7234), .Z(n6658) );
  XNOR U2934 ( .A(n6853), .B(n6658), .Z(out[1333]) );
  XNOR U2935 ( .A(in[40]), .B(n8735), .Z(n6855) );
  XOR U2936 ( .A(in[1590]), .B(n8375), .Z(n7242) );
  XOR U2937 ( .A(in[1162]), .B(n8392), .Z(n7239) );
  NAND U2938 ( .A(n7242), .B(n7239), .Z(n6659) );
  XNOR U2939 ( .A(n6855), .B(n6659), .Z(out[1334]) );
  XNOR U2940 ( .A(in[41]), .B(n8737), .Z(n6857) );
  XOR U2941 ( .A(in[1591]), .B(n8379), .Z(n7246) );
  XOR U2942 ( .A(in[1163]), .B(n8396), .Z(n7243) );
  NAND U2943 ( .A(n7246), .B(n7243), .Z(n6660) );
  XNOR U2944 ( .A(n6857), .B(n6660), .Z(out[1335]) );
  XNOR U2945 ( .A(in[42]), .B(n8739), .Z(n6859) );
  XOR U2946 ( .A(in[1592]), .B(n8387), .Z(n7250) );
  XOR U2947 ( .A(in[1164]), .B(n8400), .Z(n7247) );
  NAND U2948 ( .A(n7250), .B(n7247), .Z(n6661) );
  XNOR U2949 ( .A(n6859), .B(n6661), .Z(out[1336]) );
  XNOR U2950 ( .A(in[43]), .B(n8741), .Z(n6861) );
  XOR U2951 ( .A(in[1593]), .B(n8391), .Z(n7254) );
  XOR U2952 ( .A(in[1165]), .B(n8404), .Z(n7251) );
  NAND U2953 ( .A(n7254), .B(n7251), .Z(n6662) );
  XNOR U2954 ( .A(n6861), .B(n6662), .Z(out[1337]) );
  XNOR U2955 ( .A(in[44]), .B(n8743), .Z(n6863) );
  XOR U2956 ( .A(in[1594]), .B(n8395), .Z(n7258) );
  XOR U2957 ( .A(in[1166]), .B(n8408), .Z(n7255) );
  NAND U2958 ( .A(n7258), .B(n7255), .Z(n6663) );
  XNOR U2959 ( .A(n6863), .B(n6663), .Z(out[1338]) );
  XNOR U2960 ( .A(in[45]), .B(n8745), .Z(n6865) );
  XOR U2961 ( .A(in[1595]), .B(n8399), .Z(n7262) );
  XOR U2962 ( .A(in[1167]), .B(n8412), .Z(n7259) );
  NAND U2963 ( .A(n7262), .B(n7259), .Z(n6664) );
  XNOR U2964 ( .A(n6865), .B(n6664), .Z(out[1339]) );
  XNOR U2965 ( .A(in[670]), .B(n8711), .Z(n7429) );
  XNOR U2966 ( .A(in[604]), .B(n8543), .Z(n8606) );
  XOR U2967 ( .A(in[195]), .B(n8360), .Z(n8603) );
  NAND U2968 ( .A(n8606), .B(n8603), .Z(n6665) );
  XNOR U2969 ( .A(n7429), .B(n6665), .Z(out[133]) );
  XNOR U2970 ( .A(in[46]), .B(n8747), .Z(n6867) );
  XOR U2971 ( .A(in[1596]), .B(n8403), .Z(n7266) );
  XOR U2972 ( .A(in[1168]), .B(n8416), .Z(n7263) );
  NAND U2973 ( .A(n7266), .B(n7263), .Z(n6666) );
  XNOR U2974 ( .A(n6867), .B(n6666), .Z(out[1340]) );
  XNOR U2975 ( .A(in[47]), .B(n8749), .Z(n6869) );
  XOR U2976 ( .A(in[1597]), .B(n8407), .Z(n7270) );
  XOR U2977 ( .A(in[1169]), .B(n8420), .Z(n7267) );
  NAND U2978 ( .A(n7270), .B(n7267), .Z(n6667) );
  XNOR U2979 ( .A(n6869), .B(n6667), .Z(out[1341]) );
  XNOR U2980 ( .A(in[48]), .B(n8755), .Z(n6872) );
  XOR U2981 ( .A(in[1598]), .B(n8411), .Z(n7274) );
  XOR U2982 ( .A(in[1170]), .B(n8424), .Z(n7271) );
  NAND U2983 ( .A(n7274), .B(n7271), .Z(n6668) );
  XNOR U2984 ( .A(n6872), .B(n6668), .Z(out[1342]) );
  XNOR U2985 ( .A(in[49]), .B(n8757), .Z(n6874) );
  XOR U2986 ( .A(in[1599]), .B(n8415), .Z(n7277) );
  XNOR U2987 ( .A(in[1171]), .B(n8432), .Z(n7275) );
  NAND U2988 ( .A(n7277), .B(n7275), .Z(n6669) );
  XNOR U2989 ( .A(n6874), .B(n6669), .Z(out[1343]) );
  XOR U2990 ( .A(in[427]), .B(n8787), .Z(n6876) );
  NOR U2991 ( .A(n6741), .B(n7013), .Z(n6670) );
  XNOR U2992 ( .A(n6876), .B(n6670), .Z(out[1344]) );
  XOR U2993 ( .A(in[428]), .B(n8790), .Z(n6878) );
  NOR U2994 ( .A(n6743), .B(n7018), .Z(n6671) );
  XNOR U2995 ( .A(n6878), .B(n6671), .Z(out[1345]) );
  XOR U2996 ( .A(in[429]), .B(n8793), .Z(n6880) );
  NOR U2997 ( .A(n6746), .B(n7024), .Z(n6672) );
  XNOR U2998 ( .A(n6880), .B(n6672), .Z(out[1346]) );
  XOR U2999 ( .A(in[430]), .B(n8796), .Z(n6882) );
  NOR U3000 ( .A(n6748), .B(n7027), .Z(n6673) );
  XNOR U3001 ( .A(n6882), .B(n6673), .Z(out[1347]) );
  XOR U3002 ( .A(in[431]), .B(n8799), .Z(n6884) );
  NOR U3003 ( .A(n6750), .B(n7034), .Z(n6674) );
  XNOR U3004 ( .A(n6884), .B(n6674), .Z(out[1348]) );
  XOR U3005 ( .A(in[432]), .B(n8802), .Z(n6886) );
  NOR U3006 ( .A(n6752), .B(n7038), .Z(n6675) );
  XNOR U3007 ( .A(n6886), .B(n6675), .Z(out[1349]) );
  XNOR U3008 ( .A(in[671]), .B(n8713), .Z(n7431) );
  XNOR U3009 ( .A(in[605]), .B(n8547), .Z(n8640) );
  XOR U3010 ( .A(in[196]), .B(n8364), .Z(n8637) );
  NAND U3011 ( .A(n8640), .B(n8637), .Z(n6676) );
  XNOR U3012 ( .A(n7431), .B(n6676), .Z(out[134]) );
  XOR U3013 ( .A(in[433]), .B(n8805), .Z(n6888) );
  NOR U3014 ( .A(n6754), .B(n7042), .Z(n6677) );
  XNOR U3015 ( .A(n6888), .B(n6677), .Z(out[1350]) );
  XOR U3016 ( .A(in[434]), .B(n8808), .Z(n6890) );
  NOR U3017 ( .A(n6756), .B(n7045), .Z(n6678) );
  XNOR U3018 ( .A(n6890), .B(n6678), .Z(out[1351]) );
  XOR U3019 ( .A(in[435]), .B(n8815), .Z(n6893) );
  NOR U3020 ( .A(n6758), .B(n7051), .Z(n6679) );
  XNOR U3021 ( .A(n6893), .B(n6679), .Z(out[1352]) );
  XOR U3022 ( .A(in[436]), .B(n8818), .Z(n6895) );
  NOR U3023 ( .A(n6760), .B(n7055), .Z(n6680) );
  XNOR U3024 ( .A(n6895), .B(n6680), .Z(out[1353]) );
  XOR U3025 ( .A(in[437]), .B(n8821), .Z(n6897) );
  NOR U3026 ( .A(n6762), .B(n7059), .Z(n6681) );
  XNOR U3027 ( .A(n6897), .B(n6681), .Z(out[1354]) );
  XOR U3028 ( .A(in[438]), .B(n8824), .Z(n6899) );
  NOR U3029 ( .A(n6764), .B(n7063), .Z(n6682) );
  XNOR U3030 ( .A(n6899), .B(n6682), .Z(out[1355]) );
  XOR U3031 ( .A(in[439]), .B(n8827), .Z(n6901) );
  NOR U3032 ( .A(n6767), .B(n7067), .Z(n6683) );
  XNOR U3033 ( .A(n6901), .B(n6683), .Z(out[1356]) );
  XOR U3034 ( .A(in[440]), .B(n8830), .Z(n6903) );
  NOR U3035 ( .A(n6769), .B(n7071), .Z(n6684) );
  XNOR U3036 ( .A(n6903), .B(n6684), .Z(out[1357]) );
  XOR U3037 ( .A(in[441]), .B(n8833), .Z(n6905) );
  NOR U3038 ( .A(n6771), .B(n7076), .Z(n6685) );
  XNOR U3039 ( .A(n6905), .B(n6685), .Z(out[1358]) );
  XOR U3040 ( .A(in[442]), .B(n8836), .Z(n6907) );
  NOR U3041 ( .A(n6773), .B(n7079), .Z(n6686) );
  XNOR U3042 ( .A(n6907), .B(n6686), .Z(out[1359]) );
  XNOR U3043 ( .A(in[672]), .B(n8715), .Z(n7433) );
  XNOR U3044 ( .A(in[606]), .B(n8551), .Z(n8662) );
  XOR U3045 ( .A(in[197]), .B(n8368), .Z(n8886) );
  NAND U3046 ( .A(n8662), .B(n8886), .Z(n6687) );
  XNOR U3047 ( .A(n7433), .B(n6687), .Z(out[135]) );
  XOR U3048 ( .A(in[443]), .B(n8839), .Z(n6909) );
  NOR U3049 ( .A(n6775), .B(n7085), .Z(n6688) );
  XNOR U3050 ( .A(n6909), .B(n6688), .Z(out[1360]) );
  XOR U3051 ( .A(in[444]), .B(n8842), .Z(n6911) );
  NOR U3052 ( .A(n6777), .B(n7089), .Z(n6689) );
  XNOR U3053 ( .A(n6911), .B(n6689), .Z(out[1361]) );
  XOR U3054 ( .A(in[445]), .B(n8849), .Z(n6914) );
  NOR U3055 ( .A(n6779), .B(n7093), .Z(n6690) );
  XNOR U3056 ( .A(n6914), .B(n6690), .Z(out[1362]) );
  XOR U3057 ( .A(in[446]), .B(n8852), .Z(n6916) );
  NOR U3058 ( .A(n6781), .B(n7097), .Z(n6691) );
  XNOR U3059 ( .A(n6916), .B(n6691), .Z(out[1363]) );
  XOR U3060 ( .A(in[447]), .B(n8855), .Z(n6918) );
  NOR U3061 ( .A(n6783), .B(n7101), .Z(n6692) );
  XNOR U3062 ( .A(n6918), .B(n6692), .Z(out[1364]) );
  XOR U3063 ( .A(in[384]), .B(n8858), .Z(n6920) );
  NOR U3064 ( .A(n6785), .B(n7105), .Z(n6693) );
  XNOR U3065 ( .A(n6920), .B(n6693), .Z(out[1365]) );
  XOR U3066 ( .A(in[385]), .B(n8861), .Z(n6922) );
  NOR U3067 ( .A(n6788), .B(n7109), .Z(n6694) );
  XNOR U3068 ( .A(n6922), .B(n6694), .Z(out[1366]) );
  XOR U3069 ( .A(in[386]), .B(n8864), .Z(n6924) );
  NOR U3070 ( .A(n6790), .B(n7113), .Z(n6695) );
  XNOR U3071 ( .A(n6924), .B(n6695), .Z(out[1367]) );
  XOR U3072 ( .A(in[387]), .B(n8867), .Z(n6926) );
  NOR U3073 ( .A(n6792), .B(n7118), .Z(n6696) );
  XNOR U3074 ( .A(n6926), .B(n6696), .Z(out[1368]) );
  XOR U3075 ( .A(in[388]), .B(n8870), .Z(n6928) );
  NOR U3076 ( .A(n6794), .B(n7122), .Z(n6697) );
  XNOR U3077 ( .A(n6928), .B(n6697), .Z(out[1369]) );
  XNOR U3078 ( .A(in[673]), .B(n8717), .Z(n7435) );
  XNOR U3079 ( .A(in[607]), .B(n8555), .Z(n8684) );
  XOR U3080 ( .A(in[198]), .B(n8372), .Z(n9170) );
  NAND U3081 ( .A(n8684), .B(n9170), .Z(n6698) );
  XNOR U3082 ( .A(n7435), .B(n6698), .Z(out[136]) );
  XOR U3083 ( .A(in[389]), .B(n8873), .Z(n6930) );
  NOR U3084 ( .A(n6796), .B(n7126), .Z(n6699) );
  XNOR U3085 ( .A(n6930), .B(n6699), .Z(out[1370]) );
  XOR U3086 ( .A(in[390]), .B(n8876), .Z(n6932) );
  NOR U3087 ( .A(n6798), .B(n7130), .Z(n6700) );
  XNOR U3088 ( .A(n6932), .B(n6700), .Z(out[1371]) );
  XOR U3089 ( .A(in[391]), .B(n8887), .Z(n6936) );
  NOR U3090 ( .A(n6800), .B(n7134), .Z(n6701) );
  XNOR U3091 ( .A(n6936), .B(n6701), .Z(out[1372]) );
  XOR U3092 ( .A(in[392]), .B(n8890), .Z(n6938) );
  NOR U3093 ( .A(n6802), .B(n7138), .Z(n6702) );
  XNOR U3094 ( .A(n6938), .B(n6702), .Z(out[1373]) );
  XOR U3095 ( .A(in[393]), .B(n8893), .Z(n6940) );
  NOR U3096 ( .A(n6804), .B(n7142), .Z(n6703) );
  XNOR U3097 ( .A(n6940), .B(n6703), .Z(out[1374]) );
  XOR U3098 ( .A(in[394]), .B(n8896), .Z(n6942) );
  NOR U3099 ( .A(n6806), .B(n7145), .Z(n6704) );
  XNOR U3100 ( .A(n6942), .B(n6704), .Z(out[1375]) );
  XOR U3101 ( .A(in[395]), .B(n8899), .Z(n6944) );
  NOR U3102 ( .A(n6809), .B(n7151), .Z(n6705) );
  XNOR U3103 ( .A(n6944), .B(n6705), .Z(out[1376]) );
  XNOR U3104 ( .A(n8902), .B(in[396]), .Z(n6946) );
  NOR U3105 ( .A(n6811), .B(n7155), .Z(n6706) );
  XNOR U3106 ( .A(n6946), .B(n6706), .Z(out[1377]) );
  XNOR U3107 ( .A(n8905), .B(in[397]), .Z(n6948) );
  NOR U3108 ( .A(n6813), .B(n7160), .Z(n6707) );
  XNOR U3109 ( .A(n6948), .B(n6707), .Z(out[1378]) );
  XNOR U3110 ( .A(n8908), .B(in[398]), .Z(n6950) );
  NOR U3111 ( .A(n6815), .B(n7164), .Z(n6708) );
  XNOR U3112 ( .A(n6950), .B(n6708), .Z(out[1379]) );
  XNOR U3113 ( .A(in[674]), .B(n8719), .Z(n7437) );
  XNOR U3114 ( .A(in[608]), .B(n8563), .Z(n8706) );
  XOR U3115 ( .A(in[199]), .B(n8376), .Z(n9614) );
  NAND U3116 ( .A(n8706), .B(n9614), .Z(n6709) );
  XNOR U3117 ( .A(n7437), .B(n6709), .Z(out[137]) );
  XNOR U3118 ( .A(n8911), .B(in[399]), .Z(n6952) );
  NOR U3119 ( .A(n6817), .B(n7168), .Z(n6710) );
  XNOR U3120 ( .A(n6952), .B(n6710), .Z(out[1380]) );
  XNOR U3121 ( .A(n8914), .B(in[400]), .Z(n6954) );
  NOR U3122 ( .A(n6819), .B(n7172), .Z(n6711) );
  XNOR U3123 ( .A(n6954), .B(n6711), .Z(out[1381]) );
  XNOR U3124 ( .A(n8921), .B(in[401]), .Z(n6957) );
  NOR U3125 ( .A(n6821), .B(n7176), .Z(n6712) );
  XNOR U3126 ( .A(n6957), .B(n6712), .Z(out[1382]) );
  XNOR U3127 ( .A(n8924), .B(in[402]), .Z(n6959) );
  NOR U3128 ( .A(n6823), .B(n7180), .Z(n6713) );
  XNOR U3129 ( .A(n6959), .B(n6713), .Z(out[1383]) );
  XNOR U3130 ( .A(n8927), .B(in[403]), .Z(n6961) );
  NOR U3131 ( .A(n6825), .B(n7184), .Z(n6714) );
  XNOR U3132 ( .A(n6961), .B(n6714), .Z(out[1384]) );
  XNOR U3133 ( .A(in[404]), .B(n8930), .Z(n6963) );
  NOR U3134 ( .A(n6827), .B(n7188), .Z(n6715) );
  XNOR U3135 ( .A(n6963), .B(n6715), .Z(out[1385]) );
  XNOR U3136 ( .A(in[405]), .B(n8933), .Z(n6965) );
  NOR U3137 ( .A(n6830), .B(n7192), .Z(n6716) );
  XNOR U3138 ( .A(n6965), .B(n6716), .Z(out[1386]) );
  XNOR U3139 ( .A(in[406]), .B(n8936), .Z(n6967) );
  NOR U3140 ( .A(n6832), .B(n7196), .Z(n6717) );
  XNOR U3141 ( .A(n6967), .B(n6717), .Z(out[1387]) );
  XNOR U3142 ( .A(in[407]), .B(n8939), .Z(n6969) );
  NOR U3143 ( .A(n6834), .B(n7201), .Z(n6718) );
  XNOR U3144 ( .A(n6969), .B(n6718), .Z(out[1388]) );
  XNOR U3145 ( .A(in[408]), .B(n8942), .Z(n6971) );
  NOR U3146 ( .A(n6836), .B(n7205), .Z(n6719) );
  XNOR U3147 ( .A(n6971), .B(n6719), .Z(out[1389]) );
  XNOR U3148 ( .A(in[675]), .B(n8721), .Z(n7440) );
  XNOR U3149 ( .A(in[609]), .B(n8567), .Z(n8730) );
  NAND U3150 ( .A(n8730), .B(n8728), .Z(n6720) );
  XNOR U3151 ( .A(n7440), .B(n6720), .Z(out[138]) );
  XNOR U3152 ( .A(in[409]), .B(n8945), .Z(n6973) );
  NOR U3153 ( .A(n6838), .B(n7209), .Z(n6721) );
  XNOR U3154 ( .A(n6973), .B(n6721), .Z(out[1390]) );
  XNOR U3155 ( .A(in[410]), .B(n8948), .Z(n6975) );
  NOR U3156 ( .A(n6840), .B(n7213), .Z(n6722) );
  XNOR U3157 ( .A(n6975), .B(n6722), .Z(out[1391]) );
  XNOR U3158 ( .A(in[411]), .B(n8955), .Z(n6978) );
  NOR U3159 ( .A(n6842), .B(n7217), .Z(n6723) );
  XNOR U3160 ( .A(n6978), .B(n6723), .Z(out[1392]) );
  XNOR U3161 ( .A(in[412]), .B(n8958), .Z(n6980) );
  NOR U3162 ( .A(n6844), .B(n7221), .Z(n6724) );
  XNOR U3163 ( .A(n6980), .B(n6724), .Z(out[1393]) );
  XNOR U3164 ( .A(in[413]), .B(n8961), .Z(n6982) );
  NOR U3165 ( .A(n6846), .B(n7225), .Z(n6725) );
  XNOR U3166 ( .A(n6982), .B(n6725), .Z(out[1394]) );
  XNOR U3167 ( .A(in[414]), .B(n8964), .Z(n6984) );
  NOR U3168 ( .A(n6848), .B(n7229), .Z(n6726) );
  XNOR U3169 ( .A(n6984), .B(n6726), .Z(out[1395]) );
  XNOR U3170 ( .A(in[415]), .B(n8967), .Z(n6986) );
  NOR U3171 ( .A(n6851), .B(n7233), .Z(n6727) );
  XNOR U3172 ( .A(n6986), .B(n6727), .Z(out[1396]) );
  XNOR U3173 ( .A(in[416]), .B(n8970), .Z(n6988) );
  NOR U3174 ( .A(n6853), .B(n7237), .Z(n6728) );
  XNOR U3175 ( .A(n6988), .B(n6728), .Z(out[1397]) );
  XNOR U3176 ( .A(in[417]), .B(n8973), .Z(n6990) );
  NOR U3177 ( .A(n6855), .B(n7242), .Z(n6729) );
  XNOR U3178 ( .A(n6990), .B(n6729), .Z(out[1398]) );
  XNOR U3179 ( .A(in[418]), .B(n8976), .Z(n6992) );
  NOR U3180 ( .A(n6857), .B(n7246), .Z(n6730) );
  XNOR U3181 ( .A(n6992), .B(n6730), .Z(out[1399]) );
  XNOR U3182 ( .A(in[676]), .B(n8723), .Z(n7443) );
  XNOR U3183 ( .A(in[610]), .B(n8571), .Z(n8754) );
  NAND U3184 ( .A(n8754), .B(n8752), .Z(n6731) );
  XNOR U3185 ( .A(n7443), .B(n6731), .Z(out[139]) );
  XOR U3186 ( .A(in[203]), .B(n8396), .Z(n8812) );
  XNOR U3187 ( .A(in[1423]), .B(n8437), .Z(n8811) );
  XOR U3188 ( .A(in[1046]), .B(n8936), .Z(n7448) );
  NAND U3189 ( .A(n8811), .B(n7448), .Z(n6732) );
  XNOR U3190 ( .A(n8812), .B(n6732), .Z(out[13]) );
  XNOR U3191 ( .A(in[419]), .B(n8979), .Z(n6994) );
  NOR U3192 ( .A(n6859), .B(n7250), .Z(n6733) );
  XNOR U3193 ( .A(n6994), .B(n6733), .Z(out[1400]) );
  XOR U3194 ( .A(in[420]), .B(n8982), .Z(n6996) );
  NOR U3195 ( .A(n6861), .B(n7254), .Z(n6734) );
  XNOR U3196 ( .A(n6996), .B(n6734), .Z(out[1401]) );
  XOR U3197 ( .A(in[421]), .B(n8989), .Z(n6999) );
  NOR U3198 ( .A(n6863), .B(n7258), .Z(n6735) );
  XNOR U3199 ( .A(n6999), .B(n6735), .Z(out[1402]) );
  XOR U3200 ( .A(in[422]), .B(n8992), .Z(n7001) );
  NOR U3201 ( .A(n6865), .B(n7262), .Z(n6736) );
  XNOR U3202 ( .A(n7001), .B(n6736), .Z(out[1403]) );
  XOR U3203 ( .A(in[423]), .B(n8771), .Z(n7003) );
  NOR U3204 ( .A(n6867), .B(n7266), .Z(n6737) );
  XNOR U3205 ( .A(n7003), .B(n6737), .Z(out[1404]) );
  XOR U3206 ( .A(in[424]), .B(n8774), .Z(n7005) );
  NOR U3207 ( .A(n6869), .B(n7270), .Z(n6738) );
  XNOR U3208 ( .A(n7005), .B(n6738), .Z(out[1405]) );
  XOR U3209 ( .A(in[425]), .B(n8781), .Z(n7007) );
  NOR U3210 ( .A(n6872), .B(n7274), .Z(n6739) );
  XNOR U3211 ( .A(n7007), .B(n6739), .Z(out[1406]) );
  XOR U3212 ( .A(in[426]), .B(n8784), .Z(n7009) );
  NOR U3213 ( .A(n6874), .B(n7277), .Z(n6740) );
  XNOR U3214 ( .A(n7009), .B(n6740), .Z(out[1407]) );
  XOR U3215 ( .A(in[789]), .B(n8461), .Z(n7012) );
  NAND U3216 ( .A(n6876), .B(n6741), .Z(n6742) );
  XNOR U3217 ( .A(n7012), .B(n6742), .Z(out[1408]) );
  XOR U3218 ( .A(in[790]), .B(n8465), .Z(n7017) );
  NAND U3219 ( .A(n6878), .B(n6743), .Z(n6744) );
  XNOR U3220 ( .A(n7017), .B(n6744), .Z(out[1409]) );
  XNOR U3221 ( .A(in[677]), .B(n8725), .Z(n7446) );
  XNOR U3222 ( .A(in[611]), .B(n8575), .Z(n8780) );
  NAND U3223 ( .A(n8780), .B(n8778), .Z(n6745) );
  XNOR U3224 ( .A(n7446), .B(n6745), .Z(out[140]) );
  XOR U3225 ( .A(in[791]), .B(n8469), .Z(n7022) );
  NAND U3226 ( .A(n6880), .B(n6746), .Z(n6747) );
  XNOR U3227 ( .A(n7022), .B(n6747), .Z(out[1410]) );
  XOR U3228 ( .A(in[792]), .B(n8477), .Z(n7026) );
  NAND U3229 ( .A(n6882), .B(n6748), .Z(n6749) );
  XNOR U3230 ( .A(n7026), .B(n6749), .Z(out[1411]) );
  XOR U3231 ( .A(in[793]), .B(n8481), .Z(n7032) );
  NAND U3232 ( .A(n6884), .B(n6750), .Z(n6751) );
  XNOR U3233 ( .A(n7032), .B(n6751), .Z(out[1412]) );
  XOR U3234 ( .A(in[794]), .B(n8485), .Z(n7036) );
  NAND U3235 ( .A(n6886), .B(n6752), .Z(n6753) );
  XNOR U3236 ( .A(n7036), .B(n6753), .Z(out[1413]) );
  XOR U3237 ( .A(in[795]), .B(n8489), .Z(n7040) );
  NAND U3238 ( .A(n6888), .B(n6754), .Z(n6755) );
  XNOR U3239 ( .A(n7040), .B(n6755), .Z(out[1414]) );
  XOR U3240 ( .A(in[796]), .B(n8493), .Z(n7044) );
  NAND U3241 ( .A(n6890), .B(n6756), .Z(n6757) );
  XNOR U3242 ( .A(n7044), .B(n6757), .Z(out[1415]) );
  XOR U3243 ( .A(in[797]), .B(n8497), .Z(n7049) );
  NAND U3244 ( .A(n6893), .B(n6758), .Z(n6759) );
  XNOR U3245 ( .A(n7049), .B(n6759), .Z(out[1416]) );
  XOR U3246 ( .A(in[798]), .B(n8501), .Z(n7053) );
  NAND U3247 ( .A(n6895), .B(n6760), .Z(n6761) );
  XNOR U3248 ( .A(n7053), .B(n6761), .Z(out[1417]) );
  XOR U3249 ( .A(in[799]), .B(n8505), .Z(n7057) );
  NAND U3250 ( .A(n6897), .B(n6762), .Z(n6763) );
  XNOR U3251 ( .A(n7057), .B(n6763), .Z(out[1418]) );
  XOR U3252 ( .A(in[800]), .B(n8509), .Z(n7061) );
  NAND U3253 ( .A(n6899), .B(n6764), .Z(n6765) );
  XNOR U3254 ( .A(n7061), .B(n6765), .Z(out[1419]) );
  XNOR U3255 ( .A(in[678]), .B(n8731), .Z(n7449) );
  XNOR U3256 ( .A(in[612]), .B(n8579), .Z(n8814) );
  NAND U3257 ( .A(n8814), .B(n8812), .Z(n6766) );
  XNOR U3258 ( .A(n7449), .B(n6766), .Z(out[141]) );
  XOR U3259 ( .A(in[801]), .B(n8513), .Z(n7065) );
  NAND U3260 ( .A(n6901), .B(n6767), .Z(n6768) );
  XNOR U3261 ( .A(n7065), .B(n6768), .Z(out[1420]) );
  XOR U3262 ( .A(in[802]), .B(n8521), .Z(n7069) );
  NAND U3263 ( .A(n6903), .B(n6769), .Z(n6770) );
  XNOR U3264 ( .A(n7069), .B(n6770), .Z(out[1421]) );
  XOR U3265 ( .A(in[803]), .B(n8525), .Z(n7074) );
  NAND U3266 ( .A(n6905), .B(n6771), .Z(n6772) );
  XNOR U3267 ( .A(n7074), .B(n6772), .Z(out[1422]) );
  XOR U3268 ( .A(in[804]), .B(n8529), .Z(n7078) );
  NAND U3269 ( .A(n6907), .B(n6773), .Z(n6774) );
  XNOR U3270 ( .A(n7078), .B(n6774), .Z(out[1423]) );
  XOR U3271 ( .A(in[805]), .B(n8533), .Z(n7083) );
  NAND U3272 ( .A(n6909), .B(n6775), .Z(n6776) );
  XNOR U3273 ( .A(n7083), .B(n6776), .Z(out[1424]) );
  XNOR U3274 ( .A(in[806]), .B(n8537), .Z(n7087) );
  NAND U3275 ( .A(n6911), .B(n6777), .Z(n6778) );
  XNOR U3276 ( .A(n7087), .B(n6778), .Z(out[1425]) );
  XNOR U3277 ( .A(in[807]), .B(n8541), .Z(n7091) );
  NAND U3278 ( .A(n6914), .B(n6779), .Z(n6780) );
  XNOR U3279 ( .A(n7091), .B(n6780), .Z(out[1426]) );
  XNOR U3280 ( .A(in[808]), .B(n8545), .Z(n7095) );
  NAND U3281 ( .A(n6916), .B(n6781), .Z(n6782) );
  XNOR U3282 ( .A(n7095), .B(n6782), .Z(out[1427]) );
  XNOR U3283 ( .A(in[809]), .B(n8549), .Z(n7099) );
  NAND U3284 ( .A(n6918), .B(n6783), .Z(n6784) );
  XNOR U3285 ( .A(n7099), .B(n6784), .Z(out[1428]) );
  XNOR U3286 ( .A(in[810]), .B(n8553), .Z(n7103) );
  NAND U3287 ( .A(n6920), .B(n6785), .Z(n6786) );
  XNOR U3288 ( .A(n7103), .B(n6786), .Z(out[1429]) );
  XNOR U3289 ( .A(in[679]), .B(n8733), .Z(n7453) );
  XOR U3290 ( .A(in[613]), .B(n8583), .Z(n8848) );
  XOR U3291 ( .A(in[204]), .B(n8400), .Z(n8846) );
  NAND U3292 ( .A(n8848), .B(n8846), .Z(n6787) );
  XNOR U3293 ( .A(n7453), .B(n6787), .Z(out[142]) );
  XNOR U3294 ( .A(in[811]), .B(n8557), .Z(n7107) );
  NAND U3295 ( .A(n6922), .B(n6788), .Z(n6789) );
  XNOR U3296 ( .A(n7107), .B(n6789), .Z(out[1430]) );
  XNOR U3297 ( .A(in[812]), .B(n8565), .Z(n7111) );
  NAND U3298 ( .A(n6924), .B(n6790), .Z(n6791) );
  XNOR U3299 ( .A(n7111), .B(n6791), .Z(out[1431]) );
  XNOR U3300 ( .A(in[813]), .B(n8569), .Z(n7116) );
  NAND U3301 ( .A(n6926), .B(n6792), .Z(n6793) );
  XNOR U3302 ( .A(n7116), .B(n6793), .Z(out[1432]) );
  XNOR U3303 ( .A(in[814]), .B(n8573), .Z(n7120) );
  NAND U3304 ( .A(n6928), .B(n6794), .Z(n6795) );
  XNOR U3305 ( .A(n7120), .B(n6795), .Z(out[1433]) );
  XNOR U3306 ( .A(in[815]), .B(n8577), .Z(n7124) );
  NAND U3307 ( .A(n6930), .B(n6796), .Z(n6797) );
  XNOR U3308 ( .A(n7124), .B(n6797), .Z(out[1434]) );
  XNOR U3309 ( .A(in[816]), .B(n8581), .Z(n7128) );
  NAND U3310 ( .A(n6932), .B(n6798), .Z(n6799) );
  XNOR U3311 ( .A(n7128), .B(n6799), .Z(out[1435]) );
  XNOR U3312 ( .A(in[817]), .B(n8585), .Z(n7132) );
  NAND U3313 ( .A(n6936), .B(n6800), .Z(n6801) );
  XNOR U3314 ( .A(n7132), .B(n6801), .Z(out[1436]) );
  XNOR U3315 ( .A(in[818]), .B(n8589), .Z(n7136) );
  NAND U3316 ( .A(n6938), .B(n6802), .Z(n6803) );
  XNOR U3317 ( .A(n7136), .B(n6803), .Z(out[1437]) );
  XNOR U3318 ( .A(in[819]), .B(n8593), .Z(n7140) );
  NAND U3319 ( .A(n6940), .B(n6804), .Z(n6805) );
  XNOR U3320 ( .A(n7140), .B(n6805), .Z(out[1438]) );
  XNOR U3321 ( .A(in[820]), .B(n8597), .Z(n7144) );
  NAND U3322 ( .A(n6942), .B(n6806), .Z(n6807) );
  XNOR U3323 ( .A(n7144), .B(n6807), .Z(out[1439]) );
  XNOR U3324 ( .A(in[680]), .B(n8735), .Z(n7456) );
  XOR U3325 ( .A(in[614]), .B(n8587), .Z(n8882) );
  XOR U3326 ( .A(in[205]), .B(n8404), .Z(n8880) );
  NAND U3327 ( .A(n8882), .B(n8880), .Z(n6808) );
  XNOR U3328 ( .A(n7456), .B(n6808), .Z(out[143]) );
  XNOR U3329 ( .A(in[821]), .B(n8601), .Z(n7149) );
  NAND U3330 ( .A(n6944), .B(n6809), .Z(n6810) );
  XNOR U3331 ( .A(n7149), .B(n6810), .Z(out[1440]) );
  XNOR U3332 ( .A(in[822]), .B(n8611), .Z(n7153) );
  NAND U3333 ( .A(n6946), .B(n6811), .Z(n6812) );
  XNOR U3334 ( .A(n7153), .B(n6812), .Z(out[1441]) );
  XNOR U3335 ( .A(in[823]), .B(n8615), .Z(n7158) );
  NAND U3336 ( .A(n6948), .B(n6813), .Z(n6814) );
  XNOR U3337 ( .A(n7158), .B(n6814), .Z(out[1442]) );
  XNOR U3338 ( .A(in[824]), .B(n8619), .Z(n7162) );
  NAND U3339 ( .A(n6950), .B(n6815), .Z(n6816) );
  XNOR U3340 ( .A(n7162), .B(n6816), .Z(out[1443]) );
  XNOR U3341 ( .A(in[825]), .B(n8623), .Z(n7166) );
  NAND U3342 ( .A(n6952), .B(n6817), .Z(n6818) );
  XNOR U3343 ( .A(n7166), .B(n6818), .Z(out[1444]) );
  XNOR U3344 ( .A(in[826]), .B(n8345), .Z(n7170) );
  NAND U3345 ( .A(n6954), .B(n6819), .Z(n6820) );
  XNOR U3346 ( .A(n7170), .B(n6820), .Z(out[1445]) );
  XNOR U3347 ( .A(in[827]), .B(n8349), .Z(n7174) );
  NAND U3348 ( .A(n6957), .B(n6821), .Z(n6822) );
  XNOR U3349 ( .A(n7174), .B(n6822), .Z(out[1446]) );
  XNOR U3350 ( .A(in[828]), .B(n8353), .Z(n7178) );
  NAND U3351 ( .A(n6959), .B(n6823), .Z(n6824) );
  XNOR U3352 ( .A(n7178), .B(n6824), .Z(out[1447]) );
  XNOR U3353 ( .A(in[829]), .B(n8357), .Z(n7182) );
  NAND U3354 ( .A(n6961), .B(n6825), .Z(n6826) );
  XNOR U3355 ( .A(n7182), .B(n6826), .Z(out[1448]) );
  XNOR U3356 ( .A(in[830]), .B(n8361), .Z(n7186) );
  NAND U3357 ( .A(n6963), .B(n6827), .Z(n6828) );
  XNOR U3358 ( .A(n7186), .B(n6828), .Z(out[1449]) );
  XNOR U3359 ( .A(in[681]), .B(n8737), .Z(n7459) );
  XOR U3360 ( .A(in[615]), .B(n8591), .Z(n8920) );
  XOR U3361 ( .A(in[206]), .B(n8408), .Z(n8918) );
  NAND U3362 ( .A(n8920), .B(n8918), .Z(n6829) );
  XNOR U3363 ( .A(n7459), .B(n6829), .Z(out[144]) );
  XNOR U3364 ( .A(in[831]), .B(n8365), .Z(n7190) );
  NAND U3365 ( .A(n6965), .B(n6830), .Z(n6831) );
  XNOR U3366 ( .A(n7190), .B(n6831), .Z(out[1450]) );
  XNOR U3367 ( .A(in[768]), .B(n8369), .Z(n7194) );
  NAND U3368 ( .A(n6967), .B(n6832), .Z(n6833) );
  XNOR U3369 ( .A(n7194), .B(n6833), .Z(out[1451]) );
  XNOR U3370 ( .A(in[769]), .B(n8373), .Z(n7199) );
  NAND U3371 ( .A(n6969), .B(n6834), .Z(n6835) );
  XNOR U3372 ( .A(n7199), .B(n6835), .Z(out[1452]) );
  XOR U3373 ( .A(n8377), .B(in[770]), .Z(n7203) );
  NAND U3374 ( .A(n6971), .B(n6836), .Z(n6837) );
  XNOR U3375 ( .A(n7203), .B(n6837), .Z(out[1453]) );
  XOR U3376 ( .A(n8381), .B(in[771]), .Z(n7207) );
  NAND U3377 ( .A(n6973), .B(n6838), .Z(n6839) );
  XNOR U3378 ( .A(n7207), .B(n6839), .Z(out[1454]) );
  XOR U3379 ( .A(n8389), .B(in[772]), .Z(n7211) );
  NAND U3380 ( .A(n6975), .B(n6840), .Z(n6841) );
  XNOR U3381 ( .A(n7211), .B(n6841), .Z(out[1455]) );
  XOR U3382 ( .A(n8393), .B(in[773]), .Z(n7215) );
  NAND U3383 ( .A(n6978), .B(n6842), .Z(n6843) );
  XNOR U3384 ( .A(n7215), .B(n6843), .Z(out[1456]) );
  XOR U3385 ( .A(n8397), .B(in[774]), .Z(n7219) );
  NAND U3386 ( .A(n6980), .B(n6844), .Z(n6845) );
  XNOR U3387 ( .A(n7219), .B(n6845), .Z(out[1457]) );
  XOR U3388 ( .A(n8401), .B(in[775]), .Z(n7223) );
  NAND U3389 ( .A(n6982), .B(n6846), .Z(n6847) );
  XNOR U3390 ( .A(n7223), .B(n6847), .Z(out[1458]) );
  XOR U3391 ( .A(n8405), .B(in[776]), .Z(n7227) );
  NAND U3392 ( .A(n6984), .B(n6848), .Z(n6849) );
  XNOR U3393 ( .A(n7227), .B(n6849), .Z(out[1459]) );
  XNOR U3394 ( .A(in[682]), .B(n8739), .Z(n7462) );
  XOR U3395 ( .A(in[616]), .B(n8595), .Z(n8954) );
  XOR U3396 ( .A(in[207]), .B(n8412), .Z(n8952) );
  NAND U3397 ( .A(n8954), .B(n8952), .Z(n6850) );
  XNOR U3398 ( .A(n7462), .B(n6850), .Z(out[145]) );
  XOR U3399 ( .A(in[777]), .B(n8409), .Z(n7231) );
  NAND U3400 ( .A(n6986), .B(n6851), .Z(n6852) );
  XNOR U3401 ( .A(n7231), .B(n6852), .Z(out[1460]) );
  XOR U3402 ( .A(n8413), .B(in[778]), .Z(n7235) );
  NAND U3403 ( .A(n6988), .B(n6853), .Z(n6854) );
  XNOR U3404 ( .A(n7235), .B(n6854), .Z(out[1461]) );
  XOR U3405 ( .A(n8417), .B(in[779]), .Z(n7240) );
  NAND U3406 ( .A(n6990), .B(n6855), .Z(n6856) );
  XNOR U3407 ( .A(n7240), .B(n6856), .Z(out[1462]) );
  XOR U3408 ( .A(in[780]), .B(n8421), .Z(n7244) );
  NAND U3409 ( .A(n6992), .B(n6857), .Z(n6858) );
  XNOR U3410 ( .A(n7244), .B(n6858), .Z(out[1463]) );
  XOR U3411 ( .A(in[781]), .B(n8425), .Z(n7248) );
  NAND U3412 ( .A(n6994), .B(n6859), .Z(n6860) );
  XNOR U3413 ( .A(n7248), .B(n6860), .Z(out[1464]) );
  XOR U3414 ( .A(in[782]), .B(n8433), .Z(n7252) );
  NAND U3415 ( .A(n6996), .B(n6861), .Z(n6862) );
  XNOR U3416 ( .A(n7252), .B(n6862), .Z(out[1465]) );
  XOR U3417 ( .A(in[783]), .B(n8437), .Z(n7256) );
  NAND U3418 ( .A(n6999), .B(n6863), .Z(n6864) );
  XNOR U3419 ( .A(n7256), .B(n6864), .Z(out[1466]) );
  XOR U3420 ( .A(in[784]), .B(n8441), .Z(n7260) );
  NAND U3421 ( .A(n7001), .B(n6865), .Z(n6866) );
  XNOR U3422 ( .A(n7260), .B(n6866), .Z(out[1467]) );
  XOR U3423 ( .A(in[785]), .B(n8445), .Z(n7264) );
  NAND U3424 ( .A(n7003), .B(n6867), .Z(n6868) );
  XNOR U3425 ( .A(n7264), .B(n6868), .Z(out[1468]) );
  XOR U3426 ( .A(in[786]), .B(n8449), .Z(n7268) );
  NAND U3427 ( .A(n7005), .B(n6869), .Z(n6870) );
  XNOR U3428 ( .A(n7268), .B(n6870), .Z(out[1469]) );
  XNOR U3429 ( .A(in[683]), .B(n8741), .Z(n7465) );
  XOR U3430 ( .A(in[617]), .B(n8599), .Z(n8988) );
  XOR U3431 ( .A(in[208]), .B(n8416), .Z(n8986) );
  NAND U3432 ( .A(n8988), .B(n8986), .Z(n6871) );
  XNOR U3433 ( .A(n7465), .B(n6871), .Z(out[146]) );
  XOR U3434 ( .A(in[787]), .B(n8453), .Z(n7272) );
  NAND U3435 ( .A(n7007), .B(n6872), .Z(n6873) );
  XNOR U3436 ( .A(n7272), .B(n6873), .Z(out[1470]) );
  XOR U3437 ( .A(in[788]), .B(n8457), .Z(n7276) );
  NAND U3438 ( .A(n7009), .B(n6874), .Z(n6875) );
  XNOR U3439 ( .A(n7276), .B(n6875), .Z(out[1471]) );
  OR U3440 ( .A(n7012), .B(n6876), .Z(n6877) );
  XNOR U3441 ( .A(n7011), .B(n6877), .Z(out[1472]) );
  OR U3442 ( .A(n7017), .B(n6878), .Z(n6879) );
  XNOR U3443 ( .A(n7016), .B(n6879), .Z(out[1473]) );
  OR U3444 ( .A(n7022), .B(n6880), .Z(n6881) );
  XNOR U3445 ( .A(n7021), .B(n6881), .Z(out[1474]) );
  OR U3446 ( .A(n7026), .B(n6882), .Z(n6883) );
  XNOR U3447 ( .A(n7025), .B(n6883), .Z(out[1475]) );
  OR U3448 ( .A(n7032), .B(n6884), .Z(n6885) );
  XNOR U3449 ( .A(n7031), .B(n6885), .Z(out[1476]) );
  OR U3450 ( .A(n7036), .B(n6886), .Z(n6887) );
  XNOR U3451 ( .A(n7035), .B(n6887), .Z(out[1477]) );
  OR U3452 ( .A(n7040), .B(n6888), .Z(n6889) );
  XNOR U3453 ( .A(n7039), .B(n6889), .Z(out[1478]) );
  OR U3454 ( .A(n7044), .B(n6890), .Z(n6891) );
  XNOR U3455 ( .A(n7043), .B(n6891), .Z(out[1479]) );
  XNOR U3456 ( .A(in[684]), .B(n8743), .Z(n7468) );
  XOR U3457 ( .A(in[618]), .B(n8609), .Z(n9014) );
  XOR U3458 ( .A(in[209]), .B(n8420), .Z(n9012) );
  NAND U3459 ( .A(n9014), .B(n9012), .Z(n6892) );
  XNOR U3460 ( .A(n7468), .B(n6892), .Z(out[147]) );
  OR U3461 ( .A(n7049), .B(n6893), .Z(n6894) );
  XNOR U3462 ( .A(n7048), .B(n6894), .Z(out[1480]) );
  OR U3463 ( .A(n7053), .B(n6895), .Z(n6896) );
  XNOR U3464 ( .A(n7052), .B(n6896), .Z(out[1481]) );
  OR U3465 ( .A(n7057), .B(n6897), .Z(n6898) );
  XNOR U3466 ( .A(n7056), .B(n6898), .Z(out[1482]) );
  OR U3467 ( .A(n7061), .B(n6899), .Z(n6900) );
  XNOR U3468 ( .A(n7060), .B(n6900), .Z(out[1483]) );
  OR U3469 ( .A(n7065), .B(n6901), .Z(n6902) );
  XNOR U3470 ( .A(n7064), .B(n6902), .Z(out[1484]) );
  OR U3471 ( .A(n7069), .B(n6903), .Z(n6904) );
  XNOR U3472 ( .A(n7068), .B(n6904), .Z(out[1485]) );
  OR U3473 ( .A(n7074), .B(n6905), .Z(n6906) );
  XNOR U3474 ( .A(n7073), .B(n6906), .Z(out[1486]) );
  OR U3475 ( .A(n7078), .B(n6907), .Z(n6908) );
  XNOR U3476 ( .A(n7077), .B(n6908), .Z(out[1487]) );
  OR U3477 ( .A(n7083), .B(n6909), .Z(n6910) );
  XNOR U3478 ( .A(n7082), .B(n6910), .Z(out[1488]) );
  OR U3479 ( .A(n7087), .B(n6911), .Z(n6912) );
  XNOR U3480 ( .A(n7086), .B(n6912), .Z(out[1489]) );
  XNOR U3481 ( .A(in[685]), .B(n8745), .Z(n7471) );
  XOR U3482 ( .A(in[619]), .B(n8613), .Z(n9038) );
  XOR U3483 ( .A(in[210]), .B(n8424), .Z(n9036) );
  NAND U3484 ( .A(n9038), .B(n9036), .Z(n6913) );
  XNOR U3485 ( .A(n7471), .B(n6913), .Z(out[148]) );
  OR U3486 ( .A(n7091), .B(n6914), .Z(n6915) );
  XNOR U3487 ( .A(n7090), .B(n6915), .Z(out[1490]) );
  OR U3488 ( .A(n7095), .B(n6916), .Z(n6917) );
  XNOR U3489 ( .A(n7094), .B(n6917), .Z(out[1491]) );
  OR U3490 ( .A(n7099), .B(n6918), .Z(n6919) );
  XNOR U3491 ( .A(n7098), .B(n6919), .Z(out[1492]) );
  OR U3492 ( .A(n7103), .B(n6920), .Z(n6921) );
  XNOR U3493 ( .A(n7102), .B(n6921), .Z(out[1493]) );
  OR U3494 ( .A(n7107), .B(n6922), .Z(n6923) );
  XNOR U3495 ( .A(n7106), .B(n6923), .Z(out[1494]) );
  OR U3496 ( .A(n7111), .B(n6924), .Z(n6925) );
  XNOR U3497 ( .A(n7110), .B(n6925), .Z(out[1495]) );
  OR U3498 ( .A(n7116), .B(n6926), .Z(n6927) );
  XNOR U3499 ( .A(n7115), .B(n6927), .Z(out[1496]) );
  OR U3500 ( .A(n7120), .B(n6928), .Z(n6929) );
  XNOR U3501 ( .A(n7119), .B(n6929), .Z(out[1497]) );
  OR U3502 ( .A(n7124), .B(n6930), .Z(n6931) );
  XNOR U3503 ( .A(n7123), .B(n6931), .Z(out[1498]) );
  OR U3504 ( .A(n7128), .B(n6932), .Z(n6933) );
  XNOR U3505 ( .A(n7127), .B(n6933), .Z(out[1499]) );
  XNOR U3506 ( .A(in[686]), .B(n8747), .Z(n7473) );
  XOR U3507 ( .A(in[620]), .B(n8617), .Z(n9062) );
  XNOR U3508 ( .A(in[211]), .B(n8432), .Z(n9060) );
  NAND U3509 ( .A(n9062), .B(n9060), .Z(n6934) );
  XNOR U3510 ( .A(n7473), .B(n6934), .Z(out[149]) );
  XNOR U3511 ( .A(in[1424]), .B(n8441), .Z(n8845) );
  XOR U3512 ( .A(in[1047]), .B(n8939), .Z(n7452) );
  NAND U3513 ( .A(n8845), .B(n7452), .Z(n6935) );
  XNOR U3514 ( .A(n8846), .B(n6935), .Z(out[14]) );
  OR U3515 ( .A(n7132), .B(n6936), .Z(n6937) );
  XNOR U3516 ( .A(n7131), .B(n6937), .Z(out[1500]) );
  OR U3517 ( .A(n7136), .B(n6938), .Z(n6939) );
  XNOR U3518 ( .A(n7135), .B(n6939), .Z(out[1501]) );
  OR U3519 ( .A(n7140), .B(n6940), .Z(n6941) );
  XNOR U3520 ( .A(n7139), .B(n6941), .Z(out[1502]) );
  OR U3521 ( .A(n7144), .B(n6942), .Z(n6943) );
  XNOR U3522 ( .A(n7143), .B(n6943), .Z(out[1503]) );
  OR U3523 ( .A(n7149), .B(n6944), .Z(n6945) );
  XNOR U3524 ( .A(n7148), .B(n6945), .Z(out[1504]) );
  OR U3525 ( .A(n7153), .B(n6946), .Z(n6947) );
  XNOR U3526 ( .A(n7152), .B(n6947), .Z(out[1505]) );
  OR U3527 ( .A(n7158), .B(n6948), .Z(n6949) );
  XNOR U3528 ( .A(n7157), .B(n6949), .Z(out[1506]) );
  OR U3529 ( .A(n7162), .B(n6950), .Z(n6951) );
  XNOR U3530 ( .A(n7161), .B(n6951), .Z(out[1507]) );
  OR U3531 ( .A(n7166), .B(n6952), .Z(n6953) );
  XNOR U3532 ( .A(n7165), .B(n6953), .Z(out[1508]) );
  OR U3533 ( .A(n7170), .B(n6954), .Z(n6955) );
  XNOR U3534 ( .A(n7169), .B(n6955), .Z(out[1509]) );
  XNOR U3535 ( .A(in[687]), .B(n8749), .Z(n7476) );
  XOR U3536 ( .A(in[621]), .B(n8621), .Z(n9086) );
  XNOR U3537 ( .A(in[212]), .B(n8436), .Z(n9084) );
  NAND U3538 ( .A(n9086), .B(n9084), .Z(n6956) );
  XNOR U3539 ( .A(n7476), .B(n6956), .Z(out[150]) );
  OR U3540 ( .A(n7174), .B(n6957), .Z(n6958) );
  XNOR U3541 ( .A(n7173), .B(n6958), .Z(out[1510]) );
  OR U3542 ( .A(n7178), .B(n6959), .Z(n6960) );
  XNOR U3543 ( .A(n7177), .B(n6960), .Z(out[1511]) );
  OR U3544 ( .A(n7182), .B(n6961), .Z(n6962) );
  XNOR U3545 ( .A(n7181), .B(n6962), .Z(out[1512]) );
  OR U3546 ( .A(n7186), .B(n6963), .Z(n6964) );
  XNOR U3547 ( .A(n7185), .B(n6964), .Z(out[1513]) );
  OR U3548 ( .A(n7190), .B(n6965), .Z(n6966) );
  XNOR U3549 ( .A(n7189), .B(n6966), .Z(out[1514]) );
  OR U3550 ( .A(n7194), .B(n6967), .Z(n6968) );
  XNOR U3551 ( .A(n7193), .B(n6968), .Z(out[1515]) );
  OR U3552 ( .A(n7199), .B(n6969), .Z(n6970) );
  XNOR U3553 ( .A(n7198), .B(n6970), .Z(out[1516]) );
  OR U3554 ( .A(n7203), .B(n6971), .Z(n6972) );
  XNOR U3555 ( .A(n7202), .B(n6972), .Z(out[1517]) );
  OR U3556 ( .A(n7207), .B(n6973), .Z(n6974) );
  XNOR U3557 ( .A(n7206), .B(n6974), .Z(out[1518]) );
  OR U3558 ( .A(n7211), .B(n6975), .Z(n6976) );
  XNOR U3559 ( .A(n7210), .B(n6976), .Z(out[1519]) );
  XNOR U3560 ( .A(in[688]), .B(n8755), .Z(n7479) );
  XOR U3561 ( .A(in[622]), .B(n8343), .Z(n9110) );
  XNOR U3562 ( .A(in[213]), .B(n8440), .Z(n9108) );
  NAND U3563 ( .A(n9110), .B(n9108), .Z(n6977) );
  XNOR U3564 ( .A(n7479), .B(n6977), .Z(out[151]) );
  OR U3565 ( .A(n7215), .B(n6978), .Z(n6979) );
  XNOR U3566 ( .A(n7214), .B(n6979), .Z(out[1520]) );
  OR U3567 ( .A(n7219), .B(n6980), .Z(n6981) );
  XNOR U3568 ( .A(n7218), .B(n6981), .Z(out[1521]) );
  OR U3569 ( .A(n7223), .B(n6982), .Z(n6983) );
  XNOR U3570 ( .A(n7222), .B(n6983), .Z(out[1522]) );
  OR U3571 ( .A(n7227), .B(n6984), .Z(n6985) );
  XNOR U3572 ( .A(n7226), .B(n6985), .Z(out[1523]) );
  OR U3573 ( .A(n7231), .B(n6986), .Z(n6987) );
  XNOR U3574 ( .A(n7230), .B(n6987), .Z(out[1524]) );
  OR U3575 ( .A(n7235), .B(n6988), .Z(n6989) );
  XNOR U3576 ( .A(n7234), .B(n6989), .Z(out[1525]) );
  OR U3577 ( .A(n7240), .B(n6990), .Z(n6991) );
  XNOR U3578 ( .A(n7239), .B(n6991), .Z(out[1526]) );
  OR U3579 ( .A(n7244), .B(n6992), .Z(n6993) );
  XNOR U3580 ( .A(n7243), .B(n6993), .Z(out[1527]) );
  OR U3581 ( .A(n7248), .B(n6994), .Z(n6995) );
  XNOR U3582 ( .A(n7247), .B(n6995), .Z(out[1528]) );
  OR U3583 ( .A(n7252), .B(n6996), .Z(n6997) );
  XNOR U3584 ( .A(n7251), .B(n6997), .Z(out[1529]) );
  XNOR U3585 ( .A(in[689]), .B(n8757), .Z(n7483) );
  XOR U3586 ( .A(in[623]), .B(n8347), .Z(n9134) );
  XNOR U3587 ( .A(in[214]), .B(n8444), .Z(n9132) );
  NAND U3588 ( .A(n9134), .B(n9132), .Z(n6998) );
  XNOR U3589 ( .A(n7483), .B(n6998), .Z(out[152]) );
  OR U3590 ( .A(n7256), .B(n6999), .Z(n7000) );
  XNOR U3591 ( .A(n7255), .B(n7000), .Z(out[1530]) );
  OR U3592 ( .A(n7260), .B(n7001), .Z(n7002) );
  XNOR U3593 ( .A(n7259), .B(n7002), .Z(out[1531]) );
  OR U3594 ( .A(n7264), .B(n7003), .Z(n7004) );
  XNOR U3595 ( .A(n7263), .B(n7004), .Z(out[1532]) );
  OR U3596 ( .A(n7268), .B(n7005), .Z(n7006) );
  XNOR U3597 ( .A(n7267), .B(n7006), .Z(out[1533]) );
  OR U3598 ( .A(n7272), .B(n7007), .Z(n7008) );
  XNOR U3599 ( .A(n7271), .B(n7008), .Z(out[1534]) );
  OR U3600 ( .A(n7276), .B(n7009), .Z(n7010) );
  XNOR U3601 ( .A(n7275), .B(n7010), .Z(out[1535]) );
  ANDN U3602 ( .B(n7012), .A(n7011), .Z(n7015) );
  XOR U3603 ( .A(n7013), .B(round_const[0]), .Z(n7014) );
  XNOR U3604 ( .A(n7015), .B(n7014), .Z(out[1536]) );
  ANDN U3605 ( .B(n7017), .A(n7016), .Z(n7020) );
  XOR U3606 ( .A(n7018), .B(round_const[1]), .Z(n7019) );
  XNOR U3607 ( .A(n7020), .B(n7019), .Z(out[1537]) );
  ANDN U3608 ( .B(n7022), .A(n7021), .Z(n7023) );
  XNOR U3609 ( .A(n7024), .B(n7023), .Z(out[1538]) );
  ANDN U3610 ( .B(n7026), .A(n7025), .Z(n7029) );
  XOR U3611 ( .A(n7027), .B(round_const_3), .Z(n7028) );
  XNOR U3612 ( .A(n7029), .B(n7028), .Z(out[1539]) );
  XNOR U3613 ( .A(in[690]), .B(n8759), .Z(n7486) );
  XOR U3614 ( .A(in[624]), .B(n8351), .Z(n9166) );
  XNOR U3615 ( .A(in[215]), .B(n8448), .Z(n9164) );
  NAND U3616 ( .A(n9166), .B(n9164), .Z(n7030) );
  XNOR U3617 ( .A(n7486), .B(n7030), .Z(out[153]) );
  ANDN U3618 ( .B(n7032), .A(n7031), .Z(n7033) );
  XNOR U3619 ( .A(n7034), .B(n7033), .Z(out[1540]) );
  ANDN U3620 ( .B(n7036), .A(n7035), .Z(n7037) );
  XNOR U3621 ( .A(n7038), .B(n7037), .Z(out[1541]) );
  ANDN U3622 ( .B(n7040), .A(n7039), .Z(n7041) );
  XNOR U3623 ( .A(n7042), .B(n7041), .Z(out[1542]) );
  ANDN U3624 ( .B(n7044), .A(n7043), .Z(n7047) );
  XOR U3625 ( .A(n7045), .B(round_const_7), .Z(n7046) );
  XNOR U3626 ( .A(n7047), .B(n7046), .Z(out[1543]) );
  ANDN U3627 ( .B(n7049), .A(n7048), .Z(n7050) );
  XNOR U3628 ( .A(n7051), .B(n7050), .Z(out[1544]) );
  ANDN U3629 ( .B(n7053), .A(n7052), .Z(n7054) );
  XNOR U3630 ( .A(n7055), .B(n7054), .Z(out[1545]) );
  ANDN U3631 ( .B(n7057), .A(n7056), .Z(n7058) );
  XNOR U3632 ( .A(n7059), .B(n7058), .Z(out[1546]) );
  ANDN U3633 ( .B(n7061), .A(n7060), .Z(n7062) );
  XNOR U3634 ( .A(n7063), .B(n7062), .Z(out[1547]) );
  ANDN U3635 ( .B(n7065), .A(n7064), .Z(n7066) );
  XNOR U3636 ( .A(n7067), .B(n7066), .Z(out[1548]) );
  ANDN U3637 ( .B(n7069), .A(n7068), .Z(n7070) );
  XNOR U3638 ( .A(n7071), .B(n7070), .Z(out[1549]) );
  XNOR U3639 ( .A(in[691]), .B(n8761), .Z(n7489) );
  XOR U3640 ( .A(in[625]), .B(n8355), .Z(n9214) );
  XNOR U3641 ( .A(in[216]), .B(n8452), .Z(n9212) );
  NAND U3642 ( .A(n9214), .B(n9212), .Z(n7072) );
  XNOR U3643 ( .A(n7489), .B(n7072), .Z(out[154]) );
  ANDN U3644 ( .B(n7074), .A(n7073), .Z(n7075) );
  XNOR U3645 ( .A(n7076), .B(n7075), .Z(out[1550]) );
  ANDN U3646 ( .B(n7078), .A(n7077), .Z(n7081) );
  XOR U3647 ( .A(n7079), .B(round_const_15), .Z(n7080) );
  XNOR U3648 ( .A(n7081), .B(n7080), .Z(out[1551]) );
  ANDN U3649 ( .B(n7083), .A(n7082), .Z(n7084) );
  XNOR U3650 ( .A(n7085), .B(n7084), .Z(out[1552]) );
  ANDN U3651 ( .B(n7087), .A(n7086), .Z(n7088) );
  XNOR U3652 ( .A(n7089), .B(n7088), .Z(out[1553]) );
  ANDN U3653 ( .B(n7091), .A(n7090), .Z(n7092) );
  XNOR U3654 ( .A(n7093), .B(n7092), .Z(out[1554]) );
  ANDN U3655 ( .B(n7095), .A(n7094), .Z(n7096) );
  XNOR U3656 ( .A(n7097), .B(n7096), .Z(out[1555]) );
  ANDN U3657 ( .B(n7099), .A(n7098), .Z(n7100) );
  XNOR U3658 ( .A(n7101), .B(n7100), .Z(out[1556]) );
  ANDN U3659 ( .B(n7103), .A(n7102), .Z(n7104) );
  XNOR U3660 ( .A(n7105), .B(n7104), .Z(out[1557]) );
  ANDN U3661 ( .B(n7107), .A(n7106), .Z(n7108) );
  XNOR U3662 ( .A(n7109), .B(n7108), .Z(out[1558]) );
  ANDN U3663 ( .B(n7111), .A(n7110), .Z(n7112) );
  XNOR U3664 ( .A(n7113), .B(n7112), .Z(out[1559]) );
  XNOR U3665 ( .A(in[692]), .B(n8763), .Z(n7492) );
  XOR U3666 ( .A(in[626]), .B(n8359), .Z(n9258) );
  XNOR U3667 ( .A(in[217]), .B(n8456), .Z(n9256) );
  NAND U3668 ( .A(n9258), .B(n9256), .Z(n7114) );
  XNOR U3669 ( .A(n7492), .B(n7114), .Z(out[155]) );
  ANDN U3670 ( .B(n7116), .A(n7115), .Z(n7117) );
  XNOR U3671 ( .A(n7118), .B(n7117), .Z(out[1560]) );
  ANDN U3672 ( .B(n7120), .A(n7119), .Z(n7121) );
  XNOR U3673 ( .A(n7122), .B(n7121), .Z(out[1561]) );
  ANDN U3674 ( .B(n7124), .A(n7123), .Z(n7125) );
  XNOR U3675 ( .A(n7126), .B(n7125), .Z(out[1562]) );
  ANDN U3676 ( .B(n7128), .A(n7127), .Z(n7129) );
  XNOR U3677 ( .A(n7130), .B(n7129), .Z(out[1563]) );
  ANDN U3678 ( .B(n7132), .A(n7131), .Z(n7133) );
  XNOR U3679 ( .A(n7134), .B(n7133), .Z(out[1564]) );
  ANDN U3680 ( .B(n7136), .A(n7135), .Z(n7137) );
  XNOR U3681 ( .A(n7138), .B(n7137), .Z(out[1565]) );
  ANDN U3682 ( .B(n7140), .A(n7139), .Z(n7141) );
  XNOR U3683 ( .A(n7142), .B(n7141), .Z(out[1566]) );
  ANDN U3684 ( .B(n7144), .A(n7143), .Z(n7147) );
  XOR U3685 ( .A(n7145), .B(round_const_31), .Z(n7146) );
  XNOR U3686 ( .A(n7147), .B(n7146), .Z(out[1567]) );
  ANDN U3687 ( .B(n7149), .A(n7148), .Z(n7150) );
  XNOR U3688 ( .A(n7151), .B(n7150), .Z(out[1568]) );
  ANDN U3689 ( .B(n7153), .A(n7152), .Z(n7154) );
  XNOR U3690 ( .A(n7155), .B(n7154), .Z(out[1569]) );
  XNOR U3691 ( .A(in[693]), .B(n8765), .Z(n7495) );
  XOR U3692 ( .A(in[627]), .B(n8363), .Z(n9302) );
  XNOR U3693 ( .A(in[218]), .B(n8460), .Z(n9299) );
  NAND U3694 ( .A(n9302), .B(n9299), .Z(n7156) );
  XNOR U3695 ( .A(n7495), .B(n7156), .Z(out[156]) );
  ANDN U3696 ( .B(n7158), .A(n7157), .Z(n7159) );
  XNOR U3697 ( .A(n7160), .B(n7159), .Z(out[1570]) );
  ANDN U3698 ( .B(n7162), .A(n7161), .Z(n7163) );
  XNOR U3699 ( .A(n7164), .B(n7163), .Z(out[1571]) );
  ANDN U3700 ( .B(n7166), .A(n7165), .Z(n7167) );
  XNOR U3701 ( .A(n7168), .B(n7167), .Z(out[1572]) );
  ANDN U3702 ( .B(n7170), .A(n7169), .Z(n7171) );
  XNOR U3703 ( .A(n7172), .B(n7171), .Z(out[1573]) );
  ANDN U3704 ( .B(n7174), .A(n7173), .Z(n7175) );
  XNOR U3705 ( .A(n7176), .B(n7175), .Z(out[1574]) );
  ANDN U3706 ( .B(n7178), .A(n7177), .Z(n7179) );
  XNOR U3707 ( .A(n7180), .B(n7179), .Z(out[1575]) );
  ANDN U3708 ( .B(n7182), .A(n7181), .Z(n7183) );
  XNOR U3709 ( .A(n7184), .B(n7183), .Z(out[1576]) );
  ANDN U3710 ( .B(n7186), .A(n7185), .Z(n7187) );
  XNOR U3711 ( .A(n7188), .B(n7187), .Z(out[1577]) );
  ANDN U3712 ( .B(n7190), .A(n7189), .Z(n7191) );
  XNOR U3713 ( .A(n7192), .B(n7191), .Z(out[1578]) );
  ANDN U3714 ( .B(n7194), .A(n7193), .Z(n7195) );
  XNOR U3715 ( .A(n7196), .B(n7195), .Z(out[1579]) );
  XNOR U3716 ( .A(in[694]), .B(n8767), .Z(n7497) );
  XOR U3717 ( .A(in[628]), .B(n8367), .Z(n9346) );
  XNOR U3718 ( .A(in[219]), .B(n8464), .Z(n9343) );
  NAND U3719 ( .A(n9346), .B(n9343), .Z(n7197) );
  XNOR U3720 ( .A(n7497), .B(n7197), .Z(out[157]) );
  ANDN U3721 ( .B(n7199), .A(n7198), .Z(n7200) );
  XNOR U3722 ( .A(n7201), .B(n7200), .Z(out[1580]) );
  ANDN U3723 ( .B(n7203), .A(n7202), .Z(n7204) );
  XNOR U3724 ( .A(n7205), .B(n7204), .Z(out[1581]) );
  ANDN U3725 ( .B(n7207), .A(n7206), .Z(n7208) );
  XNOR U3726 ( .A(n7209), .B(n7208), .Z(out[1582]) );
  ANDN U3727 ( .B(n7211), .A(n7210), .Z(n7212) );
  XNOR U3728 ( .A(n7213), .B(n7212), .Z(out[1583]) );
  ANDN U3729 ( .B(n7215), .A(n7214), .Z(n7216) );
  XNOR U3730 ( .A(n7217), .B(n7216), .Z(out[1584]) );
  ANDN U3731 ( .B(n7219), .A(n7218), .Z(n7220) );
  XNOR U3732 ( .A(n7221), .B(n7220), .Z(out[1585]) );
  ANDN U3733 ( .B(n7223), .A(n7222), .Z(n7224) );
  XNOR U3734 ( .A(n7225), .B(n7224), .Z(out[1586]) );
  ANDN U3735 ( .B(n7227), .A(n7226), .Z(n7228) );
  XNOR U3736 ( .A(n7229), .B(n7228), .Z(out[1587]) );
  ANDN U3737 ( .B(n7231), .A(n7230), .Z(n7232) );
  XNOR U3738 ( .A(n7233), .B(n7232), .Z(out[1588]) );
  ANDN U3739 ( .B(n7235), .A(n7234), .Z(n7236) );
  XNOR U3740 ( .A(n7237), .B(n7236), .Z(out[1589]) );
  XNOR U3741 ( .A(in[695]), .B(n8769), .Z(n7499) );
  XOR U3742 ( .A(in[629]), .B(n8371), .Z(n9390) );
  XNOR U3743 ( .A(in[220]), .B(n8468), .Z(n9387) );
  NAND U3744 ( .A(n9390), .B(n9387), .Z(n7238) );
  XNOR U3745 ( .A(n7499), .B(n7238), .Z(out[158]) );
  ANDN U3746 ( .B(n7240), .A(n7239), .Z(n7241) );
  XNOR U3747 ( .A(n7242), .B(n7241), .Z(out[1590]) );
  ANDN U3748 ( .B(n7244), .A(n7243), .Z(n7245) );
  XNOR U3749 ( .A(n7246), .B(n7245), .Z(out[1591]) );
  ANDN U3750 ( .B(n7248), .A(n7247), .Z(n7249) );
  XNOR U3751 ( .A(n7250), .B(n7249), .Z(out[1592]) );
  ANDN U3752 ( .B(n7252), .A(n7251), .Z(n7253) );
  XNOR U3753 ( .A(n7254), .B(n7253), .Z(out[1593]) );
  ANDN U3754 ( .B(n7256), .A(n7255), .Z(n7257) );
  XNOR U3755 ( .A(n7258), .B(n7257), .Z(out[1594]) );
  ANDN U3756 ( .B(n7260), .A(n7259), .Z(n7261) );
  XNOR U3757 ( .A(n7262), .B(n7261), .Z(out[1595]) );
  ANDN U3758 ( .B(n7264), .A(n7263), .Z(n7265) );
  XNOR U3759 ( .A(n7266), .B(n7265), .Z(out[1596]) );
  ANDN U3760 ( .B(n7268), .A(n7267), .Z(n7269) );
  XNOR U3761 ( .A(n7270), .B(n7269), .Z(out[1597]) );
  ANDN U3762 ( .B(n7272), .A(n7271), .Z(n7273) );
  XNOR U3763 ( .A(n7274), .B(n7273), .Z(out[1598]) );
  ANDN U3764 ( .B(n7276), .A(n7275), .Z(n7279) );
  XOR U3765 ( .A(n7277), .B(round_const_63), .Z(n7278) );
  XNOR U3766 ( .A(n7279), .B(n7278), .Z(out[1599]) );
  XNOR U3767 ( .A(in[696]), .B(n8625), .Z(n7501) );
  XOR U3768 ( .A(in[630]), .B(n8375), .Z(n9434) );
  XNOR U3769 ( .A(in[221]), .B(n8476), .Z(n9431) );
  NAND U3770 ( .A(n9434), .B(n9431), .Z(n7280) );
  XNOR U3771 ( .A(n7501), .B(n7280), .Z(out[159]) );
  XNOR U3772 ( .A(in[1425]), .B(n8445), .Z(n8879) );
  XOR U3773 ( .A(in[1048]), .B(n8942), .Z(n7455) );
  NAND U3774 ( .A(n8879), .B(n7455), .Z(n7281) );
  XNOR U3775 ( .A(n8880), .B(n7281), .Z(out[15]) );
  XNOR U3776 ( .A(in[697]), .B(n8627), .Z(n7503) );
  XOR U3777 ( .A(in[631]), .B(n8379), .Z(n9478) );
  XNOR U3778 ( .A(in[222]), .B(n8480), .Z(n9475) );
  NAND U3779 ( .A(n9478), .B(n9475), .Z(n7282) );
  XNOR U3780 ( .A(n7503), .B(n7282), .Z(out[160]) );
  XNOR U3781 ( .A(in[698]), .B(n8629), .Z(n7505) );
  XOR U3782 ( .A(in[632]), .B(n8387), .Z(n9522) );
  XNOR U3783 ( .A(in[223]), .B(n8484), .Z(n9519) );
  NAND U3784 ( .A(n9522), .B(n9519), .Z(n7283) );
  XNOR U3785 ( .A(n7505), .B(n7283), .Z(out[161]) );
  XNOR U3786 ( .A(in[699]), .B(n8631), .Z(n7509) );
  XOR U3787 ( .A(in[633]), .B(n8391), .Z(n9566) );
  XNOR U3788 ( .A(in[224]), .B(n8488), .Z(n9563) );
  NAND U3789 ( .A(n9566), .B(n9563), .Z(n7284) );
  XNOR U3790 ( .A(n7509), .B(n7284), .Z(out[162]) );
  XNOR U3791 ( .A(in[700]), .B(n8633), .Z(n7511) );
  XOR U3792 ( .A(in[634]), .B(n8395), .Z(n9610) );
  XNOR U3793 ( .A(in[225]), .B(n8492), .Z(n9607) );
  NAND U3794 ( .A(n9610), .B(n9607), .Z(n7285) );
  XNOR U3795 ( .A(n7511), .B(n7285), .Z(out[163]) );
  XOR U3796 ( .A(in[701]), .B(n8635), .Z(n7513) );
  NOR U3797 ( .A(n7357), .B(n7638), .Z(n7286) );
  XNOR U3798 ( .A(n7513), .B(n7286), .Z(out[164]) );
  XOR U3799 ( .A(in[702]), .B(n8641), .Z(n7515) );
  NOR U3800 ( .A(n7359), .B(n7652), .Z(n7287) );
  XNOR U3801 ( .A(n7515), .B(n7287), .Z(out[165]) );
  XOR U3802 ( .A(in[703]), .B(n8643), .Z(n7517) );
  NOR U3803 ( .A(n7362), .B(n7666), .Z(n7288) );
  XNOR U3804 ( .A(n7517), .B(n7288), .Z(out[166]) );
  XOR U3805 ( .A(in[640]), .B(n8645), .Z(n7519) );
  NOR U3806 ( .A(n7364), .B(n7680), .Z(n7289) );
  XNOR U3807 ( .A(n7519), .B(n7289), .Z(out[167]) );
  XOR U3808 ( .A(in[641]), .B(n8647), .Z(n7521) );
  NOR U3809 ( .A(n7366), .B(n7696), .Z(n7290) );
  XNOR U3810 ( .A(n7521), .B(n7290), .Z(out[168]) );
  XOR U3811 ( .A(in[642]), .B(n8649), .Z(n7523) );
  NOR U3812 ( .A(n7368), .B(n7710), .Z(n7291) );
  XNOR U3813 ( .A(n7523), .B(n7291), .Z(out[169]) );
  XNOR U3814 ( .A(in[1426]), .B(n8449), .Z(n8917) );
  XOR U3815 ( .A(in[1049]), .B(n8945), .Z(n7458) );
  NAND U3816 ( .A(n8917), .B(n7458), .Z(n7292) );
  XNOR U3817 ( .A(n8918), .B(n7292), .Z(out[16]) );
  XOR U3818 ( .A(in[643]), .B(n8651), .Z(n7525) );
  NOR U3819 ( .A(n7370), .B(n7724), .Z(n7293) );
  XNOR U3820 ( .A(n7525), .B(n7293), .Z(out[170]) );
  XOR U3821 ( .A(in[644]), .B(n8653), .Z(n7527) );
  NOR U3822 ( .A(n7372), .B(n7738), .Z(n7294) );
  XNOR U3823 ( .A(n7527), .B(n7294), .Z(out[171]) );
  XOR U3824 ( .A(in[645]), .B(n8655), .Z(n7533) );
  NOR U3825 ( .A(n7374), .B(n7754), .Z(n7295) );
  XNOR U3826 ( .A(n7533), .B(n7295), .Z(out[172]) );
  XOR U3827 ( .A(in[646]), .B(n8657), .Z(n7535) );
  NOR U3828 ( .A(n7376), .B(n7778), .Z(n7296) );
  XNOR U3829 ( .A(n7535), .B(n7296), .Z(out[173]) );
  XOR U3830 ( .A(in[647]), .B(n8659), .Z(n7537) );
  NOR U3831 ( .A(n7378), .B(n7802), .Z(n7297) );
  XNOR U3832 ( .A(n7537), .B(n7297), .Z(out[174]) );
  XOR U3833 ( .A(in[648]), .B(n8663), .Z(n7539) );
  NOR U3834 ( .A(n7380), .B(n7826), .Z(n7298) );
  XNOR U3835 ( .A(n7539), .B(n7298), .Z(out[175]) );
  XOR U3836 ( .A(in[649]), .B(n8665), .Z(n7541) );
  NOR U3837 ( .A(n7383), .B(n7850), .Z(n7299) );
  XNOR U3838 ( .A(n7541), .B(n7299), .Z(out[176]) );
  XOR U3839 ( .A(in[650]), .B(n8667), .Z(n7543) );
  NOR U3840 ( .A(n7385), .B(n7874), .Z(n7300) );
  XNOR U3841 ( .A(n7543), .B(n7300), .Z(out[177]) );
  XOR U3842 ( .A(in[651]), .B(n8669), .Z(n7545) );
  NOR U3843 ( .A(n7387), .B(n7900), .Z(n7301) );
  XNOR U3844 ( .A(n7545), .B(n7301), .Z(out[178]) );
  XOR U3845 ( .A(in[652]), .B(n8671), .Z(n7547) );
  NOR U3846 ( .A(n7389), .B(n7924), .Z(n7302) );
  XNOR U3847 ( .A(n7547), .B(n7302), .Z(out[179]) );
  XNOR U3848 ( .A(in[1427]), .B(n8453), .Z(n8951) );
  XOR U3849 ( .A(in[1050]), .B(n8948), .Z(n7461) );
  NAND U3850 ( .A(n8951), .B(n7461), .Z(n7303) );
  XNOR U3851 ( .A(n8952), .B(n7303), .Z(out[17]) );
  XOR U3852 ( .A(in[653]), .B(n8673), .Z(n7549) );
  NOR U3853 ( .A(n7391), .B(n7948), .Z(n7304) );
  XNOR U3854 ( .A(n7549), .B(n7304), .Z(out[180]) );
  XOR U3855 ( .A(in[654]), .B(n8675), .Z(n7551) );
  NOR U3856 ( .A(n7393), .B(n7972), .Z(n7305) );
  XNOR U3857 ( .A(n7551), .B(n7305), .Z(out[181]) );
  XOR U3858 ( .A(in[655]), .B(n8677), .Z(n7555) );
  NOR U3859 ( .A(n7395), .B(n7996), .Z(n7306) );
  XNOR U3860 ( .A(n7555), .B(n7306), .Z(out[182]) );
  XOR U3861 ( .A(in[656]), .B(n8679), .Z(n7557) );
  NOR U3862 ( .A(n7397), .B(n8020), .Z(n7307) );
  XNOR U3863 ( .A(n7557), .B(n7307), .Z(out[183]) );
  XOR U3864 ( .A(in[657]), .B(n8681), .Z(n7559) );
  NOR U3865 ( .A(n7399), .B(n8044), .Z(n7308) );
  XNOR U3866 ( .A(n7559), .B(n7308), .Z(out[184]) );
  XOR U3867 ( .A(in[658]), .B(n8685), .Z(n7561) );
  NOR U3868 ( .A(n7401), .B(n8076), .Z(n7309) );
  XNOR U3869 ( .A(n7561), .B(n7309), .Z(out[185]) );
  XOR U3870 ( .A(in[659]), .B(n8687), .Z(n7563) );
  NOR U3871 ( .A(n7404), .B(n8120), .Z(n7310) );
  XNOR U3872 ( .A(n7563), .B(n7310), .Z(out[186]) );
  XOR U3873 ( .A(in[660]), .B(n8689), .Z(n7565) );
  NOR U3874 ( .A(n7406), .B(n8164), .Z(n7311) );
  XNOR U3875 ( .A(n7565), .B(n7311), .Z(out[187]) );
  XOR U3876 ( .A(in[661]), .B(n8691), .Z(n7567) );
  NOR U3877 ( .A(n7408), .B(n8210), .Z(n7312) );
  XNOR U3878 ( .A(n7567), .B(n7312), .Z(out[188]) );
  XOR U3879 ( .A(in[662]), .B(n8693), .Z(n7569) );
  NOR U3880 ( .A(n7410), .B(n8254), .Z(n7313) );
  XNOR U3881 ( .A(n7569), .B(n7313), .Z(out[189]) );
  XNOR U3882 ( .A(in[1428]), .B(n8457), .Z(n8985) );
  XOR U3883 ( .A(in[1051]), .B(n8955), .Z(n7464) );
  NAND U3884 ( .A(n8985), .B(n7464), .Z(n7314) );
  XNOR U3885 ( .A(n8986), .B(n7314), .Z(out[18]) );
  XOR U3886 ( .A(in[663]), .B(n8695), .Z(n7571) );
  NOR U3887 ( .A(n7412), .B(n8298), .Z(n7315) );
  XNOR U3888 ( .A(n7571), .B(n7315), .Z(out[190]) );
  XOR U3889 ( .A(in[664]), .B(n8697), .Z(n7573) );
  NOR U3890 ( .A(n7414), .B(n8342), .Z(n7316) );
  XNOR U3891 ( .A(n7573), .B(n7316), .Z(out[191]) );
  OR U3892 ( .A(n7417), .B(n8386), .Z(n7317) );
  XNOR U3893 ( .A(n7416), .B(n7317), .Z(out[192]) );
  XOR U3894 ( .A(in[1034]), .B(n8896), .Z(n7420) );
  NOR U3895 ( .A(n7419), .B(n8430), .Z(n7318) );
  XNOR U3896 ( .A(n7420), .B(n7318), .Z(out[193]) );
  XOR U3897 ( .A(in[1035]), .B(n8899), .Z(n7531) );
  NOR U3898 ( .A(n7422), .B(n8474), .Z(n7319) );
  XNOR U3899 ( .A(n7531), .B(n7319), .Z(out[194]) );
  XNOR U3900 ( .A(n8902), .B(in[1036]), .Z(n7681) );
  NOR U3901 ( .A(n7424), .B(n8518), .Z(n7320) );
  XNOR U3902 ( .A(n7681), .B(n7320), .Z(out[195]) );
  XNOR U3903 ( .A(n8905), .B(in[1037]), .Z(n7875) );
  NOR U3904 ( .A(n7427), .B(n8562), .Z(n7321) );
  XNOR U3905 ( .A(n7875), .B(n7321), .Z(out[196]) );
  XNOR U3906 ( .A(n8908), .B(in[1038]), .Z(n8165) );
  NOR U3907 ( .A(n7429), .B(n8606), .Z(n7322) );
  XNOR U3908 ( .A(n8165), .B(n7322), .Z(out[197]) );
  XNOR U3909 ( .A(n8911), .B(in[1039]), .Z(n8607) );
  NOR U3910 ( .A(n7431), .B(n8640), .Z(n7323) );
  XNOR U3911 ( .A(n8607), .B(n7323), .Z(out[198]) );
  XNOR U3912 ( .A(n8914), .B(in[1040]), .Z(n8883) );
  NOR U3913 ( .A(n7433), .B(n8662), .Z(n7324) );
  XNOR U3914 ( .A(n8883), .B(n7324), .Z(out[199]) );
  XNOR U3915 ( .A(in[1429]), .B(n8461), .Z(n9011) );
  XOR U3916 ( .A(in[1052]), .B(n8958), .Z(n7467) );
  NAND U3917 ( .A(n9011), .B(n7467), .Z(n7325) );
  XNOR U3918 ( .A(n9012), .B(n7325), .Z(out[19]) );
  XNOR U3919 ( .A(n8381), .B(in[1411]), .Z(n8427) );
  NANDN U3920 ( .A(n7420), .B(n8427), .Z(n7326) );
  XNOR U3921 ( .A(n8428), .B(n7326), .Z(out[1]) );
  XNOR U3922 ( .A(n8921), .B(in[1041]), .Z(n9167) );
  NOR U3923 ( .A(n7435), .B(n8684), .Z(n7327) );
  XNOR U3924 ( .A(n9167), .B(n7327), .Z(out[200]) );
  XNOR U3925 ( .A(n8924), .B(in[1042]), .Z(n9611) );
  NOR U3926 ( .A(n7437), .B(n8706), .Z(n7328) );
  XNOR U3927 ( .A(n9611), .B(n7328), .Z(out[201]) );
  OR U3928 ( .A(n7440), .B(n8730), .Z(n7329) );
  XNOR U3929 ( .A(n7439), .B(n7329), .Z(out[202]) );
  OR U3930 ( .A(n7443), .B(n8754), .Z(n7330) );
  XNOR U3931 ( .A(n7442), .B(n7330), .Z(out[203]) );
  OR U3932 ( .A(n7446), .B(n8780), .Z(n7331) );
  XNOR U3933 ( .A(n7445), .B(n7331), .Z(out[204]) );
  OR U3934 ( .A(n7449), .B(n8814), .Z(n7332) );
  XNOR U3935 ( .A(n7448), .B(n7332), .Z(out[205]) );
  OR U3936 ( .A(n7453), .B(n8848), .Z(n7333) );
  XNOR U3937 ( .A(n7452), .B(n7333), .Z(out[206]) );
  OR U3938 ( .A(n7456), .B(n8882), .Z(n7334) );
  XNOR U3939 ( .A(n7455), .B(n7334), .Z(out[207]) );
  OR U3940 ( .A(n7459), .B(n8920), .Z(n7335) );
  XNOR U3941 ( .A(n7458), .B(n7335), .Z(out[208]) );
  OR U3942 ( .A(n7462), .B(n8954), .Z(n7336) );
  XNOR U3943 ( .A(n7461), .B(n7336), .Z(out[209]) );
  XNOR U3944 ( .A(in[1430]), .B(n8465), .Z(n9035) );
  XOR U3945 ( .A(in[1053]), .B(n8961), .Z(n7470) );
  NAND U3946 ( .A(n9035), .B(n7470), .Z(n7337) );
  XNOR U3947 ( .A(n9036), .B(n7337), .Z(out[20]) );
  OR U3948 ( .A(n7465), .B(n8988), .Z(n7338) );
  XNOR U3949 ( .A(n7464), .B(n7338), .Z(out[210]) );
  OR U3950 ( .A(n7468), .B(n9014), .Z(n7339) );
  XNOR U3951 ( .A(n7467), .B(n7339), .Z(out[211]) );
  OR U3952 ( .A(n7471), .B(n9038), .Z(n7340) );
  XNOR U3953 ( .A(n7470), .B(n7340), .Z(out[212]) );
  XNOR U3954 ( .A(in[1054]), .B(n8964), .Z(n7474) );
  NOR U3955 ( .A(n7473), .B(n9062), .Z(n7341) );
  XNOR U3956 ( .A(n7474), .B(n7341), .Z(out[213]) );
  XNOR U3957 ( .A(in[1055]), .B(n8967), .Z(n7477) );
  NOR U3958 ( .A(n7476), .B(n9086), .Z(n7342) );
  XNOR U3959 ( .A(n7477), .B(n7342), .Z(out[214]) );
  XNOR U3960 ( .A(in[1056]), .B(n8970), .Z(n7480) );
  NOR U3961 ( .A(n7479), .B(n9110), .Z(n7343) );
  XNOR U3962 ( .A(n7480), .B(n7343), .Z(out[215]) );
  XNOR U3963 ( .A(in[1057]), .B(n8973), .Z(n7484) );
  NOR U3964 ( .A(n7483), .B(n9134), .Z(n7344) );
  XNOR U3965 ( .A(n7484), .B(n7344), .Z(out[216]) );
  XNOR U3966 ( .A(in[1058]), .B(n8976), .Z(n7487) );
  NOR U3967 ( .A(n7486), .B(n9166), .Z(n7345) );
  XNOR U3968 ( .A(n7487), .B(n7345), .Z(out[217]) );
  XNOR U3969 ( .A(in[1059]), .B(n8979), .Z(n7490) );
  NOR U3970 ( .A(n7489), .B(n9214), .Z(n7346) );
  XNOR U3971 ( .A(n7490), .B(n7346), .Z(out[218]) );
  XOR U3972 ( .A(in[1060]), .B(n8982), .Z(n7493) );
  NOR U3973 ( .A(n7492), .B(n9258), .Z(n7347) );
  XNOR U3974 ( .A(n7493), .B(n7347), .Z(out[219]) );
  XNOR U3975 ( .A(in[1431]), .B(n8469), .Z(n9059) );
  NANDN U3976 ( .A(n7474), .B(n9059), .Z(n7348) );
  XNOR U3977 ( .A(n9060), .B(n7348), .Z(out[21]) );
  XOR U3978 ( .A(in[1061]), .B(n8989), .Z(n7507) );
  NOR U3979 ( .A(n7495), .B(n9302), .Z(n7349) );
  XNOR U3980 ( .A(n7507), .B(n7349), .Z(out[220]) );
  XOR U3981 ( .A(in[1062]), .B(n8992), .Z(n7529) );
  NOR U3982 ( .A(n7497), .B(n9346), .Z(n7350) );
  XNOR U3983 ( .A(n7529), .B(n7350), .Z(out[221]) );
  XOR U3984 ( .A(in[1063]), .B(n8771), .Z(n7553) );
  NOR U3985 ( .A(n7499), .B(n9390), .Z(n7351) );
  XNOR U3986 ( .A(n7553), .B(n7351), .Z(out[222]) );
  XOR U3987 ( .A(in[1064]), .B(n8774), .Z(n7575) );
  NOR U3988 ( .A(n7501), .B(n9434), .Z(n7352) );
  XNOR U3989 ( .A(n7575), .B(n7352), .Z(out[223]) );
  XOR U3990 ( .A(in[1065]), .B(n8781), .Z(n7587) );
  NOR U3991 ( .A(n7503), .B(n9478), .Z(n7353) );
  XNOR U3992 ( .A(n7587), .B(n7353), .Z(out[224]) );
  XOR U3993 ( .A(in[1066]), .B(n8784), .Z(n7599) );
  NOR U3994 ( .A(n7505), .B(n9522), .Z(n7354) );
  XNOR U3995 ( .A(n7599), .B(n7354), .Z(out[225]) );
  XOR U3996 ( .A(in[1067]), .B(n8787), .Z(n7611) );
  NOR U3997 ( .A(n7509), .B(n9566), .Z(n7355) );
  XNOR U3998 ( .A(n7611), .B(n7355), .Z(out[226]) );
  XOR U3999 ( .A(in[1068]), .B(n8790), .Z(n7623) );
  NOR U4000 ( .A(n7511), .B(n9610), .Z(n7356) );
  XNOR U4001 ( .A(n7623), .B(n7356), .Z(out[227]) );
  XNOR U4002 ( .A(in[1069]), .B(n8793), .Z(n7636) );
  NAND U4003 ( .A(n7513), .B(n7357), .Z(n7358) );
  XNOR U4004 ( .A(n7636), .B(n7358), .Z(out[228]) );
  XNOR U4005 ( .A(in[1070]), .B(n8796), .Z(n7650) );
  NAND U4006 ( .A(n7515), .B(n7359), .Z(n7360) );
  XNOR U4007 ( .A(n7650), .B(n7360), .Z(out[229]) );
  XNOR U4008 ( .A(in[1432]), .B(n8477), .Z(n9083) );
  NANDN U4009 ( .A(n7477), .B(n9083), .Z(n7361) );
  XNOR U4010 ( .A(n9084), .B(n7361), .Z(out[22]) );
  XNOR U4011 ( .A(in[1071]), .B(n8799), .Z(n7664) );
  NAND U4012 ( .A(n7517), .B(n7362), .Z(n7363) );
  XNOR U4013 ( .A(n7664), .B(n7363), .Z(out[230]) );
  XNOR U4014 ( .A(in[1072]), .B(n8802), .Z(n7678) );
  NAND U4015 ( .A(n7519), .B(n7364), .Z(n7365) );
  XNOR U4016 ( .A(n7678), .B(n7365), .Z(out[231]) );
  XNOR U4017 ( .A(in[1073]), .B(n8805), .Z(n7694) );
  NAND U4018 ( .A(n7521), .B(n7366), .Z(n7367) );
  XNOR U4019 ( .A(n7694), .B(n7367), .Z(out[232]) );
  XNOR U4020 ( .A(in[1074]), .B(n8808), .Z(n7708) );
  NAND U4021 ( .A(n7523), .B(n7368), .Z(n7369) );
  XNOR U4022 ( .A(n7708), .B(n7369), .Z(out[233]) );
  XNOR U4023 ( .A(in[1075]), .B(n8815), .Z(n7722) );
  NAND U4024 ( .A(n7525), .B(n7370), .Z(n7371) );
  XNOR U4025 ( .A(n7722), .B(n7371), .Z(out[234]) );
  XNOR U4026 ( .A(in[1076]), .B(n8818), .Z(n7736) );
  NAND U4027 ( .A(n7527), .B(n7372), .Z(n7373) );
  XNOR U4028 ( .A(n7736), .B(n7373), .Z(out[235]) );
  XNOR U4029 ( .A(in[1077]), .B(n8821), .Z(n7752) );
  NAND U4030 ( .A(n7533), .B(n7374), .Z(n7375) );
  XNOR U4031 ( .A(n7752), .B(n7375), .Z(out[236]) );
  XNOR U4032 ( .A(in[1078]), .B(n8824), .Z(n7776) );
  NAND U4033 ( .A(n7535), .B(n7376), .Z(n7377) );
  XNOR U4034 ( .A(n7776), .B(n7377), .Z(out[237]) );
  XNOR U4035 ( .A(in[1079]), .B(n8827), .Z(n7800) );
  NAND U4036 ( .A(n7537), .B(n7378), .Z(n7379) );
  XNOR U4037 ( .A(n7800), .B(n7379), .Z(out[238]) );
  XNOR U4038 ( .A(in[1080]), .B(n8830), .Z(n7824) );
  NAND U4039 ( .A(n7539), .B(n7380), .Z(n7381) );
  XNOR U4040 ( .A(n7824), .B(n7381), .Z(out[239]) );
  XNOR U4041 ( .A(in[1433]), .B(n8481), .Z(n9107) );
  NANDN U4042 ( .A(n7480), .B(n9107), .Z(n7382) );
  XNOR U4043 ( .A(n9108), .B(n7382), .Z(out[23]) );
  XNOR U4044 ( .A(in[1081]), .B(n8833), .Z(n7848) );
  NAND U4045 ( .A(n7541), .B(n7383), .Z(n7384) );
  XNOR U4046 ( .A(n7848), .B(n7384), .Z(out[240]) );
  XNOR U4047 ( .A(in[1082]), .B(n8836), .Z(n7872) );
  NAND U4048 ( .A(n7543), .B(n7385), .Z(n7386) );
  XNOR U4049 ( .A(n7872), .B(n7386), .Z(out[241]) );
  XNOR U4050 ( .A(in[1083]), .B(n8839), .Z(n7898) );
  NAND U4051 ( .A(n7545), .B(n7387), .Z(n7388) );
  XNOR U4052 ( .A(n7898), .B(n7388), .Z(out[242]) );
  XNOR U4053 ( .A(in[1084]), .B(n8842), .Z(n7922) );
  NAND U4054 ( .A(n7547), .B(n7389), .Z(n7390) );
  XNOR U4055 ( .A(n7922), .B(n7390), .Z(out[243]) );
  XNOR U4056 ( .A(in[1085]), .B(n8849), .Z(n7946) );
  NAND U4057 ( .A(n7549), .B(n7391), .Z(n7392) );
  XNOR U4058 ( .A(n7946), .B(n7392), .Z(out[244]) );
  XNOR U4059 ( .A(in[1086]), .B(n8852), .Z(n7970) );
  NAND U4060 ( .A(n7551), .B(n7393), .Z(n7394) );
  XNOR U4061 ( .A(n7970), .B(n7394), .Z(out[245]) );
  XNOR U4062 ( .A(in[1087]), .B(n8855), .Z(n7994) );
  NAND U4063 ( .A(n7555), .B(n7395), .Z(n7396) );
  XNOR U4064 ( .A(n7994), .B(n7396), .Z(out[246]) );
  XNOR U4065 ( .A(in[1024]), .B(n8858), .Z(n8018) );
  NAND U4066 ( .A(n7557), .B(n7397), .Z(n7398) );
  XNOR U4067 ( .A(n8018), .B(n7398), .Z(out[247]) );
  XNOR U4068 ( .A(in[1025]), .B(n8861), .Z(n8042) );
  NAND U4069 ( .A(n7559), .B(n7399), .Z(n7400) );
  XNOR U4070 ( .A(n8042), .B(n7400), .Z(out[248]) );
  XNOR U4071 ( .A(in[1026]), .B(n8864), .Z(n8074) );
  NAND U4072 ( .A(n7561), .B(n7401), .Z(n7402) );
  XNOR U4073 ( .A(n8074), .B(n7402), .Z(out[249]) );
  XNOR U4074 ( .A(in[1434]), .B(n8485), .Z(n9131) );
  NANDN U4075 ( .A(n7484), .B(n9131), .Z(n7403) );
  XNOR U4076 ( .A(n9132), .B(n7403), .Z(out[24]) );
  XNOR U4077 ( .A(in[1027]), .B(n8867), .Z(n8118) );
  NAND U4078 ( .A(n7563), .B(n7404), .Z(n7405) );
  XNOR U4079 ( .A(n8118), .B(n7405), .Z(out[250]) );
  XNOR U4080 ( .A(in[1028]), .B(n8870), .Z(n8162) );
  NAND U4081 ( .A(n7565), .B(n7406), .Z(n7407) );
  XNOR U4082 ( .A(n8162), .B(n7407), .Z(out[251]) );
  XNOR U4083 ( .A(in[1029]), .B(n8873), .Z(n8208) );
  NAND U4084 ( .A(n7567), .B(n7408), .Z(n7409) );
  XNOR U4085 ( .A(n8208), .B(n7409), .Z(out[252]) );
  XNOR U4086 ( .A(in[1030]), .B(n8876), .Z(n8252) );
  NAND U4087 ( .A(n7569), .B(n7410), .Z(n7411) );
  XNOR U4088 ( .A(n8252), .B(n7411), .Z(out[253]) );
  XNOR U4089 ( .A(in[1031]), .B(n8887), .Z(n8296) );
  NAND U4090 ( .A(n7571), .B(n7412), .Z(n7413) );
  XNOR U4091 ( .A(n8296), .B(n7413), .Z(out[254]) );
  XNOR U4092 ( .A(in[1032]), .B(n8890), .Z(n8340) );
  NAND U4093 ( .A(n7573), .B(n7414), .Z(n7415) );
  XNOR U4094 ( .A(n8340), .B(n7415), .Z(out[255]) );
  ANDN U4095 ( .B(n7417), .A(n7416), .Z(n7418) );
  XNOR U4096 ( .A(n8383), .B(n7418), .Z(out[256]) );
  AND U4097 ( .A(n7420), .B(n7419), .Z(n7421) );
  XNOR U4098 ( .A(n8427), .B(n7421), .Z(out[257]) );
  XOR U4099 ( .A(n8389), .B(in[1412]), .Z(n8472) );
  NAND U4100 ( .A(n7531), .B(n7422), .Z(n7423) );
  XNOR U4101 ( .A(n8472), .B(n7423), .Z(out[258]) );
  XOR U4102 ( .A(n8393), .B(in[1413]), .Z(n8516) );
  NAND U4103 ( .A(n7681), .B(n7424), .Z(n7425) );
  XNOR U4104 ( .A(n8516), .B(n7425), .Z(out[259]) );
  XNOR U4105 ( .A(in[1435]), .B(n8489), .Z(n9163) );
  NANDN U4106 ( .A(n7487), .B(n9163), .Z(n7426) );
  XNOR U4107 ( .A(n9164), .B(n7426), .Z(out[25]) );
  XOR U4108 ( .A(n8397), .B(in[1414]), .Z(n8560) );
  NAND U4109 ( .A(n7875), .B(n7427), .Z(n7428) );
  XNOR U4110 ( .A(n8560), .B(n7428), .Z(out[260]) );
  XOR U4111 ( .A(n8401), .B(in[1415]), .Z(n8604) );
  NAND U4112 ( .A(n8165), .B(n7429), .Z(n7430) );
  XNOR U4113 ( .A(n8604), .B(n7430), .Z(out[261]) );
  XOR U4114 ( .A(n8405), .B(in[1416]), .Z(n8638) );
  NAND U4115 ( .A(n8607), .B(n7431), .Z(n7432) );
  XNOR U4116 ( .A(n8638), .B(n7432), .Z(out[262]) );
  XOR U4117 ( .A(in[1417]), .B(n8409), .Z(n8884) );
  NAND U4118 ( .A(n8883), .B(n7433), .Z(n7434) );
  XNOR U4119 ( .A(n8884), .B(n7434), .Z(out[263]) );
  XOR U4120 ( .A(n8413), .B(in[1418]), .Z(n9168) );
  NAND U4121 ( .A(n9167), .B(n7435), .Z(n7436) );
  XNOR U4122 ( .A(n9168), .B(n7436), .Z(out[264]) );
  XOR U4123 ( .A(n8417), .B(in[1419]), .Z(n9612) );
  NAND U4124 ( .A(n9611), .B(n7437), .Z(n7438) );
  XNOR U4125 ( .A(n9612), .B(n7438), .Z(out[265]) );
  ANDN U4126 ( .B(n7440), .A(n7439), .Z(n7441) );
  XNOR U4127 ( .A(n8727), .B(n7441), .Z(out[266]) );
  ANDN U4128 ( .B(n7443), .A(n7442), .Z(n7444) );
  XNOR U4129 ( .A(n8751), .B(n7444), .Z(out[267]) );
  ANDN U4130 ( .B(n7446), .A(n7445), .Z(n7447) );
  XNOR U4131 ( .A(n8777), .B(n7447), .Z(out[268]) );
  ANDN U4132 ( .B(n7449), .A(n7448), .Z(n7450) );
  XNOR U4133 ( .A(n8811), .B(n7450), .Z(out[269]) );
  XNOR U4134 ( .A(in[1436]), .B(n8493), .Z(n9211) );
  NANDN U4135 ( .A(n7490), .B(n9211), .Z(n7451) );
  XNOR U4136 ( .A(n9212), .B(n7451), .Z(out[26]) );
  ANDN U4137 ( .B(n7453), .A(n7452), .Z(n7454) );
  XNOR U4138 ( .A(n8845), .B(n7454), .Z(out[270]) );
  ANDN U4139 ( .B(n7456), .A(n7455), .Z(n7457) );
  XNOR U4140 ( .A(n8879), .B(n7457), .Z(out[271]) );
  ANDN U4141 ( .B(n7459), .A(n7458), .Z(n7460) );
  XNOR U4142 ( .A(n8917), .B(n7460), .Z(out[272]) );
  ANDN U4143 ( .B(n7462), .A(n7461), .Z(n7463) );
  XNOR U4144 ( .A(n8951), .B(n7463), .Z(out[273]) );
  ANDN U4145 ( .B(n7465), .A(n7464), .Z(n7466) );
  XNOR U4146 ( .A(n8985), .B(n7466), .Z(out[274]) );
  ANDN U4147 ( .B(n7468), .A(n7467), .Z(n7469) );
  XNOR U4148 ( .A(n9011), .B(n7469), .Z(out[275]) );
  ANDN U4149 ( .B(n7471), .A(n7470), .Z(n7472) );
  XNOR U4150 ( .A(n9035), .B(n7472), .Z(out[276]) );
  AND U4151 ( .A(n7474), .B(n7473), .Z(n7475) );
  XNOR U4152 ( .A(n9059), .B(n7475), .Z(out[277]) );
  AND U4153 ( .A(n7477), .B(n7476), .Z(n7478) );
  XNOR U4154 ( .A(n9083), .B(n7478), .Z(out[278]) );
  AND U4155 ( .A(n7480), .B(n7479), .Z(n7481) );
  XNOR U4156 ( .A(n9107), .B(n7481), .Z(out[279]) );
  XNOR U4157 ( .A(in[1437]), .B(n8497), .Z(n9255) );
  NANDN U4158 ( .A(n7493), .B(n9255), .Z(n7482) );
  XNOR U4159 ( .A(n9256), .B(n7482), .Z(out[27]) );
  AND U4160 ( .A(n7484), .B(n7483), .Z(n7485) );
  XNOR U4161 ( .A(n9131), .B(n7485), .Z(out[280]) );
  AND U4162 ( .A(n7487), .B(n7486), .Z(n7488) );
  XNOR U4163 ( .A(n9163), .B(n7488), .Z(out[281]) );
  AND U4164 ( .A(n7490), .B(n7489), .Z(n7491) );
  XNOR U4165 ( .A(n9211), .B(n7491), .Z(out[282]) );
  AND U4166 ( .A(n7493), .B(n7492), .Z(n7494) );
  XNOR U4167 ( .A(n9255), .B(n7494), .Z(out[283]) );
  XOR U4168 ( .A(in[1438]), .B(n8501), .Z(n9300) );
  NAND U4169 ( .A(n7507), .B(n7495), .Z(n7496) );
  XNOR U4170 ( .A(n9300), .B(n7496), .Z(out[284]) );
  XOR U4171 ( .A(in[1439]), .B(n8505), .Z(n9344) );
  NAND U4172 ( .A(n7529), .B(n7497), .Z(n7498) );
  XNOR U4173 ( .A(n9344), .B(n7498), .Z(out[285]) );
  XOR U4174 ( .A(in[1440]), .B(n8509), .Z(n9388) );
  NAND U4175 ( .A(n7553), .B(n7499), .Z(n7500) );
  XNOR U4176 ( .A(n9388), .B(n7500), .Z(out[286]) );
  XOR U4177 ( .A(in[1441]), .B(n8513), .Z(n9432) );
  NAND U4178 ( .A(n7575), .B(n7501), .Z(n7502) );
  XNOR U4179 ( .A(n9432), .B(n7502), .Z(out[287]) );
  XOR U4180 ( .A(in[1442]), .B(n8521), .Z(n9476) );
  NAND U4181 ( .A(n7587), .B(n7503), .Z(n7504) );
  XNOR U4182 ( .A(n9476), .B(n7504), .Z(out[288]) );
  XOR U4183 ( .A(in[1443]), .B(n8525), .Z(n9520) );
  NAND U4184 ( .A(n7599), .B(n7505), .Z(n7506) );
  XNOR U4185 ( .A(n9520), .B(n7506), .Z(out[289]) );
  OR U4186 ( .A(n9300), .B(n7507), .Z(n7508) );
  XNOR U4187 ( .A(n9299), .B(n7508), .Z(out[28]) );
  XOR U4188 ( .A(in[1444]), .B(n8529), .Z(n9564) );
  NAND U4189 ( .A(n7611), .B(n7509), .Z(n7510) );
  XNOR U4190 ( .A(n9564), .B(n7510), .Z(out[290]) );
  XOR U4191 ( .A(in[1445]), .B(n8533), .Z(n9608) );
  NAND U4192 ( .A(n7623), .B(n7511), .Z(n7512) );
  XNOR U4193 ( .A(n9608), .B(n7512), .Z(out[291]) );
  OR U4194 ( .A(n7636), .B(n7513), .Z(n7514) );
  XNOR U4195 ( .A(n7635), .B(n7514), .Z(out[292]) );
  OR U4196 ( .A(n7650), .B(n7515), .Z(n7516) );
  XNOR U4197 ( .A(n7649), .B(n7516), .Z(out[293]) );
  OR U4198 ( .A(n7664), .B(n7517), .Z(n7518) );
  XNOR U4199 ( .A(n7663), .B(n7518), .Z(out[294]) );
  OR U4200 ( .A(n7678), .B(n7519), .Z(n7520) );
  XNOR U4201 ( .A(n7677), .B(n7520), .Z(out[295]) );
  OR U4202 ( .A(n7694), .B(n7521), .Z(n7522) );
  XNOR U4203 ( .A(n7693), .B(n7522), .Z(out[296]) );
  OR U4204 ( .A(n7708), .B(n7523), .Z(n7524) );
  XNOR U4205 ( .A(n7707), .B(n7524), .Z(out[297]) );
  OR U4206 ( .A(n7722), .B(n7525), .Z(n7526) );
  XNOR U4207 ( .A(n7721), .B(n7526), .Z(out[298]) );
  OR U4208 ( .A(n7736), .B(n7527), .Z(n7528) );
  XNOR U4209 ( .A(n7735), .B(n7528), .Z(out[299]) );
  OR U4210 ( .A(n9344), .B(n7529), .Z(n7530) );
  XNOR U4211 ( .A(n9343), .B(n7530), .Z(out[29]) );
  OR U4212 ( .A(n8472), .B(n7531), .Z(n7532) );
  XNOR U4213 ( .A(n8471), .B(n7532), .Z(out[2]) );
  OR U4214 ( .A(n7752), .B(n7533), .Z(n7534) );
  XNOR U4215 ( .A(n7751), .B(n7534), .Z(out[300]) );
  OR U4216 ( .A(n7776), .B(n7535), .Z(n7536) );
  XNOR U4217 ( .A(n7775), .B(n7536), .Z(out[301]) );
  OR U4218 ( .A(n7800), .B(n7537), .Z(n7538) );
  XNOR U4219 ( .A(n7799), .B(n7538), .Z(out[302]) );
  OR U4220 ( .A(n7824), .B(n7539), .Z(n7540) );
  XNOR U4221 ( .A(n7823), .B(n7540), .Z(out[303]) );
  OR U4222 ( .A(n7848), .B(n7541), .Z(n7542) );
  XNOR U4223 ( .A(n7847), .B(n7542), .Z(out[304]) );
  OR U4224 ( .A(n7872), .B(n7543), .Z(n7544) );
  XNOR U4225 ( .A(n7871), .B(n7544), .Z(out[305]) );
  OR U4226 ( .A(n7898), .B(n7545), .Z(n7546) );
  XNOR U4227 ( .A(n7897), .B(n7546), .Z(out[306]) );
  OR U4228 ( .A(n7922), .B(n7547), .Z(n7548) );
  XNOR U4229 ( .A(n7921), .B(n7548), .Z(out[307]) );
  OR U4230 ( .A(n7946), .B(n7549), .Z(n7550) );
  XNOR U4231 ( .A(n7945), .B(n7550), .Z(out[308]) );
  OR U4232 ( .A(n7970), .B(n7551), .Z(n7552) );
  XNOR U4233 ( .A(n7969), .B(n7552), .Z(out[309]) );
  OR U4234 ( .A(n9388), .B(n7553), .Z(n7554) );
  XNOR U4235 ( .A(n9387), .B(n7554), .Z(out[30]) );
  OR U4236 ( .A(n7994), .B(n7555), .Z(n7556) );
  XNOR U4237 ( .A(n7993), .B(n7556), .Z(out[310]) );
  OR U4238 ( .A(n8018), .B(n7557), .Z(n7558) );
  XNOR U4239 ( .A(n8017), .B(n7558), .Z(out[311]) );
  OR U4240 ( .A(n8042), .B(n7559), .Z(n7560) );
  XNOR U4241 ( .A(n8041), .B(n7560), .Z(out[312]) );
  OR U4242 ( .A(n8074), .B(n7561), .Z(n7562) );
  XNOR U4243 ( .A(n8073), .B(n7562), .Z(out[313]) );
  OR U4244 ( .A(n8118), .B(n7563), .Z(n7564) );
  XNOR U4245 ( .A(n8117), .B(n7564), .Z(out[314]) );
  OR U4246 ( .A(n8162), .B(n7565), .Z(n7566) );
  XNOR U4247 ( .A(n8161), .B(n7566), .Z(out[315]) );
  OR U4248 ( .A(n8208), .B(n7567), .Z(n7568) );
  XNOR U4249 ( .A(n8207), .B(n7568), .Z(out[316]) );
  OR U4250 ( .A(n8252), .B(n7569), .Z(n7570) );
  XNOR U4251 ( .A(n8251), .B(n7570), .Z(out[317]) );
  OR U4252 ( .A(n8296), .B(n7571), .Z(n7572) );
  XNOR U4253 ( .A(n8295), .B(n7572), .Z(out[318]) );
  OR U4254 ( .A(n8340), .B(n7573), .Z(n7574) );
  XNOR U4255 ( .A(n8339), .B(n7574), .Z(out[319]) );
  OR U4256 ( .A(n9432), .B(n7575), .Z(n7576) );
  XNOR U4257 ( .A(n9431), .B(n7576), .Z(out[31]) );
  XNOR U4258 ( .A(in[72]), .B(n8890), .Z(n7747) );
  XOR U4259 ( .A(in[1317]), .B(n8725), .Z(n8060) );
  XOR U4260 ( .A(in[1244]), .B(n8543), .Z(n8057) );
  NAND U4261 ( .A(n8060), .B(n8057), .Z(n7577) );
  XNOR U4262 ( .A(n7747), .B(n7577), .Z(out[320]) );
  XNOR U4263 ( .A(in[73]), .B(n8893), .Z(n7749) );
  XOR U4264 ( .A(in[1318]), .B(n8731), .Z(n8064) );
  XOR U4265 ( .A(in[1245]), .B(n8547), .Z(n8061) );
  NAND U4266 ( .A(n8064), .B(n8061), .Z(n7578) );
  XNOR U4267 ( .A(n7749), .B(n7578), .Z(out[321]) );
  XNOR U4268 ( .A(in[74]), .B(n8896), .Z(n7755) );
  XOR U4269 ( .A(in[1319]), .B(n8733), .Z(n8068) );
  XOR U4270 ( .A(in[1246]), .B(n8551), .Z(n8065) );
  NAND U4271 ( .A(n8068), .B(n8065), .Z(n7579) );
  XNOR U4272 ( .A(n7755), .B(n7579), .Z(out[322]) );
  XNOR U4273 ( .A(in[75]), .B(n8899), .Z(n7757) );
  XOR U4274 ( .A(in[1320]), .B(n8735), .Z(n8072) );
  XOR U4275 ( .A(in[1247]), .B(n8555), .Z(n8069) );
  NAND U4276 ( .A(n8072), .B(n8069), .Z(n7580) );
  XNOR U4277 ( .A(n7757), .B(n7580), .Z(out[323]) );
  XOR U4278 ( .A(n8902), .B(in[76]), .Z(n7759) );
  XOR U4279 ( .A(in[1321]), .B(n8737), .Z(n8080) );
  XOR U4280 ( .A(in[1248]), .B(n8563), .Z(n8077) );
  NAND U4281 ( .A(n8080), .B(n8077), .Z(n7581) );
  XNOR U4282 ( .A(n7759), .B(n7581), .Z(out[324]) );
  XOR U4283 ( .A(n8905), .B(in[77]), .Z(n7761) );
  XOR U4284 ( .A(in[1322]), .B(n8739), .Z(n8084) );
  XOR U4285 ( .A(in[1249]), .B(n8567), .Z(n8081) );
  NAND U4286 ( .A(n8084), .B(n8081), .Z(n7582) );
  XNOR U4287 ( .A(n7761), .B(n7582), .Z(out[325]) );
  XOR U4288 ( .A(n8908), .B(in[78]), .Z(n7763) );
  XOR U4289 ( .A(in[1323]), .B(n8741), .Z(n8088) );
  XOR U4290 ( .A(in[1250]), .B(n8571), .Z(n8085) );
  NAND U4291 ( .A(n8088), .B(n8085), .Z(n7583) );
  XNOR U4292 ( .A(n7763), .B(n7583), .Z(out[326]) );
  XOR U4293 ( .A(n8911), .B(in[79]), .Z(n7765) );
  XOR U4294 ( .A(in[1324]), .B(n8743), .Z(n8092) );
  XOR U4295 ( .A(in[1251]), .B(n8575), .Z(n8089) );
  NAND U4296 ( .A(n8092), .B(n8089), .Z(n7584) );
  XNOR U4297 ( .A(n7765), .B(n7584), .Z(out[327]) );
  XOR U4298 ( .A(n8914), .B(in[80]), .Z(n7767) );
  XOR U4299 ( .A(in[1325]), .B(n8745), .Z(n8096) );
  XOR U4300 ( .A(in[1252]), .B(n8579), .Z(n8093) );
  NAND U4301 ( .A(n8096), .B(n8093), .Z(n7585) );
  XNOR U4302 ( .A(n7767), .B(n7585), .Z(out[328]) );
  XOR U4303 ( .A(n8921), .B(in[81]), .Z(n7769) );
  XOR U4304 ( .A(in[1326]), .B(n8747), .Z(n8100) );
  XNOR U4305 ( .A(in[1253]), .B(n8583), .Z(n8097) );
  NAND U4306 ( .A(n8100), .B(n8097), .Z(n7586) );
  XNOR U4307 ( .A(n7769), .B(n7586), .Z(out[329]) );
  OR U4308 ( .A(n9476), .B(n7587), .Z(n7588) );
  XNOR U4309 ( .A(n9475), .B(n7588), .Z(out[32]) );
  XOR U4310 ( .A(n8924), .B(in[82]), .Z(n7771) );
  XOR U4311 ( .A(in[1327]), .B(n8749), .Z(n8104) );
  XNOR U4312 ( .A(in[1254]), .B(n8587), .Z(n8101) );
  NAND U4313 ( .A(n8104), .B(n8101), .Z(n7589) );
  XNOR U4314 ( .A(n7771), .B(n7589), .Z(out[330]) );
  XOR U4315 ( .A(n8927), .B(in[83]), .Z(n7773) );
  XOR U4316 ( .A(in[1328]), .B(n8755), .Z(n8108) );
  XNOR U4317 ( .A(in[1255]), .B(n8591), .Z(n8105) );
  NAND U4318 ( .A(n8108), .B(n8105), .Z(n7590) );
  XNOR U4319 ( .A(n7773), .B(n7590), .Z(out[331]) );
  XOR U4320 ( .A(in[84]), .B(n8930), .Z(n7779) );
  XOR U4321 ( .A(in[1329]), .B(n8757), .Z(n8112) );
  XNOR U4322 ( .A(in[1256]), .B(n8595), .Z(n8109) );
  NAND U4323 ( .A(n8112), .B(n8109), .Z(n7591) );
  XNOR U4324 ( .A(n7779), .B(n7591), .Z(out[332]) );
  XOR U4325 ( .A(in[85]), .B(n8933), .Z(n7781) );
  XOR U4326 ( .A(in[1330]), .B(n8759), .Z(n8116) );
  XNOR U4327 ( .A(in[1257]), .B(n8599), .Z(n8113) );
  NAND U4328 ( .A(n8116), .B(n8113), .Z(n7592) );
  XNOR U4329 ( .A(n7781), .B(n7592), .Z(out[333]) );
  XOR U4330 ( .A(in[86]), .B(n8936), .Z(n7783) );
  XOR U4331 ( .A(in[1331]), .B(n8761), .Z(n8124) );
  XNOR U4332 ( .A(in[1258]), .B(n8609), .Z(n8121) );
  NAND U4333 ( .A(n8124), .B(n8121), .Z(n7593) );
  XNOR U4334 ( .A(n7783), .B(n7593), .Z(out[334]) );
  XOR U4335 ( .A(in[87]), .B(n8939), .Z(n7785) );
  XOR U4336 ( .A(in[1332]), .B(n8763), .Z(n8128) );
  XNOR U4337 ( .A(in[1259]), .B(n8613), .Z(n8125) );
  NAND U4338 ( .A(n8128), .B(n8125), .Z(n7594) );
  XNOR U4339 ( .A(n7785), .B(n7594), .Z(out[335]) );
  XOR U4340 ( .A(in[88]), .B(n8942), .Z(n7787) );
  XOR U4341 ( .A(in[1333]), .B(n8765), .Z(n8132) );
  XNOR U4342 ( .A(in[1260]), .B(n8617), .Z(n8129) );
  NAND U4343 ( .A(n8132), .B(n8129), .Z(n7595) );
  XNOR U4344 ( .A(n7787), .B(n7595), .Z(out[336]) );
  XOR U4345 ( .A(in[89]), .B(n8945), .Z(n7789) );
  XOR U4346 ( .A(in[1334]), .B(n8767), .Z(n8136) );
  XNOR U4347 ( .A(in[1261]), .B(n8621), .Z(n8133) );
  NAND U4348 ( .A(n8136), .B(n8133), .Z(n7596) );
  XNOR U4349 ( .A(n7789), .B(n7596), .Z(out[337]) );
  XOR U4350 ( .A(in[90]), .B(n8948), .Z(n7791) );
  XOR U4351 ( .A(in[1335]), .B(n8769), .Z(n8140) );
  XNOR U4352 ( .A(in[1262]), .B(n8343), .Z(n8137) );
  NAND U4353 ( .A(n8140), .B(n8137), .Z(n7597) );
  XNOR U4354 ( .A(n7791), .B(n7597), .Z(out[338]) );
  XOR U4355 ( .A(in[91]), .B(n8955), .Z(n7793) );
  XOR U4356 ( .A(in[1336]), .B(n8625), .Z(n8144) );
  XNOR U4357 ( .A(in[1263]), .B(n8347), .Z(n8141) );
  NAND U4358 ( .A(n8144), .B(n8141), .Z(n7598) );
  XNOR U4359 ( .A(n7793), .B(n7598), .Z(out[339]) );
  OR U4360 ( .A(n9520), .B(n7599), .Z(n7600) );
  XNOR U4361 ( .A(n9519), .B(n7600), .Z(out[33]) );
  XOR U4362 ( .A(in[92]), .B(n8958), .Z(n7795) );
  XOR U4363 ( .A(in[1337]), .B(n8627), .Z(n8148) );
  XNOR U4364 ( .A(in[1264]), .B(n8351), .Z(n8145) );
  NAND U4365 ( .A(n8148), .B(n8145), .Z(n7601) );
  XNOR U4366 ( .A(n7795), .B(n7601), .Z(out[340]) );
  XOR U4367 ( .A(in[93]), .B(n8961), .Z(n7797) );
  XOR U4368 ( .A(in[1338]), .B(n8629), .Z(n8152) );
  XNOR U4369 ( .A(in[1265]), .B(n8355), .Z(n8149) );
  NAND U4370 ( .A(n8152), .B(n8149), .Z(n7602) );
  XNOR U4371 ( .A(n7797), .B(n7602), .Z(out[341]) );
  XOR U4372 ( .A(in[94]), .B(n8964), .Z(n7803) );
  XOR U4373 ( .A(in[1339]), .B(n8631), .Z(n8156) );
  XNOR U4374 ( .A(in[1266]), .B(n8359), .Z(n8153) );
  NAND U4375 ( .A(n8156), .B(n8153), .Z(n7603) );
  XNOR U4376 ( .A(n7803), .B(n7603), .Z(out[342]) );
  XOR U4377 ( .A(in[95]), .B(n8967), .Z(n7805) );
  XOR U4378 ( .A(in[1340]), .B(n8633), .Z(n8160) );
  XNOR U4379 ( .A(in[1267]), .B(n8363), .Z(n8157) );
  NAND U4380 ( .A(n8160), .B(n8157), .Z(n7604) );
  XNOR U4381 ( .A(n7805), .B(n7604), .Z(out[343]) );
  XOR U4382 ( .A(in[96]), .B(n8970), .Z(n7807) );
  XOR U4383 ( .A(in[1341]), .B(n8635), .Z(n8170) );
  XNOR U4384 ( .A(in[1268]), .B(n8367), .Z(n8167) );
  NAND U4385 ( .A(n8170), .B(n8167), .Z(n7605) );
  XNOR U4386 ( .A(n7807), .B(n7605), .Z(out[344]) );
  XOR U4387 ( .A(in[97]), .B(n8973), .Z(n7809) );
  XOR U4388 ( .A(in[1342]), .B(n8641), .Z(n8174) );
  XNOR U4389 ( .A(in[1269]), .B(n8371), .Z(n8171) );
  NAND U4390 ( .A(n8174), .B(n8171), .Z(n7606) );
  XNOR U4391 ( .A(n7809), .B(n7606), .Z(out[345]) );
  XOR U4392 ( .A(in[98]), .B(n8976), .Z(n7811) );
  XOR U4393 ( .A(in[1343]), .B(n8643), .Z(n8178) );
  XNOR U4394 ( .A(in[1270]), .B(n8375), .Z(n8175) );
  NAND U4395 ( .A(n8178), .B(n8175), .Z(n7607) );
  XNOR U4396 ( .A(n7811), .B(n7607), .Z(out[346]) );
  XOR U4397 ( .A(in[99]), .B(n8979), .Z(n7813) );
  XOR U4398 ( .A(in[1280]), .B(n8645), .Z(n8182) );
  XNOR U4399 ( .A(in[1271]), .B(n8379), .Z(n8179) );
  NAND U4400 ( .A(n8182), .B(n8179), .Z(n7608) );
  XNOR U4401 ( .A(n7813), .B(n7608), .Z(out[347]) );
  XNOR U4402 ( .A(in[100]), .B(n8982), .Z(n7815) );
  XOR U4403 ( .A(in[1281]), .B(n8647), .Z(n8186) );
  XNOR U4404 ( .A(in[1272]), .B(n8387), .Z(n8183) );
  NAND U4405 ( .A(n8186), .B(n8183), .Z(n7609) );
  XNOR U4406 ( .A(n7815), .B(n7609), .Z(out[348]) );
  XNOR U4407 ( .A(in[101]), .B(n8989), .Z(n7817) );
  XOR U4408 ( .A(in[1282]), .B(n8649), .Z(n8190) );
  XNOR U4409 ( .A(in[1273]), .B(n8391), .Z(n8187) );
  NAND U4410 ( .A(n8190), .B(n8187), .Z(n7610) );
  XNOR U4411 ( .A(n7817), .B(n7610), .Z(out[349]) );
  OR U4412 ( .A(n9564), .B(n7611), .Z(n7612) );
  XNOR U4413 ( .A(n9563), .B(n7612), .Z(out[34]) );
  XNOR U4414 ( .A(in[102]), .B(n8992), .Z(n7819) );
  XOR U4415 ( .A(in[1283]), .B(n8651), .Z(n8194) );
  XNOR U4416 ( .A(in[1274]), .B(n8395), .Z(n8191) );
  NAND U4417 ( .A(n8194), .B(n8191), .Z(n7613) );
  XNOR U4418 ( .A(n7819), .B(n7613), .Z(out[350]) );
  XNOR U4419 ( .A(in[103]), .B(n8771), .Z(n7821) );
  XOR U4420 ( .A(in[1284]), .B(n8653), .Z(n8198) );
  XNOR U4421 ( .A(in[1275]), .B(n8399), .Z(n8195) );
  NAND U4422 ( .A(n8198), .B(n8195), .Z(n7614) );
  XNOR U4423 ( .A(n7821), .B(n7614), .Z(out[351]) );
  XNOR U4424 ( .A(in[104]), .B(n8774), .Z(n7827) );
  XOR U4425 ( .A(in[1285]), .B(n8655), .Z(n8202) );
  XNOR U4426 ( .A(in[1276]), .B(n8403), .Z(n8199) );
  NAND U4427 ( .A(n8202), .B(n8199), .Z(n7615) );
  XNOR U4428 ( .A(n7827), .B(n7615), .Z(out[352]) );
  XNOR U4429 ( .A(in[105]), .B(n8781), .Z(n7829) );
  XOR U4430 ( .A(in[1286]), .B(n8657), .Z(n8206) );
  XNOR U4431 ( .A(in[1277]), .B(n8407), .Z(n8203) );
  NAND U4432 ( .A(n8206), .B(n8203), .Z(n7616) );
  XNOR U4433 ( .A(n7829), .B(n7616), .Z(out[353]) );
  XNOR U4434 ( .A(in[106]), .B(n8784), .Z(n7831) );
  XOR U4435 ( .A(in[1287]), .B(n8659), .Z(n8214) );
  XNOR U4436 ( .A(in[1278]), .B(n8411), .Z(n8211) );
  NAND U4437 ( .A(n8214), .B(n8211), .Z(n7617) );
  XNOR U4438 ( .A(n7831), .B(n7617), .Z(out[354]) );
  XNOR U4439 ( .A(in[107]), .B(n8787), .Z(n7833) );
  XOR U4440 ( .A(in[1288]), .B(n8663), .Z(n8218) );
  XNOR U4441 ( .A(in[1279]), .B(n8415), .Z(n8215) );
  NAND U4442 ( .A(n8218), .B(n8215), .Z(n7618) );
  XNOR U4443 ( .A(n7833), .B(n7618), .Z(out[355]) );
  XNOR U4444 ( .A(in[108]), .B(n8790), .Z(n7835) );
  XOR U4445 ( .A(in[1289]), .B(n8665), .Z(n8222) );
  XNOR U4446 ( .A(in[1216]), .B(n8419), .Z(n8219) );
  NAND U4447 ( .A(n8222), .B(n8219), .Z(n7619) );
  XNOR U4448 ( .A(n7835), .B(n7619), .Z(out[356]) );
  XNOR U4449 ( .A(in[109]), .B(n8793), .Z(n7837) );
  XOR U4450 ( .A(in[1290]), .B(n8667), .Z(n8226) );
  XNOR U4451 ( .A(in[1217]), .B(n8423), .Z(n8223) );
  NAND U4452 ( .A(n8226), .B(n8223), .Z(n7620) );
  XNOR U4453 ( .A(n7837), .B(n7620), .Z(out[357]) );
  XNOR U4454 ( .A(in[110]), .B(n8796), .Z(n7839) );
  XOR U4455 ( .A(in[1291]), .B(n8669), .Z(n8230) );
  XNOR U4456 ( .A(in[1218]), .B(n8431), .Z(n8227) );
  NAND U4457 ( .A(n8230), .B(n8227), .Z(n7621) );
  XNOR U4458 ( .A(n7839), .B(n7621), .Z(out[358]) );
  XNOR U4459 ( .A(in[111]), .B(n8799), .Z(n7841) );
  XOR U4460 ( .A(in[1292]), .B(n8671), .Z(n8234) );
  XNOR U4461 ( .A(in[1219]), .B(n8435), .Z(n8231) );
  NAND U4462 ( .A(n8234), .B(n8231), .Z(n7622) );
  XNOR U4463 ( .A(n7841), .B(n7622), .Z(out[359]) );
  OR U4464 ( .A(n9608), .B(n7623), .Z(n7624) );
  XNOR U4465 ( .A(n9607), .B(n7624), .Z(out[35]) );
  XNOR U4466 ( .A(in[112]), .B(n8802), .Z(n7843) );
  XOR U4467 ( .A(in[1293]), .B(n8673), .Z(n8238) );
  XOR U4468 ( .A(in[1220]), .B(n8439), .Z(n8235) );
  NAND U4469 ( .A(n8238), .B(n8235), .Z(n7625) );
  XNOR U4470 ( .A(n7843), .B(n7625), .Z(out[360]) );
  XNOR U4471 ( .A(in[113]), .B(n8805), .Z(n7845) );
  XOR U4472 ( .A(in[1294]), .B(n8675), .Z(n8242) );
  XOR U4473 ( .A(in[1221]), .B(n8443), .Z(n8239) );
  NAND U4474 ( .A(n8242), .B(n8239), .Z(n7626) );
  XNOR U4475 ( .A(n7845), .B(n7626), .Z(out[361]) );
  XNOR U4476 ( .A(in[114]), .B(n8808), .Z(n7851) );
  XOR U4477 ( .A(in[1295]), .B(n8677), .Z(n8246) );
  XOR U4478 ( .A(in[1222]), .B(n8447), .Z(n8243) );
  NAND U4479 ( .A(n8246), .B(n8243), .Z(n7627) );
  XNOR U4480 ( .A(n7851), .B(n7627), .Z(out[362]) );
  XNOR U4481 ( .A(in[115]), .B(n8815), .Z(n7853) );
  XOR U4482 ( .A(in[1296]), .B(n8679), .Z(n8250) );
  XOR U4483 ( .A(in[1223]), .B(n8451), .Z(n8247) );
  NAND U4484 ( .A(n8250), .B(n8247), .Z(n7628) );
  XNOR U4485 ( .A(n7853), .B(n7628), .Z(out[363]) );
  XNOR U4486 ( .A(in[116]), .B(n8818), .Z(n7855) );
  XOR U4487 ( .A(in[1297]), .B(n8681), .Z(n8258) );
  XOR U4488 ( .A(in[1224]), .B(n8455), .Z(n8255) );
  NAND U4489 ( .A(n8258), .B(n8255), .Z(n7629) );
  XNOR U4490 ( .A(n7855), .B(n7629), .Z(out[364]) );
  XNOR U4491 ( .A(in[117]), .B(n8821), .Z(n7857) );
  XOR U4492 ( .A(in[1298]), .B(n8685), .Z(n8262) );
  XOR U4493 ( .A(in[1225]), .B(n8459), .Z(n8259) );
  NAND U4494 ( .A(n8262), .B(n8259), .Z(n7630) );
  XNOR U4495 ( .A(n7857), .B(n7630), .Z(out[365]) );
  XNOR U4496 ( .A(in[118]), .B(n8824), .Z(n7859) );
  XOR U4497 ( .A(in[1299]), .B(n8687), .Z(n8266) );
  XOR U4498 ( .A(in[1226]), .B(n8463), .Z(n8263) );
  NAND U4499 ( .A(n8266), .B(n8263), .Z(n7631) );
  XNOR U4500 ( .A(n7859), .B(n7631), .Z(out[366]) );
  XNOR U4501 ( .A(in[119]), .B(n8827), .Z(n7861) );
  XOR U4502 ( .A(in[1300]), .B(n8689), .Z(n8270) );
  XOR U4503 ( .A(in[1227]), .B(n8467), .Z(n8267) );
  NAND U4504 ( .A(n8270), .B(n8267), .Z(n7632) );
  XNOR U4505 ( .A(n7861), .B(n7632), .Z(out[367]) );
  XNOR U4506 ( .A(in[120]), .B(n8830), .Z(n7863) );
  XOR U4507 ( .A(in[1301]), .B(n8691), .Z(n8274) );
  XOR U4508 ( .A(in[1228]), .B(n8475), .Z(n8271) );
  NAND U4509 ( .A(n8274), .B(n8271), .Z(n7633) );
  XNOR U4510 ( .A(n7863), .B(n7633), .Z(out[368]) );
  XNOR U4511 ( .A(in[121]), .B(n8833), .Z(n7865) );
  XOR U4512 ( .A(in[1302]), .B(n8693), .Z(n8278) );
  XOR U4513 ( .A(in[1229]), .B(n8479), .Z(n8275) );
  NAND U4514 ( .A(n8278), .B(n8275), .Z(n7634) );
  XNOR U4515 ( .A(n7865), .B(n7634), .Z(out[369]) );
  ANDN U4516 ( .B(n7636), .A(n7635), .Z(n7637) );
  XNOR U4517 ( .A(n7638), .B(n7637), .Z(out[36]) );
  XNOR U4518 ( .A(in[122]), .B(n8836), .Z(n7867) );
  XOR U4519 ( .A(in[1303]), .B(n8695), .Z(n8282) );
  XOR U4520 ( .A(in[1230]), .B(n8483), .Z(n8279) );
  NAND U4521 ( .A(n8282), .B(n8279), .Z(n7639) );
  XNOR U4522 ( .A(n7867), .B(n7639), .Z(out[370]) );
  XNOR U4523 ( .A(in[123]), .B(n8839), .Z(n7869) );
  XOR U4524 ( .A(in[1304]), .B(n8697), .Z(n8286) );
  XOR U4525 ( .A(in[1231]), .B(n8487), .Z(n8283) );
  NAND U4526 ( .A(n8286), .B(n8283), .Z(n7640) );
  XNOR U4527 ( .A(n7869), .B(n7640), .Z(out[371]) );
  XNOR U4528 ( .A(in[124]), .B(n8842), .Z(n7877) );
  XOR U4529 ( .A(in[1305]), .B(n8699), .Z(n8290) );
  XOR U4530 ( .A(in[1232]), .B(n8491), .Z(n8287) );
  NAND U4531 ( .A(n8290), .B(n8287), .Z(n7641) );
  XNOR U4532 ( .A(n7877), .B(n7641), .Z(out[372]) );
  XNOR U4533 ( .A(in[125]), .B(n8849), .Z(n7879) );
  XOR U4534 ( .A(in[1306]), .B(n8701), .Z(n8294) );
  XOR U4535 ( .A(in[1233]), .B(n8495), .Z(n8291) );
  NAND U4536 ( .A(n8294), .B(n8291), .Z(n7642) );
  XNOR U4537 ( .A(n7879), .B(n7642), .Z(out[373]) );
  XNOR U4538 ( .A(in[126]), .B(n8852), .Z(n7881) );
  XOR U4539 ( .A(in[1307]), .B(n8703), .Z(n8302) );
  XOR U4540 ( .A(in[1234]), .B(n8499), .Z(n8299) );
  NAND U4541 ( .A(n8302), .B(n8299), .Z(n7643) );
  XNOR U4542 ( .A(n7881), .B(n7643), .Z(out[374]) );
  XNOR U4543 ( .A(in[127]), .B(n8855), .Z(n7883) );
  XOR U4544 ( .A(in[1308]), .B(n8707), .Z(n8306) );
  XOR U4545 ( .A(in[1235]), .B(n8503), .Z(n8303) );
  NAND U4546 ( .A(n8306), .B(n8303), .Z(n7644) );
  XNOR U4547 ( .A(n7883), .B(n7644), .Z(out[375]) );
  XNOR U4548 ( .A(in[64]), .B(n8858), .Z(n7885) );
  XOR U4549 ( .A(in[1309]), .B(n8709), .Z(n8310) );
  XOR U4550 ( .A(in[1236]), .B(n8507), .Z(n8307) );
  NAND U4551 ( .A(n8310), .B(n8307), .Z(n7645) );
  XNOR U4552 ( .A(n7885), .B(n7645), .Z(out[376]) );
  XNOR U4553 ( .A(in[65]), .B(n8861), .Z(n7887) );
  XOR U4554 ( .A(in[1310]), .B(n8711), .Z(n8314) );
  XOR U4555 ( .A(in[1237]), .B(n8511), .Z(n8311) );
  NAND U4556 ( .A(n8314), .B(n8311), .Z(n7646) );
  XNOR U4557 ( .A(n7887), .B(n7646), .Z(out[377]) );
  XNOR U4558 ( .A(in[66]), .B(n8864), .Z(n7889) );
  XOR U4559 ( .A(in[1311]), .B(n8713), .Z(n8318) );
  XOR U4560 ( .A(in[1238]), .B(n8519), .Z(n8315) );
  NAND U4561 ( .A(n8318), .B(n8315), .Z(n7647) );
  XNOR U4562 ( .A(n7889), .B(n7647), .Z(out[378]) );
  XNOR U4563 ( .A(in[67]), .B(n8867), .Z(n7891) );
  XOR U4564 ( .A(in[1312]), .B(n8715), .Z(n8322) );
  XOR U4565 ( .A(in[1239]), .B(n8523), .Z(n8319) );
  NAND U4566 ( .A(n8322), .B(n8319), .Z(n7648) );
  XNOR U4567 ( .A(n7891), .B(n7648), .Z(out[379]) );
  ANDN U4568 ( .B(n7650), .A(n7649), .Z(n7651) );
  XNOR U4569 ( .A(n7652), .B(n7651), .Z(out[37]) );
  XNOR U4570 ( .A(in[68]), .B(n8870), .Z(n7893) );
  XOR U4571 ( .A(in[1313]), .B(n8717), .Z(n8326) );
  XOR U4572 ( .A(in[1240]), .B(n8527), .Z(n8323) );
  NAND U4573 ( .A(n8326), .B(n8323), .Z(n7653) );
  XNOR U4574 ( .A(n7893), .B(n7653), .Z(out[380]) );
  XNOR U4575 ( .A(in[69]), .B(n8873), .Z(n7895) );
  XOR U4576 ( .A(in[1314]), .B(n8719), .Z(n8330) );
  XOR U4577 ( .A(in[1241]), .B(n8531), .Z(n8327) );
  NAND U4578 ( .A(n8330), .B(n8327), .Z(n7654) );
  XNOR U4579 ( .A(n7895), .B(n7654), .Z(out[381]) );
  XNOR U4580 ( .A(in[70]), .B(n8876), .Z(n7901) );
  XOR U4581 ( .A(in[1315]), .B(n8721), .Z(n8334) );
  XOR U4582 ( .A(in[1242]), .B(n8535), .Z(n8331) );
  NAND U4583 ( .A(n8334), .B(n8331), .Z(n7655) );
  XNOR U4584 ( .A(n7901), .B(n7655), .Z(out[382]) );
  XNOR U4585 ( .A(in[71]), .B(n8887), .Z(n7903) );
  XOR U4586 ( .A(in[1316]), .B(n8723), .Z(n8338) );
  XOR U4587 ( .A(in[1243]), .B(n8539), .Z(n8335) );
  NAND U4588 ( .A(n8338), .B(n8335), .Z(n7656) );
  XNOR U4589 ( .A(n7903), .B(n7656), .Z(out[383]) );
  XOR U4590 ( .A(in[497]), .B(n8585), .Z(n7905) );
  NOR U4591 ( .A(n7747), .B(n8060), .Z(n7657) );
  XNOR U4592 ( .A(n7905), .B(n7657), .Z(out[384]) );
  XOR U4593 ( .A(in[498]), .B(n8589), .Z(n7907) );
  NOR U4594 ( .A(n7749), .B(n8064), .Z(n7658) );
  XNOR U4595 ( .A(n7907), .B(n7658), .Z(out[385]) );
  XOR U4596 ( .A(in[499]), .B(n8593), .Z(n7909) );
  NOR U4597 ( .A(n7755), .B(n8068), .Z(n7659) );
  XNOR U4598 ( .A(n7909), .B(n7659), .Z(out[386]) );
  XOR U4599 ( .A(in[500]), .B(n8597), .Z(n7911) );
  NOR U4600 ( .A(n7757), .B(n8072), .Z(n7660) );
  XNOR U4601 ( .A(n7911), .B(n7660), .Z(out[387]) );
  XOR U4602 ( .A(in[501]), .B(n8601), .Z(n7913) );
  NOR U4603 ( .A(n7759), .B(n8080), .Z(n7661) );
  XNOR U4604 ( .A(n7913), .B(n7661), .Z(out[388]) );
  XOR U4605 ( .A(in[502]), .B(n8611), .Z(n7915) );
  NOR U4606 ( .A(n7761), .B(n8084), .Z(n7662) );
  XNOR U4607 ( .A(n7915), .B(n7662), .Z(out[389]) );
  ANDN U4608 ( .B(n7664), .A(n7663), .Z(n7665) );
  XNOR U4609 ( .A(n7666), .B(n7665), .Z(out[38]) );
  XOR U4610 ( .A(in[503]), .B(n8615), .Z(n7917) );
  NOR U4611 ( .A(n7763), .B(n8088), .Z(n7667) );
  XNOR U4612 ( .A(n7917), .B(n7667), .Z(out[390]) );
  XOR U4613 ( .A(in[504]), .B(n8619), .Z(n7919) );
  NOR U4614 ( .A(n7765), .B(n8092), .Z(n7668) );
  XNOR U4615 ( .A(n7919), .B(n7668), .Z(out[391]) );
  XOR U4616 ( .A(in[505]), .B(n8623), .Z(n7925) );
  NOR U4617 ( .A(n7767), .B(n8096), .Z(n7669) );
  XNOR U4618 ( .A(n7925), .B(n7669), .Z(out[392]) );
  XOR U4619 ( .A(in[506]), .B(n8345), .Z(n7927) );
  NOR U4620 ( .A(n7769), .B(n8100), .Z(n7670) );
  XNOR U4621 ( .A(n7927), .B(n7670), .Z(out[393]) );
  XOR U4622 ( .A(in[507]), .B(n8349), .Z(n7929) );
  NOR U4623 ( .A(n7771), .B(n8104), .Z(n7671) );
  XNOR U4624 ( .A(n7929), .B(n7671), .Z(out[394]) );
  XOR U4625 ( .A(in[508]), .B(n8353), .Z(n7931) );
  NOR U4626 ( .A(n7773), .B(n8108), .Z(n7672) );
  XNOR U4627 ( .A(n7931), .B(n7672), .Z(out[395]) );
  XOR U4628 ( .A(in[509]), .B(n8357), .Z(n7933) );
  NOR U4629 ( .A(n7779), .B(n8112), .Z(n7673) );
  XNOR U4630 ( .A(n7933), .B(n7673), .Z(out[396]) );
  XOR U4631 ( .A(in[510]), .B(n8361), .Z(n7935) );
  NOR U4632 ( .A(n7781), .B(n8116), .Z(n7674) );
  XNOR U4633 ( .A(n7935), .B(n7674), .Z(out[397]) );
  XOR U4634 ( .A(in[511]), .B(n8365), .Z(n7937) );
  NOR U4635 ( .A(n7783), .B(n8124), .Z(n7675) );
  XNOR U4636 ( .A(n7937), .B(n7675), .Z(out[398]) );
  XOR U4637 ( .A(in[448]), .B(n8369), .Z(n7939) );
  NOR U4638 ( .A(n7785), .B(n8128), .Z(n7676) );
  XNOR U4639 ( .A(n7939), .B(n7676), .Z(out[399]) );
  ANDN U4640 ( .B(n7678), .A(n7677), .Z(n7679) );
  XNOR U4641 ( .A(n7680), .B(n7679), .Z(out[39]) );
  OR U4642 ( .A(n8516), .B(n7681), .Z(n7682) );
  XNOR U4643 ( .A(n8515), .B(n7682), .Z(out[3]) );
  XOR U4644 ( .A(in[449]), .B(n8373), .Z(n7941) );
  NOR U4645 ( .A(n7787), .B(n8132), .Z(n7683) );
  XNOR U4646 ( .A(n7941), .B(n7683), .Z(out[400]) );
  XNOR U4647 ( .A(n8377), .B(in[450]), .Z(n7943) );
  NOR U4648 ( .A(n7789), .B(n8136), .Z(n7684) );
  XNOR U4649 ( .A(n7943), .B(n7684), .Z(out[401]) );
  XNOR U4650 ( .A(n8381), .B(in[451]), .Z(n7949) );
  NOR U4651 ( .A(n7791), .B(n8140), .Z(n7685) );
  XNOR U4652 ( .A(n7949), .B(n7685), .Z(out[402]) );
  XNOR U4653 ( .A(n8389), .B(in[452]), .Z(n7951) );
  NOR U4654 ( .A(n7793), .B(n8144), .Z(n7686) );
  XNOR U4655 ( .A(n7951), .B(n7686), .Z(out[403]) );
  XNOR U4656 ( .A(n8393), .B(in[453]), .Z(n7953) );
  NOR U4657 ( .A(n7795), .B(n8148), .Z(n7687) );
  XNOR U4658 ( .A(n7953), .B(n7687), .Z(out[404]) );
  XNOR U4659 ( .A(n8397), .B(in[454]), .Z(n7955) );
  NOR U4660 ( .A(n7797), .B(n8152), .Z(n7688) );
  XNOR U4661 ( .A(n7955), .B(n7688), .Z(out[405]) );
  XNOR U4662 ( .A(n8401), .B(in[455]), .Z(n7957) );
  NOR U4663 ( .A(n7803), .B(n8156), .Z(n7689) );
  XNOR U4664 ( .A(n7957), .B(n7689), .Z(out[406]) );
  XNOR U4665 ( .A(n8405), .B(in[456]), .Z(n7959) );
  NOR U4666 ( .A(n7805), .B(n8160), .Z(n7690) );
  XNOR U4667 ( .A(n7959), .B(n7690), .Z(out[407]) );
  XNOR U4668 ( .A(in[457]), .B(n8409), .Z(n7961) );
  NOR U4669 ( .A(n7807), .B(n8170), .Z(n7691) );
  XNOR U4670 ( .A(n7961), .B(n7691), .Z(out[408]) );
  XNOR U4671 ( .A(n8413), .B(in[458]), .Z(n7963) );
  NOR U4672 ( .A(n7809), .B(n8174), .Z(n7692) );
  XNOR U4673 ( .A(n7963), .B(n7692), .Z(out[409]) );
  ANDN U4674 ( .B(n7694), .A(n7693), .Z(n7695) );
  XNOR U4675 ( .A(n7696), .B(n7695), .Z(out[40]) );
  XNOR U4676 ( .A(n8417), .B(in[459]), .Z(n7965) );
  NOR U4677 ( .A(n7811), .B(n8178), .Z(n7697) );
  XNOR U4678 ( .A(n7965), .B(n7697), .Z(out[410]) );
  XNOR U4679 ( .A(in[460]), .B(n8421), .Z(n7967) );
  NOR U4680 ( .A(n7813), .B(n8182), .Z(n7698) );
  XNOR U4681 ( .A(n7967), .B(n7698), .Z(out[411]) );
  XNOR U4682 ( .A(in[461]), .B(n8425), .Z(n7973) );
  NOR U4683 ( .A(n7815), .B(n8186), .Z(n7699) );
  XNOR U4684 ( .A(n7973), .B(n7699), .Z(out[412]) );
  XNOR U4685 ( .A(in[462]), .B(n8433), .Z(n7975) );
  NOR U4686 ( .A(n7817), .B(n8190), .Z(n7700) );
  XNOR U4687 ( .A(n7975), .B(n7700), .Z(out[413]) );
  XNOR U4688 ( .A(in[463]), .B(n8437), .Z(n7977) );
  NOR U4689 ( .A(n7819), .B(n8194), .Z(n7701) );
  XNOR U4690 ( .A(n7977), .B(n7701), .Z(out[414]) );
  XNOR U4691 ( .A(in[464]), .B(n8441), .Z(n7979) );
  NOR U4692 ( .A(n7821), .B(n8198), .Z(n7702) );
  XNOR U4693 ( .A(n7979), .B(n7702), .Z(out[415]) );
  XNOR U4694 ( .A(in[465]), .B(n8445), .Z(n7981) );
  NOR U4695 ( .A(n7827), .B(n8202), .Z(n7703) );
  XNOR U4696 ( .A(n7981), .B(n7703), .Z(out[416]) );
  XNOR U4697 ( .A(in[466]), .B(n8449), .Z(n7983) );
  NOR U4698 ( .A(n7829), .B(n8206), .Z(n7704) );
  XNOR U4699 ( .A(n7983), .B(n7704), .Z(out[417]) );
  XNOR U4700 ( .A(in[467]), .B(n8453), .Z(n7985) );
  NOR U4701 ( .A(n7831), .B(n8214), .Z(n7705) );
  XNOR U4702 ( .A(n7985), .B(n7705), .Z(out[418]) );
  XNOR U4703 ( .A(in[468]), .B(n8457), .Z(n7987) );
  NOR U4704 ( .A(n7833), .B(n8218), .Z(n7706) );
  XNOR U4705 ( .A(n7987), .B(n7706), .Z(out[419]) );
  ANDN U4706 ( .B(n7708), .A(n7707), .Z(n7709) );
  XNOR U4707 ( .A(n7710), .B(n7709), .Z(out[41]) );
  XNOR U4708 ( .A(in[469]), .B(n8461), .Z(n7989) );
  NOR U4709 ( .A(n7835), .B(n8222), .Z(n7711) );
  XNOR U4710 ( .A(n7989), .B(n7711), .Z(out[420]) );
  XNOR U4711 ( .A(in[470]), .B(n8465), .Z(n7991) );
  NOR U4712 ( .A(n7837), .B(n8226), .Z(n7712) );
  XNOR U4713 ( .A(n7991), .B(n7712), .Z(out[421]) );
  XNOR U4714 ( .A(in[471]), .B(n8469), .Z(n7997) );
  NOR U4715 ( .A(n7839), .B(n8230), .Z(n7713) );
  XNOR U4716 ( .A(n7997), .B(n7713), .Z(out[422]) );
  XNOR U4717 ( .A(in[472]), .B(n8477), .Z(n7999) );
  NOR U4718 ( .A(n7841), .B(n8234), .Z(n7714) );
  XNOR U4719 ( .A(n7999), .B(n7714), .Z(out[423]) );
  XNOR U4720 ( .A(in[473]), .B(n8481), .Z(n8001) );
  NOR U4721 ( .A(n7843), .B(n8238), .Z(n7715) );
  XNOR U4722 ( .A(n8001), .B(n7715), .Z(out[424]) );
  XNOR U4723 ( .A(in[474]), .B(n8485), .Z(n8003) );
  NOR U4724 ( .A(n7845), .B(n8242), .Z(n7716) );
  XNOR U4725 ( .A(n8003), .B(n7716), .Z(out[425]) );
  XNOR U4726 ( .A(in[475]), .B(n8489), .Z(n8005) );
  NOR U4727 ( .A(n7851), .B(n8246), .Z(n7717) );
  XNOR U4728 ( .A(n8005), .B(n7717), .Z(out[426]) );
  XNOR U4729 ( .A(in[476]), .B(n8493), .Z(n8007) );
  NOR U4730 ( .A(n7853), .B(n8250), .Z(n7718) );
  XNOR U4731 ( .A(n8007), .B(n7718), .Z(out[427]) );
  XNOR U4732 ( .A(in[477]), .B(n8497), .Z(n8009) );
  NOR U4733 ( .A(n7855), .B(n8258), .Z(n7719) );
  XNOR U4734 ( .A(n8009), .B(n7719), .Z(out[428]) );
  XNOR U4735 ( .A(in[478]), .B(n8501), .Z(n8011) );
  NOR U4736 ( .A(n7857), .B(n8262), .Z(n7720) );
  XNOR U4737 ( .A(n8011), .B(n7720), .Z(out[429]) );
  ANDN U4738 ( .B(n7722), .A(n7721), .Z(n7723) );
  XNOR U4739 ( .A(n7724), .B(n7723), .Z(out[42]) );
  XNOR U4740 ( .A(in[479]), .B(n8505), .Z(n8013) );
  NOR U4741 ( .A(n7859), .B(n8266), .Z(n7725) );
  XNOR U4742 ( .A(n8013), .B(n7725), .Z(out[430]) );
  XNOR U4743 ( .A(in[480]), .B(n8509), .Z(n8015) );
  NOR U4744 ( .A(n7861), .B(n8270), .Z(n7726) );
  XNOR U4745 ( .A(n8015), .B(n7726), .Z(out[431]) );
  XNOR U4746 ( .A(in[481]), .B(n8513), .Z(n8021) );
  NOR U4747 ( .A(n7863), .B(n8274), .Z(n7727) );
  XNOR U4748 ( .A(n8021), .B(n7727), .Z(out[432]) );
  XNOR U4749 ( .A(in[482]), .B(n8521), .Z(n8023) );
  NOR U4750 ( .A(n7865), .B(n8278), .Z(n7728) );
  XNOR U4751 ( .A(n8023), .B(n7728), .Z(out[433]) );
  XNOR U4752 ( .A(in[483]), .B(n8525), .Z(n8025) );
  NOR U4753 ( .A(n7867), .B(n8282), .Z(n7729) );
  XNOR U4754 ( .A(n8025), .B(n7729), .Z(out[434]) );
  XNOR U4755 ( .A(in[484]), .B(n8529), .Z(n8027) );
  NOR U4756 ( .A(n7869), .B(n8286), .Z(n7730) );
  XNOR U4757 ( .A(n8027), .B(n7730), .Z(out[435]) );
  XNOR U4758 ( .A(in[485]), .B(n8533), .Z(n8029) );
  NOR U4759 ( .A(n7877), .B(n8290), .Z(n7731) );
  XNOR U4760 ( .A(n8029), .B(n7731), .Z(out[436]) );
  XOR U4761 ( .A(in[486]), .B(n8537), .Z(n8031) );
  NOR U4762 ( .A(n7879), .B(n8294), .Z(n7732) );
  XNOR U4763 ( .A(n8031), .B(n7732), .Z(out[437]) );
  XOR U4764 ( .A(in[487]), .B(n8541), .Z(n8033) );
  NOR U4765 ( .A(n7881), .B(n8302), .Z(n7733) );
  XNOR U4766 ( .A(n8033), .B(n7733), .Z(out[438]) );
  XOR U4767 ( .A(in[488]), .B(n8545), .Z(n8035) );
  NOR U4768 ( .A(n7883), .B(n8306), .Z(n7734) );
  XNOR U4769 ( .A(n8035), .B(n7734), .Z(out[439]) );
  ANDN U4770 ( .B(n7736), .A(n7735), .Z(n7737) );
  XNOR U4771 ( .A(n7738), .B(n7737), .Z(out[43]) );
  XOR U4772 ( .A(in[489]), .B(n8549), .Z(n8037) );
  NOR U4773 ( .A(n7885), .B(n8310), .Z(n7739) );
  XNOR U4774 ( .A(n8037), .B(n7739), .Z(out[440]) );
  XOR U4775 ( .A(in[490]), .B(n8553), .Z(n8039) );
  NOR U4776 ( .A(n7887), .B(n8314), .Z(n7740) );
  XNOR U4777 ( .A(n8039), .B(n7740), .Z(out[441]) );
  XOR U4778 ( .A(in[491]), .B(n8557), .Z(n8045) );
  NOR U4779 ( .A(n7889), .B(n8318), .Z(n7741) );
  XNOR U4780 ( .A(n8045), .B(n7741), .Z(out[442]) );
  XOR U4781 ( .A(in[492]), .B(n8565), .Z(n8047) );
  NOR U4782 ( .A(n7891), .B(n8322), .Z(n7742) );
  XNOR U4783 ( .A(n8047), .B(n7742), .Z(out[443]) );
  XOR U4784 ( .A(in[493]), .B(n8569), .Z(n8049) );
  NOR U4785 ( .A(n7893), .B(n8326), .Z(n7743) );
  XNOR U4786 ( .A(n8049), .B(n7743), .Z(out[444]) );
  XOR U4787 ( .A(in[494]), .B(n8573), .Z(n8051) );
  NOR U4788 ( .A(n7895), .B(n8330), .Z(n7744) );
  XNOR U4789 ( .A(n8051), .B(n7744), .Z(out[445]) );
  XOR U4790 ( .A(in[495]), .B(n8577), .Z(n8053) );
  NOR U4791 ( .A(n7901), .B(n8334), .Z(n7745) );
  XNOR U4792 ( .A(n8053), .B(n7745), .Z(out[446]) );
  XOR U4793 ( .A(in[496]), .B(n8581), .Z(n8055) );
  NOR U4794 ( .A(n7903), .B(n8338), .Z(n7746) );
  XNOR U4795 ( .A(n8055), .B(n7746), .Z(out[447]) );
  XNOR U4796 ( .A(in[886]), .B(n8584), .Z(n8058) );
  NAND U4797 ( .A(n7905), .B(n7747), .Z(n7748) );
  XNOR U4798 ( .A(n8058), .B(n7748), .Z(out[448]) );
  XNOR U4799 ( .A(in[887]), .B(n8588), .Z(n8062) );
  NAND U4800 ( .A(n7907), .B(n7749), .Z(n7750) );
  XNOR U4801 ( .A(n8062), .B(n7750), .Z(out[449]) );
  ANDN U4802 ( .B(n7752), .A(n7751), .Z(n7753) );
  XNOR U4803 ( .A(n7754), .B(n7753), .Z(out[44]) );
  XNOR U4804 ( .A(in[888]), .B(n8592), .Z(n8066) );
  NAND U4805 ( .A(n7909), .B(n7755), .Z(n7756) );
  XNOR U4806 ( .A(n8066), .B(n7756), .Z(out[450]) );
  XNOR U4807 ( .A(in[889]), .B(n8596), .Z(n8070) );
  NAND U4808 ( .A(n7911), .B(n7757), .Z(n7758) );
  XNOR U4809 ( .A(n8070), .B(n7758), .Z(out[451]) );
  XNOR U4810 ( .A(in[890]), .B(n8600), .Z(n8078) );
  NAND U4811 ( .A(n7913), .B(n7759), .Z(n7760) );
  XNOR U4812 ( .A(n8078), .B(n7760), .Z(out[452]) );
  XOR U4813 ( .A(in[891]), .B(n8610), .Z(n8082) );
  NAND U4814 ( .A(n7915), .B(n7761), .Z(n7762) );
  XNOR U4815 ( .A(n8082), .B(n7762), .Z(out[453]) );
  XOR U4816 ( .A(in[892]), .B(n8614), .Z(n8086) );
  NAND U4817 ( .A(n7917), .B(n7763), .Z(n7764) );
  XNOR U4818 ( .A(n8086), .B(n7764), .Z(out[454]) );
  XOR U4819 ( .A(in[893]), .B(n8618), .Z(n8090) );
  NAND U4820 ( .A(n7919), .B(n7765), .Z(n7766) );
  XNOR U4821 ( .A(n8090), .B(n7766), .Z(out[455]) );
  XNOR U4822 ( .A(in[894]), .B(n8622), .Z(n8094) );
  NAND U4823 ( .A(n7925), .B(n7767), .Z(n7768) );
  XNOR U4824 ( .A(n8094), .B(n7768), .Z(out[456]) );
  XOR U4825 ( .A(in[895]), .B(n8344), .Z(n8098) );
  NAND U4826 ( .A(n7927), .B(n7769), .Z(n7770) );
  XNOR U4827 ( .A(n8098), .B(n7770), .Z(out[457]) );
  XOR U4828 ( .A(in[832]), .B(n8348), .Z(n8102) );
  NAND U4829 ( .A(n7929), .B(n7771), .Z(n7772) );
  XNOR U4830 ( .A(n8102), .B(n7772), .Z(out[458]) );
  XOR U4831 ( .A(in[833]), .B(n8352), .Z(n8106) );
  NAND U4832 ( .A(n7931), .B(n7773), .Z(n7774) );
  XNOR U4833 ( .A(n8106), .B(n7774), .Z(out[459]) );
  ANDN U4834 ( .B(n7776), .A(n7775), .Z(n7777) );
  XNOR U4835 ( .A(n7778), .B(n7777), .Z(out[45]) );
  XOR U4836 ( .A(in[834]), .B(n8356), .Z(n8110) );
  NAND U4837 ( .A(n7933), .B(n7779), .Z(n7780) );
  XNOR U4838 ( .A(n8110), .B(n7780), .Z(out[460]) );
  XOR U4839 ( .A(in[835]), .B(n8360), .Z(n8114) );
  NAND U4840 ( .A(n7935), .B(n7781), .Z(n7782) );
  XNOR U4841 ( .A(n8114), .B(n7782), .Z(out[461]) );
  XOR U4842 ( .A(in[836]), .B(n8364), .Z(n8122) );
  NAND U4843 ( .A(n7937), .B(n7783), .Z(n7784) );
  XNOR U4844 ( .A(n8122), .B(n7784), .Z(out[462]) );
  XOR U4845 ( .A(in[837]), .B(n8368), .Z(n8126) );
  NAND U4846 ( .A(n7939), .B(n7785), .Z(n7786) );
  XNOR U4847 ( .A(n8126), .B(n7786), .Z(out[463]) );
  XOR U4848 ( .A(in[838]), .B(n8372), .Z(n8130) );
  NAND U4849 ( .A(n7941), .B(n7787), .Z(n7788) );
  XNOR U4850 ( .A(n8130), .B(n7788), .Z(out[464]) );
  XOR U4851 ( .A(in[839]), .B(n8376), .Z(n8134) );
  NAND U4852 ( .A(n7943), .B(n7789), .Z(n7790) );
  XNOR U4853 ( .A(n8134), .B(n7790), .Z(out[465]) );
  XOR U4854 ( .A(in[840]), .B(n8380), .Z(n8138) );
  NAND U4855 ( .A(n7949), .B(n7791), .Z(n7792) );
  XNOR U4856 ( .A(n8138), .B(n7792), .Z(out[466]) );
  XOR U4857 ( .A(in[841]), .B(n8388), .Z(n8142) );
  NAND U4858 ( .A(n7951), .B(n7793), .Z(n7794) );
  XNOR U4859 ( .A(n8142), .B(n7794), .Z(out[467]) );
  XOR U4860 ( .A(in[842]), .B(n8392), .Z(n8146) );
  NAND U4861 ( .A(n7953), .B(n7795), .Z(n7796) );
  XNOR U4862 ( .A(n8146), .B(n7796), .Z(out[468]) );
  XOR U4863 ( .A(in[843]), .B(n8396), .Z(n8150) );
  NAND U4864 ( .A(n7955), .B(n7797), .Z(n7798) );
  XNOR U4865 ( .A(n8150), .B(n7798), .Z(out[469]) );
  ANDN U4866 ( .B(n7800), .A(n7799), .Z(n7801) );
  XNOR U4867 ( .A(n7802), .B(n7801), .Z(out[46]) );
  XOR U4868 ( .A(in[844]), .B(n8400), .Z(n8154) );
  NAND U4869 ( .A(n7957), .B(n7803), .Z(n7804) );
  XNOR U4870 ( .A(n8154), .B(n7804), .Z(out[470]) );
  XOR U4871 ( .A(in[845]), .B(n8404), .Z(n8158) );
  NAND U4872 ( .A(n7959), .B(n7805), .Z(n7806) );
  XNOR U4873 ( .A(n8158), .B(n7806), .Z(out[471]) );
  XOR U4874 ( .A(in[846]), .B(n8408), .Z(n8168) );
  NAND U4875 ( .A(n7961), .B(n7807), .Z(n7808) );
  XNOR U4876 ( .A(n8168), .B(n7808), .Z(out[472]) );
  XOR U4877 ( .A(in[847]), .B(n8412), .Z(n8172) );
  NAND U4878 ( .A(n7963), .B(n7809), .Z(n7810) );
  XNOR U4879 ( .A(n8172), .B(n7810), .Z(out[473]) );
  XOR U4880 ( .A(in[848]), .B(n8416), .Z(n8176) );
  NAND U4881 ( .A(n7965), .B(n7811), .Z(n7812) );
  XNOR U4882 ( .A(n8176), .B(n7812), .Z(out[474]) );
  XOR U4883 ( .A(in[849]), .B(n8420), .Z(n8180) );
  NAND U4884 ( .A(n7967), .B(n7813), .Z(n7814) );
  XNOR U4885 ( .A(n8180), .B(n7814), .Z(out[475]) );
  XOR U4886 ( .A(in[850]), .B(n8424), .Z(n8184) );
  NAND U4887 ( .A(n7973), .B(n7815), .Z(n7816) );
  XNOR U4888 ( .A(n8184), .B(n7816), .Z(out[476]) );
  XNOR U4889 ( .A(in[851]), .B(n8432), .Z(n8188) );
  NAND U4890 ( .A(n7975), .B(n7817), .Z(n7818) );
  XNOR U4891 ( .A(n8188), .B(n7818), .Z(out[477]) );
  XNOR U4892 ( .A(in[852]), .B(n8436), .Z(n8192) );
  NAND U4893 ( .A(n7977), .B(n7819), .Z(n7820) );
  XNOR U4894 ( .A(n8192), .B(n7820), .Z(out[478]) );
  XNOR U4895 ( .A(in[853]), .B(n8440), .Z(n8196) );
  NAND U4896 ( .A(n7979), .B(n7821), .Z(n7822) );
  XNOR U4897 ( .A(n8196), .B(n7822), .Z(out[479]) );
  ANDN U4898 ( .B(n7824), .A(n7823), .Z(n7825) );
  XNOR U4899 ( .A(n7826), .B(n7825), .Z(out[47]) );
  XNOR U4900 ( .A(in[854]), .B(n8444), .Z(n8200) );
  NAND U4901 ( .A(n7981), .B(n7827), .Z(n7828) );
  XNOR U4902 ( .A(n8200), .B(n7828), .Z(out[480]) );
  XNOR U4903 ( .A(in[855]), .B(n8448), .Z(n8204) );
  NAND U4904 ( .A(n7983), .B(n7829), .Z(n7830) );
  XNOR U4905 ( .A(n8204), .B(n7830), .Z(out[481]) );
  XNOR U4906 ( .A(in[856]), .B(n8452), .Z(n8212) );
  NAND U4907 ( .A(n7985), .B(n7831), .Z(n7832) );
  XNOR U4908 ( .A(n8212), .B(n7832), .Z(out[482]) );
  XNOR U4909 ( .A(in[857]), .B(n8456), .Z(n8216) );
  NAND U4910 ( .A(n7987), .B(n7833), .Z(n7834) );
  XNOR U4911 ( .A(n8216), .B(n7834), .Z(out[483]) );
  XNOR U4912 ( .A(in[858]), .B(n8460), .Z(n8220) );
  NAND U4913 ( .A(n7989), .B(n7835), .Z(n7836) );
  XNOR U4914 ( .A(n8220), .B(n7836), .Z(out[484]) );
  XNOR U4915 ( .A(in[859]), .B(n8464), .Z(n8224) );
  NAND U4916 ( .A(n7991), .B(n7837), .Z(n7838) );
  XNOR U4917 ( .A(n8224), .B(n7838), .Z(out[485]) );
  XNOR U4918 ( .A(in[860]), .B(n8468), .Z(n8228) );
  NAND U4919 ( .A(n7997), .B(n7839), .Z(n7840) );
  XNOR U4920 ( .A(n8228), .B(n7840), .Z(out[486]) );
  XNOR U4921 ( .A(in[861]), .B(n8476), .Z(n8232) );
  NAND U4922 ( .A(n7999), .B(n7841), .Z(n7842) );
  XNOR U4923 ( .A(n8232), .B(n7842), .Z(out[487]) );
  XNOR U4924 ( .A(in[862]), .B(n8480), .Z(n8236) );
  NAND U4925 ( .A(n8001), .B(n7843), .Z(n7844) );
  XNOR U4926 ( .A(n8236), .B(n7844), .Z(out[488]) );
  XNOR U4927 ( .A(in[863]), .B(n8484), .Z(n8240) );
  NAND U4928 ( .A(n8003), .B(n7845), .Z(n7846) );
  XNOR U4929 ( .A(n8240), .B(n7846), .Z(out[489]) );
  ANDN U4930 ( .B(n7848), .A(n7847), .Z(n7849) );
  XNOR U4931 ( .A(n7850), .B(n7849), .Z(out[48]) );
  XNOR U4932 ( .A(in[864]), .B(n8488), .Z(n8244) );
  NAND U4933 ( .A(n8005), .B(n7851), .Z(n7852) );
  XNOR U4934 ( .A(n8244), .B(n7852), .Z(out[490]) );
  XNOR U4935 ( .A(in[865]), .B(n8492), .Z(n8248) );
  NAND U4936 ( .A(n8007), .B(n7853), .Z(n7854) );
  XNOR U4937 ( .A(n8248), .B(n7854), .Z(out[491]) );
  XOR U4938 ( .A(n8496), .B(in[866]), .Z(n8256) );
  NAND U4939 ( .A(n8009), .B(n7855), .Z(n7856) );
  XNOR U4940 ( .A(n8256), .B(n7856), .Z(out[492]) );
  XOR U4941 ( .A(n8500), .B(in[867]), .Z(n8260) );
  NAND U4942 ( .A(n8011), .B(n7857), .Z(n7858) );
  XNOR U4943 ( .A(n8260), .B(n7858), .Z(out[493]) );
  XOR U4944 ( .A(n8504), .B(in[868]), .Z(n8264) );
  NAND U4945 ( .A(n8013), .B(n7859), .Z(n7860) );
  XNOR U4946 ( .A(n8264), .B(n7860), .Z(out[494]) );
  XOR U4947 ( .A(n8508), .B(in[869]), .Z(n8268) );
  NAND U4948 ( .A(n8015), .B(n7861), .Z(n7862) );
  XNOR U4949 ( .A(n8268), .B(n7862), .Z(out[495]) );
  XNOR U4950 ( .A(in[870]), .B(n8512), .Z(n8272) );
  NAND U4951 ( .A(n8021), .B(n7863), .Z(n7864) );
  XNOR U4952 ( .A(n8272), .B(n7864), .Z(out[496]) );
  XNOR U4953 ( .A(in[871]), .B(n8520), .Z(n8276) );
  NAND U4954 ( .A(n8023), .B(n7865), .Z(n7866) );
  XNOR U4955 ( .A(n8276), .B(n7866), .Z(out[497]) );
  XNOR U4956 ( .A(in[872]), .B(n8524), .Z(n8280) );
  NAND U4957 ( .A(n8025), .B(n7867), .Z(n7868) );
  XNOR U4958 ( .A(n8280), .B(n7868), .Z(out[498]) );
  XNOR U4959 ( .A(in[873]), .B(n8528), .Z(n8284) );
  NAND U4960 ( .A(n8027), .B(n7869), .Z(n7870) );
  XNOR U4961 ( .A(n8284), .B(n7870), .Z(out[499]) );
  ANDN U4962 ( .B(n7872), .A(n7871), .Z(n7873) );
  XNOR U4963 ( .A(n7874), .B(n7873), .Z(out[49]) );
  OR U4964 ( .A(n8560), .B(n7875), .Z(n7876) );
  XNOR U4965 ( .A(n8559), .B(n7876), .Z(out[4]) );
  XNOR U4966 ( .A(in[874]), .B(n8532), .Z(n8288) );
  NAND U4967 ( .A(n8029), .B(n7877), .Z(n7878) );
  XNOR U4968 ( .A(n8288), .B(n7878), .Z(out[500]) );
  XNOR U4969 ( .A(in[875]), .B(n8536), .Z(n8292) );
  NAND U4970 ( .A(n8031), .B(n7879), .Z(n7880) );
  XNOR U4971 ( .A(n8292), .B(n7880), .Z(out[501]) );
  XNOR U4972 ( .A(in[876]), .B(n8540), .Z(n8300) );
  NAND U4973 ( .A(n8033), .B(n7881), .Z(n7882) );
  XNOR U4974 ( .A(n8300), .B(n7882), .Z(out[502]) );
  XNOR U4975 ( .A(in[877]), .B(n8544), .Z(n8304) );
  NAND U4976 ( .A(n8035), .B(n7883), .Z(n7884) );
  XNOR U4977 ( .A(n8304), .B(n7884), .Z(out[503]) );
  XNOR U4978 ( .A(in[878]), .B(n8548), .Z(n8308) );
  NAND U4979 ( .A(n8037), .B(n7885), .Z(n7886) );
  XNOR U4980 ( .A(n8308), .B(n7886), .Z(out[504]) );
  XNOR U4981 ( .A(in[879]), .B(n8552), .Z(n8312) );
  NAND U4982 ( .A(n8039), .B(n7887), .Z(n7888) );
  XNOR U4983 ( .A(n8312), .B(n7888), .Z(out[505]) );
  XNOR U4984 ( .A(in[880]), .B(n8556), .Z(n8316) );
  NAND U4985 ( .A(n8045), .B(n7889), .Z(n7890) );
  XNOR U4986 ( .A(n8316), .B(n7890), .Z(out[506]) );
  XNOR U4987 ( .A(in[881]), .B(n8564), .Z(n8320) );
  NAND U4988 ( .A(n8047), .B(n7891), .Z(n7892) );
  XNOR U4989 ( .A(n8320), .B(n7892), .Z(out[507]) );
  XNOR U4990 ( .A(in[882]), .B(n8568), .Z(n8324) );
  NAND U4991 ( .A(n8049), .B(n7893), .Z(n7894) );
  XNOR U4992 ( .A(n8324), .B(n7894), .Z(out[508]) );
  XNOR U4993 ( .A(in[883]), .B(n8572), .Z(n8328) );
  NAND U4994 ( .A(n8051), .B(n7895), .Z(n7896) );
  XNOR U4995 ( .A(n8328), .B(n7896), .Z(out[509]) );
  ANDN U4996 ( .B(n7898), .A(n7897), .Z(n7899) );
  XNOR U4997 ( .A(n7900), .B(n7899), .Z(out[50]) );
  XNOR U4998 ( .A(in[884]), .B(n8576), .Z(n8332) );
  NAND U4999 ( .A(n8053), .B(n7901), .Z(n7902) );
  XNOR U5000 ( .A(n8332), .B(n7902), .Z(out[510]) );
  XNOR U5001 ( .A(in[885]), .B(n8580), .Z(n8336) );
  NAND U5002 ( .A(n8055), .B(n7903), .Z(n7904) );
  XNOR U5003 ( .A(n8336), .B(n7904), .Z(out[511]) );
  OR U5004 ( .A(n8058), .B(n7905), .Z(n7906) );
  XNOR U5005 ( .A(n8057), .B(n7906), .Z(out[512]) );
  OR U5006 ( .A(n8062), .B(n7907), .Z(n7908) );
  XNOR U5007 ( .A(n8061), .B(n7908), .Z(out[513]) );
  OR U5008 ( .A(n8066), .B(n7909), .Z(n7910) );
  XNOR U5009 ( .A(n8065), .B(n7910), .Z(out[514]) );
  OR U5010 ( .A(n8070), .B(n7911), .Z(n7912) );
  XNOR U5011 ( .A(n8069), .B(n7912), .Z(out[515]) );
  OR U5012 ( .A(n8078), .B(n7913), .Z(n7914) );
  XNOR U5013 ( .A(n8077), .B(n7914), .Z(out[516]) );
  OR U5014 ( .A(n8082), .B(n7915), .Z(n7916) );
  XNOR U5015 ( .A(n8081), .B(n7916), .Z(out[517]) );
  OR U5016 ( .A(n8086), .B(n7917), .Z(n7918) );
  XNOR U5017 ( .A(n8085), .B(n7918), .Z(out[518]) );
  OR U5018 ( .A(n8090), .B(n7919), .Z(n7920) );
  XNOR U5019 ( .A(n8089), .B(n7920), .Z(out[519]) );
  ANDN U5020 ( .B(n7922), .A(n7921), .Z(n7923) );
  XNOR U5021 ( .A(n7924), .B(n7923), .Z(out[51]) );
  OR U5022 ( .A(n8094), .B(n7925), .Z(n7926) );
  XNOR U5023 ( .A(n8093), .B(n7926), .Z(out[520]) );
  OR U5024 ( .A(n8098), .B(n7927), .Z(n7928) );
  XNOR U5025 ( .A(n8097), .B(n7928), .Z(out[521]) );
  OR U5026 ( .A(n8102), .B(n7929), .Z(n7930) );
  XNOR U5027 ( .A(n8101), .B(n7930), .Z(out[522]) );
  OR U5028 ( .A(n8106), .B(n7931), .Z(n7932) );
  XNOR U5029 ( .A(n8105), .B(n7932), .Z(out[523]) );
  OR U5030 ( .A(n8110), .B(n7933), .Z(n7934) );
  XNOR U5031 ( .A(n8109), .B(n7934), .Z(out[524]) );
  OR U5032 ( .A(n8114), .B(n7935), .Z(n7936) );
  XNOR U5033 ( .A(n8113), .B(n7936), .Z(out[525]) );
  OR U5034 ( .A(n8122), .B(n7937), .Z(n7938) );
  XNOR U5035 ( .A(n8121), .B(n7938), .Z(out[526]) );
  OR U5036 ( .A(n8126), .B(n7939), .Z(n7940) );
  XNOR U5037 ( .A(n8125), .B(n7940), .Z(out[527]) );
  OR U5038 ( .A(n8130), .B(n7941), .Z(n7942) );
  XNOR U5039 ( .A(n8129), .B(n7942), .Z(out[528]) );
  OR U5040 ( .A(n8134), .B(n7943), .Z(n7944) );
  XNOR U5041 ( .A(n8133), .B(n7944), .Z(out[529]) );
  ANDN U5042 ( .B(n7946), .A(n7945), .Z(n7947) );
  XNOR U5043 ( .A(n7948), .B(n7947), .Z(out[52]) );
  OR U5044 ( .A(n8138), .B(n7949), .Z(n7950) );
  XNOR U5045 ( .A(n8137), .B(n7950), .Z(out[530]) );
  OR U5046 ( .A(n8142), .B(n7951), .Z(n7952) );
  XNOR U5047 ( .A(n8141), .B(n7952), .Z(out[531]) );
  OR U5048 ( .A(n8146), .B(n7953), .Z(n7954) );
  XNOR U5049 ( .A(n8145), .B(n7954), .Z(out[532]) );
  OR U5050 ( .A(n8150), .B(n7955), .Z(n7956) );
  XNOR U5051 ( .A(n8149), .B(n7956), .Z(out[533]) );
  OR U5052 ( .A(n8154), .B(n7957), .Z(n7958) );
  XNOR U5053 ( .A(n8153), .B(n7958), .Z(out[534]) );
  OR U5054 ( .A(n8158), .B(n7959), .Z(n7960) );
  XNOR U5055 ( .A(n8157), .B(n7960), .Z(out[535]) );
  OR U5056 ( .A(n8168), .B(n7961), .Z(n7962) );
  XNOR U5057 ( .A(n8167), .B(n7962), .Z(out[536]) );
  OR U5058 ( .A(n8172), .B(n7963), .Z(n7964) );
  XNOR U5059 ( .A(n8171), .B(n7964), .Z(out[537]) );
  OR U5060 ( .A(n8176), .B(n7965), .Z(n7966) );
  XNOR U5061 ( .A(n8175), .B(n7966), .Z(out[538]) );
  OR U5062 ( .A(n8180), .B(n7967), .Z(n7968) );
  XNOR U5063 ( .A(n8179), .B(n7968), .Z(out[539]) );
  ANDN U5064 ( .B(n7970), .A(n7969), .Z(n7971) );
  XNOR U5065 ( .A(n7972), .B(n7971), .Z(out[53]) );
  OR U5066 ( .A(n8184), .B(n7973), .Z(n7974) );
  XNOR U5067 ( .A(n8183), .B(n7974), .Z(out[540]) );
  OR U5068 ( .A(n8188), .B(n7975), .Z(n7976) );
  XNOR U5069 ( .A(n8187), .B(n7976), .Z(out[541]) );
  OR U5070 ( .A(n8192), .B(n7977), .Z(n7978) );
  XNOR U5071 ( .A(n8191), .B(n7978), .Z(out[542]) );
  OR U5072 ( .A(n8196), .B(n7979), .Z(n7980) );
  XNOR U5073 ( .A(n8195), .B(n7980), .Z(out[543]) );
  OR U5074 ( .A(n8200), .B(n7981), .Z(n7982) );
  XNOR U5075 ( .A(n8199), .B(n7982), .Z(out[544]) );
  OR U5076 ( .A(n8204), .B(n7983), .Z(n7984) );
  XNOR U5077 ( .A(n8203), .B(n7984), .Z(out[545]) );
  OR U5078 ( .A(n8212), .B(n7985), .Z(n7986) );
  XNOR U5079 ( .A(n8211), .B(n7986), .Z(out[546]) );
  OR U5080 ( .A(n8216), .B(n7987), .Z(n7988) );
  XNOR U5081 ( .A(n8215), .B(n7988), .Z(out[547]) );
  OR U5082 ( .A(n8220), .B(n7989), .Z(n7990) );
  XNOR U5083 ( .A(n8219), .B(n7990), .Z(out[548]) );
  OR U5084 ( .A(n8224), .B(n7991), .Z(n7992) );
  XNOR U5085 ( .A(n8223), .B(n7992), .Z(out[549]) );
  ANDN U5086 ( .B(n7994), .A(n7993), .Z(n7995) );
  XNOR U5087 ( .A(n7996), .B(n7995), .Z(out[54]) );
  OR U5088 ( .A(n8228), .B(n7997), .Z(n7998) );
  XNOR U5089 ( .A(n8227), .B(n7998), .Z(out[550]) );
  OR U5090 ( .A(n8232), .B(n7999), .Z(n8000) );
  XNOR U5091 ( .A(n8231), .B(n8000), .Z(out[551]) );
  OR U5092 ( .A(n8236), .B(n8001), .Z(n8002) );
  XNOR U5093 ( .A(n8235), .B(n8002), .Z(out[552]) );
  OR U5094 ( .A(n8240), .B(n8003), .Z(n8004) );
  XNOR U5095 ( .A(n8239), .B(n8004), .Z(out[553]) );
  OR U5096 ( .A(n8244), .B(n8005), .Z(n8006) );
  XNOR U5097 ( .A(n8243), .B(n8006), .Z(out[554]) );
  OR U5098 ( .A(n8248), .B(n8007), .Z(n8008) );
  XNOR U5099 ( .A(n8247), .B(n8008), .Z(out[555]) );
  OR U5100 ( .A(n8256), .B(n8009), .Z(n8010) );
  XNOR U5101 ( .A(n8255), .B(n8010), .Z(out[556]) );
  OR U5102 ( .A(n8260), .B(n8011), .Z(n8012) );
  XNOR U5103 ( .A(n8259), .B(n8012), .Z(out[557]) );
  OR U5104 ( .A(n8264), .B(n8013), .Z(n8014) );
  XNOR U5105 ( .A(n8263), .B(n8014), .Z(out[558]) );
  OR U5106 ( .A(n8268), .B(n8015), .Z(n8016) );
  XNOR U5107 ( .A(n8267), .B(n8016), .Z(out[559]) );
  ANDN U5108 ( .B(n8018), .A(n8017), .Z(n8019) );
  XNOR U5109 ( .A(n8020), .B(n8019), .Z(out[55]) );
  OR U5110 ( .A(n8272), .B(n8021), .Z(n8022) );
  XNOR U5111 ( .A(n8271), .B(n8022), .Z(out[560]) );
  OR U5112 ( .A(n8276), .B(n8023), .Z(n8024) );
  XNOR U5113 ( .A(n8275), .B(n8024), .Z(out[561]) );
  OR U5114 ( .A(n8280), .B(n8025), .Z(n8026) );
  XNOR U5115 ( .A(n8279), .B(n8026), .Z(out[562]) );
  OR U5116 ( .A(n8284), .B(n8027), .Z(n8028) );
  XNOR U5117 ( .A(n8283), .B(n8028), .Z(out[563]) );
  OR U5118 ( .A(n8288), .B(n8029), .Z(n8030) );
  XNOR U5119 ( .A(n8287), .B(n8030), .Z(out[564]) );
  OR U5120 ( .A(n8292), .B(n8031), .Z(n8032) );
  XNOR U5121 ( .A(n8291), .B(n8032), .Z(out[565]) );
  OR U5122 ( .A(n8300), .B(n8033), .Z(n8034) );
  XNOR U5123 ( .A(n8299), .B(n8034), .Z(out[566]) );
  OR U5124 ( .A(n8304), .B(n8035), .Z(n8036) );
  XNOR U5125 ( .A(n8303), .B(n8036), .Z(out[567]) );
  OR U5126 ( .A(n8308), .B(n8037), .Z(n8038) );
  XNOR U5127 ( .A(n8307), .B(n8038), .Z(out[568]) );
  OR U5128 ( .A(n8312), .B(n8039), .Z(n8040) );
  XNOR U5129 ( .A(n8311), .B(n8040), .Z(out[569]) );
  ANDN U5130 ( .B(n8042), .A(n8041), .Z(n8043) );
  XNOR U5131 ( .A(n8044), .B(n8043), .Z(out[56]) );
  OR U5132 ( .A(n8316), .B(n8045), .Z(n8046) );
  XNOR U5133 ( .A(n8315), .B(n8046), .Z(out[570]) );
  OR U5134 ( .A(n8320), .B(n8047), .Z(n8048) );
  XNOR U5135 ( .A(n8319), .B(n8048), .Z(out[571]) );
  OR U5136 ( .A(n8324), .B(n8049), .Z(n8050) );
  XNOR U5137 ( .A(n8323), .B(n8050), .Z(out[572]) );
  OR U5138 ( .A(n8328), .B(n8051), .Z(n8052) );
  XNOR U5139 ( .A(n8327), .B(n8052), .Z(out[573]) );
  OR U5140 ( .A(n8332), .B(n8053), .Z(n8054) );
  XNOR U5141 ( .A(n8331), .B(n8054), .Z(out[574]) );
  OR U5142 ( .A(n8336), .B(n8055), .Z(n8056) );
  XNOR U5143 ( .A(n8335), .B(n8056), .Z(out[575]) );
  ANDN U5144 ( .B(n8058), .A(n8057), .Z(n8059) );
  XNOR U5145 ( .A(n8060), .B(n8059), .Z(out[576]) );
  ANDN U5146 ( .B(n8062), .A(n8061), .Z(n8063) );
  XNOR U5147 ( .A(n8064), .B(n8063), .Z(out[577]) );
  ANDN U5148 ( .B(n8066), .A(n8065), .Z(n8067) );
  XNOR U5149 ( .A(n8068), .B(n8067), .Z(out[578]) );
  ANDN U5150 ( .B(n8070), .A(n8069), .Z(n8071) );
  XNOR U5151 ( .A(n8072), .B(n8071), .Z(out[579]) );
  ANDN U5152 ( .B(n8074), .A(n8073), .Z(n8075) );
  XNOR U5153 ( .A(n8076), .B(n8075), .Z(out[57]) );
  ANDN U5154 ( .B(n8078), .A(n8077), .Z(n8079) );
  XNOR U5155 ( .A(n8080), .B(n8079), .Z(out[580]) );
  ANDN U5156 ( .B(n8082), .A(n8081), .Z(n8083) );
  XNOR U5157 ( .A(n8084), .B(n8083), .Z(out[581]) );
  ANDN U5158 ( .B(n8086), .A(n8085), .Z(n8087) );
  XNOR U5159 ( .A(n8088), .B(n8087), .Z(out[582]) );
  ANDN U5160 ( .B(n8090), .A(n8089), .Z(n8091) );
  XNOR U5161 ( .A(n8092), .B(n8091), .Z(out[583]) );
  ANDN U5162 ( .B(n8094), .A(n8093), .Z(n8095) );
  XNOR U5163 ( .A(n8096), .B(n8095), .Z(out[584]) );
  ANDN U5164 ( .B(n8098), .A(n8097), .Z(n8099) );
  XNOR U5165 ( .A(n8100), .B(n8099), .Z(out[585]) );
  ANDN U5166 ( .B(n8102), .A(n8101), .Z(n8103) );
  XNOR U5167 ( .A(n8104), .B(n8103), .Z(out[586]) );
  ANDN U5168 ( .B(n8106), .A(n8105), .Z(n8107) );
  XNOR U5169 ( .A(n8108), .B(n8107), .Z(out[587]) );
  ANDN U5170 ( .B(n8110), .A(n8109), .Z(n8111) );
  XNOR U5171 ( .A(n8112), .B(n8111), .Z(out[588]) );
  ANDN U5172 ( .B(n8114), .A(n8113), .Z(n8115) );
  XNOR U5173 ( .A(n8116), .B(n8115), .Z(out[589]) );
  ANDN U5174 ( .B(n8118), .A(n8117), .Z(n8119) );
  XNOR U5175 ( .A(n8120), .B(n8119), .Z(out[58]) );
  ANDN U5176 ( .B(n8122), .A(n8121), .Z(n8123) );
  XNOR U5177 ( .A(n8124), .B(n8123), .Z(out[590]) );
  ANDN U5178 ( .B(n8126), .A(n8125), .Z(n8127) );
  XNOR U5179 ( .A(n8128), .B(n8127), .Z(out[591]) );
  ANDN U5180 ( .B(n8130), .A(n8129), .Z(n8131) );
  XNOR U5181 ( .A(n8132), .B(n8131), .Z(out[592]) );
  ANDN U5182 ( .B(n8134), .A(n8133), .Z(n8135) );
  XNOR U5183 ( .A(n8136), .B(n8135), .Z(out[593]) );
  ANDN U5184 ( .B(n8138), .A(n8137), .Z(n8139) );
  XNOR U5185 ( .A(n8140), .B(n8139), .Z(out[594]) );
  ANDN U5186 ( .B(n8142), .A(n8141), .Z(n8143) );
  XNOR U5187 ( .A(n8144), .B(n8143), .Z(out[595]) );
  ANDN U5188 ( .B(n8146), .A(n8145), .Z(n8147) );
  XNOR U5189 ( .A(n8148), .B(n8147), .Z(out[596]) );
  ANDN U5190 ( .B(n8150), .A(n8149), .Z(n8151) );
  XNOR U5191 ( .A(n8152), .B(n8151), .Z(out[597]) );
  ANDN U5192 ( .B(n8154), .A(n8153), .Z(n8155) );
  XNOR U5193 ( .A(n8156), .B(n8155), .Z(out[598]) );
  ANDN U5194 ( .B(n8158), .A(n8157), .Z(n8159) );
  XNOR U5195 ( .A(n8160), .B(n8159), .Z(out[599]) );
  ANDN U5196 ( .B(n8162), .A(n8161), .Z(n8163) );
  XNOR U5197 ( .A(n8164), .B(n8163), .Z(out[59]) );
  OR U5198 ( .A(n8604), .B(n8165), .Z(n8166) );
  XNOR U5199 ( .A(n8603), .B(n8166), .Z(out[5]) );
  ANDN U5200 ( .B(n8168), .A(n8167), .Z(n8169) );
  XNOR U5201 ( .A(n8170), .B(n8169), .Z(out[600]) );
  ANDN U5202 ( .B(n8172), .A(n8171), .Z(n8173) );
  XNOR U5203 ( .A(n8174), .B(n8173), .Z(out[601]) );
  ANDN U5204 ( .B(n8176), .A(n8175), .Z(n8177) );
  XNOR U5205 ( .A(n8178), .B(n8177), .Z(out[602]) );
  ANDN U5206 ( .B(n8180), .A(n8179), .Z(n8181) );
  XNOR U5207 ( .A(n8182), .B(n8181), .Z(out[603]) );
  ANDN U5208 ( .B(n8184), .A(n8183), .Z(n8185) );
  XNOR U5209 ( .A(n8186), .B(n8185), .Z(out[604]) );
  ANDN U5210 ( .B(n8188), .A(n8187), .Z(n8189) );
  XNOR U5211 ( .A(n8190), .B(n8189), .Z(out[605]) );
  ANDN U5212 ( .B(n8192), .A(n8191), .Z(n8193) );
  XNOR U5213 ( .A(n8194), .B(n8193), .Z(out[606]) );
  ANDN U5214 ( .B(n8196), .A(n8195), .Z(n8197) );
  XNOR U5215 ( .A(n8198), .B(n8197), .Z(out[607]) );
  ANDN U5216 ( .B(n8200), .A(n8199), .Z(n8201) );
  XNOR U5217 ( .A(n8202), .B(n8201), .Z(out[608]) );
  ANDN U5218 ( .B(n8204), .A(n8203), .Z(n8205) );
  XNOR U5219 ( .A(n8206), .B(n8205), .Z(out[609]) );
  ANDN U5220 ( .B(n8208), .A(n8207), .Z(n8209) );
  XNOR U5221 ( .A(n8210), .B(n8209), .Z(out[60]) );
  ANDN U5222 ( .B(n8212), .A(n8211), .Z(n8213) );
  XNOR U5223 ( .A(n8214), .B(n8213), .Z(out[610]) );
  ANDN U5224 ( .B(n8216), .A(n8215), .Z(n8217) );
  XNOR U5225 ( .A(n8218), .B(n8217), .Z(out[611]) );
  ANDN U5226 ( .B(n8220), .A(n8219), .Z(n8221) );
  XNOR U5227 ( .A(n8222), .B(n8221), .Z(out[612]) );
  ANDN U5228 ( .B(n8224), .A(n8223), .Z(n8225) );
  XNOR U5229 ( .A(n8226), .B(n8225), .Z(out[613]) );
  ANDN U5230 ( .B(n8228), .A(n8227), .Z(n8229) );
  XNOR U5231 ( .A(n8230), .B(n8229), .Z(out[614]) );
  ANDN U5232 ( .B(n8232), .A(n8231), .Z(n8233) );
  XNOR U5233 ( .A(n8234), .B(n8233), .Z(out[615]) );
  ANDN U5234 ( .B(n8236), .A(n8235), .Z(n8237) );
  XNOR U5235 ( .A(n8238), .B(n8237), .Z(out[616]) );
  ANDN U5236 ( .B(n8240), .A(n8239), .Z(n8241) );
  XNOR U5237 ( .A(n8242), .B(n8241), .Z(out[617]) );
  ANDN U5238 ( .B(n8244), .A(n8243), .Z(n8245) );
  XNOR U5239 ( .A(n8246), .B(n8245), .Z(out[618]) );
  ANDN U5240 ( .B(n8248), .A(n8247), .Z(n8249) );
  XNOR U5241 ( .A(n8250), .B(n8249), .Z(out[619]) );
  ANDN U5242 ( .B(n8252), .A(n8251), .Z(n8253) );
  XNOR U5243 ( .A(n8254), .B(n8253), .Z(out[61]) );
  ANDN U5244 ( .B(n8256), .A(n8255), .Z(n8257) );
  XNOR U5245 ( .A(n8258), .B(n8257), .Z(out[620]) );
  ANDN U5246 ( .B(n8260), .A(n8259), .Z(n8261) );
  XNOR U5247 ( .A(n8262), .B(n8261), .Z(out[621]) );
  ANDN U5248 ( .B(n8264), .A(n8263), .Z(n8265) );
  XNOR U5249 ( .A(n8266), .B(n8265), .Z(out[622]) );
  ANDN U5250 ( .B(n8268), .A(n8267), .Z(n8269) );
  XNOR U5251 ( .A(n8270), .B(n8269), .Z(out[623]) );
  ANDN U5252 ( .B(n8272), .A(n8271), .Z(n8273) );
  XNOR U5253 ( .A(n8274), .B(n8273), .Z(out[624]) );
  ANDN U5254 ( .B(n8276), .A(n8275), .Z(n8277) );
  XNOR U5255 ( .A(n8278), .B(n8277), .Z(out[625]) );
  ANDN U5256 ( .B(n8280), .A(n8279), .Z(n8281) );
  XNOR U5257 ( .A(n8282), .B(n8281), .Z(out[626]) );
  ANDN U5258 ( .B(n8284), .A(n8283), .Z(n8285) );
  XNOR U5259 ( .A(n8286), .B(n8285), .Z(out[627]) );
  ANDN U5260 ( .B(n8288), .A(n8287), .Z(n8289) );
  XNOR U5261 ( .A(n8290), .B(n8289), .Z(out[628]) );
  ANDN U5262 ( .B(n8292), .A(n8291), .Z(n8293) );
  XNOR U5263 ( .A(n8294), .B(n8293), .Z(out[629]) );
  ANDN U5264 ( .B(n8296), .A(n8295), .Z(n8297) );
  XNOR U5265 ( .A(n8298), .B(n8297), .Z(out[62]) );
  ANDN U5266 ( .B(n8300), .A(n8299), .Z(n8301) );
  XNOR U5267 ( .A(n8302), .B(n8301), .Z(out[630]) );
  ANDN U5268 ( .B(n8304), .A(n8303), .Z(n8305) );
  XNOR U5269 ( .A(n8306), .B(n8305), .Z(out[631]) );
  ANDN U5270 ( .B(n8308), .A(n8307), .Z(n8309) );
  XNOR U5271 ( .A(n8310), .B(n8309), .Z(out[632]) );
  ANDN U5272 ( .B(n8312), .A(n8311), .Z(n8313) );
  XNOR U5273 ( .A(n8314), .B(n8313), .Z(out[633]) );
  ANDN U5274 ( .B(n8316), .A(n8315), .Z(n8317) );
  XNOR U5275 ( .A(n8318), .B(n8317), .Z(out[634]) );
  ANDN U5276 ( .B(n8320), .A(n8319), .Z(n8321) );
  XNOR U5277 ( .A(n8322), .B(n8321), .Z(out[635]) );
  ANDN U5278 ( .B(n8324), .A(n8323), .Z(n8325) );
  XNOR U5279 ( .A(n8326), .B(n8325), .Z(out[636]) );
  ANDN U5280 ( .B(n8328), .A(n8327), .Z(n8329) );
  XNOR U5281 ( .A(n8330), .B(n8329), .Z(out[637]) );
  ANDN U5282 ( .B(n8332), .A(n8331), .Z(n8333) );
  XNOR U5283 ( .A(n8334), .B(n8333), .Z(out[638]) );
  ANDN U5284 ( .B(n8336), .A(n8335), .Z(n8337) );
  XNOR U5285 ( .A(n8338), .B(n8337), .Z(out[639]) );
  ANDN U5286 ( .B(n8340), .A(n8339), .Z(n8341) );
  XNOR U5287 ( .A(n8342), .B(n8341), .Z(out[63]) );
  XNOR U5288 ( .A(in[302]), .B(n8343), .Z(n8772) );
  XNOR U5289 ( .A(in[1535]), .B(n8344), .Z(n9150) );
  XNOR U5290 ( .A(in[1146]), .B(n8345), .Z(n9147) );
  NAND U5291 ( .A(n9150), .B(n9147), .Z(n8346) );
  XNOR U5292 ( .A(n8772), .B(n8346), .Z(out[640]) );
  XNOR U5293 ( .A(in[303]), .B(n8347), .Z(n8775) );
  XNOR U5294 ( .A(in[1472]), .B(n8348), .Z(n9154) );
  XNOR U5295 ( .A(in[1147]), .B(n8349), .Z(n9151) );
  NAND U5296 ( .A(n9154), .B(n9151), .Z(n8350) );
  XNOR U5297 ( .A(n8775), .B(n8350), .Z(out[641]) );
  XNOR U5298 ( .A(in[304]), .B(n8351), .Z(n8782) );
  XNOR U5299 ( .A(in[1473]), .B(n8352), .Z(n9158) );
  XNOR U5300 ( .A(in[1148]), .B(n8353), .Z(n9155) );
  NAND U5301 ( .A(n9158), .B(n9155), .Z(n8354) );
  XNOR U5302 ( .A(n8782), .B(n8354), .Z(out[642]) );
  XNOR U5303 ( .A(in[305]), .B(n8355), .Z(n8785) );
  XNOR U5304 ( .A(in[1474]), .B(n8356), .Z(n9162) );
  XNOR U5305 ( .A(in[1149]), .B(n8357), .Z(n9159) );
  NAND U5306 ( .A(n9162), .B(n9159), .Z(n8358) );
  XNOR U5307 ( .A(n8785), .B(n8358), .Z(out[643]) );
  XNOR U5308 ( .A(in[306]), .B(n8359), .Z(n8788) );
  XNOR U5309 ( .A(in[1475]), .B(n8360), .Z(n9174) );
  XNOR U5310 ( .A(in[1150]), .B(n8361), .Z(n9171) );
  NAND U5311 ( .A(n9174), .B(n9171), .Z(n8362) );
  XNOR U5312 ( .A(n8788), .B(n8362), .Z(out[644]) );
  XNOR U5313 ( .A(in[307]), .B(n8363), .Z(n8791) );
  XNOR U5314 ( .A(in[1476]), .B(n8364), .Z(n9178) );
  XNOR U5315 ( .A(in[1151]), .B(n8365), .Z(n9175) );
  NAND U5316 ( .A(n9178), .B(n9175), .Z(n8366) );
  XNOR U5317 ( .A(n8791), .B(n8366), .Z(out[645]) );
  XNOR U5318 ( .A(in[308]), .B(n8367), .Z(n8794) );
  XNOR U5319 ( .A(in[1477]), .B(n8368), .Z(n9182) );
  XNOR U5320 ( .A(in[1088]), .B(n8369), .Z(n9179) );
  NAND U5321 ( .A(n9182), .B(n9179), .Z(n8370) );
  XNOR U5322 ( .A(n8794), .B(n8370), .Z(out[646]) );
  XNOR U5323 ( .A(in[309]), .B(n8371), .Z(n8797) );
  XNOR U5324 ( .A(in[1478]), .B(n8372), .Z(n9186) );
  XNOR U5325 ( .A(in[1089]), .B(n8373), .Z(n9183) );
  NAND U5326 ( .A(n9186), .B(n9183), .Z(n8374) );
  XNOR U5327 ( .A(n8797), .B(n8374), .Z(out[647]) );
  XNOR U5328 ( .A(in[310]), .B(n8375), .Z(n8800) );
  XNOR U5329 ( .A(in[1479]), .B(n8376), .Z(n9190) );
  XOR U5330 ( .A(n8377), .B(in[1090]), .Z(n9187) );
  NAND U5331 ( .A(n9190), .B(n9187), .Z(n8378) );
  XNOR U5332 ( .A(n8800), .B(n8378), .Z(out[648]) );
  XNOR U5333 ( .A(in[311]), .B(n8379), .Z(n8803) );
  XNOR U5334 ( .A(in[1480]), .B(n8380), .Z(n9194) );
  XOR U5335 ( .A(n8381), .B(in[1091]), .Z(n9191) );
  NAND U5336 ( .A(n9194), .B(n9191), .Z(n8382) );
  XNOR U5337 ( .A(n8803), .B(n8382), .Z(out[649]) );
  NOR U5338 ( .A(n8384), .B(n8383), .Z(n8385) );
  XNOR U5339 ( .A(n8386), .B(n8385), .Z(out[64]) );
  XNOR U5340 ( .A(in[312]), .B(n8387), .Z(n8806) );
  XNOR U5341 ( .A(in[1481]), .B(n8388), .Z(n9198) );
  XOR U5342 ( .A(n8389), .B(in[1092]), .Z(n9195) );
  NAND U5343 ( .A(n9198), .B(n9195), .Z(n8390) );
  XNOR U5344 ( .A(n8806), .B(n8390), .Z(out[650]) );
  XNOR U5345 ( .A(in[313]), .B(n8391), .Z(n8809) );
  XNOR U5346 ( .A(in[1482]), .B(n8392), .Z(n9202) );
  XOR U5347 ( .A(n8393), .B(in[1093]), .Z(n9199) );
  NAND U5348 ( .A(n9202), .B(n9199), .Z(n8394) );
  XNOR U5349 ( .A(n8809), .B(n8394), .Z(out[651]) );
  XNOR U5350 ( .A(in[314]), .B(n8395), .Z(n8816) );
  XNOR U5351 ( .A(in[1483]), .B(n8396), .Z(n9206) );
  XOR U5352 ( .A(n8397), .B(in[1094]), .Z(n9203) );
  NAND U5353 ( .A(n9206), .B(n9203), .Z(n8398) );
  XNOR U5354 ( .A(n8816), .B(n8398), .Z(out[652]) );
  XNOR U5355 ( .A(in[315]), .B(n8399), .Z(n8819) );
  XNOR U5356 ( .A(in[1484]), .B(n8400), .Z(n9210) );
  XOR U5357 ( .A(n8401), .B(in[1095]), .Z(n9207) );
  NAND U5358 ( .A(n9210), .B(n9207), .Z(n8402) );
  XNOR U5359 ( .A(n8819), .B(n8402), .Z(out[653]) );
  XNOR U5360 ( .A(in[316]), .B(n8403), .Z(n8822) );
  XNOR U5361 ( .A(in[1485]), .B(n8404), .Z(n9218) );
  XOR U5362 ( .A(n8405), .B(in[1096]), .Z(n9215) );
  NAND U5363 ( .A(n9218), .B(n9215), .Z(n8406) );
  XNOR U5364 ( .A(n8822), .B(n8406), .Z(out[654]) );
  XNOR U5365 ( .A(in[317]), .B(n8407), .Z(n8825) );
  XNOR U5366 ( .A(in[1486]), .B(n8408), .Z(n9222) );
  XOR U5367 ( .A(in[1097]), .B(n8409), .Z(n9219) );
  NAND U5368 ( .A(n9222), .B(n9219), .Z(n8410) );
  XNOR U5369 ( .A(n8825), .B(n8410), .Z(out[655]) );
  XNOR U5370 ( .A(in[318]), .B(n8411), .Z(n8828) );
  XNOR U5371 ( .A(in[1487]), .B(n8412), .Z(n9226) );
  XOR U5372 ( .A(n8413), .B(in[1098]), .Z(n9223) );
  NAND U5373 ( .A(n9226), .B(n9223), .Z(n8414) );
  XNOR U5374 ( .A(n8828), .B(n8414), .Z(out[656]) );
  XNOR U5375 ( .A(in[319]), .B(n8415), .Z(n8831) );
  XNOR U5376 ( .A(in[1488]), .B(n8416), .Z(n9230) );
  XOR U5377 ( .A(n8417), .B(in[1099]), .Z(n9227) );
  NAND U5378 ( .A(n9230), .B(n9227), .Z(n8418) );
  XNOR U5379 ( .A(n8831), .B(n8418), .Z(out[657]) );
  XNOR U5380 ( .A(in[256]), .B(n8419), .Z(n8834) );
  XNOR U5381 ( .A(in[1489]), .B(n8420), .Z(n9234) );
  XOR U5382 ( .A(in[1100]), .B(n8421), .Z(n9231) );
  NAND U5383 ( .A(n9234), .B(n9231), .Z(n8422) );
  XNOR U5384 ( .A(n8834), .B(n8422), .Z(out[658]) );
  XNOR U5385 ( .A(in[257]), .B(n8423), .Z(n8837) );
  XNOR U5386 ( .A(in[1490]), .B(n8424), .Z(n9238) );
  XOR U5387 ( .A(in[1101]), .B(n8425), .Z(n9235) );
  NAND U5388 ( .A(n9238), .B(n9235), .Z(n8426) );
  XNOR U5389 ( .A(n8837), .B(n8426), .Z(out[659]) );
  NOR U5390 ( .A(n8428), .B(n8427), .Z(n8429) );
  XNOR U5391 ( .A(n8430), .B(n8429), .Z(out[65]) );
  XNOR U5392 ( .A(in[258]), .B(n8431), .Z(n8840) );
  XOR U5393 ( .A(in[1491]), .B(n8432), .Z(n9242) );
  XOR U5394 ( .A(in[1102]), .B(n8433), .Z(n9239) );
  NAND U5395 ( .A(n9242), .B(n9239), .Z(n8434) );
  XNOR U5396 ( .A(n8840), .B(n8434), .Z(out[660]) );
  XNOR U5397 ( .A(in[259]), .B(n8435), .Z(n8843) );
  XOR U5398 ( .A(in[1492]), .B(n8436), .Z(n9246) );
  XOR U5399 ( .A(in[1103]), .B(n8437), .Z(n9243) );
  NAND U5400 ( .A(n9246), .B(n9243), .Z(n8438) );
  XNOR U5401 ( .A(n8843), .B(n8438), .Z(out[661]) );
  XOR U5402 ( .A(in[260]), .B(n8439), .Z(n8850) );
  XOR U5403 ( .A(in[1493]), .B(n8440), .Z(n9250) );
  XOR U5404 ( .A(in[1104]), .B(n8441), .Z(n9247) );
  NAND U5405 ( .A(n9250), .B(n9247), .Z(n8442) );
  XNOR U5406 ( .A(n8850), .B(n8442), .Z(out[662]) );
  XOR U5407 ( .A(in[261]), .B(n8443), .Z(n8853) );
  XOR U5408 ( .A(in[1494]), .B(n8444), .Z(n9254) );
  XOR U5409 ( .A(in[1105]), .B(n8445), .Z(n9251) );
  NAND U5410 ( .A(n9254), .B(n9251), .Z(n8446) );
  XNOR U5411 ( .A(n8853), .B(n8446), .Z(out[663]) );
  XOR U5412 ( .A(in[262]), .B(n8447), .Z(n8856) );
  XOR U5413 ( .A(in[1495]), .B(n8448), .Z(n9262) );
  XOR U5414 ( .A(in[1106]), .B(n8449), .Z(n9259) );
  NAND U5415 ( .A(n9262), .B(n9259), .Z(n8450) );
  XNOR U5416 ( .A(n8856), .B(n8450), .Z(out[664]) );
  XOR U5417 ( .A(in[263]), .B(n8451), .Z(n8859) );
  XOR U5418 ( .A(in[1496]), .B(n8452), .Z(n9266) );
  XOR U5419 ( .A(in[1107]), .B(n8453), .Z(n9263) );
  NAND U5420 ( .A(n9266), .B(n9263), .Z(n8454) );
  XNOR U5421 ( .A(n8859), .B(n8454), .Z(out[665]) );
  XOR U5422 ( .A(in[264]), .B(n8455), .Z(n8862) );
  XOR U5423 ( .A(in[1497]), .B(n8456), .Z(n9270) );
  XOR U5424 ( .A(in[1108]), .B(n8457), .Z(n9267) );
  NAND U5425 ( .A(n9270), .B(n9267), .Z(n8458) );
  XNOR U5426 ( .A(n8862), .B(n8458), .Z(out[666]) );
  XOR U5427 ( .A(in[265]), .B(n8459), .Z(n8865) );
  XOR U5428 ( .A(in[1498]), .B(n8460), .Z(n9274) );
  XOR U5429 ( .A(in[1109]), .B(n8461), .Z(n9271) );
  NAND U5430 ( .A(n9274), .B(n9271), .Z(n8462) );
  XNOR U5431 ( .A(n8865), .B(n8462), .Z(out[667]) );
  XOR U5432 ( .A(in[266]), .B(n8463), .Z(n8868) );
  XOR U5433 ( .A(in[1499]), .B(n8464), .Z(n9278) );
  XOR U5434 ( .A(in[1110]), .B(n8465), .Z(n9275) );
  NAND U5435 ( .A(n9278), .B(n9275), .Z(n8466) );
  XNOR U5436 ( .A(n8868), .B(n8466), .Z(out[668]) );
  XOR U5437 ( .A(in[267]), .B(n8467), .Z(n8871) );
  XOR U5438 ( .A(in[1500]), .B(n8468), .Z(n9282) );
  XOR U5439 ( .A(in[1111]), .B(n8469), .Z(n9279) );
  NAND U5440 ( .A(n9282), .B(n9279), .Z(n8470) );
  XNOR U5441 ( .A(n8871), .B(n8470), .Z(out[669]) );
  ANDN U5442 ( .B(n8472), .A(n8471), .Z(n8473) );
  XNOR U5443 ( .A(n8474), .B(n8473), .Z(out[66]) );
  XOR U5444 ( .A(in[268]), .B(n8475), .Z(n8874) );
  XOR U5445 ( .A(in[1501]), .B(n8476), .Z(n9286) );
  XOR U5446 ( .A(in[1112]), .B(n8477), .Z(n9283) );
  NAND U5447 ( .A(n9286), .B(n9283), .Z(n8478) );
  XNOR U5448 ( .A(n8874), .B(n8478), .Z(out[670]) );
  XOR U5449 ( .A(in[269]), .B(n8479), .Z(n8877) );
  XOR U5450 ( .A(in[1502]), .B(n8480), .Z(n9290) );
  XOR U5451 ( .A(in[1113]), .B(n8481), .Z(n9287) );
  NAND U5452 ( .A(n9290), .B(n9287), .Z(n8482) );
  XNOR U5453 ( .A(n8877), .B(n8482), .Z(out[671]) );
  XOR U5454 ( .A(in[270]), .B(n8483), .Z(n8888) );
  XOR U5455 ( .A(in[1503]), .B(n8484), .Z(n9294) );
  XOR U5456 ( .A(in[1114]), .B(n8485), .Z(n9291) );
  NAND U5457 ( .A(n9294), .B(n9291), .Z(n8486) );
  XNOR U5458 ( .A(n8888), .B(n8486), .Z(out[672]) );
  XOR U5459 ( .A(in[271]), .B(n8487), .Z(n8891) );
  XOR U5460 ( .A(in[1504]), .B(n8488), .Z(n9298) );
  XOR U5461 ( .A(in[1115]), .B(n8489), .Z(n9295) );
  NAND U5462 ( .A(n9298), .B(n9295), .Z(n8490) );
  XNOR U5463 ( .A(n8891), .B(n8490), .Z(out[673]) );
  XOR U5464 ( .A(in[272]), .B(n8491), .Z(n8894) );
  XOR U5465 ( .A(in[1505]), .B(n8492), .Z(n9306) );
  XOR U5466 ( .A(in[1116]), .B(n8493), .Z(n9303) );
  NAND U5467 ( .A(n9306), .B(n9303), .Z(n8494) );
  XNOR U5468 ( .A(n8894), .B(n8494), .Z(out[674]) );
  XOR U5469 ( .A(in[273]), .B(n8495), .Z(n8897) );
  XNOR U5470 ( .A(n8496), .B(in[1506]), .Z(n9310) );
  XOR U5471 ( .A(in[1117]), .B(n8497), .Z(n9307) );
  NAND U5472 ( .A(n9310), .B(n9307), .Z(n8498) );
  XNOR U5473 ( .A(n8897), .B(n8498), .Z(out[675]) );
  XOR U5474 ( .A(in[274]), .B(n8499), .Z(n8900) );
  XNOR U5475 ( .A(n8500), .B(in[1507]), .Z(n9314) );
  XOR U5476 ( .A(in[1118]), .B(n8501), .Z(n9311) );
  NAND U5477 ( .A(n9314), .B(n9311), .Z(n8502) );
  XNOR U5478 ( .A(n8900), .B(n8502), .Z(out[676]) );
  XOR U5479 ( .A(in[275]), .B(n8503), .Z(n8903) );
  XNOR U5480 ( .A(n8504), .B(in[1508]), .Z(n9318) );
  XOR U5481 ( .A(in[1119]), .B(n8505), .Z(n9315) );
  NAND U5482 ( .A(n9318), .B(n9315), .Z(n8506) );
  XNOR U5483 ( .A(n8903), .B(n8506), .Z(out[677]) );
  XOR U5484 ( .A(in[276]), .B(n8507), .Z(n8906) );
  XNOR U5485 ( .A(n8508), .B(in[1509]), .Z(n9322) );
  XOR U5486 ( .A(in[1120]), .B(n8509), .Z(n9319) );
  NAND U5487 ( .A(n9322), .B(n9319), .Z(n8510) );
  XNOR U5488 ( .A(n8906), .B(n8510), .Z(out[678]) );
  XOR U5489 ( .A(in[277]), .B(n8511), .Z(n8909) );
  XOR U5490 ( .A(in[1510]), .B(n8512), .Z(n9326) );
  XOR U5491 ( .A(in[1121]), .B(n8513), .Z(n9323) );
  NAND U5492 ( .A(n9326), .B(n9323), .Z(n8514) );
  XNOR U5493 ( .A(n8909), .B(n8514), .Z(out[679]) );
  ANDN U5494 ( .B(n8516), .A(n8515), .Z(n8517) );
  XNOR U5495 ( .A(n8518), .B(n8517), .Z(out[67]) );
  XOR U5496 ( .A(in[278]), .B(n8519), .Z(n8912) );
  XOR U5497 ( .A(in[1511]), .B(n8520), .Z(n9330) );
  XOR U5498 ( .A(in[1122]), .B(n8521), .Z(n9327) );
  NAND U5499 ( .A(n9330), .B(n9327), .Z(n8522) );
  XNOR U5500 ( .A(n8912), .B(n8522), .Z(out[680]) );
  XOR U5501 ( .A(in[279]), .B(n8523), .Z(n8915) );
  XOR U5502 ( .A(in[1512]), .B(n8524), .Z(n9334) );
  XOR U5503 ( .A(in[1123]), .B(n8525), .Z(n9331) );
  NAND U5504 ( .A(n9334), .B(n9331), .Z(n8526) );
  XNOR U5505 ( .A(n8915), .B(n8526), .Z(out[681]) );
  XOR U5506 ( .A(in[280]), .B(n8527), .Z(n8922) );
  XOR U5507 ( .A(in[1513]), .B(n8528), .Z(n9338) );
  XOR U5508 ( .A(in[1124]), .B(n8529), .Z(n9335) );
  NAND U5509 ( .A(n9338), .B(n9335), .Z(n8530) );
  XNOR U5510 ( .A(n8922), .B(n8530), .Z(out[682]) );
  XOR U5511 ( .A(in[281]), .B(n8531), .Z(n8925) );
  XOR U5512 ( .A(in[1514]), .B(n8532), .Z(n9342) );
  XOR U5513 ( .A(in[1125]), .B(n8533), .Z(n9339) );
  NAND U5514 ( .A(n9342), .B(n9339), .Z(n8534) );
  XNOR U5515 ( .A(n8925), .B(n8534), .Z(out[683]) );
  XOR U5516 ( .A(in[282]), .B(n8535), .Z(n8928) );
  XOR U5517 ( .A(in[1515]), .B(n8536), .Z(n9350) );
  XNOR U5518 ( .A(in[1126]), .B(n8537), .Z(n9347) );
  NAND U5519 ( .A(n9350), .B(n9347), .Z(n8538) );
  XNOR U5520 ( .A(n8928), .B(n8538), .Z(out[684]) );
  XOR U5521 ( .A(in[283]), .B(n8539), .Z(n8931) );
  XOR U5522 ( .A(in[1516]), .B(n8540), .Z(n9354) );
  XNOR U5523 ( .A(in[1127]), .B(n8541), .Z(n9351) );
  NAND U5524 ( .A(n9354), .B(n9351), .Z(n8542) );
  XNOR U5525 ( .A(n8931), .B(n8542), .Z(out[685]) );
  XOR U5526 ( .A(in[284]), .B(n8543), .Z(n8934) );
  XOR U5527 ( .A(in[1517]), .B(n8544), .Z(n9358) );
  XNOR U5528 ( .A(in[1128]), .B(n8545), .Z(n9355) );
  NAND U5529 ( .A(n9358), .B(n9355), .Z(n8546) );
  XNOR U5530 ( .A(n8934), .B(n8546), .Z(out[686]) );
  XOR U5531 ( .A(in[285]), .B(n8547), .Z(n8937) );
  XOR U5532 ( .A(in[1518]), .B(n8548), .Z(n9362) );
  XNOR U5533 ( .A(in[1129]), .B(n8549), .Z(n9359) );
  NAND U5534 ( .A(n9362), .B(n9359), .Z(n8550) );
  XNOR U5535 ( .A(n8937), .B(n8550), .Z(out[687]) );
  XOR U5536 ( .A(in[286]), .B(n8551), .Z(n8940) );
  XOR U5537 ( .A(in[1519]), .B(n8552), .Z(n9366) );
  XNOR U5538 ( .A(in[1130]), .B(n8553), .Z(n9363) );
  NAND U5539 ( .A(n9366), .B(n9363), .Z(n8554) );
  XNOR U5540 ( .A(n8940), .B(n8554), .Z(out[688]) );
  XOR U5541 ( .A(in[287]), .B(n8555), .Z(n8943) );
  XOR U5542 ( .A(in[1520]), .B(n8556), .Z(n9370) );
  XNOR U5543 ( .A(in[1131]), .B(n8557), .Z(n9367) );
  NAND U5544 ( .A(n9370), .B(n9367), .Z(n8558) );
  XNOR U5545 ( .A(n8943), .B(n8558), .Z(out[689]) );
  ANDN U5546 ( .B(n8560), .A(n8559), .Z(n8561) );
  XNOR U5547 ( .A(n8562), .B(n8561), .Z(out[68]) );
  XOR U5548 ( .A(in[288]), .B(n8563), .Z(n8946) );
  XOR U5549 ( .A(in[1521]), .B(n8564), .Z(n9374) );
  XNOR U5550 ( .A(in[1132]), .B(n8565), .Z(n9371) );
  NAND U5551 ( .A(n9374), .B(n9371), .Z(n8566) );
  XNOR U5552 ( .A(n8946), .B(n8566), .Z(out[690]) );
  XOR U5553 ( .A(in[289]), .B(n8567), .Z(n8949) );
  XOR U5554 ( .A(in[1522]), .B(n8568), .Z(n9378) );
  XNOR U5555 ( .A(in[1133]), .B(n8569), .Z(n9375) );
  NAND U5556 ( .A(n9378), .B(n9375), .Z(n8570) );
  XNOR U5557 ( .A(n8949), .B(n8570), .Z(out[691]) );
  XOR U5558 ( .A(in[290]), .B(n8571), .Z(n8956) );
  XOR U5559 ( .A(in[1523]), .B(n8572), .Z(n9382) );
  XNOR U5560 ( .A(in[1134]), .B(n8573), .Z(n9379) );
  NAND U5561 ( .A(n9382), .B(n9379), .Z(n8574) );
  XNOR U5562 ( .A(n8956), .B(n8574), .Z(out[692]) );
  XOR U5563 ( .A(in[291]), .B(n8575), .Z(n8959) );
  XOR U5564 ( .A(in[1524]), .B(n8576), .Z(n9386) );
  XNOR U5565 ( .A(in[1135]), .B(n8577), .Z(n9383) );
  NAND U5566 ( .A(n9386), .B(n9383), .Z(n8578) );
  XNOR U5567 ( .A(n8959), .B(n8578), .Z(out[693]) );
  XOR U5568 ( .A(in[292]), .B(n8579), .Z(n8962) );
  XOR U5569 ( .A(in[1525]), .B(n8580), .Z(n9394) );
  XNOR U5570 ( .A(in[1136]), .B(n8581), .Z(n9391) );
  NAND U5571 ( .A(n9394), .B(n9391), .Z(n8582) );
  XNOR U5572 ( .A(n8962), .B(n8582), .Z(out[694]) );
  XNOR U5573 ( .A(in[293]), .B(n8583), .Z(n8965) );
  XOR U5574 ( .A(in[1526]), .B(n8584), .Z(n9398) );
  XNOR U5575 ( .A(in[1137]), .B(n8585), .Z(n9395) );
  NAND U5576 ( .A(n9398), .B(n9395), .Z(n8586) );
  XNOR U5577 ( .A(n8965), .B(n8586), .Z(out[695]) );
  XNOR U5578 ( .A(in[294]), .B(n8587), .Z(n8968) );
  XOR U5579 ( .A(in[1527]), .B(n8588), .Z(n9402) );
  XNOR U5580 ( .A(in[1138]), .B(n8589), .Z(n9399) );
  NAND U5581 ( .A(n9402), .B(n9399), .Z(n8590) );
  XNOR U5582 ( .A(n8968), .B(n8590), .Z(out[696]) );
  XNOR U5583 ( .A(in[295]), .B(n8591), .Z(n8971) );
  XOR U5584 ( .A(in[1528]), .B(n8592), .Z(n9406) );
  XNOR U5585 ( .A(in[1139]), .B(n8593), .Z(n9403) );
  NAND U5586 ( .A(n9406), .B(n9403), .Z(n8594) );
  XNOR U5587 ( .A(n8971), .B(n8594), .Z(out[697]) );
  XNOR U5588 ( .A(in[296]), .B(n8595), .Z(n8974) );
  XOR U5589 ( .A(in[1529]), .B(n8596), .Z(n9410) );
  XNOR U5590 ( .A(in[1140]), .B(n8597), .Z(n9407) );
  NAND U5591 ( .A(n9410), .B(n9407), .Z(n8598) );
  XNOR U5592 ( .A(n8974), .B(n8598), .Z(out[698]) );
  XNOR U5593 ( .A(in[297]), .B(n8599), .Z(n8977) );
  XOR U5594 ( .A(in[1530]), .B(n8600), .Z(n9414) );
  XNOR U5595 ( .A(in[1141]), .B(n8601), .Z(n9411) );
  NAND U5596 ( .A(n9414), .B(n9411), .Z(n8602) );
  XNOR U5597 ( .A(n8977), .B(n8602), .Z(out[699]) );
  ANDN U5598 ( .B(n8604), .A(n8603), .Z(n8605) );
  XNOR U5599 ( .A(n8606), .B(n8605), .Z(out[69]) );
  OR U5600 ( .A(n8638), .B(n8607), .Z(n8608) );
  XNOR U5601 ( .A(n8637), .B(n8608), .Z(out[6]) );
  XNOR U5602 ( .A(in[298]), .B(n8609), .Z(n8980) );
  XNOR U5603 ( .A(in[1531]), .B(n8610), .Z(n9418) );
  XNOR U5604 ( .A(in[1142]), .B(n8611), .Z(n9415) );
  NAND U5605 ( .A(n9418), .B(n9415), .Z(n8612) );
  XNOR U5606 ( .A(n8980), .B(n8612), .Z(out[700]) );
  XNOR U5607 ( .A(in[299]), .B(n8613), .Z(n8983) );
  XNOR U5608 ( .A(in[1532]), .B(n8614), .Z(n9422) );
  XNOR U5609 ( .A(in[1143]), .B(n8615), .Z(n9419) );
  NAND U5610 ( .A(n9422), .B(n9419), .Z(n8616) );
  XNOR U5611 ( .A(n8983), .B(n8616), .Z(out[701]) );
  XNOR U5612 ( .A(in[300]), .B(n8617), .Z(n8990) );
  XNOR U5613 ( .A(in[1533]), .B(n8618), .Z(n9426) );
  XNOR U5614 ( .A(in[1144]), .B(n8619), .Z(n9423) );
  NAND U5615 ( .A(n9426), .B(n9423), .Z(n8620) );
  XNOR U5616 ( .A(n8990), .B(n8620), .Z(out[702]) );
  XNOR U5617 ( .A(in[301]), .B(n8621), .Z(n8993) );
  XOR U5618 ( .A(in[1534]), .B(n8622), .Z(n9430) );
  XNOR U5619 ( .A(in[1145]), .B(n8623), .Z(n9427) );
  NAND U5620 ( .A(n9430), .B(n9427), .Z(n8624) );
  XNOR U5621 ( .A(n8993), .B(n8624), .Z(out[703]) );
  XOR U5622 ( .A(in[376]), .B(n8625), .Z(n8995) );
  NOR U5623 ( .A(n8772), .B(n9150), .Z(n8626) );
  XNOR U5624 ( .A(n8995), .B(n8626), .Z(out[704]) );
  XOR U5625 ( .A(in[377]), .B(n8627), .Z(n8997) );
  NOR U5626 ( .A(n8775), .B(n9154), .Z(n8628) );
  XNOR U5627 ( .A(n8997), .B(n8628), .Z(out[705]) );
  XOR U5628 ( .A(in[378]), .B(n8629), .Z(n8999) );
  NOR U5629 ( .A(n8782), .B(n9158), .Z(n8630) );
  XNOR U5630 ( .A(n8999), .B(n8630), .Z(out[706]) );
  XOR U5631 ( .A(in[379]), .B(n8631), .Z(n9001) );
  NOR U5632 ( .A(n8785), .B(n9162), .Z(n8632) );
  XNOR U5633 ( .A(n9001), .B(n8632), .Z(out[707]) );
  XOR U5634 ( .A(in[380]), .B(n8633), .Z(n9003) );
  NOR U5635 ( .A(n8788), .B(n9174), .Z(n8634) );
  XNOR U5636 ( .A(n9003), .B(n8634), .Z(out[708]) );
  XOR U5637 ( .A(in[381]), .B(n8635), .Z(n9005) );
  NOR U5638 ( .A(n8791), .B(n9178), .Z(n8636) );
  XNOR U5639 ( .A(n9005), .B(n8636), .Z(out[709]) );
  ANDN U5640 ( .B(n8638), .A(n8637), .Z(n8639) );
  XNOR U5641 ( .A(n8640), .B(n8639), .Z(out[70]) );
  XOR U5642 ( .A(in[382]), .B(n8641), .Z(n9007) );
  NOR U5643 ( .A(n8794), .B(n9182), .Z(n8642) );
  XNOR U5644 ( .A(n9007), .B(n8642), .Z(out[710]) );
  XOR U5645 ( .A(in[383]), .B(n8643), .Z(n9009) );
  NOR U5646 ( .A(n8797), .B(n9186), .Z(n8644) );
  XNOR U5647 ( .A(n9009), .B(n8644), .Z(out[711]) );
  XOR U5648 ( .A(in[320]), .B(n8645), .Z(n9015) );
  NOR U5649 ( .A(n8800), .B(n9190), .Z(n8646) );
  XNOR U5650 ( .A(n9015), .B(n8646), .Z(out[712]) );
  XOR U5651 ( .A(in[321]), .B(n8647), .Z(n9017) );
  NOR U5652 ( .A(n8803), .B(n9194), .Z(n8648) );
  XNOR U5653 ( .A(n9017), .B(n8648), .Z(out[713]) );
  XOR U5654 ( .A(in[322]), .B(n8649), .Z(n9019) );
  NOR U5655 ( .A(n8806), .B(n9198), .Z(n8650) );
  XNOR U5656 ( .A(n9019), .B(n8650), .Z(out[714]) );
  XOR U5657 ( .A(in[323]), .B(n8651), .Z(n9021) );
  NOR U5658 ( .A(n8809), .B(n9202), .Z(n8652) );
  XNOR U5659 ( .A(n9021), .B(n8652), .Z(out[715]) );
  XOR U5660 ( .A(in[324]), .B(n8653), .Z(n9023) );
  NOR U5661 ( .A(n8816), .B(n9206), .Z(n8654) );
  XNOR U5662 ( .A(n9023), .B(n8654), .Z(out[716]) );
  XOR U5663 ( .A(in[325]), .B(n8655), .Z(n9025) );
  NOR U5664 ( .A(n8819), .B(n9210), .Z(n8656) );
  XNOR U5665 ( .A(n9025), .B(n8656), .Z(out[717]) );
  XOR U5666 ( .A(in[326]), .B(n8657), .Z(n9027) );
  NOR U5667 ( .A(n8822), .B(n9218), .Z(n8658) );
  XNOR U5668 ( .A(n9027), .B(n8658), .Z(out[718]) );
  XOR U5669 ( .A(in[327]), .B(n8659), .Z(n9029) );
  NOR U5670 ( .A(n8825), .B(n9222), .Z(n8660) );
  XNOR U5671 ( .A(n9029), .B(n8660), .Z(out[719]) );
  ANDN U5672 ( .B(n8884), .A(n8886), .Z(n8661) );
  XNOR U5673 ( .A(n8662), .B(n8661), .Z(out[71]) );
  XOR U5674 ( .A(in[328]), .B(n8663), .Z(n9031) );
  NOR U5675 ( .A(n8828), .B(n9226), .Z(n8664) );
  XNOR U5676 ( .A(n9031), .B(n8664), .Z(out[720]) );
  XOR U5677 ( .A(in[329]), .B(n8665), .Z(n9033) );
  NOR U5678 ( .A(n8831), .B(n9230), .Z(n8666) );
  XNOR U5679 ( .A(n9033), .B(n8666), .Z(out[721]) );
  XOR U5680 ( .A(in[330]), .B(n8667), .Z(n9039) );
  NOR U5681 ( .A(n8834), .B(n9234), .Z(n8668) );
  XNOR U5682 ( .A(n9039), .B(n8668), .Z(out[722]) );
  XOR U5683 ( .A(in[331]), .B(n8669), .Z(n9041) );
  NOR U5684 ( .A(n8837), .B(n9238), .Z(n8670) );
  XNOR U5685 ( .A(n9041), .B(n8670), .Z(out[723]) );
  XOR U5686 ( .A(in[332]), .B(n8671), .Z(n9043) );
  NOR U5687 ( .A(n8840), .B(n9242), .Z(n8672) );
  XNOR U5688 ( .A(n9043), .B(n8672), .Z(out[724]) );
  XOR U5689 ( .A(in[333]), .B(n8673), .Z(n9045) );
  NOR U5690 ( .A(n8843), .B(n9246), .Z(n8674) );
  XNOR U5691 ( .A(n9045), .B(n8674), .Z(out[725]) );
  XOR U5692 ( .A(in[334]), .B(n8675), .Z(n9047) );
  NOR U5693 ( .A(n8850), .B(n9250), .Z(n8676) );
  XNOR U5694 ( .A(n9047), .B(n8676), .Z(out[726]) );
  XOR U5695 ( .A(in[335]), .B(n8677), .Z(n9049) );
  NOR U5696 ( .A(n8853), .B(n9254), .Z(n8678) );
  XNOR U5697 ( .A(n9049), .B(n8678), .Z(out[727]) );
  XOR U5698 ( .A(in[336]), .B(n8679), .Z(n9051) );
  NOR U5699 ( .A(n8856), .B(n9262), .Z(n8680) );
  XNOR U5700 ( .A(n9051), .B(n8680), .Z(out[728]) );
  XOR U5701 ( .A(in[337]), .B(n8681), .Z(n9053) );
  NOR U5702 ( .A(n8859), .B(n9266), .Z(n8682) );
  XNOR U5703 ( .A(n9053), .B(n8682), .Z(out[729]) );
  ANDN U5704 ( .B(n9168), .A(n9170), .Z(n8683) );
  XNOR U5705 ( .A(n8684), .B(n8683), .Z(out[72]) );
  XOR U5706 ( .A(in[338]), .B(n8685), .Z(n9055) );
  NOR U5707 ( .A(n8862), .B(n9270), .Z(n8686) );
  XNOR U5708 ( .A(n9055), .B(n8686), .Z(out[730]) );
  XOR U5709 ( .A(in[339]), .B(n8687), .Z(n9057) );
  NOR U5710 ( .A(n8865), .B(n9274), .Z(n8688) );
  XNOR U5711 ( .A(n9057), .B(n8688), .Z(out[731]) );
  XOR U5712 ( .A(in[340]), .B(n8689), .Z(n9063) );
  NOR U5713 ( .A(n8868), .B(n9278), .Z(n8690) );
  XNOR U5714 ( .A(n9063), .B(n8690), .Z(out[732]) );
  XOR U5715 ( .A(in[341]), .B(n8691), .Z(n9065) );
  NOR U5716 ( .A(n8871), .B(n9282), .Z(n8692) );
  XNOR U5717 ( .A(n9065), .B(n8692), .Z(out[733]) );
  XOR U5718 ( .A(in[342]), .B(n8693), .Z(n9067) );
  NOR U5719 ( .A(n8874), .B(n9286), .Z(n8694) );
  XNOR U5720 ( .A(n9067), .B(n8694), .Z(out[734]) );
  XOR U5721 ( .A(in[343]), .B(n8695), .Z(n9069) );
  NOR U5722 ( .A(n8877), .B(n9290), .Z(n8696) );
  XNOR U5723 ( .A(n9069), .B(n8696), .Z(out[735]) );
  XOR U5724 ( .A(in[344]), .B(n8697), .Z(n9071) );
  NOR U5725 ( .A(n8888), .B(n9294), .Z(n8698) );
  XNOR U5726 ( .A(n9071), .B(n8698), .Z(out[736]) );
  XOR U5727 ( .A(in[345]), .B(n8699), .Z(n9073) );
  NOR U5728 ( .A(n8891), .B(n9298), .Z(n8700) );
  XNOR U5729 ( .A(n9073), .B(n8700), .Z(out[737]) );
  XOR U5730 ( .A(in[346]), .B(n8701), .Z(n9075) );
  NOR U5731 ( .A(n8894), .B(n9306), .Z(n8702) );
  XNOR U5732 ( .A(n9075), .B(n8702), .Z(out[738]) );
  XOR U5733 ( .A(in[347]), .B(n8703), .Z(n9077) );
  NOR U5734 ( .A(n8897), .B(n9310), .Z(n8704) );
  XNOR U5735 ( .A(n9077), .B(n8704), .Z(out[739]) );
  ANDN U5736 ( .B(n9612), .A(n9614), .Z(n8705) );
  XNOR U5737 ( .A(n8706), .B(n8705), .Z(out[73]) );
  XOR U5738 ( .A(in[348]), .B(n8707), .Z(n9079) );
  NOR U5739 ( .A(n8900), .B(n9314), .Z(n8708) );
  XNOR U5740 ( .A(n9079), .B(n8708), .Z(out[740]) );
  XOR U5741 ( .A(in[349]), .B(n8709), .Z(n9081) );
  NOR U5742 ( .A(n8903), .B(n9318), .Z(n8710) );
  XNOR U5743 ( .A(n9081), .B(n8710), .Z(out[741]) );
  XOR U5744 ( .A(in[350]), .B(n8711), .Z(n9087) );
  NOR U5745 ( .A(n8906), .B(n9322), .Z(n8712) );
  XNOR U5746 ( .A(n9087), .B(n8712), .Z(out[742]) );
  XOR U5747 ( .A(in[351]), .B(n8713), .Z(n9089) );
  NOR U5748 ( .A(n8909), .B(n9326), .Z(n8714) );
  XNOR U5749 ( .A(n9089), .B(n8714), .Z(out[743]) );
  XOR U5750 ( .A(in[352]), .B(n8715), .Z(n9091) );
  NOR U5751 ( .A(n8912), .B(n9330), .Z(n8716) );
  XNOR U5752 ( .A(n9091), .B(n8716), .Z(out[744]) );
  XOR U5753 ( .A(in[353]), .B(n8717), .Z(n9093) );
  NOR U5754 ( .A(n8915), .B(n9334), .Z(n8718) );
  XNOR U5755 ( .A(n9093), .B(n8718), .Z(out[745]) );
  XOR U5756 ( .A(in[354]), .B(n8719), .Z(n9095) );
  NOR U5757 ( .A(n8922), .B(n9338), .Z(n8720) );
  XNOR U5758 ( .A(n9095), .B(n8720), .Z(out[746]) );
  XOR U5759 ( .A(in[355]), .B(n8721), .Z(n9097) );
  NOR U5760 ( .A(n8925), .B(n9342), .Z(n8722) );
  XNOR U5761 ( .A(n9097), .B(n8722), .Z(out[747]) );
  XOR U5762 ( .A(in[356]), .B(n8723), .Z(n9099) );
  NOR U5763 ( .A(n8928), .B(n9350), .Z(n8724) );
  XNOR U5764 ( .A(n9099), .B(n8724), .Z(out[748]) );
  XOR U5765 ( .A(in[357]), .B(n8725), .Z(n9101) );
  NOR U5766 ( .A(n8931), .B(n9354), .Z(n8726) );
  XNOR U5767 ( .A(n9101), .B(n8726), .Z(out[749]) );
  NOR U5768 ( .A(n8728), .B(n8727), .Z(n8729) );
  XNOR U5769 ( .A(n8730), .B(n8729), .Z(out[74]) );
  XOR U5770 ( .A(in[358]), .B(n8731), .Z(n9103) );
  NOR U5771 ( .A(n8934), .B(n9358), .Z(n8732) );
  XNOR U5772 ( .A(n9103), .B(n8732), .Z(out[750]) );
  XOR U5773 ( .A(in[359]), .B(n8733), .Z(n9105) );
  NOR U5774 ( .A(n8937), .B(n9362), .Z(n8734) );
  XNOR U5775 ( .A(n9105), .B(n8734), .Z(out[751]) );
  XOR U5776 ( .A(in[360]), .B(n8735), .Z(n9111) );
  NOR U5777 ( .A(n8940), .B(n9366), .Z(n8736) );
  XNOR U5778 ( .A(n9111), .B(n8736), .Z(out[752]) );
  XOR U5779 ( .A(in[361]), .B(n8737), .Z(n9113) );
  NOR U5780 ( .A(n8943), .B(n9370), .Z(n8738) );
  XNOR U5781 ( .A(n9113), .B(n8738), .Z(out[753]) );
  XOR U5782 ( .A(in[362]), .B(n8739), .Z(n9115) );
  NOR U5783 ( .A(n8946), .B(n9374), .Z(n8740) );
  XNOR U5784 ( .A(n9115), .B(n8740), .Z(out[754]) );
  XOR U5785 ( .A(in[363]), .B(n8741), .Z(n9117) );
  NOR U5786 ( .A(n8949), .B(n9378), .Z(n8742) );
  XNOR U5787 ( .A(n9117), .B(n8742), .Z(out[755]) );
  XOR U5788 ( .A(in[364]), .B(n8743), .Z(n9119) );
  NOR U5789 ( .A(n8956), .B(n9382), .Z(n8744) );
  XNOR U5790 ( .A(n9119), .B(n8744), .Z(out[756]) );
  XOR U5791 ( .A(in[365]), .B(n8745), .Z(n9121) );
  NOR U5792 ( .A(n8959), .B(n9386), .Z(n8746) );
  XNOR U5793 ( .A(n9121), .B(n8746), .Z(out[757]) );
  XOR U5794 ( .A(in[366]), .B(n8747), .Z(n9123) );
  NOR U5795 ( .A(n8962), .B(n9394), .Z(n8748) );
  XNOR U5796 ( .A(n9123), .B(n8748), .Z(out[758]) );
  XOR U5797 ( .A(in[367]), .B(n8749), .Z(n9125) );
  NOR U5798 ( .A(n8965), .B(n9398), .Z(n8750) );
  XNOR U5799 ( .A(n9125), .B(n8750), .Z(out[759]) );
  NOR U5800 ( .A(n8752), .B(n8751), .Z(n8753) );
  XNOR U5801 ( .A(n8754), .B(n8753), .Z(out[75]) );
  XOR U5802 ( .A(in[368]), .B(n8755), .Z(n9127) );
  NOR U5803 ( .A(n8968), .B(n9402), .Z(n8756) );
  XNOR U5804 ( .A(n9127), .B(n8756), .Z(out[760]) );
  XOR U5805 ( .A(in[369]), .B(n8757), .Z(n9129) );
  NOR U5806 ( .A(n8971), .B(n9406), .Z(n8758) );
  XNOR U5807 ( .A(n9129), .B(n8758), .Z(out[761]) );
  XOR U5808 ( .A(in[370]), .B(n8759), .Z(n9135) );
  NOR U5809 ( .A(n8974), .B(n9410), .Z(n8760) );
  XNOR U5810 ( .A(n9135), .B(n8760), .Z(out[762]) );
  XOR U5811 ( .A(in[371]), .B(n8761), .Z(n9137) );
  NOR U5812 ( .A(n8977), .B(n9414), .Z(n8762) );
  XNOR U5813 ( .A(n9137), .B(n8762), .Z(out[763]) );
  XOR U5814 ( .A(in[372]), .B(n8763), .Z(n9139) );
  NOR U5815 ( .A(n8980), .B(n9418), .Z(n8764) );
  XNOR U5816 ( .A(n9139), .B(n8764), .Z(out[764]) );
  XOR U5817 ( .A(in[373]), .B(n8765), .Z(n9141) );
  NOR U5818 ( .A(n8983), .B(n9422), .Z(n8766) );
  XNOR U5819 ( .A(n9141), .B(n8766), .Z(out[765]) );
  XOR U5820 ( .A(in[374]), .B(n8767), .Z(n9143) );
  NOR U5821 ( .A(n8990), .B(n9426), .Z(n8768) );
  XNOR U5822 ( .A(n9143), .B(n8768), .Z(out[766]) );
  XOR U5823 ( .A(in[375]), .B(n8769), .Z(n9145) );
  NOR U5824 ( .A(n8993), .B(n9430), .Z(n8770) );
  XNOR U5825 ( .A(n9145), .B(n8770), .Z(out[767]) );
  XNOR U5826 ( .A(in[743]), .B(n8771), .Z(n9148) );
  NAND U5827 ( .A(n8995), .B(n8772), .Z(n8773) );
  XNOR U5828 ( .A(n9148), .B(n8773), .Z(out[768]) );
  XNOR U5829 ( .A(in[744]), .B(n8774), .Z(n9152) );
  NAND U5830 ( .A(n8997), .B(n8775), .Z(n8776) );
  XNOR U5831 ( .A(n9152), .B(n8776), .Z(out[769]) );
  NOR U5832 ( .A(n8778), .B(n8777), .Z(n8779) );
  XNOR U5833 ( .A(n8780), .B(n8779), .Z(out[76]) );
  XNOR U5834 ( .A(in[745]), .B(n8781), .Z(n9156) );
  NAND U5835 ( .A(n8999), .B(n8782), .Z(n8783) );
  XNOR U5836 ( .A(n9156), .B(n8783), .Z(out[770]) );
  XNOR U5837 ( .A(in[746]), .B(n8784), .Z(n9160) );
  NAND U5838 ( .A(n9001), .B(n8785), .Z(n8786) );
  XNOR U5839 ( .A(n9160), .B(n8786), .Z(out[771]) );
  XNOR U5840 ( .A(in[747]), .B(n8787), .Z(n9172) );
  NAND U5841 ( .A(n9003), .B(n8788), .Z(n8789) );
  XNOR U5842 ( .A(n9172), .B(n8789), .Z(out[772]) );
  XNOR U5843 ( .A(in[748]), .B(n8790), .Z(n9176) );
  NAND U5844 ( .A(n9005), .B(n8791), .Z(n8792) );
  XNOR U5845 ( .A(n9176), .B(n8792), .Z(out[773]) );
  XNOR U5846 ( .A(in[749]), .B(n8793), .Z(n9180) );
  NAND U5847 ( .A(n9007), .B(n8794), .Z(n8795) );
  XNOR U5848 ( .A(n9180), .B(n8795), .Z(out[774]) );
  XNOR U5849 ( .A(in[750]), .B(n8796), .Z(n9184) );
  NAND U5850 ( .A(n9009), .B(n8797), .Z(n8798) );
  XNOR U5851 ( .A(n9184), .B(n8798), .Z(out[775]) );
  XNOR U5852 ( .A(in[751]), .B(n8799), .Z(n9188) );
  NAND U5853 ( .A(n9015), .B(n8800), .Z(n8801) );
  XNOR U5854 ( .A(n9188), .B(n8801), .Z(out[776]) );
  XNOR U5855 ( .A(in[752]), .B(n8802), .Z(n9192) );
  NAND U5856 ( .A(n9017), .B(n8803), .Z(n8804) );
  XNOR U5857 ( .A(n9192), .B(n8804), .Z(out[777]) );
  XNOR U5858 ( .A(in[753]), .B(n8805), .Z(n9196) );
  NAND U5859 ( .A(n9019), .B(n8806), .Z(n8807) );
  XNOR U5860 ( .A(n9196), .B(n8807), .Z(out[778]) );
  XNOR U5861 ( .A(in[754]), .B(n8808), .Z(n9200) );
  NAND U5862 ( .A(n9021), .B(n8809), .Z(n8810) );
  XNOR U5863 ( .A(n9200), .B(n8810), .Z(out[779]) );
  NOR U5864 ( .A(n8812), .B(n8811), .Z(n8813) );
  XNOR U5865 ( .A(n8814), .B(n8813), .Z(out[77]) );
  XNOR U5866 ( .A(in[755]), .B(n8815), .Z(n9204) );
  NAND U5867 ( .A(n9023), .B(n8816), .Z(n8817) );
  XNOR U5868 ( .A(n9204), .B(n8817), .Z(out[780]) );
  XNOR U5869 ( .A(in[756]), .B(n8818), .Z(n9208) );
  NAND U5870 ( .A(n9025), .B(n8819), .Z(n8820) );
  XNOR U5871 ( .A(n9208), .B(n8820), .Z(out[781]) );
  XNOR U5872 ( .A(in[757]), .B(n8821), .Z(n9216) );
  NAND U5873 ( .A(n9027), .B(n8822), .Z(n8823) );
  XNOR U5874 ( .A(n9216), .B(n8823), .Z(out[782]) );
  XNOR U5875 ( .A(in[758]), .B(n8824), .Z(n9220) );
  NAND U5876 ( .A(n9029), .B(n8825), .Z(n8826) );
  XNOR U5877 ( .A(n9220), .B(n8826), .Z(out[783]) );
  XNOR U5878 ( .A(in[759]), .B(n8827), .Z(n9224) );
  NAND U5879 ( .A(n9031), .B(n8828), .Z(n8829) );
  XNOR U5880 ( .A(n9224), .B(n8829), .Z(out[784]) );
  XNOR U5881 ( .A(in[760]), .B(n8830), .Z(n9228) );
  NAND U5882 ( .A(n9033), .B(n8831), .Z(n8832) );
  XNOR U5883 ( .A(n9228), .B(n8832), .Z(out[785]) );
  XNOR U5884 ( .A(in[761]), .B(n8833), .Z(n9232) );
  NAND U5885 ( .A(n9039), .B(n8834), .Z(n8835) );
  XNOR U5886 ( .A(n9232), .B(n8835), .Z(out[786]) );
  XNOR U5887 ( .A(in[762]), .B(n8836), .Z(n9236) );
  NAND U5888 ( .A(n9041), .B(n8837), .Z(n8838) );
  XNOR U5889 ( .A(n9236), .B(n8838), .Z(out[787]) );
  XNOR U5890 ( .A(in[763]), .B(n8839), .Z(n9240) );
  NAND U5891 ( .A(n9043), .B(n8840), .Z(n8841) );
  XNOR U5892 ( .A(n9240), .B(n8841), .Z(out[788]) );
  XNOR U5893 ( .A(in[764]), .B(n8842), .Z(n9244) );
  NAND U5894 ( .A(n9045), .B(n8843), .Z(n8844) );
  XNOR U5895 ( .A(n9244), .B(n8844), .Z(out[789]) );
  NOR U5896 ( .A(n8846), .B(n8845), .Z(n8847) );
  XNOR U5897 ( .A(n8848), .B(n8847), .Z(out[78]) );
  XNOR U5898 ( .A(in[765]), .B(n8849), .Z(n9248) );
  NAND U5899 ( .A(n9047), .B(n8850), .Z(n8851) );
  XNOR U5900 ( .A(n9248), .B(n8851), .Z(out[790]) );
  XNOR U5901 ( .A(in[766]), .B(n8852), .Z(n9252) );
  NAND U5902 ( .A(n9049), .B(n8853), .Z(n8854) );
  XNOR U5903 ( .A(n9252), .B(n8854), .Z(out[791]) );
  XNOR U5904 ( .A(in[767]), .B(n8855), .Z(n9260) );
  NAND U5905 ( .A(n9051), .B(n8856), .Z(n8857) );
  XNOR U5906 ( .A(n9260), .B(n8857), .Z(out[792]) );
  XNOR U5907 ( .A(in[704]), .B(n8858), .Z(n9264) );
  NAND U5908 ( .A(n9053), .B(n8859), .Z(n8860) );
  XNOR U5909 ( .A(n9264), .B(n8860), .Z(out[793]) );
  XNOR U5910 ( .A(in[705]), .B(n8861), .Z(n9268) );
  NAND U5911 ( .A(n9055), .B(n8862), .Z(n8863) );
  XNOR U5912 ( .A(n9268), .B(n8863), .Z(out[794]) );
  XNOR U5913 ( .A(in[706]), .B(n8864), .Z(n9272) );
  NAND U5914 ( .A(n9057), .B(n8865), .Z(n8866) );
  XNOR U5915 ( .A(n9272), .B(n8866), .Z(out[795]) );
  XNOR U5916 ( .A(in[707]), .B(n8867), .Z(n9276) );
  NAND U5917 ( .A(n9063), .B(n8868), .Z(n8869) );
  XNOR U5918 ( .A(n9276), .B(n8869), .Z(out[796]) );
  XNOR U5919 ( .A(in[708]), .B(n8870), .Z(n9280) );
  NAND U5920 ( .A(n9065), .B(n8871), .Z(n8872) );
  XNOR U5921 ( .A(n9280), .B(n8872), .Z(out[797]) );
  XNOR U5922 ( .A(in[709]), .B(n8873), .Z(n9284) );
  NAND U5923 ( .A(n9067), .B(n8874), .Z(n8875) );
  XNOR U5924 ( .A(n9284), .B(n8875), .Z(out[798]) );
  XNOR U5925 ( .A(in[710]), .B(n8876), .Z(n9288) );
  NAND U5926 ( .A(n9069), .B(n8877), .Z(n8878) );
  XNOR U5927 ( .A(n9288), .B(n8878), .Z(out[799]) );
  NOR U5928 ( .A(n8880), .B(n8879), .Z(n8881) );
  XNOR U5929 ( .A(n8882), .B(n8881), .Z(out[79]) );
  OR U5930 ( .A(n8884), .B(n8883), .Z(n8885) );
  XNOR U5931 ( .A(n8886), .B(n8885), .Z(out[7]) );
  XNOR U5932 ( .A(in[711]), .B(n8887), .Z(n9292) );
  NAND U5933 ( .A(n9071), .B(n8888), .Z(n8889) );
  XNOR U5934 ( .A(n9292), .B(n8889), .Z(out[800]) );
  XNOR U5935 ( .A(in[712]), .B(n8890), .Z(n9296) );
  NAND U5936 ( .A(n9073), .B(n8891), .Z(n8892) );
  XNOR U5937 ( .A(n9296), .B(n8892), .Z(out[801]) );
  XNOR U5938 ( .A(in[713]), .B(n8893), .Z(n9304) );
  NAND U5939 ( .A(n9075), .B(n8894), .Z(n8895) );
  XNOR U5940 ( .A(n9304), .B(n8895), .Z(out[802]) );
  XNOR U5941 ( .A(in[714]), .B(n8896), .Z(n9308) );
  NAND U5942 ( .A(n9077), .B(n8897), .Z(n8898) );
  XNOR U5943 ( .A(n9308), .B(n8898), .Z(out[803]) );
  XNOR U5944 ( .A(in[715]), .B(n8899), .Z(n9312) );
  NAND U5945 ( .A(n9079), .B(n8900), .Z(n8901) );
  XNOR U5946 ( .A(n9312), .B(n8901), .Z(out[804]) );
  XOR U5947 ( .A(n8902), .B(in[716]), .Z(n9316) );
  NAND U5948 ( .A(n9081), .B(n8903), .Z(n8904) );
  XNOR U5949 ( .A(n9316), .B(n8904), .Z(out[805]) );
  XOR U5950 ( .A(n8905), .B(in[717]), .Z(n9320) );
  NAND U5951 ( .A(n9087), .B(n8906), .Z(n8907) );
  XNOR U5952 ( .A(n9320), .B(n8907), .Z(out[806]) );
  XOR U5953 ( .A(n8908), .B(in[718]), .Z(n9324) );
  NAND U5954 ( .A(n9089), .B(n8909), .Z(n8910) );
  XNOR U5955 ( .A(n9324), .B(n8910), .Z(out[807]) );
  XOR U5956 ( .A(n8911), .B(in[719]), .Z(n9328) );
  NAND U5957 ( .A(n9091), .B(n8912), .Z(n8913) );
  XNOR U5958 ( .A(n9328), .B(n8913), .Z(out[808]) );
  XOR U5959 ( .A(n8914), .B(in[720]), .Z(n9332) );
  NAND U5960 ( .A(n9093), .B(n8915), .Z(n8916) );
  XNOR U5961 ( .A(n9332), .B(n8916), .Z(out[809]) );
  NOR U5962 ( .A(n8918), .B(n8917), .Z(n8919) );
  XNOR U5963 ( .A(n8920), .B(n8919), .Z(out[80]) );
  XOR U5964 ( .A(n8921), .B(in[721]), .Z(n9336) );
  NAND U5965 ( .A(n9095), .B(n8922), .Z(n8923) );
  XNOR U5966 ( .A(n9336), .B(n8923), .Z(out[810]) );
  XOR U5967 ( .A(n8924), .B(in[722]), .Z(n9340) );
  NAND U5968 ( .A(n9097), .B(n8925), .Z(n8926) );
  XNOR U5969 ( .A(n9340), .B(n8926), .Z(out[811]) );
  XOR U5970 ( .A(n8927), .B(in[723]), .Z(n9348) );
  NAND U5971 ( .A(n9099), .B(n8928), .Z(n8929) );
  XNOR U5972 ( .A(n9348), .B(n8929), .Z(out[812]) );
  XOR U5973 ( .A(in[724]), .B(n8930), .Z(n9352) );
  NAND U5974 ( .A(n9101), .B(n8931), .Z(n8932) );
  XNOR U5975 ( .A(n9352), .B(n8932), .Z(out[813]) );
  XOR U5976 ( .A(in[725]), .B(n8933), .Z(n9356) );
  NAND U5977 ( .A(n9103), .B(n8934), .Z(n8935) );
  XNOR U5978 ( .A(n9356), .B(n8935), .Z(out[814]) );
  XOR U5979 ( .A(in[726]), .B(n8936), .Z(n9360) );
  NAND U5980 ( .A(n9105), .B(n8937), .Z(n8938) );
  XNOR U5981 ( .A(n9360), .B(n8938), .Z(out[815]) );
  XOR U5982 ( .A(in[727]), .B(n8939), .Z(n9364) );
  NAND U5983 ( .A(n9111), .B(n8940), .Z(n8941) );
  XNOR U5984 ( .A(n9364), .B(n8941), .Z(out[816]) );
  XOR U5985 ( .A(in[728]), .B(n8942), .Z(n9368) );
  NAND U5986 ( .A(n9113), .B(n8943), .Z(n8944) );
  XNOR U5987 ( .A(n9368), .B(n8944), .Z(out[817]) );
  XOR U5988 ( .A(in[729]), .B(n8945), .Z(n9372) );
  NAND U5989 ( .A(n9115), .B(n8946), .Z(n8947) );
  XNOR U5990 ( .A(n9372), .B(n8947), .Z(out[818]) );
  XOR U5991 ( .A(in[730]), .B(n8948), .Z(n9376) );
  NAND U5992 ( .A(n9117), .B(n8949), .Z(n8950) );
  XNOR U5993 ( .A(n9376), .B(n8950), .Z(out[819]) );
  NOR U5994 ( .A(n8952), .B(n8951), .Z(n8953) );
  XNOR U5995 ( .A(n8954), .B(n8953), .Z(out[81]) );
  XOR U5996 ( .A(in[731]), .B(n8955), .Z(n9380) );
  NAND U5997 ( .A(n9119), .B(n8956), .Z(n8957) );
  XNOR U5998 ( .A(n9380), .B(n8957), .Z(out[820]) );
  XOR U5999 ( .A(in[732]), .B(n8958), .Z(n9384) );
  NAND U6000 ( .A(n9121), .B(n8959), .Z(n8960) );
  XNOR U6001 ( .A(n9384), .B(n8960), .Z(out[821]) );
  XOR U6002 ( .A(in[733]), .B(n8961), .Z(n9392) );
  NAND U6003 ( .A(n9123), .B(n8962), .Z(n8963) );
  XNOR U6004 ( .A(n9392), .B(n8963), .Z(out[822]) );
  XOR U6005 ( .A(in[734]), .B(n8964), .Z(n9396) );
  NAND U6006 ( .A(n9125), .B(n8965), .Z(n8966) );
  XNOR U6007 ( .A(n9396), .B(n8966), .Z(out[823]) );
  XOR U6008 ( .A(in[735]), .B(n8967), .Z(n9400) );
  NAND U6009 ( .A(n9127), .B(n8968), .Z(n8969) );
  XNOR U6010 ( .A(n9400), .B(n8969), .Z(out[824]) );
  XOR U6011 ( .A(in[736]), .B(n8970), .Z(n9404) );
  NAND U6012 ( .A(n9129), .B(n8971), .Z(n8972) );
  XNOR U6013 ( .A(n9404), .B(n8972), .Z(out[825]) );
  XOR U6014 ( .A(in[737]), .B(n8973), .Z(n9408) );
  NAND U6015 ( .A(n9135), .B(n8974), .Z(n8975) );
  XNOR U6016 ( .A(n9408), .B(n8975), .Z(out[826]) );
  XOR U6017 ( .A(in[738]), .B(n8976), .Z(n9412) );
  NAND U6018 ( .A(n9137), .B(n8977), .Z(n8978) );
  XNOR U6019 ( .A(n9412), .B(n8978), .Z(out[827]) );
  XOR U6020 ( .A(in[739]), .B(n8979), .Z(n9416) );
  NAND U6021 ( .A(n9139), .B(n8980), .Z(n8981) );
  XNOR U6022 ( .A(n9416), .B(n8981), .Z(out[828]) );
  XNOR U6023 ( .A(in[740]), .B(n8982), .Z(n9420) );
  NAND U6024 ( .A(n9141), .B(n8983), .Z(n8984) );
  XNOR U6025 ( .A(n9420), .B(n8984), .Z(out[829]) );
  NOR U6026 ( .A(n8986), .B(n8985), .Z(n8987) );
  XNOR U6027 ( .A(n8988), .B(n8987), .Z(out[82]) );
  XNOR U6028 ( .A(in[741]), .B(n8989), .Z(n9424) );
  NAND U6029 ( .A(n9143), .B(n8990), .Z(n8991) );
  XNOR U6030 ( .A(n9424), .B(n8991), .Z(out[830]) );
  XNOR U6031 ( .A(in[742]), .B(n8992), .Z(n9428) );
  NAND U6032 ( .A(n9145), .B(n8993), .Z(n8994) );
  XNOR U6033 ( .A(n9428), .B(n8994), .Z(out[831]) );
  OR U6034 ( .A(n9148), .B(n8995), .Z(n8996) );
  XNOR U6035 ( .A(n9147), .B(n8996), .Z(out[832]) );
  OR U6036 ( .A(n9152), .B(n8997), .Z(n8998) );
  XNOR U6037 ( .A(n9151), .B(n8998), .Z(out[833]) );
  OR U6038 ( .A(n9156), .B(n8999), .Z(n9000) );
  XNOR U6039 ( .A(n9155), .B(n9000), .Z(out[834]) );
  OR U6040 ( .A(n9160), .B(n9001), .Z(n9002) );
  XNOR U6041 ( .A(n9159), .B(n9002), .Z(out[835]) );
  OR U6042 ( .A(n9172), .B(n9003), .Z(n9004) );
  XNOR U6043 ( .A(n9171), .B(n9004), .Z(out[836]) );
  OR U6044 ( .A(n9176), .B(n9005), .Z(n9006) );
  XNOR U6045 ( .A(n9175), .B(n9006), .Z(out[837]) );
  OR U6046 ( .A(n9180), .B(n9007), .Z(n9008) );
  XNOR U6047 ( .A(n9179), .B(n9008), .Z(out[838]) );
  OR U6048 ( .A(n9184), .B(n9009), .Z(n9010) );
  XNOR U6049 ( .A(n9183), .B(n9010), .Z(out[839]) );
  NOR U6050 ( .A(n9012), .B(n9011), .Z(n9013) );
  XNOR U6051 ( .A(n9014), .B(n9013), .Z(out[83]) );
  OR U6052 ( .A(n9188), .B(n9015), .Z(n9016) );
  XNOR U6053 ( .A(n9187), .B(n9016), .Z(out[840]) );
  OR U6054 ( .A(n9192), .B(n9017), .Z(n9018) );
  XNOR U6055 ( .A(n9191), .B(n9018), .Z(out[841]) );
  OR U6056 ( .A(n9196), .B(n9019), .Z(n9020) );
  XNOR U6057 ( .A(n9195), .B(n9020), .Z(out[842]) );
  OR U6058 ( .A(n9200), .B(n9021), .Z(n9022) );
  XNOR U6059 ( .A(n9199), .B(n9022), .Z(out[843]) );
  OR U6060 ( .A(n9204), .B(n9023), .Z(n9024) );
  XNOR U6061 ( .A(n9203), .B(n9024), .Z(out[844]) );
  OR U6062 ( .A(n9208), .B(n9025), .Z(n9026) );
  XNOR U6063 ( .A(n9207), .B(n9026), .Z(out[845]) );
  OR U6064 ( .A(n9216), .B(n9027), .Z(n9028) );
  XNOR U6065 ( .A(n9215), .B(n9028), .Z(out[846]) );
  OR U6066 ( .A(n9220), .B(n9029), .Z(n9030) );
  XNOR U6067 ( .A(n9219), .B(n9030), .Z(out[847]) );
  OR U6068 ( .A(n9224), .B(n9031), .Z(n9032) );
  XNOR U6069 ( .A(n9223), .B(n9032), .Z(out[848]) );
  OR U6070 ( .A(n9228), .B(n9033), .Z(n9034) );
  XNOR U6071 ( .A(n9227), .B(n9034), .Z(out[849]) );
  NOR U6072 ( .A(n9036), .B(n9035), .Z(n9037) );
  XNOR U6073 ( .A(n9038), .B(n9037), .Z(out[84]) );
  OR U6074 ( .A(n9232), .B(n9039), .Z(n9040) );
  XNOR U6075 ( .A(n9231), .B(n9040), .Z(out[850]) );
  OR U6076 ( .A(n9236), .B(n9041), .Z(n9042) );
  XNOR U6077 ( .A(n9235), .B(n9042), .Z(out[851]) );
  OR U6078 ( .A(n9240), .B(n9043), .Z(n9044) );
  XNOR U6079 ( .A(n9239), .B(n9044), .Z(out[852]) );
  OR U6080 ( .A(n9244), .B(n9045), .Z(n9046) );
  XNOR U6081 ( .A(n9243), .B(n9046), .Z(out[853]) );
  OR U6082 ( .A(n9248), .B(n9047), .Z(n9048) );
  XNOR U6083 ( .A(n9247), .B(n9048), .Z(out[854]) );
  OR U6084 ( .A(n9252), .B(n9049), .Z(n9050) );
  XNOR U6085 ( .A(n9251), .B(n9050), .Z(out[855]) );
  OR U6086 ( .A(n9260), .B(n9051), .Z(n9052) );
  XNOR U6087 ( .A(n9259), .B(n9052), .Z(out[856]) );
  OR U6088 ( .A(n9264), .B(n9053), .Z(n9054) );
  XNOR U6089 ( .A(n9263), .B(n9054), .Z(out[857]) );
  OR U6090 ( .A(n9268), .B(n9055), .Z(n9056) );
  XNOR U6091 ( .A(n9267), .B(n9056), .Z(out[858]) );
  OR U6092 ( .A(n9272), .B(n9057), .Z(n9058) );
  XNOR U6093 ( .A(n9271), .B(n9058), .Z(out[859]) );
  NOR U6094 ( .A(n9060), .B(n9059), .Z(n9061) );
  XNOR U6095 ( .A(n9062), .B(n9061), .Z(out[85]) );
  OR U6096 ( .A(n9276), .B(n9063), .Z(n9064) );
  XNOR U6097 ( .A(n9275), .B(n9064), .Z(out[860]) );
  OR U6098 ( .A(n9280), .B(n9065), .Z(n9066) );
  XNOR U6099 ( .A(n9279), .B(n9066), .Z(out[861]) );
  OR U6100 ( .A(n9284), .B(n9067), .Z(n9068) );
  XNOR U6101 ( .A(n9283), .B(n9068), .Z(out[862]) );
  OR U6102 ( .A(n9288), .B(n9069), .Z(n9070) );
  XNOR U6103 ( .A(n9287), .B(n9070), .Z(out[863]) );
  OR U6104 ( .A(n9292), .B(n9071), .Z(n9072) );
  XNOR U6105 ( .A(n9291), .B(n9072), .Z(out[864]) );
  OR U6106 ( .A(n9296), .B(n9073), .Z(n9074) );
  XNOR U6107 ( .A(n9295), .B(n9074), .Z(out[865]) );
  OR U6108 ( .A(n9304), .B(n9075), .Z(n9076) );
  XNOR U6109 ( .A(n9303), .B(n9076), .Z(out[866]) );
  OR U6110 ( .A(n9308), .B(n9077), .Z(n9078) );
  XNOR U6111 ( .A(n9307), .B(n9078), .Z(out[867]) );
  OR U6112 ( .A(n9312), .B(n9079), .Z(n9080) );
  XNOR U6113 ( .A(n9311), .B(n9080), .Z(out[868]) );
  OR U6114 ( .A(n9316), .B(n9081), .Z(n9082) );
  XNOR U6115 ( .A(n9315), .B(n9082), .Z(out[869]) );
  NOR U6116 ( .A(n9084), .B(n9083), .Z(n9085) );
  XNOR U6117 ( .A(n9086), .B(n9085), .Z(out[86]) );
  OR U6118 ( .A(n9320), .B(n9087), .Z(n9088) );
  XNOR U6119 ( .A(n9319), .B(n9088), .Z(out[870]) );
  OR U6120 ( .A(n9324), .B(n9089), .Z(n9090) );
  XNOR U6121 ( .A(n9323), .B(n9090), .Z(out[871]) );
  OR U6122 ( .A(n9328), .B(n9091), .Z(n9092) );
  XNOR U6123 ( .A(n9327), .B(n9092), .Z(out[872]) );
  OR U6124 ( .A(n9332), .B(n9093), .Z(n9094) );
  XNOR U6125 ( .A(n9331), .B(n9094), .Z(out[873]) );
  OR U6126 ( .A(n9336), .B(n9095), .Z(n9096) );
  XNOR U6127 ( .A(n9335), .B(n9096), .Z(out[874]) );
  OR U6128 ( .A(n9340), .B(n9097), .Z(n9098) );
  XNOR U6129 ( .A(n9339), .B(n9098), .Z(out[875]) );
  OR U6130 ( .A(n9348), .B(n9099), .Z(n9100) );
  XNOR U6131 ( .A(n9347), .B(n9100), .Z(out[876]) );
  OR U6132 ( .A(n9352), .B(n9101), .Z(n9102) );
  XNOR U6133 ( .A(n9351), .B(n9102), .Z(out[877]) );
  OR U6134 ( .A(n9356), .B(n9103), .Z(n9104) );
  XNOR U6135 ( .A(n9355), .B(n9104), .Z(out[878]) );
  OR U6136 ( .A(n9360), .B(n9105), .Z(n9106) );
  XNOR U6137 ( .A(n9359), .B(n9106), .Z(out[879]) );
  NOR U6138 ( .A(n9108), .B(n9107), .Z(n9109) );
  XNOR U6139 ( .A(n9110), .B(n9109), .Z(out[87]) );
  OR U6140 ( .A(n9364), .B(n9111), .Z(n9112) );
  XNOR U6141 ( .A(n9363), .B(n9112), .Z(out[880]) );
  OR U6142 ( .A(n9368), .B(n9113), .Z(n9114) );
  XNOR U6143 ( .A(n9367), .B(n9114), .Z(out[881]) );
  OR U6144 ( .A(n9372), .B(n9115), .Z(n9116) );
  XNOR U6145 ( .A(n9371), .B(n9116), .Z(out[882]) );
  OR U6146 ( .A(n9376), .B(n9117), .Z(n9118) );
  XNOR U6147 ( .A(n9375), .B(n9118), .Z(out[883]) );
  OR U6148 ( .A(n9380), .B(n9119), .Z(n9120) );
  XNOR U6149 ( .A(n9379), .B(n9120), .Z(out[884]) );
  OR U6150 ( .A(n9384), .B(n9121), .Z(n9122) );
  XNOR U6151 ( .A(n9383), .B(n9122), .Z(out[885]) );
  OR U6152 ( .A(n9392), .B(n9123), .Z(n9124) );
  XNOR U6153 ( .A(n9391), .B(n9124), .Z(out[886]) );
  OR U6154 ( .A(n9396), .B(n9125), .Z(n9126) );
  XNOR U6155 ( .A(n9395), .B(n9126), .Z(out[887]) );
  OR U6156 ( .A(n9400), .B(n9127), .Z(n9128) );
  XNOR U6157 ( .A(n9399), .B(n9128), .Z(out[888]) );
  OR U6158 ( .A(n9404), .B(n9129), .Z(n9130) );
  XNOR U6159 ( .A(n9403), .B(n9130), .Z(out[889]) );
  NOR U6160 ( .A(n9132), .B(n9131), .Z(n9133) );
  XNOR U6161 ( .A(n9134), .B(n9133), .Z(out[88]) );
  OR U6162 ( .A(n9408), .B(n9135), .Z(n9136) );
  XNOR U6163 ( .A(n9407), .B(n9136), .Z(out[890]) );
  OR U6164 ( .A(n9412), .B(n9137), .Z(n9138) );
  XNOR U6165 ( .A(n9411), .B(n9138), .Z(out[891]) );
  OR U6166 ( .A(n9416), .B(n9139), .Z(n9140) );
  XNOR U6167 ( .A(n9415), .B(n9140), .Z(out[892]) );
  OR U6168 ( .A(n9420), .B(n9141), .Z(n9142) );
  XNOR U6169 ( .A(n9419), .B(n9142), .Z(out[893]) );
  OR U6170 ( .A(n9424), .B(n9143), .Z(n9144) );
  XNOR U6171 ( .A(n9423), .B(n9144), .Z(out[894]) );
  OR U6172 ( .A(n9428), .B(n9145), .Z(n9146) );
  XNOR U6173 ( .A(n9427), .B(n9146), .Z(out[895]) );
  ANDN U6174 ( .B(n9148), .A(n9147), .Z(n9149) );
  XNOR U6175 ( .A(n9150), .B(n9149), .Z(out[896]) );
  ANDN U6176 ( .B(n9152), .A(n9151), .Z(n9153) );
  XNOR U6177 ( .A(n9154), .B(n9153), .Z(out[897]) );
  ANDN U6178 ( .B(n9156), .A(n9155), .Z(n9157) );
  XNOR U6179 ( .A(n9158), .B(n9157), .Z(out[898]) );
  ANDN U6180 ( .B(n9160), .A(n9159), .Z(n9161) );
  XNOR U6181 ( .A(n9162), .B(n9161), .Z(out[899]) );
  NOR U6182 ( .A(n9164), .B(n9163), .Z(n9165) );
  XNOR U6183 ( .A(n9166), .B(n9165), .Z(out[89]) );
  OR U6184 ( .A(n9168), .B(n9167), .Z(n9169) );
  XNOR U6185 ( .A(n9170), .B(n9169), .Z(out[8]) );
  ANDN U6186 ( .B(n9172), .A(n9171), .Z(n9173) );
  XNOR U6187 ( .A(n9174), .B(n9173), .Z(out[900]) );
  ANDN U6188 ( .B(n9176), .A(n9175), .Z(n9177) );
  XNOR U6189 ( .A(n9178), .B(n9177), .Z(out[901]) );
  ANDN U6190 ( .B(n9180), .A(n9179), .Z(n9181) );
  XNOR U6191 ( .A(n9182), .B(n9181), .Z(out[902]) );
  ANDN U6192 ( .B(n9184), .A(n9183), .Z(n9185) );
  XNOR U6193 ( .A(n9186), .B(n9185), .Z(out[903]) );
  ANDN U6194 ( .B(n9188), .A(n9187), .Z(n9189) );
  XNOR U6195 ( .A(n9190), .B(n9189), .Z(out[904]) );
  ANDN U6196 ( .B(n9192), .A(n9191), .Z(n9193) );
  XNOR U6197 ( .A(n9194), .B(n9193), .Z(out[905]) );
  ANDN U6198 ( .B(n9196), .A(n9195), .Z(n9197) );
  XNOR U6199 ( .A(n9198), .B(n9197), .Z(out[906]) );
  ANDN U6200 ( .B(n9200), .A(n9199), .Z(n9201) );
  XNOR U6201 ( .A(n9202), .B(n9201), .Z(out[907]) );
  ANDN U6202 ( .B(n9204), .A(n9203), .Z(n9205) );
  XNOR U6203 ( .A(n9206), .B(n9205), .Z(out[908]) );
  ANDN U6204 ( .B(n9208), .A(n9207), .Z(n9209) );
  XNOR U6205 ( .A(n9210), .B(n9209), .Z(out[909]) );
  NOR U6206 ( .A(n9212), .B(n9211), .Z(n9213) );
  XNOR U6207 ( .A(n9214), .B(n9213), .Z(out[90]) );
  ANDN U6208 ( .B(n9216), .A(n9215), .Z(n9217) );
  XNOR U6209 ( .A(n9218), .B(n9217), .Z(out[910]) );
  ANDN U6210 ( .B(n9220), .A(n9219), .Z(n9221) );
  XNOR U6211 ( .A(n9222), .B(n9221), .Z(out[911]) );
  ANDN U6212 ( .B(n9224), .A(n9223), .Z(n9225) );
  XNOR U6213 ( .A(n9226), .B(n9225), .Z(out[912]) );
  ANDN U6214 ( .B(n9228), .A(n9227), .Z(n9229) );
  XNOR U6215 ( .A(n9230), .B(n9229), .Z(out[913]) );
  ANDN U6216 ( .B(n9232), .A(n9231), .Z(n9233) );
  XNOR U6217 ( .A(n9234), .B(n9233), .Z(out[914]) );
  ANDN U6218 ( .B(n9236), .A(n9235), .Z(n9237) );
  XNOR U6219 ( .A(n9238), .B(n9237), .Z(out[915]) );
  ANDN U6220 ( .B(n9240), .A(n9239), .Z(n9241) );
  XNOR U6221 ( .A(n9242), .B(n9241), .Z(out[916]) );
  ANDN U6222 ( .B(n9244), .A(n9243), .Z(n9245) );
  XNOR U6223 ( .A(n9246), .B(n9245), .Z(out[917]) );
  ANDN U6224 ( .B(n9248), .A(n9247), .Z(n9249) );
  XNOR U6225 ( .A(n9250), .B(n9249), .Z(out[918]) );
  ANDN U6226 ( .B(n9252), .A(n9251), .Z(n9253) );
  XNOR U6227 ( .A(n9254), .B(n9253), .Z(out[919]) );
  NOR U6228 ( .A(n9256), .B(n9255), .Z(n9257) );
  XNOR U6229 ( .A(n9258), .B(n9257), .Z(out[91]) );
  ANDN U6230 ( .B(n9260), .A(n9259), .Z(n9261) );
  XNOR U6231 ( .A(n9262), .B(n9261), .Z(out[920]) );
  ANDN U6232 ( .B(n9264), .A(n9263), .Z(n9265) );
  XNOR U6233 ( .A(n9266), .B(n9265), .Z(out[921]) );
  ANDN U6234 ( .B(n9268), .A(n9267), .Z(n9269) );
  XNOR U6235 ( .A(n9270), .B(n9269), .Z(out[922]) );
  ANDN U6236 ( .B(n9272), .A(n9271), .Z(n9273) );
  XNOR U6237 ( .A(n9274), .B(n9273), .Z(out[923]) );
  ANDN U6238 ( .B(n9276), .A(n9275), .Z(n9277) );
  XNOR U6239 ( .A(n9278), .B(n9277), .Z(out[924]) );
  ANDN U6240 ( .B(n9280), .A(n9279), .Z(n9281) );
  XNOR U6241 ( .A(n9282), .B(n9281), .Z(out[925]) );
  ANDN U6242 ( .B(n9284), .A(n9283), .Z(n9285) );
  XNOR U6243 ( .A(n9286), .B(n9285), .Z(out[926]) );
  ANDN U6244 ( .B(n9288), .A(n9287), .Z(n9289) );
  XNOR U6245 ( .A(n9290), .B(n9289), .Z(out[927]) );
  ANDN U6246 ( .B(n9292), .A(n9291), .Z(n9293) );
  XNOR U6247 ( .A(n9294), .B(n9293), .Z(out[928]) );
  ANDN U6248 ( .B(n9296), .A(n9295), .Z(n9297) );
  XNOR U6249 ( .A(n9298), .B(n9297), .Z(out[929]) );
  ANDN U6250 ( .B(n9300), .A(n9299), .Z(n9301) );
  XNOR U6251 ( .A(n9302), .B(n9301), .Z(out[92]) );
  ANDN U6252 ( .B(n9304), .A(n9303), .Z(n9305) );
  XNOR U6253 ( .A(n9306), .B(n9305), .Z(out[930]) );
  ANDN U6254 ( .B(n9308), .A(n9307), .Z(n9309) );
  XNOR U6255 ( .A(n9310), .B(n9309), .Z(out[931]) );
  ANDN U6256 ( .B(n9312), .A(n9311), .Z(n9313) );
  XNOR U6257 ( .A(n9314), .B(n9313), .Z(out[932]) );
  ANDN U6258 ( .B(n9316), .A(n9315), .Z(n9317) );
  XNOR U6259 ( .A(n9318), .B(n9317), .Z(out[933]) );
  ANDN U6260 ( .B(n9320), .A(n9319), .Z(n9321) );
  XNOR U6261 ( .A(n9322), .B(n9321), .Z(out[934]) );
  ANDN U6262 ( .B(n9324), .A(n9323), .Z(n9325) );
  XNOR U6263 ( .A(n9326), .B(n9325), .Z(out[935]) );
  ANDN U6264 ( .B(n9328), .A(n9327), .Z(n9329) );
  XNOR U6265 ( .A(n9330), .B(n9329), .Z(out[936]) );
  ANDN U6266 ( .B(n9332), .A(n9331), .Z(n9333) );
  XNOR U6267 ( .A(n9334), .B(n9333), .Z(out[937]) );
  ANDN U6268 ( .B(n9336), .A(n9335), .Z(n9337) );
  XNOR U6269 ( .A(n9338), .B(n9337), .Z(out[938]) );
  ANDN U6270 ( .B(n9340), .A(n9339), .Z(n9341) );
  XNOR U6271 ( .A(n9342), .B(n9341), .Z(out[939]) );
  ANDN U6272 ( .B(n9344), .A(n9343), .Z(n9345) );
  XNOR U6273 ( .A(n9346), .B(n9345), .Z(out[93]) );
  ANDN U6274 ( .B(n9348), .A(n9347), .Z(n9349) );
  XNOR U6275 ( .A(n9350), .B(n9349), .Z(out[940]) );
  ANDN U6276 ( .B(n9352), .A(n9351), .Z(n9353) );
  XNOR U6277 ( .A(n9354), .B(n9353), .Z(out[941]) );
  ANDN U6278 ( .B(n9356), .A(n9355), .Z(n9357) );
  XNOR U6279 ( .A(n9358), .B(n9357), .Z(out[942]) );
  ANDN U6280 ( .B(n9360), .A(n9359), .Z(n9361) );
  XNOR U6281 ( .A(n9362), .B(n9361), .Z(out[943]) );
  ANDN U6282 ( .B(n9364), .A(n9363), .Z(n9365) );
  XNOR U6283 ( .A(n9366), .B(n9365), .Z(out[944]) );
  ANDN U6284 ( .B(n9368), .A(n9367), .Z(n9369) );
  XNOR U6285 ( .A(n9370), .B(n9369), .Z(out[945]) );
  ANDN U6286 ( .B(n9372), .A(n9371), .Z(n9373) );
  XNOR U6287 ( .A(n9374), .B(n9373), .Z(out[946]) );
  ANDN U6288 ( .B(n9376), .A(n9375), .Z(n9377) );
  XNOR U6289 ( .A(n9378), .B(n9377), .Z(out[947]) );
  ANDN U6290 ( .B(n9380), .A(n9379), .Z(n9381) );
  XNOR U6291 ( .A(n9382), .B(n9381), .Z(out[948]) );
  ANDN U6292 ( .B(n9384), .A(n9383), .Z(n9385) );
  XNOR U6293 ( .A(n9386), .B(n9385), .Z(out[949]) );
  ANDN U6294 ( .B(n9388), .A(n9387), .Z(n9389) );
  XNOR U6295 ( .A(n9390), .B(n9389), .Z(out[94]) );
  ANDN U6296 ( .B(n9392), .A(n9391), .Z(n9393) );
  XNOR U6297 ( .A(n9394), .B(n9393), .Z(out[950]) );
  ANDN U6298 ( .B(n9396), .A(n9395), .Z(n9397) );
  XNOR U6299 ( .A(n9398), .B(n9397), .Z(out[951]) );
  ANDN U6300 ( .B(n9400), .A(n9399), .Z(n9401) );
  XNOR U6301 ( .A(n9402), .B(n9401), .Z(out[952]) );
  ANDN U6302 ( .B(n9404), .A(n9403), .Z(n9405) );
  XNOR U6303 ( .A(n9406), .B(n9405), .Z(out[953]) );
  ANDN U6304 ( .B(n9408), .A(n9407), .Z(n9409) );
  XNOR U6305 ( .A(n9410), .B(n9409), .Z(out[954]) );
  ANDN U6306 ( .B(n9412), .A(n9411), .Z(n9413) );
  XNOR U6307 ( .A(n9414), .B(n9413), .Z(out[955]) );
  ANDN U6308 ( .B(n9416), .A(n9415), .Z(n9417) );
  XNOR U6309 ( .A(n9418), .B(n9417), .Z(out[956]) );
  ANDN U6310 ( .B(n9420), .A(n9419), .Z(n9421) );
  XNOR U6311 ( .A(n9422), .B(n9421), .Z(out[957]) );
  ANDN U6312 ( .B(n9424), .A(n9423), .Z(n9425) );
  XNOR U6313 ( .A(n9426), .B(n9425), .Z(out[958]) );
  ANDN U6314 ( .B(n9428), .A(n9427), .Z(n9429) );
  XNOR U6315 ( .A(n9430), .B(n9429), .Z(out[959]) );
  ANDN U6316 ( .B(n9432), .A(n9431), .Z(n9433) );
  XNOR U6317 ( .A(n9434), .B(n9433), .Z(out[95]) );
  ANDN U6318 ( .B(n9436), .A(n9435), .Z(n9437) );
  XNOR U6319 ( .A(n9438), .B(n9437), .Z(out[960]) );
  ANDN U6320 ( .B(n9440), .A(n9439), .Z(n9441) );
  XNOR U6321 ( .A(n9442), .B(n9441), .Z(out[961]) );
  ANDN U6322 ( .B(n9444), .A(n9443), .Z(n9445) );
  XNOR U6323 ( .A(n9446), .B(n9445), .Z(out[962]) );
  ANDN U6324 ( .B(n9448), .A(n9447), .Z(n9449) );
  XNOR U6325 ( .A(n9450), .B(n9449), .Z(out[963]) );
  ANDN U6326 ( .B(n9452), .A(n9451), .Z(n9453) );
  XNOR U6327 ( .A(n9454), .B(n9453), .Z(out[964]) );
  ANDN U6328 ( .B(n9456), .A(n9455), .Z(n9457) );
  XNOR U6329 ( .A(n9458), .B(n9457), .Z(out[965]) );
  ANDN U6330 ( .B(n9460), .A(n9459), .Z(n9461) );
  XNOR U6331 ( .A(n9462), .B(n9461), .Z(out[966]) );
  ANDN U6332 ( .B(n9464), .A(n9463), .Z(n9465) );
  XNOR U6333 ( .A(n9466), .B(n9465), .Z(out[967]) );
  ANDN U6334 ( .B(n9468), .A(n9467), .Z(n9469) );
  XNOR U6335 ( .A(n9470), .B(n9469), .Z(out[968]) );
  ANDN U6336 ( .B(n9472), .A(n9471), .Z(n9473) );
  XNOR U6337 ( .A(n9474), .B(n9473), .Z(out[969]) );
  ANDN U6338 ( .B(n9476), .A(n9475), .Z(n9477) );
  XNOR U6339 ( .A(n9478), .B(n9477), .Z(out[96]) );
  ANDN U6340 ( .B(n9480), .A(n9479), .Z(n9481) );
  XNOR U6341 ( .A(n9482), .B(n9481), .Z(out[970]) );
  ANDN U6342 ( .B(n9484), .A(n9483), .Z(n9485) );
  XNOR U6343 ( .A(n9486), .B(n9485), .Z(out[971]) );
  ANDN U6344 ( .B(n9488), .A(n9487), .Z(n9489) );
  XNOR U6345 ( .A(n9490), .B(n9489), .Z(out[972]) );
  ANDN U6346 ( .B(n9492), .A(n9491), .Z(n9493) );
  XNOR U6347 ( .A(n9494), .B(n9493), .Z(out[973]) );
  ANDN U6348 ( .B(n9496), .A(n9495), .Z(n9497) );
  XNOR U6349 ( .A(n9498), .B(n9497), .Z(out[974]) );
  ANDN U6350 ( .B(n9500), .A(n9499), .Z(n9501) );
  XNOR U6351 ( .A(n9502), .B(n9501), .Z(out[975]) );
  ANDN U6352 ( .B(n9504), .A(n9503), .Z(n9505) );
  XNOR U6353 ( .A(n9506), .B(n9505), .Z(out[976]) );
  ANDN U6354 ( .B(n9508), .A(n9507), .Z(n9509) );
  XNOR U6355 ( .A(n9510), .B(n9509), .Z(out[977]) );
  ANDN U6356 ( .B(n9512), .A(n9511), .Z(n9513) );
  XNOR U6357 ( .A(n9514), .B(n9513), .Z(out[978]) );
  ANDN U6358 ( .B(n9516), .A(n9515), .Z(n9517) );
  XNOR U6359 ( .A(n9518), .B(n9517), .Z(out[979]) );
  ANDN U6360 ( .B(n9520), .A(n9519), .Z(n9521) );
  XNOR U6361 ( .A(n9522), .B(n9521), .Z(out[97]) );
  ANDN U6362 ( .B(n9524), .A(n9523), .Z(n9525) );
  XNOR U6363 ( .A(n9526), .B(n9525), .Z(out[980]) );
  ANDN U6364 ( .B(n9528), .A(n9527), .Z(n9529) );
  XNOR U6365 ( .A(n9530), .B(n9529), .Z(out[981]) );
  ANDN U6366 ( .B(n9532), .A(n9531), .Z(n9533) );
  XNOR U6367 ( .A(n9534), .B(n9533), .Z(out[982]) );
  ANDN U6368 ( .B(n9536), .A(n9535), .Z(n9537) );
  XNOR U6369 ( .A(n9538), .B(n9537), .Z(out[983]) );
  ANDN U6370 ( .B(n9540), .A(n9539), .Z(n9541) );
  XNOR U6371 ( .A(n9542), .B(n9541), .Z(out[984]) );
  ANDN U6372 ( .B(n9544), .A(n9543), .Z(n9545) );
  XNOR U6373 ( .A(n9546), .B(n9545), .Z(out[985]) );
  ANDN U6374 ( .B(n9548), .A(n9547), .Z(n9549) );
  XNOR U6375 ( .A(n9550), .B(n9549), .Z(out[986]) );
  ANDN U6376 ( .B(n9552), .A(n9551), .Z(n9553) );
  XNOR U6377 ( .A(n9554), .B(n9553), .Z(out[987]) );
  ANDN U6378 ( .B(n9556), .A(n9555), .Z(n9557) );
  XNOR U6379 ( .A(n9558), .B(n9557), .Z(out[988]) );
  ANDN U6380 ( .B(n9560), .A(n9559), .Z(n9561) );
  XNOR U6381 ( .A(n9562), .B(n9561), .Z(out[989]) );
  ANDN U6382 ( .B(n9564), .A(n9563), .Z(n9565) );
  XNOR U6383 ( .A(n9566), .B(n9565), .Z(out[98]) );
  ANDN U6384 ( .B(n9568), .A(n9567), .Z(n9569) );
  XNOR U6385 ( .A(n9570), .B(n9569), .Z(out[990]) );
  ANDN U6386 ( .B(n9572), .A(n9571), .Z(n9573) );
  XNOR U6387 ( .A(n9574), .B(n9573), .Z(out[991]) );
  ANDN U6388 ( .B(n9576), .A(n9575), .Z(n9577) );
  XNOR U6389 ( .A(n9578), .B(n9577), .Z(out[992]) );
  ANDN U6390 ( .B(n9580), .A(n9579), .Z(n9581) );
  XNOR U6391 ( .A(n9582), .B(n9581), .Z(out[993]) );
  ANDN U6392 ( .B(n9584), .A(n9583), .Z(n9585) );
  XNOR U6393 ( .A(n9586), .B(n9585), .Z(out[994]) );
  ANDN U6394 ( .B(n9588), .A(n9587), .Z(n9589) );
  XNOR U6395 ( .A(n9590), .B(n9589), .Z(out[995]) );
  ANDN U6396 ( .B(n9592), .A(n9591), .Z(n9593) );
  XNOR U6397 ( .A(n9594), .B(n9593), .Z(out[996]) );
  ANDN U6398 ( .B(n9596), .A(n9595), .Z(n9597) );
  XNOR U6399 ( .A(n9598), .B(n9597), .Z(out[997]) );
  ANDN U6400 ( .B(n9600), .A(n9599), .Z(n9601) );
  XNOR U6401 ( .A(n9602), .B(n9601), .Z(out[998]) );
  ANDN U6402 ( .B(n9604), .A(n9603), .Z(n9605) );
  XNOR U6403 ( .A(n9606), .B(n9605), .Z(out[999]) );
  ANDN U6404 ( .B(n9608), .A(n9607), .Z(n9609) );
  XNOR U6405 ( .A(n9610), .B(n9609), .Z(out[99]) );
  OR U6406 ( .A(n9612), .B(n9611), .Z(n9613) );
  XNOR U6407 ( .A(n9614), .B(n9613), .Z(out[9]) );
endmodule


module round_1 ( in, round_const, out );
  input [1599:0] in;
  input [63:0] round_const;
  output [1599:0] out;
  wire   round_const_63, round_const_31, round_const_15, round_const_7,
         round_const_3, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614;
  assign round_const_63 = round_const[63];
  assign round_const_31 = round_const[31];
  assign round_const_15 = round_const[15];
  assign round_const_7 = round_const[7];
  assign round_const_3 = round_const[3];

  XOR U1 ( .A(in[1469]), .B(in[509]), .Z(n4809) );
  XNOR U2 ( .A(in[829]), .B(in[189]), .Z(n4808) );
  XNOR U3 ( .A(n4809), .B(n4808), .Z(n4810) );
  XOR U4 ( .A(in[1149]), .B(n4810), .Z(n5679) );
  XOR U5 ( .A(in[1598]), .B(in[638]), .Z(n4812) );
  XNOR U6 ( .A(in[958]), .B(in[318]), .Z(n4811) );
  XNOR U7 ( .A(n4812), .B(n4811), .Z(n4813) );
  XOR U8 ( .A(in[1278]), .B(n4813), .Z(n6280) );
  XNOR U9 ( .A(n5679), .B(n6280), .Z(n8622) );
  XNOR U10 ( .A(in[254]), .B(n8622), .Z(n8384) );
  XOR U11 ( .A(in[1345]), .B(in[65]), .Z(n4815) );
  XNOR U12 ( .A(in[1025]), .B(in[385]), .Z(n4814) );
  XNOR U13 ( .A(n4815), .B(n4814), .Z(n4816) );
  XOR U14 ( .A(in[705]), .B(n4816), .Z(n6288) );
  XOR U15 ( .A(in[1474]), .B(in[514]), .Z(n4818) );
  XNOR U16 ( .A(in[834]), .B(in[194]), .Z(n4817) );
  XNOR U17 ( .A(n4818), .B(n4817), .Z(n4819) );
  XNOR U18 ( .A(in[1154]), .B(n4819), .Z(n5995) );
  XNOR U19 ( .A(n6288), .B(n5995), .Z(n8377) );
  XNOR U20 ( .A(in[1410]), .B(n8377), .Z(n8383) );
  XOR U21 ( .A(in[137]), .B(in[457]), .Z(n4821) );
  XNOR U22 ( .A(in[777]), .B(in[1417]), .Z(n4820) );
  XNOR U23 ( .A(n4821), .B(n4820), .Z(n4822) );
  XOR U24 ( .A(in[1097]), .B(n4822), .Z(n5948) );
  XOR U25 ( .A(in[328]), .B(in[8]), .Z(n4824) );
  XNOR U26 ( .A(in[968]), .B(in[648]), .Z(n4823) );
  XNOR U27 ( .A(n4824), .B(n4823), .Z(n4825) );
  XOR U28 ( .A(in[1288]), .B(n4825), .Z(n6016) );
  XNOR U29 ( .A(n5948), .B(n6016), .Z(n8893) );
  XNOR U30 ( .A(in[1033]), .B(n8893), .Z(n7416) );
  NAND U31 ( .A(n8383), .B(n7416), .Z(n4826) );
  XNOR U32 ( .A(n8384), .B(n4826), .Z(out[0]) );
  XOR U33 ( .A(in[1386]), .B(in[106]), .Z(n4828) );
  XNOR U34 ( .A(in[1066]), .B(in[746]), .Z(n4827) );
  XNOR U35 ( .A(n4828), .B(n4827), .Z(n4829) );
  XOR U36 ( .A(in[426]), .B(n4829), .Z(n5282) );
  XOR U37 ( .A(in[1515]), .B(in[555]), .Z(n4831) );
  XNOR U38 ( .A(in[875]), .B(in[235]), .Z(n4830) );
  XNOR U39 ( .A(n4831), .B(n4830), .Z(n4832) );
  XOR U40 ( .A(in[1195]), .B(n4832), .Z(n6136) );
  XNOR U41 ( .A(n5282), .B(n6136), .Z(n8557) );
  XNOR U42 ( .A(in[171]), .B(n8557), .Z(n6108) );
  XOR U43 ( .A(in[971]), .B(in[1291]), .Z(n4834) );
  XNOR U44 ( .A(in[11]), .B(in[331]), .Z(n4833) );
  XNOR U45 ( .A(n4834), .B(n4833), .Z(n4835) );
  XOR U46 ( .A(in[651]), .B(n4835), .Z(n6027) );
  XOR U47 ( .A(in[140]), .B(in[460]), .Z(n4837) );
  XNOR U48 ( .A(in[1100]), .B(in[1420]), .Z(n4836) );
  XNOR U49 ( .A(n4837), .B(n4836), .Z(n4838) );
  XNOR U50 ( .A(in[780]), .B(n4838), .Z(n5966) );
  XNOR U51 ( .A(n6027), .B(n5966), .Z(n8902) );
  XNOR U52 ( .A(in[1356]), .B(n8902), .Z(n6503) );
  XOR U53 ( .A(in[1364]), .B(in[724]), .Z(n4840) );
  XNOR U54 ( .A(in[84]), .B(in[404]), .Z(n4839) );
  XNOR U55 ( .A(n4840), .B(n4839), .Z(n4841) );
  XOR U56 ( .A(in[1044]), .B(n4841), .Z(n5584) );
  XOR U57 ( .A(in[1555]), .B(in[595]), .Z(n4843) );
  XNOR U58 ( .A(in[915]), .B(in[275]), .Z(n4842) );
  XNOR U59 ( .A(n4843), .B(n4842), .Z(n4844) );
  XOR U60 ( .A(in[1235]), .B(n4844), .Z(n5296) );
  XNOR U61 ( .A(n5584), .B(n5296), .Z(n8689) );
  XNOR U62 ( .A(in[980]), .B(n8689), .Z(n6500) );
  NAND U63 ( .A(n6503), .B(n6500), .Z(n4845) );
  XNOR U64 ( .A(n6108), .B(n4845), .Z(out[1000]) );
  XOR U65 ( .A(in[1387]), .B(in[107]), .Z(n4847) );
  XNOR U66 ( .A(in[1067]), .B(in[747]), .Z(n4846) );
  XNOR U67 ( .A(n4847), .B(n4846), .Z(n4848) );
  XOR U68 ( .A(in[427]), .B(n4848), .Z(n5293) );
  XOR U69 ( .A(in[1516]), .B(in[556]), .Z(n4850) );
  XNOR U70 ( .A(in[876]), .B(in[236]), .Z(n4849) );
  XNOR U71 ( .A(n4850), .B(n4849), .Z(n4851) );
  XOR U72 ( .A(in[1196]), .B(n4851), .Z(n6140) );
  XNOR U73 ( .A(n5293), .B(n6140), .Z(n8565) );
  XNOR U74 ( .A(in[172]), .B(n8565), .Z(n6112) );
  XOR U75 ( .A(in[972]), .B(in[12]), .Z(n4853) );
  XNOR U76 ( .A(in[1292]), .B(in[332]), .Z(n4852) );
  XNOR U77 ( .A(n4853), .B(n4852), .Z(n4854) );
  XOR U78 ( .A(in[652]), .B(n4854), .Z(n6030) );
  XOR U79 ( .A(in[141]), .B(in[461]), .Z(n4856) );
  XNOR U80 ( .A(in[1101]), .B(in[1421]), .Z(n4855) );
  XNOR U81 ( .A(n4856), .B(n4855), .Z(n4857) );
  XNOR U82 ( .A(in[781]), .B(n4857), .Z(n5971) );
  XNOR U83 ( .A(n6030), .B(n5971), .Z(n8905) );
  XNOR U84 ( .A(in[1357]), .B(n8905), .Z(n6507) );
  XOR U85 ( .A(in[1365]), .B(in[725]), .Z(n4859) );
  XNOR U86 ( .A(in[85]), .B(in[405]), .Z(n4858) );
  XNOR U87 ( .A(n4859), .B(n4858), .Z(n4860) );
  XOR U88 ( .A(in[1045]), .B(n4860), .Z(n5597) );
  XOR U89 ( .A(in[1556]), .B(in[596]), .Z(n4862) );
  XNOR U90 ( .A(in[916]), .B(in[276]), .Z(n4861) );
  XNOR U91 ( .A(n4862), .B(n4861), .Z(n4863) );
  XOR U92 ( .A(in[1236]), .B(n4863), .Z(n5311) );
  XNOR U93 ( .A(n5597), .B(n5311), .Z(n8691) );
  XNOR U94 ( .A(in[981]), .B(n8691), .Z(n6504) );
  NAND U95 ( .A(n6507), .B(n6504), .Z(n4864) );
  XNOR U96 ( .A(n6112), .B(n4864), .Z(out[1001]) );
  XOR U97 ( .A(in[1388]), .B(in[108]), .Z(n4866) );
  XNOR U98 ( .A(in[1068]), .B(in[748]), .Z(n4865) );
  XNOR U99 ( .A(n4866), .B(n4865), .Z(n4867) );
  XOR U100 ( .A(in[428]), .B(n4867), .Z(n6202) );
  XOR U101 ( .A(in[1517]), .B(in[557]), .Z(n4869) );
  XNOR U102 ( .A(in[877]), .B(in[237]), .Z(n4868) );
  XNOR U103 ( .A(n4869), .B(n4868), .Z(n4870) );
  XOR U104 ( .A(in[1197]), .B(n4870), .Z(n6144) );
  XNOR U105 ( .A(n6202), .B(n6144), .Z(n8569) );
  XNOR U106 ( .A(in[173]), .B(n8569), .Z(n6117) );
  XOR U107 ( .A(in[973]), .B(in[13]), .Z(n4872) );
  XNOR U108 ( .A(in[1293]), .B(in[333]), .Z(n4871) );
  XNOR U109 ( .A(n4872), .B(n4871), .Z(n4873) );
  XOR U110 ( .A(in[653]), .B(n4873), .Z(n6033) );
  XOR U111 ( .A(in[142]), .B(in[1422]), .Z(n4875) );
  XNOR U112 ( .A(in[1102]), .B(in[782]), .Z(n4874) );
  XNOR U113 ( .A(n4875), .B(n4874), .Z(n4876) );
  XNOR U114 ( .A(in[462]), .B(n4876), .Z(n5976) );
  XNOR U115 ( .A(n6033), .B(n5976), .Z(n8908) );
  XNOR U116 ( .A(in[1358]), .B(n8908), .Z(n6511) );
  XOR U117 ( .A(in[1366]), .B(in[726]), .Z(n4878) );
  XNOR U118 ( .A(in[86]), .B(in[406]), .Z(n4877) );
  XNOR U119 ( .A(n4878), .B(n4877), .Z(n4879) );
  XOR U120 ( .A(in[1046]), .B(n4879), .Z(n5610) );
  XOR U121 ( .A(in[1557]), .B(in[597]), .Z(n4881) );
  XNOR U122 ( .A(in[917]), .B(in[277]), .Z(n4880) );
  XNOR U123 ( .A(n4881), .B(n4880), .Z(n4882) );
  XOR U124 ( .A(in[1237]), .B(n4882), .Z(n5326) );
  XNOR U125 ( .A(n5610), .B(n5326), .Z(n8693) );
  XNOR U126 ( .A(in[982]), .B(n8693), .Z(n6508) );
  NAND U127 ( .A(n6511), .B(n6508), .Z(n4883) );
  XNOR U128 ( .A(n6117), .B(n4883), .Z(out[1002]) );
  XOR U129 ( .A(in[1389]), .B(in[109]), .Z(n4885) );
  XNOR U130 ( .A(in[1069]), .B(in[749]), .Z(n4884) );
  XNOR U131 ( .A(n4885), .B(n4884), .Z(n4886) );
  XOR U132 ( .A(in[429]), .B(n4886), .Z(n6206) );
  XOR U133 ( .A(in[1518]), .B(in[558]), .Z(n4888) );
  XNOR U134 ( .A(in[878]), .B(in[238]), .Z(n4887) );
  XNOR U135 ( .A(n4888), .B(n4887), .Z(n4889) );
  XOR U136 ( .A(in[1198]), .B(n4889), .Z(n6148) );
  XNOR U137 ( .A(n6206), .B(n6148), .Z(n8573) );
  XNOR U138 ( .A(in[174]), .B(n8573), .Z(n6121) );
  XOR U139 ( .A(in[143]), .B(in[1423]), .Z(n4891) );
  XNOR U140 ( .A(in[1103]), .B(in[783]), .Z(n4890) );
  XNOR U141 ( .A(n4891), .B(n4890), .Z(n4892) );
  XOR U142 ( .A(in[463]), .B(n4892), .Z(n5981) );
  XOR U143 ( .A(in[974]), .B(in[14]), .Z(n4894) );
  XNOR U144 ( .A(in[1294]), .B(in[334]), .Z(n4893) );
  XNOR U145 ( .A(n4894), .B(n4893), .Z(n4895) );
  XNOR U146 ( .A(in[654]), .B(n4895), .Z(n6036) );
  XNOR U147 ( .A(n5981), .B(n6036), .Z(n8911) );
  XNOR U148 ( .A(in[1359]), .B(n8911), .Z(n6515) );
  XOR U149 ( .A(in[1367]), .B(in[727]), .Z(n4897) );
  XNOR U150 ( .A(in[87]), .B(in[407]), .Z(n4896) );
  XNOR U151 ( .A(n4897), .B(n4896), .Z(n4898) );
  XOR U152 ( .A(in[1047]), .B(n4898), .Z(n5623) );
  XOR U153 ( .A(in[1558]), .B(in[598]), .Z(n4900) );
  XNOR U154 ( .A(in[918]), .B(in[278]), .Z(n4899) );
  XNOR U155 ( .A(n4900), .B(n4899), .Z(n4901) );
  XOR U156 ( .A(in[1238]), .B(n4901), .Z(n5341) );
  XNOR U157 ( .A(n5623), .B(n5341), .Z(n8695) );
  XNOR U158 ( .A(in[983]), .B(n8695), .Z(n6512) );
  NAND U159 ( .A(n6515), .B(n6512), .Z(n4902) );
  XNOR U160 ( .A(n6121), .B(n4902), .Z(out[1003]) );
  XOR U161 ( .A(in[1390]), .B(in[110]), .Z(n4904) );
  XNOR U162 ( .A(in[1070]), .B(in[750]), .Z(n4903) );
  XNOR U163 ( .A(n4904), .B(n4903), .Z(n4905) );
  XOR U164 ( .A(in[430]), .B(n4905), .Z(n6210) );
  XOR U165 ( .A(in[1519]), .B(in[559]), .Z(n4907) );
  XNOR U166 ( .A(in[879]), .B(in[239]), .Z(n4906) );
  XNOR U167 ( .A(n4907), .B(n4906), .Z(n4908) );
  XOR U168 ( .A(in[1199]), .B(n4908), .Z(n6152) );
  XNOR U169 ( .A(n6210), .B(n6152), .Z(n8577) );
  XNOR U170 ( .A(in[175]), .B(n8577), .Z(n6125) );
  XOR U171 ( .A(in[144]), .B(in[1424]), .Z(n4910) );
  XNOR U172 ( .A(in[1104]), .B(in[784]), .Z(n4909) );
  XNOR U173 ( .A(n4910), .B(n4909), .Z(n4911) );
  XOR U174 ( .A(in[464]), .B(n4911), .Z(n5986) );
  XOR U175 ( .A(in[975]), .B(in[15]), .Z(n4913) );
  XNOR U176 ( .A(in[1295]), .B(in[335]), .Z(n4912) );
  XNOR U177 ( .A(n4913), .B(n4912), .Z(n4914) );
  XNOR U178 ( .A(in[655]), .B(n4914), .Z(n6039) );
  XNOR U179 ( .A(n5986), .B(n6039), .Z(n8914) );
  XNOR U180 ( .A(in[1360]), .B(n8914), .Z(n6520) );
  XOR U181 ( .A(in[1368]), .B(in[728]), .Z(n4916) );
  XNOR U182 ( .A(in[88]), .B(in[408]), .Z(n4915) );
  XNOR U183 ( .A(n4916), .B(n4915), .Z(n4917) );
  XOR U184 ( .A(in[1048]), .B(n4917), .Z(n5636) );
  XOR U185 ( .A(in[1559]), .B(in[599]), .Z(n4919) );
  XNOR U186 ( .A(in[919]), .B(in[279]), .Z(n4918) );
  XNOR U187 ( .A(n4919), .B(n4918), .Z(n4920) );
  XOR U188 ( .A(in[1239]), .B(n4920), .Z(n5356) );
  XNOR U189 ( .A(n5636), .B(n5356), .Z(n8697) );
  XNOR U190 ( .A(in[984]), .B(n8697), .Z(n6517) );
  NAND U191 ( .A(n6520), .B(n6517), .Z(n4921) );
  XNOR U192 ( .A(n6125), .B(n4921), .Z(out[1004]) );
  XOR U193 ( .A(in[1391]), .B(in[111]), .Z(n4923) );
  XNOR U194 ( .A(in[1071]), .B(in[751]), .Z(n4922) );
  XNOR U195 ( .A(n4923), .B(n4922), .Z(n4924) );
  XOR U196 ( .A(in[431]), .B(n4924), .Z(n6214) );
  XOR U197 ( .A(in[1520]), .B(in[560]), .Z(n4926) );
  XNOR U198 ( .A(in[880]), .B(in[240]), .Z(n4925) );
  XNOR U199 ( .A(n4926), .B(n4925), .Z(n4927) );
  XOR U200 ( .A(in[1200]), .B(n4927), .Z(n6157) );
  XNOR U201 ( .A(n6214), .B(n6157), .Z(n8581) );
  XNOR U202 ( .A(in[176]), .B(n8581), .Z(n6129) );
  XOR U203 ( .A(in[145]), .B(in[1425]), .Z(n4929) );
  XNOR U204 ( .A(in[1105]), .B(in[785]), .Z(n4928) );
  XNOR U205 ( .A(n4929), .B(n4928), .Z(n4930) );
  XOR U206 ( .A(in[465]), .B(n4930), .Z(n5991) );
  XOR U207 ( .A(in[976]), .B(in[16]), .Z(n4932) );
  XNOR U208 ( .A(in[1296]), .B(in[336]), .Z(n4931) );
  XNOR U209 ( .A(n4932), .B(n4931), .Z(n4933) );
  XNOR U210 ( .A(in[656]), .B(n4933), .Z(n6042) );
  XNOR U211 ( .A(n5991), .B(n6042), .Z(n8921) );
  XNOR U212 ( .A(in[1361]), .B(n8921), .Z(n6524) );
  XOR U213 ( .A(in[1369]), .B(in[729]), .Z(n4935) );
  XNOR U214 ( .A(in[89]), .B(in[409]), .Z(n4934) );
  XNOR U215 ( .A(n4935), .B(n4934), .Z(n4936) );
  XOR U216 ( .A(in[1049]), .B(n4936), .Z(n5649) );
  XOR U217 ( .A(in[1560]), .B(in[600]), .Z(n4938) );
  XNOR U218 ( .A(in[920]), .B(in[280]), .Z(n4937) );
  XNOR U219 ( .A(n4938), .B(n4937), .Z(n4939) );
  XOR U220 ( .A(in[1240]), .B(n4939), .Z(n5371) );
  XNOR U221 ( .A(n5649), .B(n5371), .Z(n8699) );
  XNOR U222 ( .A(in[985]), .B(n8699), .Z(n6521) );
  NAND U223 ( .A(n6524), .B(n6521), .Z(n4940) );
  XNOR U224 ( .A(n6129), .B(n4940), .Z(out[1005]) );
  XOR U225 ( .A(in[1392]), .B(in[112]), .Z(n4942) );
  XNOR U226 ( .A(in[1072]), .B(in[752]), .Z(n4941) );
  XNOR U227 ( .A(n4942), .B(n4941), .Z(n4943) );
  XOR U228 ( .A(in[432]), .B(n4943), .Z(n6218) );
  XOR U229 ( .A(in[1521]), .B(in[561]), .Z(n4945) );
  XNOR U230 ( .A(in[881]), .B(in[241]), .Z(n4944) );
  XNOR U231 ( .A(n4945), .B(n4944), .Z(n4946) );
  XOR U232 ( .A(in[1201]), .B(n4946), .Z(n6161) );
  XNOR U233 ( .A(n6218), .B(n6161), .Z(n8585) );
  XNOR U234 ( .A(in[177]), .B(n8585), .Z(n6133) );
  XOR U235 ( .A(in[17]), .B(in[657]), .Z(n4948) );
  XNOR U236 ( .A(in[977]), .B(in[337]), .Z(n4947) );
  XNOR U237 ( .A(n4948), .B(n4947), .Z(n4949) );
  XOR U238 ( .A(in[1297]), .B(n4949), .Z(n6045) );
  XOR U239 ( .A(in[1426]), .B(in[466]), .Z(n4951) );
  XNOR U240 ( .A(in[786]), .B(in[146]), .Z(n4950) );
  XNOR U241 ( .A(n4951), .B(n4950), .Z(n4952) );
  XNOR U242 ( .A(in[1106]), .B(n4952), .Z(n5295) );
  XNOR U243 ( .A(n6045), .B(n5295), .Z(n8924) );
  XNOR U244 ( .A(n8924), .B(in[1362]), .Z(n6528) );
  XOR U245 ( .A(in[1370]), .B(in[730]), .Z(n4954) );
  XNOR U246 ( .A(in[90]), .B(in[410]), .Z(n4953) );
  XNOR U247 ( .A(n4954), .B(n4953), .Z(n4955) );
  XOR U248 ( .A(in[1050]), .B(n4955), .Z(n5664) );
  XOR U249 ( .A(in[1561]), .B(in[601]), .Z(n4957) );
  XNOR U250 ( .A(in[921]), .B(in[281]), .Z(n4956) );
  XNOR U251 ( .A(n4957), .B(n4956), .Z(n4958) );
  XOR U252 ( .A(in[1241]), .B(n4958), .Z(n5397) );
  XNOR U253 ( .A(n5664), .B(n5397), .Z(n8701) );
  XNOR U254 ( .A(in[986]), .B(n8701), .Z(n6525) );
  NAND U255 ( .A(n6528), .B(n6525), .Z(n4959) );
  XNOR U256 ( .A(n6133), .B(n4959), .Z(out[1006]) );
  XOR U257 ( .A(in[1393]), .B(in[113]), .Z(n4961) );
  XNOR U258 ( .A(in[1073]), .B(in[753]), .Z(n4960) );
  XNOR U259 ( .A(n4961), .B(n4960), .Z(n4962) );
  XOR U260 ( .A(in[433]), .B(n4962), .Z(n6222) );
  XOR U261 ( .A(in[1522]), .B(in[562]), .Z(n4964) );
  XNOR U262 ( .A(in[882]), .B(in[242]), .Z(n4963) );
  XNOR U263 ( .A(n4964), .B(n4963), .Z(n4965) );
  XOR U264 ( .A(in[1202]), .B(n4965), .Z(n6165) );
  XNOR U265 ( .A(n6222), .B(n6165), .Z(n8589) );
  XNOR U266 ( .A(in[178]), .B(n8589), .Z(n6137) );
  XOR U267 ( .A(in[147]), .B(in[1427]), .Z(n4967) );
  XNOR U268 ( .A(in[1107]), .B(in[787]), .Z(n4966) );
  XNOR U269 ( .A(n4967), .B(n4966), .Z(n4968) );
  XOR U270 ( .A(in[467]), .B(n4968), .Z(n5310) );
  XOR U271 ( .A(in[978]), .B(in[18]), .Z(n4970) );
  XNOR U272 ( .A(in[1298]), .B(in[338]), .Z(n4969) );
  XNOR U273 ( .A(n4970), .B(n4969), .Z(n4971) );
  XNOR U274 ( .A(in[658]), .B(n4971), .Z(n6048) );
  XNOR U275 ( .A(n5310), .B(n6048), .Z(n8927) );
  XNOR U276 ( .A(in[1363]), .B(n8927), .Z(n6532) );
  XOR U277 ( .A(in[1371]), .B(in[731]), .Z(n4973) );
  XNOR U278 ( .A(in[91]), .B(in[411]), .Z(n4972) );
  XNOR U279 ( .A(n4973), .B(n4972), .Z(n4974) );
  XOR U280 ( .A(in[1051]), .B(n4974), .Z(n5677) );
  XOR U281 ( .A(in[1562]), .B(in[602]), .Z(n4976) );
  XNOR U282 ( .A(in[922]), .B(in[282]), .Z(n4975) );
  XNOR U283 ( .A(n4976), .B(n4975), .Z(n4977) );
  XOR U284 ( .A(in[1242]), .B(n4977), .Z(n5412) );
  XNOR U285 ( .A(n5677), .B(n5412), .Z(n8703) );
  XNOR U286 ( .A(in[987]), .B(n8703), .Z(n6529) );
  NAND U287 ( .A(n6532), .B(n6529), .Z(n4978) );
  XNOR U288 ( .A(n6137), .B(n4978), .Z(out[1007]) );
  XOR U289 ( .A(in[1394]), .B(in[114]), .Z(n4980) );
  XNOR U290 ( .A(in[1074]), .B(in[754]), .Z(n4979) );
  XNOR U291 ( .A(n4980), .B(n4979), .Z(n4981) );
  XOR U292 ( .A(in[434]), .B(n4981), .Z(n6226) );
  XOR U293 ( .A(in[1523]), .B(in[563]), .Z(n4983) );
  XNOR U294 ( .A(in[883]), .B(in[243]), .Z(n4982) );
  XNOR U295 ( .A(n4983), .B(n4982), .Z(n4984) );
  XOR U296 ( .A(in[1203]), .B(n4984), .Z(n6169) );
  XNOR U297 ( .A(n6226), .B(n6169), .Z(n8593) );
  XNOR U298 ( .A(in[179]), .B(n8593), .Z(n6141) );
  XOR U299 ( .A(in[148]), .B(in[1428]), .Z(n4986) );
  XNOR U300 ( .A(in[1108]), .B(in[788]), .Z(n4985) );
  XNOR U301 ( .A(n4986), .B(n4985), .Z(n4987) );
  XOR U302 ( .A(in[468]), .B(n4987), .Z(n5325) );
  XOR U303 ( .A(in[979]), .B(in[19]), .Z(n4989) );
  XNOR U304 ( .A(in[1299]), .B(in[339]), .Z(n4988) );
  XNOR U305 ( .A(n4989), .B(n4988), .Z(n4990) );
  XNOR U306 ( .A(in[659]), .B(n4990), .Z(n6052) );
  XNOR U307 ( .A(n5325), .B(n6052), .Z(n8930) );
  XNOR U308 ( .A(in[1364]), .B(n8930), .Z(n6536) );
  XOR U309 ( .A(in[1372]), .B(in[732]), .Z(n4992) );
  XNOR U310 ( .A(in[92]), .B(in[412]), .Z(n4991) );
  XNOR U311 ( .A(n4992), .B(n4991), .Z(n4993) );
  XOR U312 ( .A(in[1052]), .B(n4993), .Z(n5697) );
  XOR U313 ( .A(in[1563]), .B(in[603]), .Z(n4995) );
  XNOR U314 ( .A(in[923]), .B(in[283]), .Z(n4994) );
  XNOR U315 ( .A(n4995), .B(n4994), .Z(n4996) );
  XOR U316 ( .A(in[1243]), .B(n4996), .Z(n5427) );
  XNOR U317 ( .A(n5697), .B(n5427), .Z(n8707) );
  XNOR U318 ( .A(in[988]), .B(n8707), .Z(n6533) );
  NAND U319 ( .A(n6536), .B(n6533), .Z(n4997) );
  XNOR U320 ( .A(n6141), .B(n4997), .Z(out[1008]) );
  XOR U321 ( .A(in[1395]), .B(in[115]), .Z(n4999) );
  XNOR U322 ( .A(in[1075]), .B(in[755]), .Z(n4998) );
  XNOR U323 ( .A(n4999), .B(n4998), .Z(n5000) );
  XOR U324 ( .A(in[435]), .B(n5000), .Z(n6230) );
  XOR U325 ( .A(in[1524]), .B(in[564]), .Z(n5002) );
  XNOR U326 ( .A(in[884]), .B(in[244]), .Z(n5001) );
  XNOR U327 ( .A(n5002), .B(n5001), .Z(n5003) );
  XOR U328 ( .A(in[1204]), .B(n5003), .Z(n6173) );
  XNOR U329 ( .A(n6230), .B(n6173), .Z(n8597) );
  XNOR U330 ( .A(in[180]), .B(n8597), .Z(n6145) );
  XOR U331 ( .A(in[340]), .B(in[660]), .Z(n5005) );
  XNOR U332 ( .A(in[20]), .B(in[1300]), .Z(n5004) );
  XNOR U333 ( .A(n5005), .B(n5004), .Z(n5006) );
  XOR U334 ( .A(in[980]), .B(n5006), .Z(n6055) );
  XOR U335 ( .A(in[149]), .B(in[1429]), .Z(n5008) );
  XNOR U336 ( .A(in[1109]), .B(in[789]), .Z(n5007) );
  XNOR U337 ( .A(n5008), .B(n5007), .Z(n5009) );
  XNOR U338 ( .A(in[469]), .B(n5009), .Z(n5340) );
  XNOR U339 ( .A(n6055), .B(n5340), .Z(n8933) );
  XNOR U340 ( .A(in[1365]), .B(n8933), .Z(n6540) );
  XOR U341 ( .A(in[1373]), .B(in[733]), .Z(n5011) );
  XNOR U342 ( .A(in[93]), .B(in[413]), .Z(n5010) );
  XNOR U343 ( .A(n5011), .B(n5010), .Z(n5012) );
  XOR U344 ( .A(in[1053]), .B(n5012), .Z(n5710) );
  XOR U345 ( .A(in[1564]), .B(in[604]), .Z(n5014) );
  XNOR U346 ( .A(in[924]), .B(in[284]), .Z(n5013) );
  XNOR U347 ( .A(n5014), .B(n5013), .Z(n5015) );
  XOR U348 ( .A(in[1244]), .B(n5015), .Z(n5442) );
  XNOR U349 ( .A(n5710), .B(n5442), .Z(n8709) );
  XNOR U350 ( .A(in[989]), .B(n8709), .Z(n6537) );
  NAND U351 ( .A(n6540), .B(n6537), .Z(n5016) );
  XNOR U352 ( .A(n6145), .B(n5016), .Z(out[1009]) );
  XOR U353 ( .A(in[1339]), .B(in[59]), .Z(n5018) );
  XNOR U354 ( .A(in[699]), .B(in[379]), .Z(n5017) );
  XNOR U355 ( .A(n5018), .B(n5017), .Z(n5019) );
  XOR U356 ( .A(in[1019]), .B(n5019), .Z(n5668) );
  XOR U357 ( .A(in[1530]), .B(in[570]), .Z(n5021) );
  XNOR U358 ( .A(in[1210]), .B(in[250]), .Z(n5020) );
  XNOR U359 ( .A(n5021), .B(n5020), .Z(n5022) );
  XOR U360 ( .A(in[890]), .B(n5022), .Z(n5134) );
  XNOR U361 ( .A(n5668), .B(n5134), .Z(n8399) );
  XNOR U362 ( .A(in[635]), .B(n8399), .Z(n7357) );
  XOR U363 ( .A(in[161]), .B(in[1441]), .Z(n5024) );
  XNOR U364 ( .A(in[801]), .B(in[1121]), .Z(n5023) );
  XNOR U365 ( .A(n5024), .B(n5023), .Z(n5025) );
  XOR U366 ( .A(in[481]), .B(n5025), .Z(n5261) );
  XOR U367 ( .A(in[1570]), .B(in[610]), .Z(n5027) );
  XNOR U368 ( .A(in[930]), .B(in[290]), .Z(n5026) );
  XNOR U369 ( .A(n5027), .B(n5026), .Z(n5028) );
  XNOR U370 ( .A(in[1250]), .B(n5028), .Z(n5144) );
  XNOR U371 ( .A(n5261), .B(n5144), .Z(n8496) );
  XNOR U372 ( .A(in[226]), .B(n8496), .Z(n7638) );
  XOR U373 ( .A(in[1510]), .B(in[550]), .Z(n5030) );
  XNOR U374 ( .A(in[870]), .B(in[230]), .Z(n5029) );
  XNOR U375 ( .A(n5030), .B(n5029), .Z(n5031) );
  XOR U376 ( .A(in[1190]), .B(n5031), .Z(n6116) );
  XOR U377 ( .A(in[1061]), .B(in[421]), .Z(n5033) );
  XNOR U378 ( .A(in[741]), .B(in[1381]), .Z(n5032) );
  XNOR U379 ( .A(n5033), .B(n5032), .Z(n5034) );
  XOR U380 ( .A(in[101]), .B(n5034), .Z(n5180) );
  XNOR U381 ( .A(n6116), .B(n5180), .Z(n8537) );
  XNOR U382 ( .A(in[1446]), .B(n8537), .Z(n7635) );
  NAND U383 ( .A(n7638), .B(n7635), .Z(n5035) );
  XNOR U384 ( .A(n7357), .B(n5035), .Z(out[100]) );
  XOR U385 ( .A(in[1396]), .B(in[116]), .Z(n5037) );
  XNOR U386 ( .A(in[1076]), .B(in[756]), .Z(n5036) );
  XNOR U387 ( .A(n5037), .B(n5036), .Z(n5038) );
  XOR U388 ( .A(in[436]), .B(n5038), .Z(n6235) );
  XOR U389 ( .A(in[1525]), .B(in[565]), .Z(n5040) );
  XNOR U390 ( .A(in[885]), .B(in[245]), .Z(n5039) );
  XNOR U391 ( .A(n5040), .B(n5039), .Z(n5041) );
  XOR U392 ( .A(in[1205]), .B(n5041), .Z(n6177) );
  XNOR U393 ( .A(n6235), .B(n6177), .Z(n8601) );
  XNOR U394 ( .A(in[181]), .B(n8601), .Z(n6149) );
  XOR U395 ( .A(in[341]), .B(in[661]), .Z(n5043) );
  XNOR U396 ( .A(in[21]), .B(in[1301]), .Z(n5042) );
  XNOR U397 ( .A(n5043), .B(n5042), .Z(n5044) );
  XOR U398 ( .A(in[981]), .B(n5044), .Z(n6058) );
  XOR U399 ( .A(in[150]), .B(in[1430]), .Z(n5046) );
  XNOR U400 ( .A(in[1110]), .B(in[790]), .Z(n5045) );
  XNOR U401 ( .A(n5046), .B(n5045), .Z(n5047) );
  XNOR U402 ( .A(in[470]), .B(n5047), .Z(n5355) );
  XNOR U403 ( .A(n6058), .B(n5355), .Z(n8936) );
  XNOR U404 ( .A(in[1366]), .B(n8936), .Z(n6544) );
  XOR U405 ( .A(in[1374]), .B(in[734]), .Z(n5049) );
  XNOR U406 ( .A(in[94]), .B(in[414]), .Z(n5048) );
  XNOR U407 ( .A(n5049), .B(n5048), .Z(n5050) );
  XOR U408 ( .A(in[1054]), .B(n5050), .Z(n5723) );
  XOR U409 ( .A(in[1565]), .B(in[605]), .Z(n5052) );
  XNOR U410 ( .A(in[925]), .B(in[285]), .Z(n5051) );
  XNOR U411 ( .A(n5052), .B(n5051), .Z(n5053) );
  XOR U412 ( .A(in[1245]), .B(n5053), .Z(n5457) );
  XNOR U413 ( .A(n5723), .B(n5457), .Z(n8711) );
  XNOR U414 ( .A(in[990]), .B(n8711), .Z(n6541) );
  NAND U415 ( .A(n6544), .B(n6541), .Z(n5054) );
  XNOR U416 ( .A(n6149), .B(n5054), .Z(out[1010]) );
  XOR U417 ( .A(in[1526]), .B(in[566]), .Z(n5056) );
  XNOR U418 ( .A(in[886]), .B(in[246]), .Z(n5055) );
  XNOR U419 ( .A(n5056), .B(n5055), .Z(n5057) );
  XOR U420 ( .A(in[1206]), .B(n5057), .Z(n6181) );
  XOR U421 ( .A(in[1397]), .B(in[117]), .Z(n5059) );
  XNOR U422 ( .A(in[1077]), .B(in[757]), .Z(n5058) );
  XNOR U423 ( .A(n5059), .B(n5058), .Z(n5060) );
  XOR U424 ( .A(in[437]), .B(n5060), .Z(n6239) );
  XNOR U425 ( .A(n6181), .B(n6239), .Z(n8611) );
  XNOR U426 ( .A(in[182]), .B(n8611), .Z(n6153) );
  XOR U427 ( .A(in[151]), .B(in[1431]), .Z(n5062) );
  XNOR U428 ( .A(in[1111]), .B(in[791]), .Z(n5061) );
  XNOR U429 ( .A(n5062), .B(n5061), .Z(n5063) );
  XOR U430 ( .A(in[471]), .B(n5063), .Z(n5370) );
  XOR U431 ( .A(in[342]), .B(in[662]), .Z(n5065) );
  XNOR U432 ( .A(in[22]), .B(in[1302]), .Z(n5064) );
  XNOR U433 ( .A(n5065), .B(n5064), .Z(n5066) );
  XNOR U434 ( .A(in[982]), .B(n5066), .Z(n6061) );
  XNOR U435 ( .A(n5370), .B(n6061), .Z(n8939) );
  XNOR U436 ( .A(in[1367]), .B(n8939), .Z(n6548) );
  XOR U437 ( .A(in[1375]), .B(in[735]), .Z(n5068) );
  XNOR U438 ( .A(in[95]), .B(in[415]), .Z(n5067) );
  XNOR U439 ( .A(n5068), .B(n5067), .Z(n5069) );
  XOR U440 ( .A(in[1055]), .B(n5069), .Z(n5736) );
  XOR U441 ( .A(in[1566]), .B(in[606]), .Z(n5071) );
  XNOR U442 ( .A(in[926]), .B(in[286]), .Z(n5070) );
  XNOR U443 ( .A(n5071), .B(n5070), .Z(n5072) );
  XOR U444 ( .A(in[1246]), .B(n5072), .Z(n5472) );
  XNOR U445 ( .A(n5736), .B(n5472), .Z(n8713) );
  XNOR U446 ( .A(in[991]), .B(n8713), .Z(n6545) );
  NAND U447 ( .A(n6548), .B(n6545), .Z(n5073) );
  XNOR U448 ( .A(n6153), .B(n5073), .Z(out[1011]) );
  XOR U449 ( .A(in[1527]), .B(in[567]), .Z(n5075) );
  XNOR U450 ( .A(in[887]), .B(in[247]), .Z(n5074) );
  XNOR U451 ( .A(n5075), .B(n5074), .Z(n5076) );
  XOR U452 ( .A(in[1207]), .B(n5076), .Z(n6185) );
  XOR U453 ( .A(in[1398]), .B(in[118]), .Z(n5078) );
  XNOR U454 ( .A(in[1078]), .B(in[758]), .Z(n5077) );
  XNOR U455 ( .A(n5078), .B(n5077), .Z(n5079) );
  XOR U456 ( .A(in[438]), .B(n5079), .Z(n6243) );
  XNOR U457 ( .A(n6185), .B(n6243), .Z(n8615) );
  XNOR U458 ( .A(in[183]), .B(n8615), .Z(n6158) );
  XOR U459 ( .A(in[343]), .B(in[663]), .Z(n5081) );
  XNOR U460 ( .A(in[23]), .B(in[1303]), .Z(n5080) );
  XNOR U461 ( .A(n5081), .B(n5080), .Z(n5082) );
  XOR U462 ( .A(in[983]), .B(n5082), .Z(n6064) );
  XOR U463 ( .A(in[152]), .B(in[1432]), .Z(n5084) );
  XNOR U464 ( .A(in[1112]), .B(in[792]), .Z(n5083) );
  XNOR U465 ( .A(n5084), .B(n5083), .Z(n5085) );
  XNOR U466 ( .A(in[472]), .B(n5085), .Z(n5396) );
  XNOR U467 ( .A(n6064), .B(n5396), .Z(n8942) );
  XNOR U468 ( .A(in[1368]), .B(n8942), .Z(n6552) );
  XOR U469 ( .A(in[1376]), .B(in[736]), .Z(n5087) );
  XNOR U470 ( .A(in[96]), .B(in[416]), .Z(n5086) );
  XNOR U471 ( .A(n5087), .B(n5086), .Z(n5088) );
  XOR U472 ( .A(in[1056]), .B(n5088), .Z(n5751) );
  XOR U473 ( .A(in[1567]), .B(in[607]), .Z(n5090) );
  XNOR U474 ( .A(in[927]), .B(in[287]), .Z(n5089) );
  XNOR U475 ( .A(n5090), .B(n5089), .Z(n5091) );
  XOR U476 ( .A(in[1247]), .B(n5091), .Z(n5487) );
  XNOR U477 ( .A(n5751), .B(n5487), .Z(n8715) );
  XNOR U478 ( .A(in[992]), .B(n8715), .Z(n6549) );
  NAND U479 ( .A(n6552), .B(n6549), .Z(n5092) );
  XNOR U480 ( .A(n6158), .B(n5092), .Z(out[1012]) );
  XOR U481 ( .A(in[1528]), .B(in[568]), .Z(n5094) );
  XNOR U482 ( .A(in[888]), .B(in[248]), .Z(n5093) );
  XNOR U483 ( .A(n5094), .B(n5093), .Z(n5095) );
  XOR U484 ( .A(in[1208]), .B(n5095), .Z(n6189) );
  XOR U485 ( .A(in[1399]), .B(in[119]), .Z(n5097) );
  XNOR U486 ( .A(in[1079]), .B(in[759]), .Z(n5096) );
  XNOR U487 ( .A(n5097), .B(n5096), .Z(n5098) );
  XOR U488 ( .A(in[439]), .B(n5098), .Z(n6247) );
  XNOR U489 ( .A(n6189), .B(n6247), .Z(n8619) );
  XNOR U490 ( .A(in[184]), .B(n8619), .Z(n6162) );
  XOR U491 ( .A(in[344]), .B(in[664]), .Z(n5100) );
  XNOR U492 ( .A(in[24]), .B(in[1304]), .Z(n5099) );
  XNOR U493 ( .A(n5100), .B(n5099), .Z(n5101) );
  XOR U494 ( .A(in[984]), .B(n5101), .Z(n6067) );
  XOR U495 ( .A(in[153]), .B(in[1433]), .Z(n5103) );
  XNOR U496 ( .A(in[1113]), .B(in[793]), .Z(n5102) );
  XNOR U497 ( .A(n5103), .B(n5102), .Z(n5104) );
  XNOR U498 ( .A(in[473]), .B(n5104), .Z(n5411) );
  XNOR U499 ( .A(n6067), .B(n5411), .Z(n8945) );
  XNOR U500 ( .A(in[1369]), .B(n8945), .Z(n6556) );
  XOR U501 ( .A(in[1377]), .B(in[737]), .Z(n5106) );
  XNOR U502 ( .A(in[97]), .B(in[417]), .Z(n5105) );
  XNOR U503 ( .A(n5106), .B(n5105), .Z(n5107) );
  XOR U504 ( .A(in[1057]), .B(n5107), .Z(n5766) );
  XOR U505 ( .A(in[1568]), .B(in[608]), .Z(n5109) );
  XNOR U506 ( .A(in[928]), .B(in[288]), .Z(n5108) );
  XNOR U507 ( .A(n5109), .B(n5108), .Z(n5110) );
  XOR U508 ( .A(in[1248]), .B(n5110), .Z(n5502) );
  XNOR U509 ( .A(n5766), .B(n5502), .Z(n8717) );
  XNOR U510 ( .A(in[993]), .B(n8717), .Z(n6553) );
  NAND U511 ( .A(n6556), .B(n6553), .Z(n5111) );
  XNOR U512 ( .A(n6162), .B(n5111), .Z(out[1013]) );
  XOR U513 ( .A(in[1529]), .B(in[569]), .Z(n5113) );
  XNOR U514 ( .A(in[889]), .B(in[249]), .Z(n5112) );
  XNOR U515 ( .A(n5113), .B(n5112), .Z(n5114) );
  XOR U516 ( .A(in[1209]), .B(n5114), .Z(n6193) );
  XOR U517 ( .A(in[1400]), .B(in[120]), .Z(n5116) );
  XNOR U518 ( .A(in[1080]), .B(in[760]), .Z(n5115) );
  XNOR U519 ( .A(n5116), .B(n5115), .Z(n5117) );
  XOR U520 ( .A(in[440]), .B(n5117), .Z(n6251) );
  XNOR U521 ( .A(n6193), .B(n6251), .Z(n8623) );
  XNOR U522 ( .A(in[185]), .B(n8623), .Z(n6166) );
  XOR U523 ( .A(in[345]), .B(in[665]), .Z(n5119) );
  XNOR U524 ( .A(in[25]), .B(in[1305]), .Z(n5118) );
  XNOR U525 ( .A(n5119), .B(n5118), .Z(n5120) );
  XOR U526 ( .A(in[985]), .B(n5120), .Z(n6070) );
  XOR U527 ( .A(in[154]), .B(in[1434]), .Z(n5122) );
  XNOR U528 ( .A(in[1114]), .B(in[794]), .Z(n5121) );
  XNOR U529 ( .A(n5122), .B(n5121), .Z(n5123) );
  XNOR U530 ( .A(in[474]), .B(n5123), .Z(n5426) );
  XNOR U531 ( .A(n6070), .B(n5426), .Z(n8948) );
  XNOR U532 ( .A(in[1370]), .B(n8948), .Z(n6561) );
  XOR U533 ( .A(in[1569]), .B(in[609]), .Z(n5125) );
  XNOR U534 ( .A(in[929]), .B(in[289]), .Z(n5124) );
  XNOR U535 ( .A(n5125), .B(n5124), .Z(n5126) );
  XOR U536 ( .A(in[1249]), .B(n5126), .Z(n5517) );
  XOR U537 ( .A(in[1378]), .B(in[738]), .Z(n5128) );
  XNOR U538 ( .A(in[98]), .B(in[418]), .Z(n5127) );
  XNOR U539 ( .A(n5128), .B(n5127), .Z(n5129) );
  XOR U540 ( .A(in[1058]), .B(n5129), .Z(n5781) );
  XNOR U541 ( .A(n5517), .B(n5781), .Z(n8719) );
  XNOR U542 ( .A(in[994]), .B(n8719), .Z(n6558) );
  NAND U543 ( .A(n6561), .B(n6558), .Z(n5130) );
  XNOR U544 ( .A(n6166), .B(n5130), .Z(out[1014]) );
  XOR U545 ( .A(in[1401]), .B(in[121]), .Z(n5132) );
  XNOR U546 ( .A(in[1081]), .B(in[761]), .Z(n5131) );
  XNOR U547 ( .A(n5132), .B(n5131), .Z(n5133) );
  XOR U548 ( .A(in[441]), .B(n5133), .Z(n6255) );
  XNOR U549 ( .A(n5134), .B(n6255), .Z(n8345) );
  XNOR U550 ( .A(in[186]), .B(n8345), .Z(n6170) );
  XOR U551 ( .A(in[155]), .B(in[1435]), .Z(n5136) );
  XNOR U552 ( .A(in[1115]), .B(in[795]), .Z(n5135) );
  XNOR U553 ( .A(n5136), .B(n5135), .Z(n5137) );
  XOR U554 ( .A(in[475]), .B(n5137), .Z(n5441) );
  XOR U555 ( .A(in[346]), .B(in[666]), .Z(n5139) );
  XNOR U556 ( .A(in[26]), .B(in[1306]), .Z(n5138) );
  XNOR U557 ( .A(n5139), .B(n5138), .Z(n5140) );
  XNOR U558 ( .A(in[986]), .B(n5140), .Z(n6073) );
  XNOR U559 ( .A(n5441), .B(n6073), .Z(n8955) );
  XNOR U560 ( .A(in[1371]), .B(n8955), .Z(n6565) );
  XOR U561 ( .A(in[1379]), .B(in[739]), .Z(n5142) );
  XNOR U562 ( .A(in[99]), .B(in[419]), .Z(n5141) );
  XNOR U563 ( .A(n5142), .B(n5141), .Z(n5143) );
  XNOR U564 ( .A(in[1059]), .B(n5143), .Z(n5796) );
  XNOR U565 ( .A(n5144), .B(n5796), .Z(n8721) );
  XNOR U566 ( .A(in[995]), .B(n8721), .Z(n6562) );
  NAND U567 ( .A(n6565), .B(n6562), .Z(n5145) );
  XNOR U568 ( .A(n6170), .B(n5145), .Z(out[1015]) );
  XOR U569 ( .A(in[1402]), .B(in[122]), .Z(n5147) );
  XNOR U570 ( .A(in[1082]), .B(in[762]), .Z(n5146) );
  XNOR U571 ( .A(n5147), .B(n5146), .Z(n5148) );
  XOR U572 ( .A(in[442]), .B(n5148), .Z(n6259) );
  XOR U573 ( .A(in[1531]), .B(in[571]), .Z(n5150) );
  XNOR U574 ( .A(in[1211]), .B(in[251]), .Z(n5149) );
  XNOR U575 ( .A(n5150), .B(n5149), .Z(n5151) );
  XOR U576 ( .A(in[891]), .B(n5151), .Z(n5223) );
  XNOR U577 ( .A(n6259), .B(n5223), .Z(n8349) );
  XNOR U578 ( .A(in[187]), .B(n8349), .Z(n6174) );
  XOR U579 ( .A(in[156]), .B(in[1436]), .Z(n5153) );
  XNOR U580 ( .A(in[1116]), .B(in[796]), .Z(n5152) );
  XNOR U581 ( .A(n5153), .B(n5152), .Z(n5154) );
  XOR U582 ( .A(in[476]), .B(n5154), .Z(n5456) );
  XOR U583 ( .A(in[347]), .B(in[667]), .Z(n5156) );
  XNOR U584 ( .A(in[27]), .B(in[1307]), .Z(n5155) );
  XNOR U585 ( .A(n5156), .B(n5155), .Z(n5157) );
  XNOR U586 ( .A(in[987]), .B(n5157), .Z(n6076) );
  XNOR U587 ( .A(n5456), .B(n6076), .Z(n8958) );
  XNOR U588 ( .A(in[1372]), .B(n8958), .Z(n6569) );
  XOR U589 ( .A(in[1060]), .B(in[420]), .Z(n5159) );
  XNOR U590 ( .A(in[740]), .B(in[1380]), .Z(n5158) );
  XNOR U591 ( .A(n5159), .B(n5158), .Z(n5160) );
  XOR U592 ( .A(in[100]), .B(n5160), .Z(n5811) );
  XOR U593 ( .A(in[1571]), .B(in[611]), .Z(n5162) );
  XNOR U594 ( .A(in[931]), .B(in[291]), .Z(n5161) );
  XNOR U595 ( .A(n5162), .B(n5161), .Z(n5163) );
  XOR U596 ( .A(in[1251]), .B(n5163), .Z(n5227) );
  XNOR U597 ( .A(n5811), .B(n5227), .Z(n8723) );
  XNOR U598 ( .A(in[996]), .B(n8723), .Z(n6566) );
  NAND U599 ( .A(n6569), .B(n6566), .Z(n5164) );
  XNOR U600 ( .A(n6174), .B(n5164), .Z(out[1016]) );
  XOR U601 ( .A(in[1403]), .B(in[123]), .Z(n5166) );
  XNOR U602 ( .A(in[1083]), .B(in[763]), .Z(n5165) );
  XNOR U603 ( .A(n5166), .B(n5165), .Z(n5167) );
  XOR U604 ( .A(in[443]), .B(n5167), .Z(n6263) );
  XOR U605 ( .A(in[1532]), .B(in[572]), .Z(n5169) );
  XNOR U606 ( .A(in[1212]), .B(in[252]), .Z(n5168) );
  XNOR U607 ( .A(n5169), .B(n5168), .Z(n5170) );
  XOR U608 ( .A(in[892]), .B(n5170), .Z(n5388) );
  XNOR U609 ( .A(n6263), .B(n5388), .Z(n8353) );
  XNOR U610 ( .A(in[188]), .B(n8353), .Z(n6178) );
  XOR U611 ( .A(in[157]), .B(in[1437]), .Z(n5172) );
  XNOR U612 ( .A(in[1117]), .B(in[797]), .Z(n5171) );
  XNOR U613 ( .A(n5172), .B(n5171), .Z(n5173) );
  XOR U614 ( .A(in[477]), .B(n5173), .Z(n5471) );
  XOR U615 ( .A(in[348]), .B(in[668]), .Z(n5175) );
  XNOR U616 ( .A(in[28]), .B(in[1308]), .Z(n5174) );
  XNOR U617 ( .A(n5175), .B(n5174), .Z(n5176) );
  XNOR U618 ( .A(in[988]), .B(n5176), .Z(n6079) );
  XNOR U619 ( .A(n5471), .B(n6079), .Z(n8961) );
  XNOR U620 ( .A(in[1373]), .B(n8961), .Z(n6573) );
  XOR U621 ( .A(in[1572]), .B(in[612]), .Z(n5178) );
  XNOR U622 ( .A(in[932]), .B(in[292]), .Z(n5177) );
  XNOR U623 ( .A(n5178), .B(n5177), .Z(n5179) );
  XOR U624 ( .A(in[1252]), .B(n5179), .Z(n5390) );
  XNOR U625 ( .A(n5180), .B(n5390), .Z(n8725) );
  XNOR U626 ( .A(in[997]), .B(n8725), .Z(n6570) );
  NAND U627 ( .A(n6573), .B(n6570), .Z(n5181) );
  XNOR U628 ( .A(n6178), .B(n5181), .Z(out[1017]) );
  XOR U629 ( .A(in[1404]), .B(in[124]), .Z(n5183) );
  XNOR U630 ( .A(in[1084]), .B(in[764]), .Z(n5182) );
  XNOR U631 ( .A(n5183), .B(n5182), .Z(n5184) );
  XOR U632 ( .A(in[444]), .B(n5184), .Z(n6267) );
  XOR U633 ( .A(in[1533]), .B(in[573]), .Z(n5186) );
  XNOR U634 ( .A(in[1213]), .B(in[253]), .Z(n5185) );
  XNOR U635 ( .A(n5186), .B(n5185), .Z(n5187) );
  XOR U636 ( .A(in[893]), .B(n5187), .Z(n5547) );
  XNOR U637 ( .A(n6267), .B(n5547), .Z(n8357) );
  XNOR U638 ( .A(in[189]), .B(n8357), .Z(n6182) );
  XOR U639 ( .A(in[158]), .B(in[1438]), .Z(n5189) );
  XNOR U640 ( .A(in[1118]), .B(in[798]), .Z(n5188) );
  XNOR U641 ( .A(n5189), .B(n5188), .Z(n5190) );
  XOR U642 ( .A(in[478]), .B(n5190), .Z(n5486) );
  XOR U643 ( .A(in[349]), .B(in[669]), .Z(n5192) );
  XNOR U644 ( .A(in[29]), .B(in[1309]), .Z(n5191) );
  XNOR U645 ( .A(n5192), .B(n5191), .Z(n5193) );
  XNOR U646 ( .A(in[989]), .B(n5193), .Z(n6083) );
  XNOR U647 ( .A(n5486), .B(n6083), .Z(n8964) );
  XNOR U648 ( .A(in[1374]), .B(n8964), .Z(n6577) );
  XOR U649 ( .A(in[1062]), .B(in[422]), .Z(n5195) );
  XNOR U650 ( .A(in[742]), .B(in[1382]), .Z(n5194) );
  XNOR U651 ( .A(n5195), .B(n5194), .Z(n5196) );
  XOR U652 ( .A(in[102]), .B(n5196), .Z(n5231) );
  XOR U653 ( .A(in[1573]), .B(in[613]), .Z(n5198) );
  XNOR U654 ( .A(in[933]), .B(in[293]), .Z(n5197) );
  XNOR U655 ( .A(n5198), .B(n5197), .Z(n5199) );
  XOR U656 ( .A(in[1253]), .B(n5199), .Z(n5549) );
  XNOR U657 ( .A(n5231), .B(n5549), .Z(n8731) );
  XNOR U658 ( .A(in[998]), .B(n8731), .Z(n6574) );
  NAND U659 ( .A(n6577), .B(n6574), .Z(n5200) );
  XNOR U660 ( .A(n6182), .B(n5200), .Z(out[1018]) );
  XOR U661 ( .A(in[1405]), .B(in[125]), .Z(n5202) );
  XNOR U662 ( .A(in[1085]), .B(in[765]), .Z(n5201) );
  XNOR U663 ( .A(n5202), .B(n5201), .Z(n5203) );
  XOR U664 ( .A(in[445]), .B(n5203), .Z(n6271) );
  XOR U665 ( .A(in[1534]), .B(in[894]), .Z(n5205) );
  XNOR U666 ( .A(in[574]), .B(in[1214]), .Z(n5204) );
  XNOR U667 ( .A(n5205), .B(n5204), .Z(n5206) );
  XOR U668 ( .A(in[254]), .B(n5206), .Z(n5684) );
  XNOR U669 ( .A(n6271), .B(n5684), .Z(n8361) );
  XNOR U670 ( .A(in[190]), .B(n8361), .Z(n6186) );
  XOR U671 ( .A(in[1439]), .B(in[479]), .Z(n5208) );
  XNOR U672 ( .A(in[799]), .B(in[159]), .Z(n5207) );
  XNOR U673 ( .A(n5208), .B(n5207), .Z(n5209) );
  XOR U674 ( .A(in[1119]), .B(n5209), .Z(n5501) );
  XOR U675 ( .A(in[350]), .B(in[670]), .Z(n5211) );
  XNOR U676 ( .A(in[30]), .B(in[1310]), .Z(n5210) );
  XNOR U677 ( .A(n5211), .B(n5210), .Z(n5212) );
  XNOR U678 ( .A(in[990]), .B(n5212), .Z(n6086) );
  XNOR U679 ( .A(n5501), .B(n6086), .Z(n8967) );
  XNOR U680 ( .A(in[1375]), .B(n8967), .Z(n6581) );
  XOR U681 ( .A(in[1063]), .B(in[423]), .Z(n5214) );
  XNOR U682 ( .A(in[743]), .B(in[1383]), .Z(n5213) );
  XNOR U683 ( .A(n5214), .B(n5213), .Z(n5215) );
  XOR U684 ( .A(in[103]), .B(n5215), .Z(n5394) );
  XOR U685 ( .A(in[1574]), .B(in[614]), .Z(n5217) );
  XNOR U686 ( .A(in[934]), .B(in[294]), .Z(n5216) );
  XNOR U687 ( .A(n5217), .B(n5216), .Z(n5218) );
  XOR U688 ( .A(in[1254]), .B(n5218), .Z(n5593) );
  XNOR U689 ( .A(n5394), .B(n5593), .Z(n8733) );
  XNOR U690 ( .A(in[999]), .B(n8733), .Z(n6578) );
  NAND U691 ( .A(n6581), .B(n6578), .Z(n5219) );
  XNOR U692 ( .A(n6186), .B(n5219), .Z(out[1019]) );
  XOR U693 ( .A(in[1340]), .B(in[60]), .Z(n5221) );
  XNOR U694 ( .A(in[700]), .B(in[380]), .Z(n5220) );
  XNOR U695 ( .A(n5221), .B(n5220), .Z(n5222) );
  XOR U696 ( .A(in[1020]), .B(n5222), .Z(n5678) );
  XNOR U697 ( .A(n5223), .B(n5678), .Z(n8403) );
  XNOR U698 ( .A(in[636]), .B(n8403), .Z(n7359) );
  XOR U699 ( .A(in[162]), .B(in[1442]), .Z(n5225) );
  XNOR U700 ( .A(in[802]), .B(in[1122]), .Z(n5224) );
  XNOR U701 ( .A(n5225), .B(n5224), .Z(n5226) );
  XNOR U702 ( .A(in[482]), .B(n5226), .Z(n5278) );
  XNOR U703 ( .A(n5227), .B(n5278), .Z(n8500) );
  XNOR U704 ( .A(in[227]), .B(n8500), .Z(n7652) );
  XOR U705 ( .A(in[1511]), .B(in[551]), .Z(n5229) );
  XNOR U706 ( .A(in[871]), .B(in[231]), .Z(n5228) );
  XNOR U707 ( .A(n5229), .B(n5228), .Z(n5230) );
  XOR U708 ( .A(in[1191]), .B(n5230), .Z(n6120) );
  XNOR U709 ( .A(n5231), .B(n6120), .Z(n8541) );
  XNOR U710 ( .A(in[1447]), .B(n8541), .Z(n7649) );
  NAND U711 ( .A(n7652), .B(n7649), .Z(n5232) );
  XNOR U712 ( .A(n7359), .B(n5232), .Z(out[101]) );
  XOR U713 ( .A(in[1406]), .B(in[126]), .Z(n5234) );
  XNOR U714 ( .A(in[1086]), .B(in[766]), .Z(n5233) );
  XNOR U715 ( .A(n5234), .B(n5233), .Z(n5235) );
  XOR U716 ( .A(in[446]), .B(n5235), .Z(n6276) );
  XOR U717 ( .A(in[1535]), .B(in[575]), .Z(n5237) );
  XNOR U718 ( .A(in[895]), .B(in[255]), .Z(n5236) );
  XNOR U719 ( .A(n5237), .B(n5236), .Z(n5238) );
  XOR U720 ( .A(in[1215]), .B(n5238), .Z(n5831) );
  XNOR U721 ( .A(n6276), .B(n5831), .Z(n8365) );
  XNOR U722 ( .A(in[191]), .B(n8365), .Z(n6190) );
  XOR U723 ( .A(in[1440]), .B(in[480]), .Z(n5240) );
  XNOR U724 ( .A(in[800]), .B(in[160]), .Z(n5239) );
  XNOR U725 ( .A(n5240), .B(n5239), .Z(n5241) );
  XOR U726 ( .A(in[1120]), .B(n5241), .Z(n5516) );
  XOR U727 ( .A(in[351]), .B(in[671]), .Z(n5243) );
  XNOR U728 ( .A(in[31]), .B(in[1311]), .Z(n5242) );
  XNOR U729 ( .A(n5243), .B(n5242), .Z(n5244) );
  XNOR U730 ( .A(in[991]), .B(n5244), .Z(n6089) );
  XNOR U731 ( .A(n5516), .B(n6089), .Z(n8970) );
  XNOR U732 ( .A(in[1376]), .B(n8970), .Z(n6585) );
  XOR U733 ( .A(in[1064]), .B(in[424]), .Z(n5246) );
  XNOR U734 ( .A(in[744]), .B(in[1384]), .Z(n5245) );
  XNOR U735 ( .A(n5246), .B(n5245), .Z(n5247) );
  XOR U736 ( .A(in[104]), .B(n5247), .Z(n5553) );
  XOR U737 ( .A(in[1575]), .B(in[615]), .Z(n5249) );
  XNOR U738 ( .A(in[935]), .B(in[295]), .Z(n5248) );
  XNOR U739 ( .A(n5249), .B(n5248), .Z(n5250) );
  XOR U740 ( .A(in[1255]), .B(n5250), .Z(n5606) );
  XNOR U741 ( .A(n5553), .B(n5606), .Z(n8735) );
  XNOR U742 ( .A(in[1000]), .B(n8735), .Z(n6582) );
  NAND U743 ( .A(n6585), .B(n6582), .Z(n5251) );
  XNOR U744 ( .A(n6190), .B(n5251), .Z(out[1020]) );
  XOR U745 ( .A(in[1407]), .B(in[127]), .Z(n5253) );
  XNOR U746 ( .A(in[1087]), .B(in[767]), .Z(n5252) );
  XNOR U747 ( .A(n5253), .B(n5252), .Z(n5254) );
  XOR U748 ( .A(in[447]), .B(n5254), .Z(n6279) );
  XOR U749 ( .A(in[1472]), .B(in[512]), .Z(n5256) );
  XNOR U750 ( .A(in[832]), .B(in[192]), .Z(n5255) );
  XNOR U751 ( .A(n5256), .B(n5255), .Z(n5257) );
  XOR U752 ( .A(in[1152]), .B(n5257), .Z(n5898) );
  XNOR U753 ( .A(n6279), .B(n5898), .Z(n8369) );
  XNOR U754 ( .A(in[128]), .B(n8369), .Z(n6194) );
  XOR U755 ( .A(in[352]), .B(in[672]), .Z(n5259) );
  XNOR U756 ( .A(in[32]), .B(in[1312]), .Z(n5258) );
  XNOR U757 ( .A(n5259), .B(n5258), .Z(n5260) );
  XNOR U758 ( .A(in[992]), .B(n5260), .Z(n6092) );
  XNOR U759 ( .A(n5261), .B(n6092), .Z(n8973) );
  XNOR U760 ( .A(in[1377]), .B(n8973), .Z(n6589) );
  XOR U761 ( .A(in[1065]), .B(in[425]), .Z(n5263) );
  XNOR U762 ( .A(in[745]), .B(in[1385]), .Z(n5262) );
  XNOR U763 ( .A(n5263), .B(n5262), .Z(n5264) );
  XOR U764 ( .A(in[105]), .B(n5264), .Z(n5688) );
  XOR U765 ( .A(in[1576]), .B(in[616]), .Z(n5266) );
  XNOR U766 ( .A(in[936]), .B(in[296]), .Z(n5265) );
  XNOR U767 ( .A(n5266), .B(n5265), .Z(n5267) );
  XOR U768 ( .A(in[1256]), .B(n5267), .Z(n5619) );
  XNOR U769 ( .A(n5688), .B(n5619), .Z(n8737) );
  XNOR U770 ( .A(in[1001]), .B(n8737), .Z(n6586) );
  NAND U771 ( .A(n6589), .B(n6586), .Z(n5268) );
  XNOR U772 ( .A(n6194), .B(n5268), .Z(out[1021]) );
  XOR U773 ( .A(in[1344]), .B(in[64]), .Z(n5270) );
  XNOR U774 ( .A(in[1024]), .B(in[384]), .Z(n5269) );
  XNOR U775 ( .A(n5270), .B(n5269), .Z(n5271) );
  XOR U776 ( .A(in[704]), .B(n5271), .Z(n6284) );
  XOR U777 ( .A(in[1473]), .B(in[513]), .Z(n5273) );
  XNOR U778 ( .A(in[833]), .B(in[193]), .Z(n5272) );
  XNOR U779 ( .A(n5273), .B(n5272), .Z(n5274) );
  XOR U780 ( .A(in[1153]), .B(n5274), .Z(n5951) );
  XNOR U781 ( .A(n6284), .B(n5951), .Z(n8373) );
  XNOR U782 ( .A(in[129]), .B(n8373), .Z(n6197) );
  XOR U783 ( .A(in[353]), .B(in[673]), .Z(n5276) );
  XNOR U784 ( .A(in[33]), .B(in[1313]), .Z(n5275) );
  XNOR U785 ( .A(n5276), .B(n5275), .Z(n5277) );
  XOR U786 ( .A(in[993]), .B(n5277), .Z(n6095) );
  XNOR U787 ( .A(n6095), .B(n5278), .Z(n8976) );
  XNOR U788 ( .A(in[1378]), .B(n8976), .Z(n6593) );
  XOR U789 ( .A(in[1577]), .B(in[617]), .Z(n5280) );
  XNOR U790 ( .A(in[937]), .B(in[297]), .Z(n5279) );
  XNOR U791 ( .A(n5280), .B(n5279), .Z(n5281) );
  XOR U792 ( .A(in[1257]), .B(n5281), .Z(n5632) );
  XNOR U793 ( .A(n5282), .B(n5632), .Z(n8739) );
  XNOR U794 ( .A(in[1002]), .B(n8739), .Z(n6590) );
  NAND U795 ( .A(n6593), .B(n6590), .Z(n5283) );
  XNOR U796 ( .A(n6197), .B(n5283), .Z(out[1022]) );
  XOR U797 ( .A(n8377), .B(in[130]), .Z(n6199) );
  XOR U798 ( .A(in[354]), .B(in[674]), .Z(n5285) );
  XNOR U799 ( .A(in[34]), .B(in[1314]), .Z(n5284) );
  XNOR U800 ( .A(n5285), .B(n5284), .Z(n5286) );
  XOR U801 ( .A(in[994]), .B(n5286), .Z(n6098) );
  XOR U802 ( .A(in[163]), .B(in[1443]), .Z(n5288) );
  XNOR U803 ( .A(in[803]), .B(in[1123]), .Z(n5287) );
  XNOR U804 ( .A(n5288), .B(n5287), .Z(n5289) );
  XNOR U805 ( .A(in[483]), .B(n5289), .Z(n5389) );
  XNOR U806 ( .A(n6098), .B(n5389), .Z(n8979) );
  XNOR U807 ( .A(in[1379]), .B(n8979), .Z(n6597) );
  XOR U808 ( .A(in[1578]), .B(in[618]), .Z(n5291) );
  XNOR U809 ( .A(in[938]), .B(in[298]), .Z(n5290) );
  XNOR U810 ( .A(n5291), .B(n5290), .Z(n5292) );
  XOR U811 ( .A(in[1258]), .B(n5292), .Z(n5645) );
  XNOR U812 ( .A(n5293), .B(n5645), .Z(n8741) );
  XNOR U813 ( .A(in[1003]), .B(n8741), .Z(n6594) );
  NAND U814 ( .A(n6597), .B(n6594), .Z(n5294) );
  XNOR U815 ( .A(n6199), .B(n5294), .Z(out[1023]) );
  XOR U816 ( .A(n5296), .B(n5295), .Z(n8432) );
  XNOR U817 ( .A(in[531]), .B(n8432), .Z(n6203) );
  XOR U818 ( .A(in[1346]), .B(in[66]), .Z(n5298) );
  XNOR U819 ( .A(in[1026]), .B(in[386]), .Z(n5297) );
  XNOR U820 ( .A(n5298), .B(n5297), .Z(n5299) );
  XOR U821 ( .A(in[706]), .B(n5299), .Z(n6292) );
  XOR U822 ( .A(in[1475]), .B(in[515]), .Z(n5301) );
  XNOR U823 ( .A(in[835]), .B(in[195]), .Z(n5300) );
  XNOR U824 ( .A(n5301), .B(n5300), .Z(n5302) );
  XNOR U825 ( .A(in[1155]), .B(n5302), .Z(n6003) );
  XNOR U826 ( .A(n6292), .B(n6003), .Z(n8381) );
  XNOR U827 ( .A(in[131]), .B(n8381), .Z(n9438) );
  XOR U828 ( .A(in[164]), .B(in[1444]), .Z(n5304) );
  XNOR U829 ( .A(in[804]), .B(in[1124]), .Z(n5303) );
  XNOR U830 ( .A(n5304), .B(n5303), .Z(n5305) );
  XOR U831 ( .A(in[484]), .B(n5305), .Z(n5548) );
  XOR U832 ( .A(in[35]), .B(in[675]), .Z(n5307) );
  XNOR U833 ( .A(in[355]), .B(in[1315]), .Z(n5306) );
  XNOR U834 ( .A(n5307), .B(n5306), .Z(n5308) );
  XOR U835 ( .A(in[995]), .B(n5308), .Z(n6101) );
  XNOR U836 ( .A(n5548), .B(n6101), .Z(n8982) );
  XNOR U837 ( .A(in[1380]), .B(n8982), .Z(n9435) );
  NAND U838 ( .A(n9438), .B(n9435), .Z(n5309) );
  XNOR U839 ( .A(n6203), .B(n5309), .Z(out[1024]) );
  XNOR U840 ( .A(n5311), .B(n5310), .Z(n8436) );
  XNOR U841 ( .A(in[532]), .B(n8436), .Z(n6207) );
  XOR U842 ( .A(in[1347]), .B(in[67]), .Z(n5313) );
  XNOR U843 ( .A(in[1027]), .B(in[387]), .Z(n5312) );
  XNOR U844 ( .A(n5313), .B(n5312), .Z(n5314) );
  XOR U845 ( .A(in[707]), .B(n5314), .Z(n6296) );
  XOR U846 ( .A(in[1476]), .B(in[516]), .Z(n5316) );
  XNOR U847 ( .A(in[836]), .B(in[196]), .Z(n5315) );
  XNOR U848 ( .A(n5316), .B(n5315), .Z(n5317) );
  XNOR U849 ( .A(in[1156]), .B(n5317), .Z(n6006) );
  XNOR U850 ( .A(n6296), .B(n6006), .Z(n8389) );
  XNOR U851 ( .A(in[132]), .B(n8389), .Z(n9442) );
  XOR U852 ( .A(in[36]), .B(in[676]), .Z(n5319) );
  XNOR U853 ( .A(in[356]), .B(in[1316]), .Z(n5318) );
  XNOR U854 ( .A(n5319), .B(n5318), .Z(n5320) );
  XOR U855 ( .A(in[996]), .B(n5320), .Z(n6104) );
  XOR U856 ( .A(in[1445]), .B(in[165]), .Z(n5322) );
  XNOR U857 ( .A(in[805]), .B(in[1125]), .Z(n5321) );
  XNOR U858 ( .A(n5322), .B(n5321), .Z(n5323) );
  XOR U859 ( .A(in[485]), .B(n5323), .Z(n5592) );
  XNOR U860 ( .A(n6104), .B(n5592), .Z(n8989) );
  XNOR U861 ( .A(in[1381]), .B(n8989), .Z(n9439) );
  NAND U862 ( .A(n9442), .B(n9439), .Z(n5324) );
  XNOR U863 ( .A(n6207), .B(n5324), .Z(out[1025]) );
  XNOR U864 ( .A(n5326), .B(n5325), .Z(n8440) );
  XNOR U865 ( .A(in[533]), .B(n8440), .Z(n6211) );
  XOR U866 ( .A(in[1348]), .B(in[68]), .Z(n5328) );
  XNOR U867 ( .A(in[1028]), .B(in[388]), .Z(n5327) );
  XNOR U868 ( .A(n5328), .B(n5327), .Z(n5329) );
  XOR U869 ( .A(in[708]), .B(n5329), .Z(n6300) );
  XOR U870 ( .A(in[1477]), .B(in[517]), .Z(n5331) );
  XNOR U871 ( .A(in[837]), .B(in[197]), .Z(n5330) );
  XNOR U872 ( .A(n5331), .B(n5330), .Z(n5332) );
  XNOR U873 ( .A(in[1157]), .B(n5332), .Z(n6009) );
  XNOR U874 ( .A(n6300), .B(n6009), .Z(n8393) );
  XNOR U875 ( .A(in[133]), .B(n8393), .Z(n9446) );
  XOR U876 ( .A(in[166]), .B(in[806]), .Z(n5334) );
  XNOR U877 ( .A(in[1126]), .B(in[486]), .Z(n5333) );
  XNOR U878 ( .A(n5334), .B(n5333), .Z(n5335) );
  XOR U879 ( .A(in[1446]), .B(n5335), .Z(n5605) );
  XOR U880 ( .A(in[37]), .B(in[677]), .Z(n5337) );
  XNOR U881 ( .A(in[357]), .B(in[1317]), .Z(n5336) );
  XNOR U882 ( .A(n5337), .B(n5336), .Z(n5338) );
  XOR U883 ( .A(in[997]), .B(n5338), .Z(n6107) );
  XNOR U884 ( .A(n5605), .B(n6107), .Z(n8992) );
  XNOR U885 ( .A(in[1382]), .B(n8992), .Z(n9443) );
  NAND U886 ( .A(n9446), .B(n9443), .Z(n5339) );
  XNOR U887 ( .A(n6211), .B(n5339), .Z(out[1026]) );
  XOR U888 ( .A(n5341), .B(n5340), .Z(n8444) );
  XNOR U889 ( .A(in[534]), .B(n8444), .Z(n6215) );
  XOR U890 ( .A(in[1349]), .B(in[69]), .Z(n5343) );
  XNOR U891 ( .A(in[1029]), .B(in[389]), .Z(n5342) );
  XNOR U892 ( .A(n5343), .B(n5342), .Z(n5344) );
  XOR U893 ( .A(in[709]), .B(n5344), .Z(n6304) );
  XOR U894 ( .A(in[1478]), .B(in[518]), .Z(n5346) );
  XNOR U895 ( .A(in[838]), .B(in[198]), .Z(n5345) );
  XNOR U896 ( .A(n5346), .B(n5345), .Z(n5347) );
  XNOR U897 ( .A(in[1158]), .B(n5347), .Z(n6012) );
  XNOR U898 ( .A(n6304), .B(n6012), .Z(n8397) );
  XNOR U899 ( .A(in[134]), .B(n8397), .Z(n9450) );
  XOR U900 ( .A(in[38]), .B(in[678]), .Z(n5349) );
  XNOR U901 ( .A(in[358]), .B(in[1318]), .Z(n5348) );
  XNOR U902 ( .A(n5349), .B(n5348), .Z(n5350) );
  XOR U903 ( .A(in[998]), .B(n5350), .Z(n6111) );
  XOR U904 ( .A(in[167]), .B(in[807]), .Z(n5352) );
  XNOR U905 ( .A(in[1127]), .B(in[487]), .Z(n5351) );
  XNOR U906 ( .A(n5352), .B(n5351), .Z(n5353) );
  XOR U907 ( .A(in[1447]), .B(n5353), .Z(n5618) );
  XNOR U908 ( .A(n6111), .B(n5618), .Z(n8771) );
  XNOR U909 ( .A(in[1383]), .B(n8771), .Z(n9447) );
  NAND U910 ( .A(n9450), .B(n9447), .Z(n5354) );
  XNOR U911 ( .A(n6215), .B(n5354), .Z(out[1027]) );
  XOR U912 ( .A(n5356), .B(n5355), .Z(n8448) );
  XNOR U913 ( .A(in[535]), .B(n8448), .Z(n6219) );
  XOR U914 ( .A(in[1350]), .B(in[70]), .Z(n5358) );
  XNOR U915 ( .A(in[1030]), .B(in[390]), .Z(n5357) );
  XNOR U916 ( .A(n5358), .B(n5357), .Z(n5359) );
  XOR U917 ( .A(in[710]), .B(n5359), .Z(n6308) );
  XOR U918 ( .A(in[199]), .B(in[1479]), .Z(n5361) );
  XNOR U919 ( .A(in[1159]), .B(in[839]), .Z(n5360) );
  XNOR U920 ( .A(n5361), .B(n5360), .Z(n5362) );
  XNOR U921 ( .A(in[519]), .B(n5362), .Z(n6015) );
  XNOR U922 ( .A(n6308), .B(n6015), .Z(n8401) );
  XNOR U923 ( .A(in[135]), .B(n8401), .Z(n9454) );
  XOR U924 ( .A(in[168]), .B(in[1448]), .Z(n5364) );
  XNOR U925 ( .A(in[1128]), .B(in[808]), .Z(n5363) );
  XNOR U926 ( .A(n5364), .B(n5363), .Z(n5365) );
  XOR U927 ( .A(in[488]), .B(n5365), .Z(n5631) );
  XOR U928 ( .A(in[39]), .B(in[679]), .Z(n5367) );
  XNOR U929 ( .A(in[359]), .B(in[1319]), .Z(n5366) );
  XNOR U930 ( .A(n5367), .B(n5366), .Z(n5368) );
  XOR U931 ( .A(in[999]), .B(n5368), .Z(n6115) );
  XNOR U932 ( .A(n5631), .B(n6115), .Z(n8774) );
  XNOR U933 ( .A(in[1384]), .B(n8774), .Z(n9451) );
  NAND U934 ( .A(n9454), .B(n9451), .Z(n5369) );
  XNOR U935 ( .A(n6219), .B(n5369), .Z(out[1028]) );
  XNOR U936 ( .A(n5371), .B(n5370), .Z(n8452) );
  XNOR U937 ( .A(in[536]), .B(n8452), .Z(n6223) );
  XOR U938 ( .A(in[1351]), .B(in[711]), .Z(n5373) );
  XNOR U939 ( .A(in[1031]), .B(in[391]), .Z(n5372) );
  XNOR U940 ( .A(n5373), .B(n5372), .Z(n5374) );
  XOR U941 ( .A(in[71]), .B(n5374), .Z(n6312) );
  XOR U942 ( .A(in[1480]), .B(in[520]), .Z(n5376) );
  XNOR U943 ( .A(in[840]), .B(in[200]), .Z(n5375) );
  XNOR U944 ( .A(n5376), .B(n5375), .Z(n5377) );
  XNOR U945 ( .A(in[1160]), .B(n5377), .Z(n6020) );
  XNOR U946 ( .A(n6312), .B(n6020), .Z(n8405) );
  XNOR U947 ( .A(in[136]), .B(n8405), .Z(n9458) );
  XOR U948 ( .A(in[680]), .B(in[1320]), .Z(n5379) );
  XNOR U949 ( .A(in[40]), .B(in[360]), .Z(n5378) );
  XNOR U950 ( .A(n5379), .B(n5378), .Z(n5380) );
  XOR U951 ( .A(in[1000]), .B(n5380), .Z(n6119) );
  XOR U952 ( .A(in[169]), .B(in[1449]), .Z(n5382) );
  XNOR U953 ( .A(in[1129]), .B(in[809]), .Z(n5381) );
  XNOR U954 ( .A(n5382), .B(n5381), .Z(n5383) );
  XOR U955 ( .A(in[489]), .B(n5383), .Z(n5644) );
  XNOR U956 ( .A(n6119), .B(n5644), .Z(n8781) );
  XNOR U957 ( .A(in[1385]), .B(n8781), .Z(n9455) );
  NAND U958 ( .A(n9458), .B(n9455), .Z(n5384) );
  XNOR U959 ( .A(n6223), .B(n5384), .Z(out[1029]) );
  XOR U960 ( .A(in[1341]), .B(in[61]), .Z(n5386) );
  XNOR U961 ( .A(in[701]), .B(in[381]), .Z(n5385) );
  XNOR U962 ( .A(n5386), .B(n5385), .Z(n5387) );
  XOR U963 ( .A(in[1021]), .B(n5387), .Z(n5701) );
  XNOR U964 ( .A(n5388), .B(n5701), .Z(n8407) );
  XNOR U965 ( .A(in[637]), .B(n8407), .Z(n7362) );
  XNOR U966 ( .A(n5390), .B(n5389), .Z(n8504) );
  XNOR U967 ( .A(in[228]), .B(n8504), .Z(n7666) );
  XOR U968 ( .A(in[1512]), .B(in[552]), .Z(n5392) );
  XNOR U969 ( .A(in[872]), .B(in[232]), .Z(n5391) );
  XNOR U970 ( .A(n5392), .B(n5391), .Z(n5393) );
  XOR U971 ( .A(in[1192]), .B(n5393), .Z(n6124) );
  XNOR U972 ( .A(n5394), .B(n6124), .Z(n8545) );
  XNOR U973 ( .A(in[1448]), .B(n8545), .Z(n7663) );
  NAND U974 ( .A(n7666), .B(n7663), .Z(n5395) );
  XNOR U975 ( .A(n7362), .B(n5395), .Z(out[102]) );
  XOR U976 ( .A(n5397), .B(n5396), .Z(n8456) );
  XNOR U977 ( .A(in[537]), .B(n8456), .Z(n6227) );
  XOR U978 ( .A(in[1352]), .B(in[712]), .Z(n5399) );
  XNOR U979 ( .A(in[1032]), .B(in[392]), .Z(n5398) );
  XNOR U980 ( .A(n5399), .B(n5398), .Z(n5400) );
  XOR U981 ( .A(in[72]), .B(n5400), .Z(n6317) );
  XOR U982 ( .A(in[1481]), .B(in[521]), .Z(n5402) );
  XNOR U983 ( .A(in[841]), .B(in[201]), .Z(n5401) );
  XNOR U984 ( .A(n5402), .B(n5401), .Z(n5403) );
  XNOR U985 ( .A(in[1161]), .B(n5403), .Z(n6023) );
  XNOR U986 ( .A(n6317), .B(n6023), .Z(n8409) );
  XNOR U987 ( .A(in[137]), .B(n8409), .Z(n9462) );
  XOR U988 ( .A(in[681]), .B(in[1321]), .Z(n5405) );
  XNOR U989 ( .A(in[41]), .B(in[361]), .Z(n5404) );
  XNOR U990 ( .A(n5405), .B(n5404), .Z(n5406) );
  XOR U991 ( .A(in[1001]), .B(n5406), .Z(n6123) );
  XOR U992 ( .A(in[170]), .B(in[1450]), .Z(n5408) );
  XNOR U993 ( .A(in[1130]), .B(in[810]), .Z(n5407) );
  XNOR U994 ( .A(n5408), .B(n5407), .Z(n5409) );
  XOR U995 ( .A(in[490]), .B(n5409), .Z(n5660) );
  XNOR U996 ( .A(n6123), .B(n5660), .Z(n8784) );
  XNOR U997 ( .A(in[1386]), .B(n8784), .Z(n9459) );
  NAND U998 ( .A(n9462), .B(n9459), .Z(n5410) );
  XNOR U999 ( .A(n6227), .B(n5410), .Z(out[1030]) );
  XOR U1000 ( .A(n5412), .B(n5411), .Z(n8460) );
  XNOR U1001 ( .A(in[538]), .B(n8460), .Z(n6231) );
  XOR U1002 ( .A(in[1353]), .B(in[393]), .Z(n5414) );
  XNOR U1003 ( .A(in[713]), .B(in[73]), .Z(n5413) );
  XNOR U1004 ( .A(n5414), .B(n5413), .Z(n5415) );
  XOR U1005 ( .A(in[1033]), .B(n5415), .Z(n6321) );
  XOR U1006 ( .A(in[1482]), .B(in[522]), .Z(n5417) );
  XNOR U1007 ( .A(in[842]), .B(in[202]), .Z(n5416) );
  XNOR U1008 ( .A(n5417), .B(n5416), .Z(n5418) );
  XNOR U1009 ( .A(in[1162]), .B(n5418), .Z(n6026) );
  XNOR U1010 ( .A(n6321), .B(n6026), .Z(n8413) );
  XNOR U1011 ( .A(in[138]), .B(n8413), .Z(n9466) );
  XOR U1012 ( .A(in[811]), .B(in[491]), .Z(n5420) );
  XNOR U1013 ( .A(in[1451]), .B(in[1131]), .Z(n5419) );
  XNOR U1014 ( .A(n5420), .B(n5419), .Z(n5421) );
  XOR U1015 ( .A(in[171]), .B(n5421), .Z(n5673) );
  XOR U1016 ( .A(in[682]), .B(in[1322]), .Z(n5423) );
  XNOR U1017 ( .A(in[42]), .B(in[362]), .Z(n5422) );
  XNOR U1018 ( .A(n5423), .B(n5422), .Z(n5424) );
  XOR U1019 ( .A(in[1002]), .B(n5424), .Z(n6128) );
  XNOR U1020 ( .A(n5673), .B(n6128), .Z(n8787) );
  XNOR U1021 ( .A(in[1387]), .B(n8787), .Z(n9463) );
  NAND U1022 ( .A(n9466), .B(n9463), .Z(n5425) );
  XNOR U1023 ( .A(n6231), .B(n5425), .Z(out[1031]) );
  XOR U1024 ( .A(n5427), .B(n5426), .Z(n8464) );
  XNOR U1025 ( .A(in[539]), .B(n8464), .Z(n6236) );
  XOR U1026 ( .A(in[1483]), .B(in[523]), .Z(n5429) );
  XNOR U1027 ( .A(in[843]), .B(in[203]), .Z(n5428) );
  XNOR U1028 ( .A(n5429), .B(n5428), .Z(n5430) );
  XOR U1029 ( .A(in[1163]), .B(n5430), .Z(n6029) );
  XOR U1030 ( .A(in[1354]), .B(in[714]), .Z(n5432) );
  XNOR U1031 ( .A(in[74]), .B(in[394]), .Z(n5431) );
  XNOR U1032 ( .A(n5432), .B(n5431), .Z(n5433) );
  XNOR U1033 ( .A(in[1034]), .B(n5433), .Z(n6325) );
  XNOR U1034 ( .A(n6029), .B(n6325), .Z(n8417) );
  XNOR U1035 ( .A(n8417), .B(in[139]), .Z(n9470) );
  XOR U1036 ( .A(in[812]), .B(in[492]), .Z(n5435) );
  XNOR U1037 ( .A(in[1452]), .B(in[1132]), .Z(n5434) );
  XNOR U1038 ( .A(n5435), .B(n5434), .Z(n5436) );
  XOR U1039 ( .A(in[172]), .B(n5436), .Z(n5693) );
  XOR U1040 ( .A(in[683]), .B(in[1323]), .Z(n5438) );
  XNOR U1041 ( .A(in[43]), .B(in[363]), .Z(n5437) );
  XNOR U1042 ( .A(n5438), .B(n5437), .Z(n5439) );
  XOR U1043 ( .A(in[1003]), .B(n5439), .Z(n6132) );
  XNOR U1044 ( .A(n5693), .B(n6132), .Z(n8790) );
  XNOR U1045 ( .A(in[1388]), .B(n8790), .Z(n9467) );
  NAND U1046 ( .A(n9470), .B(n9467), .Z(n5440) );
  XNOR U1047 ( .A(n6236), .B(n5440), .Z(out[1032]) );
  XNOR U1048 ( .A(n5442), .B(n5441), .Z(n8468) );
  XNOR U1049 ( .A(in[540]), .B(n8468), .Z(n6240) );
  XOR U1050 ( .A(in[1355]), .B(in[715]), .Z(n5444) );
  XNOR U1051 ( .A(in[1035]), .B(in[395]), .Z(n5443) );
  XNOR U1052 ( .A(n5444), .B(n5443), .Z(n5445) );
  XOR U1053 ( .A(in[75]), .B(n5445), .Z(n6329) );
  XOR U1054 ( .A(in[1484]), .B(in[524]), .Z(n5447) );
  XNOR U1055 ( .A(in[844]), .B(in[204]), .Z(n5446) );
  XNOR U1056 ( .A(n5447), .B(n5446), .Z(n5448) );
  XNOR U1057 ( .A(in[1164]), .B(n5448), .Z(n6032) );
  XNOR U1058 ( .A(n6329), .B(n6032), .Z(n8421) );
  XNOR U1059 ( .A(in[140]), .B(n8421), .Z(n9474) );
  XOR U1060 ( .A(in[813]), .B(in[493]), .Z(n5450) );
  XNOR U1061 ( .A(in[1453]), .B(in[1133]), .Z(n5449) );
  XNOR U1062 ( .A(n5450), .B(n5449), .Z(n5451) );
  XOR U1063 ( .A(in[173]), .B(n5451), .Z(n5706) );
  XOR U1064 ( .A(in[1324]), .B(in[44]), .Z(n5453) );
  XNOR U1065 ( .A(in[684]), .B(in[364]), .Z(n5452) );
  XNOR U1066 ( .A(n5453), .B(n5452), .Z(n5454) );
  XOR U1067 ( .A(in[1004]), .B(n5454), .Z(n6135) );
  XNOR U1068 ( .A(n5706), .B(n6135), .Z(n8793) );
  XNOR U1069 ( .A(in[1389]), .B(n8793), .Z(n9471) );
  NAND U1070 ( .A(n9474), .B(n9471), .Z(n5455) );
  XNOR U1071 ( .A(n6240), .B(n5455), .Z(out[1033]) );
  XNOR U1072 ( .A(n5457), .B(n5456), .Z(n8476) );
  XNOR U1073 ( .A(in[541]), .B(n8476), .Z(n6244) );
  XOR U1074 ( .A(in[76]), .B(in[1036]), .Z(n5459) );
  XNOR U1075 ( .A(in[716]), .B(in[396]), .Z(n5458) );
  XNOR U1076 ( .A(n5459), .B(n5458), .Z(n5460) );
  XOR U1077 ( .A(in[1356]), .B(n5460), .Z(n6333) );
  XOR U1078 ( .A(in[1485]), .B(in[525]), .Z(n5462) );
  XNOR U1079 ( .A(in[845]), .B(in[205]), .Z(n5461) );
  XNOR U1080 ( .A(n5462), .B(n5461), .Z(n5463) );
  XNOR U1081 ( .A(in[1165]), .B(n5463), .Z(n6035) );
  XNOR U1082 ( .A(n6333), .B(n6035), .Z(n8425) );
  XNOR U1083 ( .A(in[141]), .B(n8425), .Z(n9482) );
  XOR U1084 ( .A(in[814]), .B(in[494]), .Z(n5465) );
  XNOR U1085 ( .A(in[1454]), .B(in[1134]), .Z(n5464) );
  XNOR U1086 ( .A(n5465), .B(n5464), .Z(n5466) );
  XOR U1087 ( .A(in[174]), .B(n5466), .Z(n5719) );
  XOR U1088 ( .A(in[1325]), .B(in[45]), .Z(n5468) );
  XNOR U1089 ( .A(in[685]), .B(in[365]), .Z(n5467) );
  XNOR U1090 ( .A(n5468), .B(n5467), .Z(n5469) );
  XOR U1091 ( .A(in[1005]), .B(n5469), .Z(n6139) );
  XNOR U1092 ( .A(n5719), .B(n6139), .Z(n8796) );
  XNOR U1093 ( .A(in[1390]), .B(n8796), .Z(n9479) );
  NAND U1094 ( .A(n9482), .B(n9479), .Z(n5470) );
  XNOR U1095 ( .A(n6244), .B(n5470), .Z(out[1034]) );
  XNOR U1096 ( .A(n5472), .B(n5471), .Z(n8480) );
  XNOR U1097 ( .A(in[542]), .B(n8480), .Z(n6248) );
  XOR U1098 ( .A(in[77]), .B(in[1037]), .Z(n5474) );
  XNOR U1099 ( .A(in[717]), .B(in[397]), .Z(n5473) );
  XNOR U1100 ( .A(n5474), .B(n5473), .Z(n5475) );
  XOR U1101 ( .A(in[1357]), .B(n5475), .Z(n6337) );
  XOR U1102 ( .A(in[1486]), .B(in[526]), .Z(n5477) );
  XNOR U1103 ( .A(in[846]), .B(in[206]), .Z(n5476) );
  XNOR U1104 ( .A(n5477), .B(n5476), .Z(n5478) );
  XNOR U1105 ( .A(in[1166]), .B(n5478), .Z(n6038) );
  XNOR U1106 ( .A(n6337), .B(n6038), .Z(n8433) );
  XNOR U1107 ( .A(in[142]), .B(n8433), .Z(n9486) );
  XOR U1108 ( .A(in[1326]), .B(in[46]), .Z(n5480) );
  XNOR U1109 ( .A(in[686]), .B(in[366]), .Z(n5479) );
  XNOR U1110 ( .A(n5480), .B(n5479), .Z(n5481) );
  XOR U1111 ( .A(in[1006]), .B(n5481), .Z(n6143) );
  XOR U1112 ( .A(in[815]), .B(in[495]), .Z(n5483) );
  XNOR U1113 ( .A(in[1455]), .B(in[1135]), .Z(n5482) );
  XNOR U1114 ( .A(n5483), .B(n5482), .Z(n5484) );
  XOR U1115 ( .A(in[175]), .B(n5484), .Z(n5732) );
  XNOR U1116 ( .A(n6143), .B(n5732), .Z(n8799) );
  XNOR U1117 ( .A(in[1391]), .B(n8799), .Z(n9483) );
  NAND U1118 ( .A(n9486), .B(n9483), .Z(n5485) );
  XNOR U1119 ( .A(n6248), .B(n5485), .Z(out[1035]) );
  XNOR U1120 ( .A(n5487), .B(n5486), .Z(n8484) );
  XNOR U1121 ( .A(in[543]), .B(n8484), .Z(n6252) );
  XOR U1122 ( .A(in[78]), .B(in[1038]), .Z(n5489) );
  XNOR U1123 ( .A(in[718]), .B(in[398]), .Z(n5488) );
  XNOR U1124 ( .A(n5489), .B(n5488), .Z(n5490) );
  XOR U1125 ( .A(in[1358]), .B(n5490), .Z(n6341) );
  XOR U1126 ( .A(in[1487]), .B(in[527]), .Z(n5492) );
  XNOR U1127 ( .A(in[847]), .B(in[207]), .Z(n5491) );
  XNOR U1128 ( .A(n5492), .B(n5491), .Z(n5493) );
  XNOR U1129 ( .A(in[1167]), .B(n5493), .Z(n6041) );
  XNOR U1130 ( .A(n6341), .B(n6041), .Z(n8437) );
  XNOR U1131 ( .A(in[143]), .B(n8437), .Z(n9490) );
  XOR U1132 ( .A(in[1327]), .B(in[47]), .Z(n5495) );
  XNOR U1133 ( .A(in[687]), .B(in[367]), .Z(n5494) );
  XNOR U1134 ( .A(n5495), .B(n5494), .Z(n5496) );
  XOR U1135 ( .A(in[1007]), .B(n5496), .Z(n6147) );
  XOR U1136 ( .A(in[816]), .B(in[496]), .Z(n5498) );
  XNOR U1137 ( .A(in[1456]), .B(in[1136]), .Z(n5497) );
  XNOR U1138 ( .A(n5498), .B(n5497), .Z(n5499) );
  XOR U1139 ( .A(in[176]), .B(n5499), .Z(n5747) );
  XNOR U1140 ( .A(n6147), .B(n5747), .Z(n8802) );
  XNOR U1141 ( .A(in[1392]), .B(n8802), .Z(n9487) );
  NAND U1142 ( .A(n9490), .B(n9487), .Z(n5500) );
  XNOR U1143 ( .A(n6252), .B(n5500), .Z(out[1036]) );
  XNOR U1144 ( .A(n5502), .B(n5501), .Z(n8488) );
  XNOR U1145 ( .A(in[544]), .B(n8488), .Z(n6256) );
  XOR U1146 ( .A(in[79]), .B(in[1039]), .Z(n5504) );
  XNOR U1147 ( .A(in[719]), .B(in[399]), .Z(n5503) );
  XNOR U1148 ( .A(n5504), .B(n5503), .Z(n5505) );
  XOR U1149 ( .A(in[1359]), .B(n5505), .Z(n6345) );
  XOR U1150 ( .A(in[1488]), .B(in[528]), .Z(n5507) );
  XNOR U1151 ( .A(in[848]), .B(in[208]), .Z(n5506) );
  XNOR U1152 ( .A(n5507), .B(n5506), .Z(n5508) );
  XNOR U1153 ( .A(in[1168]), .B(n5508), .Z(n6044) );
  XNOR U1154 ( .A(n6345), .B(n6044), .Z(n8441) );
  XNOR U1155 ( .A(in[144]), .B(n8441), .Z(n9494) );
  XOR U1156 ( .A(in[1328]), .B(in[48]), .Z(n5510) );
  XNOR U1157 ( .A(in[688]), .B(in[368]), .Z(n5509) );
  XNOR U1158 ( .A(n5510), .B(n5509), .Z(n5511) );
  XOR U1159 ( .A(in[1008]), .B(n5511), .Z(n6151) );
  XOR U1160 ( .A(in[817]), .B(in[497]), .Z(n5513) );
  XNOR U1161 ( .A(in[1457]), .B(in[1137]), .Z(n5512) );
  XNOR U1162 ( .A(n5513), .B(n5512), .Z(n5514) );
  XOR U1163 ( .A(in[177]), .B(n5514), .Z(n5762) );
  XNOR U1164 ( .A(n6151), .B(n5762), .Z(n8805) );
  XNOR U1165 ( .A(in[1393]), .B(n8805), .Z(n9491) );
  NAND U1166 ( .A(n9494), .B(n9491), .Z(n5515) );
  XNOR U1167 ( .A(n6256), .B(n5515), .Z(out[1037]) );
  XNOR U1168 ( .A(n5517), .B(n5516), .Z(n8492) );
  XNOR U1169 ( .A(in[545]), .B(n8492), .Z(n6260) );
  XOR U1170 ( .A(in[80]), .B(in[1040]), .Z(n5519) );
  XNOR U1171 ( .A(in[720]), .B(in[400]), .Z(n5518) );
  XNOR U1172 ( .A(n5519), .B(n5518), .Z(n5520) );
  XOR U1173 ( .A(in[1360]), .B(n5520), .Z(n6349) );
  XOR U1174 ( .A(in[1489]), .B(in[529]), .Z(n5522) );
  XNOR U1175 ( .A(in[849]), .B(in[209]), .Z(n5521) );
  XNOR U1176 ( .A(n5522), .B(n5521), .Z(n5523) );
  XNOR U1177 ( .A(in[1169]), .B(n5523), .Z(n6047) );
  XNOR U1178 ( .A(n6349), .B(n6047), .Z(n8445) );
  XNOR U1179 ( .A(in[145]), .B(n8445), .Z(n9498) );
  XOR U1180 ( .A(in[818]), .B(in[498]), .Z(n5525) );
  XNOR U1181 ( .A(in[1458]), .B(in[1138]), .Z(n5524) );
  XNOR U1182 ( .A(n5525), .B(n5524), .Z(n5526) );
  XOR U1183 ( .A(in[178]), .B(n5526), .Z(n5777) );
  XOR U1184 ( .A(in[1329]), .B(in[49]), .Z(n5528) );
  XNOR U1185 ( .A(in[689]), .B(in[369]), .Z(n5527) );
  XNOR U1186 ( .A(n5528), .B(n5527), .Z(n5529) );
  XOR U1187 ( .A(in[1009]), .B(n5529), .Z(n6156) );
  XNOR U1188 ( .A(n5777), .B(n6156), .Z(n8808) );
  XNOR U1189 ( .A(in[1394]), .B(n8808), .Z(n9495) );
  NAND U1190 ( .A(n9498), .B(n9495), .Z(n5530) );
  XNOR U1191 ( .A(n6260), .B(n5530), .Z(out[1038]) );
  XOR U1192 ( .A(n8496), .B(in[546]), .Z(n6264) );
  XOR U1193 ( .A(in[81]), .B(in[1041]), .Z(n5532) );
  XNOR U1194 ( .A(in[721]), .B(in[401]), .Z(n5531) );
  XNOR U1195 ( .A(n5532), .B(n5531), .Z(n5533) );
  XOR U1196 ( .A(in[1361]), .B(n5533), .Z(n6353) );
  XOR U1197 ( .A(in[1490]), .B(in[530]), .Z(n5535) );
  XNOR U1198 ( .A(in[850]), .B(in[210]), .Z(n5534) );
  XNOR U1199 ( .A(n5535), .B(n5534), .Z(n5536) );
  XNOR U1200 ( .A(in[1170]), .B(n5536), .Z(n6051) );
  XNOR U1201 ( .A(n6353), .B(n6051), .Z(n8449) );
  XNOR U1202 ( .A(in[146]), .B(n8449), .Z(n9502) );
  XOR U1203 ( .A(in[1330]), .B(in[50]), .Z(n5538) );
  XNOR U1204 ( .A(in[690]), .B(in[370]), .Z(n5537) );
  XNOR U1205 ( .A(n5538), .B(n5537), .Z(n5539) );
  XOR U1206 ( .A(in[1010]), .B(n5539), .Z(n6160) );
  XOR U1207 ( .A(in[819]), .B(in[499]), .Z(n5541) );
  XNOR U1208 ( .A(in[1459]), .B(in[1139]), .Z(n5540) );
  XNOR U1209 ( .A(n5541), .B(n5540), .Z(n5542) );
  XOR U1210 ( .A(in[179]), .B(n5542), .Z(n5792) );
  XNOR U1211 ( .A(n6160), .B(n5792), .Z(n8815) );
  XNOR U1212 ( .A(in[1395]), .B(n8815), .Z(n9499) );
  NAND U1213 ( .A(n9502), .B(n9499), .Z(n5543) );
  XNOR U1214 ( .A(n6264), .B(n5543), .Z(out[1039]) );
  XOR U1215 ( .A(in[1342]), .B(in[62]), .Z(n5545) );
  XNOR U1216 ( .A(in[702]), .B(in[382]), .Z(n5544) );
  XNOR U1217 ( .A(n5545), .B(n5544), .Z(n5546) );
  XOR U1218 ( .A(in[1022]), .B(n5546), .Z(n5714) );
  XNOR U1219 ( .A(n5547), .B(n5714), .Z(n8411) );
  XNOR U1220 ( .A(in[638]), .B(n8411), .Z(n7364) );
  XOR U1221 ( .A(n5549), .B(n5548), .Z(n8508) );
  XNOR U1222 ( .A(in[229]), .B(n8508), .Z(n7680) );
  XOR U1223 ( .A(in[1513]), .B(in[553]), .Z(n5551) );
  XNOR U1224 ( .A(in[873]), .B(in[233]), .Z(n5550) );
  XNOR U1225 ( .A(n5551), .B(n5550), .Z(n5552) );
  XOR U1226 ( .A(in[1193]), .B(n5552), .Z(n6127) );
  XNOR U1227 ( .A(n5553), .B(n6127), .Z(n8549) );
  XNOR U1228 ( .A(in[1449]), .B(n8549), .Z(n7677) );
  NAND U1229 ( .A(n7680), .B(n7677), .Z(n5554) );
  XNOR U1230 ( .A(n7364), .B(n5554), .Z(out[103]) );
  XOR U1231 ( .A(n8500), .B(in[547]), .Z(n6268) );
  XOR U1232 ( .A(in[1042]), .B(in[402]), .Z(n5556) );
  XNOR U1233 ( .A(in[722]), .B(in[82]), .Z(n5555) );
  XNOR U1234 ( .A(n5556), .B(n5555), .Z(n5557) );
  XOR U1235 ( .A(in[1362]), .B(n5557), .Z(n6358) );
  XOR U1236 ( .A(in[851]), .B(in[1171]), .Z(n5559) );
  XNOR U1237 ( .A(in[1491]), .B(in[211]), .Z(n5558) );
  XNOR U1238 ( .A(n5559), .B(n5558), .Z(n5560) );
  XNOR U1239 ( .A(in[531]), .B(n5560), .Z(n6054) );
  XNOR U1240 ( .A(n6358), .B(n6054), .Z(n8453) );
  XNOR U1241 ( .A(in[147]), .B(n8453), .Z(n9506) );
  XOR U1242 ( .A(in[1331]), .B(in[51]), .Z(n5562) );
  XNOR U1243 ( .A(in[691]), .B(in[371]), .Z(n5561) );
  XNOR U1244 ( .A(n5562), .B(n5561), .Z(n5563) );
  XOR U1245 ( .A(in[1011]), .B(n5563), .Z(n6164) );
  XOR U1246 ( .A(in[820]), .B(in[500]), .Z(n5565) );
  XNOR U1247 ( .A(in[1460]), .B(in[1140]), .Z(n5564) );
  XNOR U1248 ( .A(n5565), .B(n5564), .Z(n5566) );
  XOR U1249 ( .A(in[180]), .B(n5566), .Z(n5807) );
  XNOR U1250 ( .A(n6164), .B(n5807), .Z(n8818) );
  XNOR U1251 ( .A(in[1396]), .B(n8818), .Z(n9503) );
  NAND U1252 ( .A(n9506), .B(n9503), .Z(n5567) );
  XNOR U1253 ( .A(n6268), .B(n5567), .Z(out[1040]) );
  XOR U1254 ( .A(n8504), .B(in[548]), .Z(n6272) );
  XOR U1255 ( .A(in[83]), .B(in[1043]), .Z(n5569) );
  XNOR U1256 ( .A(in[723]), .B(in[403]), .Z(n5568) );
  XNOR U1257 ( .A(n5569), .B(n5568), .Z(n5570) );
  XOR U1258 ( .A(in[1363]), .B(n5570), .Z(n6362) );
  XOR U1259 ( .A(in[852]), .B(in[1172]), .Z(n5572) );
  XNOR U1260 ( .A(in[1492]), .B(in[212]), .Z(n5571) );
  XNOR U1261 ( .A(n5572), .B(n5571), .Z(n5573) );
  XNOR U1262 ( .A(in[532]), .B(n5573), .Z(n6057) );
  XNOR U1263 ( .A(n6362), .B(n6057), .Z(n8457) );
  XNOR U1264 ( .A(in[148]), .B(n8457), .Z(n9510) );
  XOR U1265 ( .A(in[821]), .B(in[501]), .Z(n5575) );
  XNOR U1266 ( .A(in[1461]), .B(in[1141]), .Z(n5574) );
  XNOR U1267 ( .A(n5575), .B(n5574), .Z(n5576) );
  XOR U1268 ( .A(in[181]), .B(n5576), .Z(n5822) );
  XOR U1269 ( .A(in[1332]), .B(in[52]), .Z(n5578) );
  XNOR U1270 ( .A(in[692]), .B(in[372]), .Z(n5577) );
  XNOR U1271 ( .A(n5578), .B(n5577), .Z(n5579) );
  XOR U1272 ( .A(in[1012]), .B(n5579), .Z(n6168) );
  XNOR U1273 ( .A(n5822), .B(n6168), .Z(n8821) );
  XNOR U1274 ( .A(in[1397]), .B(n8821), .Z(n9507) );
  NAND U1275 ( .A(n9510), .B(n9507), .Z(n5580) );
  XNOR U1276 ( .A(n6272), .B(n5580), .Z(out[1041]) );
  XOR U1277 ( .A(n8508), .B(in[549]), .Z(n6277) );
  XOR U1278 ( .A(in[853]), .B(in[1173]), .Z(n5582) );
  XNOR U1279 ( .A(in[1493]), .B(in[213]), .Z(n5581) );
  XNOR U1280 ( .A(n5582), .B(n5581), .Z(n5583) );
  XNOR U1281 ( .A(in[533]), .B(n5583), .Z(n6060) );
  XNOR U1282 ( .A(n5584), .B(n6060), .Z(n8461) );
  XNOR U1283 ( .A(in[149]), .B(n8461), .Z(n9514) );
  XOR U1284 ( .A(in[822]), .B(in[502]), .Z(n5586) );
  XNOR U1285 ( .A(in[1462]), .B(in[1142]), .Z(n5585) );
  XNOR U1286 ( .A(n5586), .B(n5585), .Z(n5587) );
  XOR U1287 ( .A(in[182]), .B(n5587), .Z(n5836) );
  XOR U1288 ( .A(in[1333]), .B(in[53]), .Z(n5589) );
  XNOR U1289 ( .A(in[693]), .B(in[373]), .Z(n5588) );
  XNOR U1290 ( .A(n5589), .B(n5588), .Z(n5590) );
  XOR U1291 ( .A(in[1013]), .B(n5590), .Z(n6172) );
  XNOR U1292 ( .A(n5836), .B(n6172), .Z(n8824) );
  XNOR U1293 ( .A(in[1398]), .B(n8824), .Z(n9511) );
  NAND U1294 ( .A(n9514), .B(n9511), .Z(n5591) );
  XNOR U1295 ( .A(n6277), .B(n5591), .Z(out[1042]) );
  XNOR U1296 ( .A(n5593), .B(n5592), .Z(n8512) );
  XNOR U1297 ( .A(in[550]), .B(n8512), .Z(n6281) );
  XOR U1298 ( .A(in[854]), .B(in[1174]), .Z(n5595) );
  XNOR U1299 ( .A(in[1494]), .B(in[214]), .Z(n5594) );
  XNOR U1300 ( .A(n5595), .B(n5594), .Z(n5596) );
  XNOR U1301 ( .A(in[534]), .B(n5596), .Z(n6063) );
  XNOR U1302 ( .A(n5597), .B(n6063), .Z(n8465) );
  XNOR U1303 ( .A(in[150]), .B(n8465), .Z(n9518) );
  XOR U1304 ( .A(in[823]), .B(in[503]), .Z(n5599) );
  XNOR U1305 ( .A(in[1463]), .B(in[1143]), .Z(n5598) );
  XNOR U1306 ( .A(n5599), .B(n5598), .Z(n5600) );
  XOR U1307 ( .A(in[183]), .B(n5600), .Z(n5847) );
  XOR U1308 ( .A(in[1334]), .B(in[54]), .Z(n5602) );
  XNOR U1309 ( .A(in[694]), .B(in[374]), .Z(n5601) );
  XNOR U1310 ( .A(n5602), .B(n5601), .Z(n5603) );
  XOR U1311 ( .A(in[1014]), .B(n5603), .Z(n6176) );
  XNOR U1312 ( .A(n5847), .B(n6176), .Z(n8827) );
  XNOR U1313 ( .A(in[1399]), .B(n8827), .Z(n9515) );
  NAND U1314 ( .A(n9518), .B(n9515), .Z(n5604) );
  XNOR U1315 ( .A(n6281), .B(n5604), .Z(out[1043]) );
  XNOR U1316 ( .A(n5606), .B(n5605), .Z(n8520) );
  XNOR U1317 ( .A(in[551]), .B(n8520), .Z(n6285) );
  XOR U1318 ( .A(in[855]), .B(in[1175]), .Z(n5608) );
  XNOR U1319 ( .A(in[1495]), .B(in[215]), .Z(n5607) );
  XNOR U1320 ( .A(n5608), .B(n5607), .Z(n5609) );
  XNOR U1321 ( .A(in[535]), .B(n5609), .Z(n6066) );
  XNOR U1322 ( .A(n5610), .B(n6066), .Z(n8469) );
  XNOR U1323 ( .A(in[151]), .B(n8469), .Z(n9526) );
  XOR U1324 ( .A(in[1335]), .B(in[55]), .Z(n5612) );
  XNOR U1325 ( .A(in[695]), .B(in[375]), .Z(n5611) );
  XNOR U1326 ( .A(n5612), .B(n5611), .Z(n5613) );
  XOR U1327 ( .A(in[1015]), .B(n5613), .Z(n6180) );
  XOR U1328 ( .A(in[824]), .B(in[504]), .Z(n5615) );
  XNOR U1329 ( .A(in[1464]), .B(in[1144]), .Z(n5614) );
  XNOR U1330 ( .A(n5615), .B(n5614), .Z(n5616) );
  XOR U1331 ( .A(in[184]), .B(n5616), .Z(n5852) );
  XNOR U1332 ( .A(n6180), .B(n5852), .Z(n8830) );
  XNOR U1333 ( .A(in[1400]), .B(n8830), .Z(n9523) );
  NAND U1334 ( .A(n9526), .B(n9523), .Z(n5617) );
  XNOR U1335 ( .A(n6285), .B(n5617), .Z(out[1044]) );
  XNOR U1336 ( .A(n5619), .B(n5618), .Z(n8524) );
  XNOR U1337 ( .A(in[552]), .B(n8524), .Z(n6289) );
  XOR U1338 ( .A(in[856]), .B(in[1176]), .Z(n5621) );
  XNOR U1339 ( .A(in[1496]), .B(in[216]), .Z(n5620) );
  XNOR U1340 ( .A(n5621), .B(n5620), .Z(n5622) );
  XNOR U1341 ( .A(in[536]), .B(n5622), .Z(n6069) );
  XNOR U1342 ( .A(n5623), .B(n6069), .Z(n8477) );
  XNOR U1343 ( .A(in[152]), .B(n8477), .Z(n9530) );
  XOR U1344 ( .A(in[1336]), .B(in[56]), .Z(n5625) );
  XNOR U1345 ( .A(in[696]), .B(in[376]), .Z(n5624) );
  XNOR U1346 ( .A(n5625), .B(n5624), .Z(n5626) );
  XOR U1347 ( .A(in[1016]), .B(n5626), .Z(n6184) );
  XOR U1348 ( .A(in[825]), .B(in[505]), .Z(n5628) );
  XNOR U1349 ( .A(in[1465]), .B(in[1145]), .Z(n5627) );
  XNOR U1350 ( .A(n5628), .B(n5627), .Z(n5629) );
  XOR U1351 ( .A(in[185]), .B(n5629), .Z(n5863) );
  XNOR U1352 ( .A(n6184), .B(n5863), .Z(n8833) );
  XNOR U1353 ( .A(in[1401]), .B(n8833), .Z(n9527) );
  NAND U1354 ( .A(n9530), .B(n9527), .Z(n5630) );
  XNOR U1355 ( .A(n6289), .B(n5630), .Z(out[1045]) );
  XNOR U1356 ( .A(n5632), .B(n5631), .Z(n8528) );
  XNOR U1357 ( .A(in[553]), .B(n8528), .Z(n6293) );
  XOR U1358 ( .A(in[857]), .B(in[1177]), .Z(n5634) );
  XNOR U1359 ( .A(in[1497]), .B(in[217]), .Z(n5633) );
  XNOR U1360 ( .A(n5634), .B(n5633), .Z(n5635) );
  XNOR U1361 ( .A(in[537]), .B(n5635), .Z(n6072) );
  XNOR U1362 ( .A(n5636), .B(n6072), .Z(n8481) );
  XNOR U1363 ( .A(in[153]), .B(n8481), .Z(n9534) );
  XOR U1364 ( .A(in[1337]), .B(in[57]), .Z(n5638) );
  XNOR U1365 ( .A(in[697]), .B(in[377]), .Z(n5637) );
  XNOR U1366 ( .A(n5638), .B(n5637), .Z(n5639) );
  XOR U1367 ( .A(in[1017]), .B(n5639), .Z(n6188) );
  XOR U1368 ( .A(in[826]), .B(in[506]), .Z(n5641) );
  XNOR U1369 ( .A(in[1466]), .B(in[1146]), .Z(n5640) );
  XNOR U1370 ( .A(n5641), .B(n5640), .Z(n5642) );
  XOR U1371 ( .A(in[186]), .B(n5642), .Z(n5874) );
  XNOR U1372 ( .A(n6188), .B(n5874), .Z(n8836) );
  XNOR U1373 ( .A(in[1402]), .B(n8836), .Z(n9531) );
  NAND U1374 ( .A(n9534), .B(n9531), .Z(n5643) );
  XNOR U1375 ( .A(n6293), .B(n5643), .Z(out[1046]) );
  XNOR U1376 ( .A(n5645), .B(n5644), .Z(n8532) );
  XNOR U1377 ( .A(in[554]), .B(n8532), .Z(n6297) );
  XOR U1378 ( .A(in[858]), .B(in[1178]), .Z(n5647) );
  XNOR U1379 ( .A(in[1498]), .B(in[218]), .Z(n5646) );
  XNOR U1380 ( .A(n5647), .B(n5646), .Z(n5648) );
  XNOR U1381 ( .A(in[538]), .B(n5648), .Z(n6075) );
  XNOR U1382 ( .A(n5649), .B(n6075), .Z(n8485) );
  XNOR U1383 ( .A(in[154]), .B(n8485), .Z(n9538) );
  XOR U1384 ( .A(in[1338]), .B(in[58]), .Z(n5651) );
  XNOR U1385 ( .A(in[698]), .B(in[378]), .Z(n5650) );
  XNOR U1386 ( .A(n5651), .B(n5650), .Z(n5652) );
  XOR U1387 ( .A(in[1018]), .B(n5652), .Z(n6192) );
  XOR U1388 ( .A(in[827]), .B(in[507]), .Z(n5654) );
  XNOR U1389 ( .A(in[1467]), .B(in[1147]), .Z(n5653) );
  XNOR U1390 ( .A(n5654), .B(n5653), .Z(n5655) );
  XOR U1391 ( .A(in[187]), .B(n5655), .Z(n5879) );
  XNOR U1392 ( .A(n6192), .B(n5879), .Z(n8839) );
  XNOR U1393 ( .A(in[1403]), .B(n8839), .Z(n9535) );
  NAND U1394 ( .A(n9538), .B(n9535), .Z(n5656) );
  XNOR U1395 ( .A(n6297), .B(n5656), .Z(out[1047]) );
  XOR U1396 ( .A(in[1579]), .B(in[619]), .Z(n5658) );
  XNOR U1397 ( .A(in[939]), .B(in[299]), .Z(n5657) );
  XNOR U1398 ( .A(n5658), .B(n5657), .Z(n5659) );
  XOR U1399 ( .A(in[1259]), .B(n5659), .Z(n6201) );
  XNOR U1400 ( .A(n5660), .B(n6201), .Z(n8536) );
  XNOR U1401 ( .A(in[555]), .B(n8536), .Z(n6301) );
  XOR U1402 ( .A(in[859]), .B(in[1179]), .Z(n5662) );
  XNOR U1403 ( .A(in[1499]), .B(in[219]), .Z(n5661) );
  XNOR U1404 ( .A(n5662), .B(n5661), .Z(n5663) );
  XNOR U1405 ( .A(in[539]), .B(n5663), .Z(n6078) );
  XNOR U1406 ( .A(n5664), .B(n6078), .Z(n8489) );
  XNOR U1407 ( .A(in[155]), .B(n8489), .Z(n9542) );
  XOR U1408 ( .A(in[828]), .B(in[508]), .Z(n5666) );
  XNOR U1409 ( .A(in[1468]), .B(in[1148]), .Z(n5665) );
  XNOR U1410 ( .A(n5666), .B(n5665), .Z(n5667) );
  XOR U1411 ( .A(in[188]), .B(n5667), .Z(n5884) );
  XNOR U1412 ( .A(n5668), .B(n5884), .Z(n8842) );
  XNOR U1413 ( .A(in[1404]), .B(n8842), .Z(n9539) );
  NAND U1414 ( .A(n9542), .B(n9539), .Z(n5669) );
  XNOR U1415 ( .A(n6301), .B(n5669), .Z(out[1048]) );
  XOR U1416 ( .A(in[1580]), .B(in[620]), .Z(n5671) );
  XNOR U1417 ( .A(in[940]), .B(in[300]), .Z(n5670) );
  XNOR U1418 ( .A(n5671), .B(n5670), .Z(n5672) );
  XOR U1419 ( .A(in[1260]), .B(n5672), .Z(n6205) );
  XNOR U1420 ( .A(n5673), .B(n6205), .Z(n8540) );
  XNOR U1421 ( .A(in[556]), .B(n8540), .Z(n6305) );
  XOR U1422 ( .A(in[860]), .B(in[1180]), .Z(n5675) );
  XNOR U1423 ( .A(in[1500]), .B(in[220]), .Z(n5674) );
  XNOR U1424 ( .A(n5675), .B(n5674), .Z(n5676) );
  XNOR U1425 ( .A(in[540]), .B(n5676), .Z(n6082) );
  XNOR U1426 ( .A(n5677), .B(n6082), .Z(n8493) );
  XNOR U1427 ( .A(in[156]), .B(n8493), .Z(n9546) );
  XNOR U1428 ( .A(n5679), .B(n5678), .Z(n8849) );
  XNOR U1429 ( .A(in[1405]), .B(n8849), .Z(n9543) );
  NAND U1430 ( .A(n9546), .B(n9543), .Z(n5680) );
  XNOR U1431 ( .A(n6305), .B(n5680), .Z(out[1049]) );
  XOR U1432 ( .A(in[1343]), .B(in[63]), .Z(n5682) );
  XNOR U1433 ( .A(in[703]), .B(in[383]), .Z(n5681) );
  XNOR U1434 ( .A(n5682), .B(n5681), .Z(n5683) );
  XOR U1435 ( .A(in[1023]), .B(n5683), .Z(n5727) );
  XNOR U1436 ( .A(n5684), .B(n5727), .Z(n8415) );
  XNOR U1437 ( .A(in[639]), .B(n8415), .Z(n7366) );
  XOR U1438 ( .A(in[230]), .B(n8512), .Z(n7696) );
  XOR U1439 ( .A(in[874]), .B(in[1194]), .Z(n5686) );
  XNOR U1440 ( .A(in[1514]), .B(in[234]), .Z(n5685) );
  XNOR U1441 ( .A(n5686), .B(n5685), .Z(n5687) );
  XOR U1442 ( .A(in[554]), .B(n5687), .Z(n6131) );
  XNOR U1443 ( .A(n5688), .B(n6131), .Z(n8553) );
  XNOR U1444 ( .A(in[1450]), .B(n8553), .Z(n7693) );
  NAND U1445 ( .A(n7696), .B(n7693), .Z(n5689) );
  XNOR U1446 ( .A(n7366), .B(n5689), .Z(out[104]) );
  XOR U1447 ( .A(in[1581]), .B(in[621]), .Z(n5691) );
  XNOR U1448 ( .A(in[941]), .B(in[301]), .Z(n5690) );
  XNOR U1449 ( .A(n5691), .B(n5690), .Z(n5692) );
  XOR U1450 ( .A(in[1261]), .B(n5692), .Z(n6209) );
  XNOR U1451 ( .A(n5693), .B(n6209), .Z(n8544) );
  XNOR U1452 ( .A(in[557]), .B(n8544), .Z(n6309) );
  XOR U1453 ( .A(in[861]), .B(in[1181]), .Z(n5695) );
  XNOR U1454 ( .A(in[1501]), .B(in[221]), .Z(n5694) );
  XNOR U1455 ( .A(n5695), .B(n5694), .Z(n5696) );
  XNOR U1456 ( .A(in[541]), .B(n5696), .Z(n6085) );
  XNOR U1457 ( .A(n5697), .B(n6085), .Z(n8497) );
  XNOR U1458 ( .A(in[157]), .B(n8497), .Z(n9550) );
  XOR U1459 ( .A(in[830]), .B(in[510]), .Z(n5699) );
  XNOR U1460 ( .A(in[1470]), .B(in[1150]), .Z(n5698) );
  XNOR U1461 ( .A(n5699), .B(n5698), .Z(n5700) );
  XOR U1462 ( .A(in[190]), .B(n5700), .Z(n5890) );
  XNOR U1463 ( .A(n5701), .B(n5890), .Z(n8852) );
  XNOR U1464 ( .A(in[1406]), .B(n8852), .Z(n9547) );
  NAND U1465 ( .A(n9550), .B(n9547), .Z(n5702) );
  XNOR U1466 ( .A(n6309), .B(n5702), .Z(out[1050]) );
  XOR U1467 ( .A(in[1582]), .B(in[622]), .Z(n5704) );
  XNOR U1468 ( .A(in[942]), .B(in[302]), .Z(n5703) );
  XNOR U1469 ( .A(n5704), .B(n5703), .Z(n5705) );
  XOR U1470 ( .A(in[1262]), .B(n5705), .Z(n6213) );
  XNOR U1471 ( .A(n5706), .B(n6213), .Z(n8548) );
  XNOR U1472 ( .A(in[558]), .B(n8548), .Z(n6313) );
  XOR U1473 ( .A(in[862]), .B(in[1182]), .Z(n5708) );
  XNOR U1474 ( .A(in[1502]), .B(in[222]), .Z(n5707) );
  XNOR U1475 ( .A(n5708), .B(n5707), .Z(n5709) );
  XNOR U1476 ( .A(in[542]), .B(n5709), .Z(n6088) );
  XNOR U1477 ( .A(n5710), .B(n6088), .Z(n8501) );
  XNOR U1478 ( .A(in[158]), .B(n8501), .Z(n9554) );
  XOR U1479 ( .A(in[831]), .B(in[511]), .Z(n5712) );
  XNOR U1480 ( .A(in[1471]), .B(in[1151]), .Z(n5711) );
  XNOR U1481 ( .A(n5712), .B(n5711), .Z(n5713) );
  XOR U1482 ( .A(in[191]), .B(n5713), .Z(n5895) );
  XNOR U1483 ( .A(n5714), .B(n5895), .Z(n8855) );
  XNOR U1484 ( .A(in[1407]), .B(n8855), .Z(n9551) );
  NAND U1485 ( .A(n9554), .B(n9551), .Z(n5715) );
  XNOR U1486 ( .A(n6313), .B(n5715), .Z(out[1051]) );
  XOR U1487 ( .A(in[1583]), .B(in[623]), .Z(n5717) );
  XNOR U1488 ( .A(in[943]), .B(in[303]), .Z(n5716) );
  XNOR U1489 ( .A(n5717), .B(n5716), .Z(n5718) );
  XOR U1490 ( .A(in[1263]), .B(n5718), .Z(n6217) );
  XNOR U1491 ( .A(n5719), .B(n6217), .Z(n8552) );
  XNOR U1492 ( .A(in[559]), .B(n8552), .Z(n6318) );
  XOR U1493 ( .A(in[863]), .B(in[1183]), .Z(n5721) );
  XNOR U1494 ( .A(in[1503]), .B(in[223]), .Z(n5720) );
  XNOR U1495 ( .A(n5721), .B(n5720), .Z(n5722) );
  XNOR U1496 ( .A(in[543]), .B(n5722), .Z(n6091) );
  XNOR U1497 ( .A(n5723), .B(n6091), .Z(n8505) );
  XNOR U1498 ( .A(in[159]), .B(n8505), .Z(n9558) );
  XOR U1499 ( .A(in[768]), .B(in[1088]), .Z(n5725) );
  XNOR U1500 ( .A(in[448]), .B(in[1408]), .Z(n5724) );
  XNOR U1501 ( .A(n5725), .B(n5724), .Z(n5726) );
  XOR U1502 ( .A(in[128]), .B(n5726), .Z(n5903) );
  XNOR U1503 ( .A(n5727), .B(n5903), .Z(n8858) );
  XNOR U1504 ( .A(in[1344]), .B(n8858), .Z(n9555) );
  NAND U1505 ( .A(n9558), .B(n9555), .Z(n5728) );
  XNOR U1506 ( .A(n6318), .B(n5728), .Z(out[1052]) );
  XOR U1507 ( .A(in[1584]), .B(in[624]), .Z(n5730) );
  XNOR U1508 ( .A(in[944]), .B(in[304]), .Z(n5729) );
  XNOR U1509 ( .A(n5730), .B(n5729), .Z(n5731) );
  XOR U1510 ( .A(in[1264]), .B(n5731), .Z(n6221) );
  XNOR U1511 ( .A(n5732), .B(n6221), .Z(n8556) );
  XNOR U1512 ( .A(in[560]), .B(n8556), .Z(n6322) );
  XOR U1513 ( .A(in[224]), .B(in[864]), .Z(n5734) );
  XNOR U1514 ( .A(in[1184]), .B(in[1504]), .Z(n5733) );
  XNOR U1515 ( .A(n5734), .B(n5733), .Z(n5735) );
  XNOR U1516 ( .A(in[544]), .B(n5735), .Z(n6094) );
  XNOR U1517 ( .A(n5736), .B(n6094), .Z(n8509) );
  XNOR U1518 ( .A(in[160]), .B(n8509), .Z(n9562) );
  XOR U1519 ( .A(in[1280]), .B(in[640]), .Z(n5738) );
  XNOR U1520 ( .A(in[960]), .B(in[320]), .Z(n5737) );
  XNOR U1521 ( .A(n5738), .B(n5737), .Z(n5739) );
  XOR U1522 ( .A(in[0]), .B(n5739), .Z(n5830) );
  XOR U1523 ( .A(in[769]), .B(in[1089]), .Z(n5741) );
  XNOR U1524 ( .A(in[449]), .B(in[1409]), .Z(n5740) );
  XNOR U1525 ( .A(n5741), .B(n5740), .Z(n5742) );
  XOR U1526 ( .A(in[129]), .B(n5742), .Z(n5908) );
  XNOR U1527 ( .A(n5830), .B(n5908), .Z(n8861) );
  XNOR U1528 ( .A(in[1345]), .B(n8861), .Z(n9559) );
  NAND U1529 ( .A(n9562), .B(n9559), .Z(n5743) );
  XNOR U1530 ( .A(n6322), .B(n5743), .Z(out[1053]) );
  XOR U1531 ( .A(in[1585]), .B(in[625]), .Z(n5745) );
  XNOR U1532 ( .A(in[945]), .B(in[305]), .Z(n5744) );
  XNOR U1533 ( .A(n5745), .B(n5744), .Z(n5746) );
  XOR U1534 ( .A(in[1265]), .B(n5746), .Z(n6225) );
  XNOR U1535 ( .A(n5747), .B(n6225), .Z(n8564) );
  XNOR U1536 ( .A(in[561]), .B(n8564), .Z(n6326) );
  XOR U1537 ( .A(in[225]), .B(in[865]), .Z(n5749) );
  XNOR U1538 ( .A(in[1185]), .B(in[1505]), .Z(n5748) );
  XNOR U1539 ( .A(n5749), .B(n5748), .Z(n5750) );
  XNOR U1540 ( .A(in[545]), .B(n5750), .Z(n6097) );
  XNOR U1541 ( .A(n5751), .B(n6097), .Z(n8513) );
  XNOR U1542 ( .A(in[161]), .B(n8513), .Z(n9570) );
  XOR U1543 ( .A(in[1]), .B(in[641]), .Z(n5753) );
  XNOR U1544 ( .A(in[961]), .B(in[321]), .Z(n5752) );
  XNOR U1545 ( .A(n5753), .B(n5752), .Z(n5754) );
  XOR U1546 ( .A(in[1281]), .B(n5754), .Z(n5897) );
  XOR U1547 ( .A(in[1090]), .B(in[450]), .Z(n5756) );
  XNOR U1548 ( .A(in[130]), .B(in[770]), .Z(n5755) );
  XNOR U1549 ( .A(n5756), .B(n5755), .Z(n5757) );
  XOR U1550 ( .A(in[1410]), .B(n5757), .Z(n5913) );
  XNOR U1551 ( .A(n5897), .B(n5913), .Z(n8864) );
  XNOR U1552 ( .A(in[1346]), .B(n8864), .Z(n9567) );
  NAND U1553 ( .A(n9570), .B(n9567), .Z(n5758) );
  XNOR U1554 ( .A(n6326), .B(n5758), .Z(out[1054]) );
  XOR U1555 ( .A(in[1586]), .B(in[626]), .Z(n5760) );
  XNOR U1556 ( .A(in[946]), .B(in[306]), .Z(n5759) );
  XNOR U1557 ( .A(n5760), .B(n5759), .Z(n5761) );
  XOR U1558 ( .A(in[1266]), .B(n5761), .Z(n6229) );
  XNOR U1559 ( .A(n5762), .B(n6229), .Z(n8568) );
  XNOR U1560 ( .A(in[562]), .B(n8568), .Z(n6330) );
  XOR U1561 ( .A(in[1186]), .B(in[1506]), .Z(n5764) );
  XNOR U1562 ( .A(in[546]), .B(in[866]), .Z(n5763) );
  XNOR U1563 ( .A(n5764), .B(n5763), .Z(n5765) );
  XNOR U1564 ( .A(in[226]), .B(n5765), .Z(n6100) );
  XNOR U1565 ( .A(n5766), .B(n6100), .Z(n8521) );
  XNOR U1566 ( .A(in[162]), .B(n8521), .Z(n9574) );
  XOR U1567 ( .A(in[771]), .B(in[1091]), .Z(n5768) );
  XNOR U1568 ( .A(in[451]), .B(in[1411]), .Z(n5767) );
  XNOR U1569 ( .A(n5768), .B(n5767), .Z(n5769) );
  XOR U1570 ( .A(in[131]), .B(n5769), .Z(n5918) );
  XOR U1571 ( .A(in[2]), .B(in[642]), .Z(n5771) );
  XNOR U1572 ( .A(in[962]), .B(in[322]), .Z(n5770) );
  XNOR U1573 ( .A(n5771), .B(n5770), .Z(n5772) );
  XOR U1574 ( .A(in[1282]), .B(n5772), .Z(n5950) );
  XNOR U1575 ( .A(n5918), .B(n5950), .Z(n8867) );
  XNOR U1576 ( .A(in[1347]), .B(n8867), .Z(n9571) );
  NAND U1577 ( .A(n9574), .B(n9571), .Z(n5773) );
  XNOR U1578 ( .A(n6330), .B(n5773), .Z(out[1055]) );
  XOR U1579 ( .A(in[1587]), .B(in[627]), .Z(n5775) );
  XNOR U1580 ( .A(in[947]), .B(in[307]), .Z(n5774) );
  XNOR U1581 ( .A(n5775), .B(n5774), .Z(n5776) );
  XOR U1582 ( .A(in[1267]), .B(n5776), .Z(n6234) );
  XNOR U1583 ( .A(n5777), .B(n6234), .Z(n8572) );
  XNOR U1584 ( .A(in[563]), .B(n8572), .Z(n6334) );
  XOR U1585 ( .A(in[1187]), .B(in[1507]), .Z(n5779) );
  XNOR U1586 ( .A(in[547]), .B(in[867]), .Z(n5778) );
  XNOR U1587 ( .A(n5779), .B(n5778), .Z(n5780) );
  XNOR U1588 ( .A(in[227]), .B(n5780), .Z(n6103) );
  XNOR U1589 ( .A(n5781), .B(n6103), .Z(n8525) );
  XNOR U1590 ( .A(in[163]), .B(n8525), .Z(n9578) );
  XOR U1591 ( .A(in[323]), .B(in[643]), .Z(n5783) );
  XNOR U1592 ( .A(in[963]), .B(in[3]), .Z(n5782) );
  XNOR U1593 ( .A(n5783), .B(n5782), .Z(n5784) );
  XOR U1594 ( .A(in[1283]), .B(n5784), .Z(n5996) );
  XOR U1595 ( .A(in[772]), .B(in[1092]), .Z(n5786) );
  XNOR U1596 ( .A(in[452]), .B(in[1412]), .Z(n5785) );
  XNOR U1597 ( .A(n5786), .B(n5785), .Z(n5787) );
  XOR U1598 ( .A(in[132]), .B(n5787), .Z(n5923) );
  XNOR U1599 ( .A(n5996), .B(n5923), .Z(n8870) );
  XNOR U1600 ( .A(in[1348]), .B(n8870), .Z(n9575) );
  NAND U1601 ( .A(n9578), .B(n9575), .Z(n5788) );
  XNOR U1602 ( .A(n6334), .B(n5788), .Z(out[1056]) );
  XOR U1603 ( .A(in[1588]), .B(in[628]), .Z(n5790) );
  XNOR U1604 ( .A(in[948]), .B(in[308]), .Z(n5789) );
  XNOR U1605 ( .A(n5790), .B(n5789), .Z(n5791) );
  XOR U1606 ( .A(in[1268]), .B(n5791), .Z(n6238) );
  XNOR U1607 ( .A(n5792), .B(n6238), .Z(n8576) );
  XNOR U1608 ( .A(in[564]), .B(n8576), .Z(n6338) );
  XOR U1609 ( .A(in[1188]), .B(in[1508]), .Z(n5794) );
  XNOR U1610 ( .A(in[548]), .B(in[868]), .Z(n5793) );
  XNOR U1611 ( .A(n5794), .B(n5793), .Z(n5795) );
  XOR U1612 ( .A(in[228]), .B(n5795), .Z(n6106) );
  XNOR U1613 ( .A(n6106), .B(n5796), .Z(n8529) );
  XNOR U1614 ( .A(in[164]), .B(n8529), .Z(n9582) );
  XOR U1615 ( .A(in[324]), .B(in[644]), .Z(n5798) );
  XNOR U1616 ( .A(in[964]), .B(in[4]), .Z(n5797) );
  XNOR U1617 ( .A(n5798), .B(n5797), .Z(n5799) );
  XOR U1618 ( .A(in[1284]), .B(n5799), .Z(n6004) );
  XOR U1619 ( .A(in[773]), .B(in[1093]), .Z(n5801) );
  XNOR U1620 ( .A(in[453]), .B(in[1413]), .Z(n5800) );
  XNOR U1621 ( .A(n5801), .B(n5800), .Z(n5802) );
  XOR U1622 ( .A(in[133]), .B(n5802), .Z(n5928) );
  XNOR U1623 ( .A(n6004), .B(n5928), .Z(n8873) );
  XNOR U1624 ( .A(in[1349]), .B(n8873), .Z(n9579) );
  NAND U1625 ( .A(n9582), .B(n9579), .Z(n5803) );
  XNOR U1626 ( .A(n6338), .B(n5803), .Z(out[1057]) );
  XOR U1627 ( .A(in[1589]), .B(in[629]), .Z(n5805) );
  XNOR U1628 ( .A(in[949]), .B(in[309]), .Z(n5804) );
  XNOR U1629 ( .A(n5805), .B(n5804), .Z(n5806) );
  XOR U1630 ( .A(in[1269]), .B(n5806), .Z(n6242) );
  XNOR U1631 ( .A(n5807), .B(n6242), .Z(n8580) );
  XNOR U1632 ( .A(in[565]), .B(n8580), .Z(n6342) );
  XOR U1633 ( .A(in[1189]), .B(in[1509]), .Z(n5809) );
  XNOR U1634 ( .A(in[549]), .B(in[869]), .Z(n5808) );
  XNOR U1635 ( .A(n5809), .B(n5808), .Z(n5810) );
  XNOR U1636 ( .A(in[229]), .B(n5810), .Z(n6110) );
  XNOR U1637 ( .A(n5811), .B(n6110), .Z(n8533) );
  XNOR U1638 ( .A(in[165]), .B(n8533), .Z(n9586) );
  XOR U1639 ( .A(in[774]), .B(in[1094]), .Z(n5813) );
  XNOR U1640 ( .A(in[454]), .B(in[1414]), .Z(n5812) );
  XNOR U1641 ( .A(n5813), .B(n5812), .Z(n5814) );
  XOR U1642 ( .A(in[134]), .B(n5814), .Z(n5933) );
  XOR U1643 ( .A(in[325]), .B(in[645]), .Z(n5816) );
  XNOR U1644 ( .A(in[965]), .B(in[5]), .Z(n5815) );
  XNOR U1645 ( .A(n5816), .B(n5815), .Z(n5817) );
  XOR U1646 ( .A(in[1285]), .B(n5817), .Z(n6007) );
  XNOR U1647 ( .A(n5933), .B(n6007), .Z(n8876) );
  XNOR U1648 ( .A(in[1350]), .B(n8876), .Z(n9583) );
  NAND U1649 ( .A(n9586), .B(n9583), .Z(n5818) );
  XNOR U1650 ( .A(n6342), .B(n5818), .Z(out[1058]) );
  XOR U1651 ( .A(in[1590]), .B(in[630]), .Z(n5820) );
  XNOR U1652 ( .A(in[950]), .B(in[310]), .Z(n5819) );
  XNOR U1653 ( .A(n5820), .B(n5819), .Z(n5821) );
  XOR U1654 ( .A(in[1270]), .B(n5821), .Z(n6246) );
  XNOR U1655 ( .A(n5822), .B(n6246), .Z(n8584) );
  XNOR U1656 ( .A(in[566]), .B(n8584), .Z(n6346) );
  XOR U1657 ( .A(in[166]), .B(n8537), .Z(n9590) );
  XOR U1658 ( .A(in[775]), .B(in[1095]), .Z(n5824) );
  XNOR U1659 ( .A(in[455]), .B(in[1415]), .Z(n5823) );
  XNOR U1660 ( .A(n5824), .B(n5823), .Z(n5825) );
  XOR U1661 ( .A(in[135]), .B(n5825), .Z(n5938) );
  XOR U1662 ( .A(in[326]), .B(in[6]), .Z(n5827) );
  XNOR U1663 ( .A(in[966]), .B(in[646]), .Z(n5826) );
  XNOR U1664 ( .A(n5827), .B(n5826), .Z(n5828) );
  XOR U1665 ( .A(in[1286]), .B(n5828), .Z(n6010) );
  XNOR U1666 ( .A(n5938), .B(n6010), .Z(n8887) );
  XNOR U1667 ( .A(in[1351]), .B(n8887), .Z(n9587) );
  NAND U1668 ( .A(n9590), .B(n9587), .Z(n5829) );
  XNOR U1669 ( .A(n6346), .B(n5829), .Z(out[1059]) );
  XNOR U1670 ( .A(n5831), .B(n5830), .Z(n8419) );
  XNOR U1671 ( .A(in[576]), .B(n8419), .Z(n7368) );
  XOR U1672 ( .A(in[231]), .B(n8520), .Z(n7710) );
  XNOR U1673 ( .A(in[1451]), .B(n8557), .Z(n7707) );
  NAND U1674 ( .A(n7710), .B(n7707), .Z(n5832) );
  XNOR U1675 ( .A(n7368), .B(n5832), .Z(out[105]) );
  XOR U1676 ( .A(in[1591]), .B(in[631]), .Z(n5834) );
  XNOR U1677 ( .A(in[951]), .B(in[311]), .Z(n5833) );
  XNOR U1678 ( .A(n5834), .B(n5833), .Z(n5835) );
  XOR U1679 ( .A(in[1271]), .B(n5835), .Z(n6250) );
  XNOR U1680 ( .A(n5836), .B(n6250), .Z(n8588) );
  XNOR U1681 ( .A(in[567]), .B(n8588), .Z(n6350) );
  XOR U1682 ( .A(in[167]), .B(n8541), .Z(n9594) );
  XOR U1683 ( .A(in[327]), .B(in[7]), .Z(n5838) );
  XNOR U1684 ( .A(in[967]), .B(in[647]), .Z(n5837) );
  XNOR U1685 ( .A(n5838), .B(n5837), .Z(n5839) );
  XOR U1686 ( .A(in[1287]), .B(n5839), .Z(n6013) );
  XOR U1687 ( .A(in[776]), .B(in[1096]), .Z(n5841) );
  XNOR U1688 ( .A(in[456]), .B(in[1416]), .Z(n5840) );
  XNOR U1689 ( .A(n5841), .B(n5840), .Z(n5842) );
  XOR U1690 ( .A(in[136]), .B(n5842), .Z(n5943) );
  XNOR U1691 ( .A(n6013), .B(n5943), .Z(n8890) );
  XNOR U1692 ( .A(in[1352]), .B(n8890), .Z(n9591) );
  NAND U1693 ( .A(n9594), .B(n9591), .Z(n5843) );
  XNOR U1694 ( .A(n6350), .B(n5843), .Z(out[1060]) );
  XOR U1695 ( .A(in[632]), .B(in[1592]), .Z(n5845) );
  XNOR U1696 ( .A(in[1272]), .B(in[312]), .Z(n5844) );
  XNOR U1697 ( .A(n5845), .B(n5844), .Z(n5846) );
  XOR U1698 ( .A(in[952]), .B(n5846), .Z(n6254) );
  XNOR U1699 ( .A(n5847), .B(n6254), .Z(n8592) );
  XNOR U1700 ( .A(in[568]), .B(n8592), .Z(n6354) );
  XOR U1701 ( .A(in[168]), .B(n8545), .Z(n9598) );
  XNOR U1702 ( .A(in[1353]), .B(n8893), .Z(n9595) );
  NAND U1703 ( .A(n9598), .B(n9595), .Z(n5848) );
  XNOR U1704 ( .A(n6354), .B(n5848), .Z(out[1061]) );
  XOR U1705 ( .A(in[633]), .B(in[1593]), .Z(n5850) );
  XNOR U1706 ( .A(in[1273]), .B(in[313]), .Z(n5849) );
  XNOR U1707 ( .A(n5850), .B(n5849), .Z(n5851) );
  XOR U1708 ( .A(in[953]), .B(n5851), .Z(n6258) );
  XNOR U1709 ( .A(n5852), .B(n6258), .Z(n8596) );
  XNOR U1710 ( .A(in[569]), .B(n8596), .Z(n6359) );
  XOR U1711 ( .A(in[169]), .B(n8549), .Z(n9602) );
  XOR U1712 ( .A(in[329]), .B(in[969]), .Z(n5854) );
  XNOR U1713 ( .A(in[9]), .B(in[649]), .Z(n5853) );
  XNOR U1714 ( .A(n5854), .B(n5853), .Z(n5855) );
  XOR U1715 ( .A(in[1289]), .B(n5855), .Z(n6021) );
  XOR U1716 ( .A(in[778]), .B(in[1098]), .Z(n5857) );
  XNOR U1717 ( .A(in[458]), .B(in[1418]), .Z(n5856) );
  XNOR U1718 ( .A(n5857), .B(n5856), .Z(n5858) );
  XOR U1719 ( .A(in[138]), .B(n5858), .Z(n5956) );
  XNOR U1720 ( .A(n6021), .B(n5956), .Z(n8896) );
  XNOR U1721 ( .A(in[1354]), .B(n8896), .Z(n9599) );
  NAND U1722 ( .A(n9602), .B(n9599), .Z(n5859) );
  XNOR U1723 ( .A(n6359), .B(n5859), .Z(out[1062]) );
  XOR U1724 ( .A(in[634]), .B(in[1594]), .Z(n5861) );
  XNOR U1725 ( .A(in[1274]), .B(in[314]), .Z(n5860) );
  XNOR U1726 ( .A(n5861), .B(n5860), .Z(n5862) );
  XOR U1727 ( .A(in[954]), .B(n5862), .Z(n6262) );
  XNOR U1728 ( .A(n5863), .B(n6262), .Z(n8600) );
  XNOR U1729 ( .A(in[570]), .B(n8600), .Z(n6363) );
  XOR U1730 ( .A(in[170]), .B(n8553), .Z(n9606) );
  XOR U1731 ( .A(in[1290]), .B(in[650]), .Z(n5865) );
  XNOR U1732 ( .A(in[970]), .B(in[330]), .Z(n5864) );
  XNOR U1733 ( .A(n5865), .B(n5864), .Z(n5866) );
  XOR U1734 ( .A(in[10]), .B(n5866), .Z(n6024) );
  XOR U1735 ( .A(in[1419]), .B(in[779]), .Z(n5868) );
  XNOR U1736 ( .A(in[1099]), .B(in[459]), .Z(n5867) );
  XNOR U1737 ( .A(n5868), .B(n5867), .Z(n5869) );
  XOR U1738 ( .A(in[139]), .B(n5869), .Z(n5961) );
  XNOR U1739 ( .A(n6024), .B(n5961), .Z(n8899) );
  XNOR U1740 ( .A(in[1355]), .B(n8899), .Z(n9603) );
  NAND U1741 ( .A(n9606), .B(n9603), .Z(n5870) );
  XNOR U1742 ( .A(n6363), .B(n5870), .Z(out[1063]) );
  XOR U1743 ( .A(in[955]), .B(in[1275]), .Z(n5872) );
  XNOR U1744 ( .A(in[1595]), .B(in[315]), .Z(n5871) );
  XNOR U1745 ( .A(n5872), .B(n5871), .Z(n5873) );
  XNOR U1746 ( .A(in[635]), .B(n5873), .Z(n6266) );
  XNOR U1747 ( .A(n5874), .B(n6266), .Z(n8610) );
  XNOR U1748 ( .A(in[571]), .B(n8610), .Z(n6365) );
  NOR U1749 ( .A(n6108), .B(n6503), .Z(n5875) );
  XNOR U1750 ( .A(n6365), .B(n5875), .Z(out[1064]) );
  XOR U1751 ( .A(in[956]), .B(in[1276]), .Z(n5877) );
  XNOR U1752 ( .A(in[1596]), .B(in[316]), .Z(n5876) );
  XNOR U1753 ( .A(n5877), .B(n5876), .Z(n5878) );
  XNOR U1754 ( .A(in[636]), .B(n5878), .Z(n6270) );
  XNOR U1755 ( .A(n5879), .B(n6270), .Z(n8614) );
  XNOR U1756 ( .A(in[572]), .B(n8614), .Z(n6367) );
  NOR U1757 ( .A(n6112), .B(n6507), .Z(n5880) );
  XNOR U1758 ( .A(n6367), .B(n5880), .Z(out[1065]) );
  XOR U1759 ( .A(in[957]), .B(in[1277]), .Z(n5882) );
  XNOR U1760 ( .A(in[1597]), .B(in[317]), .Z(n5881) );
  XNOR U1761 ( .A(n5882), .B(n5881), .Z(n5883) );
  XNOR U1762 ( .A(in[637]), .B(n5883), .Z(n6275) );
  XNOR U1763 ( .A(n5884), .B(n6275), .Z(n8618) );
  XNOR U1764 ( .A(in[573]), .B(n8618), .Z(n6369) );
  NOR U1765 ( .A(n6117), .B(n6511), .Z(n5885) );
  XNOR U1766 ( .A(n6369), .B(n5885), .Z(out[1066]) );
  XOR U1767 ( .A(in[574]), .B(n8622), .Z(n6371) );
  NOR U1768 ( .A(n6121), .B(n6515), .Z(n5886) );
  XNOR U1769 ( .A(n6371), .B(n5886), .Z(out[1067]) );
  XOR U1770 ( .A(in[959]), .B(in[1279]), .Z(n5888) );
  XNOR U1771 ( .A(in[1599]), .B(in[319]), .Z(n5887) );
  XNOR U1772 ( .A(n5888), .B(n5887), .Z(n5889) );
  XNOR U1773 ( .A(in[639]), .B(n5889), .Z(n6283) );
  XNOR U1774 ( .A(n5890), .B(n6283), .Z(n8344) );
  XNOR U1775 ( .A(in[575]), .B(n8344), .Z(n6373) );
  NOR U1776 ( .A(n6125), .B(n6520), .Z(n5891) );
  XNOR U1777 ( .A(n6373), .B(n5891), .Z(out[1068]) );
  XOR U1778 ( .A(in[896]), .B(in[1216]), .Z(n5893) );
  XNOR U1779 ( .A(in[1536]), .B(in[256]), .Z(n5892) );
  XNOR U1780 ( .A(n5893), .B(n5892), .Z(n5894) );
  XNOR U1781 ( .A(in[576]), .B(n5894), .Z(n6287) );
  XNOR U1782 ( .A(n5895), .B(n6287), .Z(n8348) );
  XNOR U1783 ( .A(in[512]), .B(n8348), .Z(n6375) );
  NOR U1784 ( .A(n6129), .B(n6524), .Z(n5896) );
  XNOR U1785 ( .A(n6375), .B(n5896), .Z(out[1069]) );
  XNOR U1786 ( .A(n5898), .B(n5897), .Z(n8423) );
  XNOR U1787 ( .A(in[577]), .B(n8423), .Z(n7370) );
  XOR U1788 ( .A(in[232]), .B(n8524), .Z(n7724) );
  XNOR U1789 ( .A(in[1452]), .B(n8565), .Z(n7721) );
  NAND U1790 ( .A(n7724), .B(n7721), .Z(n5899) );
  XNOR U1791 ( .A(n7370), .B(n5899), .Z(out[106]) );
  XOR U1792 ( .A(in[897]), .B(in[1217]), .Z(n5901) );
  XNOR U1793 ( .A(in[1537]), .B(in[257]), .Z(n5900) );
  XNOR U1794 ( .A(n5901), .B(n5900), .Z(n5902) );
  XNOR U1795 ( .A(in[577]), .B(n5902), .Z(n6291) );
  XNOR U1796 ( .A(n5903), .B(n6291), .Z(n8352) );
  XNOR U1797 ( .A(in[513]), .B(n8352), .Z(n6377) );
  NOR U1798 ( .A(n6133), .B(n6528), .Z(n5904) );
  XNOR U1799 ( .A(n6377), .B(n5904), .Z(out[1070]) );
  XOR U1800 ( .A(in[1538]), .B(in[578]), .Z(n5906) );
  XNOR U1801 ( .A(in[898]), .B(in[258]), .Z(n5905) );
  XNOR U1802 ( .A(n5906), .B(n5905), .Z(n5907) );
  XNOR U1803 ( .A(in[1218]), .B(n5907), .Z(n6295) );
  XNOR U1804 ( .A(n5908), .B(n6295), .Z(n8356) );
  XNOR U1805 ( .A(in[514]), .B(n8356), .Z(n6379) );
  NOR U1806 ( .A(n6137), .B(n6532), .Z(n5909) );
  XNOR U1807 ( .A(n6379), .B(n5909), .Z(out[1071]) );
  XOR U1808 ( .A(in[1539]), .B(in[579]), .Z(n5911) );
  XNOR U1809 ( .A(in[899]), .B(in[259]), .Z(n5910) );
  XNOR U1810 ( .A(n5911), .B(n5910), .Z(n5912) );
  XNOR U1811 ( .A(in[1219]), .B(n5912), .Z(n6299) );
  XNOR U1812 ( .A(n5913), .B(n6299), .Z(n8360) );
  XNOR U1813 ( .A(in[515]), .B(n8360), .Z(n6383) );
  NOR U1814 ( .A(n6141), .B(n6536), .Z(n5914) );
  XNOR U1815 ( .A(n6383), .B(n5914), .Z(out[1072]) );
  XOR U1816 ( .A(in[1540]), .B(in[580]), .Z(n5916) );
  XNOR U1817 ( .A(in[900]), .B(in[260]), .Z(n5915) );
  XNOR U1818 ( .A(n5916), .B(n5915), .Z(n5917) );
  XNOR U1819 ( .A(in[1220]), .B(n5917), .Z(n6303) );
  XNOR U1820 ( .A(n5918), .B(n6303), .Z(n8364) );
  XNOR U1821 ( .A(in[516]), .B(n8364), .Z(n6385) );
  NOR U1822 ( .A(n6145), .B(n6540), .Z(n5919) );
  XNOR U1823 ( .A(n6385), .B(n5919), .Z(out[1073]) );
  XOR U1824 ( .A(in[1541]), .B(in[581]), .Z(n5921) );
  XNOR U1825 ( .A(in[901]), .B(in[261]), .Z(n5920) );
  XNOR U1826 ( .A(n5921), .B(n5920), .Z(n5922) );
  XNOR U1827 ( .A(in[1221]), .B(n5922), .Z(n6307) );
  XNOR U1828 ( .A(n5923), .B(n6307), .Z(n8368) );
  XNOR U1829 ( .A(in[517]), .B(n8368), .Z(n6387) );
  NOR U1830 ( .A(n6149), .B(n6544), .Z(n5924) );
  XNOR U1831 ( .A(n6387), .B(n5924), .Z(out[1074]) );
  XOR U1832 ( .A(in[1542]), .B(in[582]), .Z(n5926) );
  XNOR U1833 ( .A(in[902]), .B(in[262]), .Z(n5925) );
  XNOR U1834 ( .A(n5926), .B(n5925), .Z(n5927) );
  XNOR U1835 ( .A(in[1222]), .B(n5927), .Z(n6311) );
  XNOR U1836 ( .A(n5928), .B(n6311), .Z(n8372) );
  XNOR U1837 ( .A(in[518]), .B(n8372), .Z(n6389) );
  NOR U1838 ( .A(n6153), .B(n6548), .Z(n5929) );
  XNOR U1839 ( .A(n6389), .B(n5929), .Z(out[1075]) );
  XOR U1840 ( .A(in[1543]), .B(in[583]), .Z(n5931) );
  XNOR U1841 ( .A(in[903]), .B(in[263]), .Z(n5930) );
  XNOR U1842 ( .A(n5931), .B(n5930), .Z(n5932) );
  XNOR U1843 ( .A(in[1223]), .B(n5932), .Z(n6316) );
  XNOR U1844 ( .A(n5933), .B(n6316), .Z(n8376) );
  XNOR U1845 ( .A(in[519]), .B(n8376), .Z(n6391) );
  NOR U1846 ( .A(n6158), .B(n6552), .Z(n5934) );
  XNOR U1847 ( .A(n6391), .B(n5934), .Z(out[1076]) );
  XOR U1848 ( .A(in[1544]), .B(in[584]), .Z(n5936) );
  XNOR U1849 ( .A(in[904]), .B(in[264]), .Z(n5935) );
  XNOR U1850 ( .A(n5936), .B(n5935), .Z(n5937) );
  XNOR U1851 ( .A(in[1224]), .B(n5937), .Z(n6320) );
  XNOR U1852 ( .A(n5938), .B(n6320), .Z(n8380) );
  XNOR U1853 ( .A(in[520]), .B(n8380), .Z(n6393) );
  NOR U1854 ( .A(n6162), .B(n6556), .Z(n5939) );
  XNOR U1855 ( .A(n6393), .B(n5939), .Z(out[1077]) );
  XOR U1856 ( .A(in[1545]), .B(in[585]), .Z(n5941) );
  XNOR U1857 ( .A(in[905]), .B(in[265]), .Z(n5940) );
  XNOR U1858 ( .A(n5941), .B(n5940), .Z(n5942) );
  XNOR U1859 ( .A(in[1225]), .B(n5942), .Z(n6324) );
  XNOR U1860 ( .A(n5943), .B(n6324), .Z(n8388) );
  XNOR U1861 ( .A(in[521]), .B(n8388), .Z(n6395) );
  NOR U1862 ( .A(n6166), .B(n6561), .Z(n5944) );
  XNOR U1863 ( .A(n6395), .B(n5944), .Z(out[1078]) );
  XOR U1864 ( .A(in[1546]), .B(in[586]), .Z(n5946) );
  XNOR U1865 ( .A(in[906]), .B(in[266]), .Z(n5945) );
  XNOR U1866 ( .A(n5946), .B(n5945), .Z(n5947) );
  XNOR U1867 ( .A(in[1226]), .B(n5947), .Z(n6328) );
  XNOR U1868 ( .A(n5948), .B(n6328), .Z(n8392) );
  XNOR U1869 ( .A(in[522]), .B(n8392), .Z(n6397) );
  NOR U1870 ( .A(n6170), .B(n6565), .Z(n5949) );
  XNOR U1871 ( .A(n6397), .B(n5949), .Z(out[1079]) );
  XNOR U1872 ( .A(n5951), .B(n5950), .Z(n8431) );
  XNOR U1873 ( .A(in[578]), .B(n8431), .Z(n7372) );
  XOR U1874 ( .A(in[233]), .B(n8528), .Z(n7738) );
  XNOR U1875 ( .A(in[1453]), .B(n8569), .Z(n7735) );
  NAND U1876 ( .A(n7738), .B(n7735), .Z(n5952) );
  XNOR U1877 ( .A(n7372), .B(n5952), .Z(out[107]) );
  XOR U1878 ( .A(in[1547]), .B(in[587]), .Z(n5954) );
  XNOR U1879 ( .A(in[907]), .B(in[267]), .Z(n5953) );
  XNOR U1880 ( .A(n5954), .B(n5953), .Z(n5955) );
  XNOR U1881 ( .A(in[1227]), .B(n5955), .Z(n6332) );
  XNOR U1882 ( .A(n5956), .B(n6332), .Z(n8396) );
  XNOR U1883 ( .A(in[523]), .B(n8396), .Z(n6399) );
  NOR U1884 ( .A(n6174), .B(n6569), .Z(n5957) );
  XNOR U1885 ( .A(n6399), .B(n5957), .Z(out[1080]) );
  XOR U1886 ( .A(in[1548]), .B(in[588]), .Z(n5959) );
  XNOR U1887 ( .A(in[908]), .B(in[268]), .Z(n5958) );
  XNOR U1888 ( .A(n5959), .B(n5958), .Z(n5960) );
  XNOR U1889 ( .A(in[1228]), .B(n5960), .Z(n6336) );
  XNOR U1890 ( .A(n5961), .B(n6336), .Z(n8400) );
  XNOR U1891 ( .A(in[524]), .B(n8400), .Z(n6401) );
  NOR U1892 ( .A(n6178), .B(n6573), .Z(n5962) );
  XNOR U1893 ( .A(n6401), .B(n5962), .Z(out[1081]) );
  XOR U1894 ( .A(in[1549]), .B(in[589]), .Z(n5964) );
  XNOR U1895 ( .A(in[909]), .B(in[269]), .Z(n5963) );
  XNOR U1896 ( .A(n5964), .B(n5963), .Z(n5965) );
  XOR U1897 ( .A(in[1229]), .B(n5965), .Z(n6340) );
  XNOR U1898 ( .A(n6340), .B(n5966), .Z(n8404) );
  XNOR U1899 ( .A(in[525]), .B(n8404), .Z(n6404) );
  NOR U1900 ( .A(n6182), .B(n6577), .Z(n5967) );
  XNOR U1901 ( .A(n6404), .B(n5967), .Z(out[1082]) );
  XOR U1902 ( .A(in[1550]), .B(in[590]), .Z(n5969) );
  XNOR U1903 ( .A(in[910]), .B(in[270]), .Z(n5968) );
  XNOR U1904 ( .A(n5969), .B(n5968), .Z(n5970) );
  XOR U1905 ( .A(in[1230]), .B(n5970), .Z(n6344) );
  XNOR U1906 ( .A(n6344), .B(n5971), .Z(n8408) );
  XNOR U1907 ( .A(in[526]), .B(n8408), .Z(n6406) );
  NOR U1908 ( .A(n6186), .B(n6581), .Z(n5972) );
  XNOR U1909 ( .A(n6406), .B(n5972), .Z(out[1083]) );
  XOR U1910 ( .A(in[1551]), .B(in[591]), .Z(n5974) );
  XNOR U1911 ( .A(in[911]), .B(in[271]), .Z(n5973) );
  XNOR U1912 ( .A(n5974), .B(n5973), .Z(n5975) );
  XOR U1913 ( .A(in[1231]), .B(n5975), .Z(n6348) );
  XNOR U1914 ( .A(n6348), .B(n5976), .Z(n8412) );
  XNOR U1915 ( .A(in[527]), .B(n8412), .Z(n6408) );
  NOR U1916 ( .A(n6190), .B(n6585), .Z(n5977) );
  XNOR U1917 ( .A(n6408), .B(n5977), .Z(out[1084]) );
  XOR U1918 ( .A(in[1552]), .B(in[592]), .Z(n5979) );
  XNOR U1919 ( .A(in[912]), .B(in[272]), .Z(n5978) );
  XNOR U1920 ( .A(n5979), .B(n5978), .Z(n5980) );
  XNOR U1921 ( .A(in[1232]), .B(n5980), .Z(n6352) );
  XNOR U1922 ( .A(n5981), .B(n6352), .Z(n8416) );
  XNOR U1923 ( .A(in[528]), .B(n8416), .Z(n6410) );
  NOR U1924 ( .A(n6194), .B(n6589), .Z(n5982) );
  XNOR U1925 ( .A(n6410), .B(n5982), .Z(out[1085]) );
  XOR U1926 ( .A(in[1553]), .B(in[593]), .Z(n5984) );
  XNOR U1927 ( .A(in[913]), .B(in[273]), .Z(n5983) );
  XNOR U1928 ( .A(n5984), .B(n5983), .Z(n5985) );
  XNOR U1929 ( .A(in[1233]), .B(n5985), .Z(n6357) );
  XNOR U1930 ( .A(n5986), .B(n6357), .Z(n8420) );
  XNOR U1931 ( .A(in[529]), .B(n8420), .Z(n6412) );
  NOR U1932 ( .A(n6197), .B(n6593), .Z(n5987) );
  XNOR U1933 ( .A(n6412), .B(n5987), .Z(out[1086]) );
  XOR U1934 ( .A(in[1554]), .B(in[594]), .Z(n5989) );
  XNOR U1935 ( .A(in[914]), .B(in[274]), .Z(n5988) );
  XNOR U1936 ( .A(n5989), .B(n5988), .Z(n5990) );
  XNOR U1937 ( .A(in[1234]), .B(n5990), .Z(n6361) );
  XNOR U1938 ( .A(n5991), .B(n6361), .Z(n8424) );
  XNOR U1939 ( .A(in[530]), .B(n8424), .Z(n6414) );
  NOR U1940 ( .A(n6199), .B(n6597), .Z(n5992) );
  XNOR U1941 ( .A(n6414), .B(n5992), .Z(out[1087]) );
  XOR U1942 ( .A(in[957]), .B(n8407), .Z(n6416) );
  NOR U1943 ( .A(n6203), .B(n9438), .Z(n5993) );
  XNOR U1944 ( .A(n6416), .B(n5993), .Z(out[1088]) );
  XOR U1945 ( .A(in[958]), .B(n8411), .Z(n6418) );
  NOR U1946 ( .A(n6207), .B(n9442), .Z(n5994) );
  XNOR U1947 ( .A(n6418), .B(n5994), .Z(out[1089]) );
  XOR U1948 ( .A(n5996), .B(n5995), .Z(n8435) );
  XNOR U1949 ( .A(in[579]), .B(n8435), .Z(n7374) );
  XOR U1950 ( .A(in[234]), .B(n8532), .Z(n7754) );
  XNOR U1951 ( .A(in[1454]), .B(n8573), .Z(n7751) );
  NAND U1952 ( .A(n7754), .B(n7751), .Z(n5997) );
  XNOR U1953 ( .A(n7374), .B(n5997), .Z(out[108]) );
  XOR U1954 ( .A(in[959]), .B(n8415), .Z(n6420) );
  NOR U1955 ( .A(n6211), .B(n9446), .Z(n5998) );
  XNOR U1956 ( .A(n6420), .B(n5998), .Z(out[1090]) );
  XOR U1957 ( .A(in[896]), .B(n8419), .Z(n6422) );
  NOR U1958 ( .A(n6215), .B(n9450), .Z(n5999) );
  XNOR U1959 ( .A(n6422), .B(n5999), .Z(out[1091]) );
  XOR U1960 ( .A(in[897]), .B(n8423), .Z(n6425) );
  NOR U1961 ( .A(n6219), .B(n9454), .Z(n6000) );
  XNOR U1962 ( .A(n6425), .B(n6000), .Z(out[1092]) );
  XOR U1963 ( .A(in[898]), .B(n8431), .Z(n6427) );
  NOR U1964 ( .A(n6223), .B(n9458), .Z(n6001) );
  XNOR U1965 ( .A(n6427), .B(n6001), .Z(out[1093]) );
  XOR U1966 ( .A(in[899]), .B(n8435), .Z(n6429) );
  NOR U1967 ( .A(n6227), .B(n9462), .Z(n6002) );
  XNOR U1968 ( .A(n6429), .B(n6002), .Z(out[1094]) );
  XNOR U1969 ( .A(n6004), .B(n6003), .Z(n8439) );
  XNOR U1970 ( .A(in[900]), .B(n8439), .Z(n6431) );
  NOR U1971 ( .A(n6231), .B(n9466), .Z(n6005) );
  XNOR U1972 ( .A(n6431), .B(n6005), .Z(out[1095]) );
  XNOR U1973 ( .A(n6007), .B(n6006), .Z(n8443) );
  XNOR U1974 ( .A(in[901]), .B(n8443), .Z(n6433) );
  NOR U1975 ( .A(n6236), .B(n9470), .Z(n6008) );
  XNOR U1976 ( .A(n6433), .B(n6008), .Z(out[1096]) );
  XNOR U1977 ( .A(n6010), .B(n6009), .Z(n8447) );
  XNOR U1978 ( .A(in[902]), .B(n8447), .Z(n6435) );
  NOR U1979 ( .A(n6240), .B(n9474), .Z(n6011) );
  XNOR U1980 ( .A(n6435), .B(n6011), .Z(out[1097]) );
  XNOR U1981 ( .A(n6013), .B(n6012), .Z(n8451) );
  XNOR U1982 ( .A(in[903]), .B(n8451), .Z(n6437) );
  NOR U1983 ( .A(n6244), .B(n9482), .Z(n6014) );
  XNOR U1984 ( .A(n6437), .B(n6014), .Z(out[1098]) );
  XNOR U1985 ( .A(n6016), .B(n6015), .Z(n8455) );
  XNOR U1986 ( .A(in[904]), .B(n8455), .Z(n6439) );
  NOR U1987 ( .A(n6248), .B(n9486), .Z(n6017) );
  XNOR U1988 ( .A(n6439), .B(n6017), .Z(out[1099]) );
  XOR U1989 ( .A(in[580]), .B(n8439), .Z(n7376) );
  XOR U1990 ( .A(in[235]), .B(n8536), .Z(n7778) );
  XNOR U1991 ( .A(in[1455]), .B(n8577), .Z(n7775) );
  NAND U1992 ( .A(n7778), .B(n7775), .Z(n6018) );
  XNOR U1993 ( .A(n7376), .B(n6018), .Z(out[109]) );
  XOR U1994 ( .A(in[200]), .B(n8380), .Z(n8728) );
  XNOR U1995 ( .A(in[1420]), .B(n8421), .Z(n8727) );
  XOR U1996 ( .A(n8927), .B(in[1043]), .Z(n7439) );
  NAND U1997 ( .A(n8727), .B(n7439), .Z(n6019) );
  XNOR U1998 ( .A(n8728), .B(n6019), .Z(out[10]) );
  XNOR U1999 ( .A(n6021), .B(n6020), .Z(n8459) );
  XNOR U2000 ( .A(in[905]), .B(n8459), .Z(n6441) );
  NOR U2001 ( .A(n6252), .B(n9490), .Z(n6022) );
  XNOR U2002 ( .A(n6441), .B(n6022), .Z(out[1100]) );
  XNOR U2003 ( .A(n6024), .B(n6023), .Z(n8463) );
  XNOR U2004 ( .A(in[906]), .B(n8463), .Z(n6443) );
  NOR U2005 ( .A(n6256), .B(n9494), .Z(n6025) );
  XNOR U2006 ( .A(n6443), .B(n6025), .Z(out[1101]) );
  XNOR U2007 ( .A(n6027), .B(n6026), .Z(n8467) );
  XNOR U2008 ( .A(in[907]), .B(n8467), .Z(n6446) );
  NOR U2009 ( .A(n6260), .B(n9498), .Z(n6028) );
  XNOR U2010 ( .A(n6446), .B(n6028), .Z(out[1102]) );
  XOR U2011 ( .A(n6030), .B(n6029), .Z(n8475) );
  XNOR U2012 ( .A(in[908]), .B(n8475), .Z(n6448) );
  NOR U2013 ( .A(n6264), .B(n9502), .Z(n6031) );
  XNOR U2014 ( .A(n6448), .B(n6031), .Z(out[1103]) );
  XNOR U2015 ( .A(n6033), .B(n6032), .Z(n8479) );
  XNOR U2016 ( .A(in[909]), .B(n8479), .Z(n6450) );
  NOR U2017 ( .A(n6268), .B(n9506), .Z(n6034) );
  XNOR U2018 ( .A(n6450), .B(n6034), .Z(out[1104]) );
  XOR U2019 ( .A(n6036), .B(n6035), .Z(n8483) );
  XNOR U2020 ( .A(in[910]), .B(n8483), .Z(n6452) );
  NOR U2021 ( .A(n6272), .B(n9510), .Z(n6037) );
  XNOR U2022 ( .A(n6452), .B(n6037), .Z(out[1105]) );
  XOR U2023 ( .A(n6039), .B(n6038), .Z(n8487) );
  XNOR U2024 ( .A(in[911]), .B(n8487), .Z(n6454) );
  NOR U2025 ( .A(n6277), .B(n9514), .Z(n6040) );
  XNOR U2026 ( .A(n6454), .B(n6040), .Z(out[1106]) );
  XOR U2027 ( .A(n6042), .B(n6041), .Z(n8491) );
  XNOR U2028 ( .A(in[912]), .B(n8491), .Z(n6456) );
  NOR U2029 ( .A(n6281), .B(n9518), .Z(n6043) );
  XNOR U2030 ( .A(n6456), .B(n6043), .Z(out[1107]) );
  XNOR U2031 ( .A(n6045), .B(n6044), .Z(n8495) );
  XNOR U2032 ( .A(in[913]), .B(n8495), .Z(n6458) );
  NOR U2033 ( .A(n6285), .B(n9526), .Z(n6046) );
  XNOR U2034 ( .A(n6458), .B(n6046), .Z(out[1108]) );
  XOR U2035 ( .A(n6048), .B(n6047), .Z(n8499) );
  XNOR U2036 ( .A(in[914]), .B(n8499), .Z(n6460) );
  NOR U2037 ( .A(n6289), .B(n9530), .Z(n6049) );
  XNOR U2038 ( .A(n6460), .B(n6049), .Z(out[1109]) );
  XOR U2039 ( .A(in[581]), .B(n8443), .Z(n7378) );
  XOR U2040 ( .A(in[236]), .B(n8540), .Z(n7802) );
  XNOR U2041 ( .A(in[1456]), .B(n8581), .Z(n7799) );
  NAND U2042 ( .A(n7802), .B(n7799), .Z(n6050) );
  XNOR U2043 ( .A(n7378), .B(n6050), .Z(out[110]) );
  XOR U2044 ( .A(n6052), .B(n6051), .Z(n8503) );
  XNOR U2045 ( .A(in[915]), .B(n8503), .Z(n6462) );
  NOR U2046 ( .A(n6293), .B(n9534), .Z(n6053) );
  XNOR U2047 ( .A(n6462), .B(n6053), .Z(out[1110]) );
  XNOR U2048 ( .A(n6055), .B(n6054), .Z(n8507) );
  XNOR U2049 ( .A(in[916]), .B(n8507), .Z(n6464) );
  NOR U2050 ( .A(n6297), .B(n9538), .Z(n6056) );
  XNOR U2051 ( .A(n6464), .B(n6056), .Z(out[1111]) );
  XNOR U2052 ( .A(n6058), .B(n6057), .Z(n8511) );
  XNOR U2053 ( .A(in[917]), .B(n8511), .Z(n6467) );
  NOR U2054 ( .A(n6301), .B(n9542), .Z(n6059) );
  XNOR U2055 ( .A(n6467), .B(n6059), .Z(out[1112]) );
  XOR U2056 ( .A(n6061), .B(n6060), .Z(n8519) );
  XNOR U2057 ( .A(in[918]), .B(n8519), .Z(n6469) );
  NOR U2058 ( .A(n6305), .B(n9546), .Z(n6062) );
  XNOR U2059 ( .A(n6469), .B(n6062), .Z(out[1113]) );
  XNOR U2060 ( .A(n6064), .B(n6063), .Z(n8523) );
  XNOR U2061 ( .A(in[919]), .B(n8523), .Z(n6471) );
  NOR U2062 ( .A(n6309), .B(n9550), .Z(n6065) );
  XNOR U2063 ( .A(n6471), .B(n6065), .Z(out[1114]) );
  XNOR U2064 ( .A(n6067), .B(n6066), .Z(n8527) );
  XNOR U2065 ( .A(in[920]), .B(n8527), .Z(n6473) );
  NOR U2066 ( .A(n6313), .B(n9554), .Z(n6068) );
  XNOR U2067 ( .A(n6473), .B(n6068), .Z(out[1115]) );
  XNOR U2068 ( .A(n6070), .B(n6069), .Z(n8531) );
  XNOR U2069 ( .A(in[921]), .B(n8531), .Z(n6475) );
  NOR U2070 ( .A(n6318), .B(n9558), .Z(n6071) );
  XNOR U2071 ( .A(n6475), .B(n6071), .Z(out[1116]) );
  XOR U2072 ( .A(n6073), .B(n6072), .Z(n8535) );
  XNOR U2073 ( .A(in[922]), .B(n8535), .Z(n6477) );
  NOR U2074 ( .A(n6322), .B(n9562), .Z(n6074) );
  XNOR U2075 ( .A(n6477), .B(n6074), .Z(out[1117]) );
  XOR U2076 ( .A(n6076), .B(n6075), .Z(n8539) );
  XNOR U2077 ( .A(in[923]), .B(n8539), .Z(n6479) );
  NOR U2078 ( .A(n6326), .B(n9570), .Z(n6077) );
  XNOR U2079 ( .A(n6479), .B(n6077), .Z(out[1118]) );
  XOR U2080 ( .A(n6079), .B(n6078), .Z(n8543) );
  XNOR U2081 ( .A(in[924]), .B(n8543), .Z(n6481) );
  NOR U2082 ( .A(n6330), .B(n9574), .Z(n6080) );
  XNOR U2083 ( .A(n6481), .B(n6080), .Z(out[1119]) );
  XOR U2084 ( .A(in[582]), .B(n8447), .Z(n7380) );
  XOR U2085 ( .A(in[237]), .B(n8544), .Z(n7826) );
  XNOR U2086 ( .A(in[1457]), .B(n8585), .Z(n7823) );
  NAND U2087 ( .A(n7826), .B(n7823), .Z(n6081) );
  XNOR U2088 ( .A(n7380), .B(n6081), .Z(out[111]) );
  XOR U2089 ( .A(n6083), .B(n6082), .Z(n8547) );
  XNOR U2090 ( .A(in[925]), .B(n8547), .Z(n6483) );
  NOR U2091 ( .A(n6334), .B(n9578), .Z(n6084) );
  XNOR U2092 ( .A(n6483), .B(n6084), .Z(out[1120]) );
  XOR U2093 ( .A(n6086), .B(n6085), .Z(n8551) );
  XNOR U2094 ( .A(in[926]), .B(n8551), .Z(n6485) );
  NOR U2095 ( .A(n6338), .B(n9582), .Z(n6087) );
  XNOR U2096 ( .A(n6485), .B(n6087), .Z(out[1121]) );
  XOR U2097 ( .A(n6089), .B(n6088), .Z(n8555) );
  XNOR U2098 ( .A(in[927]), .B(n8555), .Z(n6488) );
  NOR U2099 ( .A(n6342), .B(n9586), .Z(n6090) );
  XNOR U2100 ( .A(n6488), .B(n6090), .Z(out[1122]) );
  XOR U2101 ( .A(n6092), .B(n6091), .Z(n8563) );
  XNOR U2102 ( .A(in[928]), .B(n8563), .Z(n6490) );
  NOR U2103 ( .A(n6346), .B(n9590), .Z(n6093) );
  XNOR U2104 ( .A(n6490), .B(n6093), .Z(out[1123]) );
  XNOR U2105 ( .A(n6095), .B(n6094), .Z(n8567) );
  XNOR U2106 ( .A(in[929]), .B(n8567), .Z(n6492) );
  NOR U2107 ( .A(n6350), .B(n9594), .Z(n6096) );
  XNOR U2108 ( .A(n6492), .B(n6096), .Z(out[1124]) );
  XNOR U2109 ( .A(n6098), .B(n6097), .Z(n8571) );
  XNOR U2110 ( .A(in[930]), .B(n8571), .Z(n6494) );
  NOR U2111 ( .A(n6354), .B(n9598), .Z(n6099) );
  XNOR U2112 ( .A(n6494), .B(n6099), .Z(out[1125]) );
  XNOR U2113 ( .A(n6101), .B(n6100), .Z(n8575) );
  XNOR U2114 ( .A(in[931]), .B(n8575), .Z(n6496) );
  NOR U2115 ( .A(n6359), .B(n9602), .Z(n6102) );
  XNOR U2116 ( .A(n6496), .B(n6102), .Z(out[1126]) );
  XNOR U2117 ( .A(n6104), .B(n6103), .Z(n8579) );
  XNOR U2118 ( .A(in[932]), .B(n8579), .Z(n6498) );
  NOR U2119 ( .A(n6363), .B(n9606), .Z(n6105) );
  XNOR U2120 ( .A(n6498), .B(n6105), .Z(out[1127]) );
  XNOR U2121 ( .A(n6107), .B(n6106), .Z(n8583) );
  XNOR U2122 ( .A(in[933]), .B(n8583), .Z(n6501) );
  NAND U2123 ( .A(n6365), .B(n6108), .Z(n6109) );
  XNOR U2124 ( .A(n6501), .B(n6109), .Z(out[1128]) );
  XOR U2125 ( .A(n6111), .B(n6110), .Z(n8587) );
  XNOR U2126 ( .A(in[934]), .B(n8587), .Z(n6505) );
  NAND U2127 ( .A(n6367), .B(n6112), .Z(n6113) );
  XNOR U2128 ( .A(n6505), .B(n6113), .Z(out[1129]) );
  XOR U2129 ( .A(in[583]), .B(n8451), .Z(n7383) );
  XOR U2130 ( .A(in[238]), .B(n8548), .Z(n7850) );
  XNOR U2131 ( .A(in[1458]), .B(n8589), .Z(n7847) );
  NAND U2132 ( .A(n7850), .B(n7847), .Z(n6114) );
  XNOR U2133 ( .A(n7383), .B(n6114), .Z(out[112]) );
  XNOR U2134 ( .A(n6116), .B(n6115), .Z(n8591) );
  XNOR U2135 ( .A(in[935]), .B(n8591), .Z(n6509) );
  NAND U2136 ( .A(n6369), .B(n6117), .Z(n6118) );
  XNOR U2137 ( .A(n6509), .B(n6118), .Z(out[1130]) );
  XNOR U2138 ( .A(n6120), .B(n6119), .Z(n8595) );
  XNOR U2139 ( .A(in[936]), .B(n8595), .Z(n6513) );
  NAND U2140 ( .A(n6371), .B(n6121), .Z(n6122) );
  XNOR U2141 ( .A(n6513), .B(n6122), .Z(out[1131]) );
  XNOR U2142 ( .A(n6124), .B(n6123), .Z(n8599) );
  XNOR U2143 ( .A(in[937]), .B(n8599), .Z(n6518) );
  NAND U2144 ( .A(n6373), .B(n6125), .Z(n6126) );
  XNOR U2145 ( .A(n6518), .B(n6126), .Z(out[1132]) );
  XNOR U2146 ( .A(n6128), .B(n6127), .Z(n8609) );
  XNOR U2147 ( .A(in[938]), .B(n8609), .Z(n6522) );
  NAND U2148 ( .A(n6375), .B(n6129), .Z(n6130) );
  XNOR U2149 ( .A(n6522), .B(n6130), .Z(out[1133]) );
  XNOR U2150 ( .A(n6132), .B(n6131), .Z(n8613) );
  XNOR U2151 ( .A(in[939]), .B(n8613), .Z(n6526) );
  NAND U2152 ( .A(n6377), .B(n6133), .Z(n6134) );
  XNOR U2153 ( .A(n6526), .B(n6134), .Z(out[1134]) );
  XNOR U2154 ( .A(n6136), .B(n6135), .Z(n8617) );
  XNOR U2155 ( .A(in[940]), .B(n8617), .Z(n6530) );
  NAND U2156 ( .A(n6379), .B(n6137), .Z(n6138) );
  XNOR U2157 ( .A(n6530), .B(n6138), .Z(out[1135]) );
  XNOR U2158 ( .A(n6140), .B(n6139), .Z(n8621) );
  XNOR U2159 ( .A(in[941]), .B(n8621), .Z(n6534) );
  NAND U2160 ( .A(n6383), .B(n6141), .Z(n6142) );
  XNOR U2161 ( .A(n6534), .B(n6142), .Z(out[1136]) );
  XNOR U2162 ( .A(n6144), .B(n6143), .Z(n8343) );
  XNOR U2163 ( .A(in[942]), .B(n8343), .Z(n6538) );
  NAND U2164 ( .A(n6385), .B(n6145), .Z(n6146) );
  XNOR U2165 ( .A(n6538), .B(n6146), .Z(out[1137]) );
  XNOR U2166 ( .A(n6148), .B(n6147), .Z(n8347) );
  XNOR U2167 ( .A(in[943]), .B(n8347), .Z(n6542) );
  NAND U2168 ( .A(n6387), .B(n6149), .Z(n6150) );
  XNOR U2169 ( .A(n6542), .B(n6150), .Z(out[1138]) );
  XNOR U2170 ( .A(n6152), .B(n6151), .Z(n8351) );
  XNOR U2171 ( .A(in[944]), .B(n8351), .Z(n6546) );
  NAND U2172 ( .A(n6389), .B(n6153), .Z(n6154) );
  XNOR U2173 ( .A(n6546), .B(n6154), .Z(out[1139]) );
  XOR U2174 ( .A(in[584]), .B(n8455), .Z(n7385) );
  XOR U2175 ( .A(in[239]), .B(n8552), .Z(n7874) );
  XNOR U2176 ( .A(in[1459]), .B(n8593), .Z(n7871) );
  NAND U2177 ( .A(n7874), .B(n7871), .Z(n6155) );
  XNOR U2178 ( .A(n7385), .B(n6155), .Z(out[113]) );
  XNOR U2179 ( .A(n6157), .B(n6156), .Z(n8355) );
  XNOR U2180 ( .A(in[945]), .B(n8355), .Z(n6550) );
  NAND U2181 ( .A(n6391), .B(n6158), .Z(n6159) );
  XNOR U2182 ( .A(n6550), .B(n6159), .Z(out[1140]) );
  XNOR U2183 ( .A(n6161), .B(n6160), .Z(n8359) );
  XNOR U2184 ( .A(in[946]), .B(n8359), .Z(n6554) );
  NAND U2185 ( .A(n6393), .B(n6162), .Z(n6163) );
  XNOR U2186 ( .A(n6554), .B(n6163), .Z(out[1141]) );
  XNOR U2187 ( .A(n6165), .B(n6164), .Z(n8363) );
  XNOR U2188 ( .A(in[947]), .B(n8363), .Z(n6559) );
  NAND U2189 ( .A(n6395), .B(n6166), .Z(n6167) );
  XNOR U2190 ( .A(n6559), .B(n6167), .Z(out[1142]) );
  XNOR U2191 ( .A(n6169), .B(n6168), .Z(n8367) );
  XNOR U2192 ( .A(in[948]), .B(n8367), .Z(n6563) );
  NAND U2193 ( .A(n6397), .B(n6170), .Z(n6171) );
  XNOR U2194 ( .A(n6563), .B(n6171), .Z(out[1143]) );
  XNOR U2195 ( .A(n6173), .B(n6172), .Z(n8371) );
  XNOR U2196 ( .A(in[949]), .B(n8371), .Z(n6567) );
  NAND U2197 ( .A(n6399), .B(n6174), .Z(n6175) );
  XNOR U2198 ( .A(n6567), .B(n6175), .Z(out[1144]) );
  XNOR U2199 ( .A(n6177), .B(n6176), .Z(n8375) );
  XNOR U2200 ( .A(in[950]), .B(n8375), .Z(n6571) );
  NAND U2201 ( .A(n6401), .B(n6178), .Z(n6179) );
  XNOR U2202 ( .A(n6571), .B(n6179), .Z(out[1145]) );
  XNOR U2203 ( .A(n6181), .B(n6180), .Z(n8379) );
  XNOR U2204 ( .A(in[951]), .B(n8379), .Z(n6575) );
  NAND U2205 ( .A(n6404), .B(n6182), .Z(n6183) );
  XNOR U2206 ( .A(n6575), .B(n6183), .Z(out[1146]) );
  XNOR U2207 ( .A(n6185), .B(n6184), .Z(n8387) );
  XNOR U2208 ( .A(in[952]), .B(n8387), .Z(n6579) );
  NAND U2209 ( .A(n6406), .B(n6186), .Z(n6187) );
  XNOR U2210 ( .A(n6579), .B(n6187), .Z(out[1147]) );
  XNOR U2211 ( .A(n6189), .B(n6188), .Z(n8391) );
  XNOR U2212 ( .A(in[953]), .B(n8391), .Z(n6583) );
  NAND U2213 ( .A(n6408), .B(n6190), .Z(n6191) );
  XNOR U2214 ( .A(n6583), .B(n6191), .Z(out[1148]) );
  XNOR U2215 ( .A(n6193), .B(n6192), .Z(n8395) );
  XNOR U2216 ( .A(in[954]), .B(n8395), .Z(n6587) );
  NAND U2217 ( .A(n6410), .B(n6194), .Z(n6195) );
  XNOR U2218 ( .A(n6587), .B(n6195), .Z(out[1149]) );
  XOR U2219 ( .A(in[585]), .B(n8459), .Z(n7387) );
  XOR U2220 ( .A(in[240]), .B(n8556), .Z(n7900) );
  XNOR U2221 ( .A(in[1460]), .B(n8597), .Z(n7897) );
  NAND U2222 ( .A(n7900), .B(n7897), .Z(n6196) );
  XNOR U2223 ( .A(n7387), .B(n6196), .Z(out[114]) );
  XNOR U2224 ( .A(in[955]), .B(n8399), .Z(n6591) );
  NAND U2225 ( .A(n6412), .B(n6197), .Z(n6198) );
  XNOR U2226 ( .A(n6591), .B(n6198), .Z(out[1150]) );
  XNOR U2227 ( .A(in[956]), .B(n8403), .Z(n6595) );
  NAND U2228 ( .A(n6414), .B(n6199), .Z(n6200) );
  XNOR U2229 ( .A(n6595), .B(n6200), .Z(out[1151]) );
  XNOR U2230 ( .A(n6202), .B(n6201), .Z(n8743) );
  XNOR U2231 ( .A(in[1004]), .B(n8743), .Z(n9436) );
  NAND U2232 ( .A(n6416), .B(n6203), .Z(n6204) );
  XNOR U2233 ( .A(n9436), .B(n6204), .Z(out[1152]) );
  XNOR U2234 ( .A(n6206), .B(n6205), .Z(n8745) );
  XNOR U2235 ( .A(in[1005]), .B(n8745), .Z(n9440) );
  NAND U2236 ( .A(n6418), .B(n6207), .Z(n6208) );
  XNOR U2237 ( .A(n9440), .B(n6208), .Z(out[1153]) );
  XNOR U2238 ( .A(n6210), .B(n6209), .Z(n8747) );
  XNOR U2239 ( .A(in[1006]), .B(n8747), .Z(n9444) );
  NAND U2240 ( .A(n6420), .B(n6211), .Z(n6212) );
  XNOR U2241 ( .A(n9444), .B(n6212), .Z(out[1154]) );
  XNOR U2242 ( .A(n6214), .B(n6213), .Z(n8749) );
  XNOR U2243 ( .A(in[1007]), .B(n8749), .Z(n9448) );
  NAND U2244 ( .A(n6422), .B(n6215), .Z(n6216) );
  XNOR U2245 ( .A(n9448), .B(n6216), .Z(out[1155]) );
  XNOR U2246 ( .A(n6218), .B(n6217), .Z(n8755) );
  XNOR U2247 ( .A(in[1008]), .B(n8755), .Z(n9452) );
  NAND U2248 ( .A(n6425), .B(n6219), .Z(n6220) );
  XNOR U2249 ( .A(n9452), .B(n6220), .Z(out[1156]) );
  XNOR U2250 ( .A(n6222), .B(n6221), .Z(n8757) );
  XNOR U2251 ( .A(in[1009]), .B(n8757), .Z(n9456) );
  NAND U2252 ( .A(n6427), .B(n6223), .Z(n6224) );
  XNOR U2253 ( .A(n9456), .B(n6224), .Z(out[1157]) );
  XNOR U2254 ( .A(n6226), .B(n6225), .Z(n8759) );
  XNOR U2255 ( .A(in[1010]), .B(n8759), .Z(n9460) );
  NAND U2256 ( .A(n6429), .B(n6227), .Z(n6228) );
  XNOR U2257 ( .A(n9460), .B(n6228), .Z(out[1158]) );
  XNOR U2258 ( .A(n6230), .B(n6229), .Z(n8761) );
  XNOR U2259 ( .A(in[1011]), .B(n8761), .Z(n9464) );
  NAND U2260 ( .A(n6431), .B(n6231), .Z(n6232) );
  XNOR U2261 ( .A(n9464), .B(n6232), .Z(out[1159]) );
  XOR U2262 ( .A(in[586]), .B(n8463), .Z(n7389) );
  XOR U2263 ( .A(in[241]), .B(n8564), .Z(n7924) );
  XNOR U2264 ( .A(in[1461]), .B(n8601), .Z(n7921) );
  NAND U2265 ( .A(n7924), .B(n7921), .Z(n6233) );
  XNOR U2266 ( .A(n7389), .B(n6233), .Z(out[115]) );
  XNOR U2267 ( .A(n6235), .B(n6234), .Z(n8763) );
  XNOR U2268 ( .A(in[1012]), .B(n8763), .Z(n9468) );
  NAND U2269 ( .A(n6433), .B(n6236), .Z(n6237) );
  XNOR U2270 ( .A(n9468), .B(n6237), .Z(out[1160]) );
  XNOR U2271 ( .A(n6239), .B(n6238), .Z(n8765) );
  XNOR U2272 ( .A(in[1013]), .B(n8765), .Z(n9472) );
  NAND U2273 ( .A(n6435), .B(n6240), .Z(n6241) );
  XNOR U2274 ( .A(n9472), .B(n6241), .Z(out[1161]) );
  XNOR U2275 ( .A(n6243), .B(n6242), .Z(n8767) );
  XNOR U2276 ( .A(in[1014]), .B(n8767), .Z(n9480) );
  NAND U2277 ( .A(n6437), .B(n6244), .Z(n6245) );
  XNOR U2278 ( .A(n9480), .B(n6245), .Z(out[1162]) );
  XNOR U2279 ( .A(n6247), .B(n6246), .Z(n8769) );
  XNOR U2280 ( .A(in[1015]), .B(n8769), .Z(n9484) );
  NAND U2281 ( .A(n6439), .B(n6248), .Z(n6249) );
  XNOR U2282 ( .A(n9484), .B(n6249), .Z(out[1163]) );
  XNOR U2283 ( .A(n6251), .B(n6250), .Z(n8625) );
  XNOR U2284 ( .A(in[1016]), .B(n8625), .Z(n9488) );
  NAND U2285 ( .A(n6441), .B(n6252), .Z(n6253) );
  XNOR U2286 ( .A(n9488), .B(n6253), .Z(out[1164]) );
  XNOR U2287 ( .A(n6255), .B(n6254), .Z(n8627) );
  XNOR U2288 ( .A(in[1017]), .B(n8627), .Z(n9492) );
  NAND U2289 ( .A(n6443), .B(n6256), .Z(n6257) );
  XNOR U2290 ( .A(n9492), .B(n6257), .Z(out[1165]) );
  XNOR U2291 ( .A(n6259), .B(n6258), .Z(n8629) );
  XNOR U2292 ( .A(in[1018]), .B(n8629), .Z(n9496) );
  NAND U2293 ( .A(n6446), .B(n6260), .Z(n6261) );
  XNOR U2294 ( .A(n9496), .B(n6261), .Z(out[1166]) );
  XNOR U2295 ( .A(n6263), .B(n6262), .Z(n8631) );
  XNOR U2296 ( .A(in[1019]), .B(n8631), .Z(n9500) );
  NAND U2297 ( .A(n6448), .B(n6264), .Z(n6265) );
  XNOR U2298 ( .A(n9500), .B(n6265), .Z(out[1167]) );
  XOR U2299 ( .A(n6267), .B(n6266), .Z(n8633) );
  XNOR U2300 ( .A(in[1020]), .B(n8633), .Z(n9504) );
  NAND U2301 ( .A(n6450), .B(n6268), .Z(n6269) );
  XNOR U2302 ( .A(n9504), .B(n6269), .Z(out[1168]) );
  XOR U2303 ( .A(n6271), .B(n6270), .Z(n8635) );
  XNOR U2304 ( .A(in[1021]), .B(n8635), .Z(n9508) );
  NAND U2305 ( .A(n6452), .B(n6272), .Z(n6273) );
  XNOR U2306 ( .A(n9508), .B(n6273), .Z(out[1169]) );
  XOR U2307 ( .A(in[587]), .B(n8467), .Z(n7391) );
  XOR U2308 ( .A(in[242]), .B(n8568), .Z(n7948) );
  XNOR U2309 ( .A(in[1462]), .B(n8611), .Z(n7945) );
  NAND U2310 ( .A(n7948), .B(n7945), .Z(n6274) );
  XNOR U2311 ( .A(n7391), .B(n6274), .Z(out[116]) );
  XOR U2312 ( .A(n6276), .B(n6275), .Z(n8641) );
  XNOR U2313 ( .A(in[1022]), .B(n8641), .Z(n9512) );
  NAND U2314 ( .A(n6454), .B(n6277), .Z(n6278) );
  XNOR U2315 ( .A(n9512), .B(n6278), .Z(out[1170]) );
  XNOR U2316 ( .A(n6280), .B(n6279), .Z(n8643) );
  XNOR U2317 ( .A(in[1023]), .B(n8643), .Z(n9516) );
  NAND U2318 ( .A(n6456), .B(n6281), .Z(n6282) );
  XNOR U2319 ( .A(n9516), .B(n6282), .Z(out[1171]) );
  XOR U2320 ( .A(n6284), .B(n6283), .Z(n8645) );
  XNOR U2321 ( .A(in[960]), .B(n8645), .Z(n9524) );
  NAND U2322 ( .A(n6458), .B(n6285), .Z(n6286) );
  XNOR U2323 ( .A(n9524), .B(n6286), .Z(out[1172]) );
  XOR U2324 ( .A(n6288), .B(n6287), .Z(n8647) );
  XNOR U2325 ( .A(in[961]), .B(n8647), .Z(n9528) );
  NAND U2326 ( .A(n6460), .B(n6289), .Z(n6290) );
  XNOR U2327 ( .A(n9528), .B(n6290), .Z(out[1173]) );
  XOR U2328 ( .A(n6292), .B(n6291), .Z(n8649) );
  XNOR U2329 ( .A(in[962]), .B(n8649), .Z(n9532) );
  NAND U2330 ( .A(n6462), .B(n6293), .Z(n6294) );
  XNOR U2331 ( .A(n9532), .B(n6294), .Z(out[1174]) );
  XOR U2332 ( .A(n6296), .B(n6295), .Z(n8651) );
  XNOR U2333 ( .A(in[963]), .B(n8651), .Z(n9536) );
  NAND U2334 ( .A(n6464), .B(n6297), .Z(n6298) );
  XNOR U2335 ( .A(n9536), .B(n6298), .Z(out[1175]) );
  XOR U2336 ( .A(n6300), .B(n6299), .Z(n8653) );
  XNOR U2337 ( .A(in[964]), .B(n8653), .Z(n9540) );
  NAND U2338 ( .A(n6467), .B(n6301), .Z(n6302) );
  XNOR U2339 ( .A(n9540), .B(n6302), .Z(out[1176]) );
  XOR U2340 ( .A(n6304), .B(n6303), .Z(n8655) );
  XNOR U2341 ( .A(in[965]), .B(n8655), .Z(n9544) );
  NAND U2342 ( .A(n6469), .B(n6305), .Z(n6306) );
  XNOR U2343 ( .A(n9544), .B(n6306), .Z(out[1177]) );
  XOR U2344 ( .A(n6308), .B(n6307), .Z(n8657) );
  XNOR U2345 ( .A(in[966]), .B(n8657), .Z(n9548) );
  NAND U2346 ( .A(n6471), .B(n6309), .Z(n6310) );
  XNOR U2347 ( .A(n9548), .B(n6310), .Z(out[1178]) );
  XOR U2348 ( .A(n6312), .B(n6311), .Z(n8659) );
  XNOR U2349 ( .A(in[967]), .B(n8659), .Z(n9552) );
  NAND U2350 ( .A(n6473), .B(n6313), .Z(n6314) );
  XNOR U2351 ( .A(n9552), .B(n6314), .Z(out[1179]) );
  XOR U2352 ( .A(in[588]), .B(n8475), .Z(n7393) );
  XOR U2353 ( .A(in[243]), .B(n8572), .Z(n7972) );
  XNOR U2354 ( .A(in[1463]), .B(n8615), .Z(n7969) );
  NAND U2355 ( .A(n7972), .B(n7969), .Z(n6315) );
  XNOR U2356 ( .A(n7393), .B(n6315), .Z(out[117]) );
  XOR U2357 ( .A(n6317), .B(n6316), .Z(n8663) );
  XNOR U2358 ( .A(in[968]), .B(n8663), .Z(n9556) );
  NAND U2359 ( .A(n6475), .B(n6318), .Z(n6319) );
  XNOR U2360 ( .A(n9556), .B(n6319), .Z(out[1180]) );
  XOR U2361 ( .A(n6321), .B(n6320), .Z(n8665) );
  XNOR U2362 ( .A(in[969]), .B(n8665), .Z(n9560) );
  NAND U2363 ( .A(n6477), .B(n6322), .Z(n6323) );
  XNOR U2364 ( .A(n9560), .B(n6323), .Z(out[1181]) );
  XNOR U2365 ( .A(n6325), .B(n6324), .Z(n8667) );
  XNOR U2366 ( .A(in[970]), .B(n8667), .Z(n9568) );
  NAND U2367 ( .A(n6479), .B(n6326), .Z(n6327) );
  XNOR U2368 ( .A(n9568), .B(n6327), .Z(out[1182]) );
  XOR U2369 ( .A(n6329), .B(n6328), .Z(n8669) );
  XNOR U2370 ( .A(in[971]), .B(n8669), .Z(n9572) );
  NAND U2371 ( .A(n6481), .B(n6330), .Z(n6331) );
  XNOR U2372 ( .A(n9572), .B(n6331), .Z(out[1183]) );
  XOR U2373 ( .A(n6333), .B(n6332), .Z(n8671) );
  XNOR U2374 ( .A(in[972]), .B(n8671), .Z(n9576) );
  NAND U2375 ( .A(n6483), .B(n6334), .Z(n6335) );
  XNOR U2376 ( .A(n9576), .B(n6335), .Z(out[1184]) );
  XOR U2377 ( .A(n6337), .B(n6336), .Z(n8673) );
  XNOR U2378 ( .A(in[973]), .B(n8673), .Z(n9580) );
  NAND U2379 ( .A(n6485), .B(n6338), .Z(n6339) );
  XNOR U2380 ( .A(n9580), .B(n6339), .Z(out[1185]) );
  XNOR U2381 ( .A(n6341), .B(n6340), .Z(n8675) );
  XNOR U2382 ( .A(in[974]), .B(n8675), .Z(n9584) );
  NAND U2383 ( .A(n6488), .B(n6342), .Z(n6343) );
  XNOR U2384 ( .A(n9584), .B(n6343), .Z(out[1186]) );
  XNOR U2385 ( .A(n6345), .B(n6344), .Z(n8677) );
  XNOR U2386 ( .A(in[975]), .B(n8677), .Z(n9588) );
  NAND U2387 ( .A(n6490), .B(n6346), .Z(n6347) );
  XNOR U2388 ( .A(n9588), .B(n6347), .Z(out[1187]) );
  XNOR U2389 ( .A(n6349), .B(n6348), .Z(n8679) );
  XNOR U2390 ( .A(in[976]), .B(n8679), .Z(n9592) );
  NAND U2391 ( .A(n6492), .B(n6350), .Z(n6351) );
  XNOR U2392 ( .A(n9592), .B(n6351), .Z(out[1188]) );
  XOR U2393 ( .A(n6353), .B(n6352), .Z(n8681) );
  XNOR U2394 ( .A(in[977]), .B(n8681), .Z(n9596) );
  NAND U2395 ( .A(n6494), .B(n6354), .Z(n6355) );
  XNOR U2396 ( .A(n9596), .B(n6355), .Z(out[1189]) );
  XOR U2397 ( .A(in[589]), .B(n8479), .Z(n7395) );
  XOR U2398 ( .A(in[244]), .B(n8576), .Z(n7996) );
  XNOR U2399 ( .A(in[1464]), .B(n8619), .Z(n7993) );
  NAND U2400 ( .A(n7996), .B(n7993), .Z(n6356) );
  XNOR U2401 ( .A(n7395), .B(n6356), .Z(out[118]) );
  XOR U2402 ( .A(n6358), .B(n6357), .Z(n8685) );
  XNOR U2403 ( .A(in[978]), .B(n8685), .Z(n9600) );
  NAND U2404 ( .A(n6496), .B(n6359), .Z(n6360) );
  XNOR U2405 ( .A(n9600), .B(n6360), .Z(out[1190]) );
  XOR U2406 ( .A(n6362), .B(n6361), .Z(n8687) );
  XNOR U2407 ( .A(in[979]), .B(n8687), .Z(n9604) );
  NAND U2408 ( .A(n6498), .B(n6363), .Z(n6364) );
  XNOR U2409 ( .A(n9604), .B(n6364), .Z(out[1191]) );
  OR U2410 ( .A(n6501), .B(n6365), .Z(n6366) );
  XNOR U2411 ( .A(n6500), .B(n6366), .Z(out[1192]) );
  OR U2412 ( .A(n6505), .B(n6367), .Z(n6368) );
  XNOR U2413 ( .A(n6504), .B(n6368), .Z(out[1193]) );
  OR U2414 ( .A(n6509), .B(n6369), .Z(n6370) );
  XNOR U2415 ( .A(n6508), .B(n6370), .Z(out[1194]) );
  OR U2416 ( .A(n6513), .B(n6371), .Z(n6372) );
  XNOR U2417 ( .A(n6512), .B(n6372), .Z(out[1195]) );
  OR U2418 ( .A(n6518), .B(n6373), .Z(n6374) );
  XNOR U2419 ( .A(n6517), .B(n6374), .Z(out[1196]) );
  OR U2420 ( .A(n6522), .B(n6375), .Z(n6376) );
  XNOR U2421 ( .A(n6521), .B(n6376), .Z(out[1197]) );
  OR U2422 ( .A(n6526), .B(n6377), .Z(n6378) );
  XNOR U2423 ( .A(n6525), .B(n6378), .Z(out[1198]) );
  OR U2424 ( .A(n6530), .B(n6379), .Z(n6380) );
  XNOR U2425 ( .A(n6529), .B(n6380), .Z(out[1199]) );
  XOR U2426 ( .A(in[590]), .B(n8483), .Z(n7397) );
  XOR U2427 ( .A(in[245]), .B(n8580), .Z(n8020) );
  XNOR U2428 ( .A(in[1465]), .B(n8623), .Z(n8017) );
  NAND U2429 ( .A(n8020), .B(n8017), .Z(n6381) );
  XNOR U2430 ( .A(n7397), .B(n6381), .Z(out[119]) );
  XOR U2431 ( .A(in[201]), .B(n8388), .Z(n8752) );
  XNOR U2432 ( .A(in[1421]), .B(n8425), .Z(n8751) );
  XOR U2433 ( .A(in[1044]), .B(n8930), .Z(n7442) );
  NAND U2434 ( .A(n8751), .B(n7442), .Z(n6382) );
  XNOR U2435 ( .A(n8752), .B(n6382), .Z(out[11]) );
  OR U2436 ( .A(n6534), .B(n6383), .Z(n6384) );
  XNOR U2437 ( .A(n6533), .B(n6384), .Z(out[1200]) );
  OR U2438 ( .A(n6538), .B(n6385), .Z(n6386) );
  XNOR U2439 ( .A(n6537), .B(n6386), .Z(out[1201]) );
  OR U2440 ( .A(n6542), .B(n6387), .Z(n6388) );
  XNOR U2441 ( .A(n6541), .B(n6388), .Z(out[1202]) );
  OR U2442 ( .A(n6546), .B(n6389), .Z(n6390) );
  XNOR U2443 ( .A(n6545), .B(n6390), .Z(out[1203]) );
  OR U2444 ( .A(n6550), .B(n6391), .Z(n6392) );
  XNOR U2445 ( .A(n6549), .B(n6392), .Z(out[1204]) );
  OR U2446 ( .A(n6554), .B(n6393), .Z(n6394) );
  XNOR U2447 ( .A(n6553), .B(n6394), .Z(out[1205]) );
  OR U2448 ( .A(n6559), .B(n6395), .Z(n6396) );
  XNOR U2449 ( .A(n6558), .B(n6396), .Z(out[1206]) );
  OR U2450 ( .A(n6563), .B(n6397), .Z(n6398) );
  XNOR U2451 ( .A(n6562), .B(n6398), .Z(out[1207]) );
  OR U2452 ( .A(n6567), .B(n6399), .Z(n6400) );
  XNOR U2453 ( .A(n6566), .B(n6400), .Z(out[1208]) );
  OR U2454 ( .A(n6571), .B(n6401), .Z(n6402) );
  XNOR U2455 ( .A(n6570), .B(n6402), .Z(out[1209]) );
  XOR U2456 ( .A(in[591]), .B(n8487), .Z(n7399) );
  XOR U2457 ( .A(in[246]), .B(n8584), .Z(n8044) );
  XNOR U2458 ( .A(in[1466]), .B(n8345), .Z(n8041) );
  NAND U2459 ( .A(n8044), .B(n8041), .Z(n6403) );
  XNOR U2460 ( .A(n7399), .B(n6403), .Z(out[120]) );
  OR U2461 ( .A(n6575), .B(n6404), .Z(n6405) );
  XNOR U2462 ( .A(n6574), .B(n6405), .Z(out[1210]) );
  OR U2463 ( .A(n6579), .B(n6406), .Z(n6407) );
  XNOR U2464 ( .A(n6578), .B(n6407), .Z(out[1211]) );
  OR U2465 ( .A(n6583), .B(n6408), .Z(n6409) );
  XNOR U2466 ( .A(n6582), .B(n6409), .Z(out[1212]) );
  OR U2467 ( .A(n6587), .B(n6410), .Z(n6411) );
  XNOR U2468 ( .A(n6586), .B(n6411), .Z(out[1213]) );
  OR U2469 ( .A(n6591), .B(n6412), .Z(n6413) );
  XNOR U2470 ( .A(n6590), .B(n6413), .Z(out[1214]) );
  OR U2471 ( .A(n6595), .B(n6414), .Z(n6415) );
  XNOR U2472 ( .A(n6594), .B(n6415), .Z(out[1215]) );
  OR U2473 ( .A(n9436), .B(n6416), .Z(n6417) );
  XNOR U2474 ( .A(n9435), .B(n6417), .Z(out[1216]) );
  OR U2475 ( .A(n9440), .B(n6418), .Z(n6419) );
  XNOR U2476 ( .A(n9439), .B(n6419), .Z(out[1217]) );
  OR U2477 ( .A(n9444), .B(n6420), .Z(n6421) );
  XNOR U2478 ( .A(n9443), .B(n6421), .Z(out[1218]) );
  OR U2479 ( .A(n9448), .B(n6422), .Z(n6423) );
  XNOR U2480 ( .A(n9447), .B(n6423), .Z(out[1219]) );
  XOR U2481 ( .A(in[592]), .B(n8491), .Z(n7401) );
  XOR U2482 ( .A(in[247]), .B(n8588), .Z(n8076) );
  XNOR U2483 ( .A(in[1467]), .B(n8349), .Z(n8073) );
  NAND U2484 ( .A(n8076), .B(n8073), .Z(n6424) );
  XNOR U2485 ( .A(n7401), .B(n6424), .Z(out[121]) );
  OR U2486 ( .A(n9452), .B(n6425), .Z(n6426) );
  XNOR U2487 ( .A(n9451), .B(n6426), .Z(out[1220]) );
  OR U2488 ( .A(n9456), .B(n6427), .Z(n6428) );
  XNOR U2489 ( .A(n9455), .B(n6428), .Z(out[1221]) );
  OR U2490 ( .A(n9460), .B(n6429), .Z(n6430) );
  XNOR U2491 ( .A(n9459), .B(n6430), .Z(out[1222]) );
  OR U2492 ( .A(n9464), .B(n6431), .Z(n6432) );
  XNOR U2493 ( .A(n9463), .B(n6432), .Z(out[1223]) );
  OR U2494 ( .A(n9468), .B(n6433), .Z(n6434) );
  XNOR U2495 ( .A(n9467), .B(n6434), .Z(out[1224]) );
  OR U2496 ( .A(n9472), .B(n6435), .Z(n6436) );
  XNOR U2497 ( .A(n9471), .B(n6436), .Z(out[1225]) );
  OR U2498 ( .A(n9480), .B(n6437), .Z(n6438) );
  XNOR U2499 ( .A(n9479), .B(n6438), .Z(out[1226]) );
  OR U2500 ( .A(n9484), .B(n6439), .Z(n6440) );
  XNOR U2501 ( .A(n9483), .B(n6440), .Z(out[1227]) );
  OR U2502 ( .A(n9488), .B(n6441), .Z(n6442) );
  XNOR U2503 ( .A(n9487), .B(n6442), .Z(out[1228]) );
  OR U2504 ( .A(n9492), .B(n6443), .Z(n6444) );
  XNOR U2505 ( .A(n9491), .B(n6444), .Z(out[1229]) );
  XOR U2506 ( .A(in[593]), .B(n8495), .Z(n7404) );
  XOR U2507 ( .A(in[248]), .B(n8592), .Z(n8120) );
  XNOR U2508 ( .A(in[1468]), .B(n8353), .Z(n8117) );
  NAND U2509 ( .A(n8120), .B(n8117), .Z(n6445) );
  XNOR U2510 ( .A(n7404), .B(n6445), .Z(out[122]) );
  OR U2511 ( .A(n9496), .B(n6446), .Z(n6447) );
  XNOR U2512 ( .A(n9495), .B(n6447), .Z(out[1230]) );
  OR U2513 ( .A(n9500), .B(n6448), .Z(n6449) );
  XNOR U2514 ( .A(n9499), .B(n6449), .Z(out[1231]) );
  OR U2515 ( .A(n9504), .B(n6450), .Z(n6451) );
  XNOR U2516 ( .A(n9503), .B(n6451), .Z(out[1232]) );
  OR U2517 ( .A(n9508), .B(n6452), .Z(n6453) );
  XNOR U2518 ( .A(n9507), .B(n6453), .Z(out[1233]) );
  OR U2519 ( .A(n9512), .B(n6454), .Z(n6455) );
  XNOR U2520 ( .A(n9511), .B(n6455), .Z(out[1234]) );
  OR U2521 ( .A(n9516), .B(n6456), .Z(n6457) );
  XNOR U2522 ( .A(n9515), .B(n6457), .Z(out[1235]) );
  OR U2523 ( .A(n9524), .B(n6458), .Z(n6459) );
  XNOR U2524 ( .A(n9523), .B(n6459), .Z(out[1236]) );
  OR U2525 ( .A(n9528), .B(n6460), .Z(n6461) );
  XNOR U2526 ( .A(n9527), .B(n6461), .Z(out[1237]) );
  OR U2527 ( .A(n9532), .B(n6462), .Z(n6463) );
  XNOR U2528 ( .A(n9531), .B(n6463), .Z(out[1238]) );
  OR U2529 ( .A(n9536), .B(n6464), .Z(n6465) );
  XNOR U2530 ( .A(n9535), .B(n6465), .Z(out[1239]) );
  XOR U2531 ( .A(in[594]), .B(n8499), .Z(n7406) );
  XOR U2532 ( .A(in[249]), .B(n8596), .Z(n8164) );
  XNOR U2533 ( .A(in[1469]), .B(n8357), .Z(n8161) );
  NAND U2534 ( .A(n8164), .B(n8161), .Z(n6466) );
  XNOR U2535 ( .A(n7406), .B(n6466), .Z(out[123]) );
  OR U2536 ( .A(n9540), .B(n6467), .Z(n6468) );
  XNOR U2537 ( .A(n9539), .B(n6468), .Z(out[1240]) );
  OR U2538 ( .A(n9544), .B(n6469), .Z(n6470) );
  XNOR U2539 ( .A(n9543), .B(n6470), .Z(out[1241]) );
  OR U2540 ( .A(n9548), .B(n6471), .Z(n6472) );
  XNOR U2541 ( .A(n9547), .B(n6472), .Z(out[1242]) );
  OR U2542 ( .A(n9552), .B(n6473), .Z(n6474) );
  XNOR U2543 ( .A(n9551), .B(n6474), .Z(out[1243]) );
  OR U2544 ( .A(n9556), .B(n6475), .Z(n6476) );
  XNOR U2545 ( .A(n9555), .B(n6476), .Z(out[1244]) );
  OR U2546 ( .A(n9560), .B(n6477), .Z(n6478) );
  XNOR U2547 ( .A(n9559), .B(n6478), .Z(out[1245]) );
  OR U2548 ( .A(n9568), .B(n6479), .Z(n6480) );
  XNOR U2549 ( .A(n9567), .B(n6480), .Z(out[1246]) );
  OR U2550 ( .A(n9572), .B(n6481), .Z(n6482) );
  XNOR U2551 ( .A(n9571), .B(n6482), .Z(out[1247]) );
  OR U2552 ( .A(n9576), .B(n6483), .Z(n6484) );
  XNOR U2553 ( .A(n9575), .B(n6484), .Z(out[1248]) );
  OR U2554 ( .A(n9580), .B(n6485), .Z(n6486) );
  XNOR U2555 ( .A(n9579), .B(n6486), .Z(out[1249]) );
  XOR U2556 ( .A(in[595]), .B(n8503), .Z(n7408) );
  XOR U2557 ( .A(in[250]), .B(n8600), .Z(n8210) );
  XNOR U2558 ( .A(in[1470]), .B(n8361), .Z(n8207) );
  NAND U2559 ( .A(n8210), .B(n8207), .Z(n6487) );
  XNOR U2560 ( .A(n7408), .B(n6487), .Z(out[124]) );
  OR U2561 ( .A(n9584), .B(n6488), .Z(n6489) );
  XNOR U2562 ( .A(n9583), .B(n6489), .Z(out[1250]) );
  OR U2563 ( .A(n9588), .B(n6490), .Z(n6491) );
  XNOR U2564 ( .A(n9587), .B(n6491), .Z(out[1251]) );
  OR U2565 ( .A(n9592), .B(n6492), .Z(n6493) );
  XNOR U2566 ( .A(n9591), .B(n6493), .Z(out[1252]) );
  OR U2567 ( .A(n9596), .B(n6494), .Z(n6495) );
  XNOR U2568 ( .A(n9595), .B(n6495), .Z(out[1253]) );
  OR U2569 ( .A(n9600), .B(n6496), .Z(n6497) );
  XNOR U2570 ( .A(n9599), .B(n6497), .Z(out[1254]) );
  OR U2571 ( .A(n9604), .B(n6498), .Z(n6499) );
  XNOR U2572 ( .A(n9603), .B(n6499), .Z(out[1255]) );
  ANDN U2573 ( .B(n6501), .A(n6500), .Z(n6502) );
  XNOR U2574 ( .A(n6503), .B(n6502), .Z(out[1256]) );
  ANDN U2575 ( .B(n6505), .A(n6504), .Z(n6506) );
  XNOR U2576 ( .A(n6507), .B(n6506), .Z(out[1257]) );
  ANDN U2577 ( .B(n6509), .A(n6508), .Z(n6510) );
  XNOR U2578 ( .A(n6511), .B(n6510), .Z(out[1258]) );
  ANDN U2579 ( .B(n6513), .A(n6512), .Z(n6514) );
  XNOR U2580 ( .A(n6515), .B(n6514), .Z(out[1259]) );
  XOR U2581 ( .A(in[596]), .B(n8507), .Z(n7410) );
  XNOR U2582 ( .A(in[251]), .B(n8610), .Z(n8254) );
  XNOR U2583 ( .A(in[1471]), .B(n8365), .Z(n8251) );
  NAND U2584 ( .A(n8254), .B(n8251), .Z(n6516) );
  XNOR U2585 ( .A(n7410), .B(n6516), .Z(out[125]) );
  ANDN U2586 ( .B(n6518), .A(n6517), .Z(n6519) );
  XNOR U2587 ( .A(n6520), .B(n6519), .Z(out[1260]) );
  ANDN U2588 ( .B(n6522), .A(n6521), .Z(n6523) );
  XNOR U2589 ( .A(n6524), .B(n6523), .Z(out[1261]) );
  ANDN U2590 ( .B(n6526), .A(n6525), .Z(n6527) );
  XNOR U2591 ( .A(n6528), .B(n6527), .Z(out[1262]) );
  ANDN U2592 ( .B(n6530), .A(n6529), .Z(n6531) );
  XNOR U2593 ( .A(n6532), .B(n6531), .Z(out[1263]) );
  ANDN U2594 ( .B(n6534), .A(n6533), .Z(n6535) );
  XNOR U2595 ( .A(n6536), .B(n6535), .Z(out[1264]) );
  ANDN U2596 ( .B(n6538), .A(n6537), .Z(n6539) );
  XNOR U2597 ( .A(n6540), .B(n6539), .Z(out[1265]) );
  ANDN U2598 ( .B(n6542), .A(n6541), .Z(n6543) );
  XNOR U2599 ( .A(n6544), .B(n6543), .Z(out[1266]) );
  ANDN U2600 ( .B(n6546), .A(n6545), .Z(n6547) );
  XNOR U2601 ( .A(n6548), .B(n6547), .Z(out[1267]) );
  ANDN U2602 ( .B(n6550), .A(n6549), .Z(n6551) );
  XNOR U2603 ( .A(n6552), .B(n6551), .Z(out[1268]) );
  ANDN U2604 ( .B(n6554), .A(n6553), .Z(n6555) );
  XNOR U2605 ( .A(n6556), .B(n6555), .Z(out[1269]) );
  XOR U2606 ( .A(in[597]), .B(n8511), .Z(n7412) );
  XNOR U2607 ( .A(in[252]), .B(n8614), .Z(n8298) );
  XNOR U2608 ( .A(in[1408]), .B(n8369), .Z(n8295) );
  NAND U2609 ( .A(n8298), .B(n8295), .Z(n6557) );
  XNOR U2610 ( .A(n7412), .B(n6557), .Z(out[126]) );
  ANDN U2611 ( .B(n6559), .A(n6558), .Z(n6560) );
  XNOR U2612 ( .A(n6561), .B(n6560), .Z(out[1270]) );
  ANDN U2613 ( .B(n6563), .A(n6562), .Z(n6564) );
  XNOR U2614 ( .A(n6565), .B(n6564), .Z(out[1271]) );
  ANDN U2615 ( .B(n6567), .A(n6566), .Z(n6568) );
  XNOR U2616 ( .A(n6569), .B(n6568), .Z(out[1272]) );
  ANDN U2617 ( .B(n6571), .A(n6570), .Z(n6572) );
  XNOR U2618 ( .A(n6573), .B(n6572), .Z(out[1273]) );
  ANDN U2619 ( .B(n6575), .A(n6574), .Z(n6576) );
  XNOR U2620 ( .A(n6577), .B(n6576), .Z(out[1274]) );
  ANDN U2621 ( .B(n6579), .A(n6578), .Z(n6580) );
  XNOR U2622 ( .A(n6581), .B(n6580), .Z(out[1275]) );
  ANDN U2623 ( .B(n6583), .A(n6582), .Z(n6584) );
  XNOR U2624 ( .A(n6585), .B(n6584), .Z(out[1276]) );
  ANDN U2625 ( .B(n6587), .A(n6586), .Z(n6588) );
  XNOR U2626 ( .A(n6589), .B(n6588), .Z(out[1277]) );
  ANDN U2627 ( .B(n6591), .A(n6590), .Z(n6592) );
  XNOR U2628 ( .A(n6593), .B(n6592), .Z(out[1278]) );
  ANDN U2629 ( .B(n6595), .A(n6594), .Z(n6596) );
  XNOR U2630 ( .A(n6597), .B(n6596), .Z(out[1279]) );
  XOR U2631 ( .A(in[598]), .B(n8519), .Z(n7414) );
  XNOR U2632 ( .A(in[253]), .B(n8618), .Z(n8342) );
  XNOR U2633 ( .A(in[1409]), .B(n8373), .Z(n8339) );
  NAND U2634 ( .A(n8342), .B(n8339), .Z(n6598) );
  XNOR U2635 ( .A(n7414), .B(n6598), .Z(out[127]) );
  XNOR U2636 ( .A(in[50]), .B(n8759), .Z(n6741) );
  XOR U2637 ( .A(in[1536]), .B(n8419), .Z(n7013) );
  XNOR U2638 ( .A(in[1172]), .B(n8436), .Z(n7011) );
  NAND U2639 ( .A(n7013), .B(n7011), .Z(n6599) );
  XNOR U2640 ( .A(n6741), .B(n6599), .Z(out[1280]) );
  XNOR U2641 ( .A(in[51]), .B(n8761), .Z(n6743) );
  XOR U2642 ( .A(in[1537]), .B(n8423), .Z(n7018) );
  XNOR U2643 ( .A(in[1173]), .B(n8440), .Z(n7016) );
  NAND U2644 ( .A(n7018), .B(n7016), .Z(n6600) );
  XNOR U2645 ( .A(n6743), .B(n6600), .Z(out[1281]) );
  XNOR U2646 ( .A(in[52]), .B(n8763), .Z(n6746) );
  XOR U2647 ( .A(in[1538]), .B(n8431), .Z(n7024) );
  XNOR U2648 ( .A(in[1174]), .B(n8444), .Z(n7021) );
  NAND U2649 ( .A(n7024), .B(n7021), .Z(n6601) );
  XNOR U2650 ( .A(n6746), .B(n6601), .Z(out[1282]) );
  XNOR U2651 ( .A(in[53]), .B(n8765), .Z(n6748) );
  XOR U2652 ( .A(in[1539]), .B(n8435), .Z(n7027) );
  XNOR U2653 ( .A(in[1175]), .B(n8448), .Z(n7025) );
  NAND U2654 ( .A(n7027), .B(n7025), .Z(n6602) );
  XNOR U2655 ( .A(n6748), .B(n6602), .Z(out[1283]) );
  XNOR U2656 ( .A(in[54]), .B(n8767), .Z(n6750) );
  XNOR U2657 ( .A(in[1540]), .B(n8439), .Z(n7034) );
  XNOR U2658 ( .A(in[1176]), .B(n8452), .Z(n7031) );
  NAND U2659 ( .A(n7034), .B(n7031), .Z(n6603) );
  XNOR U2660 ( .A(n6750), .B(n6603), .Z(out[1284]) );
  XNOR U2661 ( .A(in[55]), .B(n8769), .Z(n6752) );
  XNOR U2662 ( .A(in[1541]), .B(n8443), .Z(n7038) );
  XNOR U2663 ( .A(in[1177]), .B(n8456), .Z(n7035) );
  NAND U2664 ( .A(n7038), .B(n7035), .Z(n6604) );
  XNOR U2665 ( .A(n6752), .B(n6604), .Z(out[1285]) );
  XNOR U2666 ( .A(in[56]), .B(n8625), .Z(n6754) );
  XNOR U2667 ( .A(in[1542]), .B(n8447), .Z(n7042) );
  XNOR U2668 ( .A(in[1178]), .B(n8460), .Z(n7039) );
  NAND U2669 ( .A(n7042), .B(n7039), .Z(n6605) );
  XNOR U2670 ( .A(n6754), .B(n6605), .Z(out[1286]) );
  XNOR U2671 ( .A(in[57]), .B(n8627), .Z(n6756) );
  XNOR U2672 ( .A(in[1543]), .B(n8451), .Z(n7045) );
  XNOR U2673 ( .A(in[1179]), .B(n8464), .Z(n7043) );
  NAND U2674 ( .A(n7045), .B(n7043), .Z(n6606) );
  XNOR U2675 ( .A(n6756), .B(n6606), .Z(out[1287]) );
  XNOR U2676 ( .A(in[58]), .B(n8629), .Z(n6758) );
  XNOR U2677 ( .A(in[1544]), .B(n8455), .Z(n7051) );
  XNOR U2678 ( .A(in[1180]), .B(n8468), .Z(n7048) );
  NAND U2679 ( .A(n7051), .B(n7048), .Z(n6607) );
  XNOR U2680 ( .A(n6758), .B(n6607), .Z(out[1288]) );
  XNOR U2681 ( .A(in[59]), .B(n8631), .Z(n6760) );
  XNOR U2682 ( .A(in[1545]), .B(n8459), .Z(n7055) );
  XNOR U2683 ( .A(in[1181]), .B(n8476), .Z(n7052) );
  NAND U2684 ( .A(n7055), .B(n7052), .Z(n6608) );
  XNOR U2685 ( .A(n6760), .B(n6608), .Z(out[1289]) );
  XNOR U2686 ( .A(in[665]), .B(n8699), .Z(n7417) );
  XNOR U2687 ( .A(in[599]), .B(n8523), .Z(n8386) );
  NAND U2688 ( .A(n8386), .B(n8384), .Z(n6609) );
  XNOR U2689 ( .A(n7417), .B(n6609), .Z(out[128]) );
  XNOR U2690 ( .A(in[60]), .B(n8633), .Z(n6762) );
  XNOR U2691 ( .A(in[1546]), .B(n8463), .Z(n7059) );
  XNOR U2692 ( .A(in[1182]), .B(n8480), .Z(n7056) );
  NAND U2693 ( .A(n7059), .B(n7056), .Z(n6610) );
  XNOR U2694 ( .A(n6762), .B(n6610), .Z(out[1290]) );
  XNOR U2695 ( .A(in[61]), .B(n8635), .Z(n6764) );
  XNOR U2696 ( .A(in[1547]), .B(n8467), .Z(n7063) );
  XNOR U2697 ( .A(in[1183]), .B(n8484), .Z(n7060) );
  NAND U2698 ( .A(n7063), .B(n7060), .Z(n6611) );
  XNOR U2699 ( .A(n6764), .B(n6611), .Z(out[1291]) );
  XNOR U2700 ( .A(in[62]), .B(n8641), .Z(n6767) );
  XNOR U2701 ( .A(in[1548]), .B(n8475), .Z(n7067) );
  XNOR U2702 ( .A(in[1184]), .B(n8488), .Z(n7064) );
  NAND U2703 ( .A(n7067), .B(n7064), .Z(n6612) );
  XNOR U2704 ( .A(n6767), .B(n6612), .Z(out[1292]) );
  XNOR U2705 ( .A(in[63]), .B(n8643), .Z(n6769) );
  XNOR U2706 ( .A(in[1549]), .B(n8479), .Z(n7071) );
  XNOR U2707 ( .A(in[1185]), .B(n8492), .Z(n7068) );
  NAND U2708 ( .A(n7071), .B(n7068), .Z(n6613) );
  XNOR U2709 ( .A(n6769), .B(n6613), .Z(out[1293]) );
  XNOR U2710 ( .A(in[0]), .B(n8645), .Z(n6771) );
  XNOR U2711 ( .A(in[1550]), .B(n8483), .Z(n7076) );
  XOR U2712 ( .A(n8496), .B(in[1186]), .Z(n7073) );
  NAND U2713 ( .A(n7076), .B(n7073), .Z(n6614) );
  XNOR U2714 ( .A(n6771), .B(n6614), .Z(out[1294]) );
  XNOR U2715 ( .A(in[1]), .B(n8647), .Z(n6773) );
  XNOR U2716 ( .A(in[1551]), .B(n8487), .Z(n7079) );
  XOR U2717 ( .A(n8500), .B(in[1187]), .Z(n7077) );
  NAND U2718 ( .A(n7079), .B(n7077), .Z(n6615) );
  XNOR U2719 ( .A(n6773), .B(n6615), .Z(out[1295]) );
  XNOR U2720 ( .A(in[2]), .B(n8649), .Z(n6775) );
  XNOR U2721 ( .A(in[1552]), .B(n8491), .Z(n7085) );
  XOR U2722 ( .A(n8504), .B(in[1188]), .Z(n7082) );
  NAND U2723 ( .A(n7085), .B(n7082), .Z(n6616) );
  XNOR U2724 ( .A(n6775), .B(n6616), .Z(out[1296]) );
  XNOR U2725 ( .A(in[3]), .B(n8651), .Z(n6777) );
  XNOR U2726 ( .A(in[1553]), .B(n8495), .Z(n7089) );
  XOR U2727 ( .A(n8508), .B(in[1189]), .Z(n7086) );
  NAND U2728 ( .A(n7089), .B(n7086), .Z(n6617) );
  XNOR U2729 ( .A(n6777), .B(n6617), .Z(out[1297]) );
  XNOR U2730 ( .A(in[4]), .B(n8653), .Z(n6779) );
  XNOR U2731 ( .A(in[1554]), .B(n8499), .Z(n7093) );
  XNOR U2732 ( .A(in[1190]), .B(n8512), .Z(n7090) );
  NAND U2733 ( .A(n7093), .B(n7090), .Z(n6618) );
  XNOR U2734 ( .A(n6779), .B(n6618), .Z(out[1298]) );
  XNOR U2735 ( .A(in[5]), .B(n8655), .Z(n6781) );
  XNOR U2736 ( .A(in[1555]), .B(n8503), .Z(n7097) );
  XNOR U2737 ( .A(in[1191]), .B(n8520), .Z(n7094) );
  NAND U2738 ( .A(n7097), .B(n7094), .Z(n6619) );
  XNOR U2739 ( .A(n6781), .B(n6619), .Z(out[1299]) );
  XNOR U2740 ( .A(in[666]), .B(n8701), .Z(n7419) );
  XNOR U2741 ( .A(in[600]), .B(n8527), .Z(n8430) );
  XOR U2742 ( .A(in[255]), .B(n8344), .Z(n8428) );
  NAND U2743 ( .A(n8430), .B(n8428), .Z(n6620) );
  XNOR U2744 ( .A(n7419), .B(n6620), .Z(out[129]) );
  XOR U2745 ( .A(in[202]), .B(n8392), .Z(n8778) );
  XNOR U2746 ( .A(in[1422]), .B(n8433), .Z(n8777) );
  XOR U2747 ( .A(in[1045]), .B(n8933), .Z(n7445) );
  NAND U2748 ( .A(n8777), .B(n7445), .Z(n6621) );
  XNOR U2749 ( .A(n8778), .B(n6621), .Z(out[12]) );
  XNOR U2750 ( .A(in[6]), .B(n8657), .Z(n6783) );
  XNOR U2751 ( .A(in[1556]), .B(n8507), .Z(n7101) );
  XNOR U2752 ( .A(in[1192]), .B(n8524), .Z(n7098) );
  NAND U2753 ( .A(n7101), .B(n7098), .Z(n6622) );
  XNOR U2754 ( .A(n6783), .B(n6622), .Z(out[1300]) );
  XNOR U2755 ( .A(in[7]), .B(n8659), .Z(n6785) );
  XNOR U2756 ( .A(in[1557]), .B(n8511), .Z(n7105) );
  XNOR U2757 ( .A(in[1193]), .B(n8528), .Z(n7102) );
  NAND U2758 ( .A(n7105), .B(n7102), .Z(n6623) );
  XNOR U2759 ( .A(n6785), .B(n6623), .Z(out[1301]) );
  XNOR U2760 ( .A(in[8]), .B(n8663), .Z(n6788) );
  XNOR U2761 ( .A(in[1558]), .B(n8519), .Z(n7109) );
  XNOR U2762 ( .A(in[1194]), .B(n8532), .Z(n7106) );
  NAND U2763 ( .A(n7109), .B(n7106), .Z(n6624) );
  XNOR U2764 ( .A(n6788), .B(n6624), .Z(out[1302]) );
  XNOR U2765 ( .A(in[9]), .B(n8665), .Z(n6790) );
  XNOR U2766 ( .A(in[1559]), .B(n8523), .Z(n7113) );
  XNOR U2767 ( .A(in[1195]), .B(n8536), .Z(n7110) );
  NAND U2768 ( .A(n7113), .B(n7110), .Z(n6625) );
  XNOR U2769 ( .A(n6790), .B(n6625), .Z(out[1303]) );
  XNOR U2770 ( .A(in[10]), .B(n8667), .Z(n6792) );
  XNOR U2771 ( .A(in[1560]), .B(n8527), .Z(n7118) );
  XNOR U2772 ( .A(in[1196]), .B(n8540), .Z(n7115) );
  NAND U2773 ( .A(n7118), .B(n7115), .Z(n6626) );
  XNOR U2774 ( .A(n6792), .B(n6626), .Z(out[1304]) );
  XNOR U2775 ( .A(in[11]), .B(n8669), .Z(n6794) );
  XNOR U2776 ( .A(in[1561]), .B(n8531), .Z(n7122) );
  XNOR U2777 ( .A(in[1197]), .B(n8544), .Z(n7119) );
  NAND U2778 ( .A(n7122), .B(n7119), .Z(n6627) );
  XNOR U2779 ( .A(n6794), .B(n6627), .Z(out[1305]) );
  XNOR U2780 ( .A(in[12]), .B(n8671), .Z(n6796) );
  XNOR U2781 ( .A(in[1562]), .B(n8535), .Z(n7126) );
  XNOR U2782 ( .A(in[1198]), .B(n8548), .Z(n7123) );
  NAND U2783 ( .A(n7126), .B(n7123), .Z(n6628) );
  XNOR U2784 ( .A(n6796), .B(n6628), .Z(out[1306]) );
  XNOR U2785 ( .A(in[13]), .B(n8673), .Z(n6798) );
  XNOR U2786 ( .A(in[1563]), .B(n8539), .Z(n7130) );
  XNOR U2787 ( .A(in[1199]), .B(n8552), .Z(n7127) );
  NAND U2788 ( .A(n7130), .B(n7127), .Z(n6629) );
  XNOR U2789 ( .A(n6798), .B(n6629), .Z(out[1307]) );
  XNOR U2790 ( .A(in[14]), .B(n8675), .Z(n6800) );
  XNOR U2791 ( .A(in[1564]), .B(n8543), .Z(n7134) );
  XNOR U2792 ( .A(in[1200]), .B(n8556), .Z(n7131) );
  NAND U2793 ( .A(n7134), .B(n7131), .Z(n6630) );
  XNOR U2794 ( .A(n6800), .B(n6630), .Z(out[1308]) );
  XNOR U2795 ( .A(in[15]), .B(n8677), .Z(n6802) );
  XNOR U2796 ( .A(in[1565]), .B(n8547), .Z(n7138) );
  XNOR U2797 ( .A(in[1201]), .B(n8564), .Z(n7135) );
  NAND U2798 ( .A(n7138), .B(n7135), .Z(n6631) );
  XNOR U2799 ( .A(n6802), .B(n6631), .Z(out[1309]) );
  XNOR U2800 ( .A(in[667]), .B(n8703), .Z(n7422) );
  XNOR U2801 ( .A(in[601]), .B(n8531), .Z(n8474) );
  XOR U2802 ( .A(in[192]), .B(n8348), .Z(n8471) );
  NAND U2803 ( .A(n8474), .B(n8471), .Z(n6632) );
  XNOR U2804 ( .A(n7422), .B(n6632), .Z(out[130]) );
  XNOR U2805 ( .A(in[16]), .B(n8679), .Z(n6804) );
  XNOR U2806 ( .A(in[1566]), .B(n8551), .Z(n7142) );
  XNOR U2807 ( .A(in[1202]), .B(n8568), .Z(n7139) );
  NAND U2808 ( .A(n7142), .B(n7139), .Z(n6633) );
  XNOR U2809 ( .A(n6804), .B(n6633), .Z(out[1310]) );
  XNOR U2810 ( .A(in[17]), .B(n8681), .Z(n6806) );
  XNOR U2811 ( .A(in[1567]), .B(n8555), .Z(n7145) );
  XNOR U2812 ( .A(in[1203]), .B(n8572), .Z(n7143) );
  NAND U2813 ( .A(n7145), .B(n7143), .Z(n6634) );
  XNOR U2814 ( .A(n6806), .B(n6634), .Z(out[1311]) );
  XNOR U2815 ( .A(in[18]), .B(n8685), .Z(n6809) );
  XNOR U2816 ( .A(in[1568]), .B(n8563), .Z(n7151) );
  XNOR U2817 ( .A(in[1204]), .B(n8576), .Z(n7148) );
  NAND U2818 ( .A(n7151), .B(n7148), .Z(n6635) );
  XNOR U2819 ( .A(n6809), .B(n6635), .Z(out[1312]) );
  XNOR U2820 ( .A(in[19]), .B(n8687), .Z(n6811) );
  XNOR U2821 ( .A(in[1569]), .B(n8567), .Z(n7155) );
  XNOR U2822 ( .A(in[1205]), .B(n8580), .Z(n7152) );
  NAND U2823 ( .A(n7155), .B(n7152), .Z(n6636) );
  XNOR U2824 ( .A(n6811), .B(n6636), .Z(out[1313]) );
  XNOR U2825 ( .A(in[20]), .B(n8689), .Z(n6813) );
  XNOR U2826 ( .A(in[1570]), .B(n8571), .Z(n7160) );
  XNOR U2827 ( .A(in[1206]), .B(n8584), .Z(n7157) );
  NAND U2828 ( .A(n7160), .B(n7157), .Z(n6637) );
  XNOR U2829 ( .A(n6813), .B(n6637), .Z(out[1314]) );
  XNOR U2830 ( .A(in[21]), .B(n8691), .Z(n6815) );
  XNOR U2831 ( .A(in[1571]), .B(n8575), .Z(n7164) );
  XNOR U2832 ( .A(in[1207]), .B(n8588), .Z(n7161) );
  NAND U2833 ( .A(n7164), .B(n7161), .Z(n6638) );
  XNOR U2834 ( .A(n6815), .B(n6638), .Z(out[1315]) );
  XNOR U2835 ( .A(in[22]), .B(n8693), .Z(n6817) );
  XNOR U2836 ( .A(in[1572]), .B(n8579), .Z(n7168) );
  XNOR U2837 ( .A(in[1208]), .B(n8592), .Z(n7165) );
  NAND U2838 ( .A(n7168), .B(n7165), .Z(n6639) );
  XNOR U2839 ( .A(n6817), .B(n6639), .Z(out[1316]) );
  XNOR U2840 ( .A(in[23]), .B(n8695), .Z(n6819) );
  XOR U2841 ( .A(in[1573]), .B(n8583), .Z(n7172) );
  XNOR U2842 ( .A(in[1209]), .B(n8596), .Z(n7169) );
  NAND U2843 ( .A(n7172), .B(n7169), .Z(n6640) );
  XNOR U2844 ( .A(n6819), .B(n6640), .Z(out[1317]) );
  XNOR U2845 ( .A(in[24]), .B(n8697), .Z(n6821) );
  XOR U2846 ( .A(in[1574]), .B(n8587), .Z(n7176) );
  XNOR U2847 ( .A(in[1210]), .B(n8600), .Z(n7173) );
  NAND U2848 ( .A(n7176), .B(n7173), .Z(n6641) );
  XNOR U2849 ( .A(n6821), .B(n6641), .Z(out[1318]) );
  XNOR U2850 ( .A(in[25]), .B(n8699), .Z(n6823) );
  XOR U2851 ( .A(in[1575]), .B(n8591), .Z(n7180) );
  XOR U2852 ( .A(in[1211]), .B(n8610), .Z(n7177) );
  NAND U2853 ( .A(n7180), .B(n7177), .Z(n6642) );
  XNOR U2854 ( .A(n6823), .B(n6642), .Z(out[1319]) );
  XNOR U2855 ( .A(in[668]), .B(n8707), .Z(n7424) );
  XNOR U2856 ( .A(in[602]), .B(n8535), .Z(n8518) );
  XOR U2857 ( .A(in[193]), .B(n8352), .Z(n8515) );
  NAND U2858 ( .A(n8518), .B(n8515), .Z(n6643) );
  XNOR U2859 ( .A(n7424), .B(n6643), .Z(out[131]) );
  XNOR U2860 ( .A(in[26]), .B(n8701), .Z(n6825) );
  XOR U2861 ( .A(in[1576]), .B(n8595), .Z(n7184) );
  XOR U2862 ( .A(in[1212]), .B(n8614), .Z(n7181) );
  NAND U2863 ( .A(n7184), .B(n7181), .Z(n6644) );
  XNOR U2864 ( .A(n6825), .B(n6644), .Z(out[1320]) );
  XNOR U2865 ( .A(in[27]), .B(n8703), .Z(n6827) );
  XOR U2866 ( .A(in[1577]), .B(n8599), .Z(n7188) );
  XOR U2867 ( .A(in[1213]), .B(n8618), .Z(n7185) );
  NAND U2868 ( .A(n7188), .B(n7185), .Z(n6645) );
  XNOR U2869 ( .A(n6827), .B(n6645), .Z(out[1321]) );
  XNOR U2870 ( .A(in[28]), .B(n8707), .Z(n6830) );
  XOR U2871 ( .A(in[1578]), .B(n8609), .Z(n7192) );
  XNOR U2872 ( .A(in[1214]), .B(n8622), .Z(n7189) );
  NAND U2873 ( .A(n7192), .B(n7189), .Z(n6646) );
  XNOR U2874 ( .A(n6830), .B(n6646), .Z(out[1322]) );
  XNOR U2875 ( .A(in[29]), .B(n8709), .Z(n6832) );
  XOR U2876 ( .A(in[1579]), .B(n8613), .Z(n7196) );
  XOR U2877 ( .A(in[1215]), .B(n8344), .Z(n7193) );
  NAND U2878 ( .A(n7196), .B(n7193), .Z(n6647) );
  XNOR U2879 ( .A(n6832), .B(n6647), .Z(out[1323]) );
  XNOR U2880 ( .A(in[30]), .B(n8711), .Z(n6834) );
  XOR U2881 ( .A(in[1580]), .B(n8617), .Z(n7201) );
  XOR U2882 ( .A(in[1152]), .B(n8348), .Z(n7198) );
  NAND U2883 ( .A(n7201), .B(n7198), .Z(n6648) );
  XNOR U2884 ( .A(n6834), .B(n6648), .Z(out[1324]) );
  XNOR U2885 ( .A(in[31]), .B(n8713), .Z(n6836) );
  XOR U2886 ( .A(in[1581]), .B(n8621), .Z(n7205) );
  XOR U2887 ( .A(in[1153]), .B(n8352), .Z(n7202) );
  NAND U2888 ( .A(n7205), .B(n7202), .Z(n6649) );
  XNOR U2889 ( .A(n6836), .B(n6649), .Z(out[1325]) );
  XNOR U2890 ( .A(in[32]), .B(n8715), .Z(n6838) );
  XOR U2891 ( .A(in[1582]), .B(n8343), .Z(n7209) );
  XOR U2892 ( .A(in[1154]), .B(n8356), .Z(n7206) );
  NAND U2893 ( .A(n7209), .B(n7206), .Z(n6650) );
  XNOR U2894 ( .A(n6838), .B(n6650), .Z(out[1326]) );
  XNOR U2895 ( .A(in[33]), .B(n8717), .Z(n6840) );
  XOR U2896 ( .A(in[1583]), .B(n8347), .Z(n7213) );
  XOR U2897 ( .A(in[1155]), .B(n8360), .Z(n7210) );
  NAND U2898 ( .A(n7213), .B(n7210), .Z(n6651) );
  XNOR U2899 ( .A(n6840), .B(n6651), .Z(out[1327]) );
  XNOR U2900 ( .A(in[34]), .B(n8719), .Z(n6842) );
  XOR U2901 ( .A(in[1584]), .B(n8351), .Z(n7217) );
  XOR U2902 ( .A(in[1156]), .B(n8364), .Z(n7214) );
  NAND U2903 ( .A(n7217), .B(n7214), .Z(n6652) );
  XNOR U2904 ( .A(n6842), .B(n6652), .Z(out[1328]) );
  XNOR U2905 ( .A(in[35]), .B(n8721), .Z(n6844) );
  XOR U2906 ( .A(in[1585]), .B(n8355), .Z(n7221) );
  XOR U2907 ( .A(in[1157]), .B(n8368), .Z(n7218) );
  NAND U2908 ( .A(n7221), .B(n7218), .Z(n6653) );
  XNOR U2909 ( .A(n6844), .B(n6653), .Z(out[1329]) );
  XNOR U2910 ( .A(in[669]), .B(n8709), .Z(n7427) );
  XNOR U2911 ( .A(in[603]), .B(n8539), .Z(n8562) );
  XOR U2912 ( .A(in[194]), .B(n8356), .Z(n8559) );
  NAND U2913 ( .A(n8562), .B(n8559), .Z(n6654) );
  XNOR U2914 ( .A(n7427), .B(n6654), .Z(out[132]) );
  XNOR U2915 ( .A(in[36]), .B(n8723), .Z(n6846) );
  XOR U2916 ( .A(in[1586]), .B(n8359), .Z(n7225) );
  XOR U2917 ( .A(in[1158]), .B(n8372), .Z(n7222) );
  NAND U2918 ( .A(n7225), .B(n7222), .Z(n6655) );
  XNOR U2919 ( .A(n6846), .B(n6655), .Z(out[1330]) );
  XNOR U2920 ( .A(in[37]), .B(n8725), .Z(n6848) );
  XOR U2921 ( .A(in[1587]), .B(n8363), .Z(n7229) );
  XOR U2922 ( .A(in[1159]), .B(n8376), .Z(n7226) );
  NAND U2923 ( .A(n7229), .B(n7226), .Z(n6656) );
  XNOR U2924 ( .A(n6848), .B(n6656), .Z(out[1331]) );
  XNOR U2925 ( .A(in[38]), .B(n8731), .Z(n6851) );
  XOR U2926 ( .A(in[1588]), .B(n8367), .Z(n7233) );
  XOR U2927 ( .A(in[1160]), .B(n8380), .Z(n7230) );
  NAND U2928 ( .A(n7233), .B(n7230), .Z(n6657) );
  XNOR U2929 ( .A(n6851), .B(n6657), .Z(out[1332]) );
  XNOR U2930 ( .A(in[39]), .B(n8733), .Z(n6853) );
  XOR U2931 ( .A(in[1589]), .B(n8371), .Z(n7237) );
  XOR U2932 ( .A(in[1161]), .B(n8388), .Z(n7234) );
  NAND U2933 ( .A(n7237), .B(n7234), .Z(n6658) );
  XNOR U2934 ( .A(n6853), .B(n6658), .Z(out[1333]) );
  XNOR U2935 ( .A(in[40]), .B(n8735), .Z(n6855) );
  XOR U2936 ( .A(in[1590]), .B(n8375), .Z(n7242) );
  XOR U2937 ( .A(in[1162]), .B(n8392), .Z(n7239) );
  NAND U2938 ( .A(n7242), .B(n7239), .Z(n6659) );
  XNOR U2939 ( .A(n6855), .B(n6659), .Z(out[1334]) );
  XNOR U2940 ( .A(in[41]), .B(n8737), .Z(n6857) );
  XOR U2941 ( .A(in[1591]), .B(n8379), .Z(n7246) );
  XOR U2942 ( .A(in[1163]), .B(n8396), .Z(n7243) );
  NAND U2943 ( .A(n7246), .B(n7243), .Z(n6660) );
  XNOR U2944 ( .A(n6857), .B(n6660), .Z(out[1335]) );
  XNOR U2945 ( .A(in[42]), .B(n8739), .Z(n6859) );
  XOR U2946 ( .A(in[1592]), .B(n8387), .Z(n7250) );
  XOR U2947 ( .A(in[1164]), .B(n8400), .Z(n7247) );
  NAND U2948 ( .A(n7250), .B(n7247), .Z(n6661) );
  XNOR U2949 ( .A(n6859), .B(n6661), .Z(out[1336]) );
  XNOR U2950 ( .A(in[43]), .B(n8741), .Z(n6861) );
  XOR U2951 ( .A(in[1593]), .B(n8391), .Z(n7254) );
  XOR U2952 ( .A(in[1165]), .B(n8404), .Z(n7251) );
  NAND U2953 ( .A(n7254), .B(n7251), .Z(n6662) );
  XNOR U2954 ( .A(n6861), .B(n6662), .Z(out[1337]) );
  XNOR U2955 ( .A(in[44]), .B(n8743), .Z(n6863) );
  XOR U2956 ( .A(in[1594]), .B(n8395), .Z(n7258) );
  XOR U2957 ( .A(in[1166]), .B(n8408), .Z(n7255) );
  NAND U2958 ( .A(n7258), .B(n7255), .Z(n6663) );
  XNOR U2959 ( .A(n6863), .B(n6663), .Z(out[1338]) );
  XNOR U2960 ( .A(in[45]), .B(n8745), .Z(n6865) );
  XOR U2961 ( .A(in[1595]), .B(n8399), .Z(n7262) );
  XOR U2962 ( .A(in[1167]), .B(n8412), .Z(n7259) );
  NAND U2963 ( .A(n7262), .B(n7259), .Z(n6664) );
  XNOR U2964 ( .A(n6865), .B(n6664), .Z(out[1339]) );
  XNOR U2965 ( .A(in[670]), .B(n8711), .Z(n7429) );
  XNOR U2966 ( .A(in[604]), .B(n8543), .Z(n8606) );
  XOR U2967 ( .A(in[195]), .B(n8360), .Z(n8603) );
  NAND U2968 ( .A(n8606), .B(n8603), .Z(n6665) );
  XNOR U2969 ( .A(n7429), .B(n6665), .Z(out[133]) );
  XNOR U2970 ( .A(in[46]), .B(n8747), .Z(n6867) );
  XOR U2971 ( .A(in[1596]), .B(n8403), .Z(n7266) );
  XOR U2972 ( .A(in[1168]), .B(n8416), .Z(n7263) );
  NAND U2973 ( .A(n7266), .B(n7263), .Z(n6666) );
  XNOR U2974 ( .A(n6867), .B(n6666), .Z(out[1340]) );
  XNOR U2975 ( .A(in[47]), .B(n8749), .Z(n6869) );
  XOR U2976 ( .A(in[1597]), .B(n8407), .Z(n7270) );
  XOR U2977 ( .A(in[1169]), .B(n8420), .Z(n7267) );
  NAND U2978 ( .A(n7270), .B(n7267), .Z(n6667) );
  XNOR U2979 ( .A(n6869), .B(n6667), .Z(out[1341]) );
  XNOR U2980 ( .A(in[48]), .B(n8755), .Z(n6872) );
  XOR U2981 ( .A(in[1598]), .B(n8411), .Z(n7274) );
  XOR U2982 ( .A(in[1170]), .B(n8424), .Z(n7271) );
  NAND U2983 ( .A(n7274), .B(n7271), .Z(n6668) );
  XNOR U2984 ( .A(n6872), .B(n6668), .Z(out[1342]) );
  XNOR U2985 ( .A(in[49]), .B(n8757), .Z(n6874) );
  XOR U2986 ( .A(in[1599]), .B(n8415), .Z(n7277) );
  XNOR U2987 ( .A(in[1171]), .B(n8432), .Z(n7275) );
  NAND U2988 ( .A(n7277), .B(n7275), .Z(n6669) );
  XNOR U2989 ( .A(n6874), .B(n6669), .Z(out[1343]) );
  XOR U2990 ( .A(in[427]), .B(n8787), .Z(n6876) );
  NOR U2991 ( .A(n6741), .B(n7013), .Z(n6670) );
  XNOR U2992 ( .A(n6876), .B(n6670), .Z(out[1344]) );
  XOR U2993 ( .A(in[428]), .B(n8790), .Z(n6878) );
  NOR U2994 ( .A(n6743), .B(n7018), .Z(n6671) );
  XNOR U2995 ( .A(n6878), .B(n6671), .Z(out[1345]) );
  XOR U2996 ( .A(in[429]), .B(n8793), .Z(n6880) );
  NOR U2997 ( .A(n6746), .B(n7024), .Z(n6672) );
  XNOR U2998 ( .A(n6880), .B(n6672), .Z(out[1346]) );
  XOR U2999 ( .A(in[430]), .B(n8796), .Z(n6882) );
  NOR U3000 ( .A(n6748), .B(n7027), .Z(n6673) );
  XNOR U3001 ( .A(n6882), .B(n6673), .Z(out[1347]) );
  XOR U3002 ( .A(in[431]), .B(n8799), .Z(n6884) );
  NOR U3003 ( .A(n6750), .B(n7034), .Z(n6674) );
  XNOR U3004 ( .A(n6884), .B(n6674), .Z(out[1348]) );
  XOR U3005 ( .A(in[432]), .B(n8802), .Z(n6886) );
  NOR U3006 ( .A(n6752), .B(n7038), .Z(n6675) );
  XNOR U3007 ( .A(n6886), .B(n6675), .Z(out[1349]) );
  XNOR U3008 ( .A(in[671]), .B(n8713), .Z(n7431) );
  XNOR U3009 ( .A(in[605]), .B(n8547), .Z(n8640) );
  XOR U3010 ( .A(in[196]), .B(n8364), .Z(n8637) );
  NAND U3011 ( .A(n8640), .B(n8637), .Z(n6676) );
  XNOR U3012 ( .A(n7431), .B(n6676), .Z(out[134]) );
  XOR U3013 ( .A(in[433]), .B(n8805), .Z(n6888) );
  NOR U3014 ( .A(n6754), .B(n7042), .Z(n6677) );
  XNOR U3015 ( .A(n6888), .B(n6677), .Z(out[1350]) );
  XOR U3016 ( .A(in[434]), .B(n8808), .Z(n6890) );
  NOR U3017 ( .A(n6756), .B(n7045), .Z(n6678) );
  XNOR U3018 ( .A(n6890), .B(n6678), .Z(out[1351]) );
  XOR U3019 ( .A(in[435]), .B(n8815), .Z(n6893) );
  NOR U3020 ( .A(n6758), .B(n7051), .Z(n6679) );
  XNOR U3021 ( .A(n6893), .B(n6679), .Z(out[1352]) );
  XOR U3022 ( .A(in[436]), .B(n8818), .Z(n6895) );
  NOR U3023 ( .A(n6760), .B(n7055), .Z(n6680) );
  XNOR U3024 ( .A(n6895), .B(n6680), .Z(out[1353]) );
  XOR U3025 ( .A(in[437]), .B(n8821), .Z(n6897) );
  NOR U3026 ( .A(n6762), .B(n7059), .Z(n6681) );
  XNOR U3027 ( .A(n6897), .B(n6681), .Z(out[1354]) );
  XOR U3028 ( .A(in[438]), .B(n8824), .Z(n6899) );
  NOR U3029 ( .A(n6764), .B(n7063), .Z(n6682) );
  XNOR U3030 ( .A(n6899), .B(n6682), .Z(out[1355]) );
  XOR U3031 ( .A(in[439]), .B(n8827), .Z(n6901) );
  NOR U3032 ( .A(n6767), .B(n7067), .Z(n6683) );
  XNOR U3033 ( .A(n6901), .B(n6683), .Z(out[1356]) );
  XOR U3034 ( .A(in[440]), .B(n8830), .Z(n6903) );
  NOR U3035 ( .A(n6769), .B(n7071), .Z(n6684) );
  XNOR U3036 ( .A(n6903), .B(n6684), .Z(out[1357]) );
  XOR U3037 ( .A(in[441]), .B(n8833), .Z(n6905) );
  NOR U3038 ( .A(n6771), .B(n7076), .Z(n6685) );
  XNOR U3039 ( .A(n6905), .B(n6685), .Z(out[1358]) );
  XOR U3040 ( .A(in[442]), .B(n8836), .Z(n6907) );
  NOR U3041 ( .A(n6773), .B(n7079), .Z(n6686) );
  XNOR U3042 ( .A(n6907), .B(n6686), .Z(out[1359]) );
  XNOR U3043 ( .A(in[672]), .B(n8715), .Z(n7433) );
  XNOR U3044 ( .A(in[606]), .B(n8551), .Z(n8662) );
  XOR U3045 ( .A(in[197]), .B(n8368), .Z(n8886) );
  NAND U3046 ( .A(n8662), .B(n8886), .Z(n6687) );
  XNOR U3047 ( .A(n7433), .B(n6687), .Z(out[135]) );
  XOR U3048 ( .A(in[443]), .B(n8839), .Z(n6909) );
  NOR U3049 ( .A(n6775), .B(n7085), .Z(n6688) );
  XNOR U3050 ( .A(n6909), .B(n6688), .Z(out[1360]) );
  XOR U3051 ( .A(in[444]), .B(n8842), .Z(n6911) );
  NOR U3052 ( .A(n6777), .B(n7089), .Z(n6689) );
  XNOR U3053 ( .A(n6911), .B(n6689), .Z(out[1361]) );
  XOR U3054 ( .A(in[445]), .B(n8849), .Z(n6914) );
  NOR U3055 ( .A(n6779), .B(n7093), .Z(n6690) );
  XNOR U3056 ( .A(n6914), .B(n6690), .Z(out[1362]) );
  XOR U3057 ( .A(in[446]), .B(n8852), .Z(n6916) );
  NOR U3058 ( .A(n6781), .B(n7097), .Z(n6691) );
  XNOR U3059 ( .A(n6916), .B(n6691), .Z(out[1363]) );
  XOR U3060 ( .A(in[447]), .B(n8855), .Z(n6918) );
  NOR U3061 ( .A(n6783), .B(n7101), .Z(n6692) );
  XNOR U3062 ( .A(n6918), .B(n6692), .Z(out[1364]) );
  XOR U3063 ( .A(in[384]), .B(n8858), .Z(n6920) );
  NOR U3064 ( .A(n6785), .B(n7105), .Z(n6693) );
  XNOR U3065 ( .A(n6920), .B(n6693), .Z(out[1365]) );
  XOR U3066 ( .A(in[385]), .B(n8861), .Z(n6922) );
  NOR U3067 ( .A(n6788), .B(n7109), .Z(n6694) );
  XNOR U3068 ( .A(n6922), .B(n6694), .Z(out[1366]) );
  XOR U3069 ( .A(in[386]), .B(n8864), .Z(n6924) );
  NOR U3070 ( .A(n6790), .B(n7113), .Z(n6695) );
  XNOR U3071 ( .A(n6924), .B(n6695), .Z(out[1367]) );
  XOR U3072 ( .A(in[387]), .B(n8867), .Z(n6926) );
  NOR U3073 ( .A(n6792), .B(n7118), .Z(n6696) );
  XNOR U3074 ( .A(n6926), .B(n6696), .Z(out[1368]) );
  XOR U3075 ( .A(in[388]), .B(n8870), .Z(n6928) );
  NOR U3076 ( .A(n6794), .B(n7122), .Z(n6697) );
  XNOR U3077 ( .A(n6928), .B(n6697), .Z(out[1369]) );
  XNOR U3078 ( .A(in[673]), .B(n8717), .Z(n7435) );
  XNOR U3079 ( .A(in[607]), .B(n8555), .Z(n8684) );
  XOR U3080 ( .A(in[198]), .B(n8372), .Z(n9170) );
  NAND U3081 ( .A(n8684), .B(n9170), .Z(n6698) );
  XNOR U3082 ( .A(n7435), .B(n6698), .Z(out[136]) );
  XOR U3083 ( .A(in[389]), .B(n8873), .Z(n6930) );
  NOR U3084 ( .A(n6796), .B(n7126), .Z(n6699) );
  XNOR U3085 ( .A(n6930), .B(n6699), .Z(out[1370]) );
  XOR U3086 ( .A(in[390]), .B(n8876), .Z(n6932) );
  NOR U3087 ( .A(n6798), .B(n7130), .Z(n6700) );
  XNOR U3088 ( .A(n6932), .B(n6700), .Z(out[1371]) );
  XOR U3089 ( .A(in[391]), .B(n8887), .Z(n6936) );
  NOR U3090 ( .A(n6800), .B(n7134), .Z(n6701) );
  XNOR U3091 ( .A(n6936), .B(n6701), .Z(out[1372]) );
  XOR U3092 ( .A(in[392]), .B(n8890), .Z(n6938) );
  NOR U3093 ( .A(n6802), .B(n7138), .Z(n6702) );
  XNOR U3094 ( .A(n6938), .B(n6702), .Z(out[1373]) );
  XOR U3095 ( .A(in[393]), .B(n8893), .Z(n6940) );
  NOR U3096 ( .A(n6804), .B(n7142), .Z(n6703) );
  XNOR U3097 ( .A(n6940), .B(n6703), .Z(out[1374]) );
  XOR U3098 ( .A(in[394]), .B(n8896), .Z(n6942) );
  NOR U3099 ( .A(n6806), .B(n7145), .Z(n6704) );
  XNOR U3100 ( .A(n6942), .B(n6704), .Z(out[1375]) );
  XOR U3101 ( .A(in[395]), .B(n8899), .Z(n6944) );
  NOR U3102 ( .A(n6809), .B(n7151), .Z(n6705) );
  XNOR U3103 ( .A(n6944), .B(n6705), .Z(out[1376]) );
  XNOR U3104 ( .A(n8902), .B(in[396]), .Z(n6946) );
  NOR U3105 ( .A(n6811), .B(n7155), .Z(n6706) );
  XNOR U3106 ( .A(n6946), .B(n6706), .Z(out[1377]) );
  XNOR U3107 ( .A(n8905), .B(in[397]), .Z(n6948) );
  NOR U3108 ( .A(n6813), .B(n7160), .Z(n6707) );
  XNOR U3109 ( .A(n6948), .B(n6707), .Z(out[1378]) );
  XNOR U3110 ( .A(n8908), .B(in[398]), .Z(n6950) );
  NOR U3111 ( .A(n6815), .B(n7164), .Z(n6708) );
  XNOR U3112 ( .A(n6950), .B(n6708), .Z(out[1379]) );
  XNOR U3113 ( .A(in[674]), .B(n8719), .Z(n7437) );
  XNOR U3114 ( .A(in[608]), .B(n8563), .Z(n8706) );
  XOR U3115 ( .A(in[199]), .B(n8376), .Z(n9614) );
  NAND U3116 ( .A(n8706), .B(n9614), .Z(n6709) );
  XNOR U3117 ( .A(n7437), .B(n6709), .Z(out[137]) );
  XNOR U3118 ( .A(n8911), .B(in[399]), .Z(n6952) );
  NOR U3119 ( .A(n6817), .B(n7168), .Z(n6710) );
  XNOR U3120 ( .A(n6952), .B(n6710), .Z(out[1380]) );
  XNOR U3121 ( .A(n8914), .B(in[400]), .Z(n6954) );
  NOR U3122 ( .A(n6819), .B(n7172), .Z(n6711) );
  XNOR U3123 ( .A(n6954), .B(n6711), .Z(out[1381]) );
  XNOR U3124 ( .A(n8921), .B(in[401]), .Z(n6957) );
  NOR U3125 ( .A(n6821), .B(n7176), .Z(n6712) );
  XNOR U3126 ( .A(n6957), .B(n6712), .Z(out[1382]) );
  XNOR U3127 ( .A(n8924), .B(in[402]), .Z(n6959) );
  NOR U3128 ( .A(n6823), .B(n7180), .Z(n6713) );
  XNOR U3129 ( .A(n6959), .B(n6713), .Z(out[1383]) );
  XNOR U3130 ( .A(n8927), .B(in[403]), .Z(n6961) );
  NOR U3131 ( .A(n6825), .B(n7184), .Z(n6714) );
  XNOR U3132 ( .A(n6961), .B(n6714), .Z(out[1384]) );
  XNOR U3133 ( .A(in[404]), .B(n8930), .Z(n6963) );
  NOR U3134 ( .A(n6827), .B(n7188), .Z(n6715) );
  XNOR U3135 ( .A(n6963), .B(n6715), .Z(out[1385]) );
  XNOR U3136 ( .A(in[405]), .B(n8933), .Z(n6965) );
  NOR U3137 ( .A(n6830), .B(n7192), .Z(n6716) );
  XNOR U3138 ( .A(n6965), .B(n6716), .Z(out[1386]) );
  XNOR U3139 ( .A(in[406]), .B(n8936), .Z(n6967) );
  NOR U3140 ( .A(n6832), .B(n7196), .Z(n6717) );
  XNOR U3141 ( .A(n6967), .B(n6717), .Z(out[1387]) );
  XNOR U3142 ( .A(in[407]), .B(n8939), .Z(n6969) );
  NOR U3143 ( .A(n6834), .B(n7201), .Z(n6718) );
  XNOR U3144 ( .A(n6969), .B(n6718), .Z(out[1388]) );
  XNOR U3145 ( .A(in[408]), .B(n8942), .Z(n6971) );
  NOR U3146 ( .A(n6836), .B(n7205), .Z(n6719) );
  XNOR U3147 ( .A(n6971), .B(n6719), .Z(out[1389]) );
  XNOR U3148 ( .A(in[675]), .B(n8721), .Z(n7440) );
  XNOR U3149 ( .A(in[609]), .B(n8567), .Z(n8730) );
  NAND U3150 ( .A(n8730), .B(n8728), .Z(n6720) );
  XNOR U3151 ( .A(n7440), .B(n6720), .Z(out[138]) );
  XNOR U3152 ( .A(in[409]), .B(n8945), .Z(n6973) );
  NOR U3153 ( .A(n6838), .B(n7209), .Z(n6721) );
  XNOR U3154 ( .A(n6973), .B(n6721), .Z(out[1390]) );
  XNOR U3155 ( .A(in[410]), .B(n8948), .Z(n6975) );
  NOR U3156 ( .A(n6840), .B(n7213), .Z(n6722) );
  XNOR U3157 ( .A(n6975), .B(n6722), .Z(out[1391]) );
  XNOR U3158 ( .A(in[411]), .B(n8955), .Z(n6978) );
  NOR U3159 ( .A(n6842), .B(n7217), .Z(n6723) );
  XNOR U3160 ( .A(n6978), .B(n6723), .Z(out[1392]) );
  XNOR U3161 ( .A(in[412]), .B(n8958), .Z(n6980) );
  NOR U3162 ( .A(n6844), .B(n7221), .Z(n6724) );
  XNOR U3163 ( .A(n6980), .B(n6724), .Z(out[1393]) );
  XNOR U3164 ( .A(in[413]), .B(n8961), .Z(n6982) );
  NOR U3165 ( .A(n6846), .B(n7225), .Z(n6725) );
  XNOR U3166 ( .A(n6982), .B(n6725), .Z(out[1394]) );
  XNOR U3167 ( .A(in[414]), .B(n8964), .Z(n6984) );
  NOR U3168 ( .A(n6848), .B(n7229), .Z(n6726) );
  XNOR U3169 ( .A(n6984), .B(n6726), .Z(out[1395]) );
  XNOR U3170 ( .A(in[415]), .B(n8967), .Z(n6986) );
  NOR U3171 ( .A(n6851), .B(n7233), .Z(n6727) );
  XNOR U3172 ( .A(n6986), .B(n6727), .Z(out[1396]) );
  XNOR U3173 ( .A(in[416]), .B(n8970), .Z(n6988) );
  NOR U3174 ( .A(n6853), .B(n7237), .Z(n6728) );
  XNOR U3175 ( .A(n6988), .B(n6728), .Z(out[1397]) );
  XNOR U3176 ( .A(in[417]), .B(n8973), .Z(n6990) );
  NOR U3177 ( .A(n6855), .B(n7242), .Z(n6729) );
  XNOR U3178 ( .A(n6990), .B(n6729), .Z(out[1398]) );
  XNOR U3179 ( .A(in[418]), .B(n8976), .Z(n6992) );
  NOR U3180 ( .A(n6857), .B(n7246), .Z(n6730) );
  XNOR U3181 ( .A(n6992), .B(n6730), .Z(out[1399]) );
  XNOR U3182 ( .A(in[676]), .B(n8723), .Z(n7443) );
  XNOR U3183 ( .A(in[610]), .B(n8571), .Z(n8754) );
  NAND U3184 ( .A(n8754), .B(n8752), .Z(n6731) );
  XNOR U3185 ( .A(n7443), .B(n6731), .Z(out[139]) );
  XOR U3186 ( .A(in[203]), .B(n8396), .Z(n8812) );
  XNOR U3187 ( .A(in[1423]), .B(n8437), .Z(n8811) );
  XOR U3188 ( .A(in[1046]), .B(n8936), .Z(n7448) );
  NAND U3189 ( .A(n8811), .B(n7448), .Z(n6732) );
  XNOR U3190 ( .A(n8812), .B(n6732), .Z(out[13]) );
  XNOR U3191 ( .A(in[419]), .B(n8979), .Z(n6994) );
  NOR U3192 ( .A(n6859), .B(n7250), .Z(n6733) );
  XNOR U3193 ( .A(n6994), .B(n6733), .Z(out[1400]) );
  XOR U3194 ( .A(in[420]), .B(n8982), .Z(n6996) );
  NOR U3195 ( .A(n6861), .B(n7254), .Z(n6734) );
  XNOR U3196 ( .A(n6996), .B(n6734), .Z(out[1401]) );
  XOR U3197 ( .A(in[421]), .B(n8989), .Z(n6999) );
  NOR U3198 ( .A(n6863), .B(n7258), .Z(n6735) );
  XNOR U3199 ( .A(n6999), .B(n6735), .Z(out[1402]) );
  XOR U3200 ( .A(in[422]), .B(n8992), .Z(n7001) );
  NOR U3201 ( .A(n6865), .B(n7262), .Z(n6736) );
  XNOR U3202 ( .A(n7001), .B(n6736), .Z(out[1403]) );
  XOR U3203 ( .A(in[423]), .B(n8771), .Z(n7003) );
  NOR U3204 ( .A(n6867), .B(n7266), .Z(n6737) );
  XNOR U3205 ( .A(n7003), .B(n6737), .Z(out[1404]) );
  XOR U3206 ( .A(in[424]), .B(n8774), .Z(n7005) );
  NOR U3207 ( .A(n6869), .B(n7270), .Z(n6738) );
  XNOR U3208 ( .A(n7005), .B(n6738), .Z(out[1405]) );
  XOR U3209 ( .A(in[425]), .B(n8781), .Z(n7007) );
  NOR U3210 ( .A(n6872), .B(n7274), .Z(n6739) );
  XNOR U3211 ( .A(n7007), .B(n6739), .Z(out[1406]) );
  XOR U3212 ( .A(in[426]), .B(n8784), .Z(n7009) );
  NOR U3213 ( .A(n6874), .B(n7277), .Z(n6740) );
  XNOR U3214 ( .A(n7009), .B(n6740), .Z(out[1407]) );
  XOR U3215 ( .A(in[789]), .B(n8461), .Z(n7012) );
  NAND U3216 ( .A(n6876), .B(n6741), .Z(n6742) );
  XNOR U3217 ( .A(n7012), .B(n6742), .Z(out[1408]) );
  XOR U3218 ( .A(in[790]), .B(n8465), .Z(n7017) );
  NAND U3219 ( .A(n6878), .B(n6743), .Z(n6744) );
  XNOR U3220 ( .A(n7017), .B(n6744), .Z(out[1409]) );
  XNOR U3221 ( .A(in[677]), .B(n8725), .Z(n7446) );
  XNOR U3222 ( .A(in[611]), .B(n8575), .Z(n8780) );
  NAND U3223 ( .A(n8780), .B(n8778), .Z(n6745) );
  XNOR U3224 ( .A(n7446), .B(n6745), .Z(out[140]) );
  XOR U3225 ( .A(in[791]), .B(n8469), .Z(n7022) );
  NAND U3226 ( .A(n6880), .B(n6746), .Z(n6747) );
  XNOR U3227 ( .A(n7022), .B(n6747), .Z(out[1410]) );
  XOR U3228 ( .A(in[792]), .B(n8477), .Z(n7026) );
  NAND U3229 ( .A(n6882), .B(n6748), .Z(n6749) );
  XNOR U3230 ( .A(n7026), .B(n6749), .Z(out[1411]) );
  XOR U3231 ( .A(in[793]), .B(n8481), .Z(n7032) );
  NAND U3232 ( .A(n6884), .B(n6750), .Z(n6751) );
  XNOR U3233 ( .A(n7032), .B(n6751), .Z(out[1412]) );
  XOR U3234 ( .A(in[794]), .B(n8485), .Z(n7036) );
  NAND U3235 ( .A(n6886), .B(n6752), .Z(n6753) );
  XNOR U3236 ( .A(n7036), .B(n6753), .Z(out[1413]) );
  XOR U3237 ( .A(in[795]), .B(n8489), .Z(n7040) );
  NAND U3238 ( .A(n6888), .B(n6754), .Z(n6755) );
  XNOR U3239 ( .A(n7040), .B(n6755), .Z(out[1414]) );
  XOR U3240 ( .A(in[796]), .B(n8493), .Z(n7044) );
  NAND U3241 ( .A(n6890), .B(n6756), .Z(n6757) );
  XNOR U3242 ( .A(n7044), .B(n6757), .Z(out[1415]) );
  XOR U3243 ( .A(in[797]), .B(n8497), .Z(n7049) );
  NAND U3244 ( .A(n6893), .B(n6758), .Z(n6759) );
  XNOR U3245 ( .A(n7049), .B(n6759), .Z(out[1416]) );
  XOR U3246 ( .A(in[798]), .B(n8501), .Z(n7053) );
  NAND U3247 ( .A(n6895), .B(n6760), .Z(n6761) );
  XNOR U3248 ( .A(n7053), .B(n6761), .Z(out[1417]) );
  XOR U3249 ( .A(in[799]), .B(n8505), .Z(n7057) );
  NAND U3250 ( .A(n6897), .B(n6762), .Z(n6763) );
  XNOR U3251 ( .A(n7057), .B(n6763), .Z(out[1418]) );
  XOR U3252 ( .A(in[800]), .B(n8509), .Z(n7061) );
  NAND U3253 ( .A(n6899), .B(n6764), .Z(n6765) );
  XNOR U3254 ( .A(n7061), .B(n6765), .Z(out[1419]) );
  XNOR U3255 ( .A(in[678]), .B(n8731), .Z(n7449) );
  XNOR U3256 ( .A(in[612]), .B(n8579), .Z(n8814) );
  NAND U3257 ( .A(n8814), .B(n8812), .Z(n6766) );
  XNOR U3258 ( .A(n7449), .B(n6766), .Z(out[141]) );
  XOR U3259 ( .A(in[801]), .B(n8513), .Z(n7065) );
  NAND U3260 ( .A(n6901), .B(n6767), .Z(n6768) );
  XNOR U3261 ( .A(n7065), .B(n6768), .Z(out[1420]) );
  XOR U3262 ( .A(in[802]), .B(n8521), .Z(n7069) );
  NAND U3263 ( .A(n6903), .B(n6769), .Z(n6770) );
  XNOR U3264 ( .A(n7069), .B(n6770), .Z(out[1421]) );
  XOR U3265 ( .A(in[803]), .B(n8525), .Z(n7074) );
  NAND U3266 ( .A(n6905), .B(n6771), .Z(n6772) );
  XNOR U3267 ( .A(n7074), .B(n6772), .Z(out[1422]) );
  XOR U3268 ( .A(in[804]), .B(n8529), .Z(n7078) );
  NAND U3269 ( .A(n6907), .B(n6773), .Z(n6774) );
  XNOR U3270 ( .A(n7078), .B(n6774), .Z(out[1423]) );
  XOR U3271 ( .A(in[805]), .B(n8533), .Z(n7083) );
  NAND U3272 ( .A(n6909), .B(n6775), .Z(n6776) );
  XNOR U3273 ( .A(n7083), .B(n6776), .Z(out[1424]) );
  XNOR U3274 ( .A(in[806]), .B(n8537), .Z(n7087) );
  NAND U3275 ( .A(n6911), .B(n6777), .Z(n6778) );
  XNOR U3276 ( .A(n7087), .B(n6778), .Z(out[1425]) );
  XNOR U3277 ( .A(in[807]), .B(n8541), .Z(n7091) );
  NAND U3278 ( .A(n6914), .B(n6779), .Z(n6780) );
  XNOR U3279 ( .A(n7091), .B(n6780), .Z(out[1426]) );
  XNOR U3280 ( .A(in[808]), .B(n8545), .Z(n7095) );
  NAND U3281 ( .A(n6916), .B(n6781), .Z(n6782) );
  XNOR U3282 ( .A(n7095), .B(n6782), .Z(out[1427]) );
  XNOR U3283 ( .A(in[809]), .B(n8549), .Z(n7099) );
  NAND U3284 ( .A(n6918), .B(n6783), .Z(n6784) );
  XNOR U3285 ( .A(n7099), .B(n6784), .Z(out[1428]) );
  XNOR U3286 ( .A(in[810]), .B(n8553), .Z(n7103) );
  NAND U3287 ( .A(n6920), .B(n6785), .Z(n6786) );
  XNOR U3288 ( .A(n7103), .B(n6786), .Z(out[1429]) );
  XNOR U3289 ( .A(in[679]), .B(n8733), .Z(n7453) );
  XOR U3290 ( .A(in[613]), .B(n8583), .Z(n8848) );
  XOR U3291 ( .A(in[204]), .B(n8400), .Z(n8846) );
  NAND U3292 ( .A(n8848), .B(n8846), .Z(n6787) );
  XNOR U3293 ( .A(n7453), .B(n6787), .Z(out[142]) );
  XNOR U3294 ( .A(in[811]), .B(n8557), .Z(n7107) );
  NAND U3295 ( .A(n6922), .B(n6788), .Z(n6789) );
  XNOR U3296 ( .A(n7107), .B(n6789), .Z(out[1430]) );
  XNOR U3297 ( .A(in[812]), .B(n8565), .Z(n7111) );
  NAND U3298 ( .A(n6924), .B(n6790), .Z(n6791) );
  XNOR U3299 ( .A(n7111), .B(n6791), .Z(out[1431]) );
  XNOR U3300 ( .A(in[813]), .B(n8569), .Z(n7116) );
  NAND U3301 ( .A(n6926), .B(n6792), .Z(n6793) );
  XNOR U3302 ( .A(n7116), .B(n6793), .Z(out[1432]) );
  XNOR U3303 ( .A(in[814]), .B(n8573), .Z(n7120) );
  NAND U3304 ( .A(n6928), .B(n6794), .Z(n6795) );
  XNOR U3305 ( .A(n7120), .B(n6795), .Z(out[1433]) );
  XNOR U3306 ( .A(in[815]), .B(n8577), .Z(n7124) );
  NAND U3307 ( .A(n6930), .B(n6796), .Z(n6797) );
  XNOR U3308 ( .A(n7124), .B(n6797), .Z(out[1434]) );
  XNOR U3309 ( .A(in[816]), .B(n8581), .Z(n7128) );
  NAND U3310 ( .A(n6932), .B(n6798), .Z(n6799) );
  XNOR U3311 ( .A(n7128), .B(n6799), .Z(out[1435]) );
  XNOR U3312 ( .A(in[817]), .B(n8585), .Z(n7132) );
  NAND U3313 ( .A(n6936), .B(n6800), .Z(n6801) );
  XNOR U3314 ( .A(n7132), .B(n6801), .Z(out[1436]) );
  XNOR U3315 ( .A(in[818]), .B(n8589), .Z(n7136) );
  NAND U3316 ( .A(n6938), .B(n6802), .Z(n6803) );
  XNOR U3317 ( .A(n7136), .B(n6803), .Z(out[1437]) );
  XNOR U3318 ( .A(in[819]), .B(n8593), .Z(n7140) );
  NAND U3319 ( .A(n6940), .B(n6804), .Z(n6805) );
  XNOR U3320 ( .A(n7140), .B(n6805), .Z(out[1438]) );
  XNOR U3321 ( .A(in[820]), .B(n8597), .Z(n7144) );
  NAND U3322 ( .A(n6942), .B(n6806), .Z(n6807) );
  XNOR U3323 ( .A(n7144), .B(n6807), .Z(out[1439]) );
  XNOR U3324 ( .A(in[680]), .B(n8735), .Z(n7456) );
  XOR U3325 ( .A(in[614]), .B(n8587), .Z(n8882) );
  XOR U3326 ( .A(in[205]), .B(n8404), .Z(n8880) );
  NAND U3327 ( .A(n8882), .B(n8880), .Z(n6808) );
  XNOR U3328 ( .A(n7456), .B(n6808), .Z(out[143]) );
  XNOR U3329 ( .A(in[821]), .B(n8601), .Z(n7149) );
  NAND U3330 ( .A(n6944), .B(n6809), .Z(n6810) );
  XNOR U3331 ( .A(n7149), .B(n6810), .Z(out[1440]) );
  XNOR U3332 ( .A(in[822]), .B(n8611), .Z(n7153) );
  NAND U3333 ( .A(n6946), .B(n6811), .Z(n6812) );
  XNOR U3334 ( .A(n7153), .B(n6812), .Z(out[1441]) );
  XNOR U3335 ( .A(in[823]), .B(n8615), .Z(n7158) );
  NAND U3336 ( .A(n6948), .B(n6813), .Z(n6814) );
  XNOR U3337 ( .A(n7158), .B(n6814), .Z(out[1442]) );
  XNOR U3338 ( .A(in[824]), .B(n8619), .Z(n7162) );
  NAND U3339 ( .A(n6950), .B(n6815), .Z(n6816) );
  XNOR U3340 ( .A(n7162), .B(n6816), .Z(out[1443]) );
  XNOR U3341 ( .A(in[825]), .B(n8623), .Z(n7166) );
  NAND U3342 ( .A(n6952), .B(n6817), .Z(n6818) );
  XNOR U3343 ( .A(n7166), .B(n6818), .Z(out[1444]) );
  XNOR U3344 ( .A(in[826]), .B(n8345), .Z(n7170) );
  NAND U3345 ( .A(n6954), .B(n6819), .Z(n6820) );
  XNOR U3346 ( .A(n7170), .B(n6820), .Z(out[1445]) );
  XNOR U3347 ( .A(in[827]), .B(n8349), .Z(n7174) );
  NAND U3348 ( .A(n6957), .B(n6821), .Z(n6822) );
  XNOR U3349 ( .A(n7174), .B(n6822), .Z(out[1446]) );
  XNOR U3350 ( .A(in[828]), .B(n8353), .Z(n7178) );
  NAND U3351 ( .A(n6959), .B(n6823), .Z(n6824) );
  XNOR U3352 ( .A(n7178), .B(n6824), .Z(out[1447]) );
  XNOR U3353 ( .A(in[829]), .B(n8357), .Z(n7182) );
  NAND U3354 ( .A(n6961), .B(n6825), .Z(n6826) );
  XNOR U3355 ( .A(n7182), .B(n6826), .Z(out[1448]) );
  XNOR U3356 ( .A(in[830]), .B(n8361), .Z(n7186) );
  NAND U3357 ( .A(n6963), .B(n6827), .Z(n6828) );
  XNOR U3358 ( .A(n7186), .B(n6828), .Z(out[1449]) );
  XNOR U3359 ( .A(in[681]), .B(n8737), .Z(n7459) );
  XOR U3360 ( .A(in[615]), .B(n8591), .Z(n8920) );
  XOR U3361 ( .A(in[206]), .B(n8408), .Z(n8918) );
  NAND U3362 ( .A(n8920), .B(n8918), .Z(n6829) );
  XNOR U3363 ( .A(n7459), .B(n6829), .Z(out[144]) );
  XNOR U3364 ( .A(in[831]), .B(n8365), .Z(n7190) );
  NAND U3365 ( .A(n6965), .B(n6830), .Z(n6831) );
  XNOR U3366 ( .A(n7190), .B(n6831), .Z(out[1450]) );
  XNOR U3367 ( .A(in[768]), .B(n8369), .Z(n7194) );
  NAND U3368 ( .A(n6967), .B(n6832), .Z(n6833) );
  XNOR U3369 ( .A(n7194), .B(n6833), .Z(out[1451]) );
  XNOR U3370 ( .A(in[769]), .B(n8373), .Z(n7199) );
  NAND U3371 ( .A(n6969), .B(n6834), .Z(n6835) );
  XNOR U3372 ( .A(n7199), .B(n6835), .Z(out[1452]) );
  XOR U3373 ( .A(n8377), .B(in[770]), .Z(n7203) );
  NAND U3374 ( .A(n6971), .B(n6836), .Z(n6837) );
  XNOR U3375 ( .A(n7203), .B(n6837), .Z(out[1453]) );
  XOR U3376 ( .A(n8381), .B(in[771]), .Z(n7207) );
  NAND U3377 ( .A(n6973), .B(n6838), .Z(n6839) );
  XNOR U3378 ( .A(n7207), .B(n6839), .Z(out[1454]) );
  XOR U3379 ( .A(n8389), .B(in[772]), .Z(n7211) );
  NAND U3380 ( .A(n6975), .B(n6840), .Z(n6841) );
  XNOR U3381 ( .A(n7211), .B(n6841), .Z(out[1455]) );
  XOR U3382 ( .A(n8393), .B(in[773]), .Z(n7215) );
  NAND U3383 ( .A(n6978), .B(n6842), .Z(n6843) );
  XNOR U3384 ( .A(n7215), .B(n6843), .Z(out[1456]) );
  XOR U3385 ( .A(n8397), .B(in[774]), .Z(n7219) );
  NAND U3386 ( .A(n6980), .B(n6844), .Z(n6845) );
  XNOR U3387 ( .A(n7219), .B(n6845), .Z(out[1457]) );
  XOR U3388 ( .A(n8401), .B(in[775]), .Z(n7223) );
  NAND U3389 ( .A(n6982), .B(n6846), .Z(n6847) );
  XNOR U3390 ( .A(n7223), .B(n6847), .Z(out[1458]) );
  XOR U3391 ( .A(n8405), .B(in[776]), .Z(n7227) );
  NAND U3392 ( .A(n6984), .B(n6848), .Z(n6849) );
  XNOR U3393 ( .A(n7227), .B(n6849), .Z(out[1459]) );
  XNOR U3394 ( .A(in[682]), .B(n8739), .Z(n7462) );
  XOR U3395 ( .A(in[616]), .B(n8595), .Z(n8954) );
  XOR U3396 ( .A(in[207]), .B(n8412), .Z(n8952) );
  NAND U3397 ( .A(n8954), .B(n8952), .Z(n6850) );
  XNOR U3398 ( .A(n7462), .B(n6850), .Z(out[145]) );
  XOR U3399 ( .A(in[777]), .B(n8409), .Z(n7231) );
  NAND U3400 ( .A(n6986), .B(n6851), .Z(n6852) );
  XNOR U3401 ( .A(n7231), .B(n6852), .Z(out[1460]) );
  XOR U3402 ( .A(n8413), .B(in[778]), .Z(n7235) );
  NAND U3403 ( .A(n6988), .B(n6853), .Z(n6854) );
  XNOR U3404 ( .A(n7235), .B(n6854), .Z(out[1461]) );
  XOR U3405 ( .A(n8417), .B(in[779]), .Z(n7240) );
  NAND U3406 ( .A(n6990), .B(n6855), .Z(n6856) );
  XNOR U3407 ( .A(n7240), .B(n6856), .Z(out[1462]) );
  XOR U3408 ( .A(in[780]), .B(n8421), .Z(n7244) );
  NAND U3409 ( .A(n6992), .B(n6857), .Z(n6858) );
  XNOR U3410 ( .A(n7244), .B(n6858), .Z(out[1463]) );
  XOR U3411 ( .A(in[781]), .B(n8425), .Z(n7248) );
  NAND U3412 ( .A(n6994), .B(n6859), .Z(n6860) );
  XNOR U3413 ( .A(n7248), .B(n6860), .Z(out[1464]) );
  XOR U3414 ( .A(in[782]), .B(n8433), .Z(n7252) );
  NAND U3415 ( .A(n6996), .B(n6861), .Z(n6862) );
  XNOR U3416 ( .A(n7252), .B(n6862), .Z(out[1465]) );
  XOR U3417 ( .A(in[783]), .B(n8437), .Z(n7256) );
  NAND U3418 ( .A(n6999), .B(n6863), .Z(n6864) );
  XNOR U3419 ( .A(n7256), .B(n6864), .Z(out[1466]) );
  XOR U3420 ( .A(in[784]), .B(n8441), .Z(n7260) );
  NAND U3421 ( .A(n7001), .B(n6865), .Z(n6866) );
  XNOR U3422 ( .A(n7260), .B(n6866), .Z(out[1467]) );
  XOR U3423 ( .A(in[785]), .B(n8445), .Z(n7264) );
  NAND U3424 ( .A(n7003), .B(n6867), .Z(n6868) );
  XNOR U3425 ( .A(n7264), .B(n6868), .Z(out[1468]) );
  XOR U3426 ( .A(in[786]), .B(n8449), .Z(n7268) );
  NAND U3427 ( .A(n7005), .B(n6869), .Z(n6870) );
  XNOR U3428 ( .A(n7268), .B(n6870), .Z(out[1469]) );
  XNOR U3429 ( .A(in[683]), .B(n8741), .Z(n7465) );
  XOR U3430 ( .A(in[617]), .B(n8599), .Z(n8988) );
  XOR U3431 ( .A(in[208]), .B(n8416), .Z(n8986) );
  NAND U3432 ( .A(n8988), .B(n8986), .Z(n6871) );
  XNOR U3433 ( .A(n7465), .B(n6871), .Z(out[146]) );
  XOR U3434 ( .A(in[787]), .B(n8453), .Z(n7272) );
  NAND U3435 ( .A(n7007), .B(n6872), .Z(n6873) );
  XNOR U3436 ( .A(n7272), .B(n6873), .Z(out[1470]) );
  XOR U3437 ( .A(in[788]), .B(n8457), .Z(n7276) );
  NAND U3438 ( .A(n7009), .B(n6874), .Z(n6875) );
  XNOR U3439 ( .A(n7276), .B(n6875), .Z(out[1471]) );
  OR U3440 ( .A(n7012), .B(n6876), .Z(n6877) );
  XNOR U3441 ( .A(n7011), .B(n6877), .Z(out[1472]) );
  OR U3442 ( .A(n7017), .B(n6878), .Z(n6879) );
  XNOR U3443 ( .A(n7016), .B(n6879), .Z(out[1473]) );
  OR U3444 ( .A(n7022), .B(n6880), .Z(n6881) );
  XNOR U3445 ( .A(n7021), .B(n6881), .Z(out[1474]) );
  OR U3446 ( .A(n7026), .B(n6882), .Z(n6883) );
  XNOR U3447 ( .A(n7025), .B(n6883), .Z(out[1475]) );
  OR U3448 ( .A(n7032), .B(n6884), .Z(n6885) );
  XNOR U3449 ( .A(n7031), .B(n6885), .Z(out[1476]) );
  OR U3450 ( .A(n7036), .B(n6886), .Z(n6887) );
  XNOR U3451 ( .A(n7035), .B(n6887), .Z(out[1477]) );
  OR U3452 ( .A(n7040), .B(n6888), .Z(n6889) );
  XNOR U3453 ( .A(n7039), .B(n6889), .Z(out[1478]) );
  OR U3454 ( .A(n7044), .B(n6890), .Z(n6891) );
  XNOR U3455 ( .A(n7043), .B(n6891), .Z(out[1479]) );
  XNOR U3456 ( .A(in[684]), .B(n8743), .Z(n7468) );
  XOR U3457 ( .A(in[618]), .B(n8609), .Z(n9014) );
  XOR U3458 ( .A(in[209]), .B(n8420), .Z(n9012) );
  NAND U3459 ( .A(n9014), .B(n9012), .Z(n6892) );
  XNOR U3460 ( .A(n7468), .B(n6892), .Z(out[147]) );
  OR U3461 ( .A(n7049), .B(n6893), .Z(n6894) );
  XNOR U3462 ( .A(n7048), .B(n6894), .Z(out[1480]) );
  OR U3463 ( .A(n7053), .B(n6895), .Z(n6896) );
  XNOR U3464 ( .A(n7052), .B(n6896), .Z(out[1481]) );
  OR U3465 ( .A(n7057), .B(n6897), .Z(n6898) );
  XNOR U3466 ( .A(n7056), .B(n6898), .Z(out[1482]) );
  OR U3467 ( .A(n7061), .B(n6899), .Z(n6900) );
  XNOR U3468 ( .A(n7060), .B(n6900), .Z(out[1483]) );
  OR U3469 ( .A(n7065), .B(n6901), .Z(n6902) );
  XNOR U3470 ( .A(n7064), .B(n6902), .Z(out[1484]) );
  OR U3471 ( .A(n7069), .B(n6903), .Z(n6904) );
  XNOR U3472 ( .A(n7068), .B(n6904), .Z(out[1485]) );
  OR U3473 ( .A(n7074), .B(n6905), .Z(n6906) );
  XNOR U3474 ( .A(n7073), .B(n6906), .Z(out[1486]) );
  OR U3475 ( .A(n7078), .B(n6907), .Z(n6908) );
  XNOR U3476 ( .A(n7077), .B(n6908), .Z(out[1487]) );
  OR U3477 ( .A(n7083), .B(n6909), .Z(n6910) );
  XNOR U3478 ( .A(n7082), .B(n6910), .Z(out[1488]) );
  OR U3479 ( .A(n7087), .B(n6911), .Z(n6912) );
  XNOR U3480 ( .A(n7086), .B(n6912), .Z(out[1489]) );
  XNOR U3481 ( .A(in[685]), .B(n8745), .Z(n7471) );
  XOR U3482 ( .A(in[619]), .B(n8613), .Z(n9038) );
  XOR U3483 ( .A(in[210]), .B(n8424), .Z(n9036) );
  NAND U3484 ( .A(n9038), .B(n9036), .Z(n6913) );
  XNOR U3485 ( .A(n7471), .B(n6913), .Z(out[148]) );
  OR U3486 ( .A(n7091), .B(n6914), .Z(n6915) );
  XNOR U3487 ( .A(n7090), .B(n6915), .Z(out[1490]) );
  OR U3488 ( .A(n7095), .B(n6916), .Z(n6917) );
  XNOR U3489 ( .A(n7094), .B(n6917), .Z(out[1491]) );
  OR U3490 ( .A(n7099), .B(n6918), .Z(n6919) );
  XNOR U3491 ( .A(n7098), .B(n6919), .Z(out[1492]) );
  OR U3492 ( .A(n7103), .B(n6920), .Z(n6921) );
  XNOR U3493 ( .A(n7102), .B(n6921), .Z(out[1493]) );
  OR U3494 ( .A(n7107), .B(n6922), .Z(n6923) );
  XNOR U3495 ( .A(n7106), .B(n6923), .Z(out[1494]) );
  OR U3496 ( .A(n7111), .B(n6924), .Z(n6925) );
  XNOR U3497 ( .A(n7110), .B(n6925), .Z(out[1495]) );
  OR U3498 ( .A(n7116), .B(n6926), .Z(n6927) );
  XNOR U3499 ( .A(n7115), .B(n6927), .Z(out[1496]) );
  OR U3500 ( .A(n7120), .B(n6928), .Z(n6929) );
  XNOR U3501 ( .A(n7119), .B(n6929), .Z(out[1497]) );
  OR U3502 ( .A(n7124), .B(n6930), .Z(n6931) );
  XNOR U3503 ( .A(n7123), .B(n6931), .Z(out[1498]) );
  OR U3504 ( .A(n7128), .B(n6932), .Z(n6933) );
  XNOR U3505 ( .A(n7127), .B(n6933), .Z(out[1499]) );
  XNOR U3506 ( .A(in[686]), .B(n8747), .Z(n7473) );
  XOR U3507 ( .A(in[620]), .B(n8617), .Z(n9062) );
  XNOR U3508 ( .A(in[211]), .B(n8432), .Z(n9060) );
  NAND U3509 ( .A(n9062), .B(n9060), .Z(n6934) );
  XNOR U3510 ( .A(n7473), .B(n6934), .Z(out[149]) );
  XNOR U3511 ( .A(in[1424]), .B(n8441), .Z(n8845) );
  XOR U3512 ( .A(in[1047]), .B(n8939), .Z(n7452) );
  NAND U3513 ( .A(n8845), .B(n7452), .Z(n6935) );
  XNOR U3514 ( .A(n8846), .B(n6935), .Z(out[14]) );
  OR U3515 ( .A(n7132), .B(n6936), .Z(n6937) );
  XNOR U3516 ( .A(n7131), .B(n6937), .Z(out[1500]) );
  OR U3517 ( .A(n7136), .B(n6938), .Z(n6939) );
  XNOR U3518 ( .A(n7135), .B(n6939), .Z(out[1501]) );
  OR U3519 ( .A(n7140), .B(n6940), .Z(n6941) );
  XNOR U3520 ( .A(n7139), .B(n6941), .Z(out[1502]) );
  OR U3521 ( .A(n7144), .B(n6942), .Z(n6943) );
  XNOR U3522 ( .A(n7143), .B(n6943), .Z(out[1503]) );
  OR U3523 ( .A(n7149), .B(n6944), .Z(n6945) );
  XNOR U3524 ( .A(n7148), .B(n6945), .Z(out[1504]) );
  OR U3525 ( .A(n7153), .B(n6946), .Z(n6947) );
  XNOR U3526 ( .A(n7152), .B(n6947), .Z(out[1505]) );
  OR U3527 ( .A(n7158), .B(n6948), .Z(n6949) );
  XNOR U3528 ( .A(n7157), .B(n6949), .Z(out[1506]) );
  OR U3529 ( .A(n7162), .B(n6950), .Z(n6951) );
  XNOR U3530 ( .A(n7161), .B(n6951), .Z(out[1507]) );
  OR U3531 ( .A(n7166), .B(n6952), .Z(n6953) );
  XNOR U3532 ( .A(n7165), .B(n6953), .Z(out[1508]) );
  OR U3533 ( .A(n7170), .B(n6954), .Z(n6955) );
  XNOR U3534 ( .A(n7169), .B(n6955), .Z(out[1509]) );
  XNOR U3535 ( .A(in[687]), .B(n8749), .Z(n7476) );
  XOR U3536 ( .A(in[621]), .B(n8621), .Z(n9086) );
  XNOR U3537 ( .A(in[212]), .B(n8436), .Z(n9084) );
  NAND U3538 ( .A(n9086), .B(n9084), .Z(n6956) );
  XNOR U3539 ( .A(n7476), .B(n6956), .Z(out[150]) );
  OR U3540 ( .A(n7174), .B(n6957), .Z(n6958) );
  XNOR U3541 ( .A(n7173), .B(n6958), .Z(out[1510]) );
  OR U3542 ( .A(n7178), .B(n6959), .Z(n6960) );
  XNOR U3543 ( .A(n7177), .B(n6960), .Z(out[1511]) );
  OR U3544 ( .A(n7182), .B(n6961), .Z(n6962) );
  XNOR U3545 ( .A(n7181), .B(n6962), .Z(out[1512]) );
  OR U3546 ( .A(n7186), .B(n6963), .Z(n6964) );
  XNOR U3547 ( .A(n7185), .B(n6964), .Z(out[1513]) );
  OR U3548 ( .A(n7190), .B(n6965), .Z(n6966) );
  XNOR U3549 ( .A(n7189), .B(n6966), .Z(out[1514]) );
  OR U3550 ( .A(n7194), .B(n6967), .Z(n6968) );
  XNOR U3551 ( .A(n7193), .B(n6968), .Z(out[1515]) );
  OR U3552 ( .A(n7199), .B(n6969), .Z(n6970) );
  XNOR U3553 ( .A(n7198), .B(n6970), .Z(out[1516]) );
  OR U3554 ( .A(n7203), .B(n6971), .Z(n6972) );
  XNOR U3555 ( .A(n7202), .B(n6972), .Z(out[1517]) );
  OR U3556 ( .A(n7207), .B(n6973), .Z(n6974) );
  XNOR U3557 ( .A(n7206), .B(n6974), .Z(out[1518]) );
  OR U3558 ( .A(n7211), .B(n6975), .Z(n6976) );
  XNOR U3559 ( .A(n7210), .B(n6976), .Z(out[1519]) );
  XNOR U3560 ( .A(in[688]), .B(n8755), .Z(n7479) );
  XOR U3561 ( .A(in[622]), .B(n8343), .Z(n9110) );
  XNOR U3562 ( .A(in[213]), .B(n8440), .Z(n9108) );
  NAND U3563 ( .A(n9110), .B(n9108), .Z(n6977) );
  XNOR U3564 ( .A(n7479), .B(n6977), .Z(out[151]) );
  OR U3565 ( .A(n7215), .B(n6978), .Z(n6979) );
  XNOR U3566 ( .A(n7214), .B(n6979), .Z(out[1520]) );
  OR U3567 ( .A(n7219), .B(n6980), .Z(n6981) );
  XNOR U3568 ( .A(n7218), .B(n6981), .Z(out[1521]) );
  OR U3569 ( .A(n7223), .B(n6982), .Z(n6983) );
  XNOR U3570 ( .A(n7222), .B(n6983), .Z(out[1522]) );
  OR U3571 ( .A(n7227), .B(n6984), .Z(n6985) );
  XNOR U3572 ( .A(n7226), .B(n6985), .Z(out[1523]) );
  OR U3573 ( .A(n7231), .B(n6986), .Z(n6987) );
  XNOR U3574 ( .A(n7230), .B(n6987), .Z(out[1524]) );
  OR U3575 ( .A(n7235), .B(n6988), .Z(n6989) );
  XNOR U3576 ( .A(n7234), .B(n6989), .Z(out[1525]) );
  OR U3577 ( .A(n7240), .B(n6990), .Z(n6991) );
  XNOR U3578 ( .A(n7239), .B(n6991), .Z(out[1526]) );
  OR U3579 ( .A(n7244), .B(n6992), .Z(n6993) );
  XNOR U3580 ( .A(n7243), .B(n6993), .Z(out[1527]) );
  OR U3581 ( .A(n7248), .B(n6994), .Z(n6995) );
  XNOR U3582 ( .A(n7247), .B(n6995), .Z(out[1528]) );
  OR U3583 ( .A(n7252), .B(n6996), .Z(n6997) );
  XNOR U3584 ( .A(n7251), .B(n6997), .Z(out[1529]) );
  XNOR U3585 ( .A(in[689]), .B(n8757), .Z(n7483) );
  XOR U3586 ( .A(in[623]), .B(n8347), .Z(n9134) );
  XNOR U3587 ( .A(in[214]), .B(n8444), .Z(n9132) );
  NAND U3588 ( .A(n9134), .B(n9132), .Z(n6998) );
  XNOR U3589 ( .A(n7483), .B(n6998), .Z(out[152]) );
  OR U3590 ( .A(n7256), .B(n6999), .Z(n7000) );
  XNOR U3591 ( .A(n7255), .B(n7000), .Z(out[1530]) );
  OR U3592 ( .A(n7260), .B(n7001), .Z(n7002) );
  XNOR U3593 ( .A(n7259), .B(n7002), .Z(out[1531]) );
  OR U3594 ( .A(n7264), .B(n7003), .Z(n7004) );
  XNOR U3595 ( .A(n7263), .B(n7004), .Z(out[1532]) );
  OR U3596 ( .A(n7268), .B(n7005), .Z(n7006) );
  XNOR U3597 ( .A(n7267), .B(n7006), .Z(out[1533]) );
  OR U3598 ( .A(n7272), .B(n7007), .Z(n7008) );
  XNOR U3599 ( .A(n7271), .B(n7008), .Z(out[1534]) );
  OR U3600 ( .A(n7276), .B(n7009), .Z(n7010) );
  XNOR U3601 ( .A(n7275), .B(n7010), .Z(out[1535]) );
  ANDN U3602 ( .B(n7012), .A(n7011), .Z(n7015) );
  XOR U3603 ( .A(n7013), .B(round_const[0]), .Z(n7014) );
  XNOR U3604 ( .A(n7015), .B(n7014), .Z(out[1536]) );
  ANDN U3605 ( .B(n7017), .A(n7016), .Z(n7020) );
  XOR U3606 ( .A(n7018), .B(round_const[1]), .Z(n7019) );
  XNOR U3607 ( .A(n7020), .B(n7019), .Z(out[1537]) );
  ANDN U3608 ( .B(n7022), .A(n7021), .Z(n7023) );
  XNOR U3609 ( .A(n7024), .B(n7023), .Z(out[1538]) );
  ANDN U3610 ( .B(n7026), .A(n7025), .Z(n7029) );
  XOR U3611 ( .A(n7027), .B(round_const_3), .Z(n7028) );
  XNOR U3612 ( .A(n7029), .B(n7028), .Z(out[1539]) );
  XNOR U3613 ( .A(in[690]), .B(n8759), .Z(n7486) );
  XOR U3614 ( .A(in[624]), .B(n8351), .Z(n9166) );
  XNOR U3615 ( .A(in[215]), .B(n8448), .Z(n9164) );
  NAND U3616 ( .A(n9166), .B(n9164), .Z(n7030) );
  XNOR U3617 ( .A(n7486), .B(n7030), .Z(out[153]) );
  ANDN U3618 ( .B(n7032), .A(n7031), .Z(n7033) );
  XNOR U3619 ( .A(n7034), .B(n7033), .Z(out[1540]) );
  ANDN U3620 ( .B(n7036), .A(n7035), .Z(n7037) );
  XNOR U3621 ( .A(n7038), .B(n7037), .Z(out[1541]) );
  ANDN U3622 ( .B(n7040), .A(n7039), .Z(n7041) );
  XNOR U3623 ( .A(n7042), .B(n7041), .Z(out[1542]) );
  ANDN U3624 ( .B(n7044), .A(n7043), .Z(n7047) );
  XOR U3625 ( .A(n7045), .B(round_const_7), .Z(n7046) );
  XNOR U3626 ( .A(n7047), .B(n7046), .Z(out[1543]) );
  ANDN U3627 ( .B(n7049), .A(n7048), .Z(n7050) );
  XNOR U3628 ( .A(n7051), .B(n7050), .Z(out[1544]) );
  ANDN U3629 ( .B(n7053), .A(n7052), .Z(n7054) );
  XNOR U3630 ( .A(n7055), .B(n7054), .Z(out[1545]) );
  ANDN U3631 ( .B(n7057), .A(n7056), .Z(n7058) );
  XNOR U3632 ( .A(n7059), .B(n7058), .Z(out[1546]) );
  ANDN U3633 ( .B(n7061), .A(n7060), .Z(n7062) );
  XNOR U3634 ( .A(n7063), .B(n7062), .Z(out[1547]) );
  ANDN U3635 ( .B(n7065), .A(n7064), .Z(n7066) );
  XNOR U3636 ( .A(n7067), .B(n7066), .Z(out[1548]) );
  ANDN U3637 ( .B(n7069), .A(n7068), .Z(n7070) );
  XNOR U3638 ( .A(n7071), .B(n7070), .Z(out[1549]) );
  XNOR U3639 ( .A(in[691]), .B(n8761), .Z(n7489) );
  XOR U3640 ( .A(in[625]), .B(n8355), .Z(n9214) );
  XNOR U3641 ( .A(in[216]), .B(n8452), .Z(n9212) );
  NAND U3642 ( .A(n9214), .B(n9212), .Z(n7072) );
  XNOR U3643 ( .A(n7489), .B(n7072), .Z(out[154]) );
  ANDN U3644 ( .B(n7074), .A(n7073), .Z(n7075) );
  XNOR U3645 ( .A(n7076), .B(n7075), .Z(out[1550]) );
  ANDN U3646 ( .B(n7078), .A(n7077), .Z(n7081) );
  XOR U3647 ( .A(n7079), .B(round_const_15), .Z(n7080) );
  XNOR U3648 ( .A(n7081), .B(n7080), .Z(out[1551]) );
  ANDN U3649 ( .B(n7083), .A(n7082), .Z(n7084) );
  XNOR U3650 ( .A(n7085), .B(n7084), .Z(out[1552]) );
  ANDN U3651 ( .B(n7087), .A(n7086), .Z(n7088) );
  XNOR U3652 ( .A(n7089), .B(n7088), .Z(out[1553]) );
  ANDN U3653 ( .B(n7091), .A(n7090), .Z(n7092) );
  XNOR U3654 ( .A(n7093), .B(n7092), .Z(out[1554]) );
  ANDN U3655 ( .B(n7095), .A(n7094), .Z(n7096) );
  XNOR U3656 ( .A(n7097), .B(n7096), .Z(out[1555]) );
  ANDN U3657 ( .B(n7099), .A(n7098), .Z(n7100) );
  XNOR U3658 ( .A(n7101), .B(n7100), .Z(out[1556]) );
  ANDN U3659 ( .B(n7103), .A(n7102), .Z(n7104) );
  XNOR U3660 ( .A(n7105), .B(n7104), .Z(out[1557]) );
  ANDN U3661 ( .B(n7107), .A(n7106), .Z(n7108) );
  XNOR U3662 ( .A(n7109), .B(n7108), .Z(out[1558]) );
  ANDN U3663 ( .B(n7111), .A(n7110), .Z(n7112) );
  XNOR U3664 ( .A(n7113), .B(n7112), .Z(out[1559]) );
  XNOR U3665 ( .A(in[692]), .B(n8763), .Z(n7492) );
  XOR U3666 ( .A(in[626]), .B(n8359), .Z(n9258) );
  XNOR U3667 ( .A(in[217]), .B(n8456), .Z(n9256) );
  NAND U3668 ( .A(n9258), .B(n9256), .Z(n7114) );
  XNOR U3669 ( .A(n7492), .B(n7114), .Z(out[155]) );
  ANDN U3670 ( .B(n7116), .A(n7115), .Z(n7117) );
  XNOR U3671 ( .A(n7118), .B(n7117), .Z(out[1560]) );
  ANDN U3672 ( .B(n7120), .A(n7119), .Z(n7121) );
  XNOR U3673 ( .A(n7122), .B(n7121), .Z(out[1561]) );
  ANDN U3674 ( .B(n7124), .A(n7123), .Z(n7125) );
  XNOR U3675 ( .A(n7126), .B(n7125), .Z(out[1562]) );
  ANDN U3676 ( .B(n7128), .A(n7127), .Z(n7129) );
  XNOR U3677 ( .A(n7130), .B(n7129), .Z(out[1563]) );
  ANDN U3678 ( .B(n7132), .A(n7131), .Z(n7133) );
  XNOR U3679 ( .A(n7134), .B(n7133), .Z(out[1564]) );
  ANDN U3680 ( .B(n7136), .A(n7135), .Z(n7137) );
  XNOR U3681 ( .A(n7138), .B(n7137), .Z(out[1565]) );
  ANDN U3682 ( .B(n7140), .A(n7139), .Z(n7141) );
  XNOR U3683 ( .A(n7142), .B(n7141), .Z(out[1566]) );
  ANDN U3684 ( .B(n7144), .A(n7143), .Z(n7147) );
  XOR U3685 ( .A(n7145), .B(round_const_31), .Z(n7146) );
  XNOR U3686 ( .A(n7147), .B(n7146), .Z(out[1567]) );
  ANDN U3687 ( .B(n7149), .A(n7148), .Z(n7150) );
  XNOR U3688 ( .A(n7151), .B(n7150), .Z(out[1568]) );
  ANDN U3689 ( .B(n7153), .A(n7152), .Z(n7154) );
  XNOR U3690 ( .A(n7155), .B(n7154), .Z(out[1569]) );
  XNOR U3691 ( .A(in[693]), .B(n8765), .Z(n7495) );
  XOR U3692 ( .A(in[627]), .B(n8363), .Z(n9302) );
  XNOR U3693 ( .A(in[218]), .B(n8460), .Z(n9299) );
  NAND U3694 ( .A(n9302), .B(n9299), .Z(n7156) );
  XNOR U3695 ( .A(n7495), .B(n7156), .Z(out[156]) );
  ANDN U3696 ( .B(n7158), .A(n7157), .Z(n7159) );
  XNOR U3697 ( .A(n7160), .B(n7159), .Z(out[1570]) );
  ANDN U3698 ( .B(n7162), .A(n7161), .Z(n7163) );
  XNOR U3699 ( .A(n7164), .B(n7163), .Z(out[1571]) );
  ANDN U3700 ( .B(n7166), .A(n7165), .Z(n7167) );
  XNOR U3701 ( .A(n7168), .B(n7167), .Z(out[1572]) );
  ANDN U3702 ( .B(n7170), .A(n7169), .Z(n7171) );
  XNOR U3703 ( .A(n7172), .B(n7171), .Z(out[1573]) );
  ANDN U3704 ( .B(n7174), .A(n7173), .Z(n7175) );
  XNOR U3705 ( .A(n7176), .B(n7175), .Z(out[1574]) );
  ANDN U3706 ( .B(n7178), .A(n7177), .Z(n7179) );
  XNOR U3707 ( .A(n7180), .B(n7179), .Z(out[1575]) );
  ANDN U3708 ( .B(n7182), .A(n7181), .Z(n7183) );
  XNOR U3709 ( .A(n7184), .B(n7183), .Z(out[1576]) );
  ANDN U3710 ( .B(n7186), .A(n7185), .Z(n7187) );
  XNOR U3711 ( .A(n7188), .B(n7187), .Z(out[1577]) );
  ANDN U3712 ( .B(n7190), .A(n7189), .Z(n7191) );
  XNOR U3713 ( .A(n7192), .B(n7191), .Z(out[1578]) );
  ANDN U3714 ( .B(n7194), .A(n7193), .Z(n7195) );
  XNOR U3715 ( .A(n7196), .B(n7195), .Z(out[1579]) );
  XNOR U3716 ( .A(in[694]), .B(n8767), .Z(n7497) );
  XOR U3717 ( .A(in[628]), .B(n8367), .Z(n9346) );
  XNOR U3718 ( .A(in[219]), .B(n8464), .Z(n9343) );
  NAND U3719 ( .A(n9346), .B(n9343), .Z(n7197) );
  XNOR U3720 ( .A(n7497), .B(n7197), .Z(out[157]) );
  ANDN U3721 ( .B(n7199), .A(n7198), .Z(n7200) );
  XNOR U3722 ( .A(n7201), .B(n7200), .Z(out[1580]) );
  ANDN U3723 ( .B(n7203), .A(n7202), .Z(n7204) );
  XNOR U3724 ( .A(n7205), .B(n7204), .Z(out[1581]) );
  ANDN U3725 ( .B(n7207), .A(n7206), .Z(n7208) );
  XNOR U3726 ( .A(n7209), .B(n7208), .Z(out[1582]) );
  ANDN U3727 ( .B(n7211), .A(n7210), .Z(n7212) );
  XNOR U3728 ( .A(n7213), .B(n7212), .Z(out[1583]) );
  ANDN U3729 ( .B(n7215), .A(n7214), .Z(n7216) );
  XNOR U3730 ( .A(n7217), .B(n7216), .Z(out[1584]) );
  ANDN U3731 ( .B(n7219), .A(n7218), .Z(n7220) );
  XNOR U3732 ( .A(n7221), .B(n7220), .Z(out[1585]) );
  ANDN U3733 ( .B(n7223), .A(n7222), .Z(n7224) );
  XNOR U3734 ( .A(n7225), .B(n7224), .Z(out[1586]) );
  ANDN U3735 ( .B(n7227), .A(n7226), .Z(n7228) );
  XNOR U3736 ( .A(n7229), .B(n7228), .Z(out[1587]) );
  ANDN U3737 ( .B(n7231), .A(n7230), .Z(n7232) );
  XNOR U3738 ( .A(n7233), .B(n7232), .Z(out[1588]) );
  ANDN U3739 ( .B(n7235), .A(n7234), .Z(n7236) );
  XNOR U3740 ( .A(n7237), .B(n7236), .Z(out[1589]) );
  XNOR U3741 ( .A(in[695]), .B(n8769), .Z(n7499) );
  XOR U3742 ( .A(in[629]), .B(n8371), .Z(n9390) );
  XNOR U3743 ( .A(in[220]), .B(n8468), .Z(n9387) );
  NAND U3744 ( .A(n9390), .B(n9387), .Z(n7238) );
  XNOR U3745 ( .A(n7499), .B(n7238), .Z(out[158]) );
  ANDN U3746 ( .B(n7240), .A(n7239), .Z(n7241) );
  XNOR U3747 ( .A(n7242), .B(n7241), .Z(out[1590]) );
  ANDN U3748 ( .B(n7244), .A(n7243), .Z(n7245) );
  XNOR U3749 ( .A(n7246), .B(n7245), .Z(out[1591]) );
  ANDN U3750 ( .B(n7248), .A(n7247), .Z(n7249) );
  XNOR U3751 ( .A(n7250), .B(n7249), .Z(out[1592]) );
  ANDN U3752 ( .B(n7252), .A(n7251), .Z(n7253) );
  XNOR U3753 ( .A(n7254), .B(n7253), .Z(out[1593]) );
  ANDN U3754 ( .B(n7256), .A(n7255), .Z(n7257) );
  XNOR U3755 ( .A(n7258), .B(n7257), .Z(out[1594]) );
  ANDN U3756 ( .B(n7260), .A(n7259), .Z(n7261) );
  XNOR U3757 ( .A(n7262), .B(n7261), .Z(out[1595]) );
  ANDN U3758 ( .B(n7264), .A(n7263), .Z(n7265) );
  XNOR U3759 ( .A(n7266), .B(n7265), .Z(out[1596]) );
  ANDN U3760 ( .B(n7268), .A(n7267), .Z(n7269) );
  XNOR U3761 ( .A(n7270), .B(n7269), .Z(out[1597]) );
  ANDN U3762 ( .B(n7272), .A(n7271), .Z(n7273) );
  XNOR U3763 ( .A(n7274), .B(n7273), .Z(out[1598]) );
  ANDN U3764 ( .B(n7276), .A(n7275), .Z(n7279) );
  XOR U3765 ( .A(n7277), .B(round_const_63), .Z(n7278) );
  XNOR U3766 ( .A(n7279), .B(n7278), .Z(out[1599]) );
  XNOR U3767 ( .A(in[696]), .B(n8625), .Z(n7501) );
  XOR U3768 ( .A(in[630]), .B(n8375), .Z(n9434) );
  XNOR U3769 ( .A(in[221]), .B(n8476), .Z(n9431) );
  NAND U3770 ( .A(n9434), .B(n9431), .Z(n7280) );
  XNOR U3771 ( .A(n7501), .B(n7280), .Z(out[159]) );
  XNOR U3772 ( .A(in[1425]), .B(n8445), .Z(n8879) );
  XOR U3773 ( .A(in[1048]), .B(n8942), .Z(n7455) );
  NAND U3774 ( .A(n8879), .B(n7455), .Z(n7281) );
  XNOR U3775 ( .A(n8880), .B(n7281), .Z(out[15]) );
  XNOR U3776 ( .A(in[697]), .B(n8627), .Z(n7503) );
  XOR U3777 ( .A(in[631]), .B(n8379), .Z(n9478) );
  XNOR U3778 ( .A(in[222]), .B(n8480), .Z(n9475) );
  NAND U3779 ( .A(n9478), .B(n9475), .Z(n7282) );
  XNOR U3780 ( .A(n7503), .B(n7282), .Z(out[160]) );
  XNOR U3781 ( .A(in[698]), .B(n8629), .Z(n7505) );
  XOR U3782 ( .A(in[632]), .B(n8387), .Z(n9522) );
  XNOR U3783 ( .A(in[223]), .B(n8484), .Z(n9519) );
  NAND U3784 ( .A(n9522), .B(n9519), .Z(n7283) );
  XNOR U3785 ( .A(n7505), .B(n7283), .Z(out[161]) );
  XNOR U3786 ( .A(in[699]), .B(n8631), .Z(n7509) );
  XOR U3787 ( .A(in[633]), .B(n8391), .Z(n9566) );
  XNOR U3788 ( .A(in[224]), .B(n8488), .Z(n9563) );
  NAND U3789 ( .A(n9566), .B(n9563), .Z(n7284) );
  XNOR U3790 ( .A(n7509), .B(n7284), .Z(out[162]) );
  XNOR U3791 ( .A(in[700]), .B(n8633), .Z(n7511) );
  XOR U3792 ( .A(in[634]), .B(n8395), .Z(n9610) );
  XNOR U3793 ( .A(in[225]), .B(n8492), .Z(n9607) );
  NAND U3794 ( .A(n9610), .B(n9607), .Z(n7285) );
  XNOR U3795 ( .A(n7511), .B(n7285), .Z(out[163]) );
  XOR U3796 ( .A(in[701]), .B(n8635), .Z(n7513) );
  NOR U3797 ( .A(n7357), .B(n7638), .Z(n7286) );
  XNOR U3798 ( .A(n7513), .B(n7286), .Z(out[164]) );
  XOR U3799 ( .A(in[702]), .B(n8641), .Z(n7515) );
  NOR U3800 ( .A(n7359), .B(n7652), .Z(n7287) );
  XNOR U3801 ( .A(n7515), .B(n7287), .Z(out[165]) );
  XOR U3802 ( .A(in[703]), .B(n8643), .Z(n7517) );
  NOR U3803 ( .A(n7362), .B(n7666), .Z(n7288) );
  XNOR U3804 ( .A(n7517), .B(n7288), .Z(out[166]) );
  XOR U3805 ( .A(in[640]), .B(n8645), .Z(n7519) );
  NOR U3806 ( .A(n7364), .B(n7680), .Z(n7289) );
  XNOR U3807 ( .A(n7519), .B(n7289), .Z(out[167]) );
  XOR U3808 ( .A(in[641]), .B(n8647), .Z(n7521) );
  NOR U3809 ( .A(n7366), .B(n7696), .Z(n7290) );
  XNOR U3810 ( .A(n7521), .B(n7290), .Z(out[168]) );
  XOR U3811 ( .A(in[642]), .B(n8649), .Z(n7523) );
  NOR U3812 ( .A(n7368), .B(n7710), .Z(n7291) );
  XNOR U3813 ( .A(n7523), .B(n7291), .Z(out[169]) );
  XNOR U3814 ( .A(in[1426]), .B(n8449), .Z(n8917) );
  XOR U3815 ( .A(in[1049]), .B(n8945), .Z(n7458) );
  NAND U3816 ( .A(n8917), .B(n7458), .Z(n7292) );
  XNOR U3817 ( .A(n8918), .B(n7292), .Z(out[16]) );
  XOR U3818 ( .A(in[643]), .B(n8651), .Z(n7525) );
  NOR U3819 ( .A(n7370), .B(n7724), .Z(n7293) );
  XNOR U3820 ( .A(n7525), .B(n7293), .Z(out[170]) );
  XOR U3821 ( .A(in[644]), .B(n8653), .Z(n7527) );
  NOR U3822 ( .A(n7372), .B(n7738), .Z(n7294) );
  XNOR U3823 ( .A(n7527), .B(n7294), .Z(out[171]) );
  XOR U3824 ( .A(in[645]), .B(n8655), .Z(n7533) );
  NOR U3825 ( .A(n7374), .B(n7754), .Z(n7295) );
  XNOR U3826 ( .A(n7533), .B(n7295), .Z(out[172]) );
  XOR U3827 ( .A(in[646]), .B(n8657), .Z(n7535) );
  NOR U3828 ( .A(n7376), .B(n7778), .Z(n7296) );
  XNOR U3829 ( .A(n7535), .B(n7296), .Z(out[173]) );
  XOR U3830 ( .A(in[647]), .B(n8659), .Z(n7537) );
  NOR U3831 ( .A(n7378), .B(n7802), .Z(n7297) );
  XNOR U3832 ( .A(n7537), .B(n7297), .Z(out[174]) );
  XOR U3833 ( .A(in[648]), .B(n8663), .Z(n7539) );
  NOR U3834 ( .A(n7380), .B(n7826), .Z(n7298) );
  XNOR U3835 ( .A(n7539), .B(n7298), .Z(out[175]) );
  XOR U3836 ( .A(in[649]), .B(n8665), .Z(n7541) );
  NOR U3837 ( .A(n7383), .B(n7850), .Z(n7299) );
  XNOR U3838 ( .A(n7541), .B(n7299), .Z(out[176]) );
  XOR U3839 ( .A(in[650]), .B(n8667), .Z(n7543) );
  NOR U3840 ( .A(n7385), .B(n7874), .Z(n7300) );
  XNOR U3841 ( .A(n7543), .B(n7300), .Z(out[177]) );
  XOR U3842 ( .A(in[651]), .B(n8669), .Z(n7545) );
  NOR U3843 ( .A(n7387), .B(n7900), .Z(n7301) );
  XNOR U3844 ( .A(n7545), .B(n7301), .Z(out[178]) );
  XOR U3845 ( .A(in[652]), .B(n8671), .Z(n7547) );
  NOR U3846 ( .A(n7389), .B(n7924), .Z(n7302) );
  XNOR U3847 ( .A(n7547), .B(n7302), .Z(out[179]) );
  XNOR U3848 ( .A(in[1427]), .B(n8453), .Z(n8951) );
  XOR U3849 ( .A(in[1050]), .B(n8948), .Z(n7461) );
  NAND U3850 ( .A(n8951), .B(n7461), .Z(n7303) );
  XNOR U3851 ( .A(n8952), .B(n7303), .Z(out[17]) );
  XOR U3852 ( .A(in[653]), .B(n8673), .Z(n7549) );
  NOR U3853 ( .A(n7391), .B(n7948), .Z(n7304) );
  XNOR U3854 ( .A(n7549), .B(n7304), .Z(out[180]) );
  XOR U3855 ( .A(in[654]), .B(n8675), .Z(n7551) );
  NOR U3856 ( .A(n7393), .B(n7972), .Z(n7305) );
  XNOR U3857 ( .A(n7551), .B(n7305), .Z(out[181]) );
  XOR U3858 ( .A(in[655]), .B(n8677), .Z(n7555) );
  NOR U3859 ( .A(n7395), .B(n7996), .Z(n7306) );
  XNOR U3860 ( .A(n7555), .B(n7306), .Z(out[182]) );
  XOR U3861 ( .A(in[656]), .B(n8679), .Z(n7557) );
  NOR U3862 ( .A(n7397), .B(n8020), .Z(n7307) );
  XNOR U3863 ( .A(n7557), .B(n7307), .Z(out[183]) );
  XOR U3864 ( .A(in[657]), .B(n8681), .Z(n7559) );
  NOR U3865 ( .A(n7399), .B(n8044), .Z(n7308) );
  XNOR U3866 ( .A(n7559), .B(n7308), .Z(out[184]) );
  XOR U3867 ( .A(in[658]), .B(n8685), .Z(n7561) );
  NOR U3868 ( .A(n7401), .B(n8076), .Z(n7309) );
  XNOR U3869 ( .A(n7561), .B(n7309), .Z(out[185]) );
  XOR U3870 ( .A(in[659]), .B(n8687), .Z(n7563) );
  NOR U3871 ( .A(n7404), .B(n8120), .Z(n7310) );
  XNOR U3872 ( .A(n7563), .B(n7310), .Z(out[186]) );
  XOR U3873 ( .A(in[660]), .B(n8689), .Z(n7565) );
  NOR U3874 ( .A(n7406), .B(n8164), .Z(n7311) );
  XNOR U3875 ( .A(n7565), .B(n7311), .Z(out[187]) );
  XOR U3876 ( .A(in[661]), .B(n8691), .Z(n7567) );
  NOR U3877 ( .A(n7408), .B(n8210), .Z(n7312) );
  XNOR U3878 ( .A(n7567), .B(n7312), .Z(out[188]) );
  XOR U3879 ( .A(in[662]), .B(n8693), .Z(n7569) );
  NOR U3880 ( .A(n7410), .B(n8254), .Z(n7313) );
  XNOR U3881 ( .A(n7569), .B(n7313), .Z(out[189]) );
  XNOR U3882 ( .A(in[1428]), .B(n8457), .Z(n8985) );
  XOR U3883 ( .A(in[1051]), .B(n8955), .Z(n7464) );
  NAND U3884 ( .A(n8985), .B(n7464), .Z(n7314) );
  XNOR U3885 ( .A(n8986), .B(n7314), .Z(out[18]) );
  XOR U3886 ( .A(in[663]), .B(n8695), .Z(n7571) );
  NOR U3887 ( .A(n7412), .B(n8298), .Z(n7315) );
  XNOR U3888 ( .A(n7571), .B(n7315), .Z(out[190]) );
  XOR U3889 ( .A(in[664]), .B(n8697), .Z(n7573) );
  NOR U3890 ( .A(n7414), .B(n8342), .Z(n7316) );
  XNOR U3891 ( .A(n7573), .B(n7316), .Z(out[191]) );
  OR U3892 ( .A(n7417), .B(n8386), .Z(n7317) );
  XNOR U3893 ( .A(n7416), .B(n7317), .Z(out[192]) );
  XOR U3894 ( .A(in[1034]), .B(n8896), .Z(n7420) );
  NOR U3895 ( .A(n7419), .B(n8430), .Z(n7318) );
  XNOR U3896 ( .A(n7420), .B(n7318), .Z(out[193]) );
  XOR U3897 ( .A(in[1035]), .B(n8899), .Z(n7531) );
  NOR U3898 ( .A(n7422), .B(n8474), .Z(n7319) );
  XNOR U3899 ( .A(n7531), .B(n7319), .Z(out[194]) );
  XNOR U3900 ( .A(n8902), .B(in[1036]), .Z(n7681) );
  NOR U3901 ( .A(n7424), .B(n8518), .Z(n7320) );
  XNOR U3902 ( .A(n7681), .B(n7320), .Z(out[195]) );
  XNOR U3903 ( .A(n8905), .B(in[1037]), .Z(n7875) );
  NOR U3904 ( .A(n7427), .B(n8562), .Z(n7321) );
  XNOR U3905 ( .A(n7875), .B(n7321), .Z(out[196]) );
  XNOR U3906 ( .A(n8908), .B(in[1038]), .Z(n8165) );
  NOR U3907 ( .A(n7429), .B(n8606), .Z(n7322) );
  XNOR U3908 ( .A(n8165), .B(n7322), .Z(out[197]) );
  XNOR U3909 ( .A(n8911), .B(in[1039]), .Z(n8607) );
  NOR U3910 ( .A(n7431), .B(n8640), .Z(n7323) );
  XNOR U3911 ( .A(n8607), .B(n7323), .Z(out[198]) );
  XNOR U3912 ( .A(n8914), .B(in[1040]), .Z(n8883) );
  NOR U3913 ( .A(n7433), .B(n8662), .Z(n7324) );
  XNOR U3914 ( .A(n8883), .B(n7324), .Z(out[199]) );
  XNOR U3915 ( .A(in[1429]), .B(n8461), .Z(n9011) );
  XOR U3916 ( .A(in[1052]), .B(n8958), .Z(n7467) );
  NAND U3917 ( .A(n9011), .B(n7467), .Z(n7325) );
  XNOR U3918 ( .A(n9012), .B(n7325), .Z(out[19]) );
  XNOR U3919 ( .A(n8381), .B(in[1411]), .Z(n8427) );
  NANDN U3920 ( .A(n7420), .B(n8427), .Z(n7326) );
  XNOR U3921 ( .A(n8428), .B(n7326), .Z(out[1]) );
  XNOR U3922 ( .A(n8921), .B(in[1041]), .Z(n9167) );
  NOR U3923 ( .A(n7435), .B(n8684), .Z(n7327) );
  XNOR U3924 ( .A(n9167), .B(n7327), .Z(out[200]) );
  XNOR U3925 ( .A(n8924), .B(in[1042]), .Z(n9611) );
  NOR U3926 ( .A(n7437), .B(n8706), .Z(n7328) );
  XNOR U3927 ( .A(n9611), .B(n7328), .Z(out[201]) );
  OR U3928 ( .A(n7440), .B(n8730), .Z(n7329) );
  XNOR U3929 ( .A(n7439), .B(n7329), .Z(out[202]) );
  OR U3930 ( .A(n7443), .B(n8754), .Z(n7330) );
  XNOR U3931 ( .A(n7442), .B(n7330), .Z(out[203]) );
  OR U3932 ( .A(n7446), .B(n8780), .Z(n7331) );
  XNOR U3933 ( .A(n7445), .B(n7331), .Z(out[204]) );
  OR U3934 ( .A(n7449), .B(n8814), .Z(n7332) );
  XNOR U3935 ( .A(n7448), .B(n7332), .Z(out[205]) );
  OR U3936 ( .A(n7453), .B(n8848), .Z(n7333) );
  XNOR U3937 ( .A(n7452), .B(n7333), .Z(out[206]) );
  OR U3938 ( .A(n7456), .B(n8882), .Z(n7334) );
  XNOR U3939 ( .A(n7455), .B(n7334), .Z(out[207]) );
  OR U3940 ( .A(n7459), .B(n8920), .Z(n7335) );
  XNOR U3941 ( .A(n7458), .B(n7335), .Z(out[208]) );
  OR U3942 ( .A(n7462), .B(n8954), .Z(n7336) );
  XNOR U3943 ( .A(n7461), .B(n7336), .Z(out[209]) );
  XNOR U3944 ( .A(in[1430]), .B(n8465), .Z(n9035) );
  XOR U3945 ( .A(in[1053]), .B(n8961), .Z(n7470) );
  NAND U3946 ( .A(n9035), .B(n7470), .Z(n7337) );
  XNOR U3947 ( .A(n9036), .B(n7337), .Z(out[20]) );
  OR U3948 ( .A(n7465), .B(n8988), .Z(n7338) );
  XNOR U3949 ( .A(n7464), .B(n7338), .Z(out[210]) );
  OR U3950 ( .A(n7468), .B(n9014), .Z(n7339) );
  XNOR U3951 ( .A(n7467), .B(n7339), .Z(out[211]) );
  OR U3952 ( .A(n7471), .B(n9038), .Z(n7340) );
  XNOR U3953 ( .A(n7470), .B(n7340), .Z(out[212]) );
  XNOR U3954 ( .A(in[1054]), .B(n8964), .Z(n7474) );
  NOR U3955 ( .A(n7473), .B(n9062), .Z(n7341) );
  XNOR U3956 ( .A(n7474), .B(n7341), .Z(out[213]) );
  XNOR U3957 ( .A(in[1055]), .B(n8967), .Z(n7477) );
  NOR U3958 ( .A(n7476), .B(n9086), .Z(n7342) );
  XNOR U3959 ( .A(n7477), .B(n7342), .Z(out[214]) );
  XNOR U3960 ( .A(in[1056]), .B(n8970), .Z(n7480) );
  NOR U3961 ( .A(n7479), .B(n9110), .Z(n7343) );
  XNOR U3962 ( .A(n7480), .B(n7343), .Z(out[215]) );
  XNOR U3963 ( .A(in[1057]), .B(n8973), .Z(n7484) );
  NOR U3964 ( .A(n7483), .B(n9134), .Z(n7344) );
  XNOR U3965 ( .A(n7484), .B(n7344), .Z(out[216]) );
  XNOR U3966 ( .A(in[1058]), .B(n8976), .Z(n7487) );
  NOR U3967 ( .A(n7486), .B(n9166), .Z(n7345) );
  XNOR U3968 ( .A(n7487), .B(n7345), .Z(out[217]) );
  XNOR U3969 ( .A(in[1059]), .B(n8979), .Z(n7490) );
  NOR U3970 ( .A(n7489), .B(n9214), .Z(n7346) );
  XNOR U3971 ( .A(n7490), .B(n7346), .Z(out[218]) );
  XOR U3972 ( .A(in[1060]), .B(n8982), .Z(n7493) );
  NOR U3973 ( .A(n7492), .B(n9258), .Z(n7347) );
  XNOR U3974 ( .A(n7493), .B(n7347), .Z(out[219]) );
  XNOR U3975 ( .A(in[1431]), .B(n8469), .Z(n9059) );
  NANDN U3976 ( .A(n7474), .B(n9059), .Z(n7348) );
  XNOR U3977 ( .A(n9060), .B(n7348), .Z(out[21]) );
  XOR U3978 ( .A(in[1061]), .B(n8989), .Z(n7507) );
  NOR U3979 ( .A(n7495), .B(n9302), .Z(n7349) );
  XNOR U3980 ( .A(n7507), .B(n7349), .Z(out[220]) );
  XOR U3981 ( .A(in[1062]), .B(n8992), .Z(n7529) );
  NOR U3982 ( .A(n7497), .B(n9346), .Z(n7350) );
  XNOR U3983 ( .A(n7529), .B(n7350), .Z(out[221]) );
  XOR U3984 ( .A(in[1063]), .B(n8771), .Z(n7553) );
  NOR U3985 ( .A(n7499), .B(n9390), .Z(n7351) );
  XNOR U3986 ( .A(n7553), .B(n7351), .Z(out[222]) );
  XOR U3987 ( .A(in[1064]), .B(n8774), .Z(n7575) );
  NOR U3988 ( .A(n7501), .B(n9434), .Z(n7352) );
  XNOR U3989 ( .A(n7575), .B(n7352), .Z(out[223]) );
  XOR U3990 ( .A(in[1065]), .B(n8781), .Z(n7587) );
  NOR U3991 ( .A(n7503), .B(n9478), .Z(n7353) );
  XNOR U3992 ( .A(n7587), .B(n7353), .Z(out[224]) );
  XOR U3993 ( .A(in[1066]), .B(n8784), .Z(n7599) );
  NOR U3994 ( .A(n7505), .B(n9522), .Z(n7354) );
  XNOR U3995 ( .A(n7599), .B(n7354), .Z(out[225]) );
  XOR U3996 ( .A(in[1067]), .B(n8787), .Z(n7611) );
  NOR U3997 ( .A(n7509), .B(n9566), .Z(n7355) );
  XNOR U3998 ( .A(n7611), .B(n7355), .Z(out[226]) );
  XOR U3999 ( .A(in[1068]), .B(n8790), .Z(n7623) );
  NOR U4000 ( .A(n7511), .B(n9610), .Z(n7356) );
  XNOR U4001 ( .A(n7623), .B(n7356), .Z(out[227]) );
  XNOR U4002 ( .A(in[1069]), .B(n8793), .Z(n7636) );
  NAND U4003 ( .A(n7513), .B(n7357), .Z(n7358) );
  XNOR U4004 ( .A(n7636), .B(n7358), .Z(out[228]) );
  XNOR U4005 ( .A(in[1070]), .B(n8796), .Z(n7650) );
  NAND U4006 ( .A(n7515), .B(n7359), .Z(n7360) );
  XNOR U4007 ( .A(n7650), .B(n7360), .Z(out[229]) );
  XNOR U4008 ( .A(in[1432]), .B(n8477), .Z(n9083) );
  NANDN U4009 ( .A(n7477), .B(n9083), .Z(n7361) );
  XNOR U4010 ( .A(n9084), .B(n7361), .Z(out[22]) );
  XNOR U4011 ( .A(in[1071]), .B(n8799), .Z(n7664) );
  NAND U4012 ( .A(n7517), .B(n7362), .Z(n7363) );
  XNOR U4013 ( .A(n7664), .B(n7363), .Z(out[230]) );
  XNOR U4014 ( .A(in[1072]), .B(n8802), .Z(n7678) );
  NAND U4015 ( .A(n7519), .B(n7364), .Z(n7365) );
  XNOR U4016 ( .A(n7678), .B(n7365), .Z(out[231]) );
  XNOR U4017 ( .A(in[1073]), .B(n8805), .Z(n7694) );
  NAND U4018 ( .A(n7521), .B(n7366), .Z(n7367) );
  XNOR U4019 ( .A(n7694), .B(n7367), .Z(out[232]) );
  XNOR U4020 ( .A(in[1074]), .B(n8808), .Z(n7708) );
  NAND U4021 ( .A(n7523), .B(n7368), .Z(n7369) );
  XNOR U4022 ( .A(n7708), .B(n7369), .Z(out[233]) );
  XNOR U4023 ( .A(in[1075]), .B(n8815), .Z(n7722) );
  NAND U4024 ( .A(n7525), .B(n7370), .Z(n7371) );
  XNOR U4025 ( .A(n7722), .B(n7371), .Z(out[234]) );
  XNOR U4026 ( .A(in[1076]), .B(n8818), .Z(n7736) );
  NAND U4027 ( .A(n7527), .B(n7372), .Z(n7373) );
  XNOR U4028 ( .A(n7736), .B(n7373), .Z(out[235]) );
  XNOR U4029 ( .A(in[1077]), .B(n8821), .Z(n7752) );
  NAND U4030 ( .A(n7533), .B(n7374), .Z(n7375) );
  XNOR U4031 ( .A(n7752), .B(n7375), .Z(out[236]) );
  XNOR U4032 ( .A(in[1078]), .B(n8824), .Z(n7776) );
  NAND U4033 ( .A(n7535), .B(n7376), .Z(n7377) );
  XNOR U4034 ( .A(n7776), .B(n7377), .Z(out[237]) );
  XNOR U4035 ( .A(in[1079]), .B(n8827), .Z(n7800) );
  NAND U4036 ( .A(n7537), .B(n7378), .Z(n7379) );
  XNOR U4037 ( .A(n7800), .B(n7379), .Z(out[238]) );
  XNOR U4038 ( .A(in[1080]), .B(n8830), .Z(n7824) );
  NAND U4039 ( .A(n7539), .B(n7380), .Z(n7381) );
  XNOR U4040 ( .A(n7824), .B(n7381), .Z(out[239]) );
  XNOR U4041 ( .A(in[1433]), .B(n8481), .Z(n9107) );
  NANDN U4042 ( .A(n7480), .B(n9107), .Z(n7382) );
  XNOR U4043 ( .A(n9108), .B(n7382), .Z(out[23]) );
  XNOR U4044 ( .A(in[1081]), .B(n8833), .Z(n7848) );
  NAND U4045 ( .A(n7541), .B(n7383), .Z(n7384) );
  XNOR U4046 ( .A(n7848), .B(n7384), .Z(out[240]) );
  XNOR U4047 ( .A(in[1082]), .B(n8836), .Z(n7872) );
  NAND U4048 ( .A(n7543), .B(n7385), .Z(n7386) );
  XNOR U4049 ( .A(n7872), .B(n7386), .Z(out[241]) );
  XNOR U4050 ( .A(in[1083]), .B(n8839), .Z(n7898) );
  NAND U4051 ( .A(n7545), .B(n7387), .Z(n7388) );
  XNOR U4052 ( .A(n7898), .B(n7388), .Z(out[242]) );
  XNOR U4053 ( .A(in[1084]), .B(n8842), .Z(n7922) );
  NAND U4054 ( .A(n7547), .B(n7389), .Z(n7390) );
  XNOR U4055 ( .A(n7922), .B(n7390), .Z(out[243]) );
  XNOR U4056 ( .A(in[1085]), .B(n8849), .Z(n7946) );
  NAND U4057 ( .A(n7549), .B(n7391), .Z(n7392) );
  XNOR U4058 ( .A(n7946), .B(n7392), .Z(out[244]) );
  XNOR U4059 ( .A(in[1086]), .B(n8852), .Z(n7970) );
  NAND U4060 ( .A(n7551), .B(n7393), .Z(n7394) );
  XNOR U4061 ( .A(n7970), .B(n7394), .Z(out[245]) );
  XNOR U4062 ( .A(in[1087]), .B(n8855), .Z(n7994) );
  NAND U4063 ( .A(n7555), .B(n7395), .Z(n7396) );
  XNOR U4064 ( .A(n7994), .B(n7396), .Z(out[246]) );
  XNOR U4065 ( .A(in[1024]), .B(n8858), .Z(n8018) );
  NAND U4066 ( .A(n7557), .B(n7397), .Z(n7398) );
  XNOR U4067 ( .A(n8018), .B(n7398), .Z(out[247]) );
  XNOR U4068 ( .A(in[1025]), .B(n8861), .Z(n8042) );
  NAND U4069 ( .A(n7559), .B(n7399), .Z(n7400) );
  XNOR U4070 ( .A(n8042), .B(n7400), .Z(out[248]) );
  XNOR U4071 ( .A(in[1026]), .B(n8864), .Z(n8074) );
  NAND U4072 ( .A(n7561), .B(n7401), .Z(n7402) );
  XNOR U4073 ( .A(n8074), .B(n7402), .Z(out[249]) );
  XNOR U4074 ( .A(in[1434]), .B(n8485), .Z(n9131) );
  NANDN U4075 ( .A(n7484), .B(n9131), .Z(n7403) );
  XNOR U4076 ( .A(n9132), .B(n7403), .Z(out[24]) );
  XNOR U4077 ( .A(in[1027]), .B(n8867), .Z(n8118) );
  NAND U4078 ( .A(n7563), .B(n7404), .Z(n7405) );
  XNOR U4079 ( .A(n8118), .B(n7405), .Z(out[250]) );
  XNOR U4080 ( .A(in[1028]), .B(n8870), .Z(n8162) );
  NAND U4081 ( .A(n7565), .B(n7406), .Z(n7407) );
  XNOR U4082 ( .A(n8162), .B(n7407), .Z(out[251]) );
  XNOR U4083 ( .A(in[1029]), .B(n8873), .Z(n8208) );
  NAND U4084 ( .A(n7567), .B(n7408), .Z(n7409) );
  XNOR U4085 ( .A(n8208), .B(n7409), .Z(out[252]) );
  XNOR U4086 ( .A(in[1030]), .B(n8876), .Z(n8252) );
  NAND U4087 ( .A(n7569), .B(n7410), .Z(n7411) );
  XNOR U4088 ( .A(n8252), .B(n7411), .Z(out[253]) );
  XNOR U4089 ( .A(in[1031]), .B(n8887), .Z(n8296) );
  NAND U4090 ( .A(n7571), .B(n7412), .Z(n7413) );
  XNOR U4091 ( .A(n8296), .B(n7413), .Z(out[254]) );
  XNOR U4092 ( .A(in[1032]), .B(n8890), .Z(n8340) );
  NAND U4093 ( .A(n7573), .B(n7414), .Z(n7415) );
  XNOR U4094 ( .A(n8340), .B(n7415), .Z(out[255]) );
  ANDN U4095 ( .B(n7417), .A(n7416), .Z(n7418) );
  XNOR U4096 ( .A(n8383), .B(n7418), .Z(out[256]) );
  AND U4097 ( .A(n7420), .B(n7419), .Z(n7421) );
  XNOR U4098 ( .A(n8427), .B(n7421), .Z(out[257]) );
  XOR U4099 ( .A(n8389), .B(in[1412]), .Z(n8472) );
  NAND U4100 ( .A(n7531), .B(n7422), .Z(n7423) );
  XNOR U4101 ( .A(n8472), .B(n7423), .Z(out[258]) );
  XOR U4102 ( .A(n8393), .B(in[1413]), .Z(n8516) );
  NAND U4103 ( .A(n7681), .B(n7424), .Z(n7425) );
  XNOR U4104 ( .A(n8516), .B(n7425), .Z(out[259]) );
  XNOR U4105 ( .A(in[1435]), .B(n8489), .Z(n9163) );
  NANDN U4106 ( .A(n7487), .B(n9163), .Z(n7426) );
  XNOR U4107 ( .A(n9164), .B(n7426), .Z(out[25]) );
  XOR U4108 ( .A(n8397), .B(in[1414]), .Z(n8560) );
  NAND U4109 ( .A(n7875), .B(n7427), .Z(n7428) );
  XNOR U4110 ( .A(n8560), .B(n7428), .Z(out[260]) );
  XOR U4111 ( .A(n8401), .B(in[1415]), .Z(n8604) );
  NAND U4112 ( .A(n8165), .B(n7429), .Z(n7430) );
  XNOR U4113 ( .A(n8604), .B(n7430), .Z(out[261]) );
  XOR U4114 ( .A(n8405), .B(in[1416]), .Z(n8638) );
  NAND U4115 ( .A(n8607), .B(n7431), .Z(n7432) );
  XNOR U4116 ( .A(n8638), .B(n7432), .Z(out[262]) );
  XOR U4117 ( .A(in[1417]), .B(n8409), .Z(n8884) );
  NAND U4118 ( .A(n8883), .B(n7433), .Z(n7434) );
  XNOR U4119 ( .A(n8884), .B(n7434), .Z(out[263]) );
  XOR U4120 ( .A(n8413), .B(in[1418]), .Z(n9168) );
  NAND U4121 ( .A(n9167), .B(n7435), .Z(n7436) );
  XNOR U4122 ( .A(n9168), .B(n7436), .Z(out[264]) );
  XOR U4123 ( .A(n8417), .B(in[1419]), .Z(n9612) );
  NAND U4124 ( .A(n9611), .B(n7437), .Z(n7438) );
  XNOR U4125 ( .A(n9612), .B(n7438), .Z(out[265]) );
  ANDN U4126 ( .B(n7440), .A(n7439), .Z(n7441) );
  XNOR U4127 ( .A(n8727), .B(n7441), .Z(out[266]) );
  ANDN U4128 ( .B(n7443), .A(n7442), .Z(n7444) );
  XNOR U4129 ( .A(n8751), .B(n7444), .Z(out[267]) );
  ANDN U4130 ( .B(n7446), .A(n7445), .Z(n7447) );
  XNOR U4131 ( .A(n8777), .B(n7447), .Z(out[268]) );
  ANDN U4132 ( .B(n7449), .A(n7448), .Z(n7450) );
  XNOR U4133 ( .A(n8811), .B(n7450), .Z(out[269]) );
  XNOR U4134 ( .A(in[1436]), .B(n8493), .Z(n9211) );
  NANDN U4135 ( .A(n7490), .B(n9211), .Z(n7451) );
  XNOR U4136 ( .A(n9212), .B(n7451), .Z(out[26]) );
  ANDN U4137 ( .B(n7453), .A(n7452), .Z(n7454) );
  XNOR U4138 ( .A(n8845), .B(n7454), .Z(out[270]) );
  ANDN U4139 ( .B(n7456), .A(n7455), .Z(n7457) );
  XNOR U4140 ( .A(n8879), .B(n7457), .Z(out[271]) );
  ANDN U4141 ( .B(n7459), .A(n7458), .Z(n7460) );
  XNOR U4142 ( .A(n8917), .B(n7460), .Z(out[272]) );
  ANDN U4143 ( .B(n7462), .A(n7461), .Z(n7463) );
  XNOR U4144 ( .A(n8951), .B(n7463), .Z(out[273]) );
  ANDN U4145 ( .B(n7465), .A(n7464), .Z(n7466) );
  XNOR U4146 ( .A(n8985), .B(n7466), .Z(out[274]) );
  ANDN U4147 ( .B(n7468), .A(n7467), .Z(n7469) );
  XNOR U4148 ( .A(n9011), .B(n7469), .Z(out[275]) );
  ANDN U4149 ( .B(n7471), .A(n7470), .Z(n7472) );
  XNOR U4150 ( .A(n9035), .B(n7472), .Z(out[276]) );
  AND U4151 ( .A(n7474), .B(n7473), .Z(n7475) );
  XNOR U4152 ( .A(n9059), .B(n7475), .Z(out[277]) );
  AND U4153 ( .A(n7477), .B(n7476), .Z(n7478) );
  XNOR U4154 ( .A(n9083), .B(n7478), .Z(out[278]) );
  AND U4155 ( .A(n7480), .B(n7479), .Z(n7481) );
  XNOR U4156 ( .A(n9107), .B(n7481), .Z(out[279]) );
  XNOR U4157 ( .A(in[1437]), .B(n8497), .Z(n9255) );
  NANDN U4158 ( .A(n7493), .B(n9255), .Z(n7482) );
  XNOR U4159 ( .A(n9256), .B(n7482), .Z(out[27]) );
  AND U4160 ( .A(n7484), .B(n7483), .Z(n7485) );
  XNOR U4161 ( .A(n9131), .B(n7485), .Z(out[280]) );
  AND U4162 ( .A(n7487), .B(n7486), .Z(n7488) );
  XNOR U4163 ( .A(n9163), .B(n7488), .Z(out[281]) );
  AND U4164 ( .A(n7490), .B(n7489), .Z(n7491) );
  XNOR U4165 ( .A(n9211), .B(n7491), .Z(out[282]) );
  AND U4166 ( .A(n7493), .B(n7492), .Z(n7494) );
  XNOR U4167 ( .A(n9255), .B(n7494), .Z(out[283]) );
  XOR U4168 ( .A(in[1438]), .B(n8501), .Z(n9300) );
  NAND U4169 ( .A(n7507), .B(n7495), .Z(n7496) );
  XNOR U4170 ( .A(n9300), .B(n7496), .Z(out[284]) );
  XOR U4171 ( .A(in[1439]), .B(n8505), .Z(n9344) );
  NAND U4172 ( .A(n7529), .B(n7497), .Z(n7498) );
  XNOR U4173 ( .A(n9344), .B(n7498), .Z(out[285]) );
  XOR U4174 ( .A(in[1440]), .B(n8509), .Z(n9388) );
  NAND U4175 ( .A(n7553), .B(n7499), .Z(n7500) );
  XNOR U4176 ( .A(n9388), .B(n7500), .Z(out[286]) );
  XOR U4177 ( .A(in[1441]), .B(n8513), .Z(n9432) );
  NAND U4178 ( .A(n7575), .B(n7501), .Z(n7502) );
  XNOR U4179 ( .A(n9432), .B(n7502), .Z(out[287]) );
  XOR U4180 ( .A(in[1442]), .B(n8521), .Z(n9476) );
  NAND U4181 ( .A(n7587), .B(n7503), .Z(n7504) );
  XNOR U4182 ( .A(n9476), .B(n7504), .Z(out[288]) );
  XOR U4183 ( .A(in[1443]), .B(n8525), .Z(n9520) );
  NAND U4184 ( .A(n7599), .B(n7505), .Z(n7506) );
  XNOR U4185 ( .A(n9520), .B(n7506), .Z(out[289]) );
  OR U4186 ( .A(n9300), .B(n7507), .Z(n7508) );
  XNOR U4187 ( .A(n9299), .B(n7508), .Z(out[28]) );
  XOR U4188 ( .A(in[1444]), .B(n8529), .Z(n9564) );
  NAND U4189 ( .A(n7611), .B(n7509), .Z(n7510) );
  XNOR U4190 ( .A(n9564), .B(n7510), .Z(out[290]) );
  XOR U4191 ( .A(in[1445]), .B(n8533), .Z(n9608) );
  NAND U4192 ( .A(n7623), .B(n7511), .Z(n7512) );
  XNOR U4193 ( .A(n9608), .B(n7512), .Z(out[291]) );
  OR U4194 ( .A(n7636), .B(n7513), .Z(n7514) );
  XNOR U4195 ( .A(n7635), .B(n7514), .Z(out[292]) );
  OR U4196 ( .A(n7650), .B(n7515), .Z(n7516) );
  XNOR U4197 ( .A(n7649), .B(n7516), .Z(out[293]) );
  OR U4198 ( .A(n7664), .B(n7517), .Z(n7518) );
  XNOR U4199 ( .A(n7663), .B(n7518), .Z(out[294]) );
  OR U4200 ( .A(n7678), .B(n7519), .Z(n7520) );
  XNOR U4201 ( .A(n7677), .B(n7520), .Z(out[295]) );
  OR U4202 ( .A(n7694), .B(n7521), .Z(n7522) );
  XNOR U4203 ( .A(n7693), .B(n7522), .Z(out[296]) );
  OR U4204 ( .A(n7708), .B(n7523), .Z(n7524) );
  XNOR U4205 ( .A(n7707), .B(n7524), .Z(out[297]) );
  OR U4206 ( .A(n7722), .B(n7525), .Z(n7526) );
  XNOR U4207 ( .A(n7721), .B(n7526), .Z(out[298]) );
  OR U4208 ( .A(n7736), .B(n7527), .Z(n7528) );
  XNOR U4209 ( .A(n7735), .B(n7528), .Z(out[299]) );
  OR U4210 ( .A(n9344), .B(n7529), .Z(n7530) );
  XNOR U4211 ( .A(n9343), .B(n7530), .Z(out[29]) );
  OR U4212 ( .A(n8472), .B(n7531), .Z(n7532) );
  XNOR U4213 ( .A(n8471), .B(n7532), .Z(out[2]) );
  OR U4214 ( .A(n7752), .B(n7533), .Z(n7534) );
  XNOR U4215 ( .A(n7751), .B(n7534), .Z(out[300]) );
  OR U4216 ( .A(n7776), .B(n7535), .Z(n7536) );
  XNOR U4217 ( .A(n7775), .B(n7536), .Z(out[301]) );
  OR U4218 ( .A(n7800), .B(n7537), .Z(n7538) );
  XNOR U4219 ( .A(n7799), .B(n7538), .Z(out[302]) );
  OR U4220 ( .A(n7824), .B(n7539), .Z(n7540) );
  XNOR U4221 ( .A(n7823), .B(n7540), .Z(out[303]) );
  OR U4222 ( .A(n7848), .B(n7541), .Z(n7542) );
  XNOR U4223 ( .A(n7847), .B(n7542), .Z(out[304]) );
  OR U4224 ( .A(n7872), .B(n7543), .Z(n7544) );
  XNOR U4225 ( .A(n7871), .B(n7544), .Z(out[305]) );
  OR U4226 ( .A(n7898), .B(n7545), .Z(n7546) );
  XNOR U4227 ( .A(n7897), .B(n7546), .Z(out[306]) );
  OR U4228 ( .A(n7922), .B(n7547), .Z(n7548) );
  XNOR U4229 ( .A(n7921), .B(n7548), .Z(out[307]) );
  OR U4230 ( .A(n7946), .B(n7549), .Z(n7550) );
  XNOR U4231 ( .A(n7945), .B(n7550), .Z(out[308]) );
  OR U4232 ( .A(n7970), .B(n7551), .Z(n7552) );
  XNOR U4233 ( .A(n7969), .B(n7552), .Z(out[309]) );
  OR U4234 ( .A(n9388), .B(n7553), .Z(n7554) );
  XNOR U4235 ( .A(n9387), .B(n7554), .Z(out[30]) );
  OR U4236 ( .A(n7994), .B(n7555), .Z(n7556) );
  XNOR U4237 ( .A(n7993), .B(n7556), .Z(out[310]) );
  OR U4238 ( .A(n8018), .B(n7557), .Z(n7558) );
  XNOR U4239 ( .A(n8017), .B(n7558), .Z(out[311]) );
  OR U4240 ( .A(n8042), .B(n7559), .Z(n7560) );
  XNOR U4241 ( .A(n8041), .B(n7560), .Z(out[312]) );
  OR U4242 ( .A(n8074), .B(n7561), .Z(n7562) );
  XNOR U4243 ( .A(n8073), .B(n7562), .Z(out[313]) );
  OR U4244 ( .A(n8118), .B(n7563), .Z(n7564) );
  XNOR U4245 ( .A(n8117), .B(n7564), .Z(out[314]) );
  OR U4246 ( .A(n8162), .B(n7565), .Z(n7566) );
  XNOR U4247 ( .A(n8161), .B(n7566), .Z(out[315]) );
  OR U4248 ( .A(n8208), .B(n7567), .Z(n7568) );
  XNOR U4249 ( .A(n8207), .B(n7568), .Z(out[316]) );
  OR U4250 ( .A(n8252), .B(n7569), .Z(n7570) );
  XNOR U4251 ( .A(n8251), .B(n7570), .Z(out[317]) );
  OR U4252 ( .A(n8296), .B(n7571), .Z(n7572) );
  XNOR U4253 ( .A(n8295), .B(n7572), .Z(out[318]) );
  OR U4254 ( .A(n8340), .B(n7573), .Z(n7574) );
  XNOR U4255 ( .A(n8339), .B(n7574), .Z(out[319]) );
  OR U4256 ( .A(n9432), .B(n7575), .Z(n7576) );
  XNOR U4257 ( .A(n9431), .B(n7576), .Z(out[31]) );
  XNOR U4258 ( .A(in[72]), .B(n8890), .Z(n7747) );
  XOR U4259 ( .A(in[1317]), .B(n8725), .Z(n8060) );
  XOR U4260 ( .A(in[1244]), .B(n8543), .Z(n8057) );
  NAND U4261 ( .A(n8060), .B(n8057), .Z(n7577) );
  XNOR U4262 ( .A(n7747), .B(n7577), .Z(out[320]) );
  XNOR U4263 ( .A(in[73]), .B(n8893), .Z(n7749) );
  XOR U4264 ( .A(in[1318]), .B(n8731), .Z(n8064) );
  XOR U4265 ( .A(in[1245]), .B(n8547), .Z(n8061) );
  NAND U4266 ( .A(n8064), .B(n8061), .Z(n7578) );
  XNOR U4267 ( .A(n7749), .B(n7578), .Z(out[321]) );
  XNOR U4268 ( .A(in[74]), .B(n8896), .Z(n7755) );
  XOR U4269 ( .A(in[1319]), .B(n8733), .Z(n8068) );
  XOR U4270 ( .A(in[1246]), .B(n8551), .Z(n8065) );
  NAND U4271 ( .A(n8068), .B(n8065), .Z(n7579) );
  XNOR U4272 ( .A(n7755), .B(n7579), .Z(out[322]) );
  XNOR U4273 ( .A(in[75]), .B(n8899), .Z(n7757) );
  XOR U4274 ( .A(in[1320]), .B(n8735), .Z(n8072) );
  XOR U4275 ( .A(in[1247]), .B(n8555), .Z(n8069) );
  NAND U4276 ( .A(n8072), .B(n8069), .Z(n7580) );
  XNOR U4277 ( .A(n7757), .B(n7580), .Z(out[323]) );
  XOR U4278 ( .A(n8902), .B(in[76]), .Z(n7759) );
  XOR U4279 ( .A(in[1321]), .B(n8737), .Z(n8080) );
  XOR U4280 ( .A(in[1248]), .B(n8563), .Z(n8077) );
  NAND U4281 ( .A(n8080), .B(n8077), .Z(n7581) );
  XNOR U4282 ( .A(n7759), .B(n7581), .Z(out[324]) );
  XOR U4283 ( .A(n8905), .B(in[77]), .Z(n7761) );
  XOR U4284 ( .A(in[1322]), .B(n8739), .Z(n8084) );
  XOR U4285 ( .A(in[1249]), .B(n8567), .Z(n8081) );
  NAND U4286 ( .A(n8084), .B(n8081), .Z(n7582) );
  XNOR U4287 ( .A(n7761), .B(n7582), .Z(out[325]) );
  XOR U4288 ( .A(n8908), .B(in[78]), .Z(n7763) );
  XOR U4289 ( .A(in[1323]), .B(n8741), .Z(n8088) );
  XOR U4290 ( .A(in[1250]), .B(n8571), .Z(n8085) );
  NAND U4291 ( .A(n8088), .B(n8085), .Z(n7583) );
  XNOR U4292 ( .A(n7763), .B(n7583), .Z(out[326]) );
  XOR U4293 ( .A(n8911), .B(in[79]), .Z(n7765) );
  XOR U4294 ( .A(in[1324]), .B(n8743), .Z(n8092) );
  XOR U4295 ( .A(in[1251]), .B(n8575), .Z(n8089) );
  NAND U4296 ( .A(n8092), .B(n8089), .Z(n7584) );
  XNOR U4297 ( .A(n7765), .B(n7584), .Z(out[327]) );
  XOR U4298 ( .A(n8914), .B(in[80]), .Z(n7767) );
  XOR U4299 ( .A(in[1325]), .B(n8745), .Z(n8096) );
  XOR U4300 ( .A(in[1252]), .B(n8579), .Z(n8093) );
  NAND U4301 ( .A(n8096), .B(n8093), .Z(n7585) );
  XNOR U4302 ( .A(n7767), .B(n7585), .Z(out[328]) );
  XOR U4303 ( .A(n8921), .B(in[81]), .Z(n7769) );
  XOR U4304 ( .A(in[1326]), .B(n8747), .Z(n8100) );
  XNOR U4305 ( .A(in[1253]), .B(n8583), .Z(n8097) );
  NAND U4306 ( .A(n8100), .B(n8097), .Z(n7586) );
  XNOR U4307 ( .A(n7769), .B(n7586), .Z(out[329]) );
  OR U4308 ( .A(n9476), .B(n7587), .Z(n7588) );
  XNOR U4309 ( .A(n9475), .B(n7588), .Z(out[32]) );
  XOR U4310 ( .A(n8924), .B(in[82]), .Z(n7771) );
  XOR U4311 ( .A(in[1327]), .B(n8749), .Z(n8104) );
  XNOR U4312 ( .A(in[1254]), .B(n8587), .Z(n8101) );
  NAND U4313 ( .A(n8104), .B(n8101), .Z(n7589) );
  XNOR U4314 ( .A(n7771), .B(n7589), .Z(out[330]) );
  XOR U4315 ( .A(n8927), .B(in[83]), .Z(n7773) );
  XOR U4316 ( .A(in[1328]), .B(n8755), .Z(n8108) );
  XNOR U4317 ( .A(in[1255]), .B(n8591), .Z(n8105) );
  NAND U4318 ( .A(n8108), .B(n8105), .Z(n7590) );
  XNOR U4319 ( .A(n7773), .B(n7590), .Z(out[331]) );
  XOR U4320 ( .A(in[84]), .B(n8930), .Z(n7779) );
  XOR U4321 ( .A(in[1329]), .B(n8757), .Z(n8112) );
  XNOR U4322 ( .A(in[1256]), .B(n8595), .Z(n8109) );
  NAND U4323 ( .A(n8112), .B(n8109), .Z(n7591) );
  XNOR U4324 ( .A(n7779), .B(n7591), .Z(out[332]) );
  XOR U4325 ( .A(in[85]), .B(n8933), .Z(n7781) );
  XOR U4326 ( .A(in[1330]), .B(n8759), .Z(n8116) );
  XNOR U4327 ( .A(in[1257]), .B(n8599), .Z(n8113) );
  NAND U4328 ( .A(n8116), .B(n8113), .Z(n7592) );
  XNOR U4329 ( .A(n7781), .B(n7592), .Z(out[333]) );
  XOR U4330 ( .A(in[86]), .B(n8936), .Z(n7783) );
  XOR U4331 ( .A(in[1331]), .B(n8761), .Z(n8124) );
  XNOR U4332 ( .A(in[1258]), .B(n8609), .Z(n8121) );
  NAND U4333 ( .A(n8124), .B(n8121), .Z(n7593) );
  XNOR U4334 ( .A(n7783), .B(n7593), .Z(out[334]) );
  XOR U4335 ( .A(in[87]), .B(n8939), .Z(n7785) );
  XOR U4336 ( .A(in[1332]), .B(n8763), .Z(n8128) );
  XNOR U4337 ( .A(in[1259]), .B(n8613), .Z(n8125) );
  NAND U4338 ( .A(n8128), .B(n8125), .Z(n7594) );
  XNOR U4339 ( .A(n7785), .B(n7594), .Z(out[335]) );
  XOR U4340 ( .A(in[88]), .B(n8942), .Z(n7787) );
  XOR U4341 ( .A(in[1333]), .B(n8765), .Z(n8132) );
  XNOR U4342 ( .A(in[1260]), .B(n8617), .Z(n8129) );
  NAND U4343 ( .A(n8132), .B(n8129), .Z(n7595) );
  XNOR U4344 ( .A(n7787), .B(n7595), .Z(out[336]) );
  XOR U4345 ( .A(in[89]), .B(n8945), .Z(n7789) );
  XOR U4346 ( .A(in[1334]), .B(n8767), .Z(n8136) );
  XNOR U4347 ( .A(in[1261]), .B(n8621), .Z(n8133) );
  NAND U4348 ( .A(n8136), .B(n8133), .Z(n7596) );
  XNOR U4349 ( .A(n7789), .B(n7596), .Z(out[337]) );
  XOR U4350 ( .A(in[90]), .B(n8948), .Z(n7791) );
  XOR U4351 ( .A(in[1335]), .B(n8769), .Z(n8140) );
  XNOR U4352 ( .A(in[1262]), .B(n8343), .Z(n8137) );
  NAND U4353 ( .A(n8140), .B(n8137), .Z(n7597) );
  XNOR U4354 ( .A(n7791), .B(n7597), .Z(out[338]) );
  XOR U4355 ( .A(in[91]), .B(n8955), .Z(n7793) );
  XOR U4356 ( .A(in[1336]), .B(n8625), .Z(n8144) );
  XNOR U4357 ( .A(in[1263]), .B(n8347), .Z(n8141) );
  NAND U4358 ( .A(n8144), .B(n8141), .Z(n7598) );
  XNOR U4359 ( .A(n7793), .B(n7598), .Z(out[339]) );
  OR U4360 ( .A(n9520), .B(n7599), .Z(n7600) );
  XNOR U4361 ( .A(n9519), .B(n7600), .Z(out[33]) );
  XOR U4362 ( .A(in[92]), .B(n8958), .Z(n7795) );
  XOR U4363 ( .A(in[1337]), .B(n8627), .Z(n8148) );
  XNOR U4364 ( .A(in[1264]), .B(n8351), .Z(n8145) );
  NAND U4365 ( .A(n8148), .B(n8145), .Z(n7601) );
  XNOR U4366 ( .A(n7795), .B(n7601), .Z(out[340]) );
  XOR U4367 ( .A(in[93]), .B(n8961), .Z(n7797) );
  XOR U4368 ( .A(in[1338]), .B(n8629), .Z(n8152) );
  XNOR U4369 ( .A(in[1265]), .B(n8355), .Z(n8149) );
  NAND U4370 ( .A(n8152), .B(n8149), .Z(n7602) );
  XNOR U4371 ( .A(n7797), .B(n7602), .Z(out[341]) );
  XOR U4372 ( .A(in[94]), .B(n8964), .Z(n7803) );
  XOR U4373 ( .A(in[1339]), .B(n8631), .Z(n8156) );
  XNOR U4374 ( .A(in[1266]), .B(n8359), .Z(n8153) );
  NAND U4375 ( .A(n8156), .B(n8153), .Z(n7603) );
  XNOR U4376 ( .A(n7803), .B(n7603), .Z(out[342]) );
  XOR U4377 ( .A(in[95]), .B(n8967), .Z(n7805) );
  XOR U4378 ( .A(in[1340]), .B(n8633), .Z(n8160) );
  XNOR U4379 ( .A(in[1267]), .B(n8363), .Z(n8157) );
  NAND U4380 ( .A(n8160), .B(n8157), .Z(n7604) );
  XNOR U4381 ( .A(n7805), .B(n7604), .Z(out[343]) );
  XOR U4382 ( .A(in[96]), .B(n8970), .Z(n7807) );
  XOR U4383 ( .A(in[1341]), .B(n8635), .Z(n8170) );
  XNOR U4384 ( .A(in[1268]), .B(n8367), .Z(n8167) );
  NAND U4385 ( .A(n8170), .B(n8167), .Z(n7605) );
  XNOR U4386 ( .A(n7807), .B(n7605), .Z(out[344]) );
  XOR U4387 ( .A(in[97]), .B(n8973), .Z(n7809) );
  XOR U4388 ( .A(in[1342]), .B(n8641), .Z(n8174) );
  XNOR U4389 ( .A(in[1269]), .B(n8371), .Z(n8171) );
  NAND U4390 ( .A(n8174), .B(n8171), .Z(n7606) );
  XNOR U4391 ( .A(n7809), .B(n7606), .Z(out[345]) );
  XOR U4392 ( .A(in[98]), .B(n8976), .Z(n7811) );
  XOR U4393 ( .A(in[1343]), .B(n8643), .Z(n8178) );
  XNOR U4394 ( .A(in[1270]), .B(n8375), .Z(n8175) );
  NAND U4395 ( .A(n8178), .B(n8175), .Z(n7607) );
  XNOR U4396 ( .A(n7811), .B(n7607), .Z(out[346]) );
  XOR U4397 ( .A(in[99]), .B(n8979), .Z(n7813) );
  XOR U4398 ( .A(in[1280]), .B(n8645), .Z(n8182) );
  XNOR U4399 ( .A(in[1271]), .B(n8379), .Z(n8179) );
  NAND U4400 ( .A(n8182), .B(n8179), .Z(n7608) );
  XNOR U4401 ( .A(n7813), .B(n7608), .Z(out[347]) );
  XNOR U4402 ( .A(in[100]), .B(n8982), .Z(n7815) );
  XOR U4403 ( .A(in[1281]), .B(n8647), .Z(n8186) );
  XNOR U4404 ( .A(in[1272]), .B(n8387), .Z(n8183) );
  NAND U4405 ( .A(n8186), .B(n8183), .Z(n7609) );
  XNOR U4406 ( .A(n7815), .B(n7609), .Z(out[348]) );
  XNOR U4407 ( .A(in[101]), .B(n8989), .Z(n7817) );
  XOR U4408 ( .A(in[1282]), .B(n8649), .Z(n8190) );
  XNOR U4409 ( .A(in[1273]), .B(n8391), .Z(n8187) );
  NAND U4410 ( .A(n8190), .B(n8187), .Z(n7610) );
  XNOR U4411 ( .A(n7817), .B(n7610), .Z(out[349]) );
  OR U4412 ( .A(n9564), .B(n7611), .Z(n7612) );
  XNOR U4413 ( .A(n9563), .B(n7612), .Z(out[34]) );
  XNOR U4414 ( .A(in[102]), .B(n8992), .Z(n7819) );
  XOR U4415 ( .A(in[1283]), .B(n8651), .Z(n8194) );
  XNOR U4416 ( .A(in[1274]), .B(n8395), .Z(n8191) );
  NAND U4417 ( .A(n8194), .B(n8191), .Z(n7613) );
  XNOR U4418 ( .A(n7819), .B(n7613), .Z(out[350]) );
  XNOR U4419 ( .A(in[103]), .B(n8771), .Z(n7821) );
  XOR U4420 ( .A(in[1284]), .B(n8653), .Z(n8198) );
  XNOR U4421 ( .A(in[1275]), .B(n8399), .Z(n8195) );
  NAND U4422 ( .A(n8198), .B(n8195), .Z(n7614) );
  XNOR U4423 ( .A(n7821), .B(n7614), .Z(out[351]) );
  XNOR U4424 ( .A(in[104]), .B(n8774), .Z(n7827) );
  XOR U4425 ( .A(in[1285]), .B(n8655), .Z(n8202) );
  XNOR U4426 ( .A(in[1276]), .B(n8403), .Z(n8199) );
  NAND U4427 ( .A(n8202), .B(n8199), .Z(n7615) );
  XNOR U4428 ( .A(n7827), .B(n7615), .Z(out[352]) );
  XNOR U4429 ( .A(in[105]), .B(n8781), .Z(n7829) );
  XOR U4430 ( .A(in[1286]), .B(n8657), .Z(n8206) );
  XNOR U4431 ( .A(in[1277]), .B(n8407), .Z(n8203) );
  NAND U4432 ( .A(n8206), .B(n8203), .Z(n7616) );
  XNOR U4433 ( .A(n7829), .B(n7616), .Z(out[353]) );
  XNOR U4434 ( .A(in[106]), .B(n8784), .Z(n7831) );
  XOR U4435 ( .A(in[1287]), .B(n8659), .Z(n8214) );
  XNOR U4436 ( .A(in[1278]), .B(n8411), .Z(n8211) );
  NAND U4437 ( .A(n8214), .B(n8211), .Z(n7617) );
  XNOR U4438 ( .A(n7831), .B(n7617), .Z(out[354]) );
  XNOR U4439 ( .A(in[107]), .B(n8787), .Z(n7833) );
  XOR U4440 ( .A(in[1288]), .B(n8663), .Z(n8218) );
  XNOR U4441 ( .A(in[1279]), .B(n8415), .Z(n8215) );
  NAND U4442 ( .A(n8218), .B(n8215), .Z(n7618) );
  XNOR U4443 ( .A(n7833), .B(n7618), .Z(out[355]) );
  XNOR U4444 ( .A(in[108]), .B(n8790), .Z(n7835) );
  XOR U4445 ( .A(in[1289]), .B(n8665), .Z(n8222) );
  XNOR U4446 ( .A(in[1216]), .B(n8419), .Z(n8219) );
  NAND U4447 ( .A(n8222), .B(n8219), .Z(n7619) );
  XNOR U4448 ( .A(n7835), .B(n7619), .Z(out[356]) );
  XNOR U4449 ( .A(in[109]), .B(n8793), .Z(n7837) );
  XOR U4450 ( .A(in[1290]), .B(n8667), .Z(n8226) );
  XNOR U4451 ( .A(in[1217]), .B(n8423), .Z(n8223) );
  NAND U4452 ( .A(n8226), .B(n8223), .Z(n7620) );
  XNOR U4453 ( .A(n7837), .B(n7620), .Z(out[357]) );
  XNOR U4454 ( .A(in[110]), .B(n8796), .Z(n7839) );
  XOR U4455 ( .A(in[1291]), .B(n8669), .Z(n8230) );
  XNOR U4456 ( .A(in[1218]), .B(n8431), .Z(n8227) );
  NAND U4457 ( .A(n8230), .B(n8227), .Z(n7621) );
  XNOR U4458 ( .A(n7839), .B(n7621), .Z(out[358]) );
  XNOR U4459 ( .A(in[111]), .B(n8799), .Z(n7841) );
  XOR U4460 ( .A(in[1292]), .B(n8671), .Z(n8234) );
  XNOR U4461 ( .A(in[1219]), .B(n8435), .Z(n8231) );
  NAND U4462 ( .A(n8234), .B(n8231), .Z(n7622) );
  XNOR U4463 ( .A(n7841), .B(n7622), .Z(out[359]) );
  OR U4464 ( .A(n9608), .B(n7623), .Z(n7624) );
  XNOR U4465 ( .A(n9607), .B(n7624), .Z(out[35]) );
  XNOR U4466 ( .A(in[112]), .B(n8802), .Z(n7843) );
  XOR U4467 ( .A(in[1293]), .B(n8673), .Z(n8238) );
  XOR U4468 ( .A(in[1220]), .B(n8439), .Z(n8235) );
  NAND U4469 ( .A(n8238), .B(n8235), .Z(n7625) );
  XNOR U4470 ( .A(n7843), .B(n7625), .Z(out[360]) );
  XNOR U4471 ( .A(in[113]), .B(n8805), .Z(n7845) );
  XOR U4472 ( .A(in[1294]), .B(n8675), .Z(n8242) );
  XOR U4473 ( .A(in[1221]), .B(n8443), .Z(n8239) );
  NAND U4474 ( .A(n8242), .B(n8239), .Z(n7626) );
  XNOR U4475 ( .A(n7845), .B(n7626), .Z(out[361]) );
  XNOR U4476 ( .A(in[114]), .B(n8808), .Z(n7851) );
  XOR U4477 ( .A(in[1295]), .B(n8677), .Z(n8246) );
  XOR U4478 ( .A(in[1222]), .B(n8447), .Z(n8243) );
  NAND U4479 ( .A(n8246), .B(n8243), .Z(n7627) );
  XNOR U4480 ( .A(n7851), .B(n7627), .Z(out[362]) );
  XNOR U4481 ( .A(in[115]), .B(n8815), .Z(n7853) );
  XOR U4482 ( .A(in[1296]), .B(n8679), .Z(n8250) );
  XOR U4483 ( .A(in[1223]), .B(n8451), .Z(n8247) );
  NAND U4484 ( .A(n8250), .B(n8247), .Z(n7628) );
  XNOR U4485 ( .A(n7853), .B(n7628), .Z(out[363]) );
  XNOR U4486 ( .A(in[116]), .B(n8818), .Z(n7855) );
  XOR U4487 ( .A(in[1297]), .B(n8681), .Z(n8258) );
  XOR U4488 ( .A(in[1224]), .B(n8455), .Z(n8255) );
  NAND U4489 ( .A(n8258), .B(n8255), .Z(n7629) );
  XNOR U4490 ( .A(n7855), .B(n7629), .Z(out[364]) );
  XNOR U4491 ( .A(in[117]), .B(n8821), .Z(n7857) );
  XOR U4492 ( .A(in[1298]), .B(n8685), .Z(n8262) );
  XOR U4493 ( .A(in[1225]), .B(n8459), .Z(n8259) );
  NAND U4494 ( .A(n8262), .B(n8259), .Z(n7630) );
  XNOR U4495 ( .A(n7857), .B(n7630), .Z(out[365]) );
  XNOR U4496 ( .A(in[118]), .B(n8824), .Z(n7859) );
  XOR U4497 ( .A(in[1299]), .B(n8687), .Z(n8266) );
  XOR U4498 ( .A(in[1226]), .B(n8463), .Z(n8263) );
  NAND U4499 ( .A(n8266), .B(n8263), .Z(n7631) );
  XNOR U4500 ( .A(n7859), .B(n7631), .Z(out[366]) );
  XNOR U4501 ( .A(in[119]), .B(n8827), .Z(n7861) );
  XOR U4502 ( .A(in[1300]), .B(n8689), .Z(n8270) );
  XOR U4503 ( .A(in[1227]), .B(n8467), .Z(n8267) );
  NAND U4504 ( .A(n8270), .B(n8267), .Z(n7632) );
  XNOR U4505 ( .A(n7861), .B(n7632), .Z(out[367]) );
  XNOR U4506 ( .A(in[120]), .B(n8830), .Z(n7863) );
  XOR U4507 ( .A(in[1301]), .B(n8691), .Z(n8274) );
  XOR U4508 ( .A(in[1228]), .B(n8475), .Z(n8271) );
  NAND U4509 ( .A(n8274), .B(n8271), .Z(n7633) );
  XNOR U4510 ( .A(n7863), .B(n7633), .Z(out[368]) );
  XNOR U4511 ( .A(in[121]), .B(n8833), .Z(n7865) );
  XOR U4512 ( .A(in[1302]), .B(n8693), .Z(n8278) );
  XOR U4513 ( .A(in[1229]), .B(n8479), .Z(n8275) );
  NAND U4514 ( .A(n8278), .B(n8275), .Z(n7634) );
  XNOR U4515 ( .A(n7865), .B(n7634), .Z(out[369]) );
  ANDN U4516 ( .B(n7636), .A(n7635), .Z(n7637) );
  XNOR U4517 ( .A(n7638), .B(n7637), .Z(out[36]) );
  XNOR U4518 ( .A(in[122]), .B(n8836), .Z(n7867) );
  XOR U4519 ( .A(in[1303]), .B(n8695), .Z(n8282) );
  XOR U4520 ( .A(in[1230]), .B(n8483), .Z(n8279) );
  NAND U4521 ( .A(n8282), .B(n8279), .Z(n7639) );
  XNOR U4522 ( .A(n7867), .B(n7639), .Z(out[370]) );
  XNOR U4523 ( .A(in[123]), .B(n8839), .Z(n7869) );
  XOR U4524 ( .A(in[1304]), .B(n8697), .Z(n8286) );
  XOR U4525 ( .A(in[1231]), .B(n8487), .Z(n8283) );
  NAND U4526 ( .A(n8286), .B(n8283), .Z(n7640) );
  XNOR U4527 ( .A(n7869), .B(n7640), .Z(out[371]) );
  XNOR U4528 ( .A(in[124]), .B(n8842), .Z(n7877) );
  XOR U4529 ( .A(in[1305]), .B(n8699), .Z(n8290) );
  XOR U4530 ( .A(in[1232]), .B(n8491), .Z(n8287) );
  NAND U4531 ( .A(n8290), .B(n8287), .Z(n7641) );
  XNOR U4532 ( .A(n7877), .B(n7641), .Z(out[372]) );
  XNOR U4533 ( .A(in[125]), .B(n8849), .Z(n7879) );
  XOR U4534 ( .A(in[1306]), .B(n8701), .Z(n8294) );
  XOR U4535 ( .A(in[1233]), .B(n8495), .Z(n8291) );
  NAND U4536 ( .A(n8294), .B(n8291), .Z(n7642) );
  XNOR U4537 ( .A(n7879), .B(n7642), .Z(out[373]) );
  XNOR U4538 ( .A(in[126]), .B(n8852), .Z(n7881) );
  XOR U4539 ( .A(in[1307]), .B(n8703), .Z(n8302) );
  XOR U4540 ( .A(in[1234]), .B(n8499), .Z(n8299) );
  NAND U4541 ( .A(n8302), .B(n8299), .Z(n7643) );
  XNOR U4542 ( .A(n7881), .B(n7643), .Z(out[374]) );
  XNOR U4543 ( .A(in[127]), .B(n8855), .Z(n7883) );
  XOR U4544 ( .A(in[1308]), .B(n8707), .Z(n8306) );
  XOR U4545 ( .A(in[1235]), .B(n8503), .Z(n8303) );
  NAND U4546 ( .A(n8306), .B(n8303), .Z(n7644) );
  XNOR U4547 ( .A(n7883), .B(n7644), .Z(out[375]) );
  XNOR U4548 ( .A(in[64]), .B(n8858), .Z(n7885) );
  XOR U4549 ( .A(in[1309]), .B(n8709), .Z(n8310) );
  XOR U4550 ( .A(in[1236]), .B(n8507), .Z(n8307) );
  NAND U4551 ( .A(n8310), .B(n8307), .Z(n7645) );
  XNOR U4552 ( .A(n7885), .B(n7645), .Z(out[376]) );
  XNOR U4553 ( .A(in[65]), .B(n8861), .Z(n7887) );
  XOR U4554 ( .A(in[1310]), .B(n8711), .Z(n8314) );
  XOR U4555 ( .A(in[1237]), .B(n8511), .Z(n8311) );
  NAND U4556 ( .A(n8314), .B(n8311), .Z(n7646) );
  XNOR U4557 ( .A(n7887), .B(n7646), .Z(out[377]) );
  XNOR U4558 ( .A(in[66]), .B(n8864), .Z(n7889) );
  XOR U4559 ( .A(in[1311]), .B(n8713), .Z(n8318) );
  XOR U4560 ( .A(in[1238]), .B(n8519), .Z(n8315) );
  NAND U4561 ( .A(n8318), .B(n8315), .Z(n7647) );
  XNOR U4562 ( .A(n7889), .B(n7647), .Z(out[378]) );
  XNOR U4563 ( .A(in[67]), .B(n8867), .Z(n7891) );
  XOR U4564 ( .A(in[1312]), .B(n8715), .Z(n8322) );
  XOR U4565 ( .A(in[1239]), .B(n8523), .Z(n8319) );
  NAND U4566 ( .A(n8322), .B(n8319), .Z(n7648) );
  XNOR U4567 ( .A(n7891), .B(n7648), .Z(out[379]) );
  ANDN U4568 ( .B(n7650), .A(n7649), .Z(n7651) );
  XNOR U4569 ( .A(n7652), .B(n7651), .Z(out[37]) );
  XNOR U4570 ( .A(in[68]), .B(n8870), .Z(n7893) );
  XOR U4571 ( .A(in[1313]), .B(n8717), .Z(n8326) );
  XOR U4572 ( .A(in[1240]), .B(n8527), .Z(n8323) );
  NAND U4573 ( .A(n8326), .B(n8323), .Z(n7653) );
  XNOR U4574 ( .A(n7893), .B(n7653), .Z(out[380]) );
  XNOR U4575 ( .A(in[69]), .B(n8873), .Z(n7895) );
  XOR U4576 ( .A(in[1314]), .B(n8719), .Z(n8330) );
  XOR U4577 ( .A(in[1241]), .B(n8531), .Z(n8327) );
  NAND U4578 ( .A(n8330), .B(n8327), .Z(n7654) );
  XNOR U4579 ( .A(n7895), .B(n7654), .Z(out[381]) );
  XNOR U4580 ( .A(in[70]), .B(n8876), .Z(n7901) );
  XOR U4581 ( .A(in[1315]), .B(n8721), .Z(n8334) );
  XOR U4582 ( .A(in[1242]), .B(n8535), .Z(n8331) );
  NAND U4583 ( .A(n8334), .B(n8331), .Z(n7655) );
  XNOR U4584 ( .A(n7901), .B(n7655), .Z(out[382]) );
  XNOR U4585 ( .A(in[71]), .B(n8887), .Z(n7903) );
  XOR U4586 ( .A(in[1316]), .B(n8723), .Z(n8338) );
  XOR U4587 ( .A(in[1243]), .B(n8539), .Z(n8335) );
  NAND U4588 ( .A(n8338), .B(n8335), .Z(n7656) );
  XNOR U4589 ( .A(n7903), .B(n7656), .Z(out[383]) );
  XOR U4590 ( .A(in[497]), .B(n8585), .Z(n7905) );
  NOR U4591 ( .A(n7747), .B(n8060), .Z(n7657) );
  XNOR U4592 ( .A(n7905), .B(n7657), .Z(out[384]) );
  XOR U4593 ( .A(in[498]), .B(n8589), .Z(n7907) );
  NOR U4594 ( .A(n7749), .B(n8064), .Z(n7658) );
  XNOR U4595 ( .A(n7907), .B(n7658), .Z(out[385]) );
  XOR U4596 ( .A(in[499]), .B(n8593), .Z(n7909) );
  NOR U4597 ( .A(n7755), .B(n8068), .Z(n7659) );
  XNOR U4598 ( .A(n7909), .B(n7659), .Z(out[386]) );
  XOR U4599 ( .A(in[500]), .B(n8597), .Z(n7911) );
  NOR U4600 ( .A(n7757), .B(n8072), .Z(n7660) );
  XNOR U4601 ( .A(n7911), .B(n7660), .Z(out[387]) );
  XOR U4602 ( .A(in[501]), .B(n8601), .Z(n7913) );
  NOR U4603 ( .A(n7759), .B(n8080), .Z(n7661) );
  XNOR U4604 ( .A(n7913), .B(n7661), .Z(out[388]) );
  XOR U4605 ( .A(in[502]), .B(n8611), .Z(n7915) );
  NOR U4606 ( .A(n7761), .B(n8084), .Z(n7662) );
  XNOR U4607 ( .A(n7915), .B(n7662), .Z(out[389]) );
  ANDN U4608 ( .B(n7664), .A(n7663), .Z(n7665) );
  XNOR U4609 ( .A(n7666), .B(n7665), .Z(out[38]) );
  XOR U4610 ( .A(in[503]), .B(n8615), .Z(n7917) );
  NOR U4611 ( .A(n7763), .B(n8088), .Z(n7667) );
  XNOR U4612 ( .A(n7917), .B(n7667), .Z(out[390]) );
  XOR U4613 ( .A(in[504]), .B(n8619), .Z(n7919) );
  NOR U4614 ( .A(n7765), .B(n8092), .Z(n7668) );
  XNOR U4615 ( .A(n7919), .B(n7668), .Z(out[391]) );
  XOR U4616 ( .A(in[505]), .B(n8623), .Z(n7925) );
  NOR U4617 ( .A(n7767), .B(n8096), .Z(n7669) );
  XNOR U4618 ( .A(n7925), .B(n7669), .Z(out[392]) );
  XOR U4619 ( .A(in[506]), .B(n8345), .Z(n7927) );
  NOR U4620 ( .A(n7769), .B(n8100), .Z(n7670) );
  XNOR U4621 ( .A(n7927), .B(n7670), .Z(out[393]) );
  XOR U4622 ( .A(in[507]), .B(n8349), .Z(n7929) );
  NOR U4623 ( .A(n7771), .B(n8104), .Z(n7671) );
  XNOR U4624 ( .A(n7929), .B(n7671), .Z(out[394]) );
  XOR U4625 ( .A(in[508]), .B(n8353), .Z(n7931) );
  NOR U4626 ( .A(n7773), .B(n8108), .Z(n7672) );
  XNOR U4627 ( .A(n7931), .B(n7672), .Z(out[395]) );
  XOR U4628 ( .A(in[509]), .B(n8357), .Z(n7933) );
  NOR U4629 ( .A(n7779), .B(n8112), .Z(n7673) );
  XNOR U4630 ( .A(n7933), .B(n7673), .Z(out[396]) );
  XOR U4631 ( .A(in[510]), .B(n8361), .Z(n7935) );
  NOR U4632 ( .A(n7781), .B(n8116), .Z(n7674) );
  XNOR U4633 ( .A(n7935), .B(n7674), .Z(out[397]) );
  XOR U4634 ( .A(in[511]), .B(n8365), .Z(n7937) );
  NOR U4635 ( .A(n7783), .B(n8124), .Z(n7675) );
  XNOR U4636 ( .A(n7937), .B(n7675), .Z(out[398]) );
  XOR U4637 ( .A(in[448]), .B(n8369), .Z(n7939) );
  NOR U4638 ( .A(n7785), .B(n8128), .Z(n7676) );
  XNOR U4639 ( .A(n7939), .B(n7676), .Z(out[399]) );
  ANDN U4640 ( .B(n7678), .A(n7677), .Z(n7679) );
  XNOR U4641 ( .A(n7680), .B(n7679), .Z(out[39]) );
  OR U4642 ( .A(n8516), .B(n7681), .Z(n7682) );
  XNOR U4643 ( .A(n8515), .B(n7682), .Z(out[3]) );
  XOR U4644 ( .A(in[449]), .B(n8373), .Z(n7941) );
  NOR U4645 ( .A(n7787), .B(n8132), .Z(n7683) );
  XNOR U4646 ( .A(n7941), .B(n7683), .Z(out[400]) );
  XNOR U4647 ( .A(n8377), .B(in[450]), .Z(n7943) );
  NOR U4648 ( .A(n7789), .B(n8136), .Z(n7684) );
  XNOR U4649 ( .A(n7943), .B(n7684), .Z(out[401]) );
  XNOR U4650 ( .A(n8381), .B(in[451]), .Z(n7949) );
  NOR U4651 ( .A(n7791), .B(n8140), .Z(n7685) );
  XNOR U4652 ( .A(n7949), .B(n7685), .Z(out[402]) );
  XNOR U4653 ( .A(n8389), .B(in[452]), .Z(n7951) );
  NOR U4654 ( .A(n7793), .B(n8144), .Z(n7686) );
  XNOR U4655 ( .A(n7951), .B(n7686), .Z(out[403]) );
  XNOR U4656 ( .A(n8393), .B(in[453]), .Z(n7953) );
  NOR U4657 ( .A(n7795), .B(n8148), .Z(n7687) );
  XNOR U4658 ( .A(n7953), .B(n7687), .Z(out[404]) );
  XNOR U4659 ( .A(n8397), .B(in[454]), .Z(n7955) );
  NOR U4660 ( .A(n7797), .B(n8152), .Z(n7688) );
  XNOR U4661 ( .A(n7955), .B(n7688), .Z(out[405]) );
  XNOR U4662 ( .A(n8401), .B(in[455]), .Z(n7957) );
  NOR U4663 ( .A(n7803), .B(n8156), .Z(n7689) );
  XNOR U4664 ( .A(n7957), .B(n7689), .Z(out[406]) );
  XNOR U4665 ( .A(n8405), .B(in[456]), .Z(n7959) );
  NOR U4666 ( .A(n7805), .B(n8160), .Z(n7690) );
  XNOR U4667 ( .A(n7959), .B(n7690), .Z(out[407]) );
  XNOR U4668 ( .A(in[457]), .B(n8409), .Z(n7961) );
  NOR U4669 ( .A(n7807), .B(n8170), .Z(n7691) );
  XNOR U4670 ( .A(n7961), .B(n7691), .Z(out[408]) );
  XNOR U4671 ( .A(n8413), .B(in[458]), .Z(n7963) );
  NOR U4672 ( .A(n7809), .B(n8174), .Z(n7692) );
  XNOR U4673 ( .A(n7963), .B(n7692), .Z(out[409]) );
  ANDN U4674 ( .B(n7694), .A(n7693), .Z(n7695) );
  XNOR U4675 ( .A(n7696), .B(n7695), .Z(out[40]) );
  XNOR U4676 ( .A(n8417), .B(in[459]), .Z(n7965) );
  NOR U4677 ( .A(n7811), .B(n8178), .Z(n7697) );
  XNOR U4678 ( .A(n7965), .B(n7697), .Z(out[410]) );
  XNOR U4679 ( .A(in[460]), .B(n8421), .Z(n7967) );
  NOR U4680 ( .A(n7813), .B(n8182), .Z(n7698) );
  XNOR U4681 ( .A(n7967), .B(n7698), .Z(out[411]) );
  XNOR U4682 ( .A(in[461]), .B(n8425), .Z(n7973) );
  NOR U4683 ( .A(n7815), .B(n8186), .Z(n7699) );
  XNOR U4684 ( .A(n7973), .B(n7699), .Z(out[412]) );
  XNOR U4685 ( .A(in[462]), .B(n8433), .Z(n7975) );
  NOR U4686 ( .A(n7817), .B(n8190), .Z(n7700) );
  XNOR U4687 ( .A(n7975), .B(n7700), .Z(out[413]) );
  XNOR U4688 ( .A(in[463]), .B(n8437), .Z(n7977) );
  NOR U4689 ( .A(n7819), .B(n8194), .Z(n7701) );
  XNOR U4690 ( .A(n7977), .B(n7701), .Z(out[414]) );
  XNOR U4691 ( .A(in[464]), .B(n8441), .Z(n7979) );
  NOR U4692 ( .A(n7821), .B(n8198), .Z(n7702) );
  XNOR U4693 ( .A(n7979), .B(n7702), .Z(out[415]) );
  XNOR U4694 ( .A(in[465]), .B(n8445), .Z(n7981) );
  NOR U4695 ( .A(n7827), .B(n8202), .Z(n7703) );
  XNOR U4696 ( .A(n7981), .B(n7703), .Z(out[416]) );
  XNOR U4697 ( .A(in[466]), .B(n8449), .Z(n7983) );
  NOR U4698 ( .A(n7829), .B(n8206), .Z(n7704) );
  XNOR U4699 ( .A(n7983), .B(n7704), .Z(out[417]) );
  XNOR U4700 ( .A(in[467]), .B(n8453), .Z(n7985) );
  NOR U4701 ( .A(n7831), .B(n8214), .Z(n7705) );
  XNOR U4702 ( .A(n7985), .B(n7705), .Z(out[418]) );
  XNOR U4703 ( .A(in[468]), .B(n8457), .Z(n7987) );
  NOR U4704 ( .A(n7833), .B(n8218), .Z(n7706) );
  XNOR U4705 ( .A(n7987), .B(n7706), .Z(out[419]) );
  ANDN U4706 ( .B(n7708), .A(n7707), .Z(n7709) );
  XNOR U4707 ( .A(n7710), .B(n7709), .Z(out[41]) );
  XNOR U4708 ( .A(in[469]), .B(n8461), .Z(n7989) );
  NOR U4709 ( .A(n7835), .B(n8222), .Z(n7711) );
  XNOR U4710 ( .A(n7989), .B(n7711), .Z(out[420]) );
  XNOR U4711 ( .A(in[470]), .B(n8465), .Z(n7991) );
  NOR U4712 ( .A(n7837), .B(n8226), .Z(n7712) );
  XNOR U4713 ( .A(n7991), .B(n7712), .Z(out[421]) );
  XNOR U4714 ( .A(in[471]), .B(n8469), .Z(n7997) );
  NOR U4715 ( .A(n7839), .B(n8230), .Z(n7713) );
  XNOR U4716 ( .A(n7997), .B(n7713), .Z(out[422]) );
  XNOR U4717 ( .A(in[472]), .B(n8477), .Z(n7999) );
  NOR U4718 ( .A(n7841), .B(n8234), .Z(n7714) );
  XNOR U4719 ( .A(n7999), .B(n7714), .Z(out[423]) );
  XNOR U4720 ( .A(in[473]), .B(n8481), .Z(n8001) );
  NOR U4721 ( .A(n7843), .B(n8238), .Z(n7715) );
  XNOR U4722 ( .A(n8001), .B(n7715), .Z(out[424]) );
  XNOR U4723 ( .A(in[474]), .B(n8485), .Z(n8003) );
  NOR U4724 ( .A(n7845), .B(n8242), .Z(n7716) );
  XNOR U4725 ( .A(n8003), .B(n7716), .Z(out[425]) );
  XNOR U4726 ( .A(in[475]), .B(n8489), .Z(n8005) );
  NOR U4727 ( .A(n7851), .B(n8246), .Z(n7717) );
  XNOR U4728 ( .A(n8005), .B(n7717), .Z(out[426]) );
  XNOR U4729 ( .A(in[476]), .B(n8493), .Z(n8007) );
  NOR U4730 ( .A(n7853), .B(n8250), .Z(n7718) );
  XNOR U4731 ( .A(n8007), .B(n7718), .Z(out[427]) );
  XNOR U4732 ( .A(in[477]), .B(n8497), .Z(n8009) );
  NOR U4733 ( .A(n7855), .B(n8258), .Z(n7719) );
  XNOR U4734 ( .A(n8009), .B(n7719), .Z(out[428]) );
  XNOR U4735 ( .A(in[478]), .B(n8501), .Z(n8011) );
  NOR U4736 ( .A(n7857), .B(n8262), .Z(n7720) );
  XNOR U4737 ( .A(n8011), .B(n7720), .Z(out[429]) );
  ANDN U4738 ( .B(n7722), .A(n7721), .Z(n7723) );
  XNOR U4739 ( .A(n7724), .B(n7723), .Z(out[42]) );
  XNOR U4740 ( .A(in[479]), .B(n8505), .Z(n8013) );
  NOR U4741 ( .A(n7859), .B(n8266), .Z(n7725) );
  XNOR U4742 ( .A(n8013), .B(n7725), .Z(out[430]) );
  XNOR U4743 ( .A(in[480]), .B(n8509), .Z(n8015) );
  NOR U4744 ( .A(n7861), .B(n8270), .Z(n7726) );
  XNOR U4745 ( .A(n8015), .B(n7726), .Z(out[431]) );
  XNOR U4746 ( .A(in[481]), .B(n8513), .Z(n8021) );
  NOR U4747 ( .A(n7863), .B(n8274), .Z(n7727) );
  XNOR U4748 ( .A(n8021), .B(n7727), .Z(out[432]) );
  XNOR U4749 ( .A(in[482]), .B(n8521), .Z(n8023) );
  NOR U4750 ( .A(n7865), .B(n8278), .Z(n7728) );
  XNOR U4751 ( .A(n8023), .B(n7728), .Z(out[433]) );
  XNOR U4752 ( .A(in[483]), .B(n8525), .Z(n8025) );
  NOR U4753 ( .A(n7867), .B(n8282), .Z(n7729) );
  XNOR U4754 ( .A(n8025), .B(n7729), .Z(out[434]) );
  XNOR U4755 ( .A(in[484]), .B(n8529), .Z(n8027) );
  NOR U4756 ( .A(n7869), .B(n8286), .Z(n7730) );
  XNOR U4757 ( .A(n8027), .B(n7730), .Z(out[435]) );
  XNOR U4758 ( .A(in[485]), .B(n8533), .Z(n8029) );
  NOR U4759 ( .A(n7877), .B(n8290), .Z(n7731) );
  XNOR U4760 ( .A(n8029), .B(n7731), .Z(out[436]) );
  XOR U4761 ( .A(in[486]), .B(n8537), .Z(n8031) );
  NOR U4762 ( .A(n7879), .B(n8294), .Z(n7732) );
  XNOR U4763 ( .A(n8031), .B(n7732), .Z(out[437]) );
  XOR U4764 ( .A(in[487]), .B(n8541), .Z(n8033) );
  NOR U4765 ( .A(n7881), .B(n8302), .Z(n7733) );
  XNOR U4766 ( .A(n8033), .B(n7733), .Z(out[438]) );
  XOR U4767 ( .A(in[488]), .B(n8545), .Z(n8035) );
  NOR U4768 ( .A(n7883), .B(n8306), .Z(n7734) );
  XNOR U4769 ( .A(n8035), .B(n7734), .Z(out[439]) );
  ANDN U4770 ( .B(n7736), .A(n7735), .Z(n7737) );
  XNOR U4771 ( .A(n7738), .B(n7737), .Z(out[43]) );
  XOR U4772 ( .A(in[489]), .B(n8549), .Z(n8037) );
  NOR U4773 ( .A(n7885), .B(n8310), .Z(n7739) );
  XNOR U4774 ( .A(n8037), .B(n7739), .Z(out[440]) );
  XOR U4775 ( .A(in[490]), .B(n8553), .Z(n8039) );
  NOR U4776 ( .A(n7887), .B(n8314), .Z(n7740) );
  XNOR U4777 ( .A(n8039), .B(n7740), .Z(out[441]) );
  XOR U4778 ( .A(in[491]), .B(n8557), .Z(n8045) );
  NOR U4779 ( .A(n7889), .B(n8318), .Z(n7741) );
  XNOR U4780 ( .A(n8045), .B(n7741), .Z(out[442]) );
  XOR U4781 ( .A(in[492]), .B(n8565), .Z(n8047) );
  NOR U4782 ( .A(n7891), .B(n8322), .Z(n7742) );
  XNOR U4783 ( .A(n8047), .B(n7742), .Z(out[443]) );
  XOR U4784 ( .A(in[493]), .B(n8569), .Z(n8049) );
  NOR U4785 ( .A(n7893), .B(n8326), .Z(n7743) );
  XNOR U4786 ( .A(n8049), .B(n7743), .Z(out[444]) );
  XOR U4787 ( .A(in[494]), .B(n8573), .Z(n8051) );
  NOR U4788 ( .A(n7895), .B(n8330), .Z(n7744) );
  XNOR U4789 ( .A(n8051), .B(n7744), .Z(out[445]) );
  XOR U4790 ( .A(in[495]), .B(n8577), .Z(n8053) );
  NOR U4791 ( .A(n7901), .B(n8334), .Z(n7745) );
  XNOR U4792 ( .A(n8053), .B(n7745), .Z(out[446]) );
  XOR U4793 ( .A(in[496]), .B(n8581), .Z(n8055) );
  NOR U4794 ( .A(n7903), .B(n8338), .Z(n7746) );
  XNOR U4795 ( .A(n8055), .B(n7746), .Z(out[447]) );
  XNOR U4796 ( .A(in[886]), .B(n8584), .Z(n8058) );
  NAND U4797 ( .A(n7905), .B(n7747), .Z(n7748) );
  XNOR U4798 ( .A(n8058), .B(n7748), .Z(out[448]) );
  XNOR U4799 ( .A(in[887]), .B(n8588), .Z(n8062) );
  NAND U4800 ( .A(n7907), .B(n7749), .Z(n7750) );
  XNOR U4801 ( .A(n8062), .B(n7750), .Z(out[449]) );
  ANDN U4802 ( .B(n7752), .A(n7751), .Z(n7753) );
  XNOR U4803 ( .A(n7754), .B(n7753), .Z(out[44]) );
  XNOR U4804 ( .A(in[888]), .B(n8592), .Z(n8066) );
  NAND U4805 ( .A(n7909), .B(n7755), .Z(n7756) );
  XNOR U4806 ( .A(n8066), .B(n7756), .Z(out[450]) );
  XNOR U4807 ( .A(in[889]), .B(n8596), .Z(n8070) );
  NAND U4808 ( .A(n7911), .B(n7757), .Z(n7758) );
  XNOR U4809 ( .A(n8070), .B(n7758), .Z(out[451]) );
  XNOR U4810 ( .A(in[890]), .B(n8600), .Z(n8078) );
  NAND U4811 ( .A(n7913), .B(n7759), .Z(n7760) );
  XNOR U4812 ( .A(n8078), .B(n7760), .Z(out[452]) );
  XOR U4813 ( .A(in[891]), .B(n8610), .Z(n8082) );
  NAND U4814 ( .A(n7915), .B(n7761), .Z(n7762) );
  XNOR U4815 ( .A(n8082), .B(n7762), .Z(out[453]) );
  XOR U4816 ( .A(in[892]), .B(n8614), .Z(n8086) );
  NAND U4817 ( .A(n7917), .B(n7763), .Z(n7764) );
  XNOR U4818 ( .A(n8086), .B(n7764), .Z(out[454]) );
  XOR U4819 ( .A(in[893]), .B(n8618), .Z(n8090) );
  NAND U4820 ( .A(n7919), .B(n7765), .Z(n7766) );
  XNOR U4821 ( .A(n8090), .B(n7766), .Z(out[455]) );
  XNOR U4822 ( .A(in[894]), .B(n8622), .Z(n8094) );
  NAND U4823 ( .A(n7925), .B(n7767), .Z(n7768) );
  XNOR U4824 ( .A(n8094), .B(n7768), .Z(out[456]) );
  XOR U4825 ( .A(in[895]), .B(n8344), .Z(n8098) );
  NAND U4826 ( .A(n7927), .B(n7769), .Z(n7770) );
  XNOR U4827 ( .A(n8098), .B(n7770), .Z(out[457]) );
  XOR U4828 ( .A(in[832]), .B(n8348), .Z(n8102) );
  NAND U4829 ( .A(n7929), .B(n7771), .Z(n7772) );
  XNOR U4830 ( .A(n8102), .B(n7772), .Z(out[458]) );
  XOR U4831 ( .A(in[833]), .B(n8352), .Z(n8106) );
  NAND U4832 ( .A(n7931), .B(n7773), .Z(n7774) );
  XNOR U4833 ( .A(n8106), .B(n7774), .Z(out[459]) );
  ANDN U4834 ( .B(n7776), .A(n7775), .Z(n7777) );
  XNOR U4835 ( .A(n7778), .B(n7777), .Z(out[45]) );
  XOR U4836 ( .A(in[834]), .B(n8356), .Z(n8110) );
  NAND U4837 ( .A(n7933), .B(n7779), .Z(n7780) );
  XNOR U4838 ( .A(n8110), .B(n7780), .Z(out[460]) );
  XOR U4839 ( .A(in[835]), .B(n8360), .Z(n8114) );
  NAND U4840 ( .A(n7935), .B(n7781), .Z(n7782) );
  XNOR U4841 ( .A(n8114), .B(n7782), .Z(out[461]) );
  XOR U4842 ( .A(in[836]), .B(n8364), .Z(n8122) );
  NAND U4843 ( .A(n7937), .B(n7783), .Z(n7784) );
  XNOR U4844 ( .A(n8122), .B(n7784), .Z(out[462]) );
  XOR U4845 ( .A(in[837]), .B(n8368), .Z(n8126) );
  NAND U4846 ( .A(n7939), .B(n7785), .Z(n7786) );
  XNOR U4847 ( .A(n8126), .B(n7786), .Z(out[463]) );
  XOR U4848 ( .A(in[838]), .B(n8372), .Z(n8130) );
  NAND U4849 ( .A(n7941), .B(n7787), .Z(n7788) );
  XNOR U4850 ( .A(n8130), .B(n7788), .Z(out[464]) );
  XOR U4851 ( .A(in[839]), .B(n8376), .Z(n8134) );
  NAND U4852 ( .A(n7943), .B(n7789), .Z(n7790) );
  XNOR U4853 ( .A(n8134), .B(n7790), .Z(out[465]) );
  XOR U4854 ( .A(in[840]), .B(n8380), .Z(n8138) );
  NAND U4855 ( .A(n7949), .B(n7791), .Z(n7792) );
  XNOR U4856 ( .A(n8138), .B(n7792), .Z(out[466]) );
  XOR U4857 ( .A(in[841]), .B(n8388), .Z(n8142) );
  NAND U4858 ( .A(n7951), .B(n7793), .Z(n7794) );
  XNOR U4859 ( .A(n8142), .B(n7794), .Z(out[467]) );
  XOR U4860 ( .A(in[842]), .B(n8392), .Z(n8146) );
  NAND U4861 ( .A(n7953), .B(n7795), .Z(n7796) );
  XNOR U4862 ( .A(n8146), .B(n7796), .Z(out[468]) );
  XOR U4863 ( .A(in[843]), .B(n8396), .Z(n8150) );
  NAND U4864 ( .A(n7955), .B(n7797), .Z(n7798) );
  XNOR U4865 ( .A(n8150), .B(n7798), .Z(out[469]) );
  ANDN U4866 ( .B(n7800), .A(n7799), .Z(n7801) );
  XNOR U4867 ( .A(n7802), .B(n7801), .Z(out[46]) );
  XOR U4868 ( .A(in[844]), .B(n8400), .Z(n8154) );
  NAND U4869 ( .A(n7957), .B(n7803), .Z(n7804) );
  XNOR U4870 ( .A(n8154), .B(n7804), .Z(out[470]) );
  XOR U4871 ( .A(in[845]), .B(n8404), .Z(n8158) );
  NAND U4872 ( .A(n7959), .B(n7805), .Z(n7806) );
  XNOR U4873 ( .A(n8158), .B(n7806), .Z(out[471]) );
  XOR U4874 ( .A(in[846]), .B(n8408), .Z(n8168) );
  NAND U4875 ( .A(n7961), .B(n7807), .Z(n7808) );
  XNOR U4876 ( .A(n8168), .B(n7808), .Z(out[472]) );
  XOR U4877 ( .A(in[847]), .B(n8412), .Z(n8172) );
  NAND U4878 ( .A(n7963), .B(n7809), .Z(n7810) );
  XNOR U4879 ( .A(n8172), .B(n7810), .Z(out[473]) );
  XOR U4880 ( .A(in[848]), .B(n8416), .Z(n8176) );
  NAND U4881 ( .A(n7965), .B(n7811), .Z(n7812) );
  XNOR U4882 ( .A(n8176), .B(n7812), .Z(out[474]) );
  XOR U4883 ( .A(in[849]), .B(n8420), .Z(n8180) );
  NAND U4884 ( .A(n7967), .B(n7813), .Z(n7814) );
  XNOR U4885 ( .A(n8180), .B(n7814), .Z(out[475]) );
  XOR U4886 ( .A(in[850]), .B(n8424), .Z(n8184) );
  NAND U4887 ( .A(n7973), .B(n7815), .Z(n7816) );
  XNOR U4888 ( .A(n8184), .B(n7816), .Z(out[476]) );
  XNOR U4889 ( .A(in[851]), .B(n8432), .Z(n8188) );
  NAND U4890 ( .A(n7975), .B(n7817), .Z(n7818) );
  XNOR U4891 ( .A(n8188), .B(n7818), .Z(out[477]) );
  XNOR U4892 ( .A(in[852]), .B(n8436), .Z(n8192) );
  NAND U4893 ( .A(n7977), .B(n7819), .Z(n7820) );
  XNOR U4894 ( .A(n8192), .B(n7820), .Z(out[478]) );
  XNOR U4895 ( .A(in[853]), .B(n8440), .Z(n8196) );
  NAND U4896 ( .A(n7979), .B(n7821), .Z(n7822) );
  XNOR U4897 ( .A(n8196), .B(n7822), .Z(out[479]) );
  ANDN U4898 ( .B(n7824), .A(n7823), .Z(n7825) );
  XNOR U4899 ( .A(n7826), .B(n7825), .Z(out[47]) );
  XNOR U4900 ( .A(in[854]), .B(n8444), .Z(n8200) );
  NAND U4901 ( .A(n7981), .B(n7827), .Z(n7828) );
  XNOR U4902 ( .A(n8200), .B(n7828), .Z(out[480]) );
  XNOR U4903 ( .A(in[855]), .B(n8448), .Z(n8204) );
  NAND U4904 ( .A(n7983), .B(n7829), .Z(n7830) );
  XNOR U4905 ( .A(n8204), .B(n7830), .Z(out[481]) );
  XNOR U4906 ( .A(in[856]), .B(n8452), .Z(n8212) );
  NAND U4907 ( .A(n7985), .B(n7831), .Z(n7832) );
  XNOR U4908 ( .A(n8212), .B(n7832), .Z(out[482]) );
  XNOR U4909 ( .A(in[857]), .B(n8456), .Z(n8216) );
  NAND U4910 ( .A(n7987), .B(n7833), .Z(n7834) );
  XNOR U4911 ( .A(n8216), .B(n7834), .Z(out[483]) );
  XNOR U4912 ( .A(in[858]), .B(n8460), .Z(n8220) );
  NAND U4913 ( .A(n7989), .B(n7835), .Z(n7836) );
  XNOR U4914 ( .A(n8220), .B(n7836), .Z(out[484]) );
  XNOR U4915 ( .A(in[859]), .B(n8464), .Z(n8224) );
  NAND U4916 ( .A(n7991), .B(n7837), .Z(n7838) );
  XNOR U4917 ( .A(n8224), .B(n7838), .Z(out[485]) );
  XNOR U4918 ( .A(in[860]), .B(n8468), .Z(n8228) );
  NAND U4919 ( .A(n7997), .B(n7839), .Z(n7840) );
  XNOR U4920 ( .A(n8228), .B(n7840), .Z(out[486]) );
  XNOR U4921 ( .A(in[861]), .B(n8476), .Z(n8232) );
  NAND U4922 ( .A(n7999), .B(n7841), .Z(n7842) );
  XNOR U4923 ( .A(n8232), .B(n7842), .Z(out[487]) );
  XNOR U4924 ( .A(in[862]), .B(n8480), .Z(n8236) );
  NAND U4925 ( .A(n8001), .B(n7843), .Z(n7844) );
  XNOR U4926 ( .A(n8236), .B(n7844), .Z(out[488]) );
  XNOR U4927 ( .A(in[863]), .B(n8484), .Z(n8240) );
  NAND U4928 ( .A(n8003), .B(n7845), .Z(n7846) );
  XNOR U4929 ( .A(n8240), .B(n7846), .Z(out[489]) );
  ANDN U4930 ( .B(n7848), .A(n7847), .Z(n7849) );
  XNOR U4931 ( .A(n7850), .B(n7849), .Z(out[48]) );
  XNOR U4932 ( .A(in[864]), .B(n8488), .Z(n8244) );
  NAND U4933 ( .A(n8005), .B(n7851), .Z(n7852) );
  XNOR U4934 ( .A(n8244), .B(n7852), .Z(out[490]) );
  XNOR U4935 ( .A(in[865]), .B(n8492), .Z(n8248) );
  NAND U4936 ( .A(n8007), .B(n7853), .Z(n7854) );
  XNOR U4937 ( .A(n8248), .B(n7854), .Z(out[491]) );
  XOR U4938 ( .A(n8496), .B(in[866]), .Z(n8256) );
  NAND U4939 ( .A(n8009), .B(n7855), .Z(n7856) );
  XNOR U4940 ( .A(n8256), .B(n7856), .Z(out[492]) );
  XOR U4941 ( .A(n8500), .B(in[867]), .Z(n8260) );
  NAND U4942 ( .A(n8011), .B(n7857), .Z(n7858) );
  XNOR U4943 ( .A(n8260), .B(n7858), .Z(out[493]) );
  XOR U4944 ( .A(n8504), .B(in[868]), .Z(n8264) );
  NAND U4945 ( .A(n8013), .B(n7859), .Z(n7860) );
  XNOR U4946 ( .A(n8264), .B(n7860), .Z(out[494]) );
  XOR U4947 ( .A(n8508), .B(in[869]), .Z(n8268) );
  NAND U4948 ( .A(n8015), .B(n7861), .Z(n7862) );
  XNOR U4949 ( .A(n8268), .B(n7862), .Z(out[495]) );
  XNOR U4950 ( .A(in[870]), .B(n8512), .Z(n8272) );
  NAND U4951 ( .A(n8021), .B(n7863), .Z(n7864) );
  XNOR U4952 ( .A(n8272), .B(n7864), .Z(out[496]) );
  XNOR U4953 ( .A(in[871]), .B(n8520), .Z(n8276) );
  NAND U4954 ( .A(n8023), .B(n7865), .Z(n7866) );
  XNOR U4955 ( .A(n8276), .B(n7866), .Z(out[497]) );
  XNOR U4956 ( .A(in[872]), .B(n8524), .Z(n8280) );
  NAND U4957 ( .A(n8025), .B(n7867), .Z(n7868) );
  XNOR U4958 ( .A(n8280), .B(n7868), .Z(out[498]) );
  XNOR U4959 ( .A(in[873]), .B(n8528), .Z(n8284) );
  NAND U4960 ( .A(n8027), .B(n7869), .Z(n7870) );
  XNOR U4961 ( .A(n8284), .B(n7870), .Z(out[499]) );
  ANDN U4962 ( .B(n7872), .A(n7871), .Z(n7873) );
  XNOR U4963 ( .A(n7874), .B(n7873), .Z(out[49]) );
  OR U4964 ( .A(n8560), .B(n7875), .Z(n7876) );
  XNOR U4965 ( .A(n8559), .B(n7876), .Z(out[4]) );
  XNOR U4966 ( .A(in[874]), .B(n8532), .Z(n8288) );
  NAND U4967 ( .A(n8029), .B(n7877), .Z(n7878) );
  XNOR U4968 ( .A(n8288), .B(n7878), .Z(out[500]) );
  XNOR U4969 ( .A(in[875]), .B(n8536), .Z(n8292) );
  NAND U4970 ( .A(n8031), .B(n7879), .Z(n7880) );
  XNOR U4971 ( .A(n8292), .B(n7880), .Z(out[501]) );
  XNOR U4972 ( .A(in[876]), .B(n8540), .Z(n8300) );
  NAND U4973 ( .A(n8033), .B(n7881), .Z(n7882) );
  XNOR U4974 ( .A(n8300), .B(n7882), .Z(out[502]) );
  XNOR U4975 ( .A(in[877]), .B(n8544), .Z(n8304) );
  NAND U4976 ( .A(n8035), .B(n7883), .Z(n7884) );
  XNOR U4977 ( .A(n8304), .B(n7884), .Z(out[503]) );
  XNOR U4978 ( .A(in[878]), .B(n8548), .Z(n8308) );
  NAND U4979 ( .A(n8037), .B(n7885), .Z(n7886) );
  XNOR U4980 ( .A(n8308), .B(n7886), .Z(out[504]) );
  XNOR U4981 ( .A(in[879]), .B(n8552), .Z(n8312) );
  NAND U4982 ( .A(n8039), .B(n7887), .Z(n7888) );
  XNOR U4983 ( .A(n8312), .B(n7888), .Z(out[505]) );
  XNOR U4984 ( .A(in[880]), .B(n8556), .Z(n8316) );
  NAND U4985 ( .A(n8045), .B(n7889), .Z(n7890) );
  XNOR U4986 ( .A(n8316), .B(n7890), .Z(out[506]) );
  XNOR U4987 ( .A(in[881]), .B(n8564), .Z(n8320) );
  NAND U4988 ( .A(n8047), .B(n7891), .Z(n7892) );
  XNOR U4989 ( .A(n8320), .B(n7892), .Z(out[507]) );
  XNOR U4990 ( .A(in[882]), .B(n8568), .Z(n8324) );
  NAND U4991 ( .A(n8049), .B(n7893), .Z(n7894) );
  XNOR U4992 ( .A(n8324), .B(n7894), .Z(out[508]) );
  XNOR U4993 ( .A(in[883]), .B(n8572), .Z(n8328) );
  NAND U4994 ( .A(n8051), .B(n7895), .Z(n7896) );
  XNOR U4995 ( .A(n8328), .B(n7896), .Z(out[509]) );
  ANDN U4996 ( .B(n7898), .A(n7897), .Z(n7899) );
  XNOR U4997 ( .A(n7900), .B(n7899), .Z(out[50]) );
  XNOR U4998 ( .A(in[884]), .B(n8576), .Z(n8332) );
  NAND U4999 ( .A(n8053), .B(n7901), .Z(n7902) );
  XNOR U5000 ( .A(n8332), .B(n7902), .Z(out[510]) );
  XNOR U5001 ( .A(in[885]), .B(n8580), .Z(n8336) );
  NAND U5002 ( .A(n8055), .B(n7903), .Z(n7904) );
  XNOR U5003 ( .A(n8336), .B(n7904), .Z(out[511]) );
  OR U5004 ( .A(n8058), .B(n7905), .Z(n7906) );
  XNOR U5005 ( .A(n8057), .B(n7906), .Z(out[512]) );
  OR U5006 ( .A(n8062), .B(n7907), .Z(n7908) );
  XNOR U5007 ( .A(n8061), .B(n7908), .Z(out[513]) );
  OR U5008 ( .A(n8066), .B(n7909), .Z(n7910) );
  XNOR U5009 ( .A(n8065), .B(n7910), .Z(out[514]) );
  OR U5010 ( .A(n8070), .B(n7911), .Z(n7912) );
  XNOR U5011 ( .A(n8069), .B(n7912), .Z(out[515]) );
  OR U5012 ( .A(n8078), .B(n7913), .Z(n7914) );
  XNOR U5013 ( .A(n8077), .B(n7914), .Z(out[516]) );
  OR U5014 ( .A(n8082), .B(n7915), .Z(n7916) );
  XNOR U5015 ( .A(n8081), .B(n7916), .Z(out[517]) );
  OR U5016 ( .A(n8086), .B(n7917), .Z(n7918) );
  XNOR U5017 ( .A(n8085), .B(n7918), .Z(out[518]) );
  OR U5018 ( .A(n8090), .B(n7919), .Z(n7920) );
  XNOR U5019 ( .A(n8089), .B(n7920), .Z(out[519]) );
  ANDN U5020 ( .B(n7922), .A(n7921), .Z(n7923) );
  XNOR U5021 ( .A(n7924), .B(n7923), .Z(out[51]) );
  OR U5022 ( .A(n8094), .B(n7925), .Z(n7926) );
  XNOR U5023 ( .A(n8093), .B(n7926), .Z(out[520]) );
  OR U5024 ( .A(n8098), .B(n7927), .Z(n7928) );
  XNOR U5025 ( .A(n8097), .B(n7928), .Z(out[521]) );
  OR U5026 ( .A(n8102), .B(n7929), .Z(n7930) );
  XNOR U5027 ( .A(n8101), .B(n7930), .Z(out[522]) );
  OR U5028 ( .A(n8106), .B(n7931), .Z(n7932) );
  XNOR U5029 ( .A(n8105), .B(n7932), .Z(out[523]) );
  OR U5030 ( .A(n8110), .B(n7933), .Z(n7934) );
  XNOR U5031 ( .A(n8109), .B(n7934), .Z(out[524]) );
  OR U5032 ( .A(n8114), .B(n7935), .Z(n7936) );
  XNOR U5033 ( .A(n8113), .B(n7936), .Z(out[525]) );
  OR U5034 ( .A(n8122), .B(n7937), .Z(n7938) );
  XNOR U5035 ( .A(n8121), .B(n7938), .Z(out[526]) );
  OR U5036 ( .A(n8126), .B(n7939), .Z(n7940) );
  XNOR U5037 ( .A(n8125), .B(n7940), .Z(out[527]) );
  OR U5038 ( .A(n8130), .B(n7941), .Z(n7942) );
  XNOR U5039 ( .A(n8129), .B(n7942), .Z(out[528]) );
  OR U5040 ( .A(n8134), .B(n7943), .Z(n7944) );
  XNOR U5041 ( .A(n8133), .B(n7944), .Z(out[529]) );
  ANDN U5042 ( .B(n7946), .A(n7945), .Z(n7947) );
  XNOR U5043 ( .A(n7948), .B(n7947), .Z(out[52]) );
  OR U5044 ( .A(n8138), .B(n7949), .Z(n7950) );
  XNOR U5045 ( .A(n8137), .B(n7950), .Z(out[530]) );
  OR U5046 ( .A(n8142), .B(n7951), .Z(n7952) );
  XNOR U5047 ( .A(n8141), .B(n7952), .Z(out[531]) );
  OR U5048 ( .A(n8146), .B(n7953), .Z(n7954) );
  XNOR U5049 ( .A(n8145), .B(n7954), .Z(out[532]) );
  OR U5050 ( .A(n8150), .B(n7955), .Z(n7956) );
  XNOR U5051 ( .A(n8149), .B(n7956), .Z(out[533]) );
  OR U5052 ( .A(n8154), .B(n7957), .Z(n7958) );
  XNOR U5053 ( .A(n8153), .B(n7958), .Z(out[534]) );
  OR U5054 ( .A(n8158), .B(n7959), .Z(n7960) );
  XNOR U5055 ( .A(n8157), .B(n7960), .Z(out[535]) );
  OR U5056 ( .A(n8168), .B(n7961), .Z(n7962) );
  XNOR U5057 ( .A(n8167), .B(n7962), .Z(out[536]) );
  OR U5058 ( .A(n8172), .B(n7963), .Z(n7964) );
  XNOR U5059 ( .A(n8171), .B(n7964), .Z(out[537]) );
  OR U5060 ( .A(n8176), .B(n7965), .Z(n7966) );
  XNOR U5061 ( .A(n8175), .B(n7966), .Z(out[538]) );
  OR U5062 ( .A(n8180), .B(n7967), .Z(n7968) );
  XNOR U5063 ( .A(n8179), .B(n7968), .Z(out[539]) );
  ANDN U5064 ( .B(n7970), .A(n7969), .Z(n7971) );
  XNOR U5065 ( .A(n7972), .B(n7971), .Z(out[53]) );
  OR U5066 ( .A(n8184), .B(n7973), .Z(n7974) );
  XNOR U5067 ( .A(n8183), .B(n7974), .Z(out[540]) );
  OR U5068 ( .A(n8188), .B(n7975), .Z(n7976) );
  XNOR U5069 ( .A(n8187), .B(n7976), .Z(out[541]) );
  OR U5070 ( .A(n8192), .B(n7977), .Z(n7978) );
  XNOR U5071 ( .A(n8191), .B(n7978), .Z(out[542]) );
  OR U5072 ( .A(n8196), .B(n7979), .Z(n7980) );
  XNOR U5073 ( .A(n8195), .B(n7980), .Z(out[543]) );
  OR U5074 ( .A(n8200), .B(n7981), .Z(n7982) );
  XNOR U5075 ( .A(n8199), .B(n7982), .Z(out[544]) );
  OR U5076 ( .A(n8204), .B(n7983), .Z(n7984) );
  XNOR U5077 ( .A(n8203), .B(n7984), .Z(out[545]) );
  OR U5078 ( .A(n8212), .B(n7985), .Z(n7986) );
  XNOR U5079 ( .A(n8211), .B(n7986), .Z(out[546]) );
  OR U5080 ( .A(n8216), .B(n7987), .Z(n7988) );
  XNOR U5081 ( .A(n8215), .B(n7988), .Z(out[547]) );
  OR U5082 ( .A(n8220), .B(n7989), .Z(n7990) );
  XNOR U5083 ( .A(n8219), .B(n7990), .Z(out[548]) );
  OR U5084 ( .A(n8224), .B(n7991), .Z(n7992) );
  XNOR U5085 ( .A(n8223), .B(n7992), .Z(out[549]) );
  ANDN U5086 ( .B(n7994), .A(n7993), .Z(n7995) );
  XNOR U5087 ( .A(n7996), .B(n7995), .Z(out[54]) );
  OR U5088 ( .A(n8228), .B(n7997), .Z(n7998) );
  XNOR U5089 ( .A(n8227), .B(n7998), .Z(out[550]) );
  OR U5090 ( .A(n8232), .B(n7999), .Z(n8000) );
  XNOR U5091 ( .A(n8231), .B(n8000), .Z(out[551]) );
  OR U5092 ( .A(n8236), .B(n8001), .Z(n8002) );
  XNOR U5093 ( .A(n8235), .B(n8002), .Z(out[552]) );
  OR U5094 ( .A(n8240), .B(n8003), .Z(n8004) );
  XNOR U5095 ( .A(n8239), .B(n8004), .Z(out[553]) );
  OR U5096 ( .A(n8244), .B(n8005), .Z(n8006) );
  XNOR U5097 ( .A(n8243), .B(n8006), .Z(out[554]) );
  OR U5098 ( .A(n8248), .B(n8007), .Z(n8008) );
  XNOR U5099 ( .A(n8247), .B(n8008), .Z(out[555]) );
  OR U5100 ( .A(n8256), .B(n8009), .Z(n8010) );
  XNOR U5101 ( .A(n8255), .B(n8010), .Z(out[556]) );
  OR U5102 ( .A(n8260), .B(n8011), .Z(n8012) );
  XNOR U5103 ( .A(n8259), .B(n8012), .Z(out[557]) );
  OR U5104 ( .A(n8264), .B(n8013), .Z(n8014) );
  XNOR U5105 ( .A(n8263), .B(n8014), .Z(out[558]) );
  OR U5106 ( .A(n8268), .B(n8015), .Z(n8016) );
  XNOR U5107 ( .A(n8267), .B(n8016), .Z(out[559]) );
  ANDN U5108 ( .B(n8018), .A(n8017), .Z(n8019) );
  XNOR U5109 ( .A(n8020), .B(n8019), .Z(out[55]) );
  OR U5110 ( .A(n8272), .B(n8021), .Z(n8022) );
  XNOR U5111 ( .A(n8271), .B(n8022), .Z(out[560]) );
  OR U5112 ( .A(n8276), .B(n8023), .Z(n8024) );
  XNOR U5113 ( .A(n8275), .B(n8024), .Z(out[561]) );
  OR U5114 ( .A(n8280), .B(n8025), .Z(n8026) );
  XNOR U5115 ( .A(n8279), .B(n8026), .Z(out[562]) );
  OR U5116 ( .A(n8284), .B(n8027), .Z(n8028) );
  XNOR U5117 ( .A(n8283), .B(n8028), .Z(out[563]) );
  OR U5118 ( .A(n8288), .B(n8029), .Z(n8030) );
  XNOR U5119 ( .A(n8287), .B(n8030), .Z(out[564]) );
  OR U5120 ( .A(n8292), .B(n8031), .Z(n8032) );
  XNOR U5121 ( .A(n8291), .B(n8032), .Z(out[565]) );
  OR U5122 ( .A(n8300), .B(n8033), .Z(n8034) );
  XNOR U5123 ( .A(n8299), .B(n8034), .Z(out[566]) );
  OR U5124 ( .A(n8304), .B(n8035), .Z(n8036) );
  XNOR U5125 ( .A(n8303), .B(n8036), .Z(out[567]) );
  OR U5126 ( .A(n8308), .B(n8037), .Z(n8038) );
  XNOR U5127 ( .A(n8307), .B(n8038), .Z(out[568]) );
  OR U5128 ( .A(n8312), .B(n8039), .Z(n8040) );
  XNOR U5129 ( .A(n8311), .B(n8040), .Z(out[569]) );
  ANDN U5130 ( .B(n8042), .A(n8041), .Z(n8043) );
  XNOR U5131 ( .A(n8044), .B(n8043), .Z(out[56]) );
  OR U5132 ( .A(n8316), .B(n8045), .Z(n8046) );
  XNOR U5133 ( .A(n8315), .B(n8046), .Z(out[570]) );
  OR U5134 ( .A(n8320), .B(n8047), .Z(n8048) );
  XNOR U5135 ( .A(n8319), .B(n8048), .Z(out[571]) );
  OR U5136 ( .A(n8324), .B(n8049), .Z(n8050) );
  XNOR U5137 ( .A(n8323), .B(n8050), .Z(out[572]) );
  OR U5138 ( .A(n8328), .B(n8051), .Z(n8052) );
  XNOR U5139 ( .A(n8327), .B(n8052), .Z(out[573]) );
  OR U5140 ( .A(n8332), .B(n8053), .Z(n8054) );
  XNOR U5141 ( .A(n8331), .B(n8054), .Z(out[574]) );
  OR U5142 ( .A(n8336), .B(n8055), .Z(n8056) );
  XNOR U5143 ( .A(n8335), .B(n8056), .Z(out[575]) );
  ANDN U5144 ( .B(n8058), .A(n8057), .Z(n8059) );
  XNOR U5145 ( .A(n8060), .B(n8059), .Z(out[576]) );
  ANDN U5146 ( .B(n8062), .A(n8061), .Z(n8063) );
  XNOR U5147 ( .A(n8064), .B(n8063), .Z(out[577]) );
  ANDN U5148 ( .B(n8066), .A(n8065), .Z(n8067) );
  XNOR U5149 ( .A(n8068), .B(n8067), .Z(out[578]) );
  ANDN U5150 ( .B(n8070), .A(n8069), .Z(n8071) );
  XNOR U5151 ( .A(n8072), .B(n8071), .Z(out[579]) );
  ANDN U5152 ( .B(n8074), .A(n8073), .Z(n8075) );
  XNOR U5153 ( .A(n8076), .B(n8075), .Z(out[57]) );
  ANDN U5154 ( .B(n8078), .A(n8077), .Z(n8079) );
  XNOR U5155 ( .A(n8080), .B(n8079), .Z(out[580]) );
  ANDN U5156 ( .B(n8082), .A(n8081), .Z(n8083) );
  XNOR U5157 ( .A(n8084), .B(n8083), .Z(out[581]) );
  ANDN U5158 ( .B(n8086), .A(n8085), .Z(n8087) );
  XNOR U5159 ( .A(n8088), .B(n8087), .Z(out[582]) );
  ANDN U5160 ( .B(n8090), .A(n8089), .Z(n8091) );
  XNOR U5161 ( .A(n8092), .B(n8091), .Z(out[583]) );
  ANDN U5162 ( .B(n8094), .A(n8093), .Z(n8095) );
  XNOR U5163 ( .A(n8096), .B(n8095), .Z(out[584]) );
  ANDN U5164 ( .B(n8098), .A(n8097), .Z(n8099) );
  XNOR U5165 ( .A(n8100), .B(n8099), .Z(out[585]) );
  ANDN U5166 ( .B(n8102), .A(n8101), .Z(n8103) );
  XNOR U5167 ( .A(n8104), .B(n8103), .Z(out[586]) );
  ANDN U5168 ( .B(n8106), .A(n8105), .Z(n8107) );
  XNOR U5169 ( .A(n8108), .B(n8107), .Z(out[587]) );
  ANDN U5170 ( .B(n8110), .A(n8109), .Z(n8111) );
  XNOR U5171 ( .A(n8112), .B(n8111), .Z(out[588]) );
  ANDN U5172 ( .B(n8114), .A(n8113), .Z(n8115) );
  XNOR U5173 ( .A(n8116), .B(n8115), .Z(out[589]) );
  ANDN U5174 ( .B(n8118), .A(n8117), .Z(n8119) );
  XNOR U5175 ( .A(n8120), .B(n8119), .Z(out[58]) );
  ANDN U5176 ( .B(n8122), .A(n8121), .Z(n8123) );
  XNOR U5177 ( .A(n8124), .B(n8123), .Z(out[590]) );
  ANDN U5178 ( .B(n8126), .A(n8125), .Z(n8127) );
  XNOR U5179 ( .A(n8128), .B(n8127), .Z(out[591]) );
  ANDN U5180 ( .B(n8130), .A(n8129), .Z(n8131) );
  XNOR U5181 ( .A(n8132), .B(n8131), .Z(out[592]) );
  ANDN U5182 ( .B(n8134), .A(n8133), .Z(n8135) );
  XNOR U5183 ( .A(n8136), .B(n8135), .Z(out[593]) );
  ANDN U5184 ( .B(n8138), .A(n8137), .Z(n8139) );
  XNOR U5185 ( .A(n8140), .B(n8139), .Z(out[594]) );
  ANDN U5186 ( .B(n8142), .A(n8141), .Z(n8143) );
  XNOR U5187 ( .A(n8144), .B(n8143), .Z(out[595]) );
  ANDN U5188 ( .B(n8146), .A(n8145), .Z(n8147) );
  XNOR U5189 ( .A(n8148), .B(n8147), .Z(out[596]) );
  ANDN U5190 ( .B(n8150), .A(n8149), .Z(n8151) );
  XNOR U5191 ( .A(n8152), .B(n8151), .Z(out[597]) );
  ANDN U5192 ( .B(n8154), .A(n8153), .Z(n8155) );
  XNOR U5193 ( .A(n8156), .B(n8155), .Z(out[598]) );
  ANDN U5194 ( .B(n8158), .A(n8157), .Z(n8159) );
  XNOR U5195 ( .A(n8160), .B(n8159), .Z(out[599]) );
  ANDN U5196 ( .B(n8162), .A(n8161), .Z(n8163) );
  XNOR U5197 ( .A(n8164), .B(n8163), .Z(out[59]) );
  OR U5198 ( .A(n8604), .B(n8165), .Z(n8166) );
  XNOR U5199 ( .A(n8603), .B(n8166), .Z(out[5]) );
  ANDN U5200 ( .B(n8168), .A(n8167), .Z(n8169) );
  XNOR U5201 ( .A(n8170), .B(n8169), .Z(out[600]) );
  ANDN U5202 ( .B(n8172), .A(n8171), .Z(n8173) );
  XNOR U5203 ( .A(n8174), .B(n8173), .Z(out[601]) );
  ANDN U5204 ( .B(n8176), .A(n8175), .Z(n8177) );
  XNOR U5205 ( .A(n8178), .B(n8177), .Z(out[602]) );
  ANDN U5206 ( .B(n8180), .A(n8179), .Z(n8181) );
  XNOR U5207 ( .A(n8182), .B(n8181), .Z(out[603]) );
  ANDN U5208 ( .B(n8184), .A(n8183), .Z(n8185) );
  XNOR U5209 ( .A(n8186), .B(n8185), .Z(out[604]) );
  ANDN U5210 ( .B(n8188), .A(n8187), .Z(n8189) );
  XNOR U5211 ( .A(n8190), .B(n8189), .Z(out[605]) );
  ANDN U5212 ( .B(n8192), .A(n8191), .Z(n8193) );
  XNOR U5213 ( .A(n8194), .B(n8193), .Z(out[606]) );
  ANDN U5214 ( .B(n8196), .A(n8195), .Z(n8197) );
  XNOR U5215 ( .A(n8198), .B(n8197), .Z(out[607]) );
  ANDN U5216 ( .B(n8200), .A(n8199), .Z(n8201) );
  XNOR U5217 ( .A(n8202), .B(n8201), .Z(out[608]) );
  ANDN U5218 ( .B(n8204), .A(n8203), .Z(n8205) );
  XNOR U5219 ( .A(n8206), .B(n8205), .Z(out[609]) );
  ANDN U5220 ( .B(n8208), .A(n8207), .Z(n8209) );
  XNOR U5221 ( .A(n8210), .B(n8209), .Z(out[60]) );
  ANDN U5222 ( .B(n8212), .A(n8211), .Z(n8213) );
  XNOR U5223 ( .A(n8214), .B(n8213), .Z(out[610]) );
  ANDN U5224 ( .B(n8216), .A(n8215), .Z(n8217) );
  XNOR U5225 ( .A(n8218), .B(n8217), .Z(out[611]) );
  ANDN U5226 ( .B(n8220), .A(n8219), .Z(n8221) );
  XNOR U5227 ( .A(n8222), .B(n8221), .Z(out[612]) );
  ANDN U5228 ( .B(n8224), .A(n8223), .Z(n8225) );
  XNOR U5229 ( .A(n8226), .B(n8225), .Z(out[613]) );
  ANDN U5230 ( .B(n8228), .A(n8227), .Z(n8229) );
  XNOR U5231 ( .A(n8230), .B(n8229), .Z(out[614]) );
  ANDN U5232 ( .B(n8232), .A(n8231), .Z(n8233) );
  XNOR U5233 ( .A(n8234), .B(n8233), .Z(out[615]) );
  ANDN U5234 ( .B(n8236), .A(n8235), .Z(n8237) );
  XNOR U5235 ( .A(n8238), .B(n8237), .Z(out[616]) );
  ANDN U5236 ( .B(n8240), .A(n8239), .Z(n8241) );
  XNOR U5237 ( .A(n8242), .B(n8241), .Z(out[617]) );
  ANDN U5238 ( .B(n8244), .A(n8243), .Z(n8245) );
  XNOR U5239 ( .A(n8246), .B(n8245), .Z(out[618]) );
  ANDN U5240 ( .B(n8248), .A(n8247), .Z(n8249) );
  XNOR U5241 ( .A(n8250), .B(n8249), .Z(out[619]) );
  ANDN U5242 ( .B(n8252), .A(n8251), .Z(n8253) );
  XNOR U5243 ( .A(n8254), .B(n8253), .Z(out[61]) );
  ANDN U5244 ( .B(n8256), .A(n8255), .Z(n8257) );
  XNOR U5245 ( .A(n8258), .B(n8257), .Z(out[620]) );
  ANDN U5246 ( .B(n8260), .A(n8259), .Z(n8261) );
  XNOR U5247 ( .A(n8262), .B(n8261), .Z(out[621]) );
  ANDN U5248 ( .B(n8264), .A(n8263), .Z(n8265) );
  XNOR U5249 ( .A(n8266), .B(n8265), .Z(out[622]) );
  ANDN U5250 ( .B(n8268), .A(n8267), .Z(n8269) );
  XNOR U5251 ( .A(n8270), .B(n8269), .Z(out[623]) );
  ANDN U5252 ( .B(n8272), .A(n8271), .Z(n8273) );
  XNOR U5253 ( .A(n8274), .B(n8273), .Z(out[624]) );
  ANDN U5254 ( .B(n8276), .A(n8275), .Z(n8277) );
  XNOR U5255 ( .A(n8278), .B(n8277), .Z(out[625]) );
  ANDN U5256 ( .B(n8280), .A(n8279), .Z(n8281) );
  XNOR U5257 ( .A(n8282), .B(n8281), .Z(out[626]) );
  ANDN U5258 ( .B(n8284), .A(n8283), .Z(n8285) );
  XNOR U5259 ( .A(n8286), .B(n8285), .Z(out[627]) );
  ANDN U5260 ( .B(n8288), .A(n8287), .Z(n8289) );
  XNOR U5261 ( .A(n8290), .B(n8289), .Z(out[628]) );
  ANDN U5262 ( .B(n8292), .A(n8291), .Z(n8293) );
  XNOR U5263 ( .A(n8294), .B(n8293), .Z(out[629]) );
  ANDN U5264 ( .B(n8296), .A(n8295), .Z(n8297) );
  XNOR U5265 ( .A(n8298), .B(n8297), .Z(out[62]) );
  ANDN U5266 ( .B(n8300), .A(n8299), .Z(n8301) );
  XNOR U5267 ( .A(n8302), .B(n8301), .Z(out[630]) );
  ANDN U5268 ( .B(n8304), .A(n8303), .Z(n8305) );
  XNOR U5269 ( .A(n8306), .B(n8305), .Z(out[631]) );
  ANDN U5270 ( .B(n8308), .A(n8307), .Z(n8309) );
  XNOR U5271 ( .A(n8310), .B(n8309), .Z(out[632]) );
  ANDN U5272 ( .B(n8312), .A(n8311), .Z(n8313) );
  XNOR U5273 ( .A(n8314), .B(n8313), .Z(out[633]) );
  ANDN U5274 ( .B(n8316), .A(n8315), .Z(n8317) );
  XNOR U5275 ( .A(n8318), .B(n8317), .Z(out[634]) );
  ANDN U5276 ( .B(n8320), .A(n8319), .Z(n8321) );
  XNOR U5277 ( .A(n8322), .B(n8321), .Z(out[635]) );
  ANDN U5278 ( .B(n8324), .A(n8323), .Z(n8325) );
  XNOR U5279 ( .A(n8326), .B(n8325), .Z(out[636]) );
  ANDN U5280 ( .B(n8328), .A(n8327), .Z(n8329) );
  XNOR U5281 ( .A(n8330), .B(n8329), .Z(out[637]) );
  ANDN U5282 ( .B(n8332), .A(n8331), .Z(n8333) );
  XNOR U5283 ( .A(n8334), .B(n8333), .Z(out[638]) );
  ANDN U5284 ( .B(n8336), .A(n8335), .Z(n8337) );
  XNOR U5285 ( .A(n8338), .B(n8337), .Z(out[639]) );
  ANDN U5286 ( .B(n8340), .A(n8339), .Z(n8341) );
  XNOR U5287 ( .A(n8342), .B(n8341), .Z(out[63]) );
  XNOR U5288 ( .A(in[302]), .B(n8343), .Z(n8772) );
  XNOR U5289 ( .A(in[1535]), .B(n8344), .Z(n9150) );
  XNOR U5290 ( .A(in[1146]), .B(n8345), .Z(n9147) );
  NAND U5291 ( .A(n9150), .B(n9147), .Z(n8346) );
  XNOR U5292 ( .A(n8772), .B(n8346), .Z(out[640]) );
  XNOR U5293 ( .A(in[303]), .B(n8347), .Z(n8775) );
  XNOR U5294 ( .A(in[1472]), .B(n8348), .Z(n9154) );
  XNOR U5295 ( .A(in[1147]), .B(n8349), .Z(n9151) );
  NAND U5296 ( .A(n9154), .B(n9151), .Z(n8350) );
  XNOR U5297 ( .A(n8775), .B(n8350), .Z(out[641]) );
  XNOR U5298 ( .A(in[304]), .B(n8351), .Z(n8782) );
  XNOR U5299 ( .A(in[1473]), .B(n8352), .Z(n9158) );
  XNOR U5300 ( .A(in[1148]), .B(n8353), .Z(n9155) );
  NAND U5301 ( .A(n9158), .B(n9155), .Z(n8354) );
  XNOR U5302 ( .A(n8782), .B(n8354), .Z(out[642]) );
  XNOR U5303 ( .A(in[305]), .B(n8355), .Z(n8785) );
  XNOR U5304 ( .A(in[1474]), .B(n8356), .Z(n9162) );
  XNOR U5305 ( .A(in[1149]), .B(n8357), .Z(n9159) );
  NAND U5306 ( .A(n9162), .B(n9159), .Z(n8358) );
  XNOR U5307 ( .A(n8785), .B(n8358), .Z(out[643]) );
  XNOR U5308 ( .A(in[306]), .B(n8359), .Z(n8788) );
  XNOR U5309 ( .A(in[1475]), .B(n8360), .Z(n9174) );
  XNOR U5310 ( .A(in[1150]), .B(n8361), .Z(n9171) );
  NAND U5311 ( .A(n9174), .B(n9171), .Z(n8362) );
  XNOR U5312 ( .A(n8788), .B(n8362), .Z(out[644]) );
  XNOR U5313 ( .A(in[307]), .B(n8363), .Z(n8791) );
  XNOR U5314 ( .A(in[1476]), .B(n8364), .Z(n9178) );
  XNOR U5315 ( .A(in[1151]), .B(n8365), .Z(n9175) );
  NAND U5316 ( .A(n9178), .B(n9175), .Z(n8366) );
  XNOR U5317 ( .A(n8791), .B(n8366), .Z(out[645]) );
  XNOR U5318 ( .A(in[308]), .B(n8367), .Z(n8794) );
  XNOR U5319 ( .A(in[1477]), .B(n8368), .Z(n9182) );
  XNOR U5320 ( .A(in[1088]), .B(n8369), .Z(n9179) );
  NAND U5321 ( .A(n9182), .B(n9179), .Z(n8370) );
  XNOR U5322 ( .A(n8794), .B(n8370), .Z(out[646]) );
  XNOR U5323 ( .A(in[309]), .B(n8371), .Z(n8797) );
  XNOR U5324 ( .A(in[1478]), .B(n8372), .Z(n9186) );
  XNOR U5325 ( .A(in[1089]), .B(n8373), .Z(n9183) );
  NAND U5326 ( .A(n9186), .B(n9183), .Z(n8374) );
  XNOR U5327 ( .A(n8797), .B(n8374), .Z(out[647]) );
  XNOR U5328 ( .A(in[310]), .B(n8375), .Z(n8800) );
  XNOR U5329 ( .A(in[1479]), .B(n8376), .Z(n9190) );
  XOR U5330 ( .A(n8377), .B(in[1090]), .Z(n9187) );
  NAND U5331 ( .A(n9190), .B(n9187), .Z(n8378) );
  XNOR U5332 ( .A(n8800), .B(n8378), .Z(out[648]) );
  XNOR U5333 ( .A(in[311]), .B(n8379), .Z(n8803) );
  XNOR U5334 ( .A(in[1480]), .B(n8380), .Z(n9194) );
  XOR U5335 ( .A(n8381), .B(in[1091]), .Z(n9191) );
  NAND U5336 ( .A(n9194), .B(n9191), .Z(n8382) );
  XNOR U5337 ( .A(n8803), .B(n8382), .Z(out[649]) );
  NOR U5338 ( .A(n8384), .B(n8383), .Z(n8385) );
  XNOR U5339 ( .A(n8386), .B(n8385), .Z(out[64]) );
  XNOR U5340 ( .A(in[312]), .B(n8387), .Z(n8806) );
  XNOR U5341 ( .A(in[1481]), .B(n8388), .Z(n9198) );
  XOR U5342 ( .A(n8389), .B(in[1092]), .Z(n9195) );
  NAND U5343 ( .A(n9198), .B(n9195), .Z(n8390) );
  XNOR U5344 ( .A(n8806), .B(n8390), .Z(out[650]) );
  XNOR U5345 ( .A(in[313]), .B(n8391), .Z(n8809) );
  XNOR U5346 ( .A(in[1482]), .B(n8392), .Z(n9202) );
  XOR U5347 ( .A(n8393), .B(in[1093]), .Z(n9199) );
  NAND U5348 ( .A(n9202), .B(n9199), .Z(n8394) );
  XNOR U5349 ( .A(n8809), .B(n8394), .Z(out[651]) );
  XNOR U5350 ( .A(in[314]), .B(n8395), .Z(n8816) );
  XNOR U5351 ( .A(in[1483]), .B(n8396), .Z(n9206) );
  XOR U5352 ( .A(n8397), .B(in[1094]), .Z(n9203) );
  NAND U5353 ( .A(n9206), .B(n9203), .Z(n8398) );
  XNOR U5354 ( .A(n8816), .B(n8398), .Z(out[652]) );
  XNOR U5355 ( .A(in[315]), .B(n8399), .Z(n8819) );
  XNOR U5356 ( .A(in[1484]), .B(n8400), .Z(n9210) );
  XOR U5357 ( .A(n8401), .B(in[1095]), .Z(n9207) );
  NAND U5358 ( .A(n9210), .B(n9207), .Z(n8402) );
  XNOR U5359 ( .A(n8819), .B(n8402), .Z(out[653]) );
  XNOR U5360 ( .A(in[316]), .B(n8403), .Z(n8822) );
  XNOR U5361 ( .A(in[1485]), .B(n8404), .Z(n9218) );
  XOR U5362 ( .A(n8405), .B(in[1096]), .Z(n9215) );
  NAND U5363 ( .A(n9218), .B(n9215), .Z(n8406) );
  XNOR U5364 ( .A(n8822), .B(n8406), .Z(out[654]) );
  XNOR U5365 ( .A(in[317]), .B(n8407), .Z(n8825) );
  XNOR U5366 ( .A(in[1486]), .B(n8408), .Z(n9222) );
  XOR U5367 ( .A(in[1097]), .B(n8409), .Z(n9219) );
  NAND U5368 ( .A(n9222), .B(n9219), .Z(n8410) );
  XNOR U5369 ( .A(n8825), .B(n8410), .Z(out[655]) );
  XNOR U5370 ( .A(in[318]), .B(n8411), .Z(n8828) );
  XNOR U5371 ( .A(in[1487]), .B(n8412), .Z(n9226) );
  XOR U5372 ( .A(n8413), .B(in[1098]), .Z(n9223) );
  NAND U5373 ( .A(n9226), .B(n9223), .Z(n8414) );
  XNOR U5374 ( .A(n8828), .B(n8414), .Z(out[656]) );
  XNOR U5375 ( .A(in[319]), .B(n8415), .Z(n8831) );
  XNOR U5376 ( .A(in[1488]), .B(n8416), .Z(n9230) );
  XOR U5377 ( .A(n8417), .B(in[1099]), .Z(n9227) );
  NAND U5378 ( .A(n9230), .B(n9227), .Z(n8418) );
  XNOR U5379 ( .A(n8831), .B(n8418), .Z(out[657]) );
  XNOR U5380 ( .A(in[256]), .B(n8419), .Z(n8834) );
  XNOR U5381 ( .A(in[1489]), .B(n8420), .Z(n9234) );
  XOR U5382 ( .A(in[1100]), .B(n8421), .Z(n9231) );
  NAND U5383 ( .A(n9234), .B(n9231), .Z(n8422) );
  XNOR U5384 ( .A(n8834), .B(n8422), .Z(out[658]) );
  XNOR U5385 ( .A(in[257]), .B(n8423), .Z(n8837) );
  XNOR U5386 ( .A(in[1490]), .B(n8424), .Z(n9238) );
  XOR U5387 ( .A(in[1101]), .B(n8425), .Z(n9235) );
  NAND U5388 ( .A(n9238), .B(n9235), .Z(n8426) );
  XNOR U5389 ( .A(n8837), .B(n8426), .Z(out[659]) );
  NOR U5390 ( .A(n8428), .B(n8427), .Z(n8429) );
  XNOR U5391 ( .A(n8430), .B(n8429), .Z(out[65]) );
  XNOR U5392 ( .A(in[258]), .B(n8431), .Z(n8840) );
  XOR U5393 ( .A(in[1491]), .B(n8432), .Z(n9242) );
  XOR U5394 ( .A(in[1102]), .B(n8433), .Z(n9239) );
  NAND U5395 ( .A(n9242), .B(n9239), .Z(n8434) );
  XNOR U5396 ( .A(n8840), .B(n8434), .Z(out[660]) );
  XNOR U5397 ( .A(in[259]), .B(n8435), .Z(n8843) );
  XOR U5398 ( .A(in[1492]), .B(n8436), .Z(n9246) );
  XOR U5399 ( .A(in[1103]), .B(n8437), .Z(n9243) );
  NAND U5400 ( .A(n9246), .B(n9243), .Z(n8438) );
  XNOR U5401 ( .A(n8843), .B(n8438), .Z(out[661]) );
  XOR U5402 ( .A(in[260]), .B(n8439), .Z(n8850) );
  XOR U5403 ( .A(in[1493]), .B(n8440), .Z(n9250) );
  XOR U5404 ( .A(in[1104]), .B(n8441), .Z(n9247) );
  NAND U5405 ( .A(n9250), .B(n9247), .Z(n8442) );
  XNOR U5406 ( .A(n8850), .B(n8442), .Z(out[662]) );
  XOR U5407 ( .A(in[261]), .B(n8443), .Z(n8853) );
  XOR U5408 ( .A(in[1494]), .B(n8444), .Z(n9254) );
  XOR U5409 ( .A(in[1105]), .B(n8445), .Z(n9251) );
  NAND U5410 ( .A(n9254), .B(n9251), .Z(n8446) );
  XNOR U5411 ( .A(n8853), .B(n8446), .Z(out[663]) );
  XOR U5412 ( .A(in[262]), .B(n8447), .Z(n8856) );
  XOR U5413 ( .A(in[1495]), .B(n8448), .Z(n9262) );
  XOR U5414 ( .A(in[1106]), .B(n8449), .Z(n9259) );
  NAND U5415 ( .A(n9262), .B(n9259), .Z(n8450) );
  XNOR U5416 ( .A(n8856), .B(n8450), .Z(out[664]) );
  XOR U5417 ( .A(in[263]), .B(n8451), .Z(n8859) );
  XOR U5418 ( .A(in[1496]), .B(n8452), .Z(n9266) );
  XOR U5419 ( .A(in[1107]), .B(n8453), .Z(n9263) );
  NAND U5420 ( .A(n9266), .B(n9263), .Z(n8454) );
  XNOR U5421 ( .A(n8859), .B(n8454), .Z(out[665]) );
  XOR U5422 ( .A(in[264]), .B(n8455), .Z(n8862) );
  XOR U5423 ( .A(in[1497]), .B(n8456), .Z(n9270) );
  XOR U5424 ( .A(in[1108]), .B(n8457), .Z(n9267) );
  NAND U5425 ( .A(n9270), .B(n9267), .Z(n8458) );
  XNOR U5426 ( .A(n8862), .B(n8458), .Z(out[666]) );
  XOR U5427 ( .A(in[265]), .B(n8459), .Z(n8865) );
  XOR U5428 ( .A(in[1498]), .B(n8460), .Z(n9274) );
  XOR U5429 ( .A(in[1109]), .B(n8461), .Z(n9271) );
  NAND U5430 ( .A(n9274), .B(n9271), .Z(n8462) );
  XNOR U5431 ( .A(n8865), .B(n8462), .Z(out[667]) );
  XOR U5432 ( .A(in[266]), .B(n8463), .Z(n8868) );
  XOR U5433 ( .A(in[1499]), .B(n8464), .Z(n9278) );
  XOR U5434 ( .A(in[1110]), .B(n8465), .Z(n9275) );
  NAND U5435 ( .A(n9278), .B(n9275), .Z(n8466) );
  XNOR U5436 ( .A(n8868), .B(n8466), .Z(out[668]) );
  XOR U5437 ( .A(in[267]), .B(n8467), .Z(n8871) );
  XOR U5438 ( .A(in[1500]), .B(n8468), .Z(n9282) );
  XOR U5439 ( .A(in[1111]), .B(n8469), .Z(n9279) );
  NAND U5440 ( .A(n9282), .B(n9279), .Z(n8470) );
  XNOR U5441 ( .A(n8871), .B(n8470), .Z(out[669]) );
  ANDN U5442 ( .B(n8472), .A(n8471), .Z(n8473) );
  XNOR U5443 ( .A(n8474), .B(n8473), .Z(out[66]) );
  XOR U5444 ( .A(in[268]), .B(n8475), .Z(n8874) );
  XOR U5445 ( .A(in[1501]), .B(n8476), .Z(n9286) );
  XOR U5446 ( .A(in[1112]), .B(n8477), .Z(n9283) );
  NAND U5447 ( .A(n9286), .B(n9283), .Z(n8478) );
  XNOR U5448 ( .A(n8874), .B(n8478), .Z(out[670]) );
  XOR U5449 ( .A(in[269]), .B(n8479), .Z(n8877) );
  XOR U5450 ( .A(in[1502]), .B(n8480), .Z(n9290) );
  XOR U5451 ( .A(in[1113]), .B(n8481), .Z(n9287) );
  NAND U5452 ( .A(n9290), .B(n9287), .Z(n8482) );
  XNOR U5453 ( .A(n8877), .B(n8482), .Z(out[671]) );
  XOR U5454 ( .A(in[270]), .B(n8483), .Z(n8888) );
  XOR U5455 ( .A(in[1503]), .B(n8484), .Z(n9294) );
  XOR U5456 ( .A(in[1114]), .B(n8485), .Z(n9291) );
  NAND U5457 ( .A(n9294), .B(n9291), .Z(n8486) );
  XNOR U5458 ( .A(n8888), .B(n8486), .Z(out[672]) );
  XOR U5459 ( .A(in[271]), .B(n8487), .Z(n8891) );
  XOR U5460 ( .A(in[1504]), .B(n8488), .Z(n9298) );
  XOR U5461 ( .A(in[1115]), .B(n8489), .Z(n9295) );
  NAND U5462 ( .A(n9298), .B(n9295), .Z(n8490) );
  XNOR U5463 ( .A(n8891), .B(n8490), .Z(out[673]) );
  XOR U5464 ( .A(in[272]), .B(n8491), .Z(n8894) );
  XOR U5465 ( .A(in[1505]), .B(n8492), .Z(n9306) );
  XOR U5466 ( .A(in[1116]), .B(n8493), .Z(n9303) );
  NAND U5467 ( .A(n9306), .B(n9303), .Z(n8494) );
  XNOR U5468 ( .A(n8894), .B(n8494), .Z(out[674]) );
  XOR U5469 ( .A(in[273]), .B(n8495), .Z(n8897) );
  XNOR U5470 ( .A(n8496), .B(in[1506]), .Z(n9310) );
  XOR U5471 ( .A(in[1117]), .B(n8497), .Z(n9307) );
  NAND U5472 ( .A(n9310), .B(n9307), .Z(n8498) );
  XNOR U5473 ( .A(n8897), .B(n8498), .Z(out[675]) );
  XOR U5474 ( .A(in[274]), .B(n8499), .Z(n8900) );
  XNOR U5475 ( .A(n8500), .B(in[1507]), .Z(n9314) );
  XOR U5476 ( .A(in[1118]), .B(n8501), .Z(n9311) );
  NAND U5477 ( .A(n9314), .B(n9311), .Z(n8502) );
  XNOR U5478 ( .A(n8900), .B(n8502), .Z(out[676]) );
  XOR U5479 ( .A(in[275]), .B(n8503), .Z(n8903) );
  XNOR U5480 ( .A(n8504), .B(in[1508]), .Z(n9318) );
  XOR U5481 ( .A(in[1119]), .B(n8505), .Z(n9315) );
  NAND U5482 ( .A(n9318), .B(n9315), .Z(n8506) );
  XNOR U5483 ( .A(n8903), .B(n8506), .Z(out[677]) );
  XOR U5484 ( .A(in[276]), .B(n8507), .Z(n8906) );
  XNOR U5485 ( .A(n8508), .B(in[1509]), .Z(n9322) );
  XOR U5486 ( .A(in[1120]), .B(n8509), .Z(n9319) );
  NAND U5487 ( .A(n9322), .B(n9319), .Z(n8510) );
  XNOR U5488 ( .A(n8906), .B(n8510), .Z(out[678]) );
  XOR U5489 ( .A(in[277]), .B(n8511), .Z(n8909) );
  XOR U5490 ( .A(in[1510]), .B(n8512), .Z(n9326) );
  XOR U5491 ( .A(in[1121]), .B(n8513), .Z(n9323) );
  NAND U5492 ( .A(n9326), .B(n9323), .Z(n8514) );
  XNOR U5493 ( .A(n8909), .B(n8514), .Z(out[679]) );
  ANDN U5494 ( .B(n8516), .A(n8515), .Z(n8517) );
  XNOR U5495 ( .A(n8518), .B(n8517), .Z(out[67]) );
  XOR U5496 ( .A(in[278]), .B(n8519), .Z(n8912) );
  XOR U5497 ( .A(in[1511]), .B(n8520), .Z(n9330) );
  XOR U5498 ( .A(in[1122]), .B(n8521), .Z(n9327) );
  NAND U5499 ( .A(n9330), .B(n9327), .Z(n8522) );
  XNOR U5500 ( .A(n8912), .B(n8522), .Z(out[680]) );
  XOR U5501 ( .A(in[279]), .B(n8523), .Z(n8915) );
  XOR U5502 ( .A(in[1512]), .B(n8524), .Z(n9334) );
  XOR U5503 ( .A(in[1123]), .B(n8525), .Z(n9331) );
  NAND U5504 ( .A(n9334), .B(n9331), .Z(n8526) );
  XNOR U5505 ( .A(n8915), .B(n8526), .Z(out[681]) );
  XOR U5506 ( .A(in[280]), .B(n8527), .Z(n8922) );
  XOR U5507 ( .A(in[1513]), .B(n8528), .Z(n9338) );
  XOR U5508 ( .A(in[1124]), .B(n8529), .Z(n9335) );
  NAND U5509 ( .A(n9338), .B(n9335), .Z(n8530) );
  XNOR U5510 ( .A(n8922), .B(n8530), .Z(out[682]) );
  XOR U5511 ( .A(in[281]), .B(n8531), .Z(n8925) );
  XOR U5512 ( .A(in[1514]), .B(n8532), .Z(n9342) );
  XOR U5513 ( .A(in[1125]), .B(n8533), .Z(n9339) );
  NAND U5514 ( .A(n9342), .B(n9339), .Z(n8534) );
  XNOR U5515 ( .A(n8925), .B(n8534), .Z(out[683]) );
  XOR U5516 ( .A(in[282]), .B(n8535), .Z(n8928) );
  XOR U5517 ( .A(in[1515]), .B(n8536), .Z(n9350) );
  XNOR U5518 ( .A(in[1126]), .B(n8537), .Z(n9347) );
  NAND U5519 ( .A(n9350), .B(n9347), .Z(n8538) );
  XNOR U5520 ( .A(n8928), .B(n8538), .Z(out[684]) );
  XOR U5521 ( .A(in[283]), .B(n8539), .Z(n8931) );
  XOR U5522 ( .A(in[1516]), .B(n8540), .Z(n9354) );
  XNOR U5523 ( .A(in[1127]), .B(n8541), .Z(n9351) );
  NAND U5524 ( .A(n9354), .B(n9351), .Z(n8542) );
  XNOR U5525 ( .A(n8931), .B(n8542), .Z(out[685]) );
  XOR U5526 ( .A(in[284]), .B(n8543), .Z(n8934) );
  XOR U5527 ( .A(in[1517]), .B(n8544), .Z(n9358) );
  XNOR U5528 ( .A(in[1128]), .B(n8545), .Z(n9355) );
  NAND U5529 ( .A(n9358), .B(n9355), .Z(n8546) );
  XNOR U5530 ( .A(n8934), .B(n8546), .Z(out[686]) );
  XOR U5531 ( .A(in[285]), .B(n8547), .Z(n8937) );
  XOR U5532 ( .A(in[1518]), .B(n8548), .Z(n9362) );
  XNOR U5533 ( .A(in[1129]), .B(n8549), .Z(n9359) );
  NAND U5534 ( .A(n9362), .B(n9359), .Z(n8550) );
  XNOR U5535 ( .A(n8937), .B(n8550), .Z(out[687]) );
  XOR U5536 ( .A(in[286]), .B(n8551), .Z(n8940) );
  XOR U5537 ( .A(in[1519]), .B(n8552), .Z(n9366) );
  XNOR U5538 ( .A(in[1130]), .B(n8553), .Z(n9363) );
  NAND U5539 ( .A(n9366), .B(n9363), .Z(n8554) );
  XNOR U5540 ( .A(n8940), .B(n8554), .Z(out[688]) );
  XOR U5541 ( .A(in[287]), .B(n8555), .Z(n8943) );
  XOR U5542 ( .A(in[1520]), .B(n8556), .Z(n9370) );
  XNOR U5543 ( .A(in[1131]), .B(n8557), .Z(n9367) );
  NAND U5544 ( .A(n9370), .B(n9367), .Z(n8558) );
  XNOR U5545 ( .A(n8943), .B(n8558), .Z(out[689]) );
  ANDN U5546 ( .B(n8560), .A(n8559), .Z(n8561) );
  XNOR U5547 ( .A(n8562), .B(n8561), .Z(out[68]) );
  XOR U5548 ( .A(in[288]), .B(n8563), .Z(n8946) );
  XOR U5549 ( .A(in[1521]), .B(n8564), .Z(n9374) );
  XNOR U5550 ( .A(in[1132]), .B(n8565), .Z(n9371) );
  NAND U5551 ( .A(n9374), .B(n9371), .Z(n8566) );
  XNOR U5552 ( .A(n8946), .B(n8566), .Z(out[690]) );
  XOR U5553 ( .A(in[289]), .B(n8567), .Z(n8949) );
  XOR U5554 ( .A(in[1522]), .B(n8568), .Z(n9378) );
  XNOR U5555 ( .A(in[1133]), .B(n8569), .Z(n9375) );
  NAND U5556 ( .A(n9378), .B(n9375), .Z(n8570) );
  XNOR U5557 ( .A(n8949), .B(n8570), .Z(out[691]) );
  XOR U5558 ( .A(in[290]), .B(n8571), .Z(n8956) );
  XOR U5559 ( .A(in[1523]), .B(n8572), .Z(n9382) );
  XNOR U5560 ( .A(in[1134]), .B(n8573), .Z(n9379) );
  NAND U5561 ( .A(n9382), .B(n9379), .Z(n8574) );
  XNOR U5562 ( .A(n8956), .B(n8574), .Z(out[692]) );
  XOR U5563 ( .A(in[291]), .B(n8575), .Z(n8959) );
  XOR U5564 ( .A(in[1524]), .B(n8576), .Z(n9386) );
  XNOR U5565 ( .A(in[1135]), .B(n8577), .Z(n9383) );
  NAND U5566 ( .A(n9386), .B(n9383), .Z(n8578) );
  XNOR U5567 ( .A(n8959), .B(n8578), .Z(out[693]) );
  XOR U5568 ( .A(in[292]), .B(n8579), .Z(n8962) );
  XOR U5569 ( .A(in[1525]), .B(n8580), .Z(n9394) );
  XNOR U5570 ( .A(in[1136]), .B(n8581), .Z(n9391) );
  NAND U5571 ( .A(n9394), .B(n9391), .Z(n8582) );
  XNOR U5572 ( .A(n8962), .B(n8582), .Z(out[694]) );
  XNOR U5573 ( .A(in[293]), .B(n8583), .Z(n8965) );
  XOR U5574 ( .A(in[1526]), .B(n8584), .Z(n9398) );
  XNOR U5575 ( .A(in[1137]), .B(n8585), .Z(n9395) );
  NAND U5576 ( .A(n9398), .B(n9395), .Z(n8586) );
  XNOR U5577 ( .A(n8965), .B(n8586), .Z(out[695]) );
  XNOR U5578 ( .A(in[294]), .B(n8587), .Z(n8968) );
  XOR U5579 ( .A(in[1527]), .B(n8588), .Z(n9402) );
  XNOR U5580 ( .A(in[1138]), .B(n8589), .Z(n9399) );
  NAND U5581 ( .A(n9402), .B(n9399), .Z(n8590) );
  XNOR U5582 ( .A(n8968), .B(n8590), .Z(out[696]) );
  XNOR U5583 ( .A(in[295]), .B(n8591), .Z(n8971) );
  XOR U5584 ( .A(in[1528]), .B(n8592), .Z(n9406) );
  XNOR U5585 ( .A(in[1139]), .B(n8593), .Z(n9403) );
  NAND U5586 ( .A(n9406), .B(n9403), .Z(n8594) );
  XNOR U5587 ( .A(n8971), .B(n8594), .Z(out[697]) );
  XNOR U5588 ( .A(in[296]), .B(n8595), .Z(n8974) );
  XOR U5589 ( .A(in[1529]), .B(n8596), .Z(n9410) );
  XNOR U5590 ( .A(in[1140]), .B(n8597), .Z(n9407) );
  NAND U5591 ( .A(n9410), .B(n9407), .Z(n8598) );
  XNOR U5592 ( .A(n8974), .B(n8598), .Z(out[698]) );
  XNOR U5593 ( .A(in[297]), .B(n8599), .Z(n8977) );
  XOR U5594 ( .A(in[1530]), .B(n8600), .Z(n9414) );
  XNOR U5595 ( .A(in[1141]), .B(n8601), .Z(n9411) );
  NAND U5596 ( .A(n9414), .B(n9411), .Z(n8602) );
  XNOR U5597 ( .A(n8977), .B(n8602), .Z(out[699]) );
  ANDN U5598 ( .B(n8604), .A(n8603), .Z(n8605) );
  XNOR U5599 ( .A(n8606), .B(n8605), .Z(out[69]) );
  OR U5600 ( .A(n8638), .B(n8607), .Z(n8608) );
  XNOR U5601 ( .A(n8637), .B(n8608), .Z(out[6]) );
  XNOR U5602 ( .A(in[298]), .B(n8609), .Z(n8980) );
  XNOR U5603 ( .A(in[1531]), .B(n8610), .Z(n9418) );
  XNOR U5604 ( .A(in[1142]), .B(n8611), .Z(n9415) );
  NAND U5605 ( .A(n9418), .B(n9415), .Z(n8612) );
  XNOR U5606 ( .A(n8980), .B(n8612), .Z(out[700]) );
  XNOR U5607 ( .A(in[299]), .B(n8613), .Z(n8983) );
  XNOR U5608 ( .A(in[1532]), .B(n8614), .Z(n9422) );
  XNOR U5609 ( .A(in[1143]), .B(n8615), .Z(n9419) );
  NAND U5610 ( .A(n9422), .B(n9419), .Z(n8616) );
  XNOR U5611 ( .A(n8983), .B(n8616), .Z(out[701]) );
  XNOR U5612 ( .A(in[300]), .B(n8617), .Z(n8990) );
  XNOR U5613 ( .A(in[1533]), .B(n8618), .Z(n9426) );
  XNOR U5614 ( .A(in[1144]), .B(n8619), .Z(n9423) );
  NAND U5615 ( .A(n9426), .B(n9423), .Z(n8620) );
  XNOR U5616 ( .A(n8990), .B(n8620), .Z(out[702]) );
  XNOR U5617 ( .A(in[301]), .B(n8621), .Z(n8993) );
  XOR U5618 ( .A(in[1534]), .B(n8622), .Z(n9430) );
  XNOR U5619 ( .A(in[1145]), .B(n8623), .Z(n9427) );
  NAND U5620 ( .A(n9430), .B(n9427), .Z(n8624) );
  XNOR U5621 ( .A(n8993), .B(n8624), .Z(out[703]) );
  XOR U5622 ( .A(in[376]), .B(n8625), .Z(n8995) );
  NOR U5623 ( .A(n8772), .B(n9150), .Z(n8626) );
  XNOR U5624 ( .A(n8995), .B(n8626), .Z(out[704]) );
  XOR U5625 ( .A(in[377]), .B(n8627), .Z(n8997) );
  NOR U5626 ( .A(n8775), .B(n9154), .Z(n8628) );
  XNOR U5627 ( .A(n8997), .B(n8628), .Z(out[705]) );
  XOR U5628 ( .A(in[378]), .B(n8629), .Z(n8999) );
  NOR U5629 ( .A(n8782), .B(n9158), .Z(n8630) );
  XNOR U5630 ( .A(n8999), .B(n8630), .Z(out[706]) );
  XOR U5631 ( .A(in[379]), .B(n8631), .Z(n9001) );
  NOR U5632 ( .A(n8785), .B(n9162), .Z(n8632) );
  XNOR U5633 ( .A(n9001), .B(n8632), .Z(out[707]) );
  XOR U5634 ( .A(in[380]), .B(n8633), .Z(n9003) );
  NOR U5635 ( .A(n8788), .B(n9174), .Z(n8634) );
  XNOR U5636 ( .A(n9003), .B(n8634), .Z(out[708]) );
  XOR U5637 ( .A(in[381]), .B(n8635), .Z(n9005) );
  NOR U5638 ( .A(n8791), .B(n9178), .Z(n8636) );
  XNOR U5639 ( .A(n9005), .B(n8636), .Z(out[709]) );
  ANDN U5640 ( .B(n8638), .A(n8637), .Z(n8639) );
  XNOR U5641 ( .A(n8640), .B(n8639), .Z(out[70]) );
  XOR U5642 ( .A(in[382]), .B(n8641), .Z(n9007) );
  NOR U5643 ( .A(n8794), .B(n9182), .Z(n8642) );
  XNOR U5644 ( .A(n9007), .B(n8642), .Z(out[710]) );
  XOR U5645 ( .A(in[383]), .B(n8643), .Z(n9009) );
  NOR U5646 ( .A(n8797), .B(n9186), .Z(n8644) );
  XNOR U5647 ( .A(n9009), .B(n8644), .Z(out[711]) );
  XOR U5648 ( .A(in[320]), .B(n8645), .Z(n9015) );
  NOR U5649 ( .A(n8800), .B(n9190), .Z(n8646) );
  XNOR U5650 ( .A(n9015), .B(n8646), .Z(out[712]) );
  XOR U5651 ( .A(in[321]), .B(n8647), .Z(n9017) );
  NOR U5652 ( .A(n8803), .B(n9194), .Z(n8648) );
  XNOR U5653 ( .A(n9017), .B(n8648), .Z(out[713]) );
  XOR U5654 ( .A(in[322]), .B(n8649), .Z(n9019) );
  NOR U5655 ( .A(n8806), .B(n9198), .Z(n8650) );
  XNOR U5656 ( .A(n9019), .B(n8650), .Z(out[714]) );
  XOR U5657 ( .A(in[323]), .B(n8651), .Z(n9021) );
  NOR U5658 ( .A(n8809), .B(n9202), .Z(n8652) );
  XNOR U5659 ( .A(n9021), .B(n8652), .Z(out[715]) );
  XOR U5660 ( .A(in[324]), .B(n8653), .Z(n9023) );
  NOR U5661 ( .A(n8816), .B(n9206), .Z(n8654) );
  XNOR U5662 ( .A(n9023), .B(n8654), .Z(out[716]) );
  XOR U5663 ( .A(in[325]), .B(n8655), .Z(n9025) );
  NOR U5664 ( .A(n8819), .B(n9210), .Z(n8656) );
  XNOR U5665 ( .A(n9025), .B(n8656), .Z(out[717]) );
  XOR U5666 ( .A(in[326]), .B(n8657), .Z(n9027) );
  NOR U5667 ( .A(n8822), .B(n9218), .Z(n8658) );
  XNOR U5668 ( .A(n9027), .B(n8658), .Z(out[718]) );
  XOR U5669 ( .A(in[327]), .B(n8659), .Z(n9029) );
  NOR U5670 ( .A(n8825), .B(n9222), .Z(n8660) );
  XNOR U5671 ( .A(n9029), .B(n8660), .Z(out[719]) );
  ANDN U5672 ( .B(n8884), .A(n8886), .Z(n8661) );
  XNOR U5673 ( .A(n8662), .B(n8661), .Z(out[71]) );
  XOR U5674 ( .A(in[328]), .B(n8663), .Z(n9031) );
  NOR U5675 ( .A(n8828), .B(n9226), .Z(n8664) );
  XNOR U5676 ( .A(n9031), .B(n8664), .Z(out[720]) );
  XOR U5677 ( .A(in[329]), .B(n8665), .Z(n9033) );
  NOR U5678 ( .A(n8831), .B(n9230), .Z(n8666) );
  XNOR U5679 ( .A(n9033), .B(n8666), .Z(out[721]) );
  XOR U5680 ( .A(in[330]), .B(n8667), .Z(n9039) );
  NOR U5681 ( .A(n8834), .B(n9234), .Z(n8668) );
  XNOR U5682 ( .A(n9039), .B(n8668), .Z(out[722]) );
  XOR U5683 ( .A(in[331]), .B(n8669), .Z(n9041) );
  NOR U5684 ( .A(n8837), .B(n9238), .Z(n8670) );
  XNOR U5685 ( .A(n9041), .B(n8670), .Z(out[723]) );
  XOR U5686 ( .A(in[332]), .B(n8671), .Z(n9043) );
  NOR U5687 ( .A(n8840), .B(n9242), .Z(n8672) );
  XNOR U5688 ( .A(n9043), .B(n8672), .Z(out[724]) );
  XOR U5689 ( .A(in[333]), .B(n8673), .Z(n9045) );
  NOR U5690 ( .A(n8843), .B(n9246), .Z(n8674) );
  XNOR U5691 ( .A(n9045), .B(n8674), .Z(out[725]) );
  XOR U5692 ( .A(in[334]), .B(n8675), .Z(n9047) );
  NOR U5693 ( .A(n8850), .B(n9250), .Z(n8676) );
  XNOR U5694 ( .A(n9047), .B(n8676), .Z(out[726]) );
  XOR U5695 ( .A(in[335]), .B(n8677), .Z(n9049) );
  NOR U5696 ( .A(n8853), .B(n9254), .Z(n8678) );
  XNOR U5697 ( .A(n9049), .B(n8678), .Z(out[727]) );
  XOR U5698 ( .A(in[336]), .B(n8679), .Z(n9051) );
  NOR U5699 ( .A(n8856), .B(n9262), .Z(n8680) );
  XNOR U5700 ( .A(n9051), .B(n8680), .Z(out[728]) );
  XOR U5701 ( .A(in[337]), .B(n8681), .Z(n9053) );
  NOR U5702 ( .A(n8859), .B(n9266), .Z(n8682) );
  XNOR U5703 ( .A(n9053), .B(n8682), .Z(out[729]) );
  ANDN U5704 ( .B(n9168), .A(n9170), .Z(n8683) );
  XNOR U5705 ( .A(n8684), .B(n8683), .Z(out[72]) );
  XOR U5706 ( .A(in[338]), .B(n8685), .Z(n9055) );
  NOR U5707 ( .A(n8862), .B(n9270), .Z(n8686) );
  XNOR U5708 ( .A(n9055), .B(n8686), .Z(out[730]) );
  XOR U5709 ( .A(in[339]), .B(n8687), .Z(n9057) );
  NOR U5710 ( .A(n8865), .B(n9274), .Z(n8688) );
  XNOR U5711 ( .A(n9057), .B(n8688), .Z(out[731]) );
  XOR U5712 ( .A(in[340]), .B(n8689), .Z(n9063) );
  NOR U5713 ( .A(n8868), .B(n9278), .Z(n8690) );
  XNOR U5714 ( .A(n9063), .B(n8690), .Z(out[732]) );
  XOR U5715 ( .A(in[341]), .B(n8691), .Z(n9065) );
  NOR U5716 ( .A(n8871), .B(n9282), .Z(n8692) );
  XNOR U5717 ( .A(n9065), .B(n8692), .Z(out[733]) );
  XOR U5718 ( .A(in[342]), .B(n8693), .Z(n9067) );
  NOR U5719 ( .A(n8874), .B(n9286), .Z(n8694) );
  XNOR U5720 ( .A(n9067), .B(n8694), .Z(out[734]) );
  XOR U5721 ( .A(in[343]), .B(n8695), .Z(n9069) );
  NOR U5722 ( .A(n8877), .B(n9290), .Z(n8696) );
  XNOR U5723 ( .A(n9069), .B(n8696), .Z(out[735]) );
  XOR U5724 ( .A(in[344]), .B(n8697), .Z(n9071) );
  NOR U5725 ( .A(n8888), .B(n9294), .Z(n8698) );
  XNOR U5726 ( .A(n9071), .B(n8698), .Z(out[736]) );
  XOR U5727 ( .A(in[345]), .B(n8699), .Z(n9073) );
  NOR U5728 ( .A(n8891), .B(n9298), .Z(n8700) );
  XNOR U5729 ( .A(n9073), .B(n8700), .Z(out[737]) );
  XOR U5730 ( .A(in[346]), .B(n8701), .Z(n9075) );
  NOR U5731 ( .A(n8894), .B(n9306), .Z(n8702) );
  XNOR U5732 ( .A(n9075), .B(n8702), .Z(out[738]) );
  XOR U5733 ( .A(in[347]), .B(n8703), .Z(n9077) );
  NOR U5734 ( .A(n8897), .B(n9310), .Z(n8704) );
  XNOR U5735 ( .A(n9077), .B(n8704), .Z(out[739]) );
  ANDN U5736 ( .B(n9612), .A(n9614), .Z(n8705) );
  XNOR U5737 ( .A(n8706), .B(n8705), .Z(out[73]) );
  XOR U5738 ( .A(in[348]), .B(n8707), .Z(n9079) );
  NOR U5739 ( .A(n8900), .B(n9314), .Z(n8708) );
  XNOR U5740 ( .A(n9079), .B(n8708), .Z(out[740]) );
  XOR U5741 ( .A(in[349]), .B(n8709), .Z(n9081) );
  NOR U5742 ( .A(n8903), .B(n9318), .Z(n8710) );
  XNOR U5743 ( .A(n9081), .B(n8710), .Z(out[741]) );
  XOR U5744 ( .A(in[350]), .B(n8711), .Z(n9087) );
  NOR U5745 ( .A(n8906), .B(n9322), .Z(n8712) );
  XNOR U5746 ( .A(n9087), .B(n8712), .Z(out[742]) );
  XOR U5747 ( .A(in[351]), .B(n8713), .Z(n9089) );
  NOR U5748 ( .A(n8909), .B(n9326), .Z(n8714) );
  XNOR U5749 ( .A(n9089), .B(n8714), .Z(out[743]) );
  XOR U5750 ( .A(in[352]), .B(n8715), .Z(n9091) );
  NOR U5751 ( .A(n8912), .B(n9330), .Z(n8716) );
  XNOR U5752 ( .A(n9091), .B(n8716), .Z(out[744]) );
  XOR U5753 ( .A(in[353]), .B(n8717), .Z(n9093) );
  NOR U5754 ( .A(n8915), .B(n9334), .Z(n8718) );
  XNOR U5755 ( .A(n9093), .B(n8718), .Z(out[745]) );
  XOR U5756 ( .A(in[354]), .B(n8719), .Z(n9095) );
  NOR U5757 ( .A(n8922), .B(n9338), .Z(n8720) );
  XNOR U5758 ( .A(n9095), .B(n8720), .Z(out[746]) );
  XOR U5759 ( .A(in[355]), .B(n8721), .Z(n9097) );
  NOR U5760 ( .A(n8925), .B(n9342), .Z(n8722) );
  XNOR U5761 ( .A(n9097), .B(n8722), .Z(out[747]) );
  XOR U5762 ( .A(in[356]), .B(n8723), .Z(n9099) );
  NOR U5763 ( .A(n8928), .B(n9350), .Z(n8724) );
  XNOR U5764 ( .A(n9099), .B(n8724), .Z(out[748]) );
  XOR U5765 ( .A(in[357]), .B(n8725), .Z(n9101) );
  NOR U5766 ( .A(n8931), .B(n9354), .Z(n8726) );
  XNOR U5767 ( .A(n9101), .B(n8726), .Z(out[749]) );
  NOR U5768 ( .A(n8728), .B(n8727), .Z(n8729) );
  XNOR U5769 ( .A(n8730), .B(n8729), .Z(out[74]) );
  XOR U5770 ( .A(in[358]), .B(n8731), .Z(n9103) );
  NOR U5771 ( .A(n8934), .B(n9358), .Z(n8732) );
  XNOR U5772 ( .A(n9103), .B(n8732), .Z(out[750]) );
  XOR U5773 ( .A(in[359]), .B(n8733), .Z(n9105) );
  NOR U5774 ( .A(n8937), .B(n9362), .Z(n8734) );
  XNOR U5775 ( .A(n9105), .B(n8734), .Z(out[751]) );
  XOR U5776 ( .A(in[360]), .B(n8735), .Z(n9111) );
  NOR U5777 ( .A(n8940), .B(n9366), .Z(n8736) );
  XNOR U5778 ( .A(n9111), .B(n8736), .Z(out[752]) );
  XOR U5779 ( .A(in[361]), .B(n8737), .Z(n9113) );
  NOR U5780 ( .A(n8943), .B(n9370), .Z(n8738) );
  XNOR U5781 ( .A(n9113), .B(n8738), .Z(out[753]) );
  XOR U5782 ( .A(in[362]), .B(n8739), .Z(n9115) );
  NOR U5783 ( .A(n8946), .B(n9374), .Z(n8740) );
  XNOR U5784 ( .A(n9115), .B(n8740), .Z(out[754]) );
  XOR U5785 ( .A(in[363]), .B(n8741), .Z(n9117) );
  NOR U5786 ( .A(n8949), .B(n9378), .Z(n8742) );
  XNOR U5787 ( .A(n9117), .B(n8742), .Z(out[755]) );
  XOR U5788 ( .A(in[364]), .B(n8743), .Z(n9119) );
  NOR U5789 ( .A(n8956), .B(n9382), .Z(n8744) );
  XNOR U5790 ( .A(n9119), .B(n8744), .Z(out[756]) );
  XOR U5791 ( .A(in[365]), .B(n8745), .Z(n9121) );
  NOR U5792 ( .A(n8959), .B(n9386), .Z(n8746) );
  XNOR U5793 ( .A(n9121), .B(n8746), .Z(out[757]) );
  XOR U5794 ( .A(in[366]), .B(n8747), .Z(n9123) );
  NOR U5795 ( .A(n8962), .B(n9394), .Z(n8748) );
  XNOR U5796 ( .A(n9123), .B(n8748), .Z(out[758]) );
  XOR U5797 ( .A(in[367]), .B(n8749), .Z(n9125) );
  NOR U5798 ( .A(n8965), .B(n9398), .Z(n8750) );
  XNOR U5799 ( .A(n9125), .B(n8750), .Z(out[759]) );
  NOR U5800 ( .A(n8752), .B(n8751), .Z(n8753) );
  XNOR U5801 ( .A(n8754), .B(n8753), .Z(out[75]) );
  XOR U5802 ( .A(in[368]), .B(n8755), .Z(n9127) );
  NOR U5803 ( .A(n8968), .B(n9402), .Z(n8756) );
  XNOR U5804 ( .A(n9127), .B(n8756), .Z(out[760]) );
  XOR U5805 ( .A(in[369]), .B(n8757), .Z(n9129) );
  NOR U5806 ( .A(n8971), .B(n9406), .Z(n8758) );
  XNOR U5807 ( .A(n9129), .B(n8758), .Z(out[761]) );
  XOR U5808 ( .A(in[370]), .B(n8759), .Z(n9135) );
  NOR U5809 ( .A(n8974), .B(n9410), .Z(n8760) );
  XNOR U5810 ( .A(n9135), .B(n8760), .Z(out[762]) );
  XOR U5811 ( .A(in[371]), .B(n8761), .Z(n9137) );
  NOR U5812 ( .A(n8977), .B(n9414), .Z(n8762) );
  XNOR U5813 ( .A(n9137), .B(n8762), .Z(out[763]) );
  XOR U5814 ( .A(in[372]), .B(n8763), .Z(n9139) );
  NOR U5815 ( .A(n8980), .B(n9418), .Z(n8764) );
  XNOR U5816 ( .A(n9139), .B(n8764), .Z(out[764]) );
  XOR U5817 ( .A(in[373]), .B(n8765), .Z(n9141) );
  NOR U5818 ( .A(n8983), .B(n9422), .Z(n8766) );
  XNOR U5819 ( .A(n9141), .B(n8766), .Z(out[765]) );
  XOR U5820 ( .A(in[374]), .B(n8767), .Z(n9143) );
  NOR U5821 ( .A(n8990), .B(n9426), .Z(n8768) );
  XNOR U5822 ( .A(n9143), .B(n8768), .Z(out[766]) );
  XOR U5823 ( .A(in[375]), .B(n8769), .Z(n9145) );
  NOR U5824 ( .A(n8993), .B(n9430), .Z(n8770) );
  XNOR U5825 ( .A(n9145), .B(n8770), .Z(out[767]) );
  XNOR U5826 ( .A(in[743]), .B(n8771), .Z(n9148) );
  NAND U5827 ( .A(n8995), .B(n8772), .Z(n8773) );
  XNOR U5828 ( .A(n9148), .B(n8773), .Z(out[768]) );
  XNOR U5829 ( .A(in[744]), .B(n8774), .Z(n9152) );
  NAND U5830 ( .A(n8997), .B(n8775), .Z(n8776) );
  XNOR U5831 ( .A(n9152), .B(n8776), .Z(out[769]) );
  NOR U5832 ( .A(n8778), .B(n8777), .Z(n8779) );
  XNOR U5833 ( .A(n8780), .B(n8779), .Z(out[76]) );
  XNOR U5834 ( .A(in[745]), .B(n8781), .Z(n9156) );
  NAND U5835 ( .A(n8999), .B(n8782), .Z(n8783) );
  XNOR U5836 ( .A(n9156), .B(n8783), .Z(out[770]) );
  XNOR U5837 ( .A(in[746]), .B(n8784), .Z(n9160) );
  NAND U5838 ( .A(n9001), .B(n8785), .Z(n8786) );
  XNOR U5839 ( .A(n9160), .B(n8786), .Z(out[771]) );
  XNOR U5840 ( .A(in[747]), .B(n8787), .Z(n9172) );
  NAND U5841 ( .A(n9003), .B(n8788), .Z(n8789) );
  XNOR U5842 ( .A(n9172), .B(n8789), .Z(out[772]) );
  XNOR U5843 ( .A(in[748]), .B(n8790), .Z(n9176) );
  NAND U5844 ( .A(n9005), .B(n8791), .Z(n8792) );
  XNOR U5845 ( .A(n9176), .B(n8792), .Z(out[773]) );
  XNOR U5846 ( .A(in[749]), .B(n8793), .Z(n9180) );
  NAND U5847 ( .A(n9007), .B(n8794), .Z(n8795) );
  XNOR U5848 ( .A(n9180), .B(n8795), .Z(out[774]) );
  XNOR U5849 ( .A(in[750]), .B(n8796), .Z(n9184) );
  NAND U5850 ( .A(n9009), .B(n8797), .Z(n8798) );
  XNOR U5851 ( .A(n9184), .B(n8798), .Z(out[775]) );
  XNOR U5852 ( .A(in[751]), .B(n8799), .Z(n9188) );
  NAND U5853 ( .A(n9015), .B(n8800), .Z(n8801) );
  XNOR U5854 ( .A(n9188), .B(n8801), .Z(out[776]) );
  XNOR U5855 ( .A(in[752]), .B(n8802), .Z(n9192) );
  NAND U5856 ( .A(n9017), .B(n8803), .Z(n8804) );
  XNOR U5857 ( .A(n9192), .B(n8804), .Z(out[777]) );
  XNOR U5858 ( .A(in[753]), .B(n8805), .Z(n9196) );
  NAND U5859 ( .A(n9019), .B(n8806), .Z(n8807) );
  XNOR U5860 ( .A(n9196), .B(n8807), .Z(out[778]) );
  XNOR U5861 ( .A(in[754]), .B(n8808), .Z(n9200) );
  NAND U5862 ( .A(n9021), .B(n8809), .Z(n8810) );
  XNOR U5863 ( .A(n9200), .B(n8810), .Z(out[779]) );
  NOR U5864 ( .A(n8812), .B(n8811), .Z(n8813) );
  XNOR U5865 ( .A(n8814), .B(n8813), .Z(out[77]) );
  XNOR U5866 ( .A(in[755]), .B(n8815), .Z(n9204) );
  NAND U5867 ( .A(n9023), .B(n8816), .Z(n8817) );
  XNOR U5868 ( .A(n9204), .B(n8817), .Z(out[780]) );
  XNOR U5869 ( .A(in[756]), .B(n8818), .Z(n9208) );
  NAND U5870 ( .A(n9025), .B(n8819), .Z(n8820) );
  XNOR U5871 ( .A(n9208), .B(n8820), .Z(out[781]) );
  XNOR U5872 ( .A(in[757]), .B(n8821), .Z(n9216) );
  NAND U5873 ( .A(n9027), .B(n8822), .Z(n8823) );
  XNOR U5874 ( .A(n9216), .B(n8823), .Z(out[782]) );
  XNOR U5875 ( .A(in[758]), .B(n8824), .Z(n9220) );
  NAND U5876 ( .A(n9029), .B(n8825), .Z(n8826) );
  XNOR U5877 ( .A(n9220), .B(n8826), .Z(out[783]) );
  XNOR U5878 ( .A(in[759]), .B(n8827), .Z(n9224) );
  NAND U5879 ( .A(n9031), .B(n8828), .Z(n8829) );
  XNOR U5880 ( .A(n9224), .B(n8829), .Z(out[784]) );
  XNOR U5881 ( .A(in[760]), .B(n8830), .Z(n9228) );
  NAND U5882 ( .A(n9033), .B(n8831), .Z(n8832) );
  XNOR U5883 ( .A(n9228), .B(n8832), .Z(out[785]) );
  XNOR U5884 ( .A(in[761]), .B(n8833), .Z(n9232) );
  NAND U5885 ( .A(n9039), .B(n8834), .Z(n8835) );
  XNOR U5886 ( .A(n9232), .B(n8835), .Z(out[786]) );
  XNOR U5887 ( .A(in[762]), .B(n8836), .Z(n9236) );
  NAND U5888 ( .A(n9041), .B(n8837), .Z(n8838) );
  XNOR U5889 ( .A(n9236), .B(n8838), .Z(out[787]) );
  XNOR U5890 ( .A(in[763]), .B(n8839), .Z(n9240) );
  NAND U5891 ( .A(n9043), .B(n8840), .Z(n8841) );
  XNOR U5892 ( .A(n9240), .B(n8841), .Z(out[788]) );
  XNOR U5893 ( .A(in[764]), .B(n8842), .Z(n9244) );
  NAND U5894 ( .A(n9045), .B(n8843), .Z(n8844) );
  XNOR U5895 ( .A(n9244), .B(n8844), .Z(out[789]) );
  NOR U5896 ( .A(n8846), .B(n8845), .Z(n8847) );
  XNOR U5897 ( .A(n8848), .B(n8847), .Z(out[78]) );
  XNOR U5898 ( .A(in[765]), .B(n8849), .Z(n9248) );
  NAND U5899 ( .A(n9047), .B(n8850), .Z(n8851) );
  XNOR U5900 ( .A(n9248), .B(n8851), .Z(out[790]) );
  XNOR U5901 ( .A(in[766]), .B(n8852), .Z(n9252) );
  NAND U5902 ( .A(n9049), .B(n8853), .Z(n8854) );
  XNOR U5903 ( .A(n9252), .B(n8854), .Z(out[791]) );
  XNOR U5904 ( .A(in[767]), .B(n8855), .Z(n9260) );
  NAND U5905 ( .A(n9051), .B(n8856), .Z(n8857) );
  XNOR U5906 ( .A(n9260), .B(n8857), .Z(out[792]) );
  XNOR U5907 ( .A(in[704]), .B(n8858), .Z(n9264) );
  NAND U5908 ( .A(n9053), .B(n8859), .Z(n8860) );
  XNOR U5909 ( .A(n9264), .B(n8860), .Z(out[793]) );
  XNOR U5910 ( .A(in[705]), .B(n8861), .Z(n9268) );
  NAND U5911 ( .A(n9055), .B(n8862), .Z(n8863) );
  XNOR U5912 ( .A(n9268), .B(n8863), .Z(out[794]) );
  XNOR U5913 ( .A(in[706]), .B(n8864), .Z(n9272) );
  NAND U5914 ( .A(n9057), .B(n8865), .Z(n8866) );
  XNOR U5915 ( .A(n9272), .B(n8866), .Z(out[795]) );
  XNOR U5916 ( .A(in[707]), .B(n8867), .Z(n9276) );
  NAND U5917 ( .A(n9063), .B(n8868), .Z(n8869) );
  XNOR U5918 ( .A(n9276), .B(n8869), .Z(out[796]) );
  XNOR U5919 ( .A(in[708]), .B(n8870), .Z(n9280) );
  NAND U5920 ( .A(n9065), .B(n8871), .Z(n8872) );
  XNOR U5921 ( .A(n9280), .B(n8872), .Z(out[797]) );
  XNOR U5922 ( .A(in[709]), .B(n8873), .Z(n9284) );
  NAND U5923 ( .A(n9067), .B(n8874), .Z(n8875) );
  XNOR U5924 ( .A(n9284), .B(n8875), .Z(out[798]) );
  XNOR U5925 ( .A(in[710]), .B(n8876), .Z(n9288) );
  NAND U5926 ( .A(n9069), .B(n8877), .Z(n8878) );
  XNOR U5927 ( .A(n9288), .B(n8878), .Z(out[799]) );
  NOR U5928 ( .A(n8880), .B(n8879), .Z(n8881) );
  XNOR U5929 ( .A(n8882), .B(n8881), .Z(out[79]) );
  OR U5930 ( .A(n8884), .B(n8883), .Z(n8885) );
  XNOR U5931 ( .A(n8886), .B(n8885), .Z(out[7]) );
  XNOR U5932 ( .A(in[711]), .B(n8887), .Z(n9292) );
  NAND U5933 ( .A(n9071), .B(n8888), .Z(n8889) );
  XNOR U5934 ( .A(n9292), .B(n8889), .Z(out[800]) );
  XNOR U5935 ( .A(in[712]), .B(n8890), .Z(n9296) );
  NAND U5936 ( .A(n9073), .B(n8891), .Z(n8892) );
  XNOR U5937 ( .A(n9296), .B(n8892), .Z(out[801]) );
  XNOR U5938 ( .A(in[713]), .B(n8893), .Z(n9304) );
  NAND U5939 ( .A(n9075), .B(n8894), .Z(n8895) );
  XNOR U5940 ( .A(n9304), .B(n8895), .Z(out[802]) );
  XNOR U5941 ( .A(in[714]), .B(n8896), .Z(n9308) );
  NAND U5942 ( .A(n9077), .B(n8897), .Z(n8898) );
  XNOR U5943 ( .A(n9308), .B(n8898), .Z(out[803]) );
  XNOR U5944 ( .A(in[715]), .B(n8899), .Z(n9312) );
  NAND U5945 ( .A(n9079), .B(n8900), .Z(n8901) );
  XNOR U5946 ( .A(n9312), .B(n8901), .Z(out[804]) );
  XOR U5947 ( .A(n8902), .B(in[716]), .Z(n9316) );
  NAND U5948 ( .A(n9081), .B(n8903), .Z(n8904) );
  XNOR U5949 ( .A(n9316), .B(n8904), .Z(out[805]) );
  XOR U5950 ( .A(n8905), .B(in[717]), .Z(n9320) );
  NAND U5951 ( .A(n9087), .B(n8906), .Z(n8907) );
  XNOR U5952 ( .A(n9320), .B(n8907), .Z(out[806]) );
  XOR U5953 ( .A(n8908), .B(in[718]), .Z(n9324) );
  NAND U5954 ( .A(n9089), .B(n8909), .Z(n8910) );
  XNOR U5955 ( .A(n9324), .B(n8910), .Z(out[807]) );
  XOR U5956 ( .A(n8911), .B(in[719]), .Z(n9328) );
  NAND U5957 ( .A(n9091), .B(n8912), .Z(n8913) );
  XNOR U5958 ( .A(n9328), .B(n8913), .Z(out[808]) );
  XOR U5959 ( .A(n8914), .B(in[720]), .Z(n9332) );
  NAND U5960 ( .A(n9093), .B(n8915), .Z(n8916) );
  XNOR U5961 ( .A(n9332), .B(n8916), .Z(out[809]) );
  NOR U5962 ( .A(n8918), .B(n8917), .Z(n8919) );
  XNOR U5963 ( .A(n8920), .B(n8919), .Z(out[80]) );
  XOR U5964 ( .A(n8921), .B(in[721]), .Z(n9336) );
  NAND U5965 ( .A(n9095), .B(n8922), .Z(n8923) );
  XNOR U5966 ( .A(n9336), .B(n8923), .Z(out[810]) );
  XOR U5967 ( .A(n8924), .B(in[722]), .Z(n9340) );
  NAND U5968 ( .A(n9097), .B(n8925), .Z(n8926) );
  XNOR U5969 ( .A(n9340), .B(n8926), .Z(out[811]) );
  XOR U5970 ( .A(n8927), .B(in[723]), .Z(n9348) );
  NAND U5971 ( .A(n9099), .B(n8928), .Z(n8929) );
  XNOR U5972 ( .A(n9348), .B(n8929), .Z(out[812]) );
  XOR U5973 ( .A(in[724]), .B(n8930), .Z(n9352) );
  NAND U5974 ( .A(n9101), .B(n8931), .Z(n8932) );
  XNOR U5975 ( .A(n9352), .B(n8932), .Z(out[813]) );
  XOR U5976 ( .A(in[725]), .B(n8933), .Z(n9356) );
  NAND U5977 ( .A(n9103), .B(n8934), .Z(n8935) );
  XNOR U5978 ( .A(n9356), .B(n8935), .Z(out[814]) );
  XOR U5979 ( .A(in[726]), .B(n8936), .Z(n9360) );
  NAND U5980 ( .A(n9105), .B(n8937), .Z(n8938) );
  XNOR U5981 ( .A(n9360), .B(n8938), .Z(out[815]) );
  XOR U5982 ( .A(in[727]), .B(n8939), .Z(n9364) );
  NAND U5983 ( .A(n9111), .B(n8940), .Z(n8941) );
  XNOR U5984 ( .A(n9364), .B(n8941), .Z(out[816]) );
  XOR U5985 ( .A(in[728]), .B(n8942), .Z(n9368) );
  NAND U5986 ( .A(n9113), .B(n8943), .Z(n8944) );
  XNOR U5987 ( .A(n9368), .B(n8944), .Z(out[817]) );
  XOR U5988 ( .A(in[729]), .B(n8945), .Z(n9372) );
  NAND U5989 ( .A(n9115), .B(n8946), .Z(n8947) );
  XNOR U5990 ( .A(n9372), .B(n8947), .Z(out[818]) );
  XOR U5991 ( .A(in[730]), .B(n8948), .Z(n9376) );
  NAND U5992 ( .A(n9117), .B(n8949), .Z(n8950) );
  XNOR U5993 ( .A(n9376), .B(n8950), .Z(out[819]) );
  NOR U5994 ( .A(n8952), .B(n8951), .Z(n8953) );
  XNOR U5995 ( .A(n8954), .B(n8953), .Z(out[81]) );
  XOR U5996 ( .A(in[731]), .B(n8955), .Z(n9380) );
  NAND U5997 ( .A(n9119), .B(n8956), .Z(n8957) );
  XNOR U5998 ( .A(n9380), .B(n8957), .Z(out[820]) );
  XOR U5999 ( .A(in[732]), .B(n8958), .Z(n9384) );
  NAND U6000 ( .A(n9121), .B(n8959), .Z(n8960) );
  XNOR U6001 ( .A(n9384), .B(n8960), .Z(out[821]) );
  XOR U6002 ( .A(in[733]), .B(n8961), .Z(n9392) );
  NAND U6003 ( .A(n9123), .B(n8962), .Z(n8963) );
  XNOR U6004 ( .A(n9392), .B(n8963), .Z(out[822]) );
  XOR U6005 ( .A(in[734]), .B(n8964), .Z(n9396) );
  NAND U6006 ( .A(n9125), .B(n8965), .Z(n8966) );
  XNOR U6007 ( .A(n9396), .B(n8966), .Z(out[823]) );
  XOR U6008 ( .A(in[735]), .B(n8967), .Z(n9400) );
  NAND U6009 ( .A(n9127), .B(n8968), .Z(n8969) );
  XNOR U6010 ( .A(n9400), .B(n8969), .Z(out[824]) );
  XOR U6011 ( .A(in[736]), .B(n8970), .Z(n9404) );
  NAND U6012 ( .A(n9129), .B(n8971), .Z(n8972) );
  XNOR U6013 ( .A(n9404), .B(n8972), .Z(out[825]) );
  XOR U6014 ( .A(in[737]), .B(n8973), .Z(n9408) );
  NAND U6015 ( .A(n9135), .B(n8974), .Z(n8975) );
  XNOR U6016 ( .A(n9408), .B(n8975), .Z(out[826]) );
  XOR U6017 ( .A(in[738]), .B(n8976), .Z(n9412) );
  NAND U6018 ( .A(n9137), .B(n8977), .Z(n8978) );
  XNOR U6019 ( .A(n9412), .B(n8978), .Z(out[827]) );
  XOR U6020 ( .A(in[739]), .B(n8979), .Z(n9416) );
  NAND U6021 ( .A(n9139), .B(n8980), .Z(n8981) );
  XNOR U6022 ( .A(n9416), .B(n8981), .Z(out[828]) );
  XNOR U6023 ( .A(in[740]), .B(n8982), .Z(n9420) );
  NAND U6024 ( .A(n9141), .B(n8983), .Z(n8984) );
  XNOR U6025 ( .A(n9420), .B(n8984), .Z(out[829]) );
  NOR U6026 ( .A(n8986), .B(n8985), .Z(n8987) );
  XNOR U6027 ( .A(n8988), .B(n8987), .Z(out[82]) );
  XNOR U6028 ( .A(in[741]), .B(n8989), .Z(n9424) );
  NAND U6029 ( .A(n9143), .B(n8990), .Z(n8991) );
  XNOR U6030 ( .A(n9424), .B(n8991), .Z(out[830]) );
  XNOR U6031 ( .A(in[742]), .B(n8992), .Z(n9428) );
  NAND U6032 ( .A(n9145), .B(n8993), .Z(n8994) );
  XNOR U6033 ( .A(n9428), .B(n8994), .Z(out[831]) );
  OR U6034 ( .A(n9148), .B(n8995), .Z(n8996) );
  XNOR U6035 ( .A(n9147), .B(n8996), .Z(out[832]) );
  OR U6036 ( .A(n9152), .B(n8997), .Z(n8998) );
  XNOR U6037 ( .A(n9151), .B(n8998), .Z(out[833]) );
  OR U6038 ( .A(n9156), .B(n8999), .Z(n9000) );
  XNOR U6039 ( .A(n9155), .B(n9000), .Z(out[834]) );
  OR U6040 ( .A(n9160), .B(n9001), .Z(n9002) );
  XNOR U6041 ( .A(n9159), .B(n9002), .Z(out[835]) );
  OR U6042 ( .A(n9172), .B(n9003), .Z(n9004) );
  XNOR U6043 ( .A(n9171), .B(n9004), .Z(out[836]) );
  OR U6044 ( .A(n9176), .B(n9005), .Z(n9006) );
  XNOR U6045 ( .A(n9175), .B(n9006), .Z(out[837]) );
  OR U6046 ( .A(n9180), .B(n9007), .Z(n9008) );
  XNOR U6047 ( .A(n9179), .B(n9008), .Z(out[838]) );
  OR U6048 ( .A(n9184), .B(n9009), .Z(n9010) );
  XNOR U6049 ( .A(n9183), .B(n9010), .Z(out[839]) );
  NOR U6050 ( .A(n9012), .B(n9011), .Z(n9013) );
  XNOR U6051 ( .A(n9014), .B(n9013), .Z(out[83]) );
  OR U6052 ( .A(n9188), .B(n9015), .Z(n9016) );
  XNOR U6053 ( .A(n9187), .B(n9016), .Z(out[840]) );
  OR U6054 ( .A(n9192), .B(n9017), .Z(n9018) );
  XNOR U6055 ( .A(n9191), .B(n9018), .Z(out[841]) );
  OR U6056 ( .A(n9196), .B(n9019), .Z(n9020) );
  XNOR U6057 ( .A(n9195), .B(n9020), .Z(out[842]) );
  OR U6058 ( .A(n9200), .B(n9021), .Z(n9022) );
  XNOR U6059 ( .A(n9199), .B(n9022), .Z(out[843]) );
  OR U6060 ( .A(n9204), .B(n9023), .Z(n9024) );
  XNOR U6061 ( .A(n9203), .B(n9024), .Z(out[844]) );
  OR U6062 ( .A(n9208), .B(n9025), .Z(n9026) );
  XNOR U6063 ( .A(n9207), .B(n9026), .Z(out[845]) );
  OR U6064 ( .A(n9216), .B(n9027), .Z(n9028) );
  XNOR U6065 ( .A(n9215), .B(n9028), .Z(out[846]) );
  OR U6066 ( .A(n9220), .B(n9029), .Z(n9030) );
  XNOR U6067 ( .A(n9219), .B(n9030), .Z(out[847]) );
  OR U6068 ( .A(n9224), .B(n9031), .Z(n9032) );
  XNOR U6069 ( .A(n9223), .B(n9032), .Z(out[848]) );
  OR U6070 ( .A(n9228), .B(n9033), .Z(n9034) );
  XNOR U6071 ( .A(n9227), .B(n9034), .Z(out[849]) );
  NOR U6072 ( .A(n9036), .B(n9035), .Z(n9037) );
  XNOR U6073 ( .A(n9038), .B(n9037), .Z(out[84]) );
  OR U6074 ( .A(n9232), .B(n9039), .Z(n9040) );
  XNOR U6075 ( .A(n9231), .B(n9040), .Z(out[850]) );
  OR U6076 ( .A(n9236), .B(n9041), .Z(n9042) );
  XNOR U6077 ( .A(n9235), .B(n9042), .Z(out[851]) );
  OR U6078 ( .A(n9240), .B(n9043), .Z(n9044) );
  XNOR U6079 ( .A(n9239), .B(n9044), .Z(out[852]) );
  OR U6080 ( .A(n9244), .B(n9045), .Z(n9046) );
  XNOR U6081 ( .A(n9243), .B(n9046), .Z(out[853]) );
  OR U6082 ( .A(n9248), .B(n9047), .Z(n9048) );
  XNOR U6083 ( .A(n9247), .B(n9048), .Z(out[854]) );
  OR U6084 ( .A(n9252), .B(n9049), .Z(n9050) );
  XNOR U6085 ( .A(n9251), .B(n9050), .Z(out[855]) );
  OR U6086 ( .A(n9260), .B(n9051), .Z(n9052) );
  XNOR U6087 ( .A(n9259), .B(n9052), .Z(out[856]) );
  OR U6088 ( .A(n9264), .B(n9053), .Z(n9054) );
  XNOR U6089 ( .A(n9263), .B(n9054), .Z(out[857]) );
  OR U6090 ( .A(n9268), .B(n9055), .Z(n9056) );
  XNOR U6091 ( .A(n9267), .B(n9056), .Z(out[858]) );
  OR U6092 ( .A(n9272), .B(n9057), .Z(n9058) );
  XNOR U6093 ( .A(n9271), .B(n9058), .Z(out[859]) );
  NOR U6094 ( .A(n9060), .B(n9059), .Z(n9061) );
  XNOR U6095 ( .A(n9062), .B(n9061), .Z(out[85]) );
  OR U6096 ( .A(n9276), .B(n9063), .Z(n9064) );
  XNOR U6097 ( .A(n9275), .B(n9064), .Z(out[860]) );
  OR U6098 ( .A(n9280), .B(n9065), .Z(n9066) );
  XNOR U6099 ( .A(n9279), .B(n9066), .Z(out[861]) );
  OR U6100 ( .A(n9284), .B(n9067), .Z(n9068) );
  XNOR U6101 ( .A(n9283), .B(n9068), .Z(out[862]) );
  OR U6102 ( .A(n9288), .B(n9069), .Z(n9070) );
  XNOR U6103 ( .A(n9287), .B(n9070), .Z(out[863]) );
  OR U6104 ( .A(n9292), .B(n9071), .Z(n9072) );
  XNOR U6105 ( .A(n9291), .B(n9072), .Z(out[864]) );
  OR U6106 ( .A(n9296), .B(n9073), .Z(n9074) );
  XNOR U6107 ( .A(n9295), .B(n9074), .Z(out[865]) );
  OR U6108 ( .A(n9304), .B(n9075), .Z(n9076) );
  XNOR U6109 ( .A(n9303), .B(n9076), .Z(out[866]) );
  OR U6110 ( .A(n9308), .B(n9077), .Z(n9078) );
  XNOR U6111 ( .A(n9307), .B(n9078), .Z(out[867]) );
  OR U6112 ( .A(n9312), .B(n9079), .Z(n9080) );
  XNOR U6113 ( .A(n9311), .B(n9080), .Z(out[868]) );
  OR U6114 ( .A(n9316), .B(n9081), .Z(n9082) );
  XNOR U6115 ( .A(n9315), .B(n9082), .Z(out[869]) );
  NOR U6116 ( .A(n9084), .B(n9083), .Z(n9085) );
  XNOR U6117 ( .A(n9086), .B(n9085), .Z(out[86]) );
  OR U6118 ( .A(n9320), .B(n9087), .Z(n9088) );
  XNOR U6119 ( .A(n9319), .B(n9088), .Z(out[870]) );
  OR U6120 ( .A(n9324), .B(n9089), .Z(n9090) );
  XNOR U6121 ( .A(n9323), .B(n9090), .Z(out[871]) );
  OR U6122 ( .A(n9328), .B(n9091), .Z(n9092) );
  XNOR U6123 ( .A(n9327), .B(n9092), .Z(out[872]) );
  OR U6124 ( .A(n9332), .B(n9093), .Z(n9094) );
  XNOR U6125 ( .A(n9331), .B(n9094), .Z(out[873]) );
  OR U6126 ( .A(n9336), .B(n9095), .Z(n9096) );
  XNOR U6127 ( .A(n9335), .B(n9096), .Z(out[874]) );
  OR U6128 ( .A(n9340), .B(n9097), .Z(n9098) );
  XNOR U6129 ( .A(n9339), .B(n9098), .Z(out[875]) );
  OR U6130 ( .A(n9348), .B(n9099), .Z(n9100) );
  XNOR U6131 ( .A(n9347), .B(n9100), .Z(out[876]) );
  OR U6132 ( .A(n9352), .B(n9101), .Z(n9102) );
  XNOR U6133 ( .A(n9351), .B(n9102), .Z(out[877]) );
  OR U6134 ( .A(n9356), .B(n9103), .Z(n9104) );
  XNOR U6135 ( .A(n9355), .B(n9104), .Z(out[878]) );
  OR U6136 ( .A(n9360), .B(n9105), .Z(n9106) );
  XNOR U6137 ( .A(n9359), .B(n9106), .Z(out[879]) );
  NOR U6138 ( .A(n9108), .B(n9107), .Z(n9109) );
  XNOR U6139 ( .A(n9110), .B(n9109), .Z(out[87]) );
  OR U6140 ( .A(n9364), .B(n9111), .Z(n9112) );
  XNOR U6141 ( .A(n9363), .B(n9112), .Z(out[880]) );
  OR U6142 ( .A(n9368), .B(n9113), .Z(n9114) );
  XNOR U6143 ( .A(n9367), .B(n9114), .Z(out[881]) );
  OR U6144 ( .A(n9372), .B(n9115), .Z(n9116) );
  XNOR U6145 ( .A(n9371), .B(n9116), .Z(out[882]) );
  OR U6146 ( .A(n9376), .B(n9117), .Z(n9118) );
  XNOR U6147 ( .A(n9375), .B(n9118), .Z(out[883]) );
  OR U6148 ( .A(n9380), .B(n9119), .Z(n9120) );
  XNOR U6149 ( .A(n9379), .B(n9120), .Z(out[884]) );
  OR U6150 ( .A(n9384), .B(n9121), .Z(n9122) );
  XNOR U6151 ( .A(n9383), .B(n9122), .Z(out[885]) );
  OR U6152 ( .A(n9392), .B(n9123), .Z(n9124) );
  XNOR U6153 ( .A(n9391), .B(n9124), .Z(out[886]) );
  OR U6154 ( .A(n9396), .B(n9125), .Z(n9126) );
  XNOR U6155 ( .A(n9395), .B(n9126), .Z(out[887]) );
  OR U6156 ( .A(n9400), .B(n9127), .Z(n9128) );
  XNOR U6157 ( .A(n9399), .B(n9128), .Z(out[888]) );
  OR U6158 ( .A(n9404), .B(n9129), .Z(n9130) );
  XNOR U6159 ( .A(n9403), .B(n9130), .Z(out[889]) );
  NOR U6160 ( .A(n9132), .B(n9131), .Z(n9133) );
  XNOR U6161 ( .A(n9134), .B(n9133), .Z(out[88]) );
  OR U6162 ( .A(n9408), .B(n9135), .Z(n9136) );
  XNOR U6163 ( .A(n9407), .B(n9136), .Z(out[890]) );
  OR U6164 ( .A(n9412), .B(n9137), .Z(n9138) );
  XNOR U6165 ( .A(n9411), .B(n9138), .Z(out[891]) );
  OR U6166 ( .A(n9416), .B(n9139), .Z(n9140) );
  XNOR U6167 ( .A(n9415), .B(n9140), .Z(out[892]) );
  OR U6168 ( .A(n9420), .B(n9141), .Z(n9142) );
  XNOR U6169 ( .A(n9419), .B(n9142), .Z(out[893]) );
  OR U6170 ( .A(n9424), .B(n9143), .Z(n9144) );
  XNOR U6171 ( .A(n9423), .B(n9144), .Z(out[894]) );
  OR U6172 ( .A(n9428), .B(n9145), .Z(n9146) );
  XNOR U6173 ( .A(n9427), .B(n9146), .Z(out[895]) );
  ANDN U6174 ( .B(n9148), .A(n9147), .Z(n9149) );
  XNOR U6175 ( .A(n9150), .B(n9149), .Z(out[896]) );
  ANDN U6176 ( .B(n9152), .A(n9151), .Z(n9153) );
  XNOR U6177 ( .A(n9154), .B(n9153), .Z(out[897]) );
  ANDN U6178 ( .B(n9156), .A(n9155), .Z(n9157) );
  XNOR U6179 ( .A(n9158), .B(n9157), .Z(out[898]) );
  ANDN U6180 ( .B(n9160), .A(n9159), .Z(n9161) );
  XNOR U6181 ( .A(n9162), .B(n9161), .Z(out[899]) );
  NOR U6182 ( .A(n9164), .B(n9163), .Z(n9165) );
  XNOR U6183 ( .A(n9166), .B(n9165), .Z(out[89]) );
  OR U6184 ( .A(n9168), .B(n9167), .Z(n9169) );
  XNOR U6185 ( .A(n9170), .B(n9169), .Z(out[8]) );
  ANDN U6186 ( .B(n9172), .A(n9171), .Z(n9173) );
  XNOR U6187 ( .A(n9174), .B(n9173), .Z(out[900]) );
  ANDN U6188 ( .B(n9176), .A(n9175), .Z(n9177) );
  XNOR U6189 ( .A(n9178), .B(n9177), .Z(out[901]) );
  ANDN U6190 ( .B(n9180), .A(n9179), .Z(n9181) );
  XNOR U6191 ( .A(n9182), .B(n9181), .Z(out[902]) );
  ANDN U6192 ( .B(n9184), .A(n9183), .Z(n9185) );
  XNOR U6193 ( .A(n9186), .B(n9185), .Z(out[903]) );
  ANDN U6194 ( .B(n9188), .A(n9187), .Z(n9189) );
  XNOR U6195 ( .A(n9190), .B(n9189), .Z(out[904]) );
  ANDN U6196 ( .B(n9192), .A(n9191), .Z(n9193) );
  XNOR U6197 ( .A(n9194), .B(n9193), .Z(out[905]) );
  ANDN U6198 ( .B(n9196), .A(n9195), .Z(n9197) );
  XNOR U6199 ( .A(n9198), .B(n9197), .Z(out[906]) );
  ANDN U6200 ( .B(n9200), .A(n9199), .Z(n9201) );
  XNOR U6201 ( .A(n9202), .B(n9201), .Z(out[907]) );
  ANDN U6202 ( .B(n9204), .A(n9203), .Z(n9205) );
  XNOR U6203 ( .A(n9206), .B(n9205), .Z(out[908]) );
  ANDN U6204 ( .B(n9208), .A(n9207), .Z(n9209) );
  XNOR U6205 ( .A(n9210), .B(n9209), .Z(out[909]) );
  NOR U6206 ( .A(n9212), .B(n9211), .Z(n9213) );
  XNOR U6207 ( .A(n9214), .B(n9213), .Z(out[90]) );
  ANDN U6208 ( .B(n9216), .A(n9215), .Z(n9217) );
  XNOR U6209 ( .A(n9218), .B(n9217), .Z(out[910]) );
  ANDN U6210 ( .B(n9220), .A(n9219), .Z(n9221) );
  XNOR U6211 ( .A(n9222), .B(n9221), .Z(out[911]) );
  ANDN U6212 ( .B(n9224), .A(n9223), .Z(n9225) );
  XNOR U6213 ( .A(n9226), .B(n9225), .Z(out[912]) );
  ANDN U6214 ( .B(n9228), .A(n9227), .Z(n9229) );
  XNOR U6215 ( .A(n9230), .B(n9229), .Z(out[913]) );
  ANDN U6216 ( .B(n9232), .A(n9231), .Z(n9233) );
  XNOR U6217 ( .A(n9234), .B(n9233), .Z(out[914]) );
  ANDN U6218 ( .B(n9236), .A(n9235), .Z(n9237) );
  XNOR U6219 ( .A(n9238), .B(n9237), .Z(out[915]) );
  ANDN U6220 ( .B(n9240), .A(n9239), .Z(n9241) );
  XNOR U6221 ( .A(n9242), .B(n9241), .Z(out[916]) );
  ANDN U6222 ( .B(n9244), .A(n9243), .Z(n9245) );
  XNOR U6223 ( .A(n9246), .B(n9245), .Z(out[917]) );
  ANDN U6224 ( .B(n9248), .A(n9247), .Z(n9249) );
  XNOR U6225 ( .A(n9250), .B(n9249), .Z(out[918]) );
  ANDN U6226 ( .B(n9252), .A(n9251), .Z(n9253) );
  XNOR U6227 ( .A(n9254), .B(n9253), .Z(out[919]) );
  NOR U6228 ( .A(n9256), .B(n9255), .Z(n9257) );
  XNOR U6229 ( .A(n9258), .B(n9257), .Z(out[91]) );
  ANDN U6230 ( .B(n9260), .A(n9259), .Z(n9261) );
  XNOR U6231 ( .A(n9262), .B(n9261), .Z(out[920]) );
  ANDN U6232 ( .B(n9264), .A(n9263), .Z(n9265) );
  XNOR U6233 ( .A(n9266), .B(n9265), .Z(out[921]) );
  ANDN U6234 ( .B(n9268), .A(n9267), .Z(n9269) );
  XNOR U6235 ( .A(n9270), .B(n9269), .Z(out[922]) );
  ANDN U6236 ( .B(n9272), .A(n9271), .Z(n9273) );
  XNOR U6237 ( .A(n9274), .B(n9273), .Z(out[923]) );
  ANDN U6238 ( .B(n9276), .A(n9275), .Z(n9277) );
  XNOR U6239 ( .A(n9278), .B(n9277), .Z(out[924]) );
  ANDN U6240 ( .B(n9280), .A(n9279), .Z(n9281) );
  XNOR U6241 ( .A(n9282), .B(n9281), .Z(out[925]) );
  ANDN U6242 ( .B(n9284), .A(n9283), .Z(n9285) );
  XNOR U6243 ( .A(n9286), .B(n9285), .Z(out[926]) );
  ANDN U6244 ( .B(n9288), .A(n9287), .Z(n9289) );
  XNOR U6245 ( .A(n9290), .B(n9289), .Z(out[927]) );
  ANDN U6246 ( .B(n9292), .A(n9291), .Z(n9293) );
  XNOR U6247 ( .A(n9294), .B(n9293), .Z(out[928]) );
  ANDN U6248 ( .B(n9296), .A(n9295), .Z(n9297) );
  XNOR U6249 ( .A(n9298), .B(n9297), .Z(out[929]) );
  ANDN U6250 ( .B(n9300), .A(n9299), .Z(n9301) );
  XNOR U6251 ( .A(n9302), .B(n9301), .Z(out[92]) );
  ANDN U6252 ( .B(n9304), .A(n9303), .Z(n9305) );
  XNOR U6253 ( .A(n9306), .B(n9305), .Z(out[930]) );
  ANDN U6254 ( .B(n9308), .A(n9307), .Z(n9309) );
  XNOR U6255 ( .A(n9310), .B(n9309), .Z(out[931]) );
  ANDN U6256 ( .B(n9312), .A(n9311), .Z(n9313) );
  XNOR U6257 ( .A(n9314), .B(n9313), .Z(out[932]) );
  ANDN U6258 ( .B(n9316), .A(n9315), .Z(n9317) );
  XNOR U6259 ( .A(n9318), .B(n9317), .Z(out[933]) );
  ANDN U6260 ( .B(n9320), .A(n9319), .Z(n9321) );
  XNOR U6261 ( .A(n9322), .B(n9321), .Z(out[934]) );
  ANDN U6262 ( .B(n9324), .A(n9323), .Z(n9325) );
  XNOR U6263 ( .A(n9326), .B(n9325), .Z(out[935]) );
  ANDN U6264 ( .B(n9328), .A(n9327), .Z(n9329) );
  XNOR U6265 ( .A(n9330), .B(n9329), .Z(out[936]) );
  ANDN U6266 ( .B(n9332), .A(n9331), .Z(n9333) );
  XNOR U6267 ( .A(n9334), .B(n9333), .Z(out[937]) );
  ANDN U6268 ( .B(n9336), .A(n9335), .Z(n9337) );
  XNOR U6269 ( .A(n9338), .B(n9337), .Z(out[938]) );
  ANDN U6270 ( .B(n9340), .A(n9339), .Z(n9341) );
  XNOR U6271 ( .A(n9342), .B(n9341), .Z(out[939]) );
  ANDN U6272 ( .B(n9344), .A(n9343), .Z(n9345) );
  XNOR U6273 ( .A(n9346), .B(n9345), .Z(out[93]) );
  ANDN U6274 ( .B(n9348), .A(n9347), .Z(n9349) );
  XNOR U6275 ( .A(n9350), .B(n9349), .Z(out[940]) );
  ANDN U6276 ( .B(n9352), .A(n9351), .Z(n9353) );
  XNOR U6277 ( .A(n9354), .B(n9353), .Z(out[941]) );
  ANDN U6278 ( .B(n9356), .A(n9355), .Z(n9357) );
  XNOR U6279 ( .A(n9358), .B(n9357), .Z(out[942]) );
  ANDN U6280 ( .B(n9360), .A(n9359), .Z(n9361) );
  XNOR U6281 ( .A(n9362), .B(n9361), .Z(out[943]) );
  ANDN U6282 ( .B(n9364), .A(n9363), .Z(n9365) );
  XNOR U6283 ( .A(n9366), .B(n9365), .Z(out[944]) );
  ANDN U6284 ( .B(n9368), .A(n9367), .Z(n9369) );
  XNOR U6285 ( .A(n9370), .B(n9369), .Z(out[945]) );
  ANDN U6286 ( .B(n9372), .A(n9371), .Z(n9373) );
  XNOR U6287 ( .A(n9374), .B(n9373), .Z(out[946]) );
  ANDN U6288 ( .B(n9376), .A(n9375), .Z(n9377) );
  XNOR U6289 ( .A(n9378), .B(n9377), .Z(out[947]) );
  ANDN U6290 ( .B(n9380), .A(n9379), .Z(n9381) );
  XNOR U6291 ( .A(n9382), .B(n9381), .Z(out[948]) );
  ANDN U6292 ( .B(n9384), .A(n9383), .Z(n9385) );
  XNOR U6293 ( .A(n9386), .B(n9385), .Z(out[949]) );
  ANDN U6294 ( .B(n9388), .A(n9387), .Z(n9389) );
  XNOR U6295 ( .A(n9390), .B(n9389), .Z(out[94]) );
  ANDN U6296 ( .B(n9392), .A(n9391), .Z(n9393) );
  XNOR U6297 ( .A(n9394), .B(n9393), .Z(out[950]) );
  ANDN U6298 ( .B(n9396), .A(n9395), .Z(n9397) );
  XNOR U6299 ( .A(n9398), .B(n9397), .Z(out[951]) );
  ANDN U6300 ( .B(n9400), .A(n9399), .Z(n9401) );
  XNOR U6301 ( .A(n9402), .B(n9401), .Z(out[952]) );
  ANDN U6302 ( .B(n9404), .A(n9403), .Z(n9405) );
  XNOR U6303 ( .A(n9406), .B(n9405), .Z(out[953]) );
  ANDN U6304 ( .B(n9408), .A(n9407), .Z(n9409) );
  XNOR U6305 ( .A(n9410), .B(n9409), .Z(out[954]) );
  ANDN U6306 ( .B(n9412), .A(n9411), .Z(n9413) );
  XNOR U6307 ( .A(n9414), .B(n9413), .Z(out[955]) );
  ANDN U6308 ( .B(n9416), .A(n9415), .Z(n9417) );
  XNOR U6309 ( .A(n9418), .B(n9417), .Z(out[956]) );
  ANDN U6310 ( .B(n9420), .A(n9419), .Z(n9421) );
  XNOR U6311 ( .A(n9422), .B(n9421), .Z(out[957]) );
  ANDN U6312 ( .B(n9424), .A(n9423), .Z(n9425) );
  XNOR U6313 ( .A(n9426), .B(n9425), .Z(out[958]) );
  ANDN U6314 ( .B(n9428), .A(n9427), .Z(n9429) );
  XNOR U6315 ( .A(n9430), .B(n9429), .Z(out[959]) );
  ANDN U6316 ( .B(n9432), .A(n9431), .Z(n9433) );
  XNOR U6317 ( .A(n9434), .B(n9433), .Z(out[95]) );
  ANDN U6318 ( .B(n9436), .A(n9435), .Z(n9437) );
  XNOR U6319 ( .A(n9438), .B(n9437), .Z(out[960]) );
  ANDN U6320 ( .B(n9440), .A(n9439), .Z(n9441) );
  XNOR U6321 ( .A(n9442), .B(n9441), .Z(out[961]) );
  ANDN U6322 ( .B(n9444), .A(n9443), .Z(n9445) );
  XNOR U6323 ( .A(n9446), .B(n9445), .Z(out[962]) );
  ANDN U6324 ( .B(n9448), .A(n9447), .Z(n9449) );
  XNOR U6325 ( .A(n9450), .B(n9449), .Z(out[963]) );
  ANDN U6326 ( .B(n9452), .A(n9451), .Z(n9453) );
  XNOR U6327 ( .A(n9454), .B(n9453), .Z(out[964]) );
  ANDN U6328 ( .B(n9456), .A(n9455), .Z(n9457) );
  XNOR U6329 ( .A(n9458), .B(n9457), .Z(out[965]) );
  ANDN U6330 ( .B(n9460), .A(n9459), .Z(n9461) );
  XNOR U6331 ( .A(n9462), .B(n9461), .Z(out[966]) );
  ANDN U6332 ( .B(n9464), .A(n9463), .Z(n9465) );
  XNOR U6333 ( .A(n9466), .B(n9465), .Z(out[967]) );
  ANDN U6334 ( .B(n9468), .A(n9467), .Z(n9469) );
  XNOR U6335 ( .A(n9470), .B(n9469), .Z(out[968]) );
  ANDN U6336 ( .B(n9472), .A(n9471), .Z(n9473) );
  XNOR U6337 ( .A(n9474), .B(n9473), .Z(out[969]) );
  ANDN U6338 ( .B(n9476), .A(n9475), .Z(n9477) );
  XNOR U6339 ( .A(n9478), .B(n9477), .Z(out[96]) );
  ANDN U6340 ( .B(n9480), .A(n9479), .Z(n9481) );
  XNOR U6341 ( .A(n9482), .B(n9481), .Z(out[970]) );
  ANDN U6342 ( .B(n9484), .A(n9483), .Z(n9485) );
  XNOR U6343 ( .A(n9486), .B(n9485), .Z(out[971]) );
  ANDN U6344 ( .B(n9488), .A(n9487), .Z(n9489) );
  XNOR U6345 ( .A(n9490), .B(n9489), .Z(out[972]) );
  ANDN U6346 ( .B(n9492), .A(n9491), .Z(n9493) );
  XNOR U6347 ( .A(n9494), .B(n9493), .Z(out[973]) );
  ANDN U6348 ( .B(n9496), .A(n9495), .Z(n9497) );
  XNOR U6349 ( .A(n9498), .B(n9497), .Z(out[974]) );
  ANDN U6350 ( .B(n9500), .A(n9499), .Z(n9501) );
  XNOR U6351 ( .A(n9502), .B(n9501), .Z(out[975]) );
  ANDN U6352 ( .B(n9504), .A(n9503), .Z(n9505) );
  XNOR U6353 ( .A(n9506), .B(n9505), .Z(out[976]) );
  ANDN U6354 ( .B(n9508), .A(n9507), .Z(n9509) );
  XNOR U6355 ( .A(n9510), .B(n9509), .Z(out[977]) );
  ANDN U6356 ( .B(n9512), .A(n9511), .Z(n9513) );
  XNOR U6357 ( .A(n9514), .B(n9513), .Z(out[978]) );
  ANDN U6358 ( .B(n9516), .A(n9515), .Z(n9517) );
  XNOR U6359 ( .A(n9518), .B(n9517), .Z(out[979]) );
  ANDN U6360 ( .B(n9520), .A(n9519), .Z(n9521) );
  XNOR U6361 ( .A(n9522), .B(n9521), .Z(out[97]) );
  ANDN U6362 ( .B(n9524), .A(n9523), .Z(n9525) );
  XNOR U6363 ( .A(n9526), .B(n9525), .Z(out[980]) );
  ANDN U6364 ( .B(n9528), .A(n9527), .Z(n9529) );
  XNOR U6365 ( .A(n9530), .B(n9529), .Z(out[981]) );
  ANDN U6366 ( .B(n9532), .A(n9531), .Z(n9533) );
  XNOR U6367 ( .A(n9534), .B(n9533), .Z(out[982]) );
  ANDN U6368 ( .B(n9536), .A(n9535), .Z(n9537) );
  XNOR U6369 ( .A(n9538), .B(n9537), .Z(out[983]) );
  ANDN U6370 ( .B(n9540), .A(n9539), .Z(n9541) );
  XNOR U6371 ( .A(n9542), .B(n9541), .Z(out[984]) );
  ANDN U6372 ( .B(n9544), .A(n9543), .Z(n9545) );
  XNOR U6373 ( .A(n9546), .B(n9545), .Z(out[985]) );
  ANDN U6374 ( .B(n9548), .A(n9547), .Z(n9549) );
  XNOR U6375 ( .A(n9550), .B(n9549), .Z(out[986]) );
  ANDN U6376 ( .B(n9552), .A(n9551), .Z(n9553) );
  XNOR U6377 ( .A(n9554), .B(n9553), .Z(out[987]) );
  ANDN U6378 ( .B(n9556), .A(n9555), .Z(n9557) );
  XNOR U6379 ( .A(n9558), .B(n9557), .Z(out[988]) );
  ANDN U6380 ( .B(n9560), .A(n9559), .Z(n9561) );
  XNOR U6381 ( .A(n9562), .B(n9561), .Z(out[989]) );
  ANDN U6382 ( .B(n9564), .A(n9563), .Z(n9565) );
  XNOR U6383 ( .A(n9566), .B(n9565), .Z(out[98]) );
  ANDN U6384 ( .B(n9568), .A(n9567), .Z(n9569) );
  XNOR U6385 ( .A(n9570), .B(n9569), .Z(out[990]) );
  ANDN U6386 ( .B(n9572), .A(n9571), .Z(n9573) );
  XNOR U6387 ( .A(n9574), .B(n9573), .Z(out[991]) );
  ANDN U6388 ( .B(n9576), .A(n9575), .Z(n9577) );
  XNOR U6389 ( .A(n9578), .B(n9577), .Z(out[992]) );
  ANDN U6390 ( .B(n9580), .A(n9579), .Z(n9581) );
  XNOR U6391 ( .A(n9582), .B(n9581), .Z(out[993]) );
  ANDN U6392 ( .B(n9584), .A(n9583), .Z(n9585) );
  XNOR U6393 ( .A(n9586), .B(n9585), .Z(out[994]) );
  ANDN U6394 ( .B(n9588), .A(n9587), .Z(n9589) );
  XNOR U6395 ( .A(n9590), .B(n9589), .Z(out[995]) );
  ANDN U6396 ( .B(n9592), .A(n9591), .Z(n9593) );
  XNOR U6397 ( .A(n9594), .B(n9593), .Z(out[996]) );
  ANDN U6398 ( .B(n9596), .A(n9595), .Z(n9597) );
  XNOR U6399 ( .A(n9598), .B(n9597), .Z(out[997]) );
  ANDN U6400 ( .B(n9600), .A(n9599), .Z(n9601) );
  XNOR U6401 ( .A(n9602), .B(n9601), .Z(out[998]) );
  ANDN U6402 ( .B(n9604), .A(n9603), .Z(n9605) );
  XNOR U6403 ( .A(n9606), .B(n9605), .Z(out[999]) );
  ANDN U6404 ( .B(n9608), .A(n9607), .Z(n9609) );
  XNOR U6405 ( .A(n9610), .B(n9609), .Z(out[99]) );
  OR U6406 ( .A(n9612), .B(n9611), .Z(n9613) );
  XNOR U6407 ( .A(n9614), .B(n9613), .Z(out[9]) );
endmodule


module sha3_seq_CC12 ( clk, rst, in, out );
  input [575:0] in;
  output [1599:0] out;
  input clk, rst;
  wire   init, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74,
         N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123,
         N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134,
         N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145,
         N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156,
         N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167,
         N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189,
         N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200,
         N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211,
         N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222,
         N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233,
         N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244,
         N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255,
         N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266,
         N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277,
         N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288,
         N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299,
         N300, N301, N302, N303, N304, N305, N306, N307, N308, N309, N310,
         N311, N312, N313, N314, N315, N316, N317, N318, N319, N320, N321,
         N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332,
         N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343,
         N344, N345, N346, N347, N348, N349, N350, N351, N352, N353, N354,
         N355, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365,
         N366, N367, N368, N369, N370, N371, N372, N373, N374, N375, N376,
         N377, N378, N379, N380, N381, N382, N383, N384, N385, N386, N387,
         N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398,
         N399, N400, N401, N402, N403, N404, N405, N406, N407, N408, N409,
         N410, N411, N412, N413, N414, N415, N416, N417, N418, N419, N420,
         N421, N422, N423, N424, N425, N426, N427, N428, N429, N430, N431,
         N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, N442,
         N443, N444, N445, N446, N447, N448, N449, N450, N451, N452, N453,
         N454, N455, N456, N457, N458, N459, N460, N461, N462, N463, N464,
         N465, N466, N467, N468, N469, N470, N471, N472, N473, N474, N475,
         N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, N486,
         N487, N488, N489, N490, N491, N492, N493, N494, N495, N496, N497,
         N498, N499, N500, N501, N502, N503, N504, N505, N506, N507, N508,
         N509, N510, N511, N512, N513, N514, N515, N516, N517, N518, N519,
         N520, N521, N522, N523, N524, N525, N526, N527, N528, N529, N530,
         N531, N532, N533, N534, N535, N536, N537, N538, N539, N540, N541,
         N542, N543, N544, N545, N546, N547, N548, N549, N550, N551, N552,
         N553, N554, N555, N556, N557, N558, N559, N560, N561, N562, N563,
         N564, N565, N566, N567, N568, N569, N570, N571, N572, N573, N574,
         N575, N576, N577, N578, N579, N580, N581, N582, N583, N584, N585,
         N586, N587, N588, N589, N590, N591, N592, N593, N594, N595, N596,
         N597, N598, N599, N600, N601, N602, N603, N604, N605, N606, N607,
         N608, N609, N610, N611, N612, N613, N614, N615, N616, N617, N618,
         N619, N620, N621, N622, N623, N624, N625, N626, N627, N628, N629,
         N630, N631, N632, N633, N634, N635, N636, N637, N638, N639, N640,
         N641, N642, N643, N644, N645, N646, N647, N648, N649, N650, N651,
         N652, N653, N654, N655, N656, N657, N658, N659, N660, N661, N662,
         N663, N664, N665, N666, N667, N668, N669, N670, N671, N672, N673,
         N674, N675, N676, N677, N678, N679, N680, N681, N682, N683, N684,
         N685, N686, N687, N688, N689, N690, N691, N692, N693, N694, N695,
         N696, N697, N698, N699, N700, N701, N702, N703, N704, N705, N706,
         N707, N708, N709, N710, N711, N712, N713, N714, N715, N716, N717,
         N718, N719, N720, N721, N722, N723, N724, N725, N726, N727, N728,
         N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739,
         N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750,
         N751, N752, N753, N754, N755, N756, N757, N758, N759, N760, N761,
         N762, N763, N764, N765, N766, N767, N768, N769, N770, N771, N772,
         N773, N774, N775, N776, N777, N778, N779, N780, N781, N782, N783,
         N784, N785, N786, N787, N788, N789, N790, N791, N792, N793, N794,
         N795, N796, N797, N798, N799, N800, N801, N802, N803, N804, N805,
         N806, N807, N808, N809, N810, N811, N812, N813, N814, N815, N816,
         N817, N818, N819, N820, N821, N822, N823, N824, N825, N826, N827,
         N828, N829, N830, N831, N832, N833, N834, N835, N836, N837, N838,
         N839, N840, N841, N842, N843, N844, N845, N846, N847, N848, N849,
         N850, N851, N852, N853, N854, N855, N856, N857, N858, N859, N860,
         N861, N862, N863, N864, N865, N866, N867, N868, N869, N870, N871,
         N872, N873, N874, N875, N876, N877, N878, N879, N880, N881, N882,
         N883, N884, N885, N886, N887, N888, N889, N890, N891, N892, N893,
         N894, N895, N896, N897, N898, N899, N900, N901, N902, N903, N904,
         N905, N906, N907, N908, N909, N910, N911, N912, N913, N914, N915,
         N916, N917, N918, N919, N920, N921, N922, N923, N924, N925, N926,
         N927, N928, N929, N930, N931, N932, N933, N934, N935, N936, N937,
         N938, N939, N940, N941, N942, N943, N944, N945, N946, N947, N948,
         N949, N950, N951, N952, N953, N954, N955, N956, N957, N958, N959,
         N960, N961, N962, N963, N964, N965, N966, N967, N968, N969, N970,
         N971, N972, N973, N974, N975, N976, N977, N978, N979, N980, N981,
         N982, N983, N984, N985, N986, N987, N988, N989, N990, N991, N992,
         N993, N994, N995, N996, N997, N998, N999, N1000, N1001, N1002, N1003,
         N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013,
         N1014, N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022, N1023,
         N1024, N1025, N1026, N1027, N1028, N1029, N1030, N1031, N1032, N1033,
         N1034, N1035, N1036, N1037, N1038, N1039, N1040, N1041, N1042, N1043,
         N1044, N1045, N1046, N1047, N1048, N1049, N1050, N1051, N1052, N1053,
         N1054, N1055, N1056, N1057, N1058, N1059, N1060, N1061, N1062, N1063,
         N1064, N1065, N1066, N1067, N1068, N1069, N1070, N1071, N1072, N1073,
         N1074, N1075, N1076, N1077, N1078, N1079, N1080, N1081, N1082, N1083,
         N1084, N1085, N1086, N1087, N1088, N1089, N1090, N1091, N1092, N1093,
         N1094, N1095, N1096, N1097, N1098, N1099, N1100, N1101, N1102, N1103,
         N1104, N1105, N1106, N1107, N1108, N1109, N1110, N1111, N1112, N1113,
         N1114, N1115, N1116, N1117, N1118, N1119, N1120, N1121, N1122, N1123,
         N1124, N1125, N1126, N1127, N1128, N1129, N1130, N1131, N1132, N1133,
         N1134, N1135, N1136, N1137, N1138, N1139, N1140, N1141, N1142, N1143,
         N1144, N1145, N1146, N1147, N1148, N1149, N1150, N1151, N1152, N1153,
         N1154, N1155, N1156, N1157, N1158, N1159, N1160, N1161, N1162, N1163,
         N1164, N1165, N1166, N1167, N1168, N1169, N1170, N1171, N1172, N1173,
         N1174, N1175, N1176, N1177, N1178, N1179, N1180, N1181, N1182, N1183,
         N1184, N1185, N1186, N1187, N1188, N1189, N1190, N1191, N1192, N1193,
         N1194, N1195, N1196, N1197, N1198, N1199, N1200, N1201, N1202, N1203,
         N1204, N1205, N1206, N1207, N1208, N1209, N1210, N1211, N1212, N1213,
         N1214, N1215, N1216, N1217, N1218, N1219, N1220, N1221, N1222, N1223,
         N1224, N1225, N1226, N1227, N1228, N1229, N1230, N1231, N1232, N1233,
         N1234, N1235, N1236, N1237, N1238, N1239, N1240, N1241, N1242, N1243,
         N1244, N1245, N1246, N1247, N1248, N1249, N1250, N1251, N1252, N1253,
         N1254, N1255, N1256, N1257, N1258, N1259, N1260, N1261, N1262, N1263,
         N1264, N1265, N1266, N1267, N1268, N1269, N1270, N1271, N1272, N1273,
         N1274, N1275, N1276, N1277, N1278, N1279, N1280, N1281, N1282, N1283,
         N1284, N1285, N1286, N1287, N1288, N1289, N1290, N1291, N1292, N1293,
         N1294, N1295, N1296, N1297, N1298, N1299, N1300, N1301, N1302, N1303,
         N1304, N1305, N1306, N1307, N1308, N1309, N1310, N1311, N1312, N1313,
         N1314, N1315, N1316, N1317, N1318, N1319, N1320, N1321, N1322, N1323,
         N1324, N1325, N1326, N1327, N1328, N1329, N1330, N1331, N1332, N1333,
         N1334, N1335, N1336, N1337, N1338, N1339, N1340, N1341, N1342, N1343,
         N1344, N1345, N1346, N1347, N1348, N1349, N1350, N1351, N1352, N1353,
         N1354, N1355, N1356, N1357, N1358, N1359, N1360, N1361, N1362, N1363,
         N1364, N1365, N1366, N1367, N1368, N1369, N1370, N1371, N1372, N1373,
         N1374, N1375, N1376, N1377, N1378, N1379, N1380, N1381, N1382, N1383,
         N1384, N1385, N1386, N1387, N1388, N1389, N1390, N1391, N1392, N1393,
         N1394, N1395, N1396, N1397, N1398, N1399, N1400, N1401, N1402, N1403,
         N1404, N1405, N1406, N1407, N1408, N1409, N1410, N1411, N1412, N1413,
         N1414, N1415, N1416, N1417, N1418, N1419, N1420, N1421, N1422, N1423,
         N1424, N1425, N1426, N1427, N1428, N1429, N1430, N1431, N1432, N1433,
         N1434, N1435, N1436, N1437, N1438, N1439, N1440, N1441, N1442, N1443,
         N1444, N1445, N1446, N1447, N1448, N1449, N1450, N1451, N1452, N1453,
         N1454, N1455, N1456, N1457, N1458, N1459, N1460, N1461, N1462, N1463,
         N1464, N1465, N1466, N1467, N1468, N1469, N1470, N1471, N1472, N1473,
         N1474, N1475, N1476, N1477, N1478, N1479, N1480, N1481, N1482, N1483,
         N1484, N1485, N1486, N1487, N1488, N1489, N1490, N1491, N1492, N1493,
         N1494, N1495, N1496, N1497, N1498, N1499, N1500, N1501, N1502, N1503,
         N1504, N1505, N1506, N1507, N1508, N1509, N1510, N1511, N1512, N1513,
         N1514, N1515, N1516, N1517, N1518, N1519, N1520, N1521, N1522, N1523,
         N1524, N1525, N1526, N1527, N1528, N1529, N1530, N1531, N1532, N1533,
         N1534, N1535, N1536, N1537, N1538, N1539, N1540, N1541, N1542, N1543,
         N1544, N1545, N1546, N1547, N1548, N1549, N1550, N1551, N1552, N1553,
         N1554, N1555, N1556, N1557, N1558, N1559, N1560, N1561, N1562, N1563,
         N1564, N1565, N1566, N1567, N1568, N1569, N1570, N1571, N1572, N1573,
         N1574, N1575, N1576, N1577, N1578, N1579, N1580, N1581, N1582, N1583,
         N1584, N1585, N1586, N1587, N1588, N1589, N1590, N1591, N1592, N1593,
         N1594, N1595, N1596, N1597, N1598, N1599, N1600, N1601, N1602, N1603,
         N1604, N1605, N1606, N1607, N1608, N1609, N1610, N1611, N1612, N1613,
         N1614, N1615, N1616, N1617, \round_in[1][1599] , \round_in[1][1598] ,
         \round_in[1][1597] , \round_in[1][1596] , \round_in[1][1595] ,
         \round_in[1][1594] , \round_in[1][1593] , \round_in[1][1592] ,
         \round_in[1][1591] , \round_in[1][1590] , \round_in[1][1589] ,
         \round_in[1][1588] , \round_in[1][1587] , \round_in[1][1586] ,
         \round_in[1][1585] , \round_in[1][1584] , \round_in[1][1583] ,
         \round_in[1][1582] , \round_in[1][1581] , \round_in[1][1580] ,
         \round_in[1][1579] , \round_in[1][1578] , \round_in[1][1577] ,
         \round_in[1][1576] , \round_in[1][1575] , \round_in[1][1574] ,
         \round_in[1][1573] , \round_in[1][1572] , \round_in[1][1571] ,
         \round_in[1][1570] , \round_in[1][1569] , \round_in[1][1568] ,
         \round_in[1][1567] , \round_in[1][1566] , \round_in[1][1565] ,
         \round_in[1][1564] , \round_in[1][1563] , \round_in[1][1562] ,
         \round_in[1][1561] , \round_in[1][1560] , \round_in[1][1559] ,
         \round_in[1][1558] , \round_in[1][1557] , \round_in[1][1556] ,
         \round_in[1][1555] , \round_in[1][1554] , \round_in[1][1553] ,
         \round_in[1][1552] , \round_in[1][1551] , \round_in[1][1550] ,
         \round_in[1][1549] , \round_in[1][1548] , \round_in[1][1547] ,
         \round_in[1][1546] , \round_in[1][1545] , \round_in[1][1544] ,
         \round_in[1][1543] , \round_in[1][1542] , \round_in[1][1541] ,
         \round_in[1][1540] , \round_in[1][1539] , \round_in[1][1538] ,
         \round_in[1][1537] , \round_in[1][1536] , \round_in[1][1535] ,
         \round_in[1][1534] , \round_in[1][1533] , \round_in[1][1532] ,
         \round_in[1][1531] , \round_in[1][1530] , \round_in[1][1529] ,
         \round_in[1][1528] , \round_in[1][1527] , \round_in[1][1526] ,
         \round_in[1][1525] , \round_in[1][1524] , \round_in[1][1523] ,
         \round_in[1][1522] , \round_in[1][1521] , \round_in[1][1520] ,
         \round_in[1][1519] , \round_in[1][1518] , \round_in[1][1517] ,
         \round_in[1][1516] , \round_in[1][1515] , \round_in[1][1514] ,
         \round_in[1][1513] , \round_in[1][1512] , \round_in[1][1511] ,
         \round_in[1][1510] , \round_in[1][1509] , \round_in[1][1508] ,
         \round_in[1][1507] , \round_in[1][1506] , \round_in[1][1505] ,
         \round_in[1][1504] , \round_in[1][1503] , \round_in[1][1502] ,
         \round_in[1][1501] , \round_in[1][1500] , \round_in[1][1499] ,
         \round_in[1][1498] , \round_in[1][1497] , \round_in[1][1496] ,
         \round_in[1][1495] , \round_in[1][1494] , \round_in[1][1493] ,
         \round_in[1][1492] , \round_in[1][1491] , \round_in[1][1490] ,
         \round_in[1][1489] , \round_in[1][1488] , \round_in[1][1487] ,
         \round_in[1][1486] , \round_in[1][1485] , \round_in[1][1484] ,
         \round_in[1][1483] , \round_in[1][1482] , \round_in[1][1481] ,
         \round_in[1][1480] , \round_in[1][1479] , \round_in[1][1478] ,
         \round_in[1][1477] , \round_in[1][1476] , \round_in[1][1475] ,
         \round_in[1][1474] , \round_in[1][1473] , \round_in[1][1472] ,
         \round_in[1][1471] , \round_in[1][1470] , \round_in[1][1469] ,
         \round_in[1][1468] , \round_in[1][1467] , \round_in[1][1466] ,
         \round_in[1][1465] , \round_in[1][1464] , \round_in[1][1463] ,
         \round_in[1][1462] , \round_in[1][1461] , \round_in[1][1460] ,
         \round_in[1][1459] , \round_in[1][1458] , \round_in[1][1457] ,
         \round_in[1][1456] , \round_in[1][1455] , \round_in[1][1454] ,
         \round_in[1][1453] , \round_in[1][1452] , \round_in[1][1451] ,
         \round_in[1][1450] , \round_in[1][1449] , \round_in[1][1448] ,
         \round_in[1][1447] , \round_in[1][1446] , \round_in[1][1445] ,
         \round_in[1][1444] , \round_in[1][1443] , \round_in[1][1442] ,
         \round_in[1][1441] , \round_in[1][1440] , \round_in[1][1439] ,
         \round_in[1][1438] , \round_in[1][1437] , \round_in[1][1436] ,
         \round_in[1][1435] , \round_in[1][1434] , \round_in[1][1433] ,
         \round_in[1][1432] , \round_in[1][1431] , \round_in[1][1430] ,
         \round_in[1][1429] , \round_in[1][1428] , \round_in[1][1427] ,
         \round_in[1][1426] , \round_in[1][1425] , \round_in[1][1424] ,
         \round_in[1][1423] , \round_in[1][1422] , \round_in[1][1421] ,
         \round_in[1][1420] , \round_in[1][1419] , \round_in[1][1418] ,
         \round_in[1][1417] , \round_in[1][1416] , \round_in[1][1415] ,
         \round_in[1][1414] , \round_in[1][1413] , \round_in[1][1412] ,
         \round_in[1][1411] , \round_in[1][1410] , \round_in[1][1409] ,
         \round_in[1][1408] , \round_in[1][1407] , \round_in[1][1406] ,
         \round_in[1][1405] , \round_in[1][1404] , \round_in[1][1403] ,
         \round_in[1][1402] , \round_in[1][1401] , \round_in[1][1400] ,
         \round_in[1][1399] , \round_in[1][1398] , \round_in[1][1397] ,
         \round_in[1][1396] , \round_in[1][1395] , \round_in[1][1394] ,
         \round_in[1][1393] , \round_in[1][1392] , \round_in[1][1391] ,
         \round_in[1][1390] , \round_in[1][1389] , \round_in[1][1388] ,
         \round_in[1][1387] , \round_in[1][1386] , \round_in[1][1385] ,
         \round_in[1][1384] , \round_in[1][1383] , \round_in[1][1382] ,
         \round_in[1][1381] , \round_in[1][1380] , \round_in[1][1379] ,
         \round_in[1][1378] , \round_in[1][1377] , \round_in[1][1376] ,
         \round_in[1][1375] , \round_in[1][1374] , \round_in[1][1373] ,
         \round_in[1][1372] , \round_in[1][1371] , \round_in[1][1370] ,
         \round_in[1][1369] , \round_in[1][1368] , \round_in[1][1367] ,
         \round_in[1][1366] , \round_in[1][1365] , \round_in[1][1364] ,
         \round_in[1][1363] , \round_in[1][1362] , \round_in[1][1361] ,
         \round_in[1][1360] , \round_in[1][1359] , \round_in[1][1358] ,
         \round_in[1][1357] , \round_in[1][1356] , \round_in[1][1355] ,
         \round_in[1][1354] , \round_in[1][1353] , \round_in[1][1352] ,
         \round_in[1][1351] , \round_in[1][1350] , \round_in[1][1349] ,
         \round_in[1][1348] , \round_in[1][1347] , \round_in[1][1346] ,
         \round_in[1][1345] , \round_in[1][1344] , \round_in[1][1343] ,
         \round_in[1][1342] , \round_in[1][1341] , \round_in[1][1340] ,
         \round_in[1][1339] , \round_in[1][1338] , \round_in[1][1337] ,
         \round_in[1][1336] , \round_in[1][1335] , \round_in[1][1334] ,
         \round_in[1][1333] , \round_in[1][1332] , \round_in[1][1331] ,
         \round_in[1][1330] , \round_in[1][1329] , \round_in[1][1328] ,
         \round_in[1][1327] , \round_in[1][1326] , \round_in[1][1325] ,
         \round_in[1][1324] , \round_in[1][1323] , \round_in[1][1322] ,
         \round_in[1][1321] , \round_in[1][1320] , \round_in[1][1319] ,
         \round_in[1][1318] , \round_in[1][1317] , \round_in[1][1316] ,
         \round_in[1][1315] , \round_in[1][1314] , \round_in[1][1313] ,
         \round_in[1][1312] , \round_in[1][1311] , \round_in[1][1310] ,
         \round_in[1][1309] , \round_in[1][1308] , \round_in[1][1307] ,
         \round_in[1][1306] , \round_in[1][1305] , \round_in[1][1304] ,
         \round_in[1][1303] , \round_in[1][1302] , \round_in[1][1301] ,
         \round_in[1][1300] , \round_in[1][1299] , \round_in[1][1298] ,
         \round_in[1][1297] , \round_in[1][1296] , \round_in[1][1295] ,
         \round_in[1][1294] , \round_in[1][1293] , \round_in[1][1292] ,
         \round_in[1][1291] , \round_in[1][1290] , \round_in[1][1289] ,
         \round_in[1][1288] , \round_in[1][1287] , \round_in[1][1286] ,
         \round_in[1][1285] , \round_in[1][1284] , \round_in[1][1283] ,
         \round_in[1][1282] , \round_in[1][1281] , \round_in[1][1280] ,
         \round_in[1][1279] , \round_in[1][1278] , \round_in[1][1277] ,
         \round_in[1][1276] , \round_in[1][1275] , \round_in[1][1274] ,
         \round_in[1][1273] , \round_in[1][1272] , \round_in[1][1271] ,
         \round_in[1][1270] , \round_in[1][1269] , \round_in[1][1268] ,
         \round_in[1][1267] , \round_in[1][1266] , \round_in[1][1265] ,
         \round_in[1][1264] , \round_in[1][1263] , \round_in[1][1262] ,
         \round_in[1][1261] , \round_in[1][1260] , \round_in[1][1259] ,
         \round_in[1][1258] , \round_in[1][1257] , \round_in[1][1256] ,
         \round_in[1][1255] , \round_in[1][1254] , \round_in[1][1253] ,
         \round_in[1][1252] , \round_in[1][1251] , \round_in[1][1250] ,
         \round_in[1][1249] , \round_in[1][1248] , \round_in[1][1247] ,
         \round_in[1][1246] , \round_in[1][1245] , \round_in[1][1244] ,
         \round_in[1][1243] , \round_in[1][1242] , \round_in[1][1241] ,
         \round_in[1][1240] , \round_in[1][1239] , \round_in[1][1238] ,
         \round_in[1][1237] , \round_in[1][1236] , \round_in[1][1235] ,
         \round_in[1][1234] , \round_in[1][1233] , \round_in[1][1232] ,
         \round_in[1][1231] , \round_in[1][1230] , \round_in[1][1229] ,
         \round_in[1][1228] , \round_in[1][1227] , \round_in[1][1226] ,
         \round_in[1][1225] , \round_in[1][1224] , \round_in[1][1223] ,
         \round_in[1][1222] , \round_in[1][1221] , \round_in[1][1220] ,
         \round_in[1][1219] , \round_in[1][1218] , \round_in[1][1217] ,
         \round_in[1][1216] , \round_in[1][1215] , \round_in[1][1214] ,
         \round_in[1][1213] , \round_in[1][1212] , \round_in[1][1211] ,
         \round_in[1][1210] , \round_in[1][1209] , \round_in[1][1208] ,
         \round_in[1][1207] , \round_in[1][1206] , \round_in[1][1205] ,
         \round_in[1][1204] , \round_in[1][1203] , \round_in[1][1202] ,
         \round_in[1][1201] , \round_in[1][1200] , \round_in[1][1199] ,
         \round_in[1][1198] , \round_in[1][1197] , \round_in[1][1196] ,
         \round_in[1][1195] , \round_in[1][1194] , \round_in[1][1193] ,
         \round_in[1][1192] , \round_in[1][1191] , \round_in[1][1190] ,
         \round_in[1][1189] , \round_in[1][1188] , \round_in[1][1187] ,
         \round_in[1][1186] , \round_in[1][1185] , \round_in[1][1184] ,
         \round_in[1][1183] , \round_in[1][1182] , \round_in[1][1181] ,
         \round_in[1][1180] , \round_in[1][1179] , \round_in[1][1178] ,
         \round_in[1][1177] , \round_in[1][1176] , \round_in[1][1175] ,
         \round_in[1][1174] , \round_in[1][1173] , \round_in[1][1172] ,
         \round_in[1][1171] , \round_in[1][1170] , \round_in[1][1169] ,
         \round_in[1][1168] , \round_in[1][1167] , \round_in[1][1166] ,
         \round_in[1][1165] , \round_in[1][1164] , \round_in[1][1163] ,
         \round_in[1][1162] , \round_in[1][1161] , \round_in[1][1160] ,
         \round_in[1][1159] , \round_in[1][1158] , \round_in[1][1157] ,
         \round_in[1][1156] , \round_in[1][1155] , \round_in[1][1154] ,
         \round_in[1][1153] , \round_in[1][1152] , \round_in[1][1151] ,
         \round_in[1][1150] , \round_in[1][1149] , \round_in[1][1148] ,
         \round_in[1][1147] , \round_in[1][1146] , \round_in[1][1145] ,
         \round_in[1][1144] , \round_in[1][1143] , \round_in[1][1142] ,
         \round_in[1][1141] , \round_in[1][1140] , \round_in[1][1139] ,
         \round_in[1][1138] , \round_in[1][1137] , \round_in[1][1136] ,
         \round_in[1][1135] , \round_in[1][1134] , \round_in[1][1133] ,
         \round_in[1][1132] , \round_in[1][1131] , \round_in[1][1130] ,
         \round_in[1][1129] , \round_in[1][1128] , \round_in[1][1127] ,
         \round_in[1][1126] , \round_in[1][1125] , \round_in[1][1124] ,
         \round_in[1][1123] , \round_in[1][1122] , \round_in[1][1121] ,
         \round_in[1][1120] , \round_in[1][1119] , \round_in[1][1118] ,
         \round_in[1][1117] , \round_in[1][1116] , \round_in[1][1115] ,
         \round_in[1][1114] , \round_in[1][1113] , \round_in[1][1112] ,
         \round_in[1][1111] , \round_in[1][1110] , \round_in[1][1109] ,
         \round_in[1][1108] , \round_in[1][1107] , \round_in[1][1106] ,
         \round_in[1][1105] , \round_in[1][1104] , \round_in[1][1103] ,
         \round_in[1][1102] , \round_in[1][1101] , \round_in[1][1100] ,
         \round_in[1][1099] , \round_in[1][1098] , \round_in[1][1097] ,
         \round_in[1][1096] , \round_in[1][1095] , \round_in[1][1094] ,
         \round_in[1][1093] , \round_in[1][1092] , \round_in[1][1091] ,
         \round_in[1][1090] , \round_in[1][1089] , \round_in[1][1088] ,
         \round_in[1][1087] , \round_in[1][1086] , \round_in[1][1085] ,
         \round_in[1][1084] , \round_in[1][1083] , \round_in[1][1082] ,
         \round_in[1][1081] , \round_in[1][1080] , \round_in[1][1079] ,
         \round_in[1][1078] , \round_in[1][1077] , \round_in[1][1076] ,
         \round_in[1][1075] , \round_in[1][1074] , \round_in[1][1073] ,
         \round_in[1][1072] , \round_in[1][1071] , \round_in[1][1070] ,
         \round_in[1][1069] , \round_in[1][1068] , \round_in[1][1067] ,
         \round_in[1][1066] , \round_in[1][1065] , \round_in[1][1064] ,
         \round_in[1][1063] , \round_in[1][1062] , \round_in[1][1061] ,
         \round_in[1][1060] , \round_in[1][1059] , \round_in[1][1058] ,
         \round_in[1][1057] , \round_in[1][1056] , \round_in[1][1055] ,
         \round_in[1][1054] , \round_in[1][1053] , \round_in[1][1052] ,
         \round_in[1][1051] , \round_in[1][1050] , \round_in[1][1049] ,
         \round_in[1][1048] , \round_in[1][1047] , \round_in[1][1046] ,
         \round_in[1][1045] , \round_in[1][1044] , \round_in[1][1043] ,
         \round_in[1][1042] , \round_in[1][1041] , \round_in[1][1040] ,
         \round_in[1][1039] , \round_in[1][1038] , \round_in[1][1037] ,
         \round_in[1][1036] , \round_in[1][1035] , \round_in[1][1034] ,
         \round_in[1][1033] , \round_in[1][1032] , \round_in[1][1031] ,
         \round_in[1][1030] , \round_in[1][1029] , \round_in[1][1028] ,
         \round_in[1][1027] , \round_in[1][1026] , \round_in[1][1025] ,
         \round_in[1][1024] , \round_in[1][1023] , \round_in[1][1022] ,
         \round_in[1][1021] , \round_in[1][1020] , \round_in[1][1019] ,
         \round_in[1][1018] , \round_in[1][1017] , \round_in[1][1016] ,
         \round_in[1][1015] , \round_in[1][1014] , \round_in[1][1013] ,
         \round_in[1][1012] , \round_in[1][1011] , \round_in[1][1010] ,
         \round_in[1][1009] , \round_in[1][1008] , \round_in[1][1007] ,
         \round_in[1][1006] , \round_in[1][1005] , \round_in[1][1004] ,
         \round_in[1][1003] , \round_in[1][1002] , \round_in[1][1001] ,
         \round_in[1][1000] , \round_in[1][999] , \round_in[1][998] ,
         \round_in[1][997] , \round_in[1][996] , \round_in[1][995] ,
         \round_in[1][994] , \round_in[1][993] , \round_in[1][992] ,
         \round_in[1][991] , \round_in[1][990] , \round_in[1][989] ,
         \round_in[1][988] , \round_in[1][987] , \round_in[1][986] ,
         \round_in[1][985] , \round_in[1][984] , \round_in[1][983] ,
         \round_in[1][982] , \round_in[1][981] , \round_in[1][980] ,
         \round_in[1][979] , \round_in[1][978] , \round_in[1][977] ,
         \round_in[1][976] , \round_in[1][975] , \round_in[1][974] ,
         \round_in[1][973] , \round_in[1][972] , \round_in[1][971] ,
         \round_in[1][970] , \round_in[1][969] , \round_in[1][968] ,
         \round_in[1][967] , \round_in[1][966] , \round_in[1][965] ,
         \round_in[1][964] , \round_in[1][963] , \round_in[1][962] ,
         \round_in[1][961] , \round_in[1][960] , \round_in[1][959] ,
         \round_in[1][958] , \round_in[1][957] , \round_in[1][956] ,
         \round_in[1][955] , \round_in[1][954] , \round_in[1][953] ,
         \round_in[1][952] , \round_in[1][951] , \round_in[1][950] ,
         \round_in[1][949] , \round_in[1][948] , \round_in[1][947] ,
         \round_in[1][946] , \round_in[1][945] , \round_in[1][944] ,
         \round_in[1][943] , \round_in[1][942] , \round_in[1][941] ,
         \round_in[1][940] , \round_in[1][939] , \round_in[1][938] ,
         \round_in[1][937] , \round_in[1][936] , \round_in[1][935] ,
         \round_in[1][934] , \round_in[1][933] , \round_in[1][932] ,
         \round_in[1][931] , \round_in[1][930] , \round_in[1][929] ,
         \round_in[1][928] , \round_in[1][927] , \round_in[1][926] ,
         \round_in[1][925] , \round_in[1][924] , \round_in[1][923] ,
         \round_in[1][922] , \round_in[1][921] , \round_in[1][920] ,
         \round_in[1][919] , \round_in[1][918] , \round_in[1][917] ,
         \round_in[1][916] , \round_in[1][915] , \round_in[1][914] ,
         \round_in[1][913] , \round_in[1][912] , \round_in[1][911] ,
         \round_in[1][910] , \round_in[1][909] , \round_in[1][908] ,
         \round_in[1][907] , \round_in[1][906] , \round_in[1][905] ,
         \round_in[1][904] , \round_in[1][903] , \round_in[1][902] ,
         \round_in[1][901] , \round_in[1][900] , \round_in[1][899] ,
         \round_in[1][898] , \round_in[1][897] , \round_in[1][896] ,
         \round_in[1][895] , \round_in[1][894] , \round_in[1][893] ,
         \round_in[1][892] , \round_in[1][891] , \round_in[1][890] ,
         \round_in[1][889] , \round_in[1][888] , \round_in[1][887] ,
         \round_in[1][886] , \round_in[1][885] , \round_in[1][884] ,
         \round_in[1][883] , \round_in[1][882] , \round_in[1][881] ,
         \round_in[1][880] , \round_in[1][879] , \round_in[1][878] ,
         \round_in[1][877] , \round_in[1][876] , \round_in[1][875] ,
         \round_in[1][874] , \round_in[1][873] , \round_in[1][872] ,
         \round_in[1][871] , \round_in[1][870] , \round_in[1][869] ,
         \round_in[1][868] , \round_in[1][867] , \round_in[1][866] ,
         \round_in[1][865] , \round_in[1][864] , \round_in[1][863] ,
         \round_in[1][862] , \round_in[1][861] , \round_in[1][860] ,
         \round_in[1][859] , \round_in[1][858] , \round_in[1][857] ,
         \round_in[1][856] , \round_in[1][855] , \round_in[1][854] ,
         \round_in[1][853] , \round_in[1][852] , \round_in[1][851] ,
         \round_in[1][850] , \round_in[1][849] , \round_in[1][848] ,
         \round_in[1][847] , \round_in[1][846] , \round_in[1][845] ,
         \round_in[1][844] , \round_in[1][843] , \round_in[1][842] ,
         \round_in[1][841] , \round_in[1][840] , \round_in[1][839] ,
         \round_in[1][838] , \round_in[1][837] , \round_in[1][836] ,
         \round_in[1][835] , \round_in[1][834] , \round_in[1][833] ,
         \round_in[1][832] , \round_in[1][831] , \round_in[1][830] ,
         \round_in[1][829] , \round_in[1][828] , \round_in[1][827] ,
         \round_in[1][826] , \round_in[1][825] , \round_in[1][824] ,
         \round_in[1][823] , \round_in[1][822] , \round_in[1][821] ,
         \round_in[1][820] , \round_in[1][819] , \round_in[1][818] ,
         \round_in[1][817] , \round_in[1][816] , \round_in[1][815] ,
         \round_in[1][814] , \round_in[1][813] , \round_in[1][812] ,
         \round_in[1][811] , \round_in[1][810] , \round_in[1][809] ,
         \round_in[1][808] , \round_in[1][807] , \round_in[1][806] ,
         \round_in[1][805] , \round_in[1][804] , \round_in[1][803] ,
         \round_in[1][802] , \round_in[1][801] , \round_in[1][800] ,
         \round_in[1][799] , \round_in[1][798] , \round_in[1][797] ,
         \round_in[1][796] , \round_in[1][795] , \round_in[1][794] ,
         \round_in[1][793] , \round_in[1][792] , \round_in[1][791] ,
         \round_in[1][790] , \round_in[1][789] , \round_in[1][788] ,
         \round_in[1][787] , \round_in[1][786] , \round_in[1][785] ,
         \round_in[1][784] , \round_in[1][783] , \round_in[1][782] ,
         \round_in[1][781] , \round_in[1][780] , \round_in[1][779] ,
         \round_in[1][778] , \round_in[1][777] , \round_in[1][776] ,
         \round_in[1][775] , \round_in[1][774] , \round_in[1][773] ,
         \round_in[1][772] , \round_in[1][771] , \round_in[1][770] ,
         \round_in[1][769] , \round_in[1][768] , \round_in[1][767] ,
         \round_in[1][766] , \round_in[1][765] , \round_in[1][764] ,
         \round_in[1][763] , \round_in[1][762] , \round_in[1][761] ,
         \round_in[1][760] , \round_in[1][759] , \round_in[1][758] ,
         \round_in[1][757] , \round_in[1][756] , \round_in[1][755] ,
         \round_in[1][754] , \round_in[1][753] , \round_in[1][752] ,
         \round_in[1][751] , \round_in[1][750] , \round_in[1][749] ,
         \round_in[1][748] , \round_in[1][747] , \round_in[1][746] ,
         \round_in[1][745] , \round_in[1][744] , \round_in[1][743] ,
         \round_in[1][742] , \round_in[1][741] , \round_in[1][740] ,
         \round_in[1][739] , \round_in[1][738] , \round_in[1][737] ,
         \round_in[1][736] , \round_in[1][735] , \round_in[1][734] ,
         \round_in[1][733] , \round_in[1][732] , \round_in[1][731] ,
         \round_in[1][730] , \round_in[1][729] , \round_in[1][728] ,
         \round_in[1][727] , \round_in[1][726] , \round_in[1][725] ,
         \round_in[1][724] , \round_in[1][723] , \round_in[1][722] ,
         \round_in[1][721] , \round_in[1][720] , \round_in[1][719] ,
         \round_in[1][718] , \round_in[1][717] , \round_in[1][716] ,
         \round_in[1][715] , \round_in[1][714] , \round_in[1][713] ,
         \round_in[1][712] , \round_in[1][711] , \round_in[1][710] ,
         \round_in[1][709] , \round_in[1][708] , \round_in[1][707] ,
         \round_in[1][706] , \round_in[1][705] , \round_in[1][704] ,
         \round_in[1][703] , \round_in[1][702] , \round_in[1][701] ,
         \round_in[1][700] , \round_in[1][699] , \round_in[1][698] ,
         \round_in[1][697] , \round_in[1][696] , \round_in[1][695] ,
         \round_in[1][694] , \round_in[1][693] , \round_in[1][692] ,
         \round_in[1][691] , \round_in[1][690] , \round_in[1][689] ,
         \round_in[1][688] , \round_in[1][687] , \round_in[1][686] ,
         \round_in[1][685] , \round_in[1][684] , \round_in[1][683] ,
         \round_in[1][682] , \round_in[1][681] , \round_in[1][680] ,
         \round_in[1][679] , \round_in[1][678] , \round_in[1][677] ,
         \round_in[1][676] , \round_in[1][675] , \round_in[1][674] ,
         \round_in[1][673] , \round_in[1][672] , \round_in[1][671] ,
         \round_in[1][670] , \round_in[1][669] , \round_in[1][668] ,
         \round_in[1][667] , \round_in[1][666] , \round_in[1][665] ,
         \round_in[1][664] , \round_in[1][663] , \round_in[1][662] ,
         \round_in[1][661] , \round_in[1][660] , \round_in[1][659] ,
         \round_in[1][658] , \round_in[1][657] , \round_in[1][656] ,
         \round_in[1][655] , \round_in[1][654] , \round_in[1][653] ,
         \round_in[1][652] , \round_in[1][651] , \round_in[1][650] ,
         \round_in[1][649] , \round_in[1][648] , \round_in[1][647] ,
         \round_in[1][646] , \round_in[1][645] , \round_in[1][644] ,
         \round_in[1][643] , \round_in[1][642] , \round_in[1][641] ,
         \round_in[1][640] , \round_in[1][639] , \round_in[1][638] ,
         \round_in[1][637] , \round_in[1][636] , \round_in[1][635] ,
         \round_in[1][634] , \round_in[1][633] , \round_in[1][632] ,
         \round_in[1][631] , \round_in[1][630] , \round_in[1][629] ,
         \round_in[1][628] , \round_in[1][627] , \round_in[1][626] ,
         \round_in[1][625] , \round_in[1][624] , \round_in[1][623] ,
         \round_in[1][622] , \round_in[1][621] , \round_in[1][620] ,
         \round_in[1][619] , \round_in[1][618] , \round_in[1][617] ,
         \round_in[1][616] , \round_in[1][615] , \round_in[1][614] ,
         \round_in[1][613] , \round_in[1][612] , \round_in[1][611] ,
         \round_in[1][610] , \round_in[1][609] , \round_in[1][608] ,
         \round_in[1][607] , \round_in[1][606] , \round_in[1][605] ,
         \round_in[1][604] , \round_in[1][603] , \round_in[1][602] ,
         \round_in[1][601] , \round_in[1][600] , \round_in[1][599] ,
         \round_in[1][598] , \round_in[1][597] , \round_in[1][596] ,
         \round_in[1][595] , \round_in[1][594] , \round_in[1][593] ,
         \round_in[1][592] , \round_in[1][591] , \round_in[1][590] ,
         \round_in[1][589] , \round_in[1][588] , \round_in[1][587] ,
         \round_in[1][586] , \round_in[1][585] , \round_in[1][584] ,
         \round_in[1][583] , \round_in[1][582] , \round_in[1][581] ,
         \round_in[1][580] , \round_in[1][579] , \round_in[1][578] ,
         \round_in[1][577] , \round_in[1][576] , \round_in[1][575] ,
         \round_in[1][574] , \round_in[1][573] , \round_in[1][572] ,
         \round_in[1][571] , \round_in[1][570] , \round_in[1][569] ,
         \round_in[1][568] , \round_in[1][567] , \round_in[1][566] ,
         \round_in[1][565] , \round_in[1][564] , \round_in[1][563] ,
         \round_in[1][562] , \round_in[1][561] , \round_in[1][560] ,
         \round_in[1][559] , \round_in[1][558] , \round_in[1][557] ,
         \round_in[1][556] , \round_in[1][555] , \round_in[1][554] ,
         \round_in[1][553] , \round_in[1][552] , \round_in[1][551] ,
         \round_in[1][550] , \round_in[1][549] , \round_in[1][548] ,
         \round_in[1][547] , \round_in[1][546] , \round_in[1][545] ,
         \round_in[1][544] , \round_in[1][543] , \round_in[1][542] ,
         \round_in[1][541] , \round_in[1][540] , \round_in[1][539] ,
         \round_in[1][538] , \round_in[1][537] , \round_in[1][536] ,
         \round_in[1][535] , \round_in[1][534] , \round_in[1][533] ,
         \round_in[1][532] , \round_in[1][531] , \round_in[1][530] ,
         \round_in[1][529] , \round_in[1][528] , \round_in[1][527] ,
         \round_in[1][526] , \round_in[1][525] , \round_in[1][524] ,
         \round_in[1][523] , \round_in[1][522] , \round_in[1][521] ,
         \round_in[1][520] , \round_in[1][519] , \round_in[1][518] ,
         \round_in[1][517] , \round_in[1][516] , \round_in[1][515] ,
         \round_in[1][514] , \round_in[1][513] , \round_in[1][512] ,
         \round_in[1][511] , \round_in[1][510] , \round_in[1][509] ,
         \round_in[1][508] , \round_in[1][507] , \round_in[1][506] ,
         \round_in[1][505] , \round_in[1][504] , \round_in[1][503] ,
         \round_in[1][502] , \round_in[1][501] , \round_in[1][500] ,
         \round_in[1][499] , \round_in[1][498] , \round_in[1][497] ,
         \round_in[1][496] , \round_in[1][495] , \round_in[1][494] ,
         \round_in[1][493] , \round_in[1][492] , \round_in[1][491] ,
         \round_in[1][490] , \round_in[1][489] , \round_in[1][488] ,
         \round_in[1][487] , \round_in[1][486] , \round_in[1][485] ,
         \round_in[1][484] , \round_in[1][483] , \round_in[1][482] ,
         \round_in[1][481] , \round_in[1][480] , \round_in[1][479] ,
         \round_in[1][478] , \round_in[1][477] , \round_in[1][476] ,
         \round_in[1][475] , \round_in[1][474] , \round_in[1][473] ,
         \round_in[1][472] , \round_in[1][471] , \round_in[1][470] ,
         \round_in[1][469] , \round_in[1][468] , \round_in[1][467] ,
         \round_in[1][466] , \round_in[1][465] , \round_in[1][464] ,
         \round_in[1][463] , \round_in[1][462] , \round_in[1][461] ,
         \round_in[1][460] , \round_in[1][459] , \round_in[1][458] ,
         \round_in[1][457] , \round_in[1][456] , \round_in[1][455] ,
         \round_in[1][454] , \round_in[1][453] , \round_in[1][452] ,
         \round_in[1][451] , \round_in[1][450] , \round_in[1][449] ,
         \round_in[1][448] , \round_in[1][447] , \round_in[1][446] ,
         \round_in[1][445] , \round_in[1][444] , \round_in[1][443] ,
         \round_in[1][442] , \round_in[1][441] , \round_in[1][440] ,
         \round_in[1][439] , \round_in[1][438] , \round_in[1][437] ,
         \round_in[1][436] , \round_in[1][435] , \round_in[1][434] ,
         \round_in[1][433] , \round_in[1][432] , \round_in[1][431] ,
         \round_in[1][430] , \round_in[1][429] , \round_in[1][428] ,
         \round_in[1][427] , \round_in[1][426] , \round_in[1][425] ,
         \round_in[1][424] , \round_in[1][423] , \round_in[1][422] ,
         \round_in[1][421] , \round_in[1][420] , \round_in[1][419] ,
         \round_in[1][418] , \round_in[1][417] , \round_in[1][416] ,
         \round_in[1][415] , \round_in[1][414] , \round_in[1][413] ,
         \round_in[1][412] , \round_in[1][411] , \round_in[1][410] ,
         \round_in[1][409] , \round_in[1][408] , \round_in[1][407] ,
         \round_in[1][406] , \round_in[1][405] , \round_in[1][404] ,
         \round_in[1][403] , \round_in[1][402] , \round_in[1][401] ,
         \round_in[1][400] , \round_in[1][399] , \round_in[1][398] ,
         \round_in[1][397] , \round_in[1][396] , \round_in[1][395] ,
         \round_in[1][394] , \round_in[1][393] , \round_in[1][392] ,
         \round_in[1][391] , \round_in[1][390] , \round_in[1][389] ,
         \round_in[1][388] , \round_in[1][387] , \round_in[1][386] ,
         \round_in[1][385] , \round_in[1][384] , \round_in[1][383] ,
         \round_in[1][382] , \round_in[1][381] , \round_in[1][380] ,
         \round_in[1][379] , \round_in[1][378] , \round_in[1][377] ,
         \round_in[1][376] , \round_in[1][375] , \round_in[1][374] ,
         \round_in[1][373] , \round_in[1][372] , \round_in[1][371] ,
         \round_in[1][370] , \round_in[1][369] , \round_in[1][368] ,
         \round_in[1][367] , \round_in[1][366] , \round_in[1][365] ,
         \round_in[1][364] , \round_in[1][363] , \round_in[1][362] ,
         \round_in[1][361] , \round_in[1][360] , \round_in[1][359] ,
         \round_in[1][358] , \round_in[1][357] , \round_in[1][356] ,
         \round_in[1][355] , \round_in[1][354] , \round_in[1][353] ,
         \round_in[1][352] , \round_in[1][351] , \round_in[1][350] ,
         \round_in[1][349] , \round_in[1][348] , \round_in[1][347] ,
         \round_in[1][346] , \round_in[1][345] , \round_in[1][344] ,
         \round_in[1][343] , \round_in[1][342] , \round_in[1][341] ,
         \round_in[1][340] , \round_in[1][339] , \round_in[1][338] ,
         \round_in[1][337] , \round_in[1][336] , \round_in[1][335] ,
         \round_in[1][334] , \round_in[1][333] , \round_in[1][332] ,
         \round_in[1][331] , \round_in[1][330] , \round_in[1][329] ,
         \round_in[1][328] , \round_in[1][327] , \round_in[1][326] ,
         \round_in[1][325] , \round_in[1][324] , \round_in[1][323] ,
         \round_in[1][322] , \round_in[1][321] , \round_in[1][320] ,
         \round_in[1][319] , \round_in[1][318] , \round_in[1][317] ,
         \round_in[1][316] , \round_in[1][315] , \round_in[1][314] ,
         \round_in[1][313] , \round_in[1][312] , \round_in[1][311] ,
         \round_in[1][310] , \round_in[1][309] , \round_in[1][308] ,
         \round_in[1][307] , \round_in[1][306] , \round_in[1][305] ,
         \round_in[1][304] , \round_in[1][303] , \round_in[1][302] ,
         \round_in[1][301] , \round_in[1][300] , \round_in[1][299] ,
         \round_in[1][298] , \round_in[1][297] , \round_in[1][296] ,
         \round_in[1][295] , \round_in[1][294] , \round_in[1][293] ,
         \round_in[1][292] , \round_in[1][291] , \round_in[1][290] ,
         \round_in[1][289] , \round_in[1][288] , \round_in[1][287] ,
         \round_in[1][286] , \round_in[1][285] , \round_in[1][284] ,
         \round_in[1][283] , \round_in[1][282] , \round_in[1][281] ,
         \round_in[1][280] , \round_in[1][279] , \round_in[1][278] ,
         \round_in[1][277] , \round_in[1][276] , \round_in[1][275] ,
         \round_in[1][274] , \round_in[1][273] , \round_in[1][272] ,
         \round_in[1][271] , \round_in[1][270] , \round_in[1][269] ,
         \round_in[1][268] , \round_in[1][267] , \round_in[1][266] ,
         \round_in[1][265] , \round_in[1][264] , \round_in[1][263] ,
         \round_in[1][262] , \round_in[1][261] , \round_in[1][260] ,
         \round_in[1][259] , \round_in[1][258] , \round_in[1][257] ,
         \round_in[1][256] , \round_in[1][255] , \round_in[1][254] ,
         \round_in[1][253] , \round_in[1][252] , \round_in[1][251] ,
         \round_in[1][250] , \round_in[1][249] , \round_in[1][248] ,
         \round_in[1][247] , \round_in[1][246] , \round_in[1][245] ,
         \round_in[1][244] , \round_in[1][243] , \round_in[1][242] ,
         \round_in[1][241] , \round_in[1][240] , \round_in[1][239] ,
         \round_in[1][238] , \round_in[1][237] , \round_in[1][236] ,
         \round_in[1][235] , \round_in[1][234] , \round_in[1][233] ,
         \round_in[1][232] , \round_in[1][231] , \round_in[1][230] ,
         \round_in[1][229] , \round_in[1][228] , \round_in[1][227] ,
         \round_in[1][226] , \round_in[1][225] , \round_in[1][224] ,
         \round_in[1][223] , \round_in[1][222] , \round_in[1][221] ,
         \round_in[1][220] , \round_in[1][219] , \round_in[1][218] ,
         \round_in[1][217] , \round_in[1][216] , \round_in[1][215] ,
         \round_in[1][214] , \round_in[1][213] , \round_in[1][212] ,
         \round_in[1][211] , \round_in[1][210] , \round_in[1][209] ,
         \round_in[1][208] , \round_in[1][207] , \round_in[1][206] ,
         \round_in[1][205] , \round_in[1][204] , \round_in[1][203] ,
         \round_in[1][202] , \round_in[1][201] , \round_in[1][200] ,
         \round_in[1][199] , \round_in[1][198] , \round_in[1][197] ,
         \round_in[1][196] , \round_in[1][195] , \round_in[1][194] ,
         \round_in[1][193] , \round_in[1][192] , \round_in[1][191] ,
         \round_in[1][190] , \round_in[1][189] , \round_in[1][188] ,
         \round_in[1][187] , \round_in[1][186] , \round_in[1][185] ,
         \round_in[1][184] , \round_in[1][183] , \round_in[1][182] ,
         \round_in[1][181] , \round_in[1][180] , \round_in[1][179] ,
         \round_in[1][178] , \round_in[1][177] , \round_in[1][176] ,
         \round_in[1][175] , \round_in[1][174] , \round_in[1][173] ,
         \round_in[1][172] , \round_in[1][171] , \round_in[1][170] ,
         \round_in[1][169] , \round_in[1][168] , \round_in[1][167] ,
         \round_in[1][166] , \round_in[1][165] , \round_in[1][164] ,
         \round_in[1][163] , \round_in[1][162] , \round_in[1][161] ,
         \round_in[1][160] , \round_in[1][159] , \round_in[1][158] ,
         \round_in[1][157] , \round_in[1][156] , \round_in[1][155] ,
         \round_in[1][154] , \round_in[1][153] , \round_in[1][152] ,
         \round_in[1][151] , \round_in[1][150] , \round_in[1][149] ,
         \round_in[1][148] , \round_in[1][147] , \round_in[1][146] ,
         \round_in[1][145] , \round_in[1][144] , \round_in[1][143] ,
         \round_in[1][142] , \round_in[1][141] , \round_in[1][140] ,
         \round_in[1][139] , \round_in[1][138] , \round_in[1][137] ,
         \round_in[1][136] , \round_in[1][135] , \round_in[1][134] ,
         \round_in[1][133] , \round_in[1][132] , \round_in[1][131] ,
         \round_in[1][130] , \round_in[1][129] , \round_in[1][128] ,
         \round_in[1][127] , \round_in[1][126] , \round_in[1][125] ,
         \round_in[1][124] , \round_in[1][123] , \round_in[1][122] ,
         \round_in[1][121] , \round_in[1][120] , \round_in[1][119] ,
         \round_in[1][118] , \round_in[1][117] , \round_in[1][116] ,
         \round_in[1][115] , \round_in[1][114] , \round_in[1][113] ,
         \round_in[1][112] , \round_in[1][111] , \round_in[1][110] ,
         \round_in[1][109] , \round_in[1][108] , \round_in[1][107] ,
         \round_in[1][106] , \round_in[1][105] , \round_in[1][104] ,
         \round_in[1][103] , \round_in[1][102] , \round_in[1][101] ,
         \round_in[1][100] , \round_in[1][99] , \round_in[1][98] ,
         \round_in[1][97] , \round_in[1][96] , \round_in[1][95] ,
         \round_in[1][94] , \round_in[1][93] , \round_in[1][92] ,
         \round_in[1][91] , \round_in[1][90] , \round_in[1][89] ,
         \round_in[1][88] , \round_in[1][87] , \round_in[1][86] ,
         \round_in[1][85] , \round_in[1][84] , \round_in[1][83] ,
         \round_in[1][82] , \round_in[1][81] , \round_in[1][80] ,
         \round_in[1][79] , \round_in[1][78] , \round_in[1][77] ,
         \round_in[1][76] , \round_in[1][75] , \round_in[1][74] ,
         \round_in[1][73] , \round_in[1][72] , \round_in[1][71] ,
         \round_in[1][70] , \round_in[1][69] , \round_in[1][68] ,
         \round_in[1][67] , \round_in[1][66] , \round_in[1][65] ,
         \round_in[1][64] , \round_in[1][63] , \round_in[1][62] ,
         \round_in[1][61] , \round_in[1][60] , \round_in[1][59] ,
         \round_in[1][58] , \round_in[1][57] , \round_in[1][56] ,
         \round_in[1][55] , \round_in[1][54] , \round_in[1][53] ,
         \round_in[1][52] , \round_in[1][51] , \round_in[1][50] ,
         \round_in[1][49] , \round_in[1][48] , \round_in[1][47] ,
         \round_in[1][46] , \round_in[1][45] , \round_in[1][44] ,
         \round_in[1][43] , \round_in[1][42] , \round_in[1][41] ,
         \round_in[1][40] , \round_in[1][39] , \round_in[1][38] ,
         \round_in[1][37] , \round_in[1][36] , \round_in[1][35] ,
         \round_in[1][34] , \round_in[1][33] , \round_in[1][32] ,
         \round_in[1][31] , \round_in[1][30] , \round_in[1][29] ,
         \round_in[1][28] , \round_in[1][27] , \round_in[1][26] ,
         \round_in[1][25] , \round_in[1][24] , \round_in[1][23] ,
         \round_in[1][22] , \round_in[1][21] , \round_in[1][20] ,
         \round_in[1][19] , \round_in[1][18] , \round_in[1][17] ,
         \round_in[1][16] , \round_in[1][15] , \round_in[1][14] ,
         \round_in[1][13] , \round_in[1][12] , \round_in[1][11] ,
         \round_in[1][10] , \round_in[1][9] , \round_in[1][8] ,
         \round_in[1][7] , \round_in[1][6] , \round_in[1][5] ,
         \round_in[1][4] , \round_in[1][3] , \round_in[1][2] ,
         \round_in[1][1] , \round_in[1][0] , \round_in[0][1599] ,
         \round_in[0][1598] , \round_in[0][1597] , \round_in[0][1596] ,
         \round_in[0][1595] , \round_in[0][1594] , \round_in[0][1593] ,
         \round_in[0][1592] , \round_in[0][1591] , \round_in[0][1590] ,
         \round_in[0][1589] , \round_in[0][1588] , \round_in[0][1587] ,
         \round_in[0][1586] , \round_in[0][1585] , \round_in[0][1584] ,
         \round_in[0][1583] , \round_in[0][1582] , \round_in[0][1581] ,
         \round_in[0][1580] , \round_in[0][1579] , \round_in[0][1578] ,
         \round_in[0][1577] , \round_in[0][1576] , \round_in[0][1575] ,
         \round_in[0][1574] , \round_in[0][1573] , \round_in[0][1572] ,
         \round_in[0][1571] , \round_in[0][1570] , \round_in[0][1569] ,
         \round_in[0][1568] , \round_in[0][1567] , \round_in[0][1566] ,
         \round_in[0][1565] , \round_in[0][1564] , \round_in[0][1563] ,
         \round_in[0][1562] , \round_in[0][1561] , \round_in[0][1560] ,
         \round_in[0][1559] , \round_in[0][1558] , \round_in[0][1557] ,
         \round_in[0][1556] , \round_in[0][1555] , \round_in[0][1554] ,
         \round_in[0][1553] , \round_in[0][1552] , \round_in[0][1551] ,
         \round_in[0][1550] , \round_in[0][1549] , \round_in[0][1548] ,
         \round_in[0][1547] , \round_in[0][1546] , \round_in[0][1545] ,
         \round_in[0][1544] , \round_in[0][1543] , \round_in[0][1542] ,
         \round_in[0][1541] , \round_in[0][1540] , \round_in[0][1539] ,
         \round_in[0][1538] , \round_in[0][1537] , \round_in[0][1536] ,
         \round_in[0][1535] , \round_in[0][1534] , \round_in[0][1533] ,
         \round_in[0][1532] , \round_in[0][1531] , \round_in[0][1530] ,
         \round_in[0][1529] , \round_in[0][1528] , \round_in[0][1527] ,
         \round_in[0][1526] , \round_in[0][1525] , \round_in[0][1524] ,
         \round_in[0][1523] , \round_in[0][1522] , \round_in[0][1521] ,
         \round_in[0][1520] , \round_in[0][1519] , \round_in[0][1518] ,
         \round_in[0][1517] , \round_in[0][1516] , \round_in[0][1515] ,
         \round_in[0][1514] , \round_in[0][1513] , \round_in[0][1512] ,
         \round_in[0][1511] , \round_in[0][1510] , \round_in[0][1509] ,
         \round_in[0][1508] , \round_in[0][1507] , \round_in[0][1506] ,
         \round_in[0][1505] , \round_in[0][1504] , \round_in[0][1503] ,
         \round_in[0][1502] , \round_in[0][1501] , \round_in[0][1500] ,
         \round_in[0][1499] , \round_in[0][1498] , \round_in[0][1497] ,
         \round_in[0][1496] , \round_in[0][1495] , \round_in[0][1494] ,
         \round_in[0][1493] , \round_in[0][1492] , \round_in[0][1491] ,
         \round_in[0][1490] , \round_in[0][1489] , \round_in[0][1488] ,
         \round_in[0][1487] , \round_in[0][1486] , \round_in[0][1485] ,
         \round_in[0][1484] , \round_in[0][1483] , \round_in[0][1482] ,
         \round_in[0][1481] , \round_in[0][1480] , \round_in[0][1479] ,
         \round_in[0][1478] , \round_in[0][1477] , \round_in[0][1476] ,
         \round_in[0][1475] , \round_in[0][1474] , \round_in[0][1473] ,
         \round_in[0][1472] , \round_in[0][1471] , \round_in[0][1470] ,
         \round_in[0][1469] , \round_in[0][1468] , \round_in[0][1467] ,
         \round_in[0][1466] , \round_in[0][1465] , \round_in[0][1464] ,
         \round_in[0][1463] , \round_in[0][1462] , \round_in[0][1461] ,
         \round_in[0][1460] , \round_in[0][1459] , \round_in[0][1458] ,
         \round_in[0][1457] , \round_in[0][1456] , \round_in[0][1455] ,
         \round_in[0][1454] , \round_in[0][1453] , \round_in[0][1452] ,
         \round_in[0][1451] , \round_in[0][1450] , \round_in[0][1449] ,
         \round_in[0][1448] , \round_in[0][1447] , \round_in[0][1446] ,
         \round_in[0][1445] , \round_in[0][1444] , \round_in[0][1443] ,
         \round_in[0][1442] , \round_in[0][1441] , \round_in[0][1440] ,
         \round_in[0][1439] , \round_in[0][1438] , \round_in[0][1437] ,
         \round_in[0][1436] , \round_in[0][1435] , \round_in[0][1434] ,
         \round_in[0][1433] , \round_in[0][1432] , \round_in[0][1431] ,
         \round_in[0][1430] , \round_in[0][1429] , \round_in[0][1428] ,
         \round_in[0][1427] , \round_in[0][1426] , \round_in[0][1425] ,
         \round_in[0][1424] , \round_in[0][1423] , \round_in[0][1422] ,
         \round_in[0][1421] , \round_in[0][1420] , \round_in[0][1419] ,
         \round_in[0][1418] , \round_in[0][1417] , \round_in[0][1416] ,
         \round_in[0][1415] , \round_in[0][1414] , \round_in[0][1413] ,
         \round_in[0][1412] , \round_in[0][1411] , \round_in[0][1410] ,
         \round_in[0][1409] , \round_in[0][1408] , \round_in[0][1407] ,
         \round_in[0][1406] , \round_in[0][1405] , \round_in[0][1404] ,
         \round_in[0][1403] , \round_in[0][1402] , \round_in[0][1401] ,
         \round_in[0][1400] , \round_in[0][1399] , \round_in[0][1398] ,
         \round_in[0][1397] , \round_in[0][1396] , \round_in[0][1395] ,
         \round_in[0][1394] , \round_in[0][1393] , \round_in[0][1392] ,
         \round_in[0][1391] , \round_in[0][1390] , \round_in[0][1389] ,
         \round_in[0][1388] , \round_in[0][1387] , \round_in[0][1386] ,
         \round_in[0][1385] , \round_in[0][1384] , \round_in[0][1383] ,
         \round_in[0][1382] , \round_in[0][1381] , \round_in[0][1380] ,
         \round_in[0][1379] , \round_in[0][1378] , \round_in[0][1377] ,
         \round_in[0][1376] , \round_in[0][1375] , \round_in[0][1374] ,
         \round_in[0][1373] , \round_in[0][1372] , \round_in[0][1371] ,
         \round_in[0][1370] , \round_in[0][1369] , \round_in[0][1368] ,
         \round_in[0][1367] , \round_in[0][1366] , \round_in[0][1365] ,
         \round_in[0][1364] , \round_in[0][1363] , \round_in[0][1362] ,
         \round_in[0][1361] , \round_in[0][1360] , \round_in[0][1359] ,
         \round_in[0][1358] , \round_in[0][1357] , \round_in[0][1356] ,
         \round_in[0][1355] , \round_in[0][1354] , \round_in[0][1353] ,
         \round_in[0][1352] , \round_in[0][1351] , \round_in[0][1350] ,
         \round_in[0][1349] , \round_in[0][1348] , \round_in[0][1347] ,
         \round_in[0][1346] , \round_in[0][1345] , \round_in[0][1344] ,
         \round_in[0][1343] , \round_in[0][1342] , \round_in[0][1341] ,
         \round_in[0][1340] , \round_in[0][1339] , \round_in[0][1338] ,
         \round_in[0][1337] , \round_in[0][1336] , \round_in[0][1335] ,
         \round_in[0][1334] , \round_in[0][1333] , \round_in[0][1332] ,
         \round_in[0][1331] , \round_in[0][1330] , \round_in[0][1329] ,
         \round_in[0][1328] , \round_in[0][1327] , \round_in[0][1326] ,
         \round_in[0][1325] , \round_in[0][1324] , \round_in[0][1323] ,
         \round_in[0][1322] , \round_in[0][1321] , \round_in[0][1320] ,
         \round_in[0][1319] , \round_in[0][1318] , \round_in[0][1317] ,
         \round_in[0][1316] , \round_in[0][1315] , \round_in[0][1314] ,
         \round_in[0][1313] , \round_in[0][1312] , \round_in[0][1311] ,
         \round_in[0][1310] , \round_in[0][1309] , \round_in[0][1308] ,
         \round_in[0][1307] , \round_in[0][1306] , \round_in[0][1305] ,
         \round_in[0][1304] , \round_in[0][1303] , \round_in[0][1302] ,
         \round_in[0][1301] , \round_in[0][1300] , \round_in[0][1299] ,
         \round_in[0][1298] , \round_in[0][1297] , \round_in[0][1296] ,
         \round_in[0][1295] , \round_in[0][1294] , \round_in[0][1293] ,
         \round_in[0][1292] , \round_in[0][1291] , \round_in[0][1290] ,
         \round_in[0][1289] , \round_in[0][1288] , \round_in[0][1287] ,
         \round_in[0][1286] , \round_in[0][1285] , \round_in[0][1284] ,
         \round_in[0][1283] , \round_in[0][1282] , \round_in[0][1281] ,
         \round_in[0][1280] , \round_in[0][1279] , \round_in[0][1278] ,
         \round_in[0][1277] , \round_in[0][1276] , \round_in[0][1275] ,
         \round_in[0][1274] , \round_in[0][1273] , \round_in[0][1272] ,
         \round_in[0][1271] , \round_in[0][1270] , \round_in[0][1269] ,
         \round_in[0][1268] , \round_in[0][1267] , \round_in[0][1266] ,
         \round_in[0][1265] , \round_in[0][1264] , \round_in[0][1263] ,
         \round_in[0][1262] , \round_in[0][1261] , \round_in[0][1260] ,
         \round_in[0][1259] , \round_in[0][1258] , \round_in[0][1257] ,
         \round_in[0][1256] , \round_in[0][1255] , \round_in[0][1254] ,
         \round_in[0][1253] , \round_in[0][1252] , \round_in[0][1251] ,
         \round_in[0][1250] , \round_in[0][1249] , \round_in[0][1248] ,
         \round_in[0][1247] , \round_in[0][1246] , \round_in[0][1245] ,
         \round_in[0][1244] , \round_in[0][1243] , \round_in[0][1242] ,
         \round_in[0][1241] , \round_in[0][1240] , \round_in[0][1239] ,
         \round_in[0][1238] , \round_in[0][1237] , \round_in[0][1236] ,
         \round_in[0][1235] , \round_in[0][1234] , \round_in[0][1233] ,
         \round_in[0][1232] , \round_in[0][1231] , \round_in[0][1230] ,
         \round_in[0][1229] , \round_in[0][1228] , \round_in[0][1227] ,
         \round_in[0][1226] , \round_in[0][1225] , \round_in[0][1224] ,
         \round_in[0][1223] , \round_in[0][1222] , \round_in[0][1221] ,
         \round_in[0][1220] , \round_in[0][1219] , \round_in[0][1218] ,
         \round_in[0][1217] , \round_in[0][1216] , \round_in[0][1215] ,
         \round_in[0][1214] , \round_in[0][1213] , \round_in[0][1212] ,
         \round_in[0][1211] , \round_in[0][1210] , \round_in[0][1209] ,
         \round_in[0][1208] , \round_in[0][1207] , \round_in[0][1206] ,
         \round_in[0][1205] , \round_in[0][1204] , \round_in[0][1203] ,
         \round_in[0][1202] , \round_in[0][1201] , \round_in[0][1200] ,
         \round_in[0][1199] , \round_in[0][1198] , \round_in[0][1197] ,
         \round_in[0][1196] , \round_in[0][1195] , \round_in[0][1194] ,
         \round_in[0][1193] , \round_in[0][1192] , \round_in[0][1191] ,
         \round_in[0][1190] , \round_in[0][1189] , \round_in[0][1188] ,
         \round_in[0][1187] , \round_in[0][1186] , \round_in[0][1185] ,
         \round_in[0][1184] , \round_in[0][1183] , \round_in[0][1182] ,
         \round_in[0][1181] , \round_in[0][1180] , \round_in[0][1179] ,
         \round_in[0][1178] , \round_in[0][1177] , \round_in[0][1176] ,
         \round_in[0][1175] , \round_in[0][1174] , \round_in[0][1173] ,
         \round_in[0][1172] , \round_in[0][1171] , \round_in[0][1170] ,
         \round_in[0][1169] , \round_in[0][1168] , \round_in[0][1167] ,
         \round_in[0][1166] , \round_in[0][1165] , \round_in[0][1164] ,
         \round_in[0][1163] , \round_in[0][1162] , \round_in[0][1161] ,
         \round_in[0][1160] , \round_in[0][1159] , \round_in[0][1158] ,
         \round_in[0][1157] , \round_in[0][1156] , \round_in[0][1155] ,
         \round_in[0][1154] , \round_in[0][1153] , \round_in[0][1152] ,
         \round_in[0][1151] , \round_in[0][1150] , \round_in[0][1149] ,
         \round_in[0][1148] , \round_in[0][1147] , \round_in[0][1146] ,
         \round_in[0][1145] , \round_in[0][1144] , \round_in[0][1143] ,
         \round_in[0][1142] , \round_in[0][1141] , \round_in[0][1140] ,
         \round_in[0][1139] , \round_in[0][1138] , \round_in[0][1137] ,
         \round_in[0][1136] , \round_in[0][1135] , \round_in[0][1134] ,
         \round_in[0][1133] , \round_in[0][1132] , \round_in[0][1131] ,
         \round_in[0][1130] , \round_in[0][1129] , \round_in[0][1128] ,
         \round_in[0][1127] , \round_in[0][1126] , \round_in[0][1125] ,
         \round_in[0][1124] , \round_in[0][1123] , \round_in[0][1122] ,
         \round_in[0][1121] , \round_in[0][1120] , \round_in[0][1119] ,
         \round_in[0][1118] , \round_in[0][1117] , \round_in[0][1116] ,
         \round_in[0][1115] , \round_in[0][1114] , \round_in[0][1113] ,
         \round_in[0][1112] , \round_in[0][1111] , \round_in[0][1110] ,
         \round_in[0][1109] , \round_in[0][1108] , \round_in[0][1107] ,
         \round_in[0][1106] , \round_in[0][1105] , \round_in[0][1104] ,
         \round_in[0][1103] , \round_in[0][1102] , \round_in[0][1101] ,
         \round_in[0][1100] , \round_in[0][1099] , \round_in[0][1098] ,
         \round_in[0][1097] , \round_in[0][1096] , \round_in[0][1095] ,
         \round_in[0][1094] , \round_in[0][1093] , \round_in[0][1092] ,
         \round_in[0][1091] , \round_in[0][1090] , \round_in[0][1089] ,
         \round_in[0][1088] , \round_in[0][1087] , \round_in[0][1086] ,
         \round_in[0][1085] , \round_in[0][1084] , \round_in[0][1083] ,
         \round_in[0][1082] , \round_in[0][1081] , \round_in[0][1080] ,
         \round_in[0][1079] , \round_in[0][1078] , \round_in[0][1077] ,
         \round_in[0][1076] , \round_in[0][1075] , \round_in[0][1074] ,
         \round_in[0][1073] , \round_in[0][1072] , \round_in[0][1071] ,
         \round_in[0][1070] , \round_in[0][1069] , \round_in[0][1068] ,
         \round_in[0][1067] , \round_in[0][1066] , \round_in[0][1065] ,
         \round_in[0][1064] , \round_in[0][1063] , \round_in[0][1062] ,
         \round_in[0][1061] , \round_in[0][1060] , \round_in[0][1059] ,
         \round_in[0][1058] , \round_in[0][1057] , \round_in[0][1056] ,
         \round_in[0][1055] , \round_in[0][1054] , \round_in[0][1053] ,
         \round_in[0][1052] , \round_in[0][1051] , \round_in[0][1050] ,
         \round_in[0][1049] , \round_in[0][1048] , \round_in[0][1047] ,
         \round_in[0][1046] , \round_in[0][1045] , \round_in[0][1044] ,
         \round_in[0][1043] , \round_in[0][1042] , \round_in[0][1041] ,
         \round_in[0][1040] , \round_in[0][1039] , \round_in[0][1038] ,
         \round_in[0][1037] , \round_in[0][1036] , \round_in[0][1035] ,
         \round_in[0][1034] , \round_in[0][1033] , \round_in[0][1032] ,
         \round_in[0][1031] , \round_in[0][1030] , \round_in[0][1029] ,
         \round_in[0][1028] , \round_in[0][1027] , \round_in[0][1026] ,
         \round_in[0][1025] , \round_in[0][1024] , \round_in[0][1023] ,
         \round_in[0][1022] , \round_in[0][1021] , \round_in[0][1020] ,
         \round_in[0][1019] , \round_in[0][1018] , \round_in[0][1017] ,
         \round_in[0][1016] , \round_in[0][1015] , \round_in[0][1014] ,
         \round_in[0][1013] , \round_in[0][1012] , \round_in[0][1011] ,
         \round_in[0][1010] , \round_in[0][1009] , \round_in[0][1008] ,
         \round_in[0][1007] , \round_in[0][1006] , \round_in[0][1005] ,
         \round_in[0][1004] , \round_in[0][1003] , \round_in[0][1002] ,
         \round_in[0][1001] , \round_in[0][1000] , \round_in[0][999] ,
         \round_in[0][998] , \round_in[0][997] , \round_in[0][996] ,
         \round_in[0][995] , \round_in[0][994] , \round_in[0][993] ,
         \round_in[0][992] , \round_in[0][991] , \round_in[0][990] ,
         \round_in[0][989] , \round_in[0][988] , \round_in[0][987] ,
         \round_in[0][986] , \round_in[0][985] , \round_in[0][984] ,
         \round_in[0][983] , \round_in[0][982] , \round_in[0][981] ,
         \round_in[0][980] , \round_in[0][979] , \round_in[0][978] ,
         \round_in[0][977] , \round_in[0][976] , \round_in[0][975] ,
         \round_in[0][974] , \round_in[0][973] , \round_in[0][972] ,
         \round_in[0][971] , \round_in[0][970] , \round_in[0][969] ,
         \round_in[0][968] , \round_in[0][967] , \round_in[0][966] ,
         \round_in[0][965] , \round_in[0][964] , \round_in[0][963] ,
         \round_in[0][962] , \round_in[0][961] , \round_in[0][960] ,
         \round_in[0][959] , \round_in[0][958] , \round_in[0][957] ,
         \round_in[0][956] , \round_in[0][955] , \round_in[0][954] ,
         \round_in[0][953] , \round_in[0][952] , \round_in[0][951] ,
         \round_in[0][950] , \round_in[0][949] , \round_in[0][948] ,
         \round_in[0][947] , \round_in[0][946] , \round_in[0][945] ,
         \round_in[0][944] , \round_in[0][943] , \round_in[0][942] ,
         \round_in[0][941] , \round_in[0][940] , \round_in[0][939] ,
         \round_in[0][938] , \round_in[0][937] , \round_in[0][936] ,
         \round_in[0][935] , \round_in[0][934] , \round_in[0][933] ,
         \round_in[0][932] , \round_in[0][931] , \round_in[0][930] ,
         \round_in[0][929] , \round_in[0][928] , \round_in[0][927] ,
         \round_in[0][926] , \round_in[0][925] , \round_in[0][924] ,
         \round_in[0][923] , \round_in[0][922] , \round_in[0][921] ,
         \round_in[0][920] , \round_in[0][919] , \round_in[0][918] ,
         \round_in[0][917] , \round_in[0][916] , \round_in[0][915] ,
         \round_in[0][914] , \round_in[0][913] , \round_in[0][912] ,
         \round_in[0][911] , \round_in[0][910] , \round_in[0][909] ,
         \round_in[0][908] , \round_in[0][907] , \round_in[0][906] ,
         \round_in[0][905] , \round_in[0][904] , \round_in[0][903] ,
         \round_in[0][902] , \round_in[0][901] , \round_in[0][900] ,
         \round_in[0][899] , \round_in[0][898] , \round_in[0][897] ,
         \round_in[0][896] , \round_in[0][895] , \round_in[0][894] ,
         \round_in[0][893] , \round_in[0][892] , \round_in[0][891] ,
         \round_in[0][890] , \round_in[0][889] , \round_in[0][888] ,
         \round_in[0][887] , \round_in[0][886] , \round_in[0][885] ,
         \round_in[0][884] , \round_in[0][883] , \round_in[0][882] ,
         \round_in[0][881] , \round_in[0][880] , \round_in[0][879] ,
         \round_in[0][878] , \round_in[0][877] , \round_in[0][876] ,
         \round_in[0][875] , \round_in[0][874] , \round_in[0][873] ,
         \round_in[0][872] , \round_in[0][871] , \round_in[0][870] ,
         \round_in[0][869] , \round_in[0][868] , \round_in[0][867] ,
         \round_in[0][866] , \round_in[0][865] , \round_in[0][864] ,
         \round_in[0][863] , \round_in[0][862] , \round_in[0][861] ,
         \round_in[0][860] , \round_in[0][859] , \round_in[0][858] ,
         \round_in[0][857] , \round_in[0][856] , \round_in[0][855] ,
         \round_in[0][854] , \round_in[0][853] , \round_in[0][852] ,
         \round_in[0][851] , \round_in[0][850] , \round_in[0][849] ,
         \round_in[0][848] , \round_in[0][847] , \round_in[0][846] ,
         \round_in[0][845] , \round_in[0][844] , \round_in[0][843] ,
         \round_in[0][842] , \round_in[0][841] , \round_in[0][840] ,
         \round_in[0][839] , \round_in[0][838] , \round_in[0][837] ,
         \round_in[0][836] , \round_in[0][835] , \round_in[0][834] ,
         \round_in[0][833] , \round_in[0][832] , \round_in[0][831] ,
         \round_in[0][830] , \round_in[0][829] , \round_in[0][828] ,
         \round_in[0][827] , \round_in[0][826] , \round_in[0][825] ,
         \round_in[0][824] , \round_in[0][823] , \round_in[0][822] ,
         \round_in[0][821] , \round_in[0][820] , \round_in[0][819] ,
         \round_in[0][818] , \round_in[0][817] , \round_in[0][816] ,
         \round_in[0][815] , \round_in[0][814] , \round_in[0][813] ,
         \round_in[0][812] , \round_in[0][811] , \round_in[0][810] ,
         \round_in[0][809] , \round_in[0][808] , \round_in[0][807] ,
         \round_in[0][806] , \round_in[0][805] , \round_in[0][804] ,
         \round_in[0][803] , \round_in[0][802] , \round_in[0][801] ,
         \round_in[0][800] , \round_in[0][799] , \round_in[0][798] ,
         \round_in[0][797] , \round_in[0][796] , \round_in[0][795] ,
         \round_in[0][794] , \round_in[0][793] , \round_in[0][792] ,
         \round_in[0][791] , \round_in[0][790] , \round_in[0][789] ,
         \round_in[0][788] , \round_in[0][787] , \round_in[0][786] ,
         \round_in[0][785] , \round_in[0][784] , \round_in[0][783] ,
         \round_in[0][782] , \round_in[0][781] , \round_in[0][780] ,
         \round_in[0][779] , \round_in[0][778] , \round_in[0][777] ,
         \round_in[0][776] , \round_in[0][775] , \round_in[0][774] ,
         \round_in[0][773] , \round_in[0][772] , \round_in[0][771] ,
         \round_in[0][770] , \round_in[0][769] , \round_in[0][768] ,
         \round_in[0][767] , \round_in[0][766] , \round_in[0][765] ,
         \round_in[0][764] , \round_in[0][763] , \round_in[0][762] ,
         \round_in[0][761] , \round_in[0][760] , \round_in[0][759] ,
         \round_in[0][758] , \round_in[0][757] , \round_in[0][756] ,
         \round_in[0][755] , \round_in[0][754] , \round_in[0][753] ,
         \round_in[0][752] , \round_in[0][751] , \round_in[0][750] ,
         \round_in[0][749] , \round_in[0][748] , \round_in[0][747] ,
         \round_in[0][746] , \round_in[0][745] , \round_in[0][744] ,
         \round_in[0][743] , \round_in[0][742] , \round_in[0][741] ,
         \round_in[0][740] , \round_in[0][739] , \round_in[0][738] ,
         \round_in[0][737] , \round_in[0][736] , \round_in[0][735] ,
         \round_in[0][734] , \round_in[0][733] , \round_in[0][732] ,
         \round_in[0][731] , \round_in[0][730] , \round_in[0][729] ,
         \round_in[0][728] , \round_in[0][727] , \round_in[0][726] ,
         \round_in[0][725] , \round_in[0][724] , \round_in[0][723] ,
         \round_in[0][722] , \round_in[0][721] , \round_in[0][720] ,
         \round_in[0][719] , \round_in[0][718] , \round_in[0][717] ,
         \round_in[0][716] , \round_in[0][715] , \round_in[0][714] ,
         \round_in[0][713] , \round_in[0][712] , \round_in[0][711] ,
         \round_in[0][710] , \round_in[0][709] , \round_in[0][708] ,
         \round_in[0][707] , \round_in[0][706] , \round_in[0][705] ,
         \round_in[0][704] , \round_in[0][703] , \round_in[0][702] ,
         \round_in[0][701] , \round_in[0][700] , \round_in[0][699] ,
         \round_in[0][698] , \round_in[0][697] , \round_in[0][696] ,
         \round_in[0][695] , \round_in[0][694] , \round_in[0][693] ,
         \round_in[0][692] , \round_in[0][691] , \round_in[0][690] ,
         \round_in[0][689] , \round_in[0][688] , \round_in[0][687] ,
         \round_in[0][686] , \round_in[0][685] , \round_in[0][684] ,
         \round_in[0][683] , \round_in[0][682] , \round_in[0][681] ,
         \round_in[0][680] , \round_in[0][679] , \round_in[0][678] ,
         \round_in[0][677] , \round_in[0][676] , \round_in[0][675] ,
         \round_in[0][674] , \round_in[0][673] , \round_in[0][672] ,
         \round_in[0][671] , \round_in[0][670] , \round_in[0][669] ,
         \round_in[0][668] , \round_in[0][667] , \round_in[0][666] ,
         \round_in[0][665] , \round_in[0][664] , \round_in[0][663] ,
         \round_in[0][662] , \round_in[0][661] , \round_in[0][660] ,
         \round_in[0][659] , \round_in[0][658] , \round_in[0][657] ,
         \round_in[0][656] , \round_in[0][655] , \round_in[0][654] ,
         \round_in[0][653] , \round_in[0][652] , \round_in[0][651] ,
         \round_in[0][650] , \round_in[0][649] , \round_in[0][648] ,
         \round_in[0][647] , \round_in[0][646] , \round_in[0][645] ,
         \round_in[0][644] , \round_in[0][643] , \round_in[0][642] ,
         \round_in[0][641] , \round_in[0][640] , \round_in[0][639] ,
         \round_in[0][638] , \round_in[0][637] , \round_in[0][636] ,
         \round_in[0][635] , \round_in[0][634] , \round_in[0][633] ,
         \round_in[0][632] , \round_in[0][631] , \round_in[0][630] ,
         \round_in[0][629] , \round_in[0][628] , \round_in[0][627] ,
         \round_in[0][626] , \round_in[0][625] , \round_in[0][624] ,
         \round_in[0][623] , \round_in[0][622] , \round_in[0][621] ,
         \round_in[0][620] , \round_in[0][619] , \round_in[0][618] ,
         \round_in[0][617] , \round_in[0][616] , \round_in[0][615] ,
         \round_in[0][614] , \round_in[0][613] , \round_in[0][612] ,
         \round_in[0][611] , \round_in[0][610] , \round_in[0][609] ,
         \round_in[0][608] , \round_in[0][607] , \round_in[0][606] ,
         \round_in[0][605] , \round_in[0][604] , \round_in[0][603] ,
         \round_in[0][602] , \round_in[0][601] , \round_in[0][600] ,
         \round_in[0][599] , \round_in[0][598] , \round_in[0][597] ,
         \round_in[0][596] , \round_in[0][595] , \round_in[0][594] ,
         \round_in[0][593] , \round_in[0][592] , \round_in[0][591] ,
         \round_in[0][590] , \round_in[0][589] , \round_in[0][588] ,
         \round_in[0][587] , \round_in[0][586] , \round_in[0][585] ,
         \round_in[0][584] , \round_in[0][583] , \round_in[0][582] ,
         \round_in[0][581] , \round_in[0][580] , \round_in[0][579] ,
         \round_in[0][578] , \round_in[0][577] , \round_in[0][576] ,
         \round_in[0][575] , \round_in[0][574] , \round_in[0][573] ,
         \round_in[0][572] , \round_in[0][571] , \round_in[0][570] ,
         \round_in[0][569] , \round_in[0][568] , \round_in[0][567] ,
         \round_in[0][566] , \round_in[0][565] , \round_in[0][564] ,
         \round_in[0][563] , \round_in[0][562] , \round_in[0][561] ,
         \round_in[0][560] , \round_in[0][559] , \round_in[0][558] ,
         \round_in[0][557] , \round_in[0][556] , \round_in[0][555] ,
         \round_in[0][554] , \round_in[0][553] , \round_in[0][552] ,
         \round_in[0][551] , \round_in[0][550] , \round_in[0][549] ,
         \round_in[0][548] , \round_in[0][547] , \round_in[0][546] ,
         \round_in[0][545] , \round_in[0][544] , \round_in[0][543] ,
         \round_in[0][542] , \round_in[0][541] , \round_in[0][540] ,
         \round_in[0][539] , \round_in[0][538] , \round_in[0][537] ,
         \round_in[0][536] , \round_in[0][535] , \round_in[0][534] ,
         \round_in[0][533] , \round_in[0][532] , \round_in[0][531] ,
         \round_in[0][530] , \round_in[0][529] , \round_in[0][528] ,
         \round_in[0][527] , \round_in[0][526] , \round_in[0][525] ,
         \round_in[0][524] , \round_in[0][523] , \round_in[0][522] ,
         \round_in[0][521] , \round_in[0][520] , \round_in[0][519] ,
         \round_in[0][518] , \round_in[0][517] , \round_in[0][516] ,
         \round_in[0][515] , \round_in[0][514] , \round_in[0][513] ,
         \round_in[0][512] , \round_in[0][511] , \round_in[0][510] ,
         \round_in[0][509] , \round_in[0][508] , \round_in[0][507] ,
         \round_in[0][506] , \round_in[0][505] , \round_in[0][504] ,
         \round_in[0][503] , \round_in[0][502] , \round_in[0][501] ,
         \round_in[0][500] , \round_in[0][499] , \round_in[0][498] ,
         \round_in[0][497] , \round_in[0][496] , \round_in[0][495] ,
         \round_in[0][494] , \round_in[0][493] , \round_in[0][492] ,
         \round_in[0][491] , \round_in[0][490] , \round_in[0][489] ,
         \round_in[0][488] , \round_in[0][487] , \round_in[0][486] ,
         \round_in[0][485] , \round_in[0][484] , \round_in[0][483] ,
         \round_in[0][482] , \round_in[0][481] , \round_in[0][480] ,
         \round_in[0][479] , \round_in[0][478] , \round_in[0][477] ,
         \round_in[0][476] , \round_in[0][475] , \round_in[0][474] ,
         \round_in[0][473] , \round_in[0][472] , \round_in[0][471] ,
         \round_in[0][470] , \round_in[0][469] , \round_in[0][468] ,
         \round_in[0][467] , \round_in[0][466] , \round_in[0][465] ,
         \round_in[0][464] , \round_in[0][463] , \round_in[0][462] ,
         \round_in[0][461] , \round_in[0][460] , \round_in[0][459] ,
         \round_in[0][458] , \round_in[0][457] , \round_in[0][456] ,
         \round_in[0][455] , \round_in[0][454] , \round_in[0][453] ,
         \round_in[0][452] , \round_in[0][451] , \round_in[0][450] ,
         \round_in[0][449] , \round_in[0][448] , \round_in[0][447] ,
         \round_in[0][446] , \round_in[0][445] , \round_in[0][444] ,
         \round_in[0][443] , \round_in[0][442] , \round_in[0][441] ,
         \round_in[0][440] , \round_in[0][439] , \round_in[0][438] ,
         \round_in[0][437] , \round_in[0][436] , \round_in[0][435] ,
         \round_in[0][434] , \round_in[0][433] , \round_in[0][432] ,
         \round_in[0][431] , \round_in[0][430] , \round_in[0][429] ,
         \round_in[0][428] , \round_in[0][427] , \round_in[0][426] ,
         \round_in[0][425] , \round_in[0][424] , \round_in[0][423] ,
         \round_in[0][422] , \round_in[0][421] , \round_in[0][420] ,
         \round_in[0][419] , \round_in[0][418] , \round_in[0][417] ,
         \round_in[0][416] , \round_in[0][415] , \round_in[0][414] ,
         \round_in[0][413] , \round_in[0][412] , \round_in[0][411] ,
         \round_in[0][410] , \round_in[0][409] , \round_in[0][408] ,
         \round_in[0][407] , \round_in[0][406] , \round_in[0][405] ,
         \round_in[0][404] , \round_in[0][403] , \round_in[0][402] ,
         \round_in[0][401] , \round_in[0][400] , \round_in[0][399] ,
         \round_in[0][398] , \round_in[0][397] , \round_in[0][396] ,
         \round_in[0][395] , \round_in[0][394] , \round_in[0][393] ,
         \round_in[0][392] , \round_in[0][391] , \round_in[0][390] ,
         \round_in[0][389] , \round_in[0][388] , \round_in[0][387] ,
         \round_in[0][386] , \round_in[0][385] , \round_in[0][384] ,
         \round_in[0][383] , \round_in[0][382] , \round_in[0][381] ,
         \round_in[0][380] , \round_in[0][379] , \round_in[0][378] ,
         \round_in[0][377] , \round_in[0][376] , \round_in[0][375] ,
         \round_in[0][374] , \round_in[0][373] , \round_in[0][372] ,
         \round_in[0][371] , \round_in[0][370] , \round_in[0][369] ,
         \round_in[0][368] , \round_in[0][367] , \round_in[0][366] ,
         \round_in[0][365] , \round_in[0][364] , \round_in[0][363] ,
         \round_in[0][362] , \round_in[0][361] , \round_in[0][360] ,
         \round_in[0][359] , \round_in[0][358] , \round_in[0][357] ,
         \round_in[0][356] , \round_in[0][355] , \round_in[0][354] ,
         \round_in[0][353] , \round_in[0][352] , \round_in[0][351] ,
         \round_in[0][350] , \round_in[0][349] , \round_in[0][348] ,
         \round_in[0][347] , \round_in[0][346] , \round_in[0][345] ,
         \round_in[0][344] , \round_in[0][343] , \round_in[0][342] ,
         \round_in[0][341] , \round_in[0][340] , \round_in[0][339] ,
         \round_in[0][338] , \round_in[0][337] , \round_in[0][336] ,
         \round_in[0][335] , \round_in[0][334] , \round_in[0][333] ,
         \round_in[0][332] , \round_in[0][331] , \round_in[0][330] ,
         \round_in[0][329] , \round_in[0][328] , \round_in[0][327] ,
         \round_in[0][326] , \round_in[0][325] , \round_in[0][324] ,
         \round_in[0][323] , \round_in[0][322] , \round_in[0][321] ,
         \round_in[0][320] , \round_in[0][319] , \round_in[0][318] ,
         \round_in[0][317] , \round_in[0][316] , \round_in[0][315] ,
         \round_in[0][314] , \round_in[0][313] , \round_in[0][312] ,
         \round_in[0][311] , \round_in[0][310] , \round_in[0][309] ,
         \round_in[0][308] , \round_in[0][307] , \round_in[0][306] ,
         \round_in[0][305] , \round_in[0][304] , \round_in[0][303] ,
         \round_in[0][302] , \round_in[0][301] , \round_in[0][300] ,
         \round_in[0][299] , \round_in[0][298] , \round_in[0][297] ,
         \round_in[0][296] , \round_in[0][295] , \round_in[0][294] ,
         \round_in[0][293] , \round_in[0][292] , \round_in[0][291] ,
         \round_in[0][290] , \round_in[0][289] , \round_in[0][288] ,
         \round_in[0][287] , \round_in[0][286] , \round_in[0][285] ,
         \round_in[0][284] , \round_in[0][283] , \round_in[0][282] ,
         \round_in[0][281] , \round_in[0][280] , \round_in[0][279] ,
         \round_in[0][278] , \round_in[0][277] , \round_in[0][276] ,
         \round_in[0][275] , \round_in[0][274] , \round_in[0][273] ,
         \round_in[0][272] , \round_in[0][271] , \round_in[0][270] ,
         \round_in[0][269] , \round_in[0][268] , \round_in[0][267] ,
         \round_in[0][266] , \round_in[0][265] , \round_in[0][264] ,
         \round_in[0][263] , \round_in[0][262] , \round_in[0][261] ,
         \round_in[0][260] , \round_in[0][259] , \round_in[0][258] ,
         \round_in[0][257] , \round_in[0][256] , \round_in[0][255] ,
         \round_in[0][254] , \round_in[0][253] , \round_in[0][252] ,
         \round_in[0][251] , \round_in[0][250] , \round_in[0][249] ,
         \round_in[0][248] , \round_in[0][247] , \round_in[0][246] ,
         \round_in[0][245] , \round_in[0][244] , \round_in[0][243] ,
         \round_in[0][242] , \round_in[0][241] , \round_in[0][240] ,
         \round_in[0][239] , \round_in[0][238] , \round_in[0][237] ,
         \round_in[0][236] , \round_in[0][235] , \round_in[0][234] ,
         \round_in[0][233] , \round_in[0][232] , \round_in[0][231] ,
         \round_in[0][230] , \round_in[0][229] , \round_in[0][228] ,
         \round_in[0][227] , \round_in[0][226] , \round_in[0][225] ,
         \round_in[0][224] , \round_in[0][223] , \round_in[0][222] ,
         \round_in[0][221] , \round_in[0][220] , \round_in[0][219] ,
         \round_in[0][218] , \round_in[0][217] , \round_in[0][216] ,
         \round_in[0][215] , \round_in[0][214] , \round_in[0][213] ,
         \round_in[0][212] , \round_in[0][211] , \round_in[0][210] ,
         \round_in[0][209] , \round_in[0][208] , \round_in[0][207] ,
         \round_in[0][206] , \round_in[0][205] , \round_in[0][204] ,
         \round_in[0][203] , \round_in[0][202] , \round_in[0][201] ,
         \round_in[0][200] , \round_in[0][199] , \round_in[0][198] ,
         \round_in[0][197] , \round_in[0][196] , \round_in[0][195] ,
         \round_in[0][194] , \round_in[0][193] , \round_in[0][192] ,
         \round_in[0][191] , \round_in[0][190] , \round_in[0][189] ,
         \round_in[0][188] , \round_in[0][187] , \round_in[0][186] ,
         \round_in[0][185] , \round_in[0][184] , \round_in[0][183] ,
         \round_in[0][182] , \round_in[0][181] , \round_in[0][180] ,
         \round_in[0][179] , \round_in[0][178] , \round_in[0][177] ,
         \round_in[0][176] , \round_in[0][175] , \round_in[0][174] ,
         \round_in[0][173] , \round_in[0][172] , \round_in[0][171] ,
         \round_in[0][170] , \round_in[0][169] , \round_in[0][168] ,
         \round_in[0][167] , \round_in[0][166] , \round_in[0][165] ,
         \round_in[0][164] , \round_in[0][163] , \round_in[0][162] ,
         \round_in[0][161] , \round_in[0][160] , \round_in[0][159] ,
         \round_in[0][158] , \round_in[0][157] , \round_in[0][156] ,
         \round_in[0][155] , \round_in[0][154] , \round_in[0][153] ,
         \round_in[0][152] , \round_in[0][151] , \round_in[0][150] ,
         \round_in[0][149] , \round_in[0][148] , \round_in[0][147] ,
         \round_in[0][146] , \round_in[0][145] , \round_in[0][144] ,
         \round_in[0][143] , \round_in[0][142] , \round_in[0][141] ,
         \round_in[0][140] , \round_in[0][139] , \round_in[0][138] ,
         \round_in[0][137] , \round_in[0][136] , \round_in[0][135] ,
         \round_in[0][134] , \round_in[0][133] , \round_in[0][132] ,
         \round_in[0][131] , \round_in[0][130] , \round_in[0][129] ,
         \round_in[0][128] , \round_in[0][127] , \round_in[0][126] ,
         \round_in[0][125] , \round_in[0][124] , \round_in[0][123] ,
         \round_in[0][122] , \round_in[0][121] , \round_in[0][120] ,
         \round_in[0][119] , \round_in[0][118] , \round_in[0][117] ,
         \round_in[0][116] , \round_in[0][115] , \round_in[0][114] ,
         \round_in[0][113] , \round_in[0][112] , \round_in[0][111] ,
         \round_in[0][110] , \round_in[0][109] , \round_in[0][108] ,
         \round_in[0][107] , \round_in[0][106] , \round_in[0][105] ,
         \round_in[0][104] , \round_in[0][103] , \round_in[0][102] ,
         \round_in[0][101] , \round_in[0][100] , \round_in[0][99] ,
         \round_in[0][98] , \round_in[0][97] , \round_in[0][96] ,
         \round_in[0][95] , \round_in[0][94] , \round_in[0][93] ,
         \round_in[0][92] , \round_in[0][91] , \round_in[0][90] ,
         \round_in[0][89] , \round_in[0][88] , \round_in[0][87] ,
         \round_in[0][86] , \round_in[0][85] , \round_in[0][84] ,
         \round_in[0][83] , \round_in[0][82] , \round_in[0][81] ,
         \round_in[0][80] , \round_in[0][79] , \round_in[0][78] ,
         \round_in[0][77] , \round_in[0][76] , \round_in[0][75] ,
         \round_in[0][74] , \round_in[0][73] , \round_in[0][72] ,
         \round_in[0][71] , \round_in[0][70] , \round_in[0][69] ,
         \round_in[0][68] , \round_in[0][67] , \round_in[0][66] ,
         \round_in[0][65] , \round_in[0][64] , \round_in[0][63] ,
         \round_in[0][62] , \round_in[0][61] , \round_in[0][60] ,
         \round_in[0][59] , \round_in[0][58] , \round_in[0][57] ,
         \round_in[0][56] , \round_in[0][55] , \round_in[0][54] ,
         \round_in[0][53] , \round_in[0][52] , \round_in[0][51] ,
         \round_in[0][50] , \round_in[0][49] , \round_in[0][48] ,
         \round_in[0][47] , \round_in[0][46] , \round_in[0][45] ,
         \round_in[0][44] , \round_in[0][43] , \round_in[0][42] ,
         \round_in[0][41] , \round_in[0][40] , \round_in[0][39] ,
         \round_in[0][38] , \round_in[0][37] , \round_in[0][36] ,
         \round_in[0][35] , \round_in[0][34] , \round_in[0][33] ,
         \round_in[0][32] , \round_in[0][31] , \round_in[0][30] ,
         \round_in[0][29] , \round_in[0][28] , \round_in[0][27] ,
         \round_in[0][26] , \round_in[0][25] , \round_in[0][24] ,
         \round_in[0][23] , \round_in[0][22] , \round_in[0][21] ,
         \round_in[0][20] , \round_in[0][19] , \round_in[0][18] ,
         \round_in[0][17] , \round_in[0][16] , \round_in[0][15] ,
         \round_in[0][14] , \round_in[0][13] , \round_in[0][12] ,
         \round_in[0][11] , \round_in[0][10] , \round_in[0][9] ,
         \round_in[0][8] , \round_in[0][7] , \round_in[0][6] ,
         \round_in[0][5] , \round_in[0][4] , \round_in[0][3] ,
         \round_in[0][2] , \round_in[0][1] , \round_in[0][0] , \rc[1][63] ,
         \rc[1][31] , \rc[1][15] , \rc[1][7] , \rc[1][3] , \rc[1][1] ,
         \rc[0][0] , \RCONST[0].rconst_/N67 , \RCONST[0].rconst_/N57 ,
         \RCONST[0].rconst_/N48 , \RCONST[0].rconst_/N37 ,
         \RCONST[0].rconst_/N28 , \RCONST[0].rconst_/N18 ,
         \RCONST[1].rconst_/N10 , n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968;
  wire   [11:0] rc_i;
  wire   [1599:0] round_reg;

  round_0 \ROUND[0].round_  ( .in({\round_in[0][1599] , \round_in[0][1598] , 
        \round_in[0][1597] , \round_in[0][1596] , \round_in[0][1595] , 
        \round_in[0][1594] , \round_in[0][1593] , \round_in[0][1592] , 
        \round_in[0][1591] , \round_in[0][1590] , \round_in[0][1589] , 
        \round_in[0][1588] , \round_in[0][1587] , \round_in[0][1586] , 
        \round_in[0][1585] , \round_in[0][1584] , \round_in[0][1583] , 
        \round_in[0][1582] , \round_in[0][1581] , \round_in[0][1580] , 
        \round_in[0][1579] , \round_in[0][1578] , \round_in[0][1577] , 
        \round_in[0][1576] , \round_in[0][1575] , \round_in[0][1574] , 
        \round_in[0][1573] , \round_in[0][1572] , \round_in[0][1571] , 
        \round_in[0][1570] , \round_in[0][1569] , \round_in[0][1568] , 
        \round_in[0][1567] , \round_in[0][1566] , \round_in[0][1565] , 
        \round_in[0][1564] , \round_in[0][1563] , \round_in[0][1562] , 
        \round_in[0][1561] , \round_in[0][1560] , \round_in[0][1559] , 
        \round_in[0][1558] , \round_in[0][1557] , \round_in[0][1556] , 
        \round_in[0][1555] , \round_in[0][1554] , \round_in[0][1553] , 
        \round_in[0][1552] , \round_in[0][1551] , \round_in[0][1550] , 
        \round_in[0][1549] , \round_in[0][1548] , \round_in[0][1547] , 
        \round_in[0][1546] , \round_in[0][1545] , \round_in[0][1544] , 
        \round_in[0][1543] , \round_in[0][1542] , \round_in[0][1541] , 
        \round_in[0][1540] , \round_in[0][1539] , \round_in[0][1538] , 
        \round_in[0][1537] , \round_in[0][1536] , \round_in[0][1535] , 
        \round_in[0][1534] , \round_in[0][1533] , \round_in[0][1532] , 
        \round_in[0][1531] , \round_in[0][1530] , \round_in[0][1529] , 
        \round_in[0][1528] , \round_in[0][1527] , \round_in[0][1526] , 
        \round_in[0][1525] , \round_in[0][1524] , \round_in[0][1523] , 
        \round_in[0][1522] , \round_in[0][1521] , \round_in[0][1520] , 
        \round_in[0][1519] , \round_in[0][1518] , \round_in[0][1517] , 
        \round_in[0][1516] , \round_in[0][1515] , \round_in[0][1514] , 
        \round_in[0][1513] , \round_in[0][1512] , \round_in[0][1511] , 
        \round_in[0][1510] , \round_in[0][1509] , \round_in[0][1508] , 
        \round_in[0][1507] , \round_in[0][1506] , \round_in[0][1505] , 
        \round_in[0][1504] , \round_in[0][1503] , \round_in[0][1502] , 
        \round_in[0][1501] , \round_in[0][1500] , \round_in[0][1499] , 
        \round_in[0][1498] , \round_in[0][1497] , \round_in[0][1496] , 
        \round_in[0][1495] , \round_in[0][1494] , \round_in[0][1493] , 
        \round_in[0][1492] , \round_in[0][1491] , \round_in[0][1490] , 
        \round_in[0][1489] , \round_in[0][1488] , \round_in[0][1487] , 
        \round_in[0][1486] , \round_in[0][1485] , \round_in[0][1484] , 
        \round_in[0][1483] , \round_in[0][1482] , \round_in[0][1481] , 
        \round_in[0][1480] , \round_in[0][1479] , \round_in[0][1478] , 
        \round_in[0][1477] , \round_in[0][1476] , \round_in[0][1475] , 
        \round_in[0][1474] , \round_in[0][1473] , \round_in[0][1472] , 
        \round_in[0][1471] , \round_in[0][1470] , \round_in[0][1469] , 
        \round_in[0][1468] , \round_in[0][1467] , \round_in[0][1466] , 
        \round_in[0][1465] , \round_in[0][1464] , \round_in[0][1463] , 
        \round_in[0][1462] , \round_in[0][1461] , \round_in[0][1460] , 
        \round_in[0][1459] , \round_in[0][1458] , \round_in[0][1457] , 
        \round_in[0][1456] , \round_in[0][1455] , \round_in[0][1454] , 
        \round_in[0][1453] , \round_in[0][1452] , \round_in[0][1451] , 
        \round_in[0][1450] , \round_in[0][1449] , \round_in[0][1448] , 
        \round_in[0][1447] , \round_in[0][1446] , \round_in[0][1445] , 
        \round_in[0][1444] , \round_in[0][1443] , \round_in[0][1442] , 
        \round_in[0][1441] , \round_in[0][1440] , \round_in[0][1439] , 
        \round_in[0][1438] , \round_in[0][1437] , \round_in[0][1436] , 
        \round_in[0][1435] , \round_in[0][1434] , \round_in[0][1433] , 
        \round_in[0][1432] , \round_in[0][1431] , \round_in[0][1430] , 
        \round_in[0][1429] , \round_in[0][1428] , \round_in[0][1427] , 
        \round_in[0][1426] , \round_in[0][1425] , \round_in[0][1424] , 
        \round_in[0][1423] , \round_in[0][1422] , \round_in[0][1421] , 
        \round_in[0][1420] , \round_in[0][1419] , \round_in[0][1418] , 
        \round_in[0][1417] , \round_in[0][1416] , \round_in[0][1415] , 
        \round_in[0][1414] , \round_in[0][1413] , \round_in[0][1412] , 
        \round_in[0][1411] , \round_in[0][1410] , \round_in[0][1409] , 
        \round_in[0][1408] , \round_in[0][1407] , \round_in[0][1406] , 
        \round_in[0][1405] , \round_in[0][1404] , \round_in[0][1403] , 
        \round_in[0][1402] , \round_in[0][1401] , \round_in[0][1400] , 
        \round_in[0][1399] , \round_in[0][1398] , \round_in[0][1397] , 
        \round_in[0][1396] , \round_in[0][1395] , \round_in[0][1394] , 
        \round_in[0][1393] , \round_in[0][1392] , \round_in[0][1391] , 
        \round_in[0][1390] , \round_in[0][1389] , \round_in[0][1388] , 
        \round_in[0][1387] , \round_in[0][1386] , \round_in[0][1385] , 
        \round_in[0][1384] , \round_in[0][1383] , \round_in[0][1382] , 
        \round_in[0][1381] , \round_in[0][1380] , \round_in[0][1379] , 
        \round_in[0][1378] , \round_in[0][1377] , \round_in[0][1376] , 
        \round_in[0][1375] , \round_in[0][1374] , \round_in[0][1373] , 
        \round_in[0][1372] , \round_in[0][1371] , \round_in[0][1370] , 
        \round_in[0][1369] , \round_in[0][1368] , \round_in[0][1367] , 
        \round_in[0][1366] , \round_in[0][1365] , \round_in[0][1364] , 
        \round_in[0][1363] , \round_in[0][1362] , \round_in[0][1361] , 
        \round_in[0][1360] , \round_in[0][1359] , \round_in[0][1358] , 
        \round_in[0][1357] , \round_in[0][1356] , \round_in[0][1355] , 
        \round_in[0][1354] , \round_in[0][1353] , \round_in[0][1352] , 
        \round_in[0][1351] , \round_in[0][1350] , \round_in[0][1349] , 
        \round_in[0][1348] , \round_in[0][1347] , \round_in[0][1346] , 
        \round_in[0][1345] , \round_in[0][1344] , \round_in[0][1343] , 
        \round_in[0][1342] , \round_in[0][1341] , \round_in[0][1340] , 
        \round_in[0][1339] , \round_in[0][1338] , \round_in[0][1337] , 
        \round_in[0][1336] , \round_in[0][1335] , \round_in[0][1334] , 
        \round_in[0][1333] , \round_in[0][1332] , \round_in[0][1331] , 
        \round_in[0][1330] , \round_in[0][1329] , \round_in[0][1328] , 
        \round_in[0][1327] , \round_in[0][1326] , \round_in[0][1325] , 
        \round_in[0][1324] , \round_in[0][1323] , \round_in[0][1322] , 
        \round_in[0][1321] , \round_in[0][1320] , \round_in[0][1319] , 
        \round_in[0][1318] , \round_in[0][1317] , \round_in[0][1316] , 
        \round_in[0][1315] , \round_in[0][1314] , \round_in[0][1313] , 
        \round_in[0][1312] , \round_in[0][1311] , \round_in[0][1310] , 
        \round_in[0][1309] , \round_in[0][1308] , \round_in[0][1307] , 
        \round_in[0][1306] , \round_in[0][1305] , \round_in[0][1304] , 
        \round_in[0][1303] , \round_in[0][1302] , \round_in[0][1301] , 
        \round_in[0][1300] , \round_in[0][1299] , \round_in[0][1298] , 
        \round_in[0][1297] , \round_in[0][1296] , \round_in[0][1295] , 
        \round_in[0][1294] , \round_in[0][1293] , \round_in[0][1292] , 
        \round_in[0][1291] , \round_in[0][1290] , \round_in[0][1289] , 
        \round_in[0][1288] , \round_in[0][1287] , \round_in[0][1286] , 
        \round_in[0][1285] , \round_in[0][1284] , \round_in[0][1283] , 
        \round_in[0][1282] , \round_in[0][1281] , \round_in[0][1280] , 
        \round_in[0][1279] , \round_in[0][1278] , \round_in[0][1277] , 
        \round_in[0][1276] , \round_in[0][1275] , \round_in[0][1274] , 
        \round_in[0][1273] , \round_in[0][1272] , \round_in[0][1271] , 
        \round_in[0][1270] , \round_in[0][1269] , \round_in[0][1268] , 
        \round_in[0][1267] , \round_in[0][1266] , \round_in[0][1265] , 
        \round_in[0][1264] , \round_in[0][1263] , \round_in[0][1262] , 
        \round_in[0][1261] , \round_in[0][1260] , \round_in[0][1259] , 
        \round_in[0][1258] , \round_in[0][1257] , \round_in[0][1256] , 
        \round_in[0][1255] , \round_in[0][1254] , \round_in[0][1253] , 
        \round_in[0][1252] , \round_in[0][1251] , \round_in[0][1250] , 
        \round_in[0][1249] , \round_in[0][1248] , \round_in[0][1247] , 
        \round_in[0][1246] , \round_in[0][1245] , \round_in[0][1244] , 
        \round_in[0][1243] , \round_in[0][1242] , \round_in[0][1241] , 
        \round_in[0][1240] , \round_in[0][1239] , \round_in[0][1238] , 
        \round_in[0][1237] , \round_in[0][1236] , \round_in[0][1235] , 
        \round_in[0][1234] , \round_in[0][1233] , \round_in[0][1232] , 
        \round_in[0][1231] , \round_in[0][1230] , \round_in[0][1229] , 
        \round_in[0][1228] , \round_in[0][1227] , \round_in[0][1226] , 
        \round_in[0][1225] , \round_in[0][1224] , \round_in[0][1223] , 
        \round_in[0][1222] , \round_in[0][1221] , \round_in[0][1220] , 
        \round_in[0][1219] , \round_in[0][1218] , \round_in[0][1217] , 
        \round_in[0][1216] , \round_in[0][1215] , \round_in[0][1214] , 
        \round_in[0][1213] , \round_in[0][1212] , \round_in[0][1211] , 
        \round_in[0][1210] , \round_in[0][1209] , \round_in[0][1208] , 
        \round_in[0][1207] , \round_in[0][1206] , \round_in[0][1205] , 
        \round_in[0][1204] , \round_in[0][1203] , \round_in[0][1202] , 
        \round_in[0][1201] , \round_in[0][1200] , \round_in[0][1199] , 
        \round_in[0][1198] , \round_in[0][1197] , \round_in[0][1196] , 
        \round_in[0][1195] , \round_in[0][1194] , \round_in[0][1193] , 
        \round_in[0][1192] , \round_in[0][1191] , \round_in[0][1190] , 
        \round_in[0][1189] , \round_in[0][1188] , \round_in[0][1187] , 
        \round_in[0][1186] , \round_in[0][1185] , \round_in[0][1184] , 
        \round_in[0][1183] , \round_in[0][1182] , \round_in[0][1181] , 
        \round_in[0][1180] , \round_in[0][1179] , \round_in[0][1178] , 
        \round_in[0][1177] , \round_in[0][1176] , \round_in[0][1175] , 
        \round_in[0][1174] , \round_in[0][1173] , \round_in[0][1172] , 
        \round_in[0][1171] , \round_in[0][1170] , \round_in[0][1169] , 
        \round_in[0][1168] , \round_in[0][1167] , \round_in[0][1166] , 
        \round_in[0][1165] , \round_in[0][1164] , \round_in[0][1163] , 
        \round_in[0][1162] , \round_in[0][1161] , \round_in[0][1160] , 
        \round_in[0][1159] , \round_in[0][1158] , \round_in[0][1157] , 
        \round_in[0][1156] , \round_in[0][1155] , \round_in[0][1154] , 
        \round_in[0][1153] , \round_in[0][1152] , \round_in[0][1151] , 
        \round_in[0][1150] , \round_in[0][1149] , \round_in[0][1148] , 
        \round_in[0][1147] , \round_in[0][1146] , \round_in[0][1145] , 
        \round_in[0][1144] , \round_in[0][1143] , \round_in[0][1142] , 
        \round_in[0][1141] , \round_in[0][1140] , \round_in[0][1139] , 
        \round_in[0][1138] , \round_in[0][1137] , \round_in[0][1136] , 
        \round_in[0][1135] , \round_in[0][1134] , \round_in[0][1133] , 
        \round_in[0][1132] , \round_in[0][1131] , \round_in[0][1130] , 
        \round_in[0][1129] , \round_in[0][1128] , \round_in[0][1127] , 
        \round_in[0][1126] , \round_in[0][1125] , \round_in[0][1124] , 
        \round_in[0][1123] , \round_in[0][1122] , \round_in[0][1121] , 
        \round_in[0][1120] , \round_in[0][1119] , \round_in[0][1118] , 
        \round_in[0][1117] , \round_in[0][1116] , \round_in[0][1115] , 
        \round_in[0][1114] , \round_in[0][1113] , \round_in[0][1112] , 
        \round_in[0][1111] , \round_in[0][1110] , \round_in[0][1109] , 
        \round_in[0][1108] , \round_in[0][1107] , \round_in[0][1106] , 
        \round_in[0][1105] , \round_in[0][1104] , \round_in[0][1103] , 
        \round_in[0][1102] , \round_in[0][1101] , \round_in[0][1100] , 
        \round_in[0][1099] , \round_in[0][1098] , \round_in[0][1097] , 
        \round_in[0][1096] , \round_in[0][1095] , \round_in[0][1094] , 
        \round_in[0][1093] , \round_in[0][1092] , \round_in[0][1091] , 
        \round_in[0][1090] , \round_in[0][1089] , \round_in[0][1088] , 
        \round_in[0][1087] , \round_in[0][1086] , \round_in[0][1085] , 
        \round_in[0][1084] , \round_in[0][1083] , \round_in[0][1082] , 
        \round_in[0][1081] , \round_in[0][1080] , \round_in[0][1079] , 
        \round_in[0][1078] , \round_in[0][1077] , \round_in[0][1076] , 
        \round_in[0][1075] , \round_in[0][1074] , \round_in[0][1073] , 
        \round_in[0][1072] , \round_in[0][1071] , \round_in[0][1070] , 
        \round_in[0][1069] , \round_in[0][1068] , \round_in[0][1067] , 
        \round_in[0][1066] , \round_in[0][1065] , \round_in[0][1064] , 
        \round_in[0][1063] , \round_in[0][1062] , \round_in[0][1061] , 
        \round_in[0][1060] , \round_in[0][1059] , \round_in[0][1058] , 
        \round_in[0][1057] , \round_in[0][1056] , \round_in[0][1055] , 
        \round_in[0][1054] , \round_in[0][1053] , \round_in[0][1052] , 
        \round_in[0][1051] , \round_in[0][1050] , \round_in[0][1049] , 
        \round_in[0][1048] , \round_in[0][1047] , \round_in[0][1046] , 
        \round_in[0][1045] , \round_in[0][1044] , \round_in[0][1043] , 
        \round_in[0][1042] , \round_in[0][1041] , \round_in[0][1040] , 
        \round_in[0][1039] , \round_in[0][1038] , \round_in[0][1037] , 
        \round_in[0][1036] , \round_in[0][1035] , \round_in[0][1034] , 
        \round_in[0][1033] , \round_in[0][1032] , \round_in[0][1031] , 
        \round_in[0][1030] , \round_in[0][1029] , \round_in[0][1028] , 
        \round_in[0][1027] , \round_in[0][1026] , \round_in[0][1025] , 
        \round_in[0][1024] , \round_in[0][1023] , \round_in[0][1022] , 
        \round_in[0][1021] , \round_in[0][1020] , \round_in[0][1019] , 
        \round_in[0][1018] , \round_in[0][1017] , \round_in[0][1016] , 
        \round_in[0][1015] , \round_in[0][1014] , \round_in[0][1013] , 
        \round_in[0][1012] , \round_in[0][1011] , \round_in[0][1010] , 
        \round_in[0][1009] , \round_in[0][1008] , \round_in[0][1007] , 
        \round_in[0][1006] , \round_in[0][1005] , \round_in[0][1004] , 
        \round_in[0][1003] , \round_in[0][1002] , \round_in[0][1001] , 
        \round_in[0][1000] , \round_in[0][999] , \round_in[0][998] , 
        \round_in[0][997] , \round_in[0][996] , \round_in[0][995] , 
        \round_in[0][994] , \round_in[0][993] , \round_in[0][992] , 
        \round_in[0][991] , \round_in[0][990] , \round_in[0][989] , 
        \round_in[0][988] , \round_in[0][987] , \round_in[0][986] , 
        \round_in[0][985] , \round_in[0][984] , \round_in[0][983] , 
        \round_in[0][982] , \round_in[0][981] , \round_in[0][980] , 
        \round_in[0][979] , \round_in[0][978] , \round_in[0][977] , 
        \round_in[0][976] , \round_in[0][975] , \round_in[0][974] , 
        \round_in[0][973] , \round_in[0][972] , \round_in[0][971] , 
        \round_in[0][970] , \round_in[0][969] , \round_in[0][968] , 
        \round_in[0][967] , \round_in[0][966] , \round_in[0][965] , 
        \round_in[0][964] , \round_in[0][963] , \round_in[0][962] , 
        \round_in[0][961] , \round_in[0][960] , \round_in[0][959] , 
        \round_in[0][958] , \round_in[0][957] , \round_in[0][956] , 
        \round_in[0][955] , \round_in[0][954] , \round_in[0][953] , 
        \round_in[0][952] , \round_in[0][951] , \round_in[0][950] , 
        \round_in[0][949] , \round_in[0][948] , \round_in[0][947] , 
        \round_in[0][946] , \round_in[0][945] , \round_in[0][944] , 
        \round_in[0][943] , \round_in[0][942] , \round_in[0][941] , 
        \round_in[0][940] , \round_in[0][939] , \round_in[0][938] , 
        \round_in[0][937] , \round_in[0][936] , \round_in[0][935] , 
        \round_in[0][934] , \round_in[0][933] , \round_in[0][932] , 
        \round_in[0][931] , \round_in[0][930] , \round_in[0][929] , 
        \round_in[0][928] , \round_in[0][927] , \round_in[0][926] , 
        \round_in[0][925] , \round_in[0][924] , \round_in[0][923] , 
        \round_in[0][922] , \round_in[0][921] , \round_in[0][920] , 
        \round_in[0][919] , \round_in[0][918] , \round_in[0][917] , 
        \round_in[0][916] , \round_in[0][915] , \round_in[0][914] , 
        \round_in[0][913] , \round_in[0][912] , \round_in[0][911] , 
        \round_in[0][910] , \round_in[0][909] , \round_in[0][908] , 
        \round_in[0][907] , \round_in[0][906] , \round_in[0][905] , 
        \round_in[0][904] , \round_in[0][903] , \round_in[0][902] , 
        \round_in[0][901] , \round_in[0][900] , \round_in[0][899] , 
        \round_in[0][898] , \round_in[0][897] , \round_in[0][896] , 
        \round_in[0][895] , \round_in[0][894] , \round_in[0][893] , 
        \round_in[0][892] , \round_in[0][891] , \round_in[0][890] , 
        \round_in[0][889] , \round_in[0][888] , \round_in[0][887] , 
        \round_in[0][886] , \round_in[0][885] , \round_in[0][884] , 
        \round_in[0][883] , \round_in[0][882] , \round_in[0][881] , 
        \round_in[0][880] , \round_in[0][879] , \round_in[0][878] , 
        \round_in[0][877] , \round_in[0][876] , \round_in[0][875] , 
        \round_in[0][874] , \round_in[0][873] , \round_in[0][872] , 
        \round_in[0][871] , \round_in[0][870] , \round_in[0][869] , 
        \round_in[0][868] , \round_in[0][867] , \round_in[0][866] , 
        \round_in[0][865] , \round_in[0][864] , \round_in[0][863] , 
        \round_in[0][862] , \round_in[0][861] , \round_in[0][860] , 
        \round_in[0][859] , \round_in[0][858] , \round_in[0][857] , 
        \round_in[0][856] , \round_in[0][855] , \round_in[0][854] , 
        \round_in[0][853] , \round_in[0][852] , \round_in[0][851] , 
        \round_in[0][850] , \round_in[0][849] , \round_in[0][848] , 
        \round_in[0][847] , \round_in[0][846] , \round_in[0][845] , 
        \round_in[0][844] , \round_in[0][843] , \round_in[0][842] , 
        \round_in[0][841] , \round_in[0][840] , \round_in[0][839] , 
        \round_in[0][838] , \round_in[0][837] , \round_in[0][836] , 
        \round_in[0][835] , \round_in[0][834] , \round_in[0][833] , 
        \round_in[0][832] , \round_in[0][831] , \round_in[0][830] , 
        \round_in[0][829] , \round_in[0][828] , \round_in[0][827] , 
        \round_in[0][826] , \round_in[0][825] , \round_in[0][824] , 
        \round_in[0][823] , \round_in[0][822] , \round_in[0][821] , 
        \round_in[0][820] , \round_in[0][819] , \round_in[0][818] , 
        \round_in[0][817] , \round_in[0][816] , \round_in[0][815] , 
        \round_in[0][814] , \round_in[0][813] , \round_in[0][812] , 
        \round_in[0][811] , \round_in[0][810] , \round_in[0][809] , 
        \round_in[0][808] , \round_in[0][807] , \round_in[0][806] , 
        \round_in[0][805] , \round_in[0][804] , \round_in[0][803] , 
        \round_in[0][802] , \round_in[0][801] , \round_in[0][800] , 
        \round_in[0][799] , \round_in[0][798] , \round_in[0][797] , 
        \round_in[0][796] , \round_in[0][795] , \round_in[0][794] , 
        \round_in[0][793] , \round_in[0][792] , \round_in[0][791] , 
        \round_in[0][790] , \round_in[0][789] , \round_in[0][788] , 
        \round_in[0][787] , \round_in[0][786] , \round_in[0][785] , 
        \round_in[0][784] , \round_in[0][783] , \round_in[0][782] , 
        \round_in[0][781] , \round_in[0][780] , \round_in[0][779] , 
        \round_in[0][778] , \round_in[0][777] , \round_in[0][776] , 
        \round_in[0][775] , \round_in[0][774] , \round_in[0][773] , 
        \round_in[0][772] , \round_in[0][771] , \round_in[0][770] , 
        \round_in[0][769] , \round_in[0][768] , \round_in[0][767] , 
        \round_in[0][766] , \round_in[0][765] , \round_in[0][764] , 
        \round_in[0][763] , \round_in[0][762] , \round_in[0][761] , 
        \round_in[0][760] , \round_in[0][759] , \round_in[0][758] , 
        \round_in[0][757] , \round_in[0][756] , \round_in[0][755] , 
        \round_in[0][754] , \round_in[0][753] , \round_in[0][752] , 
        \round_in[0][751] , \round_in[0][750] , \round_in[0][749] , 
        \round_in[0][748] , \round_in[0][747] , \round_in[0][746] , 
        \round_in[0][745] , \round_in[0][744] , \round_in[0][743] , 
        \round_in[0][742] , \round_in[0][741] , \round_in[0][740] , 
        \round_in[0][739] , \round_in[0][738] , \round_in[0][737] , 
        \round_in[0][736] , \round_in[0][735] , \round_in[0][734] , 
        \round_in[0][733] , \round_in[0][732] , \round_in[0][731] , 
        \round_in[0][730] , \round_in[0][729] , \round_in[0][728] , 
        \round_in[0][727] , \round_in[0][726] , \round_in[0][725] , 
        \round_in[0][724] , \round_in[0][723] , \round_in[0][722] , 
        \round_in[0][721] , \round_in[0][720] , \round_in[0][719] , 
        \round_in[0][718] , \round_in[0][717] , \round_in[0][716] , 
        \round_in[0][715] , \round_in[0][714] , \round_in[0][713] , 
        \round_in[0][712] , \round_in[0][711] , \round_in[0][710] , 
        \round_in[0][709] , \round_in[0][708] , \round_in[0][707] , 
        \round_in[0][706] , \round_in[0][705] , \round_in[0][704] , 
        \round_in[0][703] , \round_in[0][702] , \round_in[0][701] , 
        \round_in[0][700] , \round_in[0][699] , \round_in[0][698] , 
        \round_in[0][697] , \round_in[0][696] , \round_in[0][695] , 
        \round_in[0][694] , \round_in[0][693] , \round_in[0][692] , 
        \round_in[0][691] , \round_in[0][690] , \round_in[0][689] , 
        \round_in[0][688] , \round_in[0][687] , \round_in[0][686] , 
        \round_in[0][685] , \round_in[0][684] , \round_in[0][683] , 
        \round_in[0][682] , \round_in[0][681] , \round_in[0][680] , 
        \round_in[0][679] , \round_in[0][678] , \round_in[0][677] , 
        \round_in[0][676] , \round_in[0][675] , \round_in[0][674] , 
        \round_in[0][673] , \round_in[0][672] , \round_in[0][671] , 
        \round_in[0][670] , \round_in[0][669] , \round_in[0][668] , 
        \round_in[0][667] , \round_in[0][666] , \round_in[0][665] , 
        \round_in[0][664] , \round_in[0][663] , \round_in[0][662] , 
        \round_in[0][661] , \round_in[0][660] , \round_in[0][659] , 
        \round_in[0][658] , \round_in[0][657] , \round_in[0][656] , 
        \round_in[0][655] , \round_in[0][654] , \round_in[0][653] , 
        \round_in[0][652] , \round_in[0][651] , \round_in[0][650] , 
        \round_in[0][649] , \round_in[0][648] , \round_in[0][647] , 
        \round_in[0][646] , \round_in[0][645] , \round_in[0][644] , 
        \round_in[0][643] , \round_in[0][642] , \round_in[0][641] , 
        \round_in[0][640] , \round_in[0][639] , \round_in[0][638] , 
        \round_in[0][637] , \round_in[0][636] , \round_in[0][635] , 
        \round_in[0][634] , \round_in[0][633] , \round_in[0][632] , 
        \round_in[0][631] , \round_in[0][630] , \round_in[0][629] , 
        \round_in[0][628] , \round_in[0][627] , \round_in[0][626] , 
        \round_in[0][625] , \round_in[0][624] , \round_in[0][623] , 
        \round_in[0][622] , \round_in[0][621] , \round_in[0][620] , 
        \round_in[0][619] , \round_in[0][618] , \round_in[0][617] , 
        \round_in[0][616] , \round_in[0][615] , \round_in[0][614] , 
        \round_in[0][613] , \round_in[0][612] , \round_in[0][611] , 
        \round_in[0][610] , \round_in[0][609] , \round_in[0][608] , 
        \round_in[0][607] , \round_in[0][606] , \round_in[0][605] , 
        \round_in[0][604] , \round_in[0][603] , \round_in[0][602] , 
        \round_in[0][601] , \round_in[0][600] , \round_in[0][599] , 
        \round_in[0][598] , \round_in[0][597] , \round_in[0][596] , 
        \round_in[0][595] , \round_in[0][594] , \round_in[0][593] , 
        \round_in[0][592] , \round_in[0][591] , \round_in[0][590] , 
        \round_in[0][589] , \round_in[0][588] , \round_in[0][587] , 
        \round_in[0][586] , \round_in[0][585] , \round_in[0][584] , 
        \round_in[0][583] , \round_in[0][582] , \round_in[0][581] , 
        \round_in[0][580] , \round_in[0][579] , \round_in[0][578] , 
        \round_in[0][577] , \round_in[0][576] , \round_in[0][575] , 
        \round_in[0][574] , \round_in[0][573] , \round_in[0][572] , 
        \round_in[0][571] , \round_in[0][570] , \round_in[0][569] , 
        \round_in[0][568] , \round_in[0][567] , \round_in[0][566] , 
        \round_in[0][565] , \round_in[0][564] , \round_in[0][563] , 
        \round_in[0][562] , \round_in[0][561] , \round_in[0][560] , 
        \round_in[0][559] , \round_in[0][558] , \round_in[0][557] , 
        \round_in[0][556] , \round_in[0][555] , \round_in[0][554] , 
        \round_in[0][553] , \round_in[0][552] , \round_in[0][551] , 
        \round_in[0][550] , \round_in[0][549] , \round_in[0][548] , 
        \round_in[0][547] , \round_in[0][546] , \round_in[0][545] , 
        \round_in[0][544] , \round_in[0][543] , \round_in[0][542] , 
        \round_in[0][541] , \round_in[0][540] , \round_in[0][539] , 
        \round_in[0][538] , \round_in[0][537] , \round_in[0][536] , 
        \round_in[0][535] , \round_in[0][534] , \round_in[0][533] , 
        \round_in[0][532] , \round_in[0][531] , \round_in[0][530] , 
        \round_in[0][529] , \round_in[0][528] , \round_in[0][527] , 
        \round_in[0][526] , \round_in[0][525] , \round_in[0][524] , 
        \round_in[0][523] , \round_in[0][522] , \round_in[0][521] , 
        \round_in[0][520] , \round_in[0][519] , \round_in[0][518] , 
        \round_in[0][517] , \round_in[0][516] , \round_in[0][515] , 
        \round_in[0][514] , \round_in[0][513] , \round_in[0][512] , 
        \round_in[0][511] , \round_in[0][510] , \round_in[0][509] , 
        \round_in[0][508] , \round_in[0][507] , \round_in[0][506] , 
        \round_in[0][505] , \round_in[0][504] , \round_in[0][503] , 
        \round_in[0][502] , \round_in[0][501] , \round_in[0][500] , 
        \round_in[0][499] , \round_in[0][498] , \round_in[0][497] , 
        \round_in[0][496] , \round_in[0][495] , \round_in[0][494] , 
        \round_in[0][493] , \round_in[0][492] , \round_in[0][491] , 
        \round_in[0][490] , \round_in[0][489] , \round_in[0][488] , 
        \round_in[0][487] , \round_in[0][486] , \round_in[0][485] , 
        \round_in[0][484] , \round_in[0][483] , \round_in[0][482] , 
        \round_in[0][481] , \round_in[0][480] , \round_in[0][479] , 
        \round_in[0][478] , \round_in[0][477] , \round_in[0][476] , 
        \round_in[0][475] , \round_in[0][474] , \round_in[0][473] , 
        \round_in[0][472] , \round_in[0][471] , \round_in[0][470] , 
        \round_in[0][469] , \round_in[0][468] , \round_in[0][467] , 
        \round_in[0][466] , \round_in[0][465] , \round_in[0][464] , 
        \round_in[0][463] , \round_in[0][462] , \round_in[0][461] , 
        \round_in[0][460] , \round_in[0][459] , \round_in[0][458] , 
        \round_in[0][457] , \round_in[0][456] , \round_in[0][455] , 
        \round_in[0][454] , \round_in[0][453] , \round_in[0][452] , 
        \round_in[0][451] , \round_in[0][450] , \round_in[0][449] , 
        \round_in[0][448] , \round_in[0][447] , \round_in[0][446] , 
        \round_in[0][445] , \round_in[0][444] , \round_in[0][443] , 
        \round_in[0][442] , \round_in[0][441] , \round_in[0][440] , 
        \round_in[0][439] , \round_in[0][438] , \round_in[0][437] , 
        \round_in[0][436] , \round_in[0][435] , \round_in[0][434] , 
        \round_in[0][433] , \round_in[0][432] , \round_in[0][431] , 
        \round_in[0][430] , \round_in[0][429] , \round_in[0][428] , 
        \round_in[0][427] , \round_in[0][426] , \round_in[0][425] , 
        \round_in[0][424] , \round_in[0][423] , \round_in[0][422] , 
        \round_in[0][421] , \round_in[0][420] , \round_in[0][419] , 
        \round_in[0][418] , \round_in[0][417] , \round_in[0][416] , 
        \round_in[0][415] , \round_in[0][414] , \round_in[0][413] , 
        \round_in[0][412] , \round_in[0][411] , \round_in[0][410] , 
        \round_in[0][409] , \round_in[0][408] , \round_in[0][407] , 
        \round_in[0][406] , \round_in[0][405] , \round_in[0][404] , 
        \round_in[0][403] , \round_in[0][402] , \round_in[0][401] , 
        \round_in[0][400] , \round_in[0][399] , \round_in[0][398] , 
        \round_in[0][397] , \round_in[0][396] , \round_in[0][395] , 
        \round_in[0][394] , \round_in[0][393] , \round_in[0][392] , 
        \round_in[0][391] , \round_in[0][390] , \round_in[0][389] , 
        \round_in[0][388] , \round_in[0][387] , \round_in[0][386] , 
        \round_in[0][385] , \round_in[0][384] , \round_in[0][383] , 
        \round_in[0][382] , \round_in[0][381] , \round_in[0][380] , 
        \round_in[0][379] , \round_in[0][378] , \round_in[0][377] , 
        \round_in[0][376] , \round_in[0][375] , \round_in[0][374] , 
        \round_in[0][373] , \round_in[0][372] , \round_in[0][371] , 
        \round_in[0][370] , \round_in[0][369] , \round_in[0][368] , 
        \round_in[0][367] , \round_in[0][366] , \round_in[0][365] , 
        \round_in[0][364] , \round_in[0][363] , \round_in[0][362] , 
        \round_in[0][361] , \round_in[0][360] , \round_in[0][359] , 
        \round_in[0][358] , \round_in[0][357] , \round_in[0][356] , 
        \round_in[0][355] , \round_in[0][354] , \round_in[0][353] , 
        \round_in[0][352] , \round_in[0][351] , \round_in[0][350] , 
        \round_in[0][349] , \round_in[0][348] , \round_in[0][347] , 
        \round_in[0][346] , \round_in[0][345] , \round_in[0][344] , 
        \round_in[0][343] , \round_in[0][342] , \round_in[0][341] , 
        \round_in[0][340] , \round_in[0][339] , \round_in[0][338] , 
        \round_in[0][337] , \round_in[0][336] , \round_in[0][335] , 
        \round_in[0][334] , \round_in[0][333] , \round_in[0][332] , 
        \round_in[0][331] , \round_in[0][330] , \round_in[0][329] , 
        \round_in[0][328] , \round_in[0][327] , \round_in[0][326] , 
        \round_in[0][325] , \round_in[0][324] , \round_in[0][323] , 
        \round_in[0][322] , \round_in[0][321] , \round_in[0][320] , 
        \round_in[0][319] , \round_in[0][318] , \round_in[0][317] , 
        \round_in[0][316] , \round_in[0][315] , \round_in[0][314] , 
        \round_in[0][313] , \round_in[0][312] , \round_in[0][311] , 
        \round_in[0][310] , \round_in[0][309] , \round_in[0][308] , 
        \round_in[0][307] , \round_in[0][306] , \round_in[0][305] , 
        \round_in[0][304] , \round_in[0][303] , \round_in[0][302] , 
        \round_in[0][301] , \round_in[0][300] , \round_in[0][299] , 
        \round_in[0][298] , \round_in[0][297] , \round_in[0][296] , 
        \round_in[0][295] , \round_in[0][294] , \round_in[0][293] , 
        \round_in[0][292] , \round_in[0][291] , \round_in[0][290] , 
        \round_in[0][289] , \round_in[0][288] , \round_in[0][287] , 
        \round_in[0][286] , \round_in[0][285] , \round_in[0][284] , 
        \round_in[0][283] , \round_in[0][282] , \round_in[0][281] , 
        \round_in[0][280] , \round_in[0][279] , \round_in[0][278] , 
        \round_in[0][277] , \round_in[0][276] , \round_in[0][275] , 
        \round_in[0][274] , \round_in[0][273] , \round_in[0][272] , 
        \round_in[0][271] , \round_in[0][270] , \round_in[0][269] , 
        \round_in[0][268] , \round_in[0][267] , \round_in[0][266] , 
        \round_in[0][265] , \round_in[0][264] , \round_in[0][263] , 
        \round_in[0][262] , \round_in[0][261] , \round_in[0][260] , 
        \round_in[0][259] , \round_in[0][258] , \round_in[0][257] , 
        \round_in[0][256] , \round_in[0][255] , \round_in[0][254] , 
        \round_in[0][253] , \round_in[0][252] , \round_in[0][251] , 
        \round_in[0][250] , \round_in[0][249] , \round_in[0][248] , 
        \round_in[0][247] , \round_in[0][246] , \round_in[0][245] , 
        \round_in[0][244] , \round_in[0][243] , \round_in[0][242] , 
        \round_in[0][241] , \round_in[0][240] , \round_in[0][239] , 
        \round_in[0][238] , \round_in[0][237] , \round_in[0][236] , 
        \round_in[0][235] , \round_in[0][234] , \round_in[0][233] , 
        \round_in[0][232] , \round_in[0][231] , \round_in[0][230] , 
        \round_in[0][229] , \round_in[0][228] , \round_in[0][227] , 
        \round_in[0][226] , \round_in[0][225] , \round_in[0][224] , 
        \round_in[0][223] , \round_in[0][222] , \round_in[0][221] , 
        \round_in[0][220] , \round_in[0][219] , \round_in[0][218] , 
        \round_in[0][217] , \round_in[0][216] , \round_in[0][215] , 
        \round_in[0][214] , \round_in[0][213] , \round_in[0][212] , 
        \round_in[0][211] , \round_in[0][210] , \round_in[0][209] , 
        \round_in[0][208] , \round_in[0][207] , \round_in[0][206] , 
        \round_in[0][205] , \round_in[0][204] , \round_in[0][203] , 
        \round_in[0][202] , \round_in[0][201] , \round_in[0][200] , 
        \round_in[0][199] , \round_in[0][198] , \round_in[0][197] , 
        \round_in[0][196] , \round_in[0][195] , \round_in[0][194] , 
        \round_in[0][193] , \round_in[0][192] , \round_in[0][191] , 
        \round_in[0][190] , \round_in[0][189] , \round_in[0][188] , 
        \round_in[0][187] , \round_in[0][186] , \round_in[0][185] , 
        \round_in[0][184] , \round_in[0][183] , \round_in[0][182] , 
        \round_in[0][181] , \round_in[0][180] , \round_in[0][179] , 
        \round_in[0][178] , \round_in[0][177] , \round_in[0][176] , 
        \round_in[0][175] , \round_in[0][174] , \round_in[0][173] , 
        \round_in[0][172] , \round_in[0][171] , \round_in[0][170] , 
        \round_in[0][169] , \round_in[0][168] , \round_in[0][167] , 
        \round_in[0][166] , \round_in[0][165] , \round_in[0][164] , 
        \round_in[0][163] , \round_in[0][162] , \round_in[0][161] , 
        \round_in[0][160] , \round_in[0][159] , \round_in[0][158] , 
        \round_in[0][157] , \round_in[0][156] , \round_in[0][155] , 
        \round_in[0][154] , \round_in[0][153] , \round_in[0][152] , 
        \round_in[0][151] , \round_in[0][150] , \round_in[0][149] , 
        \round_in[0][148] , \round_in[0][147] , \round_in[0][146] , 
        \round_in[0][145] , \round_in[0][144] , \round_in[0][143] , 
        \round_in[0][142] , \round_in[0][141] , \round_in[0][140] , 
        \round_in[0][139] , \round_in[0][138] , \round_in[0][137] , 
        \round_in[0][136] , \round_in[0][135] , \round_in[0][134] , 
        \round_in[0][133] , \round_in[0][132] , \round_in[0][131] , 
        \round_in[0][130] , \round_in[0][129] , \round_in[0][128] , 
        \round_in[0][127] , \round_in[0][126] , \round_in[0][125] , 
        \round_in[0][124] , \round_in[0][123] , \round_in[0][122] , 
        \round_in[0][121] , \round_in[0][120] , \round_in[0][119] , 
        \round_in[0][118] , \round_in[0][117] , \round_in[0][116] , 
        \round_in[0][115] , \round_in[0][114] , \round_in[0][113] , 
        \round_in[0][112] , \round_in[0][111] , \round_in[0][110] , 
        \round_in[0][109] , \round_in[0][108] , \round_in[0][107] , 
        \round_in[0][106] , \round_in[0][105] , \round_in[0][104] , 
        \round_in[0][103] , \round_in[0][102] , \round_in[0][101] , 
        \round_in[0][100] , \round_in[0][99] , \round_in[0][98] , 
        \round_in[0][97] , \round_in[0][96] , \round_in[0][95] , 
        \round_in[0][94] , \round_in[0][93] , \round_in[0][92] , 
        \round_in[0][91] , \round_in[0][90] , \round_in[0][89] , 
        \round_in[0][88] , \round_in[0][87] , \round_in[0][86] , 
        \round_in[0][85] , \round_in[0][84] , \round_in[0][83] , 
        \round_in[0][82] , \round_in[0][81] , \round_in[0][80] , 
        \round_in[0][79] , \round_in[0][78] , \round_in[0][77] , 
        \round_in[0][76] , \round_in[0][75] , \round_in[0][74] , 
        \round_in[0][73] , \round_in[0][72] , \round_in[0][71] , 
        \round_in[0][70] , \round_in[0][69] , \round_in[0][68] , 
        \round_in[0][67] , \round_in[0][66] , \round_in[0][65] , 
        \round_in[0][64] , \round_in[0][63] , \round_in[0][62] , 
        \round_in[0][61] , \round_in[0][60] , \round_in[0][59] , 
        \round_in[0][58] , \round_in[0][57] , \round_in[0][56] , 
        \round_in[0][55] , \round_in[0][54] , \round_in[0][53] , 
        \round_in[0][52] , \round_in[0][51] , \round_in[0][50] , 
        \round_in[0][49] , \round_in[0][48] , \round_in[0][47] , 
        \round_in[0][46] , \round_in[0][45] , \round_in[0][44] , 
        \round_in[0][43] , \round_in[0][42] , \round_in[0][41] , 
        \round_in[0][40] , \round_in[0][39] , \round_in[0][38] , 
        \round_in[0][37] , \round_in[0][36] , \round_in[0][35] , 
        \round_in[0][34] , \round_in[0][33] , \round_in[0][32] , 
        \round_in[0][31] , \round_in[0][30] , \round_in[0][29] , 
        \round_in[0][28] , \round_in[0][27] , \round_in[0][26] , 
        \round_in[0][25] , \round_in[0][24] , \round_in[0][23] , 
        \round_in[0][22] , \round_in[0][21] , \round_in[0][20] , 
        \round_in[0][19] , \round_in[0][18] , \round_in[0][17] , 
        \round_in[0][16] , \round_in[0][15] , \round_in[0][14] , 
        \round_in[0][13] , \round_in[0][12] , \round_in[0][11] , 
        \round_in[0][10] , \round_in[0][9] , \round_in[0][8] , 
        \round_in[0][7] , \round_in[0][6] , \round_in[0][5] , \round_in[0][4] , 
        \round_in[0][3] , \round_in[0][2] , \round_in[0][1] , \round_in[0][0] }), .round_const({\RCONST[0].rconst_/N67 , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, \RCONST[0].rconst_/N57 , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \RCONST[0].rconst_/N48 , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \RCONST[0].rconst_/N37 , 1'b0, 1'b0, 1'b0, \RCONST[0].rconst_/N28 , 
        1'b0, \RCONST[0].rconst_/N18 , \rc[0][0] }), .out({\round_in[1][1599] , 
        \round_in[1][1598] , \round_in[1][1597] , \round_in[1][1596] , 
        \round_in[1][1595] , \round_in[1][1594] , \round_in[1][1593] , 
        \round_in[1][1592] , \round_in[1][1591] , \round_in[1][1590] , 
        \round_in[1][1589] , \round_in[1][1588] , \round_in[1][1587] , 
        \round_in[1][1586] , \round_in[1][1585] , \round_in[1][1584] , 
        \round_in[1][1583] , \round_in[1][1582] , \round_in[1][1581] , 
        \round_in[1][1580] , \round_in[1][1579] , \round_in[1][1578] , 
        \round_in[1][1577] , \round_in[1][1576] , \round_in[1][1575] , 
        \round_in[1][1574] , \round_in[1][1573] , \round_in[1][1572] , 
        \round_in[1][1571] , \round_in[1][1570] , \round_in[1][1569] , 
        \round_in[1][1568] , \round_in[1][1567] , \round_in[1][1566] , 
        \round_in[1][1565] , \round_in[1][1564] , \round_in[1][1563] , 
        \round_in[1][1562] , \round_in[1][1561] , \round_in[1][1560] , 
        \round_in[1][1559] , \round_in[1][1558] , \round_in[1][1557] , 
        \round_in[1][1556] , \round_in[1][1555] , \round_in[1][1554] , 
        \round_in[1][1553] , \round_in[1][1552] , \round_in[1][1551] , 
        \round_in[1][1550] , \round_in[1][1549] , \round_in[1][1548] , 
        \round_in[1][1547] , \round_in[1][1546] , \round_in[1][1545] , 
        \round_in[1][1544] , \round_in[1][1543] , \round_in[1][1542] , 
        \round_in[1][1541] , \round_in[1][1540] , \round_in[1][1539] , 
        \round_in[1][1538] , \round_in[1][1537] , \round_in[1][1536] , 
        \round_in[1][1535] , \round_in[1][1534] , \round_in[1][1533] , 
        \round_in[1][1532] , \round_in[1][1531] , \round_in[1][1530] , 
        \round_in[1][1529] , \round_in[1][1528] , \round_in[1][1527] , 
        \round_in[1][1526] , \round_in[1][1525] , \round_in[1][1524] , 
        \round_in[1][1523] , \round_in[1][1522] , \round_in[1][1521] , 
        \round_in[1][1520] , \round_in[1][1519] , \round_in[1][1518] , 
        \round_in[1][1517] , \round_in[1][1516] , \round_in[1][1515] , 
        \round_in[1][1514] , \round_in[1][1513] , \round_in[1][1512] , 
        \round_in[1][1511] , \round_in[1][1510] , \round_in[1][1509] , 
        \round_in[1][1508] , \round_in[1][1507] , \round_in[1][1506] , 
        \round_in[1][1505] , \round_in[1][1504] , \round_in[1][1503] , 
        \round_in[1][1502] , \round_in[1][1501] , \round_in[1][1500] , 
        \round_in[1][1499] , \round_in[1][1498] , \round_in[1][1497] , 
        \round_in[1][1496] , \round_in[1][1495] , \round_in[1][1494] , 
        \round_in[1][1493] , \round_in[1][1492] , \round_in[1][1491] , 
        \round_in[1][1490] , \round_in[1][1489] , \round_in[1][1488] , 
        \round_in[1][1487] , \round_in[1][1486] , \round_in[1][1485] , 
        \round_in[1][1484] , \round_in[1][1483] , \round_in[1][1482] , 
        \round_in[1][1481] , \round_in[1][1480] , \round_in[1][1479] , 
        \round_in[1][1478] , \round_in[1][1477] , \round_in[1][1476] , 
        \round_in[1][1475] , \round_in[1][1474] , \round_in[1][1473] , 
        \round_in[1][1472] , \round_in[1][1471] , \round_in[1][1470] , 
        \round_in[1][1469] , \round_in[1][1468] , \round_in[1][1467] , 
        \round_in[1][1466] , \round_in[1][1465] , \round_in[1][1464] , 
        \round_in[1][1463] , \round_in[1][1462] , \round_in[1][1461] , 
        \round_in[1][1460] , \round_in[1][1459] , \round_in[1][1458] , 
        \round_in[1][1457] , \round_in[1][1456] , \round_in[1][1455] , 
        \round_in[1][1454] , \round_in[1][1453] , \round_in[1][1452] , 
        \round_in[1][1451] , \round_in[1][1450] , \round_in[1][1449] , 
        \round_in[1][1448] , \round_in[1][1447] , \round_in[1][1446] , 
        \round_in[1][1445] , \round_in[1][1444] , \round_in[1][1443] , 
        \round_in[1][1442] , \round_in[1][1441] , \round_in[1][1440] , 
        \round_in[1][1439] , \round_in[1][1438] , \round_in[1][1437] , 
        \round_in[1][1436] , \round_in[1][1435] , \round_in[1][1434] , 
        \round_in[1][1433] , \round_in[1][1432] , \round_in[1][1431] , 
        \round_in[1][1430] , \round_in[1][1429] , \round_in[1][1428] , 
        \round_in[1][1427] , \round_in[1][1426] , \round_in[1][1425] , 
        \round_in[1][1424] , \round_in[1][1423] , \round_in[1][1422] , 
        \round_in[1][1421] , \round_in[1][1420] , \round_in[1][1419] , 
        \round_in[1][1418] , \round_in[1][1417] , \round_in[1][1416] , 
        \round_in[1][1415] , \round_in[1][1414] , \round_in[1][1413] , 
        \round_in[1][1412] , \round_in[1][1411] , \round_in[1][1410] , 
        \round_in[1][1409] , \round_in[1][1408] , \round_in[1][1407] , 
        \round_in[1][1406] , \round_in[1][1405] , \round_in[1][1404] , 
        \round_in[1][1403] , \round_in[1][1402] , \round_in[1][1401] , 
        \round_in[1][1400] , \round_in[1][1399] , \round_in[1][1398] , 
        \round_in[1][1397] , \round_in[1][1396] , \round_in[1][1395] , 
        \round_in[1][1394] , \round_in[1][1393] , \round_in[1][1392] , 
        \round_in[1][1391] , \round_in[1][1390] , \round_in[1][1389] , 
        \round_in[1][1388] , \round_in[1][1387] , \round_in[1][1386] , 
        \round_in[1][1385] , \round_in[1][1384] , \round_in[1][1383] , 
        \round_in[1][1382] , \round_in[1][1381] , \round_in[1][1380] , 
        \round_in[1][1379] , \round_in[1][1378] , \round_in[1][1377] , 
        \round_in[1][1376] , \round_in[1][1375] , \round_in[1][1374] , 
        \round_in[1][1373] , \round_in[1][1372] , \round_in[1][1371] , 
        \round_in[1][1370] , \round_in[1][1369] , \round_in[1][1368] , 
        \round_in[1][1367] , \round_in[1][1366] , \round_in[1][1365] , 
        \round_in[1][1364] , \round_in[1][1363] , \round_in[1][1362] , 
        \round_in[1][1361] , \round_in[1][1360] , \round_in[1][1359] , 
        \round_in[1][1358] , \round_in[1][1357] , \round_in[1][1356] , 
        \round_in[1][1355] , \round_in[1][1354] , \round_in[1][1353] , 
        \round_in[1][1352] , \round_in[1][1351] , \round_in[1][1350] , 
        \round_in[1][1349] , \round_in[1][1348] , \round_in[1][1347] , 
        \round_in[1][1346] , \round_in[1][1345] , \round_in[1][1344] , 
        \round_in[1][1343] , \round_in[1][1342] , \round_in[1][1341] , 
        \round_in[1][1340] , \round_in[1][1339] , \round_in[1][1338] , 
        \round_in[1][1337] , \round_in[1][1336] , \round_in[1][1335] , 
        \round_in[1][1334] , \round_in[1][1333] , \round_in[1][1332] , 
        \round_in[1][1331] , \round_in[1][1330] , \round_in[1][1329] , 
        \round_in[1][1328] , \round_in[1][1327] , \round_in[1][1326] , 
        \round_in[1][1325] , \round_in[1][1324] , \round_in[1][1323] , 
        \round_in[1][1322] , \round_in[1][1321] , \round_in[1][1320] , 
        \round_in[1][1319] , \round_in[1][1318] , \round_in[1][1317] , 
        \round_in[1][1316] , \round_in[1][1315] , \round_in[1][1314] , 
        \round_in[1][1313] , \round_in[1][1312] , \round_in[1][1311] , 
        \round_in[1][1310] , \round_in[1][1309] , \round_in[1][1308] , 
        \round_in[1][1307] , \round_in[1][1306] , \round_in[1][1305] , 
        \round_in[1][1304] , \round_in[1][1303] , \round_in[1][1302] , 
        \round_in[1][1301] , \round_in[1][1300] , \round_in[1][1299] , 
        \round_in[1][1298] , \round_in[1][1297] , \round_in[1][1296] , 
        \round_in[1][1295] , \round_in[1][1294] , \round_in[1][1293] , 
        \round_in[1][1292] , \round_in[1][1291] , \round_in[1][1290] , 
        \round_in[1][1289] , \round_in[1][1288] , \round_in[1][1287] , 
        \round_in[1][1286] , \round_in[1][1285] , \round_in[1][1284] , 
        \round_in[1][1283] , \round_in[1][1282] , \round_in[1][1281] , 
        \round_in[1][1280] , \round_in[1][1279] , \round_in[1][1278] , 
        \round_in[1][1277] , \round_in[1][1276] , \round_in[1][1275] , 
        \round_in[1][1274] , \round_in[1][1273] , \round_in[1][1272] , 
        \round_in[1][1271] , \round_in[1][1270] , \round_in[1][1269] , 
        \round_in[1][1268] , \round_in[1][1267] , \round_in[1][1266] , 
        \round_in[1][1265] , \round_in[1][1264] , \round_in[1][1263] , 
        \round_in[1][1262] , \round_in[1][1261] , \round_in[1][1260] , 
        \round_in[1][1259] , \round_in[1][1258] , \round_in[1][1257] , 
        \round_in[1][1256] , \round_in[1][1255] , \round_in[1][1254] , 
        \round_in[1][1253] , \round_in[1][1252] , \round_in[1][1251] , 
        \round_in[1][1250] , \round_in[1][1249] , \round_in[1][1248] , 
        \round_in[1][1247] , \round_in[1][1246] , \round_in[1][1245] , 
        \round_in[1][1244] , \round_in[1][1243] , \round_in[1][1242] , 
        \round_in[1][1241] , \round_in[1][1240] , \round_in[1][1239] , 
        \round_in[1][1238] , \round_in[1][1237] , \round_in[1][1236] , 
        \round_in[1][1235] , \round_in[1][1234] , \round_in[1][1233] , 
        \round_in[1][1232] , \round_in[1][1231] , \round_in[1][1230] , 
        \round_in[1][1229] , \round_in[1][1228] , \round_in[1][1227] , 
        \round_in[1][1226] , \round_in[1][1225] , \round_in[1][1224] , 
        \round_in[1][1223] , \round_in[1][1222] , \round_in[1][1221] , 
        \round_in[1][1220] , \round_in[1][1219] , \round_in[1][1218] , 
        \round_in[1][1217] , \round_in[1][1216] , \round_in[1][1215] , 
        \round_in[1][1214] , \round_in[1][1213] , \round_in[1][1212] , 
        \round_in[1][1211] , \round_in[1][1210] , \round_in[1][1209] , 
        \round_in[1][1208] , \round_in[1][1207] , \round_in[1][1206] , 
        \round_in[1][1205] , \round_in[1][1204] , \round_in[1][1203] , 
        \round_in[1][1202] , \round_in[1][1201] , \round_in[1][1200] , 
        \round_in[1][1199] , \round_in[1][1198] , \round_in[1][1197] , 
        \round_in[1][1196] , \round_in[1][1195] , \round_in[1][1194] , 
        \round_in[1][1193] , \round_in[1][1192] , \round_in[1][1191] , 
        \round_in[1][1190] , \round_in[1][1189] , \round_in[1][1188] , 
        \round_in[1][1187] , \round_in[1][1186] , \round_in[1][1185] , 
        \round_in[1][1184] , \round_in[1][1183] , \round_in[1][1182] , 
        \round_in[1][1181] , \round_in[1][1180] , \round_in[1][1179] , 
        \round_in[1][1178] , \round_in[1][1177] , \round_in[1][1176] , 
        \round_in[1][1175] , \round_in[1][1174] , \round_in[1][1173] , 
        \round_in[1][1172] , \round_in[1][1171] , \round_in[1][1170] , 
        \round_in[1][1169] , \round_in[1][1168] , \round_in[1][1167] , 
        \round_in[1][1166] , \round_in[1][1165] , \round_in[1][1164] , 
        \round_in[1][1163] , \round_in[1][1162] , \round_in[1][1161] , 
        \round_in[1][1160] , \round_in[1][1159] , \round_in[1][1158] , 
        \round_in[1][1157] , \round_in[1][1156] , \round_in[1][1155] , 
        \round_in[1][1154] , \round_in[1][1153] , \round_in[1][1152] , 
        \round_in[1][1151] , \round_in[1][1150] , \round_in[1][1149] , 
        \round_in[1][1148] , \round_in[1][1147] , \round_in[1][1146] , 
        \round_in[1][1145] , \round_in[1][1144] , \round_in[1][1143] , 
        \round_in[1][1142] , \round_in[1][1141] , \round_in[1][1140] , 
        \round_in[1][1139] , \round_in[1][1138] , \round_in[1][1137] , 
        \round_in[1][1136] , \round_in[1][1135] , \round_in[1][1134] , 
        \round_in[1][1133] , \round_in[1][1132] , \round_in[1][1131] , 
        \round_in[1][1130] , \round_in[1][1129] , \round_in[1][1128] , 
        \round_in[1][1127] , \round_in[1][1126] , \round_in[1][1125] , 
        \round_in[1][1124] , \round_in[1][1123] , \round_in[1][1122] , 
        \round_in[1][1121] , \round_in[1][1120] , \round_in[1][1119] , 
        \round_in[1][1118] , \round_in[1][1117] , \round_in[1][1116] , 
        \round_in[1][1115] , \round_in[1][1114] , \round_in[1][1113] , 
        \round_in[1][1112] , \round_in[1][1111] , \round_in[1][1110] , 
        \round_in[1][1109] , \round_in[1][1108] , \round_in[1][1107] , 
        \round_in[1][1106] , \round_in[1][1105] , \round_in[1][1104] , 
        \round_in[1][1103] , \round_in[1][1102] , \round_in[1][1101] , 
        \round_in[1][1100] , \round_in[1][1099] , \round_in[1][1098] , 
        \round_in[1][1097] , \round_in[1][1096] , \round_in[1][1095] , 
        \round_in[1][1094] , \round_in[1][1093] , \round_in[1][1092] , 
        \round_in[1][1091] , \round_in[1][1090] , \round_in[1][1089] , 
        \round_in[1][1088] , \round_in[1][1087] , \round_in[1][1086] , 
        \round_in[1][1085] , \round_in[1][1084] , \round_in[1][1083] , 
        \round_in[1][1082] , \round_in[1][1081] , \round_in[1][1080] , 
        \round_in[1][1079] , \round_in[1][1078] , \round_in[1][1077] , 
        \round_in[1][1076] , \round_in[1][1075] , \round_in[1][1074] , 
        \round_in[1][1073] , \round_in[1][1072] , \round_in[1][1071] , 
        \round_in[1][1070] , \round_in[1][1069] , \round_in[1][1068] , 
        \round_in[1][1067] , \round_in[1][1066] , \round_in[1][1065] , 
        \round_in[1][1064] , \round_in[1][1063] , \round_in[1][1062] , 
        \round_in[1][1061] , \round_in[1][1060] , \round_in[1][1059] , 
        \round_in[1][1058] , \round_in[1][1057] , \round_in[1][1056] , 
        \round_in[1][1055] , \round_in[1][1054] , \round_in[1][1053] , 
        \round_in[1][1052] , \round_in[1][1051] , \round_in[1][1050] , 
        \round_in[1][1049] , \round_in[1][1048] , \round_in[1][1047] , 
        \round_in[1][1046] , \round_in[1][1045] , \round_in[1][1044] , 
        \round_in[1][1043] , \round_in[1][1042] , \round_in[1][1041] , 
        \round_in[1][1040] , \round_in[1][1039] , \round_in[1][1038] , 
        \round_in[1][1037] , \round_in[1][1036] , \round_in[1][1035] , 
        \round_in[1][1034] , \round_in[1][1033] , \round_in[1][1032] , 
        \round_in[1][1031] , \round_in[1][1030] , \round_in[1][1029] , 
        \round_in[1][1028] , \round_in[1][1027] , \round_in[1][1026] , 
        \round_in[1][1025] , \round_in[1][1024] , \round_in[1][1023] , 
        \round_in[1][1022] , \round_in[1][1021] , \round_in[1][1020] , 
        \round_in[1][1019] , \round_in[1][1018] , \round_in[1][1017] , 
        \round_in[1][1016] , \round_in[1][1015] , \round_in[1][1014] , 
        \round_in[1][1013] , \round_in[1][1012] , \round_in[1][1011] , 
        \round_in[1][1010] , \round_in[1][1009] , \round_in[1][1008] , 
        \round_in[1][1007] , \round_in[1][1006] , \round_in[1][1005] , 
        \round_in[1][1004] , \round_in[1][1003] , \round_in[1][1002] , 
        \round_in[1][1001] , \round_in[1][1000] , \round_in[1][999] , 
        \round_in[1][998] , \round_in[1][997] , \round_in[1][996] , 
        \round_in[1][995] , \round_in[1][994] , \round_in[1][993] , 
        \round_in[1][992] , \round_in[1][991] , \round_in[1][990] , 
        \round_in[1][989] , \round_in[1][988] , \round_in[1][987] , 
        \round_in[1][986] , \round_in[1][985] , \round_in[1][984] , 
        \round_in[1][983] , \round_in[1][982] , \round_in[1][981] , 
        \round_in[1][980] , \round_in[1][979] , \round_in[1][978] , 
        \round_in[1][977] , \round_in[1][976] , \round_in[1][975] , 
        \round_in[1][974] , \round_in[1][973] , \round_in[1][972] , 
        \round_in[1][971] , \round_in[1][970] , \round_in[1][969] , 
        \round_in[1][968] , \round_in[1][967] , \round_in[1][966] , 
        \round_in[1][965] , \round_in[1][964] , \round_in[1][963] , 
        \round_in[1][962] , \round_in[1][961] , \round_in[1][960] , 
        \round_in[1][959] , \round_in[1][958] , \round_in[1][957] , 
        \round_in[1][956] , \round_in[1][955] , \round_in[1][954] , 
        \round_in[1][953] , \round_in[1][952] , \round_in[1][951] , 
        \round_in[1][950] , \round_in[1][949] , \round_in[1][948] , 
        \round_in[1][947] , \round_in[1][946] , \round_in[1][945] , 
        \round_in[1][944] , \round_in[1][943] , \round_in[1][942] , 
        \round_in[1][941] , \round_in[1][940] , \round_in[1][939] , 
        \round_in[1][938] , \round_in[1][937] , \round_in[1][936] , 
        \round_in[1][935] , \round_in[1][934] , \round_in[1][933] , 
        \round_in[1][932] , \round_in[1][931] , \round_in[1][930] , 
        \round_in[1][929] , \round_in[1][928] , \round_in[1][927] , 
        \round_in[1][926] , \round_in[1][925] , \round_in[1][924] , 
        \round_in[1][923] , \round_in[1][922] , \round_in[1][921] , 
        \round_in[1][920] , \round_in[1][919] , \round_in[1][918] , 
        \round_in[1][917] , \round_in[1][916] , \round_in[1][915] , 
        \round_in[1][914] , \round_in[1][913] , \round_in[1][912] , 
        \round_in[1][911] , \round_in[1][910] , \round_in[1][909] , 
        \round_in[1][908] , \round_in[1][907] , \round_in[1][906] , 
        \round_in[1][905] , \round_in[1][904] , \round_in[1][903] , 
        \round_in[1][902] , \round_in[1][901] , \round_in[1][900] , 
        \round_in[1][899] , \round_in[1][898] , \round_in[1][897] , 
        \round_in[1][896] , \round_in[1][895] , \round_in[1][894] , 
        \round_in[1][893] , \round_in[1][892] , \round_in[1][891] , 
        \round_in[1][890] , \round_in[1][889] , \round_in[1][888] , 
        \round_in[1][887] , \round_in[1][886] , \round_in[1][885] , 
        \round_in[1][884] , \round_in[1][883] , \round_in[1][882] , 
        \round_in[1][881] , \round_in[1][880] , \round_in[1][879] , 
        \round_in[1][878] , \round_in[1][877] , \round_in[1][876] , 
        \round_in[1][875] , \round_in[1][874] , \round_in[1][873] , 
        \round_in[1][872] , \round_in[1][871] , \round_in[1][870] , 
        \round_in[1][869] , \round_in[1][868] , \round_in[1][867] , 
        \round_in[1][866] , \round_in[1][865] , \round_in[1][864] , 
        \round_in[1][863] , \round_in[1][862] , \round_in[1][861] , 
        \round_in[1][860] , \round_in[1][859] , \round_in[1][858] , 
        \round_in[1][857] , \round_in[1][856] , \round_in[1][855] , 
        \round_in[1][854] , \round_in[1][853] , \round_in[1][852] , 
        \round_in[1][851] , \round_in[1][850] , \round_in[1][849] , 
        \round_in[1][848] , \round_in[1][847] , \round_in[1][846] , 
        \round_in[1][845] , \round_in[1][844] , \round_in[1][843] , 
        \round_in[1][842] , \round_in[1][841] , \round_in[1][840] , 
        \round_in[1][839] , \round_in[1][838] , \round_in[1][837] , 
        \round_in[1][836] , \round_in[1][835] , \round_in[1][834] , 
        \round_in[1][833] , \round_in[1][832] , \round_in[1][831] , 
        \round_in[1][830] , \round_in[1][829] , \round_in[1][828] , 
        \round_in[1][827] , \round_in[1][826] , \round_in[1][825] , 
        \round_in[1][824] , \round_in[1][823] , \round_in[1][822] , 
        \round_in[1][821] , \round_in[1][820] , \round_in[1][819] , 
        \round_in[1][818] , \round_in[1][817] , \round_in[1][816] , 
        \round_in[1][815] , \round_in[1][814] , \round_in[1][813] , 
        \round_in[1][812] , \round_in[1][811] , \round_in[1][810] , 
        \round_in[1][809] , \round_in[1][808] , \round_in[1][807] , 
        \round_in[1][806] , \round_in[1][805] , \round_in[1][804] , 
        \round_in[1][803] , \round_in[1][802] , \round_in[1][801] , 
        \round_in[1][800] , \round_in[1][799] , \round_in[1][798] , 
        \round_in[1][797] , \round_in[1][796] , \round_in[1][795] , 
        \round_in[1][794] , \round_in[1][793] , \round_in[1][792] , 
        \round_in[1][791] , \round_in[1][790] , \round_in[1][789] , 
        \round_in[1][788] , \round_in[1][787] , \round_in[1][786] , 
        \round_in[1][785] , \round_in[1][784] , \round_in[1][783] , 
        \round_in[1][782] , \round_in[1][781] , \round_in[1][780] , 
        \round_in[1][779] , \round_in[1][778] , \round_in[1][777] , 
        \round_in[1][776] , \round_in[1][775] , \round_in[1][774] , 
        \round_in[1][773] , \round_in[1][772] , \round_in[1][771] , 
        \round_in[1][770] , \round_in[1][769] , \round_in[1][768] , 
        \round_in[1][767] , \round_in[1][766] , \round_in[1][765] , 
        \round_in[1][764] , \round_in[1][763] , \round_in[1][762] , 
        \round_in[1][761] , \round_in[1][760] , \round_in[1][759] , 
        \round_in[1][758] , \round_in[1][757] , \round_in[1][756] , 
        \round_in[1][755] , \round_in[1][754] , \round_in[1][753] , 
        \round_in[1][752] , \round_in[1][751] , \round_in[1][750] , 
        \round_in[1][749] , \round_in[1][748] , \round_in[1][747] , 
        \round_in[1][746] , \round_in[1][745] , \round_in[1][744] , 
        \round_in[1][743] , \round_in[1][742] , \round_in[1][741] , 
        \round_in[1][740] , \round_in[1][739] , \round_in[1][738] , 
        \round_in[1][737] , \round_in[1][736] , \round_in[1][735] , 
        \round_in[1][734] , \round_in[1][733] , \round_in[1][732] , 
        \round_in[1][731] , \round_in[1][730] , \round_in[1][729] , 
        \round_in[1][728] , \round_in[1][727] , \round_in[1][726] , 
        \round_in[1][725] , \round_in[1][724] , \round_in[1][723] , 
        \round_in[1][722] , \round_in[1][721] , \round_in[1][720] , 
        \round_in[1][719] , \round_in[1][718] , \round_in[1][717] , 
        \round_in[1][716] , \round_in[1][715] , \round_in[1][714] , 
        \round_in[1][713] , \round_in[1][712] , \round_in[1][711] , 
        \round_in[1][710] , \round_in[1][709] , \round_in[1][708] , 
        \round_in[1][707] , \round_in[1][706] , \round_in[1][705] , 
        \round_in[1][704] , \round_in[1][703] , \round_in[1][702] , 
        \round_in[1][701] , \round_in[1][700] , \round_in[1][699] , 
        \round_in[1][698] , \round_in[1][697] , \round_in[1][696] , 
        \round_in[1][695] , \round_in[1][694] , \round_in[1][693] , 
        \round_in[1][692] , \round_in[1][691] , \round_in[1][690] , 
        \round_in[1][689] , \round_in[1][688] , \round_in[1][687] , 
        \round_in[1][686] , \round_in[1][685] , \round_in[1][684] , 
        \round_in[1][683] , \round_in[1][682] , \round_in[1][681] , 
        \round_in[1][680] , \round_in[1][679] , \round_in[1][678] , 
        \round_in[1][677] , \round_in[1][676] , \round_in[1][675] , 
        \round_in[1][674] , \round_in[1][673] , \round_in[1][672] , 
        \round_in[1][671] , \round_in[1][670] , \round_in[1][669] , 
        \round_in[1][668] , \round_in[1][667] , \round_in[1][666] , 
        \round_in[1][665] , \round_in[1][664] , \round_in[1][663] , 
        \round_in[1][662] , \round_in[1][661] , \round_in[1][660] , 
        \round_in[1][659] , \round_in[1][658] , \round_in[1][657] , 
        \round_in[1][656] , \round_in[1][655] , \round_in[1][654] , 
        \round_in[1][653] , \round_in[1][652] , \round_in[1][651] , 
        \round_in[1][650] , \round_in[1][649] , \round_in[1][648] , 
        \round_in[1][647] , \round_in[1][646] , \round_in[1][645] , 
        \round_in[1][644] , \round_in[1][643] , \round_in[1][642] , 
        \round_in[1][641] , \round_in[1][640] , \round_in[1][639] , 
        \round_in[1][638] , \round_in[1][637] , \round_in[1][636] , 
        \round_in[1][635] , \round_in[1][634] , \round_in[1][633] , 
        \round_in[1][632] , \round_in[1][631] , \round_in[1][630] , 
        \round_in[1][629] , \round_in[1][628] , \round_in[1][627] , 
        \round_in[1][626] , \round_in[1][625] , \round_in[1][624] , 
        \round_in[1][623] , \round_in[1][622] , \round_in[1][621] , 
        \round_in[1][620] , \round_in[1][619] , \round_in[1][618] , 
        \round_in[1][617] , \round_in[1][616] , \round_in[1][615] , 
        \round_in[1][614] , \round_in[1][613] , \round_in[1][612] , 
        \round_in[1][611] , \round_in[1][610] , \round_in[1][609] , 
        \round_in[1][608] , \round_in[1][607] , \round_in[1][606] , 
        \round_in[1][605] , \round_in[1][604] , \round_in[1][603] , 
        \round_in[1][602] , \round_in[1][601] , \round_in[1][600] , 
        \round_in[1][599] , \round_in[1][598] , \round_in[1][597] , 
        \round_in[1][596] , \round_in[1][595] , \round_in[1][594] , 
        \round_in[1][593] , \round_in[1][592] , \round_in[1][591] , 
        \round_in[1][590] , \round_in[1][589] , \round_in[1][588] , 
        \round_in[1][587] , \round_in[1][586] , \round_in[1][585] , 
        \round_in[1][584] , \round_in[1][583] , \round_in[1][582] , 
        \round_in[1][581] , \round_in[1][580] , \round_in[1][579] , 
        \round_in[1][578] , \round_in[1][577] , \round_in[1][576] , 
        \round_in[1][575] , \round_in[1][574] , \round_in[1][573] , 
        \round_in[1][572] , \round_in[1][571] , \round_in[1][570] , 
        \round_in[1][569] , \round_in[1][568] , \round_in[1][567] , 
        \round_in[1][566] , \round_in[1][565] , \round_in[1][564] , 
        \round_in[1][563] , \round_in[1][562] , \round_in[1][561] , 
        \round_in[1][560] , \round_in[1][559] , \round_in[1][558] , 
        \round_in[1][557] , \round_in[1][556] , \round_in[1][555] , 
        \round_in[1][554] , \round_in[1][553] , \round_in[1][552] , 
        \round_in[1][551] , \round_in[1][550] , \round_in[1][549] , 
        \round_in[1][548] , \round_in[1][547] , \round_in[1][546] , 
        \round_in[1][545] , \round_in[1][544] , \round_in[1][543] , 
        \round_in[1][542] , \round_in[1][541] , \round_in[1][540] , 
        \round_in[1][539] , \round_in[1][538] , \round_in[1][537] , 
        \round_in[1][536] , \round_in[1][535] , \round_in[1][534] , 
        \round_in[1][533] , \round_in[1][532] , \round_in[1][531] , 
        \round_in[1][530] , \round_in[1][529] , \round_in[1][528] , 
        \round_in[1][527] , \round_in[1][526] , \round_in[1][525] , 
        \round_in[1][524] , \round_in[1][523] , \round_in[1][522] , 
        \round_in[1][521] , \round_in[1][520] , \round_in[1][519] , 
        \round_in[1][518] , \round_in[1][517] , \round_in[1][516] , 
        \round_in[1][515] , \round_in[1][514] , \round_in[1][513] , 
        \round_in[1][512] , \round_in[1][511] , \round_in[1][510] , 
        \round_in[1][509] , \round_in[1][508] , \round_in[1][507] , 
        \round_in[1][506] , \round_in[1][505] , \round_in[1][504] , 
        \round_in[1][503] , \round_in[1][502] , \round_in[1][501] , 
        \round_in[1][500] , \round_in[1][499] , \round_in[1][498] , 
        \round_in[1][497] , \round_in[1][496] , \round_in[1][495] , 
        \round_in[1][494] , \round_in[1][493] , \round_in[1][492] , 
        \round_in[1][491] , \round_in[1][490] , \round_in[1][489] , 
        \round_in[1][488] , \round_in[1][487] , \round_in[1][486] , 
        \round_in[1][485] , \round_in[1][484] , \round_in[1][483] , 
        \round_in[1][482] , \round_in[1][481] , \round_in[1][480] , 
        \round_in[1][479] , \round_in[1][478] , \round_in[1][477] , 
        \round_in[1][476] , \round_in[1][475] , \round_in[1][474] , 
        \round_in[1][473] , \round_in[1][472] , \round_in[1][471] , 
        \round_in[1][470] , \round_in[1][469] , \round_in[1][468] , 
        \round_in[1][467] , \round_in[1][466] , \round_in[1][465] , 
        \round_in[1][464] , \round_in[1][463] , \round_in[1][462] , 
        \round_in[1][461] , \round_in[1][460] , \round_in[1][459] , 
        \round_in[1][458] , \round_in[1][457] , \round_in[1][456] , 
        \round_in[1][455] , \round_in[1][454] , \round_in[1][453] , 
        \round_in[1][452] , \round_in[1][451] , \round_in[1][450] , 
        \round_in[1][449] , \round_in[1][448] , \round_in[1][447] , 
        \round_in[1][446] , \round_in[1][445] , \round_in[1][444] , 
        \round_in[1][443] , \round_in[1][442] , \round_in[1][441] , 
        \round_in[1][440] , \round_in[1][439] , \round_in[1][438] , 
        \round_in[1][437] , \round_in[1][436] , \round_in[1][435] , 
        \round_in[1][434] , \round_in[1][433] , \round_in[1][432] , 
        \round_in[1][431] , \round_in[1][430] , \round_in[1][429] , 
        \round_in[1][428] , \round_in[1][427] , \round_in[1][426] , 
        \round_in[1][425] , \round_in[1][424] , \round_in[1][423] , 
        \round_in[1][422] , \round_in[1][421] , \round_in[1][420] , 
        \round_in[1][419] , \round_in[1][418] , \round_in[1][417] , 
        \round_in[1][416] , \round_in[1][415] , \round_in[1][414] , 
        \round_in[1][413] , \round_in[1][412] , \round_in[1][411] , 
        \round_in[1][410] , \round_in[1][409] , \round_in[1][408] , 
        \round_in[1][407] , \round_in[1][406] , \round_in[1][405] , 
        \round_in[1][404] , \round_in[1][403] , \round_in[1][402] , 
        \round_in[1][401] , \round_in[1][400] , \round_in[1][399] , 
        \round_in[1][398] , \round_in[1][397] , \round_in[1][396] , 
        \round_in[1][395] , \round_in[1][394] , \round_in[1][393] , 
        \round_in[1][392] , \round_in[1][391] , \round_in[1][390] , 
        \round_in[1][389] , \round_in[1][388] , \round_in[1][387] , 
        \round_in[1][386] , \round_in[1][385] , \round_in[1][384] , 
        \round_in[1][383] , \round_in[1][382] , \round_in[1][381] , 
        \round_in[1][380] , \round_in[1][379] , \round_in[1][378] , 
        \round_in[1][377] , \round_in[1][376] , \round_in[1][375] , 
        \round_in[1][374] , \round_in[1][373] , \round_in[1][372] , 
        \round_in[1][371] , \round_in[1][370] , \round_in[1][369] , 
        \round_in[1][368] , \round_in[1][367] , \round_in[1][366] , 
        \round_in[1][365] , \round_in[1][364] , \round_in[1][363] , 
        \round_in[1][362] , \round_in[1][361] , \round_in[1][360] , 
        \round_in[1][359] , \round_in[1][358] , \round_in[1][357] , 
        \round_in[1][356] , \round_in[1][355] , \round_in[1][354] , 
        \round_in[1][353] , \round_in[1][352] , \round_in[1][351] , 
        \round_in[1][350] , \round_in[1][349] , \round_in[1][348] , 
        \round_in[1][347] , \round_in[1][346] , \round_in[1][345] , 
        \round_in[1][344] , \round_in[1][343] , \round_in[1][342] , 
        \round_in[1][341] , \round_in[1][340] , \round_in[1][339] , 
        \round_in[1][338] , \round_in[1][337] , \round_in[1][336] , 
        \round_in[1][335] , \round_in[1][334] , \round_in[1][333] , 
        \round_in[1][332] , \round_in[1][331] , \round_in[1][330] , 
        \round_in[1][329] , \round_in[1][328] , \round_in[1][327] , 
        \round_in[1][326] , \round_in[1][325] , \round_in[1][324] , 
        \round_in[1][323] , \round_in[1][322] , \round_in[1][321] , 
        \round_in[1][320] , \round_in[1][319] , \round_in[1][318] , 
        \round_in[1][317] , \round_in[1][316] , \round_in[1][315] , 
        \round_in[1][314] , \round_in[1][313] , \round_in[1][312] , 
        \round_in[1][311] , \round_in[1][310] , \round_in[1][309] , 
        \round_in[1][308] , \round_in[1][307] , \round_in[1][306] , 
        \round_in[1][305] , \round_in[1][304] , \round_in[1][303] , 
        \round_in[1][302] , \round_in[1][301] , \round_in[1][300] , 
        \round_in[1][299] , \round_in[1][298] , \round_in[1][297] , 
        \round_in[1][296] , \round_in[1][295] , \round_in[1][294] , 
        \round_in[1][293] , \round_in[1][292] , \round_in[1][291] , 
        \round_in[1][290] , \round_in[1][289] , \round_in[1][288] , 
        \round_in[1][287] , \round_in[1][286] , \round_in[1][285] , 
        \round_in[1][284] , \round_in[1][283] , \round_in[1][282] , 
        \round_in[1][281] , \round_in[1][280] , \round_in[1][279] , 
        \round_in[1][278] , \round_in[1][277] , \round_in[1][276] , 
        \round_in[1][275] , \round_in[1][274] , \round_in[1][273] , 
        \round_in[1][272] , \round_in[1][271] , \round_in[1][270] , 
        \round_in[1][269] , \round_in[1][268] , \round_in[1][267] , 
        \round_in[1][266] , \round_in[1][265] , \round_in[1][264] , 
        \round_in[1][263] , \round_in[1][262] , \round_in[1][261] , 
        \round_in[1][260] , \round_in[1][259] , \round_in[1][258] , 
        \round_in[1][257] , \round_in[1][256] , \round_in[1][255] , 
        \round_in[1][254] , \round_in[1][253] , \round_in[1][252] , 
        \round_in[1][251] , \round_in[1][250] , \round_in[1][249] , 
        \round_in[1][248] , \round_in[1][247] , \round_in[1][246] , 
        \round_in[1][245] , \round_in[1][244] , \round_in[1][243] , 
        \round_in[1][242] , \round_in[1][241] , \round_in[1][240] , 
        \round_in[1][239] , \round_in[1][238] , \round_in[1][237] , 
        \round_in[1][236] , \round_in[1][235] , \round_in[1][234] , 
        \round_in[1][233] , \round_in[1][232] , \round_in[1][231] , 
        \round_in[1][230] , \round_in[1][229] , \round_in[1][228] , 
        \round_in[1][227] , \round_in[1][226] , \round_in[1][225] , 
        \round_in[1][224] , \round_in[1][223] , \round_in[1][222] , 
        \round_in[1][221] , \round_in[1][220] , \round_in[1][219] , 
        \round_in[1][218] , \round_in[1][217] , \round_in[1][216] , 
        \round_in[1][215] , \round_in[1][214] , \round_in[1][213] , 
        \round_in[1][212] , \round_in[1][211] , \round_in[1][210] , 
        \round_in[1][209] , \round_in[1][208] , \round_in[1][207] , 
        \round_in[1][206] , \round_in[1][205] , \round_in[1][204] , 
        \round_in[1][203] , \round_in[1][202] , \round_in[1][201] , 
        \round_in[1][200] , \round_in[1][199] , \round_in[1][198] , 
        \round_in[1][197] , \round_in[1][196] , \round_in[1][195] , 
        \round_in[1][194] , \round_in[1][193] , \round_in[1][192] , 
        \round_in[1][191] , \round_in[1][190] , \round_in[1][189] , 
        \round_in[1][188] , \round_in[1][187] , \round_in[1][186] , 
        \round_in[1][185] , \round_in[1][184] , \round_in[1][183] , 
        \round_in[1][182] , \round_in[1][181] , \round_in[1][180] , 
        \round_in[1][179] , \round_in[1][178] , \round_in[1][177] , 
        \round_in[1][176] , \round_in[1][175] , \round_in[1][174] , 
        \round_in[1][173] , \round_in[1][172] , \round_in[1][171] , 
        \round_in[1][170] , \round_in[1][169] , \round_in[1][168] , 
        \round_in[1][167] , \round_in[1][166] , \round_in[1][165] , 
        \round_in[1][164] , \round_in[1][163] , \round_in[1][162] , 
        \round_in[1][161] , \round_in[1][160] , \round_in[1][159] , 
        \round_in[1][158] , \round_in[1][157] , \round_in[1][156] , 
        \round_in[1][155] , \round_in[1][154] , \round_in[1][153] , 
        \round_in[1][152] , \round_in[1][151] , \round_in[1][150] , 
        \round_in[1][149] , \round_in[1][148] , \round_in[1][147] , 
        \round_in[1][146] , \round_in[1][145] , \round_in[1][144] , 
        \round_in[1][143] , \round_in[1][142] , \round_in[1][141] , 
        \round_in[1][140] , \round_in[1][139] , \round_in[1][138] , 
        \round_in[1][137] , \round_in[1][136] , \round_in[1][135] , 
        \round_in[1][134] , \round_in[1][133] , \round_in[1][132] , 
        \round_in[1][131] , \round_in[1][130] , \round_in[1][129] , 
        \round_in[1][128] , \round_in[1][127] , \round_in[1][126] , 
        \round_in[1][125] , \round_in[1][124] , \round_in[1][123] , 
        \round_in[1][122] , \round_in[1][121] , \round_in[1][120] , 
        \round_in[1][119] , \round_in[1][118] , \round_in[1][117] , 
        \round_in[1][116] , \round_in[1][115] , \round_in[1][114] , 
        \round_in[1][113] , \round_in[1][112] , \round_in[1][111] , 
        \round_in[1][110] , \round_in[1][109] , \round_in[1][108] , 
        \round_in[1][107] , \round_in[1][106] , \round_in[1][105] , 
        \round_in[1][104] , \round_in[1][103] , \round_in[1][102] , 
        \round_in[1][101] , \round_in[1][100] , \round_in[1][99] , 
        \round_in[1][98] , \round_in[1][97] , \round_in[1][96] , 
        \round_in[1][95] , \round_in[1][94] , \round_in[1][93] , 
        \round_in[1][92] , \round_in[1][91] , \round_in[1][90] , 
        \round_in[1][89] , \round_in[1][88] , \round_in[1][87] , 
        \round_in[1][86] , \round_in[1][85] , \round_in[1][84] , 
        \round_in[1][83] , \round_in[1][82] , \round_in[1][81] , 
        \round_in[1][80] , \round_in[1][79] , \round_in[1][78] , 
        \round_in[1][77] , \round_in[1][76] , \round_in[1][75] , 
        \round_in[1][74] , \round_in[1][73] , \round_in[1][72] , 
        \round_in[1][71] , \round_in[1][70] , \round_in[1][69] , 
        \round_in[1][68] , \round_in[1][67] , \round_in[1][66] , 
        \round_in[1][65] , \round_in[1][64] , \round_in[1][63] , 
        \round_in[1][62] , \round_in[1][61] , \round_in[1][60] , 
        \round_in[1][59] , \round_in[1][58] , \round_in[1][57] , 
        \round_in[1][56] , \round_in[1][55] , \round_in[1][54] , 
        \round_in[1][53] , \round_in[1][52] , \round_in[1][51] , 
        \round_in[1][50] , \round_in[1][49] , \round_in[1][48] , 
        \round_in[1][47] , \round_in[1][46] , \round_in[1][45] , 
        \round_in[1][44] , \round_in[1][43] , \round_in[1][42] , 
        \round_in[1][41] , \round_in[1][40] , \round_in[1][39] , 
        \round_in[1][38] , \round_in[1][37] , \round_in[1][36] , 
        \round_in[1][35] , \round_in[1][34] , \round_in[1][33] , 
        \round_in[1][32] , \round_in[1][31] , \round_in[1][30] , 
        \round_in[1][29] , \round_in[1][28] , \round_in[1][27] , 
        \round_in[1][26] , \round_in[1][25] , \round_in[1][24] , 
        \round_in[1][23] , \round_in[1][22] , \round_in[1][21] , 
        \round_in[1][20] , \round_in[1][19] , \round_in[1][18] , 
        \round_in[1][17] , \round_in[1][16] , \round_in[1][15] , 
        \round_in[1][14] , \round_in[1][13] , \round_in[1][12] , 
        \round_in[1][11] , \round_in[1][10] , \round_in[1][9] , 
        \round_in[1][8] , \round_in[1][7] , \round_in[1][6] , \round_in[1][5] , 
        \round_in[1][4] , \round_in[1][3] , \round_in[1][2] , \round_in[1][1] , 
        \round_in[1][0] }) );
  round_1 \ROUND[1].round_  ( .in({\round_in[1][1599] , \round_in[1][1598] , 
        \round_in[1][1597] , \round_in[1][1596] , \round_in[1][1595] , 
        \round_in[1][1594] , \round_in[1][1593] , \round_in[1][1592] , 
        \round_in[1][1591] , \round_in[1][1590] , \round_in[1][1589] , 
        \round_in[1][1588] , \round_in[1][1587] , \round_in[1][1586] , 
        \round_in[1][1585] , \round_in[1][1584] , \round_in[1][1583] , 
        \round_in[1][1582] , \round_in[1][1581] , \round_in[1][1580] , 
        \round_in[1][1579] , \round_in[1][1578] , \round_in[1][1577] , 
        \round_in[1][1576] , \round_in[1][1575] , \round_in[1][1574] , 
        \round_in[1][1573] , \round_in[1][1572] , \round_in[1][1571] , 
        \round_in[1][1570] , \round_in[1][1569] , \round_in[1][1568] , 
        \round_in[1][1567] , \round_in[1][1566] , \round_in[1][1565] , 
        \round_in[1][1564] , \round_in[1][1563] , \round_in[1][1562] , 
        \round_in[1][1561] , \round_in[1][1560] , \round_in[1][1559] , 
        \round_in[1][1558] , \round_in[1][1557] , \round_in[1][1556] , 
        \round_in[1][1555] , \round_in[1][1554] , \round_in[1][1553] , 
        \round_in[1][1552] , \round_in[1][1551] , \round_in[1][1550] , 
        \round_in[1][1549] , \round_in[1][1548] , \round_in[1][1547] , 
        \round_in[1][1546] , \round_in[1][1545] , \round_in[1][1544] , 
        \round_in[1][1543] , \round_in[1][1542] , \round_in[1][1541] , 
        \round_in[1][1540] , \round_in[1][1539] , \round_in[1][1538] , 
        \round_in[1][1537] , \round_in[1][1536] , \round_in[1][1535] , 
        \round_in[1][1534] , \round_in[1][1533] , \round_in[1][1532] , 
        \round_in[1][1531] , \round_in[1][1530] , \round_in[1][1529] , 
        \round_in[1][1528] , \round_in[1][1527] , \round_in[1][1526] , 
        \round_in[1][1525] , \round_in[1][1524] , \round_in[1][1523] , 
        \round_in[1][1522] , \round_in[1][1521] , \round_in[1][1520] , 
        \round_in[1][1519] , \round_in[1][1518] , \round_in[1][1517] , 
        \round_in[1][1516] , \round_in[1][1515] , \round_in[1][1514] , 
        \round_in[1][1513] , \round_in[1][1512] , \round_in[1][1511] , 
        \round_in[1][1510] , \round_in[1][1509] , \round_in[1][1508] , 
        \round_in[1][1507] , \round_in[1][1506] , \round_in[1][1505] , 
        \round_in[1][1504] , \round_in[1][1503] , \round_in[1][1502] , 
        \round_in[1][1501] , \round_in[1][1500] , \round_in[1][1499] , 
        \round_in[1][1498] , \round_in[1][1497] , \round_in[1][1496] , 
        \round_in[1][1495] , \round_in[1][1494] , \round_in[1][1493] , 
        \round_in[1][1492] , \round_in[1][1491] , \round_in[1][1490] , 
        \round_in[1][1489] , \round_in[1][1488] , \round_in[1][1487] , 
        \round_in[1][1486] , \round_in[1][1485] , \round_in[1][1484] , 
        \round_in[1][1483] , \round_in[1][1482] , \round_in[1][1481] , 
        \round_in[1][1480] , \round_in[1][1479] , \round_in[1][1478] , 
        \round_in[1][1477] , \round_in[1][1476] , \round_in[1][1475] , 
        \round_in[1][1474] , \round_in[1][1473] , \round_in[1][1472] , 
        \round_in[1][1471] , \round_in[1][1470] , \round_in[1][1469] , 
        \round_in[1][1468] , \round_in[1][1467] , \round_in[1][1466] , 
        \round_in[1][1465] , \round_in[1][1464] , \round_in[1][1463] , 
        \round_in[1][1462] , \round_in[1][1461] , \round_in[1][1460] , 
        \round_in[1][1459] , \round_in[1][1458] , \round_in[1][1457] , 
        \round_in[1][1456] , \round_in[1][1455] , \round_in[1][1454] , 
        \round_in[1][1453] , \round_in[1][1452] , \round_in[1][1451] , 
        \round_in[1][1450] , \round_in[1][1449] , \round_in[1][1448] , 
        \round_in[1][1447] , \round_in[1][1446] , \round_in[1][1445] , 
        \round_in[1][1444] , \round_in[1][1443] , \round_in[1][1442] , 
        \round_in[1][1441] , \round_in[1][1440] , \round_in[1][1439] , 
        \round_in[1][1438] , \round_in[1][1437] , \round_in[1][1436] , 
        \round_in[1][1435] , \round_in[1][1434] , \round_in[1][1433] , 
        \round_in[1][1432] , \round_in[1][1431] , \round_in[1][1430] , 
        \round_in[1][1429] , \round_in[1][1428] , \round_in[1][1427] , 
        \round_in[1][1426] , \round_in[1][1425] , \round_in[1][1424] , 
        \round_in[1][1423] , \round_in[1][1422] , \round_in[1][1421] , 
        \round_in[1][1420] , \round_in[1][1419] , \round_in[1][1418] , 
        \round_in[1][1417] , \round_in[1][1416] , \round_in[1][1415] , 
        \round_in[1][1414] , \round_in[1][1413] , \round_in[1][1412] , 
        \round_in[1][1411] , \round_in[1][1410] , \round_in[1][1409] , 
        \round_in[1][1408] , \round_in[1][1407] , \round_in[1][1406] , 
        \round_in[1][1405] , \round_in[1][1404] , \round_in[1][1403] , 
        \round_in[1][1402] , \round_in[1][1401] , \round_in[1][1400] , 
        \round_in[1][1399] , \round_in[1][1398] , \round_in[1][1397] , 
        \round_in[1][1396] , \round_in[1][1395] , \round_in[1][1394] , 
        \round_in[1][1393] , \round_in[1][1392] , \round_in[1][1391] , 
        \round_in[1][1390] , \round_in[1][1389] , \round_in[1][1388] , 
        \round_in[1][1387] , \round_in[1][1386] , \round_in[1][1385] , 
        \round_in[1][1384] , \round_in[1][1383] , \round_in[1][1382] , 
        \round_in[1][1381] , \round_in[1][1380] , \round_in[1][1379] , 
        \round_in[1][1378] , \round_in[1][1377] , \round_in[1][1376] , 
        \round_in[1][1375] , \round_in[1][1374] , \round_in[1][1373] , 
        \round_in[1][1372] , \round_in[1][1371] , \round_in[1][1370] , 
        \round_in[1][1369] , \round_in[1][1368] , \round_in[1][1367] , 
        \round_in[1][1366] , \round_in[1][1365] , \round_in[1][1364] , 
        \round_in[1][1363] , \round_in[1][1362] , \round_in[1][1361] , 
        \round_in[1][1360] , \round_in[1][1359] , \round_in[1][1358] , 
        \round_in[1][1357] , \round_in[1][1356] , \round_in[1][1355] , 
        \round_in[1][1354] , \round_in[1][1353] , \round_in[1][1352] , 
        \round_in[1][1351] , \round_in[1][1350] , \round_in[1][1349] , 
        \round_in[1][1348] , \round_in[1][1347] , \round_in[1][1346] , 
        \round_in[1][1345] , \round_in[1][1344] , \round_in[1][1343] , 
        \round_in[1][1342] , \round_in[1][1341] , \round_in[1][1340] , 
        \round_in[1][1339] , \round_in[1][1338] , \round_in[1][1337] , 
        \round_in[1][1336] , \round_in[1][1335] , \round_in[1][1334] , 
        \round_in[1][1333] , \round_in[1][1332] , \round_in[1][1331] , 
        \round_in[1][1330] , \round_in[1][1329] , \round_in[1][1328] , 
        \round_in[1][1327] , \round_in[1][1326] , \round_in[1][1325] , 
        \round_in[1][1324] , \round_in[1][1323] , \round_in[1][1322] , 
        \round_in[1][1321] , \round_in[1][1320] , \round_in[1][1319] , 
        \round_in[1][1318] , \round_in[1][1317] , \round_in[1][1316] , 
        \round_in[1][1315] , \round_in[1][1314] , \round_in[1][1313] , 
        \round_in[1][1312] , \round_in[1][1311] , \round_in[1][1310] , 
        \round_in[1][1309] , \round_in[1][1308] , \round_in[1][1307] , 
        \round_in[1][1306] , \round_in[1][1305] , \round_in[1][1304] , 
        \round_in[1][1303] , \round_in[1][1302] , \round_in[1][1301] , 
        \round_in[1][1300] , \round_in[1][1299] , \round_in[1][1298] , 
        \round_in[1][1297] , \round_in[1][1296] , \round_in[1][1295] , 
        \round_in[1][1294] , \round_in[1][1293] , \round_in[1][1292] , 
        \round_in[1][1291] , \round_in[1][1290] , \round_in[1][1289] , 
        \round_in[1][1288] , \round_in[1][1287] , \round_in[1][1286] , 
        \round_in[1][1285] , \round_in[1][1284] , \round_in[1][1283] , 
        \round_in[1][1282] , \round_in[1][1281] , \round_in[1][1280] , 
        \round_in[1][1279] , \round_in[1][1278] , \round_in[1][1277] , 
        \round_in[1][1276] , \round_in[1][1275] , \round_in[1][1274] , 
        \round_in[1][1273] , \round_in[1][1272] , \round_in[1][1271] , 
        \round_in[1][1270] , \round_in[1][1269] , \round_in[1][1268] , 
        \round_in[1][1267] , \round_in[1][1266] , \round_in[1][1265] , 
        \round_in[1][1264] , \round_in[1][1263] , \round_in[1][1262] , 
        \round_in[1][1261] , \round_in[1][1260] , \round_in[1][1259] , 
        \round_in[1][1258] , \round_in[1][1257] , \round_in[1][1256] , 
        \round_in[1][1255] , \round_in[1][1254] , \round_in[1][1253] , 
        \round_in[1][1252] , \round_in[1][1251] , \round_in[1][1250] , 
        \round_in[1][1249] , \round_in[1][1248] , \round_in[1][1247] , 
        \round_in[1][1246] , \round_in[1][1245] , \round_in[1][1244] , 
        \round_in[1][1243] , \round_in[1][1242] , \round_in[1][1241] , 
        \round_in[1][1240] , \round_in[1][1239] , \round_in[1][1238] , 
        \round_in[1][1237] , \round_in[1][1236] , \round_in[1][1235] , 
        \round_in[1][1234] , \round_in[1][1233] , \round_in[1][1232] , 
        \round_in[1][1231] , \round_in[1][1230] , \round_in[1][1229] , 
        \round_in[1][1228] , \round_in[1][1227] , \round_in[1][1226] , 
        \round_in[1][1225] , \round_in[1][1224] , \round_in[1][1223] , 
        \round_in[1][1222] , \round_in[1][1221] , \round_in[1][1220] , 
        \round_in[1][1219] , \round_in[1][1218] , \round_in[1][1217] , 
        \round_in[1][1216] , \round_in[1][1215] , \round_in[1][1214] , 
        \round_in[1][1213] , \round_in[1][1212] , \round_in[1][1211] , 
        \round_in[1][1210] , \round_in[1][1209] , \round_in[1][1208] , 
        \round_in[1][1207] , \round_in[1][1206] , \round_in[1][1205] , 
        \round_in[1][1204] , \round_in[1][1203] , \round_in[1][1202] , 
        \round_in[1][1201] , \round_in[1][1200] , \round_in[1][1199] , 
        \round_in[1][1198] , \round_in[1][1197] , \round_in[1][1196] , 
        \round_in[1][1195] , \round_in[1][1194] , \round_in[1][1193] , 
        \round_in[1][1192] , \round_in[1][1191] , \round_in[1][1190] , 
        \round_in[1][1189] , \round_in[1][1188] , \round_in[1][1187] , 
        \round_in[1][1186] , \round_in[1][1185] , \round_in[1][1184] , 
        \round_in[1][1183] , \round_in[1][1182] , \round_in[1][1181] , 
        \round_in[1][1180] , \round_in[1][1179] , \round_in[1][1178] , 
        \round_in[1][1177] , \round_in[1][1176] , \round_in[1][1175] , 
        \round_in[1][1174] , \round_in[1][1173] , \round_in[1][1172] , 
        \round_in[1][1171] , \round_in[1][1170] , \round_in[1][1169] , 
        \round_in[1][1168] , \round_in[1][1167] , \round_in[1][1166] , 
        \round_in[1][1165] , \round_in[1][1164] , \round_in[1][1163] , 
        \round_in[1][1162] , \round_in[1][1161] , \round_in[1][1160] , 
        \round_in[1][1159] , \round_in[1][1158] , \round_in[1][1157] , 
        \round_in[1][1156] , \round_in[1][1155] , \round_in[1][1154] , 
        \round_in[1][1153] , \round_in[1][1152] , \round_in[1][1151] , 
        \round_in[1][1150] , \round_in[1][1149] , \round_in[1][1148] , 
        \round_in[1][1147] , \round_in[1][1146] , \round_in[1][1145] , 
        \round_in[1][1144] , \round_in[1][1143] , \round_in[1][1142] , 
        \round_in[1][1141] , \round_in[1][1140] , \round_in[1][1139] , 
        \round_in[1][1138] , \round_in[1][1137] , \round_in[1][1136] , 
        \round_in[1][1135] , \round_in[1][1134] , \round_in[1][1133] , 
        \round_in[1][1132] , \round_in[1][1131] , \round_in[1][1130] , 
        \round_in[1][1129] , \round_in[1][1128] , \round_in[1][1127] , 
        \round_in[1][1126] , \round_in[1][1125] , \round_in[1][1124] , 
        \round_in[1][1123] , \round_in[1][1122] , \round_in[1][1121] , 
        \round_in[1][1120] , \round_in[1][1119] , \round_in[1][1118] , 
        \round_in[1][1117] , \round_in[1][1116] , \round_in[1][1115] , 
        \round_in[1][1114] , \round_in[1][1113] , \round_in[1][1112] , 
        \round_in[1][1111] , \round_in[1][1110] , \round_in[1][1109] , 
        \round_in[1][1108] , \round_in[1][1107] , \round_in[1][1106] , 
        \round_in[1][1105] , \round_in[1][1104] , \round_in[1][1103] , 
        \round_in[1][1102] , \round_in[1][1101] , \round_in[1][1100] , 
        \round_in[1][1099] , \round_in[1][1098] , \round_in[1][1097] , 
        \round_in[1][1096] , \round_in[1][1095] , \round_in[1][1094] , 
        \round_in[1][1093] , \round_in[1][1092] , \round_in[1][1091] , 
        \round_in[1][1090] , \round_in[1][1089] , \round_in[1][1088] , 
        \round_in[1][1087] , \round_in[1][1086] , \round_in[1][1085] , 
        \round_in[1][1084] , \round_in[1][1083] , \round_in[1][1082] , 
        \round_in[1][1081] , \round_in[1][1080] , \round_in[1][1079] , 
        \round_in[1][1078] , \round_in[1][1077] , \round_in[1][1076] , 
        \round_in[1][1075] , \round_in[1][1074] , \round_in[1][1073] , 
        \round_in[1][1072] , \round_in[1][1071] , \round_in[1][1070] , 
        \round_in[1][1069] , \round_in[1][1068] , \round_in[1][1067] , 
        \round_in[1][1066] , \round_in[1][1065] , \round_in[1][1064] , 
        \round_in[1][1063] , \round_in[1][1062] , \round_in[1][1061] , 
        \round_in[1][1060] , \round_in[1][1059] , \round_in[1][1058] , 
        \round_in[1][1057] , \round_in[1][1056] , \round_in[1][1055] , 
        \round_in[1][1054] , \round_in[1][1053] , \round_in[1][1052] , 
        \round_in[1][1051] , \round_in[1][1050] , \round_in[1][1049] , 
        \round_in[1][1048] , \round_in[1][1047] , \round_in[1][1046] , 
        \round_in[1][1045] , \round_in[1][1044] , \round_in[1][1043] , 
        \round_in[1][1042] , \round_in[1][1041] , \round_in[1][1040] , 
        \round_in[1][1039] , \round_in[1][1038] , \round_in[1][1037] , 
        \round_in[1][1036] , \round_in[1][1035] , \round_in[1][1034] , 
        \round_in[1][1033] , \round_in[1][1032] , \round_in[1][1031] , 
        \round_in[1][1030] , \round_in[1][1029] , \round_in[1][1028] , 
        \round_in[1][1027] , \round_in[1][1026] , \round_in[1][1025] , 
        \round_in[1][1024] , \round_in[1][1023] , \round_in[1][1022] , 
        \round_in[1][1021] , \round_in[1][1020] , \round_in[1][1019] , 
        \round_in[1][1018] , \round_in[1][1017] , \round_in[1][1016] , 
        \round_in[1][1015] , \round_in[1][1014] , \round_in[1][1013] , 
        \round_in[1][1012] , \round_in[1][1011] , \round_in[1][1010] , 
        \round_in[1][1009] , \round_in[1][1008] , \round_in[1][1007] , 
        \round_in[1][1006] , \round_in[1][1005] , \round_in[1][1004] , 
        \round_in[1][1003] , \round_in[1][1002] , \round_in[1][1001] , 
        \round_in[1][1000] , \round_in[1][999] , \round_in[1][998] , 
        \round_in[1][997] , \round_in[1][996] , \round_in[1][995] , 
        \round_in[1][994] , \round_in[1][993] , \round_in[1][992] , 
        \round_in[1][991] , \round_in[1][990] , \round_in[1][989] , 
        \round_in[1][988] , \round_in[1][987] , \round_in[1][986] , 
        \round_in[1][985] , \round_in[1][984] , \round_in[1][983] , 
        \round_in[1][982] , \round_in[1][981] , \round_in[1][980] , 
        \round_in[1][979] , \round_in[1][978] , \round_in[1][977] , 
        \round_in[1][976] , \round_in[1][975] , \round_in[1][974] , 
        \round_in[1][973] , \round_in[1][972] , \round_in[1][971] , 
        \round_in[1][970] , \round_in[1][969] , \round_in[1][968] , 
        \round_in[1][967] , \round_in[1][966] , \round_in[1][965] , 
        \round_in[1][964] , \round_in[1][963] , \round_in[1][962] , 
        \round_in[1][961] , \round_in[1][960] , \round_in[1][959] , 
        \round_in[1][958] , \round_in[1][957] , \round_in[1][956] , 
        \round_in[1][955] , \round_in[1][954] , \round_in[1][953] , 
        \round_in[1][952] , \round_in[1][951] , \round_in[1][950] , 
        \round_in[1][949] , \round_in[1][948] , \round_in[1][947] , 
        \round_in[1][946] , \round_in[1][945] , \round_in[1][944] , 
        \round_in[1][943] , \round_in[1][942] , \round_in[1][941] , 
        \round_in[1][940] , \round_in[1][939] , \round_in[1][938] , 
        \round_in[1][937] , \round_in[1][936] , \round_in[1][935] , 
        \round_in[1][934] , \round_in[1][933] , \round_in[1][932] , 
        \round_in[1][931] , \round_in[1][930] , \round_in[1][929] , 
        \round_in[1][928] , \round_in[1][927] , \round_in[1][926] , 
        \round_in[1][925] , \round_in[1][924] , \round_in[1][923] , 
        \round_in[1][922] , \round_in[1][921] , \round_in[1][920] , 
        \round_in[1][919] , \round_in[1][918] , \round_in[1][917] , 
        \round_in[1][916] , \round_in[1][915] , \round_in[1][914] , 
        \round_in[1][913] , \round_in[1][912] , \round_in[1][911] , 
        \round_in[1][910] , \round_in[1][909] , \round_in[1][908] , 
        \round_in[1][907] , \round_in[1][906] , \round_in[1][905] , 
        \round_in[1][904] , \round_in[1][903] , \round_in[1][902] , 
        \round_in[1][901] , \round_in[1][900] , \round_in[1][899] , 
        \round_in[1][898] , \round_in[1][897] , \round_in[1][896] , 
        \round_in[1][895] , \round_in[1][894] , \round_in[1][893] , 
        \round_in[1][892] , \round_in[1][891] , \round_in[1][890] , 
        \round_in[1][889] , \round_in[1][888] , \round_in[1][887] , 
        \round_in[1][886] , \round_in[1][885] , \round_in[1][884] , 
        \round_in[1][883] , \round_in[1][882] , \round_in[1][881] , 
        \round_in[1][880] , \round_in[1][879] , \round_in[1][878] , 
        \round_in[1][877] , \round_in[1][876] , \round_in[1][875] , 
        \round_in[1][874] , \round_in[1][873] , \round_in[1][872] , 
        \round_in[1][871] , \round_in[1][870] , \round_in[1][869] , 
        \round_in[1][868] , \round_in[1][867] , \round_in[1][866] , 
        \round_in[1][865] , \round_in[1][864] , \round_in[1][863] , 
        \round_in[1][862] , \round_in[1][861] , \round_in[1][860] , 
        \round_in[1][859] , \round_in[1][858] , \round_in[1][857] , 
        \round_in[1][856] , \round_in[1][855] , \round_in[1][854] , 
        \round_in[1][853] , \round_in[1][852] , \round_in[1][851] , 
        \round_in[1][850] , \round_in[1][849] , \round_in[1][848] , 
        \round_in[1][847] , \round_in[1][846] , \round_in[1][845] , 
        \round_in[1][844] , \round_in[1][843] , \round_in[1][842] , 
        \round_in[1][841] , \round_in[1][840] , \round_in[1][839] , 
        \round_in[1][838] , \round_in[1][837] , \round_in[1][836] , 
        \round_in[1][835] , \round_in[1][834] , \round_in[1][833] , 
        \round_in[1][832] , \round_in[1][831] , \round_in[1][830] , 
        \round_in[1][829] , \round_in[1][828] , \round_in[1][827] , 
        \round_in[1][826] , \round_in[1][825] , \round_in[1][824] , 
        \round_in[1][823] , \round_in[1][822] , \round_in[1][821] , 
        \round_in[1][820] , \round_in[1][819] , \round_in[1][818] , 
        \round_in[1][817] , \round_in[1][816] , \round_in[1][815] , 
        \round_in[1][814] , \round_in[1][813] , \round_in[1][812] , 
        \round_in[1][811] , \round_in[1][810] , \round_in[1][809] , 
        \round_in[1][808] , \round_in[1][807] , \round_in[1][806] , 
        \round_in[1][805] , \round_in[1][804] , \round_in[1][803] , 
        \round_in[1][802] , \round_in[1][801] , \round_in[1][800] , 
        \round_in[1][799] , \round_in[1][798] , \round_in[1][797] , 
        \round_in[1][796] , \round_in[1][795] , \round_in[1][794] , 
        \round_in[1][793] , \round_in[1][792] , \round_in[1][791] , 
        \round_in[1][790] , \round_in[1][789] , \round_in[1][788] , 
        \round_in[1][787] , \round_in[1][786] , \round_in[1][785] , 
        \round_in[1][784] , \round_in[1][783] , \round_in[1][782] , 
        \round_in[1][781] , \round_in[1][780] , \round_in[1][779] , 
        \round_in[1][778] , \round_in[1][777] , \round_in[1][776] , 
        \round_in[1][775] , \round_in[1][774] , \round_in[1][773] , 
        \round_in[1][772] , \round_in[1][771] , \round_in[1][770] , 
        \round_in[1][769] , \round_in[1][768] , \round_in[1][767] , 
        \round_in[1][766] , \round_in[1][765] , \round_in[1][764] , 
        \round_in[1][763] , \round_in[1][762] , \round_in[1][761] , 
        \round_in[1][760] , \round_in[1][759] , \round_in[1][758] , 
        \round_in[1][757] , \round_in[1][756] , \round_in[1][755] , 
        \round_in[1][754] , \round_in[1][753] , \round_in[1][752] , 
        \round_in[1][751] , \round_in[1][750] , \round_in[1][749] , 
        \round_in[1][748] , \round_in[1][747] , \round_in[1][746] , 
        \round_in[1][745] , \round_in[1][744] , \round_in[1][743] , 
        \round_in[1][742] , \round_in[1][741] , \round_in[1][740] , 
        \round_in[1][739] , \round_in[1][738] , \round_in[1][737] , 
        \round_in[1][736] , \round_in[1][735] , \round_in[1][734] , 
        \round_in[1][733] , \round_in[1][732] , \round_in[1][731] , 
        \round_in[1][730] , \round_in[1][729] , \round_in[1][728] , 
        \round_in[1][727] , \round_in[1][726] , \round_in[1][725] , 
        \round_in[1][724] , \round_in[1][723] , \round_in[1][722] , 
        \round_in[1][721] , \round_in[1][720] , \round_in[1][719] , 
        \round_in[1][718] , \round_in[1][717] , \round_in[1][716] , 
        \round_in[1][715] , \round_in[1][714] , \round_in[1][713] , 
        \round_in[1][712] , \round_in[1][711] , \round_in[1][710] , 
        \round_in[1][709] , \round_in[1][708] , \round_in[1][707] , 
        \round_in[1][706] , \round_in[1][705] , \round_in[1][704] , 
        \round_in[1][703] , \round_in[1][702] , \round_in[1][701] , 
        \round_in[1][700] , \round_in[1][699] , \round_in[1][698] , 
        \round_in[1][697] , \round_in[1][696] , \round_in[1][695] , 
        \round_in[1][694] , \round_in[1][693] , \round_in[1][692] , 
        \round_in[1][691] , \round_in[1][690] , \round_in[1][689] , 
        \round_in[1][688] , \round_in[1][687] , \round_in[1][686] , 
        \round_in[1][685] , \round_in[1][684] , \round_in[1][683] , 
        \round_in[1][682] , \round_in[1][681] , \round_in[1][680] , 
        \round_in[1][679] , \round_in[1][678] , \round_in[1][677] , 
        \round_in[1][676] , \round_in[1][675] , \round_in[1][674] , 
        \round_in[1][673] , \round_in[1][672] , \round_in[1][671] , 
        \round_in[1][670] , \round_in[1][669] , \round_in[1][668] , 
        \round_in[1][667] , \round_in[1][666] , \round_in[1][665] , 
        \round_in[1][664] , \round_in[1][663] , \round_in[1][662] , 
        \round_in[1][661] , \round_in[1][660] , \round_in[1][659] , 
        \round_in[1][658] , \round_in[1][657] , \round_in[1][656] , 
        \round_in[1][655] , \round_in[1][654] , \round_in[1][653] , 
        \round_in[1][652] , \round_in[1][651] , \round_in[1][650] , 
        \round_in[1][649] , \round_in[1][648] , \round_in[1][647] , 
        \round_in[1][646] , \round_in[1][645] , \round_in[1][644] , 
        \round_in[1][643] , \round_in[1][642] , \round_in[1][641] , 
        \round_in[1][640] , \round_in[1][639] , \round_in[1][638] , 
        \round_in[1][637] , \round_in[1][636] , \round_in[1][635] , 
        \round_in[1][634] , \round_in[1][633] , \round_in[1][632] , 
        \round_in[1][631] , \round_in[1][630] , \round_in[1][629] , 
        \round_in[1][628] , \round_in[1][627] , \round_in[1][626] , 
        \round_in[1][625] , \round_in[1][624] , \round_in[1][623] , 
        \round_in[1][622] , \round_in[1][621] , \round_in[1][620] , 
        \round_in[1][619] , \round_in[1][618] , \round_in[1][617] , 
        \round_in[1][616] , \round_in[1][615] , \round_in[1][614] , 
        \round_in[1][613] , \round_in[1][612] , \round_in[1][611] , 
        \round_in[1][610] , \round_in[1][609] , \round_in[1][608] , 
        \round_in[1][607] , \round_in[1][606] , \round_in[1][605] , 
        \round_in[1][604] , \round_in[1][603] , \round_in[1][602] , 
        \round_in[1][601] , \round_in[1][600] , \round_in[1][599] , 
        \round_in[1][598] , \round_in[1][597] , \round_in[1][596] , 
        \round_in[1][595] , \round_in[1][594] , \round_in[1][593] , 
        \round_in[1][592] , \round_in[1][591] , \round_in[1][590] , 
        \round_in[1][589] , \round_in[1][588] , \round_in[1][587] , 
        \round_in[1][586] , \round_in[1][585] , \round_in[1][584] , 
        \round_in[1][583] , \round_in[1][582] , \round_in[1][581] , 
        \round_in[1][580] , \round_in[1][579] , \round_in[1][578] , 
        \round_in[1][577] , \round_in[1][576] , \round_in[1][575] , 
        \round_in[1][574] , \round_in[1][573] , \round_in[1][572] , 
        \round_in[1][571] , \round_in[1][570] , \round_in[1][569] , 
        \round_in[1][568] , \round_in[1][567] , \round_in[1][566] , 
        \round_in[1][565] , \round_in[1][564] , \round_in[1][563] , 
        \round_in[1][562] , \round_in[1][561] , \round_in[1][560] , 
        \round_in[1][559] , \round_in[1][558] , \round_in[1][557] , 
        \round_in[1][556] , \round_in[1][555] , \round_in[1][554] , 
        \round_in[1][553] , \round_in[1][552] , \round_in[1][551] , 
        \round_in[1][550] , \round_in[1][549] , \round_in[1][548] , 
        \round_in[1][547] , \round_in[1][546] , \round_in[1][545] , 
        \round_in[1][544] , \round_in[1][543] , \round_in[1][542] , 
        \round_in[1][541] , \round_in[1][540] , \round_in[1][539] , 
        \round_in[1][538] , \round_in[1][537] , \round_in[1][536] , 
        \round_in[1][535] , \round_in[1][534] , \round_in[1][533] , 
        \round_in[1][532] , \round_in[1][531] , \round_in[1][530] , 
        \round_in[1][529] , \round_in[1][528] , \round_in[1][527] , 
        \round_in[1][526] , \round_in[1][525] , \round_in[1][524] , 
        \round_in[1][523] , \round_in[1][522] , \round_in[1][521] , 
        \round_in[1][520] , \round_in[1][519] , \round_in[1][518] , 
        \round_in[1][517] , \round_in[1][516] , \round_in[1][515] , 
        \round_in[1][514] , \round_in[1][513] , \round_in[1][512] , 
        \round_in[1][511] , \round_in[1][510] , \round_in[1][509] , 
        \round_in[1][508] , \round_in[1][507] , \round_in[1][506] , 
        \round_in[1][505] , \round_in[1][504] , \round_in[1][503] , 
        \round_in[1][502] , \round_in[1][501] , \round_in[1][500] , 
        \round_in[1][499] , \round_in[1][498] , \round_in[1][497] , 
        \round_in[1][496] , \round_in[1][495] , \round_in[1][494] , 
        \round_in[1][493] , \round_in[1][492] , \round_in[1][491] , 
        \round_in[1][490] , \round_in[1][489] , \round_in[1][488] , 
        \round_in[1][487] , \round_in[1][486] , \round_in[1][485] , 
        \round_in[1][484] , \round_in[1][483] , \round_in[1][482] , 
        \round_in[1][481] , \round_in[1][480] , \round_in[1][479] , 
        \round_in[1][478] , \round_in[1][477] , \round_in[1][476] , 
        \round_in[1][475] , \round_in[1][474] , \round_in[1][473] , 
        \round_in[1][472] , \round_in[1][471] , \round_in[1][470] , 
        \round_in[1][469] , \round_in[1][468] , \round_in[1][467] , 
        \round_in[1][466] , \round_in[1][465] , \round_in[1][464] , 
        \round_in[1][463] , \round_in[1][462] , \round_in[1][461] , 
        \round_in[1][460] , \round_in[1][459] , \round_in[1][458] , 
        \round_in[1][457] , \round_in[1][456] , \round_in[1][455] , 
        \round_in[1][454] , \round_in[1][453] , \round_in[1][452] , 
        \round_in[1][451] , \round_in[1][450] , \round_in[1][449] , 
        \round_in[1][448] , \round_in[1][447] , \round_in[1][446] , 
        \round_in[1][445] , \round_in[1][444] , \round_in[1][443] , 
        \round_in[1][442] , \round_in[1][441] , \round_in[1][440] , 
        \round_in[1][439] , \round_in[1][438] , \round_in[1][437] , 
        \round_in[1][436] , \round_in[1][435] , \round_in[1][434] , 
        \round_in[1][433] , \round_in[1][432] , \round_in[1][431] , 
        \round_in[1][430] , \round_in[1][429] , \round_in[1][428] , 
        \round_in[1][427] , \round_in[1][426] , \round_in[1][425] , 
        \round_in[1][424] , \round_in[1][423] , \round_in[1][422] , 
        \round_in[1][421] , \round_in[1][420] , \round_in[1][419] , 
        \round_in[1][418] , \round_in[1][417] , \round_in[1][416] , 
        \round_in[1][415] , \round_in[1][414] , \round_in[1][413] , 
        \round_in[1][412] , \round_in[1][411] , \round_in[1][410] , 
        \round_in[1][409] , \round_in[1][408] , \round_in[1][407] , 
        \round_in[1][406] , \round_in[1][405] , \round_in[1][404] , 
        \round_in[1][403] , \round_in[1][402] , \round_in[1][401] , 
        \round_in[1][400] , \round_in[1][399] , \round_in[1][398] , 
        \round_in[1][397] , \round_in[1][396] , \round_in[1][395] , 
        \round_in[1][394] , \round_in[1][393] , \round_in[1][392] , 
        \round_in[1][391] , \round_in[1][390] , \round_in[1][389] , 
        \round_in[1][388] , \round_in[1][387] , \round_in[1][386] , 
        \round_in[1][385] , \round_in[1][384] , \round_in[1][383] , 
        \round_in[1][382] , \round_in[1][381] , \round_in[1][380] , 
        \round_in[1][379] , \round_in[1][378] , \round_in[1][377] , 
        \round_in[1][376] , \round_in[1][375] , \round_in[1][374] , 
        \round_in[1][373] , \round_in[1][372] , \round_in[1][371] , 
        \round_in[1][370] , \round_in[1][369] , \round_in[1][368] , 
        \round_in[1][367] , \round_in[1][366] , \round_in[1][365] , 
        \round_in[1][364] , \round_in[1][363] , \round_in[1][362] , 
        \round_in[1][361] , \round_in[1][360] , \round_in[1][359] , 
        \round_in[1][358] , \round_in[1][357] , \round_in[1][356] , 
        \round_in[1][355] , \round_in[1][354] , \round_in[1][353] , 
        \round_in[1][352] , \round_in[1][351] , \round_in[1][350] , 
        \round_in[1][349] , \round_in[1][348] , \round_in[1][347] , 
        \round_in[1][346] , \round_in[1][345] , \round_in[1][344] , 
        \round_in[1][343] , \round_in[1][342] , \round_in[1][341] , 
        \round_in[1][340] , \round_in[1][339] , \round_in[1][338] , 
        \round_in[1][337] , \round_in[1][336] , \round_in[1][335] , 
        \round_in[1][334] , \round_in[1][333] , \round_in[1][332] , 
        \round_in[1][331] , \round_in[1][330] , \round_in[1][329] , 
        \round_in[1][328] , \round_in[1][327] , \round_in[1][326] , 
        \round_in[1][325] , \round_in[1][324] , \round_in[1][323] , 
        \round_in[1][322] , \round_in[1][321] , \round_in[1][320] , 
        \round_in[1][319] , \round_in[1][318] , \round_in[1][317] , 
        \round_in[1][316] , \round_in[1][315] , \round_in[1][314] , 
        \round_in[1][313] , \round_in[1][312] , \round_in[1][311] , 
        \round_in[1][310] , \round_in[1][309] , \round_in[1][308] , 
        \round_in[1][307] , \round_in[1][306] , \round_in[1][305] , 
        \round_in[1][304] , \round_in[1][303] , \round_in[1][302] , 
        \round_in[1][301] , \round_in[1][300] , \round_in[1][299] , 
        \round_in[1][298] , \round_in[1][297] , \round_in[1][296] , 
        \round_in[1][295] , \round_in[1][294] , \round_in[1][293] , 
        \round_in[1][292] , \round_in[1][291] , \round_in[1][290] , 
        \round_in[1][289] , \round_in[1][288] , \round_in[1][287] , 
        \round_in[1][286] , \round_in[1][285] , \round_in[1][284] , 
        \round_in[1][283] , \round_in[1][282] , \round_in[1][281] , 
        \round_in[1][280] , \round_in[1][279] , \round_in[1][278] , 
        \round_in[1][277] , \round_in[1][276] , \round_in[1][275] , 
        \round_in[1][274] , \round_in[1][273] , \round_in[1][272] , 
        \round_in[1][271] , \round_in[1][270] , \round_in[1][269] , 
        \round_in[1][268] , \round_in[1][267] , \round_in[1][266] , 
        \round_in[1][265] , \round_in[1][264] , \round_in[1][263] , 
        \round_in[1][262] , \round_in[1][261] , \round_in[1][260] , 
        \round_in[1][259] , \round_in[1][258] , \round_in[1][257] , 
        \round_in[1][256] , \round_in[1][255] , \round_in[1][254] , 
        \round_in[1][253] , \round_in[1][252] , \round_in[1][251] , 
        \round_in[1][250] , \round_in[1][249] , \round_in[1][248] , 
        \round_in[1][247] , \round_in[1][246] , \round_in[1][245] , 
        \round_in[1][244] , \round_in[1][243] , \round_in[1][242] , 
        \round_in[1][241] , \round_in[1][240] , \round_in[1][239] , 
        \round_in[1][238] , \round_in[1][237] , \round_in[1][236] , 
        \round_in[1][235] , \round_in[1][234] , \round_in[1][233] , 
        \round_in[1][232] , \round_in[1][231] , \round_in[1][230] , 
        \round_in[1][229] , \round_in[1][228] , \round_in[1][227] , 
        \round_in[1][226] , \round_in[1][225] , \round_in[1][224] , 
        \round_in[1][223] , \round_in[1][222] , \round_in[1][221] , 
        \round_in[1][220] , \round_in[1][219] , \round_in[1][218] , 
        \round_in[1][217] , \round_in[1][216] , \round_in[1][215] , 
        \round_in[1][214] , \round_in[1][213] , \round_in[1][212] , 
        \round_in[1][211] , \round_in[1][210] , \round_in[1][209] , 
        \round_in[1][208] , \round_in[1][207] , \round_in[1][206] , 
        \round_in[1][205] , \round_in[1][204] , \round_in[1][203] , 
        \round_in[1][202] , \round_in[1][201] , \round_in[1][200] , 
        \round_in[1][199] , \round_in[1][198] , \round_in[1][197] , 
        \round_in[1][196] , \round_in[1][195] , \round_in[1][194] , 
        \round_in[1][193] , \round_in[1][192] , \round_in[1][191] , 
        \round_in[1][190] , \round_in[1][189] , \round_in[1][188] , 
        \round_in[1][187] , \round_in[1][186] , \round_in[1][185] , 
        \round_in[1][184] , \round_in[1][183] , \round_in[1][182] , 
        \round_in[1][181] , \round_in[1][180] , \round_in[1][179] , 
        \round_in[1][178] , \round_in[1][177] , \round_in[1][176] , 
        \round_in[1][175] , \round_in[1][174] , \round_in[1][173] , 
        \round_in[1][172] , \round_in[1][171] , \round_in[1][170] , 
        \round_in[1][169] , \round_in[1][168] , \round_in[1][167] , 
        \round_in[1][166] , \round_in[1][165] , \round_in[1][164] , 
        \round_in[1][163] , \round_in[1][162] , \round_in[1][161] , 
        \round_in[1][160] , \round_in[1][159] , \round_in[1][158] , 
        \round_in[1][157] , \round_in[1][156] , \round_in[1][155] , 
        \round_in[1][154] , \round_in[1][153] , \round_in[1][152] , 
        \round_in[1][151] , \round_in[1][150] , \round_in[1][149] , 
        \round_in[1][148] , \round_in[1][147] , \round_in[1][146] , 
        \round_in[1][145] , \round_in[1][144] , \round_in[1][143] , 
        \round_in[1][142] , \round_in[1][141] , \round_in[1][140] , 
        \round_in[1][139] , \round_in[1][138] , \round_in[1][137] , 
        \round_in[1][136] , \round_in[1][135] , \round_in[1][134] , 
        \round_in[1][133] , \round_in[1][132] , \round_in[1][131] , 
        \round_in[1][130] , \round_in[1][129] , \round_in[1][128] , 
        \round_in[1][127] , \round_in[1][126] , \round_in[1][125] , 
        \round_in[1][124] , \round_in[1][123] , \round_in[1][122] , 
        \round_in[1][121] , \round_in[1][120] , \round_in[1][119] , 
        \round_in[1][118] , \round_in[1][117] , \round_in[1][116] , 
        \round_in[1][115] , \round_in[1][114] , \round_in[1][113] , 
        \round_in[1][112] , \round_in[1][111] , \round_in[1][110] , 
        \round_in[1][109] , \round_in[1][108] , \round_in[1][107] , 
        \round_in[1][106] , \round_in[1][105] , \round_in[1][104] , 
        \round_in[1][103] , \round_in[1][102] , \round_in[1][101] , 
        \round_in[1][100] , \round_in[1][99] , \round_in[1][98] , 
        \round_in[1][97] , \round_in[1][96] , \round_in[1][95] , 
        \round_in[1][94] , \round_in[1][93] , \round_in[1][92] , 
        \round_in[1][91] , \round_in[1][90] , \round_in[1][89] , 
        \round_in[1][88] , \round_in[1][87] , \round_in[1][86] , 
        \round_in[1][85] , \round_in[1][84] , \round_in[1][83] , 
        \round_in[1][82] , \round_in[1][81] , \round_in[1][80] , 
        \round_in[1][79] , \round_in[1][78] , \round_in[1][77] , 
        \round_in[1][76] , \round_in[1][75] , \round_in[1][74] , 
        \round_in[1][73] , \round_in[1][72] , \round_in[1][71] , 
        \round_in[1][70] , \round_in[1][69] , \round_in[1][68] , 
        \round_in[1][67] , \round_in[1][66] , \round_in[1][65] , 
        \round_in[1][64] , \round_in[1][63] , \round_in[1][62] , 
        \round_in[1][61] , \round_in[1][60] , \round_in[1][59] , 
        \round_in[1][58] , \round_in[1][57] , \round_in[1][56] , 
        \round_in[1][55] , \round_in[1][54] , \round_in[1][53] , 
        \round_in[1][52] , \round_in[1][51] , \round_in[1][50] , 
        \round_in[1][49] , \round_in[1][48] , \round_in[1][47] , 
        \round_in[1][46] , \round_in[1][45] , \round_in[1][44] , 
        \round_in[1][43] , \round_in[1][42] , \round_in[1][41] , 
        \round_in[1][40] , \round_in[1][39] , \round_in[1][38] , 
        \round_in[1][37] , \round_in[1][36] , \round_in[1][35] , 
        \round_in[1][34] , \round_in[1][33] , \round_in[1][32] , 
        \round_in[1][31] , \round_in[1][30] , \round_in[1][29] , 
        \round_in[1][28] , \round_in[1][27] , \round_in[1][26] , 
        \round_in[1][25] , \round_in[1][24] , \round_in[1][23] , 
        \round_in[1][22] , \round_in[1][21] , \round_in[1][20] , 
        \round_in[1][19] , \round_in[1][18] , \round_in[1][17] , 
        \round_in[1][16] , \round_in[1][15] , \round_in[1][14] , 
        \round_in[1][13] , \round_in[1][12] , \round_in[1][11] , 
        \round_in[1][10] , \round_in[1][9] , \round_in[1][8] , 
        \round_in[1][7] , \round_in[1][6] , \round_in[1][5] , \round_in[1][4] , 
        \round_in[1][3] , \round_in[1][2] , \round_in[1][1] , \round_in[1][0] }), .round_const({\rc[1][63] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \rc[1][31] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \rc[1][15] , 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, \rc[1][7] , 1'b0, 1'b0, 1'b0, \rc[1][3] , 1'b0, 
        \rc[1][1] , \RCONST[1].rconst_/N10 }), .out(out) );
  DFF init_reg ( .D(n2792), .CLK(clk), .RST(1'b0), .Q(init) );
  DFF \rc_i_reg[0]  ( .D(N6), .CLK(clk), .RST(1'b0), .Q(rc_i[0]) );
  DFF \rc_i_reg[1]  ( .D(N7), .CLK(clk), .RST(1'b0), .Q(rc_i[1]) );
  DFF \rc_i_reg[2]  ( .D(N8), .CLK(clk), .RST(1'b0), .Q(rc_i[2]) );
  DFF \rc_i_reg[3]  ( .D(N9), .CLK(clk), .RST(1'b0), .Q(rc_i[3]) );
  DFF \rc_i_reg[4]  ( .D(N10), .CLK(clk), .RST(1'b0), .Q(rc_i[4]) );
  DFF \rc_i_reg[5]  ( .D(N11), .CLK(clk), .RST(1'b0), .Q(rc_i[5]) );
  DFF \rc_i_reg[6]  ( .D(N12), .CLK(clk), .RST(1'b0), .Q(rc_i[6]) );
  DFF \rc_i_reg[7]  ( .D(N13), .CLK(clk), .RST(1'b0), .Q(rc_i[7]) );
  DFF \rc_i_reg[8]  ( .D(N14), .CLK(clk), .RST(1'b0), .Q(rc_i[8]) );
  DFF \rc_i_reg[9]  ( .D(N15), .CLK(clk), .RST(1'b0), .Q(rc_i[9]) );
  DFF \rc_i_reg[10]  ( .D(N16), .CLK(clk), .RST(1'b0), .Q(rc_i[10]) );
  DFF \rc_i_reg[11]  ( .D(N17), .CLK(clk), .RST(1'b0), .Q(rc_i[11]) );
  DFF \round_reg_reg[0]  ( .D(N18), .CLK(clk), .RST(1'b0), .Q(round_reg[0]) );
  DFF \round_reg_reg[1]  ( .D(N19), .CLK(clk), .RST(1'b0), .Q(round_reg[1]) );
  DFF \round_reg_reg[2]  ( .D(N20), .CLK(clk), .RST(1'b0), .Q(round_reg[2]) );
  DFF \round_reg_reg[3]  ( .D(N21), .CLK(clk), .RST(1'b0), .Q(round_reg[3]) );
  DFF \round_reg_reg[4]  ( .D(N22), .CLK(clk), .RST(1'b0), .Q(round_reg[4]) );
  DFF \round_reg_reg[5]  ( .D(N23), .CLK(clk), .RST(1'b0), .Q(round_reg[5]) );
  DFF \round_reg_reg[6]  ( .D(N24), .CLK(clk), .RST(1'b0), .Q(round_reg[6]) );
  DFF \round_reg_reg[7]  ( .D(N25), .CLK(clk), .RST(1'b0), .Q(round_reg[7]) );
  DFF \round_reg_reg[8]  ( .D(N26), .CLK(clk), .RST(1'b0), .Q(round_reg[8]) );
  DFF \round_reg_reg[9]  ( .D(N27), .CLK(clk), .RST(1'b0), .Q(round_reg[9]) );
  DFF \round_reg_reg[10]  ( .D(N28), .CLK(clk), .RST(1'b0), .Q(round_reg[10])
         );
  DFF \round_reg_reg[11]  ( .D(N29), .CLK(clk), .RST(1'b0), .Q(round_reg[11])
         );
  DFF \round_reg_reg[12]  ( .D(N30), .CLK(clk), .RST(1'b0), .Q(round_reg[12])
         );
  DFF \round_reg_reg[13]  ( .D(N31), .CLK(clk), .RST(1'b0), .Q(round_reg[13])
         );
  DFF \round_reg_reg[14]  ( .D(N32), .CLK(clk), .RST(1'b0), .Q(round_reg[14])
         );
  DFF \round_reg_reg[15]  ( .D(N33), .CLK(clk), .RST(1'b0), .Q(round_reg[15])
         );
  DFF \round_reg_reg[16]  ( .D(N34), .CLK(clk), .RST(1'b0), .Q(round_reg[16])
         );
  DFF \round_reg_reg[17]  ( .D(N35), .CLK(clk), .RST(1'b0), .Q(round_reg[17])
         );
  DFF \round_reg_reg[18]  ( .D(N36), .CLK(clk), .RST(1'b0), .Q(round_reg[18])
         );
  DFF \round_reg_reg[19]  ( .D(N37), .CLK(clk), .RST(1'b0), .Q(round_reg[19])
         );
  DFF \round_reg_reg[20]  ( .D(N38), .CLK(clk), .RST(1'b0), .Q(round_reg[20])
         );
  DFF \round_reg_reg[21]  ( .D(N39), .CLK(clk), .RST(1'b0), .Q(round_reg[21])
         );
  DFF \round_reg_reg[22]  ( .D(N40), .CLK(clk), .RST(1'b0), .Q(round_reg[22])
         );
  DFF \round_reg_reg[23]  ( .D(N41), .CLK(clk), .RST(1'b0), .Q(round_reg[23])
         );
  DFF \round_reg_reg[24]  ( .D(N42), .CLK(clk), .RST(1'b0), .Q(round_reg[24])
         );
  DFF \round_reg_reg[25]  ( .D(N43), .CLK(clk), .RST(1'b0), .Q(round_reg[25])
         );
  DFF \round_reg_reg[26]  ( .D(N44), .CLK(clk), .RST(1'b0), .Q(round_reg[26])
         );
  DFF \round_reg_reg[27]  ( .D(N45), .CLK(clk), .RST(1'b0), .Q(round_reg[27])
         );
  DFF \round_reg_reg[28]  ( .D(N46), .CLK(clk), .RST(1'b0), .Q(round_reg[28])
         );
  DFF \round_reg_reg[29]  ( .D(N47), .CLK(clk), .RST(1'b0), .Q(round_reg[29])
         );
  DFF \round_reg_reg[30]  ( .D(N48), .CLK(clk), .RST(1'b0), .Q(round_reg[30])
         );
  DFF \round_reg_reg[31]  ( .D(N49), .CLK(clk), .RST(1'b0), .Q(round_reg[31])
         );
  DFF \round_reg_reg[32]  ( .D(N50), .CLK(clk), .RST(1'b0), .Q(round_reg[32])
         );
  DFF \round_reg_reg[33]  ( .D(N51), .CLK(clk), .RST(1'b0), .Q(round_reg[33])
         );
  DFF \round_reg_reg[34]  ( .D(N52), .CLK(clk), .RST(1'b0), .Q(round_reg[34])
         );
  DFF \round_reg_reg[35]  ( .D(N53), .CLK(clk), .RST(1'b0), .Q(round_reg[35])
         );
  DFF \round_reg_reg[36]  ( .D(N54), .CLK(clk), .RST(1'b0), .Q(round_reg[36])
         );
  DFF \round_reg_reg[37]  ( .D(N55), .CLK(clk), .RST(1'b0), .Q(round_reg[37])
         );
  DFF \round_reg_reg[38]  ( .D(N56), .CLK(clk), .RST(1'b0), .Q(round_reg[38])
         );
  DFF \round_reg_reg[39]  ( .D(N57), .CLK(clk), .RST(1'b0), .Q(round_reg[39])
         );
  DFF \round_reg_reg[40]  ( .D(N58), .CLK(clk), .RST(1'b0), .Q(round_reg[40])
         );
  DFF \round_reg_reg[41]  ( .D(N59), .CLK(clk), .RST(1'b0), .Q(round_reg[41])
         );
  DFF \round_reg_reg[42]  ( .D(N60), .CLK(clk), .RST(1'b0), .Q(round_reg[42])
         );
  DFF \round_reg_reg[43]  ( .D(N61), .CLK(clk), .RST(1'b0), .Q(round_reg[43])
         );
  DFF \round_reg_reg[44]  ( .D(N62), .CLK(clk), .RST(1'b0), .Q(round_reg[44])
         );
  DFF \round_reg_reg[45]  ( .D(N63), .CLK(clk), .RST(1'b0), .Q(round_reg[45])
         );
  DFF \round_reg_reg[46]  ( .D(N64), .CLK(clk), .RST(1'b0), .Q(round_reg[46])
         );
  DFF \round_reg_reg[47]  ( .D(N65), .CLK(clk), .RST(1'b0), .Q(round_reg[47])
         );
  DFF \round_reg_reg[48]  ( .D(N66), .CLK(clk), .RST(1'b0), .Q(round_reg[48])
         );
  DFF \round_reg_reg[49]  ( .D(N67), .CLK(clk), .RST(1'b0), .Q(round_reg[49])
         );
  DFF \round_reg_reg[50]  ( .D(N68), .CLK(clk), .RST(1'b0), .Q(round_reg[50])
         );
  DFF \round_reg_reg[51]  ( .D(N69), .CLK(clk), .RST(1'b0), .Q(round_reg[51])
         );
  DFF \round_reg_reg[52]  ( .D(N70), .CLK(clk), .RST(1'b0), .Q(round_reg[52])
         );
  DFF \round_reg_reg[53]  ( .D(N71), .CLK(clk), .RST(1'b0), .Q(round_reg[53])
         );
  DFF \round_reg_reg[54]  ( .D(N72), .CLK(clk), .RST(1'b0), .Q(round_reg[54])
         );
  DFF \round_reg_reg[55]  ( .D(N73), .CLK(clk), .RST(1'b0), .Q(round_reg[55])
         );
  DFF \round_reg_reg[56]  ( .D(N74), .CLK(clk), .RST(1'b0), .Q(round_reg[56])
         );
  DFF \round_reg_reg[57]  ( .D(N75), .CLK(clk), .RST(1'b0), .Q(round_reg[57])
         );
  DFF \round_reg_reg[58]  ( .D(N76), .CLK(clk), .RST(1'b0), .Q(round_reg[58])
         );
  DFF \round_reg_reg[59]  ( .D(N77), .CLK(clk), .RST(1'b0), .Q(round_reg[59])
         );
  DFF \round_reg_reg[60]  ( .D(N78), .CLK(clk), .RST(1'b0), .Q(round_reg[60])
         );
  DFF \round_reg_reg[61]  ( .D(N79), .CLK(clk), .RST(1'b0), .Q(round_reg[61])
         );
  DFF \round_reg_reg[62]  ( .D(N80), .CLK(clk), .RST(1'b0), .Q(round_reg[62])
         );
  DFF \round_reg_reg[63]  ( .D(N81), .CLK(clk), .RST(1'b0), .Q(round_reg[63])
         );
  DFF \round_reg_reg[64]  ( .D(N82), .CLK(clk), .RST(1'b0), .Q(round_reg[64])
         );
  DFF \round_reg_reg[65]  ( .D(N83), .CLK(clk), .RST(1'b0), .Q(round_reg[65])
         );
  DFF \round_reg_reg[66]  ( .D(N84), .CLK(clk), .RST(1'b0), .Q(round_reg[66])
         );
  DFF \round_reg_reg[67]  ( .D(N85), .CLK(clk), .RST(1'b0), .Q(round_reg[67])
         );
  DFF \round_reg_reg[68]  ( .D(N86), .CLK(clk), .RST(1'b0), .Q(round_reg[68])
         );
  DFF \round_reg_reg[69]  ( .D(N87), .CLK(clk), .RST(1'b0), .Q(round_reg[69])
         );
  DFF \round_reg_reg[70]  ( .D(N88), .CLK(clk), .RST(1'b0), .Q(round_reg[70])
         );
  DFF \round_reg_reg[71]  ( .D(N89), .CLK(clk), .RST(1'b0), .Q(round_reg[71])
         );
  DFF \round_reg_reg[72]  ( .D(N90), .CLK(clk), .RST(1'b0), .Q(round_reg[72])
         );
  DFF \round_reg_reg[73]  ( .D(N91), .CLK(clk), .RST(1'b0), .Q(round_reg[73])
         );
  DFF \round_reg_reg[74]  ( .D(N92), .CLK(clk), .RST(1'b0), .Q(round_reg[74])
         );
  DFF \round_reg_reg[75]  ( .D(N93), .CLK(clk), .RST(1'b0), .Q(round_reg[75])
         );
  DFF \round_reg_reg[76]  ( .D(N94), .CLK(clk), .RST(1'b0), .Q(round_reg[76])
         );
  DFF \round_reg_reg[77]  ( .D(N95), .CLK(clk), .RST(1'b0), .Q(round_reg[77])
         );
  DFF \round_reg_reg[78]  ( .D(N96), .CLK(clk), .RST(1'b0), .Q(round_reg[78])
         );
  DFF \round_reg_reg[79]  ( .D(N97), .CLK(clk), .RST(1'b0), .Q(round_reg[79])
         );
  DFF \round_reg_reg[80]  ( .D(N98), .CLK(clk), .RST(1'b0), .Q(round_reg[80])
         );
  DFF \round_reg_reg[81]  ( .D(N99), .CLK(clk), .RST(1'b0), .Q(round_reg[81])
         );
  DFF \round_reg_reg[82]  ( .D(N100), .CLK(clk), .RST(1'b0), .Q(round_reg[82])
         );
  DFF \round_reg_reg[83]  ( .D(N101), .CLK(clk), .RST(1'b0), .Q(round_reg[83])
         );
  DFF \round_reg_reg[84]  ( .D(N102), .CLK(clk), .RST(1'b0), .Q(round_reg[84])
         );
  DFF \round_reg_reg[85]  ( .D(N103), .CLK(clk), .RST(1'b0), .Q(round_reg[85])
         );
  DFF \round_reg_reg[86]  ( .D(N104), .CLK(clk), .RST(1'b0), .Q(round_reg[86])
         );
  DFF \round_reg_reg[87]  ( .D(N105), .CLK(clk), .RST(1'b0), .Q(round_reg[87])
         );
  DFF \round_reg_reg[88]  ( .D(N106), .CLK(clk), .RST(1'b0), .Q(round_reg[88])
         );
  DFF \round_reg_reg[89]  ( .D(N107), .CLK(clk), .RST(1'b0), .Q(round_reg[89])
         );
  DFF \round_reg_reg[90]  ( .D(N108), .CLK(clk), .RST(1'b0), .Q(round_reg[90])
         );
  DFF \round_reg_reg[91]  ( .D(N109), .CLK(clk), .RST(1'b0), .Q(round_reg[91])
         );
  DFF \round_reg_reg[92]  ( .D(N110), .CLK(clk), .RST(1'b0), .Q(round_reg[92])
         );
  DFF \round_reg_reg[93]  ( .D(N111), .CLK(clk), .RST(1'b0), .Q(round_reg[93])
         );
  DFF \round_reg_reg[94]  ( .D(N112), .CLK(clk), .RST(1'b0), .Q(round_reg[94])
         );
  DFF \round_reg_reg[95]  ( .D(N113), .CLK(clk), .RST(1'b0), .Q(round_reg[95])
         );
  DFF \round_reg_reg[96]  ( .D(N114), .CLK(clk), .RST(1'b0), .Q(round_reg[96])
         );
  DFF \round_reg_reg[97]  ( .D(N115), .CLK(clk), .RST(1'b0), .Q(round_reg[97])
         );
  DFF \round_reg_reg[98]  ( .D(N116), .CLK(clk), .RST(1'b0), .Q(round_reg[98])
         );
  DFF \round_reg_reg[99]  ( .D(N117), .CLK(clk), .RST(1'b0), .Q(round_reg[99])
         );
  DFF \round_reg_reg[100]  ( .D(N118), .CLK(clk), .RST(1'b0), .Q(
        round_reg[100]) );
  DFF \round_reg_reg[101]  ( .D(N119), .CLK(clk), .RST(1'b0), .Q(
        round_reg[101]) );
  DFF \round_reg_reg[102]  ( .D(N120), .CLK(clk), .RST(1'b0), .Q(
        round_reg[102]) );
  DFF \round_reg_reg[103]  ( .D(N121), .CLK(clk), .RST(1'b0), .Q(
        round_reg[103]) );
  DFF \round_reg_reg[104]  ( .D(N122), .CLK(clk), .RST(1'b0), .Q(
        round_reg[104]) );
  DFF \round_reg_reg[105]  ( .D(N123), .CLK(clk), .RST(1'b0), .Q(
        round_reg[105]) );
  DFF \round_reg_reg[106]  ( .D(N124), .CLK(clk), .RST(1'b0), .Q(
        round_reg[106]) );
  DFF \round_reg_reg[107]  ( .D(N125), .CLK(clk), .RST(1'b0), .Q(
        round_reg[107]) );
  DFF \round_reg_reg[108]  ( .D(N126), .CLK(clk), .RST(1'b0), .Q(
        round_reg[108]) );
  DFF \round_reg_reg[109]  ( .D(N127), .CLK(clk), .RST(1'b0), .Q(
        round_reg[109]) );
  DFF \round_reg_reg[110]  ( .D(N128), .CLK(clk), .RST(1'b0), .Q(
        round_reg[110]) );
  DFF \round_reg_reg[111]  ( .D(N129), .CLK(clk), .RST(1'b0), .Q(
        round_reg[111]) );
  DFF \round_reg_reg[112]  ( .D(N130), .CLK(clk), .RST(1'b0), .Q(
        round_reg[112]) );
  DFF \round_reg_reg[113]  ( .D(N131), .CLK(clk), .RST(1'b0), .Q(
        round_reg[113]) );
  DFF \round_reg_reg[114]  ( .D(N132), .CLK(clk), .RST(1'b0), .Q(
        round_reg[114]) );
  DFF \round_reg_reg[115]  ( .D(N133), .CLK(clk), .RST(1'b0), .Q(
        round_reg[115]) );
  DFF \round_reg_reg[116]  ( .D(N134), .CLK(clk), .RST(1'b0), .Q(
        round_reg[116]) );
  DFF \round_reg_reg[117]  ( .D(N135), .CLK(clk), .RST(1'b0), .Q(
        round_reg[117]) );
  DFF \round_reg_reg[118]  ( .D(N136), .CLK(clk), .RST(1'b0), .Q(
        round_reg[118]) );
  DFF \round_reg_reg[119]  ( .D(N137), .CLK(clk), .RST(1'b0), .Q(
        round_reg[119]) );
  DFF \round_reg_reg[120]  ( .D(N138), .CLK(clk), .RST(1'b0), .Q(
        round_reg[120]) );
  DFF \round_reg_reg[121]  ( .D(N139), .CLK(clk), .RST(1'b0), .Q(
        round_reg[121]) );
  DFF \round_reg_reg[122]  ( .D(N140), .CLK(clk), .RST(1'b0), .Q(
        round_reg[122]) );
  DFF \round_reg_reg[123]  ( .D(N141), .CLK(clk), .RST(1'b0), .Q(
        round_reg[123]) );
  DFF \round_reg_reg[124]  ( .D(N142), .CLK(clk), .RST(1'b0), .Q(
        round_reg[124]) );
  DFF \round_reg_reg[125]  ( .D(N143), .CLK(clk), .RST(1'b0), .Q(
        round_reg[125]) );
  DFF \round_reg_reg[126]  ( .D(N144), .CLK(clk), .RST(1'b0), .Q(
        round_reg[126]) );
  DFF \round_reg_reg[127]  ( .D(N145), .CLK(clk), .RST(1'b0), .Q(
        round_reg[127]) );
  DFF \round_reg_reg[128]  ( .D(N146), .CLK(clk), .RST(1'b0), .Q(
        round_reg[128]) );
  DFF \round_reg_reg[129]  ( .D(N147), .CLK(clk), .RST(1'b0), .Q(
        round_reg[129]) );
  DFF \round_reg_reg[130]  ( .D(N148), .CLK(clk), .RST(1'b0), .Q(
        round_reg[130]) );
  DFF \round_reg_reg[131]  ( .D(N149), .CLK(clk), .RST(1'b0), .Q(
        round_reg[131]) );
  DFF \round_reg_reg[132]  ( .D(N150), .CLK(clk), .RST(1'b0), .Q(
        round_reg[132]) );
  DFF \round_reg_reg[133]  ( .D(N151), .CLK(clk), .RST(1'b0), .Q(
        round_reg[133]) );
  DFF \round_reg_reg[134]  ( .D(N152), .CLK(clk), .RST(1'b0), .Q(
        round_reg[134]) );
  DFF \round_reg_reg[135]  ( .D(N153), .CLK(clk), .RST(1'b0), .Q(
        round_reg[135]) );
  DFF \round_reg_reg[136]  ( .D(N154), .CLK(clk), .RST(1'b0), .Q(
        round_reg[136]) );
  DFF \round_reg_reg[137]  ( .D(N155), .CLK(clk), .RST(1'b0), .Q(
        round_reg[137]) );
  DFF \round_reg_reg[138]  ( .D(N156), .CLK(clk), .RST(1'b0), .Q(
        round_reg[138]) );
  DFF \round_reg_reg[139]  ( .D(N157), .CLK(clk), .RST(1'b0), .Q(
        round_reg[139]) );
  DFF \round_reg_reg[140]  ( .D(N158), .CLK(clk), .RST(1'b0), .Q(
        round_reg[140]) );
  DFF \round_reg_reg[141]  ( .D(N159), .CLK(clk), .RST(1'b0), .Q(
        round_reg[141]) );
  DFF \round_reg_reg[142]  ( .D(N160), .CLK(clk), .RST(1'b0), .Q(
        round_reg[142]) );
  DFF \round_reg_reg[143]  ( .D(N161), .CLK(clk), .RST(1'b0), .Q(
        round_reg[143]) );
  DFF \round_reg_reg[144]  ( .D(N162), .CLK(clk), .RST(1'b0), .Q(
        round_reg[144]) );
  DFF \round_reg_reg[145]  ( .D(N163), .CLK(clk), .RST(1'b0), .Q(
        round_reg[145]) );
  DFF \round_reg_reg[146]  ( .D(N164), .CLK(clk), .RST(1'b0), .Q(
        round_reg[146]) );
  DFF \round_reg_reg[147]  ( .D(N165), .CLK(clk), .RST(1'b0), .Q(
        round_reg[147]) );
  DFF \round_reg_reg[148]  ( .D(N166), .CLK(clk), .RST(1'b0), .Q(
        round_reg[148]) );
  DFF \round_reg_reg[149]  ( .D(N167), .CLK(clk), .RST(1'b0), .Q(
        round_reg[149]) );
  DFF \round_reg_reg[150]  ( .D(N168), .CLK(clk), .RST(1'b0), .Q(
        round_reg[150]) );
  DFF \round_reg_reg[151]  ( .D(N169), .CLK(clk), .RST(1'b0), .Q(
        round_reg[151]) );
  DFF \round_reg_reg[152]  ( .D(N170), .CLK(clk), .RST(1'b0), .Q(
        round_reg[152]) );
  DFF \round_reg_reg[153]  ( .D(N171), .CLK(clk), .RST(1'b0), .Q(
        round_reg[153]) );
  DFF \round_reg_reg[154]  ( .D(N172), .CLK(clk), .RST(1'b0), .Q(
        round_reg[154]) );
  DFF \round_reg_reg[155]  ( .D(N173), .CLK(clk), .RST(1'b0), .Q(
        round_reg[155]) );
  DFF \round_reg_reg[156]  ( .D(N174), .CLK(clk), .RST(1'b0), .Q(
        round_reg[156]) );
  DFF \round_reg_reg[157]  ( .D(N175), .CLK(clk), .RST(1'b0), .Q(
        round_reg[157]) );
  DFF \round_reg_reg[158]  ( .D(N176), .CLK(clk), .RST(1'b0), .Q(
        round_reg[158]) );
  DFF \round_reg_reg[159]  ( .D(N177), .CLK(clk), .RST(1'b0), .Q(
        round_reg[159]) );
  DFF \round_reg_reg[160]  ( .D(N178), .CLK(clk), .RST(1'b0), .Q(
        round_reg[160]) );
  DFF \round_reg_reg[161]  ( .D(N179), .CLK(clk), .RST(1'b0), .Q(
        round_reg[161]) );
  DFF \round_reg_reg[162]  ( .D(N180), .CLK(clk), .RST(1'b0), .Q(
        round_reg[162]) );
  DFF \round_reg_reg[163]  ( .D(N181), .CLK(clk), .RST(1'b0), .Q(
        round_reg[163]) );
  DFF \round_reg_reg[164]  ( .D(N182), .CLK(clk), .RST(1'b0), .Q(
        round_reg[164]) );
  DFF \round_reg_reg[165]  ( .D(N183), .CLK(clk), .RST(1'b0), .Q(
        round_reg[165]) );
  DFF \round_reg_reg[166]  ( .D(N184), .CLK(clk), .RST(1'b0), .Q(
        round_reg[166]) );
  DFF \round_reg_reg[167]  ( .D(N185), .CLK(clk), .RST(1'b0), .Q(
        round_reg[167]) );
  DFF \round_reg_reg[168]  ( .D(N186), .CLK(clk), .RST(1'b0), .Q(
        round_reg[168]) );
  DFF \round_reg_reg[169]  ( .D(N187), .CLK(clk), .RST(1'b0), .Q(
        round_reg[169]) );
  DFF \round_reg_reg[170]  ( .D(N188), .CLK(clk), .RST(1'b0), .Q(
        round_reg[170]) );
  DFF \round_reg_reg[171]  ( .D(N189), .CLK(clk), .RST(1'b0), .Q(
        round_reg[171]) );
  DFF \round_reg_reg[172]  ( .D(N190), .CLK(clk), .RST(1'b0), .Q(
        round_reg[172]) );
  DFF \round_reg_reg[173]  ( .D(N191), .CLK(clk), .RST(1'b0), .Q(
        round_reg[173]) );
  DFF \round_reg_reg[174]  ( .D(N192), .CLK(clk), .RST(1'b0), .Q(
        round_reg[174]) );
  DFF \round_reg_reg[175]  ( .D(N193), .CLK(clk), .RST(1'b0), .Q(
        round_reg[175]) );
  DFF \round_reg_reg[176]  ( .D(N194), .CLK(clk), .RST(1'b0), .Q(
        round_reg[176]) );
  DFF \round_reg_reg[177]  ( .D(N195), .CLK(clk), .RST(1'b0), .Q(
        round_reg[177]) );
  DFF \round_reg_reg[178]  ( .D(N196), .CLK(clk), .RST(1'b0), .Q(
        round_reg[178]) );
  DFF \round_reg_reg[179]  ( .D(N197), .CLK(clk), .RST(1'b0), .Q(
        round_reg[179]) );
  DFF \round_reg_reg[180]  ( .D(N198), .CLK(clk), .RST(1'b0), .Q(
        round_reg[180]) );
  DFF \round_reg_reg[181]  ( .D(N199), .CLK(clk), .RST(1'b0), .Q(
        round_reg[181]) );
  DFF \round_reg_reg[182]  ( .D(N200), .CLK(clk), .RST(1'b0), .Q(
        round_reg[182]) );
  DFF \round_reg_reg[183]  ( .D(N201), .CLK(clk), .RST(1'b0), .Q(
        round_reg[183]) );
  DFF \round_reg_reg[184]  ( .D(N202), .CLK(clk), .RST(1'b0), .Q(
        round_reg[184]) );
  DFF \round_reg_reg[185]  ( .D(N203), .CLK(clk), .RST(1'b0), .Q(
        round_reg[185]) );
  DFF \round_reg_reg[186]  ( .D(N204), .CLK(clk), .RST(1'b0), .Q(
        round_reg[186]) );
  DFF \round_reg_reg[187]  ( .D(N205), .CLK(clk), .RST(1'b0), .Q(
        round_reg[187]) );
  DFF \round_reg_reg[188]  ( .D(N206), .CLK(clk), .RST(1'b0), .Q(
        round_reg[188]) );
  DFF \round_reg_reg[189]  ( .D(N207), .CLK(clk), .RST(1'b0), .Q(
        round_reg[189]) );
  DFF \round_reg_reg[190]  ( .D(N208), .CLK(clk), .RST(1'b0), .Q(
        round_reg[190]) );
  DFF \round_reg_reg[191]  ( .D(N209), .CLK(clk), .RST(1'b0), .Q(
        round_reg[191]) );
  DFF \round_reg_reg[192]  ( .D(N210), .CLK(clk), .RST(1'b0), .Q(
        round_reg[192]) );
  DFF \round_reg_reg[193]  ( .D(N211), .CLK(clk), .RST(1'b0), .Q(
        round_reg[193]) );
  DFF \round_reg_reg[194]  ( .D(N212), .CLK(clk), .RST(1'b0), .Q(
        round_reg[194]) );
  DFF \round_reg_reg[195]  ( .D(N213), .CLK(clk), .RST(1'b0), .Q(
        round_reg[195]) );
  DFF \round_reg_reg[196]  ( .D(N214), .CLK(clk), .RST(1'b0), .Q(
        round_reg[196]) );
  DFF \round_reg_reg[197]  ( .D(N215), .CLK(clk), .RST(1'b0), .Q(
        round_reg[197]) );
  DFF \round_reg_reg[198]  ( .D(N216), .CLK(clk), .RST(1'b0), .Q(
        round_reg[198]) );
  DFF \round_reg_reg[199]  ( .D(N217), .CLK(clk), .RST(1'b0), .Q(
        round_reg[199]) );
  DFF \round_reg_reg[200]  ( .D(N218), .CLK(clk), .RST(1'b0), .Q(
        round_reg[200]) );
  DFF \round_reg_reg[201]  ( .D(N219), .CLK(clk), .RST(1'b0), .Q(
        round_reg[201]) );
  DFF \round_reg_reg[202]  ( .D(N220), .CLK(clk), .RST(1'b0), .Q(
        round_reg[202]) );
  DFF \round_reg_reg[203]  ( .D(N221), .CLK(clk), .RST(1'b0), .Q(
        round_reg[203]) );
  DFF \round_reg_reg[204]  ( .D(N222), .CLK(clk), .RST(1'b0), .Q(
        round_reg[204]) );
  DFF \round_reg_reg[205]  ( .D(N223), .CLK(clk), .RST(1'b0), .Q(
        round_reg[205]) );
  DFF \round_reg_reg[206]  ( .D(N224), .CLK(clk), .RST(1'b0), .Q(
        round_reg[206]) );
  DFF \round_reg_reg[207]  ( .D(N225), .CLK(clk), .RST(1'b0), .Q(
        round_reg[207]) );
  DFF \round_reg_reg[208]  ( .D(N226), .CLK(clk), .RST(1'b0), .Q(
        round_reg[208]) );
  DFF \round_reg_reg[209]  ( .D(N227), .CLK(clk), .RST(1'b0), .Q(
        round_reg[209]) );
  DFF \round_reg_reg[210]  ( .D(N228), .CLK(clk), .RST(1'b0), .Q(
        round_reg[210]) );
  DFF \round_reg_reg[211]  ( .D(N229), .CLK(clk), .RST(1'b0), .Q(
        round_reg[211]) );
  DFF \round_reg_reg[212]  ( .D(N230), .CLK(clk), .RST(1'b0), .Q(
        round_reg[212]) );
  DFF \round_reg_reg[213]  ( .D(N231), .CLK(clk), .RST(1'b0), .Q(
        round_reg[213]) );
  DFF \round_reg_reg[214]  ( .D(N232), .CLK(clk), .RST(1'b0), .Q(
        round_reg[214]) );
  DFF \round_reg_reg[215]  ( .D(N233), .CLK(clk), .RST(1'b0), .Q(
        round_reg[215]) );
  DFF \round_reg_reg[216]  ( .D(N234), .CLK(clk), .RST(1'b0), .Q(
        round_reg[216]) );
  DFF \round_reg_reg[217]  ( .D(N235), .CLK(clk), .RST(1'b0), .Q(
        round_reg[217]) );
  DFF \round_reg_reg[218]  ( .D(N236), .CLK(clk), .RST(1'b0), .Q(
        round_reg[218]) );
  DFF \round_reg_reg[219]  ( .D(N237), .CLK(clk), .RST(1'b0), .Q(
        round_reg[219]) );
  DFF \round_reg_reg[220]  ( .D(N238), .CLK(clk), .RST(1'b0), .Q(
        round_reg[220]) );
  DFF \round_reg_reg[221]  ( .D(N239), .CLK(clk), .RST(1'b0), .Q(
        round_reg[221]) );
  DFF \round_reg_reg[222]  ( .D(N240), .CLK(clk), .RST(1'b0), .Q(
        round_reg[222]) );
  DFF \round_reg_reg[223]  ( .D(N241), .CLK(clk), .RST(1'b0), .Q(
        round_reg[223]) );
  DFF \round_reg_reg[224]  ( .D(N242), .CLK(clk), .RST(1'b0), .Q(
        round_reg[224]) );
  DFF \round_reg_reg[225]  ( .D(N243), .CLK(clk), .RST(1'b0), .Q(
        round_reg[225]) );
  DFF \round_reg_reg[226]  ( .D(N244), .CLK(clk), .RST(1'b0), .Q(
        round_reg[226]) );
  DFF \round_reg_reg[227]  ( .D(N245), .CLK(clk), .RST(1'b0), .Q(
        round_reg[227]) );
  DFF \round_reg_reg[228]  ( .D(N246), .CLK(clk), .RST(1'b0), .Q(
        round_reg[228]) );
  DFF \round_reg_reg[229]  ( .D(N247), .CLK(clk), .RST(1'b0), .Q(
        round_reg[229]) );
  DFF \round_reg_reg[230]  ( .D(N248), .CLK(clk), .RST(1'b0), .Q(
        round_reg[230]) );
  DFF \round_reg_reg[231]  ( .D(N249), .CLK(clk), .RST(1'b0), .Q(
        round_reg[231]) );
  DFF \round_reg_reg[232]  ( .D(N250), .CLK(clk), .RST(1'b0), .Q(
        round_reg[232]) );
  DFF \round_reg_reg[233]  ( .D(N251), .CLK(clk), .RST(1'b0), .Q(
        round_reg[233]) );
  DFF \round_reg_reg[234]  ( .D(N252), .CLK(clk), .RST(1'b0), .Q(
        round_reg[234]) );
  DFF \round_reg_reg[235]  ( .D(N253), .CLK(clk), .RST(1'b0), .Q(
        round_reg[235]) );
  DFF \round_reg_reg[236]  ( .D(N254), .CLK(clk), .RST(1'b0), .Q(
        round_reg[236]) );
  DFF \round_reg_reg[237]  ( .D(N255), .CLK(clk), .RST(1'b0), .Q(
        round_reg[237]) );
  DFF \round_reg_reg[238]  ( .D(N256), .CLK(clk), .RST(1'b0), .Q(
        round_reg[238]) );
  DFF \round_reg_reg[239]  ( .D(N257), .CLK(clk), .RST(1'b0), .Q(
        round_reg[239]) );
  DFF \round_reg_reg[240]  ( .D(N258), .CLK(clk), .RST(1'b0), .Q(
        round_reg[240]) );
  DFF \round_reg_reg[241]  ( .D(N259), .CLK(clk), .RST(1'b0), .Q(
        round_reg[241]) );
  DFF \round_reg_reg[242]  ( .D(N260), .CLK(clk), .RST(1'b0), .Q(
        round_reg[242]) );
  DFF \round_reg_reg[243]  ( .D(N261), .CLK(clk), .RST(1'b0), .Q(
        round_reg[243]) );
  DFF \round_reg_reg[244]  ( .D(N262), .CLK(clk), .RST(1'b0), .Q(
        round_reg[244]) );
  DFF \round_reg_reg[245]  ( .D(N263), .CLK(clk), .RST(1'b0), .Q(
        round_reg[245]) );
  DFF \round_reg_reg[246]  ( .D(N264), .CLK(clk), .RST(1'b0), .Q(
        round_reg[246]) );
  DFF \round_reg_reg[247]  ( .D(N265), .CLK(clk), .RST(1'b0), .Q(
        round_reg[247]) );
  DFF \round_reg_reg[248]  ( .D(N266), .CLK(clk), .RST(1'b0), .Q(
        round_reg[248]) );
  DFF \round_reg_reg[249]  ( .D(N267), .CLK(clk), .RST(1'b0), .Q(
        round_reg[249]) );
  DFF \round_reg_reg[250]  ( .D(N268), .CLK(clk), .RST(1'b0), .Q(
        round_reg[250]) );
  DFF \round_reg_reg[251]  ( .D(N269), .CLK(clk), .RST(1'b0), .Q(
        round_reg[251]) );
  DFF \round_reg_reg[252]  ( .D(N270), .CLK(clk), .RST(1'b0), .Q(
        round_reg[252]) );
  DFF \round_reg_reg[253]  ( .D(N271), .CLK(clk), .RST(1'b0), .Q(
        round_reg[253]) );
  DFF \round_reg_reg[254]  ( .D(N272), .CLK(clk), .RST(1'b0), .Q(
        round_reg[254]) );
  DFF \round_reg_reg[255]  ( .D(N273), .CLK(clk), .RST(1'b0), .Q(
        round_reg[255]) );
  DFF \round_reg_reg[256]  ( .D(N274), .CLK(clk), .RST(1'b0), .Q(
        round_reg[256]) );
  DFF \round_reg_reg[257]  ( .D(N275), .CLK(clk), .RST(1'b0), .Q(
        round_reg[257]) );
  DFF \round_reg_reg[258]  ( .D(N276), .CLK(clk), .RST(1'b0), .Q(
        round_reg[258]) );
  DFF \round_reg_reg[259]  ( .D(N277), .CLK(clk), .RST(1'b0), .Q(
        round_reg[259]) );
  DFF \round_reg_reg[260]  ( .D(N278), .CLK(clk), .RST(1'b0), .Q(
        round_reg[260]) );
  DFF \round_reg_reg[261]  ( .D(N279), .CLK(clk), .RST(1'b0), .Q(
        round_reg[261]) );
  DFF \round_reg_reg[262]  ( .D(N280), .CLK(clk), .RST(1'b0), .Q(
        round_reg[262]) );
  DFF \round_reg_reg[263]  ( .D(N281), .CLK(clk), .RST(1'b0), .Q(
        round_reg[263]) );
  DFF \round_reg_reg[264]  ( .D(N282), .CLK(clk), .RST(1'b0), .Q(
        round_reg[264]) );
  DFF \round_reg_reg[265]  ( .D(N283), .CLK(clk), .RST(1'b0), .Q(
        round_reg[265]) );
  DFF \round_reg_reg[266]  ( .D(N284), .CLK(clk), .RST(1'b0), .Q(
        round_reg[266]) );
  DFF \round_reg_reg[267]  ( .D(N285), .CLK(clk), .RST(1'b0), .Q(
        round_reg[267]) );
  DFF \round_reg_reg[268]  ( .D(N286), .CLK(clk), .RST(1'b0), .Q(
        round_reg[268]) );
  DFF \round_reg_reg[269]  ( .D(N287), .CLK(clk), .RST(1'b0), .Q(
        round_reg[269]) );
  DFF \round_reg_reg[270]  ( .D(N288), .CLK(clk), .RST(1'b0), .Q(
        round_reg[270]) );
  DFF \round_reg_reg[271]  ( .D(N289), .CLK(clk), .RST(1'b0), .Q(
        round_reg[271]) );
  DFF \round_reg_reg[272]  ( .D(N290), .CLK(clk), .RST(1'b0), .Q(
        round_reg[272]) );
  DFF \round_reg_reg[273]  ( .D(N291), .CLK(clk), .RST(1'b0), .Q(
        round_reg[273]) );
  DFF \round_reg_reg[274]  ( .D(N292), .CLK(clk), .RST(1'b0), .Q(
        round_reg[274]) );
  DFF \round_reg_reg[275]  ( .D(N293), .CLK(clk), .RST(1'b0), .Q(
        round_reg[275]) );
  DFF \round_reg_reg[276]  ( .D(N294), .CLK(clk), .RST(1'b0), .Q(
        round_reg[276]) );
  DFF \round_reg_reg[277]  ( .D(N295), .CLK(clk), .RST(1'b0), .Q(
        round_reg[277]) );
  DFF \round_reg_reg[278]  ( .D(N296), .CLK(clk), .RST(1'b0), .Q(
        round_reg[278]) );
  DFF \round_reg_reg[279]  ( .D(N297), .CLK(clk), .RST(1'b0), .Q(
        round_reg[279]) );
  DFF \round_reg_reg[280]  ( .D(N298), .CLK(clk), .RST(1'b0), .Q(
        round_reg[280]) );
  DFF \round_reg_reg[281]  ( .D(N299), .CLK(clk), .RST(1'b0), .Q(
        round_reg[281]) );
  DFF \round_reg_reg[282]  ( .D(N300), .CLK(clk), .RST(1'b0), .Q(
        round_reg[282]) );
  DFF \round_reg_reg[283]  ( .D(N301), .CLK(clk), .RST(1'b0), .Q(
        round_reg[283]) );
  DFF \round_reg_reg[284]  ( .D(N302), .CLK(clk), .RST(1'b0), .Q(
        round_reg[284]) );
  DFF \round_reg_reg[285]  ( .D(N303), .CLK(clk), .RST(1'b0), .Q(
        round_reg[285]) );
  DFF \round_reg_reg[286]  ( .D(N304), .CLK(clk), .RST(1'b0), .Q(
        round_reg[286]) );
  DFF \round_reg_reg[287]  ( .D(N305), .CLK(clk), .RST(1'b0), .Q(
        round_reg[287]) );
  DFF \round_reg_reg[288]  ( .D(N306), .CLK(clk), .RST(1'b0), .Q(
        round_reg[288]) );
  DFF \round_reg_reg[289]  ( .D(N307), .CLK(clk), .RST(1'b0), .Q(
        round_reg[289]) );
  DFF \round_reg_reg[290]  ( .D(N308), .CLK(clk), .RST(1'b0), .Q(
        round_reg[290]) );
  DFF \round_reg_reg[291]  ( .D(N309), .CLK(clk), .RST(1'b0), .Q(
        round_reg[291]) );
  DFF \round_reg_reg[292]  ( .D(N310), .CLK(clk), .RST(1'b0), .Q(
        round_reg[292]) );
  DFF \round_reg_reg[293]  ( .D(N311), .CLK(clk), .RST(1'b0), .Q(
        round_reg[293]) );
  DFF \round_reg_reg[294]  ( .D(N312), .CLK(clk), .RST(1'b0), .Q(
        round_reg[294]) );
  DFF \round_reg_reg[295]  ( .D(N313), .CLK(clk), .RST(1'b0), .Q(
        round_reg[295]) );
  DFF \round_reg_reg[296]  ( .D(N314), .CLK(clk), .RST(1'b0), .Q(
        round_reg[296]) );
  DFF \round_reg_reg[297]  ( .D(N315), .CLK(clk), .RST(1'b0), .Q(
        round_reg[297]) );
  DFF \round_reg_reg[298]  ( .D(N316), .CLK(clk), .RST(1'b0), .Q(
        round_reg[298]) );
  DFF \round_reg_reg[299]  ( .D(N317), .CLK(clk), .RST(1'b0), .Q(
        round_reg[299]) );
  DFF \round_reg_reg[300]  ( .D(N318), .CLK(clk), .RST(1'b0), .Q(
        round_reg[300]) );
  DFF \round_reg_reg[301]  ( .D(N319), .CLK(clk), .RST(1'b0), .Q(
        round_reg[301]) );
  DFF \round_reg_reg[302]  ( .D(N320), .CLK(clk), .RST(1'b0), .Q(
        round_reg[302]) );
  DFF \round_reg_reg[303]  ( .D(N321), .CLK(clk), .RST(1'b0), .Q(
        round_reg[303]) );
  DFF \round_reg_reg[304]  ( .D(N322), .CLK(clk), .RST(1'b0), .Q(
        round_reg[304]) );
  DFF \round_reg_reg[305]  ( .D(N323), .CLK(clk), .RST(1'b0), .Q(
        round_reg[305]) );
  DFF \round_reg_reg[306]  ( .D(N324), .CLK(clk), .RST(1'b0), .Q(
        round_reg[306]) );
  DFF \round_reg_reg[307]  ( .D(N325), .CLK(clk), .RST(1'b0), .Q(
        round_reg[307]) );
  DFF \round_reg_reg[308]  ( .D(N326), .CLK(clk), .RST(1'b0), .Q(
        round_reg[308]) );
  DFF \round_reg_reg[309]  ( .D(N327), .CLK(clk), .RST(1'b0), .Q(
        round_reg[309]) );
  DFF \round_reg_reg[310]  ( .D(N328), .CLK(clk), .RST(1'b0), .Q(
        round_reg[310]) );
  DFF \round_reg_reg[311]  ( .D(N329), .CLK(clk), .RST(1'b0), .Q(
        round_reg[311]) );
  DFF \round_reg_reg[312]  ( .D(N330), .CLK(clk), .RST(1'b0), .Q(
        round_reg[312]) );
  DFF \round_reg_reg[313]  ( .D(N331), .CLK(clk), .RST(1'b0), .Q(
        round_reg[313]) );
  DFF \round_reg_reg[314]  ( .D(N332), .CLK(clk), .RST(1'b0), .Q(
        round_reg[314]) );
  DFF \round_reg_reg[315]  ( .D(N333), .CLK(clk), .RST(1'b0), .Q(
        round_reg[315]) );
  DFF \round_reg_reg[316]  ( .D(N334), .CLK(clk), .RST(1'b0), .Q(
        round_reg[316]) );
  DFF \round_reg_reg[317]  ( .D(N335), .CLK(clk), .RST(1'b0), .Q(
        round_reg[317]) );
  DFF \round_reg_reg[318]  ( .D(N336), .CLK(clk), .RST(1'b0), .Q(
        round_reg[318]) );
  DFF \round_reg_reg[319]  ( .D(N337), .CLK(clk), .RST(1'b0), .Q(
        round_reg[319]) );
  DFF \round_reg_reg[320]  ( .D(N338), .CLK(clk), .RST(1'b0), .Q(
        round_reg[320]) );
  DFF \round_reg_reg[321]  ( .D(N339), .CLK(clk), .RST(1'b0), .Q(
        round_reg[321]) );
  DFF \round_reg_reg[322]  ( .D(N340), .CLK(clk), .RST(1'b0), .Q(
        round_reg[322]) );
  DFF \round_reg_reg[323]  ( .D(N341), .CLK(clk), .RST(1'b0), .Q(
        round_reg[323]) );
  DFF \round_reg_reg[324]  ( .D(N342), .CLK(clk), .RST(1'b0), .Q(
        round_reg[324]) );
  DFF \round_reg_reg[325]  ( .D(N343), .CLK(clk), .RST(1'b0), .Q(
        round_reg[325]) );
  DFF \round_reg_reg[326]  ( .D(N344), .CLK(clk), .RST(1'b0), .Q(
        round_reg[326]) );
  DFF \round_reg_reg[327]  ( .D(N345), .CLK(clk), .RST(1'b0), .Q(
        round_reg[327]) );
  DFF \round_reg_reg[328]  ( .D(N346), .CLK(clk), .RST(1'b0), .Q(
        round_reg[328]) );
  DFF \round_reg_reg[329]  ( .D(N347), .CLK(clk), .RST(1'b0), .Q(
        round_reg[329]) );
  DFF \round_reg_reg[330]  ( .D(N348), .CLK(clk), .RST(1'b0), .Q(
        round_reg[330]) );
  DFF \round_reg_reg[331]  ( .D(N349), .CLK(clk), .RST(1'b0), .Q(
        round_reg[331]) );
  DFF \round_reg_reg[332]  ( .D(N350), .CLK(clk), .RST(1'b0), .Q(
        round_reg[332]) );
  DFF \round_reg_reg[333]  ( .D(N351), .CLK(clk), .RST(1'b0), .Q(
        round_reg[333]) );
  DFF \round_reg_reg[334]  ( .D(N352), .CLK(clk), .RST(1'b0), .Q(
        round_reg[334]) );
  DFF \round_reg_reg[335]  ( .D(N353), .CLK(clk), .RST(1'b0), .Q(
        round_reg[335]) );
  DFF \round_reg_reg[336]  ( .D(N354), .CLK(clk), .RST(1'b0), .Q(
        round_reg[336]) );
  DFF \round_reg_reg[337]  ( .D(N355), .CLK(clk), .RST(1'b0), .Q(
        round_reg[337]) );
  DFF \round_reg_reg[338]  ( .D(N356), .CLK(clk), .RST(1'b0), .Q(
        round_reg[338]) );
  DFF \round_reg_reg[339]  ( .D(N357), .CLK(clk), .RST(1'b0), .Q(
        round_reg[339]) );
  DFF \round_reg_reg[340]  ( .D(N358), .CLK(clk), .RST(1'b0), .Q(
        round_reg[340]) );
  DFF \round_reg_reg[341]  ( .D(N359), .CLK(clk), .RST(1'b0), .Q(
        round_reg[341]) );
  DFF \round_reg_reg[342]  ( .D(N360), .CLK(clk), .RST(1'b0), .Q(
        round_reg[342]) );
  DFF \round_reg_reg[343]  ( .D(N361), .CLK(clk), .RST(1'b0), .Q(
        round_reg[343]) );
  DFF \round_reg_reg[344]  ( .D(N362), .CLK(clk), .RST(1'b0), .Q(
        round_reg[344]) );
  DFF \round_reg_reg[345]  ( .D(N363), .CLK(clk), .RST(1'b0), .Q(
        round_reg[345]) );
  DFF \round_reg_reg[346]  ( .D(N364), .CLK(clk), .RST(1'b0), .Q(
        round_reg[346]) );
  DFF \round_reg_reg[347]  ( .D(N365), .CLK(clk), .RST(1'b0), .Q(
        round_reg[347]) );
  DFF \round_reg_reg[348]  ( .D(N366), .CLK(clk), .RST(1'b0), .Q(
        round_reg[348]) );
  DFF \round_reg_reg[349]  ( .D(N367), .CLK(clk), .RST(1'b0), .Q(
        round_reg[349]) );
  DFF \round_reg_reg[350]  ( .D(N368), .CLK(clk), .RST(1'b0), .Q(
        round_reg[350]) );
  DFF \round_reg_reg[351]  ( .D(N369), .CLK(clk), .RST(1'b0), .Q(
        round_reg[351]) );
  DFF \round_reg_reg[352]  ( .D(N370), .CLK(clk), .RST(1'b0), .Q(
        round_reg[352]) );
  DFF \round_reg_reg[353]  ( .D(N371), .CLK(clk), .RST(1'b0), .Q(
        round_reg[353]) );
  DFF \round_reg_reg[354]  ( .D(N372), .CLK(clk), .RST(1'b0), .Q(
        round_reg[354]) );
  DFF \round_reg_reg[355]  ( .D(N373), .CLK(clk), .RST(1'b0), .Q(
        round_reg[355]) );
  DFF \round_reg_reg[356]  ( .D(N374), .CLK(clk), .RST(1'b0), .Q(
        round_reg[356]) );
  DFF \round_reg_reg[357]  ( .D(N375), .CLK(clk), .RST(1'b0), .Q(
        round_reg[357]) );
  DFF \round_reg_reg[358]  ( .D(N376), .CLK(clk), .RST(1'b0), .Q(
        round_reg[358]) );
  DFF \round_reg_reg[359]  ( .D(N377), .CLK(clk), .RST(1'b0), .Q(
        round_reg[359]) );
  DFF \round_reg_reg[360]  ( .D(N378), .CLK(clk), .RST(1'b0), .Q(
        round_reg[360]) );
  DFF \round_reg_reg[361]  ( .D(N379), .CLK(clk), .RST(1'b0), .Q(
        round_reg[361]) );
  DFF \round_reg_reg[362]  ( .D(N380), .CLK(clk), .RST(1'b0), .Q(
        round_reg[362]) );
  DFF \round_reg_reg[363]  ( .D(N381), .CLK(clk), .RST(1'b0), .Q(
        round_reg[363]) );
  DFF \round_reg_reg[364]  ( .D(N382), .CLK(clk), .RST(1'b0), .Q(
        round_reg[364]) );
  DFF \round_reg_reg[365]  ( .D(N383), .CLK(clk), .RST(1'b0), .Q(
        round_reg[365]) );
  DFF \round_reg_reg[366]  ( .D(N384), .CLK(clk), .RST(1'b0), .Q(
        round_reg[366]) );
  DFF \round_reg_reg[367]  ( .D(N385), .CLK(clk), .RST(1'b0), .Q(
        round_reg[367]) );
  DFF \round_reg_reg[368]  ( .D(N386), .CLK(clk), .RST(1'b0), .Q(
        round_reg[368]) );
  DFF \round_reg_reg[369]  ( .D(N387), .CLK(clk), .RST(1'b0), .Q(
        round_reg[369]) );
  DFF \round_reg_reg[370]  ( .D(N388), .CLK(clk), .RST(1'b0), .Q(
        round_reg[370]) );
  DFF \round_reg_reg[371]  ( .D(N389), .CLK(clk), .RST(1'b0), .Q(
        round_reg[371]) );
  DFF \round_reg_reg[372]  ( .D(N390), .CLK(clk), .RST(1'b0), .Q(
        round_reg[372]) );
  DFF \round_reg_reg[373]  ( .D(N391), .CLK(clk), .RST(1'b0), .Q(
        round_reg[373]) );
  DFF \round_reg_reg[374]  ( .D(N392), .CLK(clk), .RST(1'b0), .Q(
        round_reg[374]) );
  DFF \round_reg_reg[375]  ( .D(N393), .CLK(clk), .RST(1'b0), .Q(
        round_reg[375]) );
  DFF \round_reg_reg[376]  ( .D(N394), .CLK(clk), .RST(1'b0), .Q(
        round_reg[376]) );
  DFF \round_reg_reg[377]  ( .D(N395), .CLK(clk), .RST(1'b0), .Q(
        round_reg[377]) );
  DFF \round_reg_reg[378]  ( .D(N396), .CLK(clk), .RST(1'b0), .Q(
        round_reg[378]) );
  DFF \round_reg_reg[379]  ( .D(N397), .CLK(clk), .RST(1'b0), .Q(
        round_reg[379]) );
  DFF \round_reg_reg[380]  ( .D(N398), .CLK(clk), .RST(1'b0), .Q(
        round_reg[380]) );
  DFF \round_reg_reg[381]  ( .D(N399), .CLK(clk), .RST(1'b0), .Q(
        round_reg[381]) );
  DFF \round_reg_reg[382]  ( .D(N400), .CLK(clk), .RST(1'b0), .Q(
        round_reg[382]) );
  DFF \round_reg_reg[383]  ( .D(N401), .CLK(clk), .RST(1'b0), .Q(
        round_reg[383]) );
  DFF \round_reg_reg[384]  ( .D(N402), .CLK(clk), .RST(1'b0), .Q(
        round_reg[384]) );
  DFF \round_reg_reg[385]  ( .D(N403), .CLK(clk), .RST(1'b0), .Q(
        round_reg[385]) );
  DFF \round_reg_reg[386]  ( .D(N404), .CLK(clk), .RST(1'b0), .Q(
        round_reg[386]) );
  DFF \round_reg_reg[387]  ( .D(N405), .CLK(clk), .RST(1'b0), .Q(
        round_reg[387]) );
  DFF \round_reg_reg[388]  ( .D(N406), .CLK(clk), .RST(1'b0), .Q(
        round_reg[388]) );
  DFF \round_reg_reg[389]  ( .D(N407), .CLK(clk), .RST(1'b0), .Q(
        round_reg[389]) );
  DFF \round_reg_reg[390]  ( .D(N408), .CLK(clk), .RST(1'b0), .Q(
        round_reg[390]) );
  DFF \round_reg_reg[391]  ( .D(N409), .CLK(clk), .RST(1'b0), .Q(
        round_reg[391]) );
  DFF \round_reg_reg[392]  ( .D(N410), .CLK(clk), .RST(1'b0), .Q(
        round_reg[392]) );
  DFF \round_reg_reg[393]  ( .D(N411), .CLK(clk), .RST(1'b0), .Q(
        round_reg[393]) );
  DFF \round_reg_reg[394]  ( .D(N412), .CLK(clk), .RST(1'b0), .Q(
        round_reg[394]) );
  DFF \round_reg_reg[395]  ( .D(N413), .CLK(clk), .RST(1'b0), .Q(
        round_reg[395]) );
  DFF \round_reg_reg[396]  ( .D(N414), .CLK(clk), .RST(1'b0), .Q(
        round_reg[396]) );
  DFF \round_reg_reg[397]  ( .D(N415), .CLK(clk), .RST(1'b0), .Q(
        round_reg[397]) );
  DFF \round_reg_reg[398]  ( .D(N416), .CLK(clk), .RST(1'b0), .Q(
        round_reg[398]) );
  DFF \round_reg_reg[399]  ( .D(N417), .CLK(clk), .RST(1'b0), .Q(
        round_reg[399]) );
  DFF \round_reg_reg[400]  ( .D(N418), .CLK(clk), .RST(1'b0), .Q(
        round_reg[400]) );
  DFF \round_reg_reg[401]  ( .D(N419), .CLK(clk), .RST(1'b0), .Q(
        round_reg[401]) );
  DFF \round_reg_reg[402]  ( .D(N420), .CLK(clk), .RST(1'b0), .Q(
        round_reg[402]) );
  DFF \round_reg_reg[403]  ( .D(N421), .CLK(clk), .RST(1'b0), .Q(
        round_reg[403]) );
  DFF \round_reg_reg[404]  ( .D(N422), .CLK(clk), .RST(1'b0), .Q(
        round_reg[404]) );
  DFF \round_reg_reg[405]  ( .D(N423), .CLK(clk), .RST(1'b0), .Q(
        round_reg[405]) );
  DFF \round_reg_reg[406]  ( .D(N424), .CLK(clk), .RST(1'b0), .Q(
        round_reg[406]) );
  DFF \round_reg_reg[407]  ( .D(N425), .CLK(clk), .RST(1'b0), .Q(
        round_reg[407]) );
  DFF \round_reg_reg[408]  ( .D(N426), .CLK(clk), .RST(1'b0), .Q(
        round_reg[408]) );
  DFF \round_reg_reg[409]  ( .D(N427), .CLK(clk), .RST(1'b0), .Q(
        round_reg[409]) );
  DFF \round_reg_reg[410]  ( .D(N428), .CLK(clk), .RST(1'b0), .Q(
        round_reg[410]) );
  DFF \round_reg_reg[411]  ( .D(N429), .CLK(clk), .RST(1'b0), .Q(
        round_reg[411]) );
  DFF \round_reg_reg[412]  ( .D(N430), .CLK(clk), .RST(1'b0), .Q(
        round_reg[412]) );
  DFF \round_reg_reg[413]  ( .D(N431), .CLK(clk), .RST(1'b0), .Q(
        round_reg[413]) );
  DFF \round_reg_reg[414]  ( .D(N432), .CLK(clk), .RST(1'b0), .Q(
        round_reg[414]) );
  DFF \round_reg_reg[415]  ( .D(N433), .CLK(clk), .RST(1'b0), .Q(
        round_reg[415]) );
  DFF \round_reg_reg[416]  ( .D(N434), .CLK(clk), .RST(1'b0), .Q(
        round_reg[416]) );
  DFF \round_reg_reg[417]  ( .D(N435), .CLK(clk), .RST(1'b0), .Q(
        round_reg[417]) );
  DFF \round_reg_reg[418]  ( .D(N436), .CLK(clk), .RST(1'b0), .Q(
        round_reg[418]) );
  DFF \round_reg_reg[419]  ( .D(N437), .CLK(clk), .RST(1'b0), .Q(
        round_reg[419]) );
  DFF \round_reg_reg[420]  ( .D(N438), .CLK(clk), .RST(1'b0), .Q(
        round_reg[420]) );
  DFF \round_reg_reg[421]  ( .D(N439), .CLK(clk), .RST(1'b0), .Q(
        round_reg[421]) );
  DFF \round_reg_reg[422]  ( .D(N440), .CLK(clk), .RST(1'b0), .Q(
        round_reg[422]) );
  DFF \round_reg_reg[423]  ( .D(N441), .CLK(clk), .RST(1'b0), .Q(
        round_reg[423]) );
  DFF \round_reg_reg[424]  ( .D(N442), .CLK(clk), .RST(1'b0), .Q(
        round_reg[424]) );
  DFF \round_reg_reg[425]  ( .D(N443), .CLK(clk), .RST(1'b0), .Q(
        round_reg[425]) );
  DFF \round_reg_reg[426]  ( .D(N444), .CLK(clk), .RST(1'b0), .Q(
        round_reg[426]) );
  DFF \round_reg_reg[427]  ( .D(N445), .CLK(clk), .RST(1'b0), .Q(
        round_reg[427]) );
  DFF \round_reg_reg[428]  ( .D(N446), .CLK(clk), .RST(1'b0), .Q(
        round_reg[428]) );
  DFF \round_reg_reg[429]  ( .D(N447), .CLK(clk), .RST(1'b0), .Q(
        round_reg[429]) );
  DFF \round_reg_reg[430]  ( .D(N448), .CLK(clk), .RST(1'b0), .Q(
        round_reg[430]) );
  DFF \round_reg_reg[431]  ( .D(N449), .CLK(clk), .RST(1'b0), .Q(
        round_reg[431]) );
  DFF \round_reg_reg[432]  ( .D(N450), .CLK(clk), .RST(1'b0), .Q(
        round_reg[432]) );
  DFF \round_reg_reg[433]  ( .D(N451), .CLK(clk), .RST(1'b0), .Q(
        round_reg[433]) );
  DFF \round_reg_reg[434]  ( .D(N452), .CLK(clk), .RST(1'b0), .Q(
        round_reg[434]) );
  DFF \round_reg_reg[435]  ( .D(N453), .CLK(clk), .RST(1'b0), .Q(
        round_reg[435]) );
  DFF \round_reg_reg[436]  ( .D(N454), .CLK(clk), .RST(1'b0), .Q(
        round_reg[436]) );
  DFF \round_reg_reg[437]  ( .D(N455), .CLK(clk), .RST(1'b0), .Q(
        round_reg[437]) );
  DFF \round_reg_reg[438]  ( .D(N456), .CLK(clk), .RST(1'b0), .Q(
        round_reg[438]) );
  DFF \round_reg_reg[439]  ( .D(N457), .CLK(clk), .RST(1'b0), .Q(
        round_reg[439]) );
  DFF \round_reg_reg[440]  ( .D(N458), .CLK(clk), .RST(1'b0), .Q(
        round_reg[440]) );
  DFF \round_reg_reg[441]  ( .D(N459), .CLK(clk), .RST(1'b0), .Q(
        round_reg[441]) );
  DFF \round_reg_reg[442]  ( .D(N460), .CLK(clk), .RST(1'b0), .Q(
        round_reg[442]) );
  DFF \round_reg_reg[443]  ( .D(N461), .CLK(clk), .RST(1'b0), .Q(
        round_reg[443]) );
  DFF \round_reg_reg[444]  ( .D(N462), .CLK(clk), .RST(1'b0), .Q(
        round_reg[444]) );
  DFF \round_reg_reg[445]  ( .D(N463), .CLK(clk), .RST(1'b0), .Q(
        round_reg[445]) );
  DFF \round_reg_reg[446]  ( .D(N464), .CLK(clk), .RST(1'b0), .Q(
        round_reg[446]) );
  DFF \round_reg_reg[447]  ( .D(N465), .CLK(clk), .RST(1'b0), .Q(
        round_reg[447]) );
  DFF \round_reg_reg[448]  ( .D(N466), .CLK(clk), .RST(1'b0), .Q(
        round_reg[448]) );
  DFF \round_reg_reg[449]  ( .D(N467), .CLK(clk), .RST(1'b0), .Q(
        round_reg[449]) );
  DFF \round_reg_reg[450]  ( .D(N468), .CLK(clk), .RST(1'b0), .Q(
        round_reg[450]) );
  DFF \round_reg_reg[451]  ( .D(N469), .CLK(clk), .RST(1'b0), .Q(
        round_reg[451]) );
  DFF \round_reg_reg[452]  ( .D(N470), .CLK(clk), .RST(1'b0), .Q(
        round_reg[452]) );
  DFF \round_reg_reg[453]  ( .D(N471), .CLK(clk), .RST(1'b0), .Q(
        round_reg[453]) );
  DFF \round_reg_reg[454]  ( .D(N472), .CLK(clk), .RST(1'b0), .Q(
        round_reg[454]) );
  DFF \round_reg_reg[455]  ( .D(N473), .CLK(clk), .RST(1'b0), .Q(
        round_reg[455]) );
  DFF \round_reg_reg[456]  ( .D(N474), .CLK(clk), .RST(1'b0), .Q(
        round_reg[456]) );
  DFF \round_reg_reg[457]  ( .D(N475), .CLK(clk), .RST(1'b0), .Q(
        round_reg[457]) );
  DFF \round_reg_reg[458]  ( .D(N476), .CLK(clk), .RST(1'b0), .Q(
        round_reg[458]) );
  DFF \round_reg_reg[459]  ( .D(N477), .CLK(clk), .RST(1'b0), .Q(
        round_reg[459]) );
  DFF \round_reg_reg[460]  ( .D(N478), .CLK(clk), .RST(1'b0), .Q(
        round_reg[460]) );
  DFF \round_reg_reg[461]  ( .D(N479), .CLK(clk), .RST(1'b0), .Q(
        round_reg[461]) );
  DFF \round_reg_reg[462]  ( .D(N480), .CLK(clk), .RST(1'b0), .Q(
        round_reg[462]) );
  DFF \round_reg_reg[463]  ( .D(N481), .CLK(clk), .RST(1'b0), .Q(
        round_reg[463]) );
  DFF \round_reg_reg[464]  ( .D(N482), .CLK(clk), .RST(1'b0), .Q(
        round_reg[464]) );
  DFF \round_reg_reg[465]  ( .D(N483), .CLK(clk), .RST(1'b0), .Q(
        round_reg[465]) );
  DFF \round_reg_reg[466]  ( .D(N484), .CLK(clk), .RST(1'b0), .Q(
        round_reg[466]) );
  DFF \round_reg_reg[467]  ( .D(N485), .CLK(clk), .RST(1'b0), .Q(
        round_reg[467]) );
  DFF \round_reg_reg[468]  ( .D(N486), .CLK(clk), .RST(1'b0), .Q(
        round_reg[468]) );
  DFF \round_reg_reg[469]  ( .D(N487), .CLK(clk), .RST(1'b0), .Q(
        round_reg[469]) );
  DFF \round_reg_reg[470]  ( .D(N488), .CLK(clk), .RST(1'b0), .Q(
        round_reg[470]) );
  DFF \round_reg_reg[471]  ( .D(N489), .CLK(clk), .RST(1'b0), .Q(
        round_reg[471]) );
  DFF \round_reg_reg[472]  ( .D(N490), .CLK(clk), .RST(1'b0), .Q(
        round_reg[472]) );
  DFF \round_reg_reg[473]  ( .D(N491), .CLK(clk), .RST(1'b0), .Q(
        round_reg[473]) );
  DFF \round_reg_reg[474]  ( .D(N492), .CLK(clk), .RST(1'b0), .Q(
        round_reg[474]) );
  DFF \round_reg_reg[475]  ( .D(N493), .CLK(clk), .RST(1'b0), .Q(
        round_reg[475]) );
  DFF \round_reg_reg[476]  ( .D(N494), .CLK(clk), .RST(1'b0), .Q(
        round_reg[476]) );
  DFF \round_reg_reg[477]  ( .D(N495), .CLK(clk), .RST(1'b0), .Q(
        round_reg[477]) );
  DFF \round_reg_reg[478]  ( .D(N496), .CLK(clk), .RST(1'b0), .Q(
        round_reg[478]) );
  DFF \round_reg_reg[479]  ( .D(N497), .CLK(clk), .RST(1'b0), .Q(
        round_reg[479]) );
  DFF \round_reg_reg[480]  ( .D(N498), .CLK(clk), .RST(1'b0), .Q(
        round_reg[480]) );
  DFF \round_reg_reg[481]  ( .D(N499), .CLK(clk), .RST(1'b0), .Q(
        round_reg[481]) );
  DFF \round_reg_reg[482]  ( .D(N500), .CLK(clk), .RST(1'b0), .Q(
        round_reg[482]) );
  DFF \round_reg_reg[483]  ( .D(N501), .CLK(clk), .RST(1'b0), .Q(
        round_reg[483]) );
  DFF \round_reg_reg[484]  ( .D(N502), .CLK(clk), .RST(1'b0), .Q(
        round_reg[484]) );
  DFF \round_reg_reg[485]  ( .D(N503), .CLK(clk), .RST(1'b0), .Q(
        round_reg[485]) );
  DFF \round_reg_reg[486]  ( .D(N504), .CLK(clk), .RST(1'b0), .Q(
        round_reg[486]) );
  DFF \round_reg_reg[487]  ( .D(N505), .CLK(clk), .RST(1'b0), .Q(
        round_reg[487]) );
  DFF \round_reg_reg[488]  ( .D(N506), .CLK(clk), .RST(1'b0), .Q(
        round_reg[488]) );
  DFF \round_reg_reg[489]  ( .D(N507), .CLK(clk), .RST(1'b0), .Q(
        round_reg[489]) );
  DFF \round_reg_reg[490]  ( .D(N508), .CLK(clk), .RST(1'b0), .Q(
        round_reg[490]) );
  DFF \round_reg_reg[491]  ( .D(N509), .CLK(clk), .RST(1'b0), .Q(
        round_reg[491]) );
  DFF \round_reg_reg[492]  ( .D(N510), .CLK(clk), .RST(1'b0), .Q(
        round_reg[492]) );
  DFF \round_reg_reg[493]  ( .D(N511), .CLK(clk), .RST(1'b0), .Q(
        round_reg[493]) );
  DFF \round_reg_reg[494]  ( .D(N512), .CLK(clk), .RST(1'b0), .Q(
        round_reg[494]) );
  DFF \round_reg_reg[495]  ( .D(N513), .CLK(clk), .RST(1'b0), .Q(
        round_reg[495]) );
  DFF \round_reg_reg[496]  ( .D(N514), .CLK(clk), .RST(1'b0), .Q(
        round_reg[496]) );
  DFF \round_reg_reg[497]  ( .D(N515), .CLK(clk), .RST(1'b0), .Q(
        round_reg[497]) );
  DFF \round_reg_reg[498]  ( .D(N516), .CLK(clk), .RST(1'b0), .Q(
        round_reg[498]) );
  DFF \round_reg_reg[499]  ( .D(N517), .CLK(clk), .RST(1'b0), .Q(
        round_reg[499]) );
  DFF \round_reg_reg[500]  ( .D(N518), .CLK(clk), .RST(1'b0), .Q(
        round_reg[500]) );
  DFF \round_reg_reg[501]  ( .D(N519), .CLK(clk), .RST(1'b0), .Q(
        round_reg[501]) );
  DFF \round_reg_reg[502]  ( .D(N520), .CLK(clk), .RST(1'b0), .Q(
        round_reg[502]) );
  DFF \round_reg_reg[503]  ( .D(N521), .CLK(clk), .RST(1'b0), .Q(
        round_reg[503]) );
  DFF \round_reg_reg[504]  ( .D(N522), .CLK(clk), .RST(1'b0), .Q(
        round_reg[504]) );
  DFF \round_reg_reg[505]  ( .D(N523), .CLK(clk), .RST(1'b0), .Q(
        round_reg[505]) );
  DFF \round_reg_reg[506]  ( .D(N524), .CLK(clk), .RST(1'b0), .Q(
        round_reg[506]) );
  DFF \round_reg_reg[507]  ( .D(N525), .CLK(clk), .RST(1'b0), .Q(
        round_reg[507]) );
  DFF \round_reg_reg[508]  ( .D(N526), .CLK(clk), .RST(1'b0), .Q(
        round_reg[508]) );
  DFF \round_reg_reg[509]  ( .D(N527), .CLK(clk), .RST(1'b0), .Q(
        round_reg[509]) );
  DFF \round_reg_reg[510]  ( .D(N528), .CLK(clk), .RST(1'b0), .Q(
        round_reg[510]) );
  DFF \round_reg_reg[511]  ( .D(N529), .CLK(clk), .RST(1'b0), .Q(
        round_reg[511]) );
  DFF \round_reg_reg[512]  ( .D(N530), .CLK(clk), .RST(1'b0), .Q(
        round_reg[512]) );
  DFF \round_reg_reg[513]  ( .D(N531), .CLK(clk), .RST(1'b0), .Q(
        round_reg[513]) );
  DFF \round_reg_reg[514]  ( .D(N532), .CLK(clk), .RST(1'b0), .Q(
        round_reg[514]) );
  DFF \round_reg_reg[515]  ( .D(N533), .CLK(clk), .RST(1'b0), .Q(
        round_reg[515]) );
  DFF \round_reg_reg[516]  ( .D(N534), .CLK(clk), .RST(1'b0), .Q(
        round_reg[516]) );
  DFF \round_reg_reg[517]  ( .D(N535), .CLK(clk), .RST(1'b0), .Q(
        round_reg[517]) );
  DFF \round_reg_reg[518]  ( .D(N536), .CLK(clk), .RST(1'b0), .Q(
        round_reg[518]) );
  DFF \round_reg_reg[519]  ( .D(N537), .CLK(clk), .RST(1'b0), .Q(
        round_reg[519]) );
  DFF \round_reg_reg[520]  ( .D(N538), .CLK(clk), .RST(1'b0), .Q(
        round_reg[520]) );
  DFF \round_reg_reg[521]  ( .D(N539), .CLK(clk), .RST(1'b0), .Q(
        round_reg[521]) );
  DFF \round_reg_reg[522]  ( .D(N540), .CLK(clk), .RST(1'b0), .Q(
        round_reg[522]) );
  DFF \round_reg_reg[523]  ( .D(N541), .CLK(clk), .RST(1'b0), .Q(
        round_reg[523]) );
  DFF \round_reg_reg[524]  ( .D(N542), .CLK(clk), .RST(1'b0), .Q(
        round_reg[524]) );
  DFF \round_reg_reg[525]  ( .D(N543), .CLK(clk), .RST(1'b0), .Q(
        round_reg[525]) );
  DFF \round_reg_reg[526]  ( .D(N544), .CLK(clk), .RST(1'b0), .Q(
        round_reg[526]) );
  DFF \round_reg_reg[527]  ( .D(N545), .CLK(clk), .RST(1'b0), .Q(
        round_reg[527]) );
  DFF \round_reg_reg[528]  ( .D(N546), .CLK(clk), .RST(1'b0), .Q(
        round_reg[528]) );
  DFF \round_reg_reg[529]  ( .D(N547), .CLK(clk), .RST(1'b0), .Q(
        round_reg[529]) );
  DFF \round_reg_reg[530]  ( .D(N548), .CLK(clk), .RST(1'b0), .Q(
        round_reg[530]) );
  DFF \round_reg_reg[531]  ( .D(N549), .CLK(clk), .RST(1'b0), .Q(
        round_reg[531]) );
  DFF \round_reg_reg[532]  ( .D(N550), .CLK(clk), .RST(1'b0), .Q(
        round_reg[532]) );
  DFF \round_reg_reg[533]  ( .D(N551), .CLK(clk), .RST(1'b0), .Q(
        round_reg[533]) );
  DFF \round_reg_reg[534]  ( .D(N552), .CLK(clk), .RST(1'b0), .Q(
        round_reg[534]) );
  DFF \round_reg_reg[535]  ( .D(N553), .CLK(clk), .RST(1'b0), .Q(
        round_reg[535]) );
  DFF \round_reg_reg[536]  ( .D(N554), .CLK(clk), .RST(1'b0), .Q(
        round_reg[536]) );
  DFF \round_reg_reg[537]  ( .D(N555), .CLK(clk), .RST(1'b0), .Q(
        round_reg[537]) );
  DFF \round_reg_reg[538]  ( .D(N556), .CLK(clk), .RST(1'b0), .Q(
        round_reg[538]) );
  DFF \round_reg_reg[539]  ( .D(N557), .CLK(clk), .RST(1'b0), .Q(
        round_reg[539]) );
  DFF \round_reg_reg[540]  ( .D(N558), .CLK(clk), .RST(1'b0), .Q(
        round_reg[540]) );
  DFF \round_reg_reg[541]  ( .D(N559), .CLK(clk), .RST(1'b0), .Q(
        round_reg[541]) );
  DFF \round_reg_reg[542]  ( .D(N560), .CLK(clk), .RST(1'b0), .Q(
        round_reg[542]) );
  DFF \round_reg_reg[543]  ( .D(N561), .CLK(clk), .RST(1'b0), .Q(
        round_reg[543]) );
  DFF \round_reg_reg[544]  ( .D(N562), .CLK(clk), .RST(1'b0), .Q(
        round_reg[544]) );
  DFF \round_reg_reg[545]  ( .D(N563), .CLK(clk), .RST(1'b0), .Q(
        round_reg[545]) );
  DFF \round_reg_reg[546]  ( .D(N564), .CLK(clk), .RST(1'b0), .Q(
        round_reg[546]) );
  DFF \round_reg_reg[547]  ( .D(N565), .CLK(clk), .RST(1'b0), .Q(
        round_reg[547]) );
  DFF \round_reg_reg[548]  ( .D(N566), .CLK(clk), .RST(1'b0), .Q(
        round_reg[548]) );
  DFF \round_reg_reg[549]  ( .D(N567), .CLK(clk), .RST(1'b0), .Q(
        round_reg[549]) );
  DFF \round_reg_reg[550]  ( .D(N568), .CLK(clk), .RST(1'b0), .Q(
        round_reg[550]) );
  DFF \round_reg_reg[551]  ( .D(N569), .CLK(clk), .RST(1'b0), .Q(
        round_reg[551]) );
  DFF \round_reg_reg[552]  ( .D(N570), .CLK(clk), .RST(1'b0), .Q(
        round_reg[552]) );
  DFF \round_reg_reg[553]  ( .D(N571), .CLK(clk), .RST(1'b0), .Q(
        round_reg[553]) );
  DFF \round_reg_reg[554]  ( .D(N572), .CLK(clk), .RST(1'b0), .Q(
        round_reg[554]) );
  DFF \round_reg_reg[555]  ( .D(N573), .CLK(clk), .RST(1'b0), .Q(
        round_reg[555]) );
  DFF \round_reg_reg[556]  ( .D(N574), .CLK(clk), .RST(1'b0), .Q(
        round_reg[556]) );
  DFF \round_reg_reg[557]  ( .D(N575), .CLK(clk), .RST(1'b0), .Q(
        round_reg[557]) );
  DFF \round_reg_reg[558]  ( .D(N576), .CLK(clk), .RST(1'b0), .Q(
        round_reg[558]) );
  DFF \round_reg_reg[559]  ( .D(N577), .CLK(clk), .RST(1'b0), .Q(
        round_reg[559]) );
  DFF \round_reg_reg[560]  ( .D(N578), .CLK(clk), .RST(1'b0), .Q(
        round_reg[560]) );
  DFF \round_reg_reg[561]  ( .D(N579), .CLK(clk), .RST(1'b0), .Q(
        round_reg[561]) );
  DFF \round_reg_reg[562]  ( .D(N580), .CLK(clk), .RST(1'b0), .Q(
        round_reg[562]) );
  DFF \round_reg_reg[563]  ( .D(N581), .CLK(clk), .RST(1'b0), .Q(
        round_reg[563]) );
  DFF \round_reg_reg[564]  ( .D(N582), .CLK(clk), .RST(1'b0), .Q(
        round_reg[564]) );
  DFF \round_reg_reg[565]  ( .D(N583), .CLK(clk), .RST(1'b0), .Q(
        round_reg[565]) );
  DFF \round_reg_reg[566]  ( .D(N584), .CLK(clk), .RST(1'b0), .Q(
        round_reg[566]) );
  DFF \round_reg_reg[567]  ( .D(N585), .CLK(clk), .RST(1'b0), .Q(
        round_reg[567]) );
  DFF \round_reg_reg[568]  ( .D(N586), .CLK(clk), .RST(1'b0), .Q(
        round_reg[568]) );
  DFF \round_reg_reg[569]  ( .D(N587), .CLK(clk), .RST(1'b0), .Q(
        round_reg[569]) );
  DFF \round_reg_reg[570]  ( .D(N588), .CLK(clk), .RST(1'b0), .Q(
        round_reg[570]) );
  DFF \round_reg_reg[571]  ( .D(N589), .CLK(clk), .RST(1'b0), .Q(
        round_reg[571]) );
  DFF \round_reg_reg[572]  ( .D(N590), .CLK(clk), .RST(1'b0), .Q(
        round_reg[572]) );
  DFF \round_reg_reg[573]  ( .D(N591), .CLK(clk), .RST(1'b0), .Q(
        round_reg[573]) );
  DFF \round_reg_reg[574]  ( .D(N592), .CLK(clk), .RST(1'b0), .Q(
        round_reg[574]) );
  DFF \round_reg_reg[575]  ( .D(N593), .CLK(clk), .RST(1'b0), .Q(
        round_reg[575]) );
  DFF \round_reg_reg[576]  ( .D(N594), .CLK(clk), .RST(1'b0), .Q(
        round_reg[576]) );
  DFF \round_reg_reg[577]  ( .D(N595), .CLK(clk), .RST(1'b0), .Q(
        round_reg[577]) );
  DFF \round_reg_reg[578]  ( .D(N596), .CLK(clk), .RST(1'b0), .Q(
        round_reg[578]) );
  DFF \round_reg_reg[579]  ( .D(N597), .CLK(clk), .RST(1'b0), .Q(
        round_reg[579]) );
  DFF \round_reg_reg[580]  ( .D(N598), .CLK(clk), .RST(1'b0), .Q(
        round_reg[580]) );
  DFF \round_reg_reg[581]  ( .D(N599), .CLK(clk), .RST(1'b0), .Q(
        round_reg[581]) );
  DFF \round_reg_reg[582]  ( .D(N600), .CLK(clk), .RST(1'b0), .Q(
        round_reg[582]) );
  DFF \round_reg_reg[583]  ( .D(N601), .CLK(clk), .RST(1'b0), .Q(
        round_reg[583]) );
  DFF \round_reg_reg[584]  ( .D(N602), .CLK(clk), .RST(1'b0), .Q(
        round_reg[584]) );
  DFF \round_reg_reg[585]  ( .D(N603), .CLK(clk), .RST(1'b0), .Q(
        round_reg[585]) );
  DFF \round_reg_reg[586]  ( .D(N604), .CLK(clk), .RST(1'b0), .Q(
        round_reg[586]) );
  DFF \round_reg_reg[587]  ( .D(N605), .CLK(clk), .RST(1'b0), .Q(
        round_reg[587]) );
  DFF \round_reg_reg[588]  ( .D(N606), .CLK(clk), .RST(1'b0), .Q(
        round_reg[588]) );
  DFF \round_reg_reg[589]  ( .D(N607), .CLK(clk), .RST(1'b0), .Q(
        round_reg[589]) );
  DFF \round_reg_reg[590]  ( .D(N608), .CLK(clk), .RST(1'b0), .Q(
        round_reg[590]) );
  DFF \round_reg_reg[591]  ( .D(N609), .CLK(clk), .RST(1'b0), .Q(
        round_reg[591]) );
  DFF \round_reg_reg[592]  ( .D(N610), .CLK(clk), .RST(1'b0), .Q(
        round_reg[592]) );
  DFF \round_reg_reg[593]  ( .D(N611), .CLK(clk), .RST(1'b0), .Q(
        round_reg[593]) );
  DFF \round_reg_reg[594]  ( .D(N612), .CLK(clk), .RST(1'b0), .Q(
        round_reg[594]) );
  DFF \round_reg_reg[595]  ( .D(N613), .CLK(clk), .RST(1'b0), .Q(
        round_reg[595]) );
  DFF \round_reg_reg[596]  ( .D(N614), .CLK(clk), .RST(1'b0), .Q(
        round_reg[596]) );
  DFF \round_reg_reg[597]  ( .D(N615), .CLK(clk), .RST(1'b0), .Q(
        round_reg[597]) );
  DFF \round_reg_reg[598]  ( .D(N616), .CLK(clk), .RST(1'b0), .Q(
        round_reg[598]) );
  DFF \round_reg_reg[599]  ( .D(N617), .CLK(clk), .RST(1'b0), .Q(
        round_reg[599]) );
  DFF \round_reg_reg[600]  ( .D(N618), .CLK(clk), .RST(1'b0), .Q(
        round_reg[600]) );
  DFF \round_reg_reg[601]  ( .D(N619), .CLK(clk), .RST(1'b0), .Q(
        round_reg[601]) );
  DFF \round_reg_reg[602]  ( .D(N620), .CLK(clk), .RST(1'b0), .Q(
        round_reg[602]) );
  DFF \round_reg_reg[603]  ( .D(N621), .CLK(clk), .RST(1'b0), .Q(
        round_reg[603]) );
  DFF \round_reg_reg[604]  ( .D(N622), .CLK(clk), .RST(1'b0), .Q(
        round_reg[604]) );
  DFF \round_reg_reg[605]  ( .D(N623), .CLK(clk), .RST(1'b0), .Q(
        round_reg[605]) );
  DFF \round_reg_reg[606]  ( .D(N624), .CLK(clk), .RST(1'b0), .Q(
        round_reg[606]) );
  DFF \round_reg_reg[607]  ( .D(N625), .CLK(clk), .RST(1'b0), .Q(
        round_reg[607]) );
  DFF \round_reg_reg[608]  ( .D(N626), .CLK(clk), .RST(1'b0), .Q(
        round_reg[608]) );
  DFF \round_reg_reg[609]  ( .D(N627), .CLK(clk), .RST(1'b0), .Q(
        round_reg[609]) );
  DFF \round_reg_reg[610]  ( .D(N628), .CLK(clk), .RST(1'b0), .Q(
        round_reg[610]) );
  DFF \round_reg_reg[611]  ( .D(N629), .CLK(clk), .RST(1'b0), .Q(
        round_reg[611]) );
  DFF \round_reg_reg[612]  ( .D(N630), .CLK(clk), .RST(1'b0), .Q(
        round_reg[612]) );
  DFF \round_reg_reg[613]  ( .D(N631), .CLK(clk), .RST(1'b0), .Q(
        round_reg[613]) );
  DFF \round_reg_reg[614]  ( .D(N632), .CLK(clk), .RST(1'b0), .Q(
        round_reg[614]) );
  DFF \round_reg_reg[615]  ( .D(N633), .CLK(clk), .RST(1'b0), .Q(
        round_reg[615]) );
  DFF \round_reg_reg[616]  ( .D(N634), .CLK(clk), .RST(1'b0), .Q(
        round_reg[616]) );
  DFF \round_reg_reg[617]  ( .D(N635), .CLK(clk), .RST(1'b0), .Q(
        round_reg[617]) );
  DFF \round_reg_reg[618]  ( .D(N636), .CLK(clk), .RST(1'b0), .Q(
        round_reg[618]) );
  DFF \round_reg_reg[619]  ( .D(N637), .CLK(clk), .RST(1'b0), .Q(
        round_reg[619]) );
  DFF \round_reg_reg[620]  ( .D(N638), .CLK(clk), .RST(1'b0), .Q(
        round_reg[620]) );
  DFF \round_reg_reg[621]  ( .D(N639), .CLK(clk), .RST(1'b0), .Q(
        round_reg[621]) );
  DFF \round_reg_reg[622]  ( .D(N640), .CLK(clk), .RST(1'b0), .Q(
        round_reg[622]) );
  DFF \round_reg_reg[623]  ( .D(N641), .CLK(clk), .RST(1'b0), .Q(
        round_reg[623]) );
  DFF \round_reg_reg[624]  ( .D(N642), .CLK(clk), .RST(1'b0), .Q(
        round_reg[624]) );
  DFF \round_reg_reg[625]  ( .D(N643), .CLK(clk), .RST(1'b0), .Q(
        round_reg[625]) );
  DFF \round_reg_reg[626]  ( .D(N644), .CLK(clk), .RST(1'b0), .Q(
        round_reg[626]) );
  DFF \round_reg_reg[627]  ( .D(N645), .CLK(clk), .RST(1'b0), .Q(
        round_reg[627]) );
  DFF \round_reg_reg[628]  ( .D(N646), .CLK(clk), .RST(1'b0), .Q(
        round_reg[628]) );
  DFF \round_reg_reg[629]  ( .D(N647), .CLK(clk), .RST(1'b0), .Q(
        round_reg[629]) );
  DFF \round_reg_reg[630]  ( .D(N648), .CLK(clk), .RST(1'b0), .Q(
        round_reg[630]) );
  DFF \round_reg_reg[631]  ( .D(N649), .CLK(clk), .RST(1'b0), .Q(
        round_reg[631]) );
  DFF \round_reg_reg[632]  ( .D(N650), .CLK(clk), .RST(1'b0), .Q(
        round_reg[632]) );
  DFF \round_reg_reg[633]  ( .D(N651), .CLK(clk), .RST(1'b0), .Q(
        round_reg[633]) );
  DFF \round_reg_reg[634]  ( .D(N652), .CLK(clk), .RST(1'b0), .Q(
        round_reg[634]) );
  DFF \round_reg_reg[635]  ( .D(N653), .CLK(clk), .RST(1'b0), .Q(
        round_reg[635]) );
  DFF \round_reg_reg[636]  ( .D(N654), .CLK(clk), .RST(1'b0), .Q(
        round_reg[636]) );
  DFF \round_reg_reg[637]  ( .D(N655), .CLK(clk), .RST(1'b0), .Q(
        round_reg[637]) );
  DFF \round_reg_reg[638]  ( .D(N656), .CLK(clk), .RST(1'b0), .Q(
        round_reg[638]) );
  DFF \round_reg_reg[639]  ( .D(N657), .CLK(clk), .RST(1'b0), .Q(
        round_reg[639]) );
  DFF \round_reg_reg[640]  ( .D(N658), .CLK(clk), .RST(1'b0), .Q(
        round_reg[640]) );
  DFF \round_reg_reg[641]  ( .D(N659), .CLK(clk), .RST(1'b0), .Q(
        round_reg[641]) );
  DFF \round_reg_reg[642]  ( .D(N660), .CLK(clk), .RST(1'b0), .Q(
        round_reg[642]) );
  DFF \round_reg_reg[643]  ( .D(N661), .CLK(clk), .RST(1'b0), .Q(
        round_reg[643]) );
  DFF \round_reg_reg[644]  ( .D(N662), .CLK(clk), .RST(1'b0), .Q(
        round_reg[644]) );
  DFF \round_reg_reg[645]  ( .D(N663), .CLK(clk), .RST(1'b0), .Q(
        round_reg[645]) );
  DFF \round_reg_reg[646]  ( .D(N664), .CLK(clk), .RST(1'b0), .Q(
        round_reg[646]) );
  DFF \round_reg_reg[647]  ( .D(N665), .CLK(clk), .RST(1'b0), .Q(
        round_reg[647]) );
  DFF \round_reg_reg[648]  ( .D(N666), .CLK(clk), .RST(1'b0), .Q(
        round_reg[648]) );
  DFF \round_reg_reg[649]  ( .D(N667), .CLK(clk), .RST(1'b0), .Q(
        round_reg[649]) );
  DFF \round_reg_reg[650]  ( .D(N668), .CLK(clk), .RST(1'b0), .Q(
        round_reg[650]) );
  DFF \round_reg_reg[651]  ( .D(N669), .CLK(clk), .RST(1'b0), .Q(
        round_reg[651]) );
  DFF \round_reg_reg[652]  ( .D(N670), .CLK(clk), .RST(1'b0), .Q(
        round_reg[652]) );
  DFF \round_reg_reg[653]  ( .D(N671), .CLK(clk), .RST(1'b0), .Q(
        round_reg[653]) );
  DFF \round_reg_reg[654]  ( .D(N672), .CLK(clk), .RST(1'b0), .Q(
        round_reg[654]) );
  DFF \round_reg_reg[655]  ( .D(N673), .CLK(clk), .RST(1'b0), .Q(
        round_reg[655]) );
  DFF \round_reg_reg[656]  ( .D(N674), .CLK(clk), .RST(1'b0), .Q(
        round_reg[656]) );
  DFF \round_reg_reg[657]  ( .D(N675), .CLK(clk), .RST(1'b0), .Q(
        round_reg[657]) );
  DFF \round_reg_reg[658]  ( .D(N676), .CLK(clk), .RST(1'b0), .Q(
        round_reg[658]) );
  DFF \round_reg_reg[659]  ( .D(N677), .CLK(clk), .RST(1'b0), .Q(
        round_reg[659]) );
  DFF \round_reg_reg[660]  ( .D(N678), .CLK(clk), .RST(1'b0), .Q(
        round_reg[660]) );
  DFF \round_reg_reg[661]  ( .D(N679), .CLK(clk), .RST(1'b0), .Q(
        round_reg[661]) );
  DFF \round_reg_reg[662]  ( .D(N680), .CLK(clk), .RST(1'b0), .Q(
        round_reg[662]) );
  DFF \round_reg_reg[663]  ( .D(N681), .CLK(clk), .RST(1'b0), .Q(
        round_reg[663]) );
  DFF \round_reg_reg[664]  ( .D(N682), .CLK(clk), .RST(1'b0), .Q(
        round_reg[664]) );
  DFF \round_reg_reg[665]  ( .D(N683), .CLK(clk), .RST(1'b0), .Q(
        round_reg[665]) );
  DFF \round_reg_reg[666]  ( .D(N684), .CLK(clk), .RST(1'b0), .Q(
        round_reg[666]) );
  DFF \round_reg_reg[667]  ( .D(N685), .CLK(clk), .RST(1'b0), .Q(
        round_reg[667]) );
  DFF \round_reg_reg[668]  ( .D(N686), .CLK(clk), .RST(1'b0), .Q(
        round_reg[668]) );
  DFF \round_reg_reg[669]  ( .D(N687), .CLK(clk), .RST(1'b0), .Q(
        round_reg[669]) );
  DFF \round_reg_reg[670]  ( .D(N688), .CLK(clk), .RST(1'b0), .Q(
        round_reg[670]) );
  DFF \round_reg_reg[671]  ( .D(N689), .CLK(clk), .RST(1'b0), .Q(
        round_reg[671]) );
  DFF \round_reg_reg[672]  ( .D(N690), .CLK(clk), .RST(1'b0), .Q(
        round_reg[672]) );
  DFF \round_reg_reg[673]  ( .D(N691), .CLK(clk), .RST(1'b0), .Q(
        round_reg[673]) );
  DFF \round_reg_reg[674]  ( .D(N692), .CLK(clk), .RST(1'b0), .Q(
        round_reg[674]) );
  DFF \round_reg_reg[675]  ( .D(N693), .CLK(clk), .RST(1'b0), .Q(
        round_reg[675]) );
  DFF \round_reg_reg[676]  ( .D(N694), .CLK(clk), .RST(1'b0), .Q(
        round_reg[676]) );
  DFF \round_reg_reg[677]  ( .D(N695), .CLK(clk), .RST(1'b0), .Q(
        round_reg[677]) );
  DFF \round_reg_reg[678]  ( .D(N696), .CLK(clk), .RST(1'b0), .Q(
        round_reg[678]) );
  DFF \round_reg_reg[679]  ( .D(N697), .CLK(clk), .RST(1'b0), .Q(
        round_reg[679]) );
  DFF \round_reg_reg[680]  ( .D(N698), .CLK(clk), .RST(1'b0), .Q(
        round_reg[680]) );
  DFF \round_reg_reg[681]  ( .D(N699), .CLK(clk), .RST(1'b0), .Q(
        round_reg[681]) );
  DFF \round_reg_reg[682]  ( .D(N700), .CLK(clk), .RST(1'b0), .Q(
        round_reg[682]) );
  DFF \round_reg_reg[683]  ( .D(N701), .CLK(clk), .RST(1'b0), .Q(
        round_reg[683]) );
  DFF \round_reg_reg[684]  ( .D(N702), .CLK(clk), .RST(1'b0), .Q(
        round_reg[684]) );
  DFF \round_reg_reg[685]  ( .D(N703), .CLK(clk), .RST(1'b0), .Q(
        round_reg[685]) );
  DFF \round_reg_reg[686]  ( .D(N704), .CLK(clk), .RST(1'b0), .Q(
        round_reg[686]) );
  DFF \round_reg_reg[687]  ( .D(N705), .CLK(clk), .RST(1'b0), .Q(
        round_reg[687]) );
  DFF \round_reg_reg[688]  ( .D(N706), .CLK(clk), .RST(1'b0), .Q(
        round_reg[688]) );
  DFF \round_reg_reg[689]  ( .D(N707), .CLK(clk), .RST(1'b0), .Q(
        round_reg[689]) );
  DFF \round_reg_reg[690]  ( .D(N708), .CLK(clk), .RST(1'b0), .Q(
        round_reg[690]) );
  DFF \round_reg_reg[691]  ( .D(N709), .CLK(clk), .RST(1'b0), .Q(
        round_reg[691]) );
  DFF \round_reg_reg[692]  ( .D(N710), .CLK(clk), .RST(1'b0), .Q(
        round_reg[692]) );
  DFF \round_reg_reg[693]  ( .D(N711), .CLK(clk), .RST(1'b0), .Q(
        round_reg[693]) );
  DFF \round_reg_reg[694]  ( .D(N712), .CLK(clk), .RST(1'b0), .Q(
        round_reg[694]) );
  DFF \round_reg_reg[695]  ( .D(N713), .CLK(clk), .RST(1'b0), .Q(
        round_reg[695]) );
  DFF \round_reg_reg[696]  ( .D(N714), .CLK(clk), .RST(1'b0), .Q(
        round_reg[696]) );
  DFF \round_reg_reg[697]  ( .D(N715), .CLK(clk), .RST(1'b0), .Q(
        round_reg[697]) );
  DFF \round_reg_reg[698]  ( .D(N716), .CLK(clk), .RST(1'b0), .Q(
        round_reg[698]) );
  DFF \round_reg_reg[699]  ( .D(N717), .CLK(clk), .RST(1'b0), .Q(
        round_reg[699]) );
  DFF \round_reg_reg[700]  ( .D(N718), .CLK(clk), .RST(1'b0), .Q(
        round_reg[700]) );
  DFF \round_reg_reg[701]  ( .D(N719), .CLK(clk), .RST(1'b0), .Q(
        round_reg[701]) );
  DFF \round_reg_reg[702]  ( .D(N720), .CLK(clk), .RST(1'b0), .Q(
        round_reg[702]) );
  DFF \round_reg_reg[703]  ( .D(N721), .CLK(clk), .RST(1'b0), .Q(
        round_reg[703]) );
  DFF \round_reg_reg[704]  ( .D(N722), .CLK(clk), .RST(1'b0), .Q(
        round_reg[704]) );
  DFF \round_reg_reg[705]  ( .D(N723), .CLK(clk), .RST(1'b0), .Q(
        round_reg[705]) );
  DFF \round_reg_reg[706]  ( .D(N724), .CLK(clk), .RST(1'b0), .Q(
        round_reg[706]) );
  DFF \round_reg_reg[707]  ( .D(N725), .CLK(clk), .RST(1'b0), .Q(
        round_reg[707]) );
  DFF \round_reg_reg[708]  ( .D(N726), .CLK(clk), .RST(1'b0), .Q(
        round_reg[708]) );
  DFF \round_reg_reg[709]  ( .D(N727), .CLK(clk), .RST(1'b0), .Q(
        round_reg[709]) );
  DFF \round_reg_reg[710]  ( .D(N728), .CLK(clk), .RST(1'b0), .Q(
        round_reg[710]) );
  DFF \round_reg_reg[711]  ( .D(N729), .CLK(clk), .RST(1'b0), .Q(
        round_reg[711]) );
  DFF \round_reg_reg[712]  ( .D(N730), .CLK(clk), .RST(1'b0), .Q(
        round_reg[712]) );
  DFF \round_reg_reg[713]  ( .D(N731), .CLK(clk), .RST(1'b0), .Q(
        round_reg[713]) );
  DFF \round_reg_reg[714]  ( .D(N732), .CLK(clk), .RST(1'b0), .Q(
        round_reg[714]) );
  DFF \round_reg_reg[715]  ( .D(N733), .CLK(clk), .RST(1'b0), .Q(
        round_reg[715]) );
  DFF \round_reg_reg[716]  ( .D(N734), .CLK(clk), .RST(1'b0), .Q(
        round_reg[716]) );
  DFF \round_reg_reg[717]  ( .D(N735), .CLK(clk), .RST(1'b0), .Q(
        round_reg[717]) );
  DFF \round_reg_reg[718]  ( .D(N736), .CLK(clk), .RST(1'b0), .Q(
        round_reg[718]) );
  DFF \round_reg_reg[719]  ( .D(N737), .CLK(clk), .RST(1'b0), .Q(
        round_reg[719]) );
  DFF \round_reg_reg[720]  ( .D(N738), .CLK(clk), .RST(1'b0), .Q(
        round_reg[720]) );
  DFF \round_reg_reg[721]  ( .D(N739), .CLK(clk), .RST(1'b0), .Q(
        round_reg[721]) );
  DFF \round_reg_reg[722]  ( .D(N740), .CLK(clk), .RST(1'b0), .Q(
        round_reg[722]) );
  DFF \round_reg_reg[723]  ( .D(N741), .CLK(clk), .RST(1'b0), .Q(
        round_reg[723]) );
  DFF \round_reg_reg[724]  ( .D(N742), .CLK(clk), .RST(1'b0), .Q(
        round_reg[724]) );
  DFF \round_reg_reg[725]  ( .D(N743), .CLK(clk), .RST(1'b0), .Q(
        round_reg[725]) );
  DFF \round_reg_reg[726]  ( .D(N744), .CLK(clk), .RST(1'b0), .Q(
        round_reg[726]) );
  DFF \round_reg_reg[727]  ( .D(N745), .CLK(clk), .RST(1'b0), .Q(
        round_reg[727]) );
  DFF \round_reg_reg[728]  ( .D(N746), .CLK(clk), .RST(1'b0), .Q(
        round_reg[728]) );
  DFF \round_reg_reg[729]  ( .D(N747), .CLK(clk), .RST(1'b0), .Q(
        round_reg[729]) );
  DFF \round_reg_reg[730]  ( .D(N748), .CLK(clk), .RST(1'b0), .Q(
        round_reg[730]) );
  DFF \round_reg_reg[731]  ( .D(N749), .CLK(clk), .RST(1'b0), .Q(
        round_reg[731]) );
  DFF \round_reg_reg[732]  ( .D(N750), .CLK(clk), .RST(1'b0), .Q(
        round_reg[732]) );
  DFF \round_reg_reg[733]  ( .D(N751), .CLK(clk), .RST(1'b0), .Q(
        round_reg[733]) );
  DFF \round_reg_reg[734]  ( .D(N752), .CLK(clk), .RST(1'b0), .Q(
        round_reg[734]) );
  DFF \round_reg_reg[735]  ( .D(N753), .CLK(clk), .RST(1'b0), .Q(
        round_reg[735]) );
  DFF \round_reg_reg[736]  ( .D(N754), .CLK(clk), .RST(1'b0), .Q(
        round_reg[736]) );
  DFF \round_reg_reg[737]  ( .D(N755), .CLK(clk), .RST(1'b0), .Q(
        round_reg[737]) );
  DFF \round_reg_reg[738]  ( .D(N756), .CLK(clk), .RST(1'b0), .Q(
        round_reg[738]) );
  DFF \round_reg_reg[739]  ( .D(N757), .CLK(clk), .RST(1'b0), .Q(
        round_reg[739]) );
  DFF \round_reg_reg[740]  ( .D(N758), .CLK(clk), .RST(1'b0), .Q(
        round_reg[740]) );
  DFF \round_reg_reg[741]  ( .D(N759), .CLK(clk), .RST(1'b0), .Q(
        round_reg[741]) );
  DFF \round_reg_reg[742]  ( .D(N760), .CLK(clk), .RST(1'b0), .Q(
        round_reg[742]) );
  DFF \round_reg_reg[743]  ( .D(N761), .CLK(clk), .RST(1'b0), .Q(
        round_reg[743]) );
  DFF \round_reg_reg[744]  ( .D(N762), .CLK(clk), .RST(1'b0), .Q(
        round_reg[744]) );
  DFF \round_reg_reg[745]  ( .D(N763), .CLK(clk), .RST(1'b0), .Q(
        round_reg[745]) );
  DFF \round_reg_reg[746]  ( .D(N764), .CLK(clk), .RST(1'b0), .Q(
        round_reg[746]) );
  DFF \round_reg_reg[747]  ( .D(N765), .CLK(clk), .RST(1'b0), .Q(
        round_reg[747]) );
  DFF \round_reg_reg[748]  ( .D(N766), .CLK(clk), .RST(1'b0), .Q(
        round_reg[748]) );
  DFF \round_reg_reg[749]  ( .D(N767), .CLK(clk), .RST(1'b0), .Q(
        round_reg[749]) );
  DFF \round_reg_reg[750]  ( .D(N768), .CLK(clk), .RST(1'b0), .Q(
        round_reg[750]) );
  DFF \round_reg_reg[751]  ( .D(N769), .CLK(clk), .RST(1'b0), .Q(
        round_reg[751]) );
  DFF \round_reg_reg[752]  ( .D(N770), .CLK(clk), .RST(1'b0), .Q(
        round_reg[752]) );
  DFF \round_reg_reg[753]  ( .D(N771), .CLK(clk), .RST(1'b0), .Q(
        round_reg[753]) );
  DFF \round_reg_reg[754]  ( .D(N772), .CLK(clk), .RST(1'b0), .Q(
        round_reg[754]) );
  DFF \round_reg_reg[755]  ( .D(N773), .CLK(clk), .RST(1'b0), .Q(
        round_reg[755]) );
  DFF \round_reg_reg[756]  ( .D(N774), .CLK(clk), .RST(1'b0), .Q(
        round_reg[756]) );
  DFF \round_reg_reg[757]  ( .D(N775), .CLK(clk), .RST(1'b0), .Q(
        round_reg[757]) );
  DFF \round_reg_reg[758]  ( .D(N776), .CLK(clk), .RST(1'b0), .Q(
        round_reg[758]) );
  DFF \round_reg_reg[759]  ( .D(N777), .CLK(clk), .RST(1'b0), .Q(
        round_reg[759]) );
  DFF \round_reg_reg[760]  ( .D(N778), .CLK(clk), .RST(1'b0), .Q(
        round_reg[760]) );
  DFF \round_reg_reg[761]  ( .D(N779), .CLK(clk), .RST(1'b0), .Q(
        round_reg[761]) );
  DFF \round_reg_reg[762]  ( .D(N780), .CLK(clk), .RST(1'b0), .Q(
        round_reg[762]) );
  DFF \round_reg_reg[763]  ( .D(N781), .CLK(clk), .RST(1'b0), .Q(
        round_reg[763]) );
  DFF \round_reg_reg[764]  ( .D(N782), .CLK(clk), .RST(1'b0), .Q(
        round_reg[764]) );
  DFF \round_reg_reg[765]  ( .D(N783), .CLK(clk), .RST(1'b0), .Q(
        round_reg[765]) );
  DFF \round_reg_reg[766]  ( .D(N784), .CLK(clk), .RST(1'b0), .Q(
        round_reg[766]) );
  DFF \round_reg_reg[767]  ( .D(N785), .CLK(clk), .RST(1'b0), .Q(
        round_reg[767]) );
  DFF \round_reg_reg[768]  ( .D(N786), .CLK(clk), .RST(1'b0), .Q(
        round_reg[768]) );
  DFF \round_reg_reg[769]  ( .D(N787), .CLK(clk), .RST(1'b0), .Q(
        round_reg[769]) );
  DFF \round_reg_reg[770]  ( .D(N788), .CLK(clk), .RST(1'b0), .Q(
        round_reg[770]) );
  DFF \round_reg_reg[771]  ( .D(N789), .CLK(clk), .RST(1'b0), .Q(
        round_reg[771]) );
  DFF \round_reg_reg[772]  ( .D(N790), .CLK(clk), .RST(1'b0), .Q(
        round_reg[772]) );
  DFF \round_reg_reg[773]  ( .D(N791), .CLK(clk), .RST(1'b0), .Q(
        round_reg[773]) );
  DFF \round_reg_reg[774]  ( .D(N792), .CLK(clk), .RST(1'b0), .Q(
        round_reg[774]) );
  DFF \round_reg_reg[775]  ( .D(N793), .CLK(clk), .RST(1'b0), .Q(
        round_reg[775]) );
  DFF \round_reg_reg[776]  ( .D(N794), .CLK(clk), .RST(1'b0), .Q(
        round_reg[776]) );
  DFF \round_reg_reg[777]  ( .D(N795), .CLK(clk), .RST(1'b0), .Q(
        round_reg[777]) );
  DFF \round_reg_reg[778]  ( .D(N796), .CLK(clk), .RST(1'b0), .Q(
        round_reg[778]) );
  DFF \round_reg_reg[779]  ( .D(N797), .CLK(clk), .RST(1'b0), .Q(
        round_reg[779]) );
  DFF \round_reg_reg[780]  ( .D(N798), .CLK(clk), .RST(1'b0), .Q(
        round_reg[780]) );
  DFF \round_reg_reg[781]  ( .D(N799), .CLK(clk), .RST(1'b0), .Q(
        round_reg[781]) );
  DFF \round_reg_reg[782]  ( .D(N800), .CLK(clk), .RST(1'b0), .Q(
        round_reg[782]) );
  DFF \round_reg_reg[783]  ( .D(N801), .CLK(clk), .RST(1'b0), .Q(
        round_reg[783]) );
  DFF \round_reg_reg[784]  ( .D(N802), .CLK(clk), .RST(1'b0), .Q(
        round_reg[784]) );
  DFF \round_reg_reg[785]  ( .D(N803), .CLK(clk), .RST(1'b0), .Q(
        round_reg[785]) );
  DFF \round_reg_reg[786]  ( .D(N804), .CLK(clk), .RST(1'b0), .Q(
        round_reg[786]) );
  DFF \round_reg_reg[787]  ( .D(N805), .CLK(clk), .RST(1'b0), .Q(
        round_reg[787]) );
  DFF \round_reg_reg[788]  ( .D(N806), .CLK(clk), .RST(1'b0), .Q(
        round_reg[788]) );
  DFF \round_reg_reg[789]  ( .D(N807), .CLK(clk), .RST(1'b0), .Q(
        round_reg[789]) );
  DFF \round_reg_reg[790]  ( .D(N808), .CLK(clk), .RST(1'b0), .Q(
        round_reg[790]) );
  DFF \round_reg_reg[791]  ( .D(N809), .CLK(clk), .RST(1'b0), .Q(
        round_reg[791]) );
  DFF \round_reg_reg[792]  ( .D(N810), .CLK(clk), .RST(1'b0), .Q(
        round_reg[792]) );
  DFF \round_reg_reg[793]  ( .D(N811), .CLK(clk), .RST(1'b0), .Q(
        round_reg[793]) );
  DFF \round_reg_reg[794]  ( .D(N812), .CLK(clk), .RST(1'b0), .Q(
        round_reg[794]) );
  DFF \round_reg_reg[795]  ( .D(N813), .CLK(clk), .RST(1'b0), .Q(
        round_reg[795]) );
  DFF \round_reg_reg[796]  ( .D(N814), .CLK(clk), .RST(1'b0), .Q(
        round_reg[796]) );
  DFF \round_reg_reg[797]  ( .D(N815), .CLK(clk), .RST(1'b0), .Q(
        round_reg[797]) );
  DFF \round_reg_reg[798]  ( .D(N816), .CLK(clk), .RST(1'b0), .Q(
        round_reg[798]) );
  DFF \round_reg_reg[799]  ( .D(N817), .CLK(clk), .RST(1'b0), .Q(
        round_reg[799]) );
  DFF \round_reg_reg[800]  ( .D(N818), .CLK(clk), .RST(1'b0), .Q(
        round_reg[800]) );
  DFF \round_reg_reg[801]  ( .D(N819), .CLK(clk), .RST(1'b0), .Q(
        round_reg[801]) );
  DFF \round_reg_reg[802]  ( .D(N820), .CLK(clk), .RST(1'b0), .Q(
        round_reg[802]) );
  DFF \round_reg_reg[803]  ( .D(N821), .CLK(clk), .RST(1'b0), .Q(
        round_reg[803]) );
  DFF \round_reg_reg[804]  ( .D(N822), .CLK(clk), .RST(1'b0), .Q(
        round_reg[804]) );
  DFF \round_reg_reg[805]  ( .D(N823), .CLK(clk), .RST(1'b0), .Q(
        round_reg[805]) );
  DFF \round_reg_reg[806]  ( .D(N824), .CLK(clk), .RST(1'b0), .Q(
        round_reg[806]) );
  DFF \round_reg_reg[807]  ( .D(N825), .CLK(clk), .RST(1'b0), .Q(
        round_reg[807]) );
  DFF \round_reg_reg[808]  ( .D(N826), .CLK(clk), .RST(1'b0), .Q(
        round_reg[808]) );
  DFF \round_reg_reg[809]  ( .D(N827), .CLK(clk), .RST(1'b0), .Q(
        round_reg[809]) );
  DFF \round_reg_reg[810]  ( .D(N828), .CLK(clk), .RST(1'b0), .Q(
        round_reg[810]) );
  DFF \round_reg_reg[811]  ( .D(N829), .CLK(clk), .RST(1'b0), .Q(
        round_reg[811]) );
  DFF \round_reg_reg[812]  ( .D(N830), .CLK(clk), .RST(1'b0), .Q(
        round_reg[812]) );
  DFF \round_reg_reg[813]  ( .D(N831), .CLK(clk), .RST(1'b0), .Q(
        round_reg[813]) );
  DFF \round_reg_reg[814]  ( .D(N832), .CLK(clk), .RST(1'b0), .Q(
        round_reg[814]) );
  DFF \round_reg_reg[815]  ( .D(N833), .CLK(clk), .RST(1'b0), .Q(
        round_reg[815]) );
  DFF \round_reg_reg[816]  ( .D(N834), .CLK(clk), .RST(1'b0), .Q(
        round_reg[816]) );
  DFF \round_reg_reg[817]  ( .D(N835), .CLK(clk), .RST(1'b0), .Q(
        round_reg[817]) );
  DFF \round_reg_reg[818]  ( .D(N836), .CLK(clk), .RST(1'b0), .Q(
        round_reg[818]) );
  DFF \round_reg_reg[819]  ( .D(N837), .CLK(clk), .RST(1'b0), .Q(
        round_reg[819]) );
  DFF \round_reg_reg[820]  ( .D(N838), .CLK(clk), .RST(1'b0), .Q(
        round_reg[820]) );
  DFF \round_reg_reg[821]  ( .D(N839), .CLK(clk), .RST(1'b0), .Q(
        round_reg[821]) );
  DFF \round_reg_reg[822]  ( .D(N840), .CLK(clk), .RST(1'b0), .Q(
        round_reg[822]) );
  DFF \round_reg_reg[823]  ( .D(N841), .CLK(clk), .RST(1'b0), .Q(
        round_reg[823]) );
  DFF \round_reg_reg[824]  ( .D(N842), .CLK(clk), .RST(1'b0), .Q(
        round_reg[824]) );
  DFF \round_reg_reg[825]  ( .D(N843), .CLK(clk), .RST(1'b0), .Q(
        round_reg[825]) );
  DFF \round_reg_reg[826]  ( .D(N844), .CLK(clk), .RST(1'b0), .Q(
        round_reg[826]) );
  DFF \round_reg_reg[827]  ( .D(N845), .CLK(clk), .RST(1'b0), .Q(
        round_reg[827]) );
  DFF \round_reg_reg[828]  ( .D(N846), .CLK(clk), .RST(1'b0), .Q(
        round_reg[828]) );
  DFF \round_reg_reg[829]  ( .D(N847), .CLK(clk), .RST(1'b0), .Q(
        round_reg[829]) );
  DFF \round_reg_reg[830]  ( .D(N848), .CLK(clk), .RST(1'b0), .Q(
        round_reg[830]) );
  DFF \round_reg_reg[831]  ( .D(N849), .CLK(clk), .RST(1'b0), .Q(
        round_reg[831]) );
  DFF \round_reg_reg[832]  ( .D(N850), .CLK(clk), .RST(1'b0), .Q(
        round_reg[832]) );
  DFF \round_reg_reg[833]  ( .D(N851), .CLK(clk), .RST(1'b0), .Q(
        round_reg[833]) );
  DFF \round_reg_reg[834]  ( .D(N852), .CLK(clk), .RST(1'b0), .Q(
        round_reg[834]) );
  DFF \round_reg_reg[835]  ( .D(N853), .CLK(clk), .RST(1'b0), .Q(
        round_reg[835]) );
  DFF \round_reg_reg[836]  ( .D(N854), .CLK(clk), .RST(1'b0), .Q(
        round_reg[836]) );
  DFF \round_reg_reg[837]  ( .D(N855), .CLK(clk), .RST(1'b0), .Q(
        round_reg[837]) );
  DFF \round_reg_reg[838]  ( .D(N856), .CLK(clk), .RST(1'b0), .Q(
        round_reg[838]) );
  DFF \round_reg_reg[839]  ( .D(N857), .CLK(clk), .RST(1'b0), .Q(
        round_reg[839]) );
  DFF \round_reg_reg[840]  ( .D(N858), .CLK(clk), .RST(1'b0), .Q(
        round_reg[840]) );
  DFF \round_reg_reg[841]  ( .D(N859), .CLK(clk), .RST(1'b0), .Q(
        round_reg[841]) );
  DFF \round_reg_reg[842]  ( .D(N860), .CLK(clk), .RST(1'b0), .Q(
        round_reg[842]) );
  DFF \round_reg_reg[843]  ( .D(N861), .CLK(clk), .RST(1'b0), .Q(
        round_reg[843]) );
  DFF \round_reg_reg[844]  ( .D(N862), .CLK(clk), .RST(1'b0), .Q(
        round_reg[844]) );
  DFF \round_reg_reg[845]  ( .D(N863), .CLK(clk), .RST(1'b0), .Q(
        round_reg[845]) );
  DFF \round_reg_reg[846]  ( .D(N864), .CLK(clk), .RST(1'b0), .Q(
        round_reg[846]) );
  DFF \round_reg_reg[847]  ( .D(N865), .CLK(clk), .RST(1'b0), .Q(
        round_reg[847]) );
  DFF \round_reg_reg[848]  ( .D(N866), .CLK(clk), .RST(1'b0), .Q(
        round_reg[848]) );
  DFF \round_reg_reg[849]  ( .D(N867), .CLK(clk), .RST(1'b0), .Q(
        round_reg[849]) );
  DFF \round_reg_reg[850]  ( .D(N868), .CLK(clk), .RST(1'b0), .Q(
        round_reg[850]) );
  DFF \round_reg_reg[851]  ( .D(N869), .CLK(clk), .RST(1'b0), .Q(
        round_reg[851]) );
  DFF \round_reg_reg[852]  ( .D(N870), .CLK(clk), .RST(1'b0), .Q(
        round_reg[852]) );
  DFF \round_reg_reg[853]  ( .D(N871), .CLK(clk), .RST(1'b0), .Q(
        round_reg[853]) );
  DFF \round_reg_reg[854]  ( .D(N872), .CLK(clk), .RST(1'b0), .Q(
        round_reg[854]) );
  DFF \round_reg_reg[855]  ( .D(N873), .CLK(clk), .RST(1'b0), .Q(
        round_reg[855]) );
  DFF \round_reg_reg[856]  ( .D(N874), .CLK(clk), .RST(1'b0), .Q(
        round_reg[856]) );
  DFF \round_reg_reg[857]  ( .D(N875), .CLK(clk), .RST(1'b0), .Q(
        round_reg[857]) );
  DFF \round_reg_reg[858]  ( .D(N876), .CLK(clk), .RST(1'b0), .Q(
        round_reg[858]) );
  DFF \round_reg_reg[859]  ( .D(N877), .CLK(clk), .RST(1'b0), .Q(
        round_reg[859]) );
  DFF \round_reg_reg[860]  ( .D(N878), .CLK(clk), .RST(1'b0), .Q(
        round_reg[860]) );
  DFF \round_reg_reg[861]  ( .D(N879), .CLK(clk), .RST(1'b0), .Q(
        round_reg[861]) );
  DFF \round_reg_reg[862]  ( .D(N880), .CLK(clk), .RST(1'b0), .Q(
        round_reg[862]) );
  DFF \round_reg_reg[863]  ( .D(N881), .CLK(clk), .RST(1'b0), .Q(
        round_reg[863]) );
  DFF \round_reg_reg[864]  ( .D(N882), .CLK(clk), .RST(1'b0), .Q(
        round_reg[864]) );
  DFF \round_reg_reg[865]  ( .D(N883), .CLK(clk), .RST(1'b0), .Q(
        round_reg[865]) );
  DFF \round_reg_reg[866]  ( .D(N884), .CLK(clk), .RST(1'b0), .Q(
        round_reg[866]) );
  DFF \round_reg_reg[867]  ( .D(N885), .CLK(clk), .RST(1'b0), .Q(
        round_reg[867]) );
  DFF \round_reg_reg[868]  ( .D(N886), .CLK(clk), .RST(1'b0), .Q(
        round_reg[868]) );
  DFF \round_reg_reg[869]  ( .D(N887), .CLK(clk), .RST(1'b0), .Q(
        round_reg[869]) );
  DFF \round_reg_reg[870]  ( .D(N888), .CLK(clk), .RST(1'b0), .Q(
        round_reg[870]) );
  DFF \round_reg_reg[871]  ( .D(N889), .CLK(clk), .RST(1'b0), .Q(
        round_reg[871]) );
  DFF \round_reg_reg[872]  ( .D(N890), .CLK(clk), .RST(1'b0), .Q(
        round_reg[872]) );
  DFF \round_reg_reg[873]  ( .D(N891), .CLK(clk), .RST(1'b0), .Q(
        round_reg[873]) );
  DFF \round_reg_reg[874]  ( .D(N892), .CLK(clk), .RST(1'b0), .Q(
        round_reg[874]) );
  DFF \round_reg_reg[875]  ( .D(N893), .CLK(clk), .RST(1'b0), .Q(
        round_reg[875]) );
  DFF \round_reg_reg[876]  ( .D(N894), .CLK(clk), .RST(1'b0), .Q(
        round_reg[876]) );
  DFF \round_reg_reg[877]  ( .D(N895), .CLK(clk), .RST(1'b0), .Q(
        round_reg[877]) );
  DFF \round_reg_reg[878]  ( .D(N896), .CLK(clk), .RST(1'b0), .Q(
        round_reg[878]) );
  DFF \round_reg_reg[879]  ( .D(N897), .CLK(clk), .RST(1'b0), .Q(
        round_reg[879]) );
  DFF \round_reg_reg[880]  ( .D(N898), .CLK(clk), .RST(1'b0), .Q(
        round_reg[880]) );
  DFF \round_reg_reg[881]  ( .D(N899), .CLK(clk), .RST(1'b0), .Q(
        round_reg[881]) );
  DFF \round_reg_reg[882]  ( .D(N900), .CLK(clk), .RST(1'b0), .Q(
        round_reg[882]) );
  DFF \round_reg_reg[883]  ( .D(N901), .CLK(clk), .RST(1'b0), .Q(
        round_reg[883]) );
  DFF \round_reg_reg[884]  ( .D(N902), .CLK(clk), .RST(1'b0), .Q(
        round_reg[884]) );
  DFF \round_reg_reg[885]  ( .D(N903), .CLK(clk), .RST(1'b0), .Q(
        round_reg[885]) );
  DFF \round_reg_reg[886]  ( .D(N904), .CLK(clk), .RST(1'b0), .Q(
        round_reg[886]) );
  DFF \round_reg_reg[887]  ( .D(N905), .CLK(clk), .RST(1'b0), .Q(
        round_reg[887]) );
  DFF \round_reg_reg[888]  ( .D(N906), .CLK(clk), .RST(1'b0), .Q(
        round_reg[888]) );
  DFF \round_reg_reg[889]  ( .D(N907), .CLK(clk), .RST(1'b0), .Q(
        round_reg[889]) );
  DFF \round_reg_reg[890]  ( .D(N908), .CLK(clk), .RST(1'b0), .Q(
        round_reg[890]) );
  DFF \round_reg_reg[891]  ( .D(N909), .CLK(clk), .RST(1'b0), .Q(
        round_reg[891]) );
  DFF \round_reg_reg[892]  ( .D(N910), .CLK(clk), .RST(1'b0), .Q(
        round_reg[892]) );
  DFF \round_reg_reg[893]  ( .D(N911), .CLK(clk), .RST(1'b0), .Q(
        round_reg[893]) );
  DFF \round_reg_reg[894]  ( .D(N912), .CLK(clk), .RST(1'b0), .Q(
        round_reg[894]) );
  DFF \round_reg_reg[895]  ( .D(N913), .CLK(clk), .RST(1'b0), .Q(
        round_reg[895]) );
  DFF \round_reg_reg[896]  ( .D(N914), .CLK(clk), .RST(1'b0), .Q(
        round_reg[896]) );
  DFF \round_reg_reg[897]  ( .D(N915), .CLK(clk), .RST(1'b0), .Q(
        round_reg[897]) );
  DFF \round_reg_reg[898]  ( .D(N916), .CLK(clk), .RST(1'b0), .Q(
        round_reg[898]) );
  DFF \round_reg_reg[899]  ( .D(N917), .CLK(clk), .RST(1'b0), .Q(
        round_reg[899]) );
  DFF \round_reg_reg[900]  ( .D(N918), .CLK(clk), .RST(1'b0), .Q(
        round_reg[900]) );
  DFF \round_reg_reg[901]  ( .D(N919), .CLK(clk), .RST(1'b0), .Q(
        round_reg[901]) );
  DFF \round_reg_reg[902]  ( .D(N920), .CLK(clk), .RST(1'b0), .Q(
        round_reg[902]) );
  DFF \round_reg_reg[903]  ( .D(N921), .CLK(clk), .RST(1'b0), .Q(
        round_reg[903]) );
  DFF \round_reg_reg[904]  ( .D(N922), .CLK(clk), .RST(1'b0), .Q(
        round_reg[904]) );
  DFF \round_reg_reg[905]  ( .D(N923), .CLK(clk), .RST(1'b0), .Q(
        round_reg[905]) );
  DFF \round_reg_reg[906]  ( .D(N924), .CLK(clk), .RST(1'b0), .Q(
        round_reg[906]) );
  DFF \round_reg_reg[907]  ( .D(N925), .CLK(clk), .RST(1'b0), .Q(
        round_reg[907]) );
  DFF \round_reg_reg[908]  ( .D(N926), .CLK(clk), .RST(1'b0), .Q(
        round_reg[908]) );
  DFF \round_reg_reg[909]  ( .D(N927), .CLK(clk), .RST(1'b0), .Q(
        round_reg[909]) );
  DFF \round_reg_reg[910]  ( .D(N928), .CLK(clk), .RST(1'b0), .Q(
        round_reg[910]) );
  DFF \round_reg_reg[911]  ( .D(N929), .CLK(clk), .RST(1'b0), .Q(
        round_reg[911]) );
  DFF \round_reg_reg[912]  ( .D(N930), .CLK(clk), .RST(1'b0), .Q(
        round_reg[912]) );
  DFF \round_reg_reg[913]  ( .D(N931), .CLK(clk), .RST(1'b0), .Q(
        round_reg[913]) );
  DFF \round_reg_reg[914]  ( .D(N932), .CLK(clk), .RST(1'b0), .Q(
        round_reg[914]) );
  DFF \round_reg_reg[915]  ( .D(N933), .CLK(clk), .RST(1'b0), .Q(
        round_reg[915]) );
  DFF \round_reg_reg[916]  ( .D(N934), .CLK(clk), .RST(1'b0), .Q(
        round_reg[916]) );
  DFF \round_reg_reg[917]  ( .D(N935), .CLK(clk), .RST(1'b0), .Q(
        round_reg[917]) );
  DFF \round_reg_reg[918]  ( .D(N936), .CLK(clk), .RST(1'b0), .Q(
        round_reg[918]) );
  DFF \round_reg_reg[919]  ( .D(N937), .CLK(clk), .RST(1'b0), .Q(
        round_reg[919]) );
  DFF \round_reg_reg[920]  ( .D(N938), .CLK(clk), .RST(1'b0), .Q(
        round_reg[920]) );
  DFF \round_reg_reg[921]  ( .D(N939), .CLK(clk), .RST(1'b0), .Q(
        round_reg[921]) );
  DFF \round_reg_reg[922]  ( .D(N940), .CLK(clk), .RST(1'b0), .Q(
        round_reg[922]) );
  DFF \round_reg_reg[923]  ( .D(N941), .CLK(clk), .RST(1'b0), .Q(
        round_reg[923]) );
  DFF \round_reg_reg[924]  ( .D(N942), .CLK(clk), .RST(1'b0), .Q(
        round_reg[924]) );
  DFF \round_reg_reg[925]  ( .D(N943), .CLK(clk), .RST(1'b0), .Q(
        round_reg[925]) );
  DFF \round_reg_reg[926]  ( .D(N944), .CLK(clk), .RST(1'b0), .Q(
        round_reg[926]) );
  DFF \round_reg_reg[927]  ( .D(N945), .CLK(clk), .RST(1'b0), .Q(
        round_reg[927]) );
  DFF \round_reg_reg[928]  ( .D(N946), .CLK(clk), .RST(1'b0), .Q(
        round_reg[928]) );
  DFF \round_reg_reg[929]  ( .D(N947), .CLK(clk), .RST(1'b0), .Q(
        round_reg[929]) );
  DFF \round_reg_reg[930]  ( .D(N948), .CLK(clk), .RST(1'b0), .Q(
        round_reg[930]) );
  DFF \round_reg_reg[931]  ( .D(N949), .CLK(clk), .RST(1'b0), .Q(
        round_reg[931]) );
  DFF \round_reg_reg[932]  ( .D(N950), .CLK(clk), .RST(1'b0), .Q(
        round_reg[932]) );
  DFF \round_reg_reg[933]  ( .D(N951), .CLK(clk), .RST(1'b0), .Q(
        round_reg[933]) );
  DFF \round_reg_reg[934]  ( .D(N952), .CLK(clk), .RST(1'b0), .Q(
        round_reg[934]) );
  DFF \round_reg_reg[935]  ( .D(N953), .CLK(clk), .RST(1'b0), .Q(
        round_reg[935]) );
  DFF \round_reg_reg[936]  ( .D(N954), .CLK(clk), .RST(1'b0), .Q(
        round_reg[936]) );
  DFF \round_reg_reg[937]  ( .D(N955), .CLK(clk), .RST(1'b0), .Q(
        round_reg[937]) );
  DFF \round_reg_reg[938]  ( .D(N956), .CLK(clk), .RST(1'b0), .Q(
        round_reg[938]) );
  DFF \round_reg_reg[939]  ( .D(N957), .CLK(clk), .RST(1'b0), .Q(
        round_reg[939]) );
  DFF \round_reg_reg[940]  ( .D(N958), .CLK(clk), .RST(1'b0), .Q(
        round_reg[940]) );
  DFF \round_reg_reg[941]  ( .D(N959), .CLK(clk), .RST(1'b0), .Q(
        round_reg[941]) );
  DFF \round_reg_reg[942]  ( .D(N960), .CLK(clk), .RST(1'b0), .Q(
        round_reg[942]) );
  DFF \round_reg_reg[943]  ( .D(N961), .CLK(clk), .RST(1'b0), .Q(
        round_reg[943]) );
  DFF \round_reg_reg[944]  ( .D(N962), .CLK(clk), .RST(1'b0), .Q(
        round_reg[944]) );
  DFF \round_reg_reg[945]  ( .D(N963), .CLK(clk), .RST(1'b0), .Q(
        round_reg[945]) );
  DFF \round_reg_reg[946]  ( .D(N964), .CLK(clk), .RST(1'b0), .Q(
        round_reg[946]) );
  DFF \round_reg_reg[947]  ( .D(N965), .CLK(clk), .RST(1'b0), .Q(
        round_reg[947]) );
  DFF \round_reg_reg[948]  ( .D(N966), .CLK(clk), .RST(1'b0), .Q(
        round_reg[948]) );
  DFF \round_reg_reg[949]  ( .D(N967), .CLK(clk), .RST(1'b0), .Q(
        round_reg[949]) );
  DFF \round_reg_reg[950]  ( .D(N968), .CLK(clk), .RST(1'b0), .Q(
        round_reg[950]) );
  DFF \round_reg_reg[951]  ( .D(N969), .CLK(clk), .RST(1'b0), .Q(
        round_reg[951]) );
  DFF \round_reg_reg[952]  ( .D(N970), .CLK(clk), .RST(1'b0), .Q(
        round_reg[952]) );
  DFF \round_reg_reg[953]  ( .D(N971), .CLK(clk), .RST(1'b0), .Q(
        round_reg[953]) );
  DFF \round_reg_reg[954]  ( .D(N972), .CLK(clk), .RST(1'b0), .Q(
        round_reg[954]) );
  DFF \round_reg_reg[955]  ( .D(N973), .CLK(clk), .RST(1'b0), .Q(
        round_reg[955]) );
  DFF \round_reg_reg[956]  ( .D(N974), .CLK(clk), .RST(1'b0), .Q(
        round_reg[956]) );
  DFF \round_reg_reg[957]  ( .D(N975), .CLK(clk), .RST(1'b0), .Q(
        round_reg[957]) );
  DFF \round_reg_reg[958]  ( .D(N976), .CLK(clk), .RST(1'b0), .Q(
        round_reg[958]) );
  DFF \round_reg_reg[959]  ( .D(N977), .CLK(clk), .RST(1'b0), .Q(
        round_reg[959]) );
  DFF \round_reg_reg[960]  ( .D(N978), .CLK(clk), .RST(1'b0), .Q(
        round_reg[960]) );
  DFF \round_reg_reg[961]  ( .D(N979), .CLK(clk), .RST(1'b0), .Q(
        round_reg[961]) );
  DFF \round_reg_reg[962]  ( .D(N980), .CLK(clk), .RST(1'b0), .Q(
        round_reg[962]) );
  DFF \round_reg_reg[963]  ( .D(N981), .CLK(clk), .RST(1'b0), .Q(
        round_reg[963]) );
  DFF \round_reg_reg[964]  ( .D(N982), .CLK(clk), .RST(1'b0), .Q(
        round_reg[964]) );
  DFF \round_reg_reg[965]  ( .D(N983), .CLK(clk), .RST(1'b0), .Q(
        round_reg[965]) );
  DFF \round_reg_reg[966]  ( .D(N984), .CLK(clk), .RST(1'b0), .Q(
        round_reg[966]) );
  DFF \round_reg_reg[967]  ( .D(N985), .CLK(clk), .RST(1'b0), .Q(
        round_reg[967]) );
  DFF \round_reg_reg[968]  ( .D(N986), .CLK(clk), .RST(1'b0), .Q(
        round_reg[968]) );
  DFF \round_reg_reg[969]  ( .D(N987), .CLK(clk), .RST(1'b0), .Q(
        round_reg[969]) );
  DFF \round_reg_reg[970]  ( .D(N988), .CLK(clk), .RST(1'b0), .Q(
        round_reg[970]) );
  DFF \round_reg_reg[971]  ( .D(N989), .CLK(clk), .RST(1'b0), .Q(
        round_reg[971]) );
  DFF \round_reg_reg[972]  ( .D(N990), .CLK(clk), .RST(1'b0), .Q(
        round_reg[972]) );
  DFF \round_reg_reg[973]  ( .D(N991), .CLK(clk), .RST(1'b0), .Q(
        round_reg[973]) );
  DFF \round_reg_reg[974]  ( .D(N992), .CLK(clk), .RST(1'b0), .Q(
        round_reg[974]) );
  DFF \round_reg_reg[975]  ( .D(N993), .CLK(clk), .RST(1'b0), .Q(
        round_reg[975]) );
  DFF \round_reg_reg[976]  ( .D(N994), .CLK(clk), .RST(1'b0), .Q(
        round_reg[976]) );
  DFF \round_reg_reg[977]  ( .D(N995), .CLK(clk), .RST(1'b0), .Q(
        round_reg[977]) );
  DFF \round_reg_reg[978]  ( .D(N996), .CLK(clk), .RST(1'b0), .Q(
        round_reg[978]) );
  DFF \round_reg_reg[979]  ( .D(N997), .CLK(clk), .RST(1'b0), .Q(
        round_reg[979]) );
  DFF \round_reg_reg[980]  ( .D(N998), .CLK(clk), .RST(1'b0), .Q(
        round_reg[980]) );
  DFF \round_reg_reg[981]  ( .D(N999), .CLK(clk), .RST(1'b0), .Q(
        round_reg[981]) );
  DFF \round_reg_reg[982]  ( .D(N1000), .CLK(clk), .RST(1'b0), .Q(
        round_reg[982]) );
  DFF \round_reg_reg[983]  ( .D(N1001), .CLK(clk), .RST(1'b0), .Q(
        round_reg[983]) );
  DFF \round_reg_reg[984]  ( .D(N1002), .CLK(clk), .RST(1'b0), .Q(
        round_reg[984]) );
  DFF \round_reg_reg[985]  ( .D(N1003), .CLK(clk), .RST(1'b0), .Q(
        round_reg[985]) );
  DFF \round_reg_reg[986]  ( .D(N1004), .CLK(clk), .RST(1'b0), .Q(
        round_reg[986]) );
  DFF \round_reg_reg[987]  ( .D(N1005), .CLK(clk), .RST(1'b0), .Q(
        round_reg[987]) );
  DFF \round_reg_reg[988]  ( .D(N1006), .CLK(clk), .RST(1'b0), .Q(
        round_reg[988]) );
  DFF \round_reg_reg[989]  ( .D(N1007), .CLK(clk), .RST(1'b0), .Q(
        round_reg[989]) );
  DFF \round_reg_reg[990]  ( .D(N1008), .CLK(clk), .RST(1'b0), .Q(
        round_reg[990]) );
  DFF \round_reg_reg[991]  ( .D(N1009), .CLK(clk), .RST(1'b0), .Q(
        round_reg[991]) );
  DFF \round_reg_reg[992]  ( .D(N1010), .CLK(clk), .RST(1'b0), .Q(
        round_reg[992]) );
  DFF \round_reg_reg[993]  ( .D(N1011), .CLK(clk), .RST(1'b0), .Q(
        round_reg[993]) );
  DFF \round_reg_reg[994]  ( .D(N1012), .CLK(clk), .RST(1'b0), .Q(
        round_reg[994]) );
  DFF \round_reg_reg[995]  ( .D(N1013), .CLK(clk), .RST(1'b0), .Q(
        round_reg[995]) );
  DFF \round_reg_reg[996]  ( .D(N1014), .CLK(clk), .RST(1'b0), .Q(
        round_reg[996]) );
  DFF \round_reg_reg[997]  ( .D(N1015), .CLK(clk), .RST(1'b0), .Q(
        round_reg[997]) );
  DFF \round_reg_reg[998]  ( .D(N1016), .CLK(clk), .RST(1'b0), .Q(
        round_reg[998]) );
  DFF \round_reg_reg[999]  ( .D(N1017), .CLK(clk), .RST(1'b0), .Q(
        round_reg[999]) );
  DFF \round_reg_reg[1000]  ( .D(N1018), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1000]) );
  DFF \round_reg_reg[1001]  ( .D(N1019), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1001]) );
  DFF \round_reg_reg[1002]  ( .D(N1020), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1002]) );
  DFF \round_reg_reg[1003]  ( .D(N1021), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1003]) );
  DFF \round_reg_reg[1004]  ( .D(N1022), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1004]) );
  DFF \round_reg_reg[1005]  ( .D(N1023), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1005]) );
  DFF \round_reg_reg[1006]  ( .D(N1024), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1006]) );
  DFF \round_reg_reg[1007]  ( .D(N1025), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1007]) );
  DFF \round_reg_reg[1008]  ( .D(N1026), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1008]) );
  DFF \round_reg_reg[1009]  ( .D(N1027), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1009]) );
  DFF \round_reg_reg[1010]  ( .D(N1028), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1010]) );
  DFF \round_reg_reg[1011]  ( .D(N1029), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1011]) );
  DFF \round_reg_reg[1012]  ( .D(N1030), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1012]) );
  DFF \round_reg_reg[1013]  ( .D(N1031), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1013]) );
  DFF \round_reg_reg[1014]  ( .D(N1032), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1014]) );
  DFF \round_reg_reg[1015]  ( .D(N1033), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1015]) );
  DFF \round_reg_reg[1016]  ( .D(N1034), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1016]) );
  DFF \round_reg_reg[1017]  ( .D(N1035), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1017]) );
  DFF \round_reg_reg[1018]  ( .D(N1036), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1018]) );
  DFF \round_reg_reg[1019]  ( .D(N1037), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1019]) );
  DFF \round_reg_reg[1020]  ( .D(N1038), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1020]) );
  DFF \round_reg_reg[1021]  ( .D(N1039), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1021]) );
  DFF \round_reg_reg[1022]  ( .D(N1040), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1022]) );
  DFF \round_reg_reg[1023]  ( .D(N1041), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1023]) );
  DFF \round_reg_reg[1024]  ( .D(N1042), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1024]) );
  DFF \round_reg_reg[1025]  ( .D(N1043), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1025]) );
  DFF \round_reg_reg[1026]  ( .D(N1044), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1026]) );
  DFF \round_reg_reg[1027]  ( .D(N1045), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1027]) );
  DFF \round_reg_reg[1028]  ( .D(N1046), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1028]) );
  DFF \round_reg_reg[1029]  ( .D(N1047), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1029]) );
  DFF \round_reg_reg[1030]  ( .D(N1048), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1030]) );
  DFF \round_reg_reg[1031]  ( .D(N1049), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1031]) );
  DFF \round_reg_reg[1032]  ( .D(N1050), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1032]) );
  DFF \round_reg_reg[1033]  ( .D(N1051), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1033]) );
  DFF \round_reg_reg[1034]  ( .D(N1052), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1034]) );
  DFF \round_reg_reg[1035]  ( .D(N1053), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1035]) );
  DFF \round_reg_reg[1036]  ( .D(N1054), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1036]) );
  DFF \round_reg_reg[1037]  ( .D(N1055), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1037]) );
  DFF \round_reg_reg[1038]  ( .D(N1056), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1038]) );
  DFF \round_reg_reg[1039]  ( .D(N1057), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1039]) );
  DFF \round_reg_reg[1040]  ( .D(N1058), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1040]) );
  DFF \round_reg_reg[1041]  ( .D(N1059), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1041]) );
  DFF \round_reg_reg[1042]  ( .D(N1060), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1042]) );
  DFF \round_reg_reg[1043]  ( .D(N1061), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1043]) );
  DFF \round_reg_reg[1044]  ( .D(N1062), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1044]) );
  DFF \round_reg_reg[1045]  ( .D(N1063), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1045]) );
  DFF \round_reg_reg[1046]  ( .D(N1064), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1046]) );
  DFF \round_reg_reg[1047]  ( .D(N1065), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1047]) );
  DFF \round_reg_reg[1048]  ( .D(N1066), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1048]) );
  DFF \round_reg_reg[1049]  ( .D(N1067), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1049]) );
  DFF \round_reg_reg[1050]  ( .D(N1068), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1050]) );
  DFF \round_reg_reg[1051]  ( .D(N1069), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1051]) );
  DFF \round_reg_reg[1052]  ( .D(N1070), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1052]) );
  DFF \round_reg_reg[1053]  ( .D(N1071), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1053]) );
  DFF \round_reg_reg[1054]  ( .D(N1072), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1054]) );
  DFF \round_reg_reg[1055]  ( .D(N1073), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1055]) );
  DFF \round_reg_reg[1056]  ( .D(N1074), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1056]) );
  DFF \round_reg_reg[1057]  ( .D(N1075), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1057]) );
  DFF \round_reg_reg[1058]  ( .D(N1076), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1058]) );
  DFF \round_reg_reg[1059]  ( .D(N1077), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1059]) );
  DFF \round_reg_reg[1060]  ( .D(N1078), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1060]) );
  DFF \round_reg_reg[1061]  ( .D(N1079), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1061]) );
  DFF \round_reg_reg[1062]  ( .D(N1080), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1062]) );
  DFF \round_reg_reg[1063]  ( .D(N1081), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1063]) );
  DFF \round_reg_reg[1064]  ( .D(N1082), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1064]) );
  DFF \round_reg_reg[1065]  ( .D(N1083), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1065]) );
  DFF \round_reg_reg[1066]  ( .D(N1084), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1066]) );
  DFF \round_reg_reg[1067]  ( .D(N1085), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1067]) );
  DFF \round_reg_reg[1068]  ( .D(N1086), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1068]) );
  DFF \round_reg_reg[1069]  ( .D(N1087), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1069]) );
  DFF \round_reg_reg[1070]  ( .D(N1088), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1070]) );
  DFF \round_reg_reg[1071]  ( .D(N1089), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1071]) );
  DFF \round_reg_reg[1072]  ( .D(N1090), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1072]) );
  DFF \round_reg_reg[1073]  ( .D(N1091), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1073]) );
  DFF \round_reg_reg[1074]  ( .D(N1092), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1074]) );
  DFF \round_reg_reg[1075]  ( .D(N1093), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1075]) );
  DFF \round_reg_reg[1076]  ( .D(N1094), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1076]) );
  DFF \round_reg_reg[1077]  ( .D(N1095), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1077]) );
  DFF \round_reg_reg[1078]  ( .D(N1096), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1078]) );
  DFF \round_reg_reg[1079]  ( .D(N1097), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1079]) );
  DFF \round_reg_reg[1080]  ( .D(N1098), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1080]) );
  DFF \round_reg_reg[1081]  ( .D(N1099), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1081]) );
  DFF \round_reg_reg[1082]  ( .D(N1100), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1082]) );
  DFF \round_reg_reg[1083]  ( .D(N1101), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1083]) );
  DFF \round_reg_reg[1084]  ( .D(N1102), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1084]) );
  DFF \round_reg_reg[1085]  ( .D(N1103), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1085]) );
  DFF \round_reg_reg[1086]  ( .D(N1104), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1086]) );
  DFF \round_reg_reg[1087]  ( .D(N1105), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1087]) );
  DFF \round_reg_reg[1088]  ( .D(N1106), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1088]) );
  DFF \round_reg_reg[1089]  ( .D(N1107), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1089]) );
  DFF \round_reg_reg[1090]  ( .D(N1108), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1090]) );
  DFF \round_reg_reg[1091]  ( .D(N1109), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1091]) );
  DFF \round_reg_reg[1092]  ( .D(N1110), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1092]) );
  DFF \round_reg_reg[1093]  ( .D(N1111), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1093]) );
  DFF \round_reg_reg[1094]  ( .D(N1112), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1094]) );
  DFF \round_reg_reg[1095]  ( .D(N1113), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1095]) );
  DFF \round_reg_reg[1096]  ( .D(N1114), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1096]) );
  DFF \round_reg_reg[1097]  ( .D(N1115), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1097]) );
  DFF \round_reg_reg[1098]  ( .D(N1116), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1098]) );
  DFF \round_reg_reg[1099]  ( .D(N1117), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1099]) );
  DFF \round_reg_reg[1100]  ( .D(N1118), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1100]) );
  DFF \round_reg_reg[1101]  ( .D(N1119), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1101]) );
  DFF \round_reg_reg[1102]  ( .D(N1120), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1102]) );
  DFF \round_reg_reg[1103]  ( .D(N1121), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1103]) );
  DFF \round_reg_reg[1104]  ( .D(N1122), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1104]) );
  DFF \round_reg_reg[1105]  ( .D(N1123), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1105]) );
  DFF \round_reg_reg[1106]  ( .D(N1124), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1106]) );
  DFF \round_reg_reg[1107]  ( .D(N1125), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1107]) );
  DFF \round_reg_reg[1108]  ( .D(N1126), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1108]) );
  DFF \round_reg_reg[1109]  ( .D(N1127), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1109]) );
  DFF \round_reg_reg[1110]  ( .D(N1128), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1110]) );
  DFF \round_reg_reg[1111]  ( .D(N1129), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1111]) );
  DFF \round_reg_reg[1112]  ( .D(N1130), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1112]) );
  DFF \round_reg_reg[1113]  ( .D(N1131), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1113]) );
  DFF \round_reg_reg[1114]  ( .D(N1132), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1114]) );
  DFF \round_reg_reg[1115]  ( .D(N1133), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1115]) );
  DFF \round_reg_reg[1116]  ( .D(N1134), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1116]) );
  DFF \round_reg_reg[1117]  ( .D(N1135), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1117]) );
  DFF \round_reg_reg[1118]  ( .D(N1136), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1118]) );
  DFF \round_reg_reg[1119]  ( .D(N1137), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1119]) );
  DFF \round_reg_reg[1120]  ( .D(N1138), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1120]) );
  DFF \round_reg_reg[1121]  ( .D(N1139), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1121]) );
  DFF \round_reg_reg[1122]  ( .D(N1140), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1122]) );
  DFF \round_reg_reg[1123]  ( .D(N1141), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1123]) );
  DFF \round_reg_reg[1124]  ( .D(N1142), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1124]) );
  DFF \round_reg_reg[1125]  ( .D(N1143), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1125]) );
  DFF \round_reg_reg[1126]  ( .D(N1144), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1126]) );
  DFF \round_reg_reg[1127]  ( .D(N1145), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1127]) );
  DFF \round_reg_reg[1128]  ( .D(N1146), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1128]) );
  DFF \round_reg_reg[1129]  ( .D(N1147), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1129]) );
  DFF \round_reg_reg[1130]  ( .D(N1148), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1130]) );
  DFF \round_reg_reg[1131]  ( .D(N1149), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1131]) );
  DFF \round_reg_reg[1132]  ( .D(N1150), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1132]) );
  DFF \round_reg_reg[1133]  ( .D(N1151), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1133]) );
  DFF \round_reg_reg[1134]  ( .D(N1152), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1134]) );
  DFF \round_reg_reg[1135]  ( .D(N1153), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1135]) );
  DFF \round_reg_reg[1136]  ( .D(N1154), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1136]) );
  DFF \round_reg_reg[1137]  ( .D(N1155), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1137]) );
  DFF \round_reg_reg[1138]  ( .D(N1156), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1138]) );
  DFF \round_reg_reg[1139]  ( .D(N1157), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1139]) );
  DFF \round_reg_reg[1140]  ( .D(N1158), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1140]) );
  DFF \round_reg_reg[1141]  ( .D(N1159), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1141]) );
  DFF \round_reg_reg[1142]  ( .D(N1160), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1142]) );
  DFF \round_reg_reg[1143]  ( .D(N1161), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1143]) );
  DFF \round_reg_reg[1144]  ( .D(N1162), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1144]) );
  DFF \round_reg_reg[1145]  ( .D(N1163), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1145]) );
  DFF \round_reg_reg[1146]  ( .D(N1164), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1146]) );
  DFF \round_reg_reg[1147]  ( .D(N1165), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1147]) );
  DFF \round_reg_reg[1148]  ( .D(N1166), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1148]) );
  DFF \round_reg_reg[1149]  ( .D(N1167), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1149]) );
  DFF \round_reg_reg[1150]  ( .D(N1168), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1150]) );
  DFF \round_reg_reg[1151]  ( .D(N1169), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1151]) );
  DFF \round_reg_reg[1152]  ( .D(N1170), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1152]) );
  DFF \round_reg_reg[1153]  ( .D(N1171), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1153]) );
  DFF \round_reg_reg[1154]  ( .D(N1172), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1154]) );
  DFF \round_reg_reg[1155]  ( .D(N1173), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1155]) );
  DFF \round_reg_reg[1156]  ( .D(N1174), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1156]) );
  DFF \round_reg_reg[1157]  ( .D(N1175), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1157]) );
  DFF \round_reg_reg[1158]  ( .D(N1176), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1158]) );
  DFF \round_reg_reg[1159]  ( .D(N1177), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1159]) );
  DFF \round_reg_reg[1160]  ( .D(N1178), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1160]) );
  DFF \round_reg_reg[1161]  ( .D(N1179), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1161]) );
  DFF \round_reg_reg[1162]  ( .D(N1180), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1162]) );
  DFF \round_reg_reg[1163]  ( .D(N1181), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1163]) );
  DFF \round_reg_reg[1164]  ( .D(N1182), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1164]) );
  DFF \round_reg_reg[1165]  ( .D(N1183), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1165]) );
  DFF \round_reg_reg[1166]  ( .D(N1184), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1166]) );
  DFF \round_reg_reg[1167]  ( .D(N1185), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1167]) );
  DFF \round_reg_reg[1168]  ( .D(N1186), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1168]) );
  DFF \round_reg_reg[1169]  ( .D(N1187), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1169]) );
  DFF \round_reg_reg[1170]  ( .D(N1188), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1170]) );
  DFF \round_reg_reg[1171]  ( .D(N1189), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1171]) );
  DFF \round_reg_reg[1172]  ( .D(N1190), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1172]) );
  DFF \round_reg_reg[1173]  ( .D(N1191), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1173]) );
  DFF \round_reg_reg[1174]  ( .D(N1192), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1174]) );
  DFF \round_reg_reg[1175]  ( .D(N1193), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1175]) );
  DFF \round_reg_reg[1176]  ( .D(N1194), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1176]) );
  DFF \round_reg_reg[1177]  ( .D(N1195), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1177]) );
  DFF \round_reg_reg[1178]  ( .D(N1196), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1178]) );
  DFF \round_reg_reg[1179]  ( .D(N1197), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1179]) );
  DFF \round_reg_reg[1180]  ( .D(N1198), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1180]) );
  DFF \round_reg_reg[1181]  ( .D(N1199), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1181]) );
  DFF \round_reg_reg[1182]  ( .D(N1200), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1182]) );
  DFF \round_reg_reg[1183]  ( .D(N1201), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1183]) );
  DFF \round_reg_reg[1184]  ( .D(N1202), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1184]) );
  DFF \round_reg_reg[1185]  ( .D(N1203), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1185]) );
  DFF \round_reg_reg[1186]  ( .D(N1204), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1186]) );
  DFF \round_reg_reg[1187]  ( .D(N1205), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1187]) );
  DFF \round_reg_reg[1188]  ( .D(N1206), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1188]) );
  DFF \round_reg_reg[1189]  ( .D(N1207), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1189]) );
  DFF \round_reg_reg[1190]  ( .D(N1208), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1190]) );
  DFF \round_reg_reg[1191]  ( .D(N1209), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1191]) );
  DFF \round_reg_reg[1192]  ( .D(N1210), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1192]) );
  DFF \round_reg_reg[1193]  ( .D(N1211), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1193]) );
  DFF \round_reg_reg[1194]  ( .D(N1212), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1194]) );
  DFF \round_reg_reg[1195]  ( .D(N1213), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1195]) );
  DFF \round_reg_reg[1196]  ( .D(N1214), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1196]) );
  DFF \round_reg_reg[1197]  ( .D(N1215), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1197]) );
  DFF \round_reg_reg[1198]  ( .D(N1216), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1198]) );
  DFF \round_reg_reg[1199]  ( .D(N1217), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1199]) );
  DFF \round_reg_reg[1200]  ( .D(N1218), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1200]) );
  DFF \round_reg_reg[1201]  ( .D(N1219), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1201]) );
  DFF \round_reg_reg[1202]  ( .D(N1220), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1202]) );
  DFF \round_reg_reg[1203]  ( .D(N1221), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1203]) );
  DFF \round_reg_reg[1204]  ( .D(N1222), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1204]) );
  DFF \round_reg_reg[1205]  ( .D(N1223), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1205]) );
  DFF \round_reg_reg[1206]  ( .D(N1224), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1206]) );
  DFF \round_reg_reg[1207]  ( .D(N1225), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1207]) );
  DFF \round_reg_reg[1208]  ( .D(N1226), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1208]) );
  DFF \round_reg_reg[1209]  ( .D(N1227), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1209]) );
  DFF \round_reg_reg[1210]  ( .D(N1228), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1210]) );
  DFF \round_reg_reg[1211]  ( .D(N1229), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1211]) );
  DFF \round_reg_reg[1212]  ( .D(N1230), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1212]) );
  DFF \round_reg_reg[1213]  ( .D(N1231), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1213]) );
  DFF \round_reg_reg[1214]  ( .D(N1232), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1214]) );
  DFF \round_reg_reg[1215]  ( .D(N1233), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1215]) );
  DFF \round_reg_reg[1216]  ( .D(N1234), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1216]) );
  DFF \round_reg_reg[1217]  ( .D(N1235), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1217]) );
  DFF \round_reg_reg[1218]  ( .D(N1236), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1218]) );
  DFF \round_reg_reg[1219]  ( .D(N1237), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1219]) );
  DFF \round_reg_reg[1220]  ( .D(N1238), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1220]) );
  DFF \round_reg_reg[1221]  ( .D(N1239), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1221]) );
  DFF \round_reg_reg[1222]  ( .D(N1240), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1222]) );
  DFF \round_reg_reg[1223]  ( .D(N1241), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1223]) );
  DFF \round_reg_reg[1224]  ( .D(N1242), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1224]) );
  DFF \round_reg_reg[1225]  ( .D(N1243), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1225]) );
  DFF \round_reg_reg[1226]  ( .D(N1244), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1226]) );
  DFF \round_reg_reg[1227]  ( .D(N1245), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1227]) );
  DFF \round_reg_reg[1228]  ( .D(N1246), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1228]) );
  DFF \round_reg_reg[1229]  ( .D(N1247), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1229]) );
  DFF \round_reg_reg[1230]  ( .D(N1248), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1230]) );
  DFF \round_reg_reg[1231]  ( .D(N1249), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1231]) );
  DFF \round_reg_reg[1232]  ( .D(N1250), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1232]) );
  DFF \round_reg_reg[1233]  ( .D(N1251), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1233]) );
  DFF \round_reg_reg[1234]  ( .D(N1252), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1234]) );
  DFF \round_reg_reg[1235]  ( .D(N1253), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1235]) );
  DFF \round_reg_reg[1236]  ( .D(N1254), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1236]) );
  DFF \round_reg_reg[1237]  ( .D(N1255), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1237]) );
  DFF \round_reg_reg[1238]  ( .D(N1256), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1238]) );
  DFF \round_reg_reg[1239]  ( .D(N1257), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1239]) );
  DFF \round_reg_reg[1240]  ( .D(N1258), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1240]) );
  DFF \round_reg_reg[1241]  ( .D(N1259), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1241]) );
  DFF \round_reg_reg[1242]  ( .D(N1260), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1242]) );
  DFF \round_reg_reg[1243]  ( .D(N1261), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1243]) );
  DFF \round_reg_reg[1244]  ( .D(N1262), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1244]) );
  DFF \round_reg_reg[1245]  ( .D(N1263), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1245]) );
  DFF \round_reg_reg[1246]  ( .D(N1264), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1246]) );
  DFF \round_reg_reg[1247]  ( .D(N1265), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1247]) );
  DFF \round_reg_reg[1248]  ( .D(N1266), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1248]) );
  DFF \round_reg_reg[1249]  ( .D(N1267), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1249]) );
  DFF \round_reg_reg[1250]  ( .D(N1268), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1250]) );
  DFF \round_reg_reg[1251]  ( .D(N1269), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1251]) );
  DFF \round_reg_reg[1252]  ( .D(N1270), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1252]) );
  DFF \round_reg_reg[1253]  ( .D(N1271), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1253]) );
  DFF \round_reg_reg[1254]  ( .D(N1272), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1254]) );
  DFF \round_reg_reg[1255]  ( .D(N1273), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1255]) );
  DFF \round_reg_reg[1256]  ( .D(N1274), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1256]) );
  DFF \round_reg_reg[1257]  ( .D(N1275), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1257]) );
  DFF \round_reg_reg[1258]  ( .D(N1276), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1258]) );
  DFF \round_reg_reg[1259]  ( .D(N1277), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1259]) );
  DFF \round_reg_reg[1260]  ( .D(N1278), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1260]) );
  DFF \round_reg_reg[1261]  ( .D(N1279), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1261]) );
  DFF \round_reg_reg[1262]  ( .D(N1280), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1262]) );
  DFF \round_reg_reg[1263]  ( .D(N1281), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1263]) );
  DFF \round_reg_reg[1264]  ( .D(N1282), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1264]) );
  DFF \round_reg_reg[1265]  ( .D(N1283), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1265]) );
  DFF \round_reg_reg[1266]  ( .D(N1284), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1266]) );
  DFF \round_reg_reg[1267]  ( .D(N1285), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1267]) );
  DFF \round_reg_reg[1268]  ( .D(N1286), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1268]) );
  DFF \round_reg_reg[1269]  ( .D(N1287), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1269]) );
  DFF \round_reg_reg[1270]  ( .D(N1288), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1270]) );
  DFF \round_reg_reg[1271]  ( .D(N1289), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1271]) );
  DFF \round_reg_reg[1272]  ( .D(N1290), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1272]) );
  DFF \round_reg_reg[1273]  ( .D(N1291), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1273]) );
  DFF \round_reg_reg[1274]  ( .D(N1292), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1274]) );
  DFF \round_reg_reg[1275]  ( .D(N1293), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1275]) );
  DFF \round_reg_reg[1276]  ( .D(N1294), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1276]) );
  DFF \round_reg_reg[1277]  ( .D(N1295), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1277]) );
  DFF \round_reg_reg[1278]  ( .D(N1296), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1278]) );
  DFF \round_reg_reg[1279]  ( .D(N1297), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1279]) );
  DFF \round_reg_reg[1280]  ( .D(N1298), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1280]) );
  DFF \round_reg_reg[1281]  ( .D(N1299), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1281]) );
  DFF \round_reg_reg[1282]  ( .D(N1300), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1282]) );
  DFF \round_reg_reg[1283]  ( .D(N1301), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1283]) );
  DFF \round_reg_reg[1284]  ( .D(N1302), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1284]) );
  DFF \round_reg_reg[1285]  ( .D(N1303), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1285]) );
  DFF \round_reg_reg[1286]  ( .D(N1304), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1286]) );
  DFF \round_reg_reg[1287]  ( .D(N1305), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1287]) );
  DFF \round_reg_reg[1288]  ( .D(N1306), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1288]) );
  DFF \round_reg_reg[1289]  ( .D(N1307), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1289]) );
  DFF \round_reg_reg[1290]  ( .D(N1308), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1290]) );
  DFF \round_reg_reg[1291]  ( .D(N1309), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1291]) );
  DFF \round_reg_reg[1292]  ( .D(N1310), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1292]) );
  DFF \round_reg_reg[1293]  ( .D(N1311), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1293]) );
  DFF \round_reg_reg[1294]  ( .D(N1312), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1294]) );
  DFF \round_reg_reg[1295]  ( .D(N1313), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1295]) );
  DFF \round_reg_reg[1296]  ( .D(N1314), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1296]) );
  DFF \round_reg_reg[1297]  ( .D(N1315), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1297]) );
  DFF \round_reg_reg[1298]  ( .D(N1316), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1298]) );
  DFF \round_reg_reg[1299]  ( .D(N1317), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1299]) );
  DFF \round_reg_reg[1300]  ( .D(N1318), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1300]) );
  DFF \round_reg_reg[1301]  ( .D(N1319), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1301]) );
  DFF \round_reg_reg[1302]  ( .D(N1320), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1302]) );
  DFF \round_reg_reg[1303]  ( .D(N1321), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1303]) );
  DFF \round_reg_reg[1304]  ( .D(N1322), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1304]) );
  DFF \round_reg_reg[1305]  ( .D(N1323), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1305]) );
  DFF \round_reg_reg[1306]  ( .D(N1324), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1306]) );
  DFF \round_reg_reg[1307]  ( .D(N1325), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1307]) );
  DFF \round_reg_reg[1308]  ( .D(N1326), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1308]) );
  DFF \round_reg_reg[1309]  ( .D(N1327), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1309]) );
  DFF \round_reg_reg[1310]  ( .D(N1328), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1310]) );
  DFF \round_reg_reg[1311]  ( .D(N1329), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1311]) );
  DFF \round_reg_reg[1312]  ( .D(N1330), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1312]) );
  DFF \round_reg_reg[1313]  ( .D(N1331), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1313]) );
  DFF \round_reg_reg[1314]  ( .D(N1332), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1314]) );
  DFF \round_reg_reg[1315]  ( .D(N1333), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1315]) );
  DFF \round_reg_reg[1316]  ( .D(N1334), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1316]) );
  DFF \round_reg_reg[1317]  ( .D(N1335), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1317]) );
  DFF \round_reg_reg[1318]  ( .D(N1336), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1318]) );
  DFF \round_reg_reg[1319]  ( .D(N1337), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1319]) );
  DFF \round_reg_reg[1320]  ( .D(N1338), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1320]) );
  DFF \round_reg_reg[1321]  ( .D(N1339), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1321]) );
  DFF \round_reg_reg[1322]  ( .D(N1340), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1322]) );
  DFF \round_reg_reg[1323]  ( .D(N1341), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1323]) );
  DFF \round_reg_reg[1324]  ( .D(N1342), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1324]) );
  DFF \round_reg_reg[1325]  ( .D(N1343), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1325]) );
  DFF \round_reg_reg[1326]  ( .D(N1344), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1326]) );
  DFF \round_reg_reg[1327]  ( .D(N1345), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1327]) );
  DFF \round_reg_reg[1328]  ( .D(N1346), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1328]) );
  DFF \round_reg_reg[1329]  ( .D(N1347), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1329]) );
  DFF \round_reg_reg[1330]  ( .D(N1348), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1330]) );
  DFF \round_reg_reg[1331]  ( .D(N1349), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1331]) );
  DFF \round_reg_reg[1332]  ( .D(N1350), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1332]) );
  DFF \round_reg_reg[1333]  ( .D(N1351), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1333]) );
  DFF \round_reg_reg[1334]  ( .D(N1352), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1334]) );
  DFF \round_reg_reg[1335]  ( .D(N1353), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1335]) );
  DFF \round_reg_reg[1336]  ( .D(N1354), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1336]) );
  DFF \round_reg_reg[1337]  ( .D(N1355), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1337]) );
  DFF \round_reg_reg[1338]  ( .D(N1356), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1338]) );
  DFF \round_reg_reg[1339]  ( .D(N1357), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1339]) );
  DFF \round_reg_reg[1340]  ( .D(N1358), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1340]) );
  DFF \round_reg_reg[1341]  ( .D(N1359), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1341]) );
  DFF \round_reg_reg[1342]  ( .D(N1360), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1342]) );
  DFF \round_reg_reg[1343]  ( .D(N1361), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1343]) );
  DFF \round_reg_reg[1344]  ( .D(N1362), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1344]) );
  DFF \round_reg_reg[1345]  ( .D(N1363), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1345]) );
  DFF \round_reg_reg[1346]  ( .D(N1364), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1346]) );
  DFF \round_reg_reg[1347]  ( .D(N1365), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1347]) );
  DFF \round_reg_reg[1348]  ( .D(N1366), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1348]) );
  DFF \round_reg_reg[1349]  ( .D(N1367), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1349]) );
  DFF \round_reg_reg[1350]  ( .D(N1368), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1350]) );
  DFF \round_reg_reg[1351]  ( .D(N1369), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1351]) );
  DFF \round_reg_reg[1352]  ( .D(N1370), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1352]) );
  DFF \round_reg_reg[1353]  ( .D(N1371), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1353]) );
  DFF \round_reg_reg[1354]  ( .D(N1372), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1354]) );
  DFF \round_reg_reg[1355]  ( .D(N1373), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1355]) );
  DFF \round_reg_reg[1356]  ( .D(N1374), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1356]) );
  DFF \round_reg_reg[1357]  ( .D(N1375), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1357]) );
  DFF \round_reg_reg[1358]  ( .D(N1376), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1358]) );
  DFF \round_reg_reg[1359]  ( .D(N1377), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1359]) );
  DFF \round_reg_reg[1360]  ( .D(N1378), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1360]) );
  DFF \round_reg_reg[1361]  ( .D(N1379), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1361]) );
  DFF \round_reg_reg[1362]  ( .D(N1380), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1362]) );
  DFF \round_reg_reg[1363]  ( .D(N1381), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1363]) );
  DFF \round_reg_reg[1364]  ( .D(N1382), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1364]) );
  DFF \round_reg_reg[1365]  ( .D(N1383), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1365]) );
  DFF \round_reg_reg[1366]  ( .D(N1384), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1366]) );
  DFF \round_reg_reg[1367]  ( .D(N1385), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1367]) );
  DFF \round_reg_reg[1368]  ( .D(N1386), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1368]) );
  DFF \round_reg_reg[1369]  ( .D(N1387), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1369]) );
  DFF \round_reg_reg[1370]  ( .D(N1388), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1370]) );
  DFF \round_reg_reg[1371]  ( .D(N1389), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1371]) );
  DFF \round_reg_reg[1372]  ( .D(N1390), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1372]) );
  DFF \round_reg_reg[1373]  ( .D(N1391), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1373]) );
  DFF \round_reg_reg[1374]  ( .D(N1392), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1374]) );
  DFF \round_reg_reg[1375]  ( .D(N1393), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1375]) );
  DFF \round_reg_reg[1376]  ( .D(N1394), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1376]) );
  DFF \round_reg_reg[1377]  ( .D(N1395), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1377]) );
  DFF \round_reg_reg[1378]  ( .D(N1396), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1378]) );
  DFF \round_reg_reg[1379]  ( .D(N1397), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1379]) );
  DFF \round_reg_reg[1380]  ( .D(N1398), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1380]) );
  DFF \round_reg_reg[1381]  ( .D(N1399), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1381]) );
  DFF \round_reg_reg[1382]  ( .D(N1400), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1382]) );
  DFF \round_reg_reg[1383]  ( .D(N1401), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1383]) );
  DFF \round_reg_reg[1384]  ( .D(N1402), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1384]) );
  DFF \round_reg_reg[1385]  ( .D(N1403), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1385]) );
  DFF \round_reg_reg[1386]  ( .D(N1404), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1386]) );
  DFF \round_reg_reg[1387]  ( .D(N1405), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1387]) );
  DFF \round_reg_reg[1388]  ( .D(N1406), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1388]) );
  DFF \round_reg_reg[1389]  ( .D(N1407), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1389]) );
  DFF \round_reg_reg[1390]  ( .D(N1408), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1390]) );
  DFF \round_reg_reg[1391]  ( .D(N1409), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1391]) );
  DFF \round_reg_reg[1392]  ( .D(N1410), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1392]) );
  DFF \round_reg_reg[1393]  ( .D(N1411), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1393]) );
  DFF \round_reg_reg[1394]  ( .D(N1412), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1394]) );
  DFF \round_reg_reg[1395]  ( .D(N1413), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1395]) );
  DFF \round_reg_reg[1396]  ( .D(N1414), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1396]) );
  DFF \round_reg_reg[1397]  ( .D(N1415), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1397]) );
  DFF \round_reg_reg[1398]  ( .D(N1416), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1398]) );
  DFF \round_reg_reg[1399]  ( .D(N1417), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1399]) );
  DFF \round_reg_reg[1400]  ( .D(N1418), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1400]) );
  DFF \round_reg_reg[1401]  ( .D(N1419), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1401]) );
  DFF \round_reg_reg[1402]  ( .D(N1420), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1402]) );
  DFF \round_reg_reg[1403]  ( .D(N1421), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1403]) );
  DFF \round_reg_reg[1404]  ( .D(N1422), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1404]) );
  DFF \round_reg_reg[1405]  ( .D(N1423), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1405]) );
  DFF \round_reg_reg[1406]  ( .D(N1424), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1406]) );
  DFF \round_reg_reg[1407]  ( .D(N1425), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1407]) );
  DFF \round_reg_reg[1408]  ( .D(N1426), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1408]) );
  DFF \round_reg_reg[1409]  ( .D(N1427), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1409]) );
  DFF \round_reg_reg[1410]  ( .D(N1428), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1410]) );
  DFF \round_reg_reg[1411]  ( .D(N1429), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1411]) );
  DFF \round_reg_reg[1412]  ( .D(N1430), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1412]) );
  DFF \round_reg_reg[1413]  ( .D(N1431), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1413]) );
  DFF \round_reg_reg[1414]  ( .D(N1432), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1414]) );
  DFF \round_reg_reg[1415]  ( .D(N1433), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1415]) );
  DFF \round_reg_reg[1416]  ( .D(N1434), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1416]) );
  DFF \round_reg_reg[1417]  ( .D(N1435), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1417]) );
  DFF \round_reg_reg[1418]  ( .D(N1436), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1418]) );
  DFF \round_reg_reg[1419]  ( .D(N1437), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1419]) );
  DFF \round_reg_reg[1420]  ( .D(N1438), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1420]) );
  DFF \round_reg_reg[1421]  ( .D(N1439), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1421]) );
  DFF \round_reg_reg[1422]  ( .D(N1440), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1422]) );
  DFF \round_reg_reg[1423]  ( .D(N1441), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1423]) );
  DFF \round_reg_reg[1424]  ( .D(N1442), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1424]) );
  DFF \round_reg_reg[1425]  ( .D(N1443), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1425]) );
  DFF \round_reg_reg[1426]  ( .D(N1444), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1426]) );
  DFF \round_reg_reg[1427]  ( .D(N1445), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1427]) );
  DFF \round_reg_reg[1428]  ( .D(N1446), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1428]) );
  DFF \round_reg_reg[1429]  ( .D(N1447), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1429]) );
  DFF \round_reg_reg[1430]  ( .D(N1448), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1430]) );
  DFF \round_reg_reg[1431]  ( .D(N1449), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1431]) );
  DFF \round_reg_reg[1432]  ( .D(N1450), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1432]) );
  DFF \round_reg_reg[1433]  ( .D(N1451), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1433]) );
  DFF \round_reg_reg[1434]  ( .D(N1452), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1434]) );
  DFF \round_reg_reg[1435]  ( .D(N1453), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1435]) );
  DFF \round_reg_reg[1436]  ( .D(N1454), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1436]) );
  DFF \round_reg_reg[1437]  ( .D(N1455), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1437]) );
  DFF \round_reg_reg[1438]  ( .D(N1456), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1438]) );
  DFF \round_reg_reg[1439]  ( .D(N1457), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1439]) );
  DFF \round_reg_reg[1440]  ( .D(N1458), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1440]) );
  DFF \round_reg_reg[1441]  ( .D(N1459), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1441]) );
  DFF \round_reg_reg[1442]  ( .D(N1460), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1442]) );
  DFF \round_reg_reg[1443]  ( .D(N1461), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1443]) );
  DFF \round_reg_reg[1444]  ( .D(N1462), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1444]) );
  DFF \round_reg_reg[1445]  ( .D(N1463), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1445]) );
  DFF \round_reg_reg[1446]  ( .D(N1464), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1446]) );
  DFF \round_reg_reg[1447]  ( .D(N1465), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1447]) );
  DFF \round_reg_reg[1448]  ( .D(N1466), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1448]) );
  DFF \round_reg_reg[1449]  ( .D(N1467), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1449]) );
  DFF \round_reg_reg[1450]  ( .D(N1468), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1450]) );
  DFF \round_reg_reg[1451]  ( .D(N1469), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1451]) );
  DFF \round_reg_reg[1452]  ( .D(N1470), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1452]) );
  DFF \round_reg_reg[1453]  ( .D(N1471), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1453]) );
  DFF \round_reg_reg[1454]  ( .D(N1472), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1454]) );
  DFF \round_reg_reg[1455]  ( .D(N1473), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1455]) );
  DFF \round_reg_reg[1456]  ( .D(N1474), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1456]) );
  DFF \round_reg_reg[1457]  ( .D(N1475), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1457]) );
  DFF \round_reg_reg[1458]  ( .D(N1476), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1458]) );
  DFF \round_reg_reg[1459]  ( .D(N1477), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1459]) );
  DFF \round_reg_reg[1460]  ( .D(N1478), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1460]) );
  DFF \round_reg_reg[1461]  ( .D(N1479), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1461]) );
  DFF \round_reg_reg[1462]  ( .D(N1480), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1462]) );
  DFF \round_reg_reg[1463]  ( .D(N1481), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1463]) );
  DFF \round_reg_reg[1464]  ( .D(N1482), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1464]) );
  DFF \round_reg_reg[1465]  ( .D(N1483), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1465]) );
  DFF \round_reg_reg[1466]  ( .D(N1484), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1466]) );
  DFF \round_reg_reg[1467]  ( .D(N1485), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1467]) );
  DFF \round_reg_reg[1468]  ( .D(N1486), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1468]) );
  DFF \round_reg_reg[1469]  ( .D(N1487), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1469]) );
  DFF \round_reg_reg[1470]  ( .D(N1488), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1470]) );
  DFF \round_reg_reg[1471]  ( .D(N1489), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1471]) );
  DFF \round_reg_reg[1472]  ( .D(N1490), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1472]) );
  DFF \round_reg_reg[1473]  ( .D(N1491), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1473]) );
  DFF \round_reg_reg[1474]  ( .D(N1492), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1474]) );
  DFF \round_reg_reg[1475]  ( .D(N1493), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1475]) );
  DFF \round_reg_reg[1476]  ( .D(N1494), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1476]) );
  DFF \round_reg_reg[1477]  ( .D(N1495), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1477]) );
  DFF \round_reg_reg[1478]  ( .D(N1496), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1478]) );
  DFF \round_reg_reg[1479]  ( .D(N1497), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1479]) );
  DFF \round_reg_reg[1480]  ( .D(N1498), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1480]) );
  DFF \round_reg_reg[1481]  ( .D(N1499), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1481]) );
  DFF \round_reg_reg[1482]  ( .D(N1500), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1482]) );
  DFF \round_reg_reg[1483]  ( .D(N1501), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1483]) );
  DFF \round_reg_reg[1484]  ( .D(N1502), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1484]) );
  DFF \round_reg_reg[1485]  ( .D(N1503), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1485]) );
  DFF \round_reg_reg[1486]  ( .D(N1504), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1486]) );
  DFF \round_reg_reg[1487]  ( .D(N1505), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1487]) );
  DFF \round_reg_reg[1488]  ( .D(N1506), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1488]) );
  DFF \round_reg_reg[1489]  ( .D(N1507), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1489]) );
  DFF \round_reg_reg[1490]  ( .D(N1508), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1490]) );
  DFF \round_reg_reg[1491]  ( .D(N1509), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1491]) );
  DFF \round_reg_reg[1492]  ( .D(N1510), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1492]) );
  DFF \round_reg_reg[1493]  ( .D(N1511), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1493]) );
  DFF \round_reg_reg[1494]  ( .D(N1512), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1494]) );
  DFF \round_reg_reg[1495]  ( .D(N1513), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1495]) );
  DFF \round_reg_reg[1496]  ( .D(N1514), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1496]) );
  DFF \round_reg_reg[1497]  ( .D(N1515), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1497]) );
  DFF \round_reg_reg[1498]  ( .D(N1516), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1498]) );
  DFF \round_reg_reg[1499]  ( .D(N1517), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1499]) );
  DFF \round_reg_reg[1500]  ( .D(N1518), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1500]) );
  DFF \round_reg_reg[1501]  ( .D(N1519), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1501]) );
  DFF \round_reg_reg[1502]  ( .D(N1520), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1502]) );
  DFF \round_reg_reg[1503]  ( .D(N1521), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1503]) );
  DFF \round_reg_reg[1504]  ( .D(N1522), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1504]) );
  DFF \round_reg_reg[1505]  ( .D(N1523), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1505]) );
  DFF \round_reg_reg[1506]  ( .D(N1524), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1506]) );
  DFF \round_reg_reg[1507]  ( .D(N1525), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1507]) );
  DFF \round_reg_reg[1508]  ( .D(N1526), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1508]) );
  DFF \round_reg_reg[1509]  ( .D(N1527), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1509]) );
  DFF \round_reg_reg[1510]  ( .D(N1528), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1510]) );
  DFF \round_reg_reg[1511]  ( .D(N1529), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1511]) );
  DFF \round_reg_reg[1512]  ( .D(N1530), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1512]) );
  DFF \round_reg_reg[1513]  ( .D(N1531), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1513]) );
  DFF \round_reg_reg[1514]  ( .D(N1532), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1514]) );
  DFF \round_reg_reg[1515]  ( .D(N1533), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1515]) );
  DFF \round_reg_reg[1516]  ( .D(N1534), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1516]) );
  DFF \round_reg_reg[1517]  ( .D(N1535), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1517]) );
  DFF \round_reg_reg[1518]  ( .D(N1536), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1518]) );
  DFF \round_reg_reg[1519]  ( .D(N1537), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1519]) );
  DFF \round_reg_reg[1520]  ( .D(N1538), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1520]) );
  DFF \round_reg_reg[1521]  ( .D(N1539), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1521]) );
  DFF \round_reg_reg[1522]  ( .D(N1540), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1522]) );
  DFF \round_reg_reg[1523]  ( .D(N1541), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1523]) );
  DFF \round_reg_reg[1524]  ( .D(N1542), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1524]) );
  DFF \round_reg_reg[1525]  ( .D(N1543), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1525]) );
  DFF \round_reg_reg[1526]  ( .D(N1544), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1526]) );
  DFF \round_reg_reg[1527]  ( .D(N1545), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1527]) );
  DFF \round_reg_reg[1528]  ( .D(N1546), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1528]) );
  DFF \round_reg_reg[1529]  ( .D(N1547), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1529]) );
  DFF \round_reg_reg[1530]  ( .D(N1548), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1530]) );
  DFF \round_reg_reg[1531]  ( .D(N1549), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1531]) );
  DFF \round_reg_reg[1532]  ( .D(N1550), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1532]) );
  DFF \round_reg_reg[1533]  ( .D(N1551), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1533]) );
  DFF \round_reg_reg[1534]  ( .D(N1552), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1534]) );
  DFF \round_reg_reg[1535]  ( .D(N1553), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1535]) );
  DFF \round_reg_reg[1536]  ( .D(N1554), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1536]) );
  DFF \round_reg_reg[1537]  ( .D(N1555), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1537]) );
  DFF \round_reg_reg[1538]  ( .D(N1556), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1538]) );
  DFF \round_reg_reg[1539]  ( .D(N1557), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1539]) );
  DFF \round_reg_reg[1540]  ( .D(N1558), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1540]) );
  DFF \round_reg_reg[1541]  ( .D(N1559), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1541]) );
  DFF \round_reg_reg[1542]  ( .D(N1560), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1542]) );
  DFF \round_reg_reg[1543]  ( .D(N1561), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1543]) );
  DFF \round_reg_reg[1544]  ( .D(N1562), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1544]) );
  DFF \round_reg_reg[1545]  ( .D(N1563), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1545]) );
  DFF \round_reg_reg[1546]  ( .D(N1564), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1546]) );
  DFF \round_reg_reg[1547]  ( .D(N1565), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1547]) );
  DFF \round_reg_reg[1548]  ( .D(N1566), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1548]) );
  DFF \round_reg_reg[1549]  ( .D(N1567), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1549]) );
  DFF \round_reg_reg[1550]  ( .D(N1568), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1550]) );
  DFF \round_reg_reg[1551]  ( .D(N1569), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1551]) );
  DFF \round_reg_reg[1552]  ( .D(N1570), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1552]) );
  DFF \round_reg_reg[1553]  ( .D(N1571), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1553]) );
  DFF \round_reg_reg[1554]  ( .D(N1572), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1554]) );
  DFF \round_reg_reg[1555]  ( .D(N1573), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1555]) );
  DFF \round_reg_reg[1556]  ( .D(N1574), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1556]) );
  DFF \round_reg_reg[1557]  ( .D(N1575), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1557]) );
  DFF \round_reg_reg[1558]  ( .D(N1576), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1558]) );
  DFF \round_reg_reg[1559]  ( .D(N1577), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1559]) );
  DFF \round_reg_reg[1560]  ( .D(N1578), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1560]) );
  DFF \round_reg_reg[1561]  ( .D(N1579), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1561]) );
  DFF \round_reg_reg[1562]  ( .D(N1580), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1562]) );
  DFF \round_reg_reg[1563]  ( .D(N1581), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1563]) );
  DFF \round_reg_reg[1564]  ( .D(N1582), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1564]) );
  DFF \round_reg_reg[1565]  ( .D(N1583), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1565]) );
  DFF \round_reg_reg[1566]  ( .D(N1584), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1566]) );
  DFF \round_reg_reg[1567]  ( .D(N1585), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1567]) );
  DFF \round_reg_reg[1568]  ( .D(N1586), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1568]) );
  DFF \round_reg_reg[1569]  ( .D(N1587), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1569]) );
  DFF \round_reg_reg[1570]  ( .D(N1588), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1570]) );
  DFF \round_reg_reg[1571]  ( .D(N1589), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1571]) );
  DFF \round_reg_reg[1572]  ( .D(N1590), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1572]) );
  DFF \round_reg_reg[1573]  ( .D(N1591), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1573]) );
  DFF \round_reg_reg[1574]  ( .D(N1592), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1574]) );
  DFF \round_reg_reg[1575]  ( .D(N1593), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1575]) );
  DFF \round_reg_reg[1576]  ( .D(N1594), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1576]) );
  DFF \round_reg_reg[1577]  ( .D(N1595), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1577]) );
  DFF \round_reg_reg[1578]  ( .D(N1596), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1578]) );
  DFF \round_reg_reg[1579]  ( .D(N1597), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1579]) );
  DFF \round_reg_reg[1580]  ( .D(N1598), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1580]) );
  DFF \round_reg_reg[1581]  ( .D(N1599), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1581]) );
  DFF \round_reg_reg[1582]  ( .D(N1600), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1582]) );
  DFF \round_reg_reg[1583]  ( .D(N1601), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1583]) );
  DFF \round_reg_reg[1584]  ( .D(N1602), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1584]) );
  DFF \round_reg_reg[1585]  ( .D(N1603), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1585]) );
  DFF \round_reg_reg[1586]  ( .D(N1604), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1586]) );
  DFF \round_reg_reg[1587]  ( .D(N1605), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1587]) );
  DFF \round_reg_reg[1588]  ( .D(N1606), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1588]) );
  DFF \round_reg_reg[1589]  ( .D(N1607), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1589]) );
  DFF \round_reg_reg[1590]  ( .D(N1608), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1590]) );
  DFF \round_reg_reg[1591]  ( .D(N1609), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1591]) );
  DFF \round_reg_reg[1592]  ( .D(N1610), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1592]) );
  DFF \round_reg_reg[1593]  ( .D(N1611), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1593]) );
  DFF \round_reg_reg[1594]  ( .D(N1612), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1594]) );
  DFF \round_reg_reg[1595]  ( .D(N1613), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1595]) );
  DFF \round_reg_reg[1596]  ( .D(N1614), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1596]) );
  DFF \round_reg_reg[1597]  ( .D(N1615), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1597]) );
  DFF \round_reg_reg[1598]  ( .D(N1616), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1598]) );
  DFF \round_reg_reg[1599]  ( .D(N1617), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1599]) );
  IV U6020 ( .A(rst), .Z(n2792) );
  ANDN U6021 ( .B(rc_i[3]), .A(rst), .Z(N10) );
  ANDN U6022 ( .B(out[82]), .A(rst), .Z(N100) );
  ANDN U6023 ( .B(out[982]), .A(rst), .Z(N1000) );
  ANDN U6024 ( .B(out[983]), .A(rst), .Z(N1001) );
  ANDN U6025 ( .B(out[984]), .A(rst), .Z(N1002) );
  ANDN U6026 ( .B(out[985]), .A(rst), .Z(N1003) );
  ANDN U6027 ( .B(out[986]), .A(rst), .Z(N1004) );
  ANDN U6028 ( .B(out[987]), .A(rst), .Z(N1005) );
  ANDN U6029 ( .B(out[988]), .A(rst), .Z(N1006) );
  ANDN U6030 ( .B(out[989]), .A(rst), .Z(N1007) );
  ANDN U6031 ( .B(out[990]), .A(rst), .Z(N1008) );
  ANDN U6032 ( .B(out[991]), .A(rst), .Z(N1009) );
  ANDN U6033 ( .B(out[83]), .A(rst), .Z(N101) );
  ANDN U6034 ( .B(out[992]), .A(rst), .Z(N1010) );
  ANDN U6035 ( .B(out[993]), .A(rst), .Z(N1011) );
  ANDN U6036 ( .B(out[994]), .A(rst), .Z(N1012) );
  ANDN U6037 ( .B(out[995]), .A(rst), .Z(N1013) );
  ANDN U6038 ( .B(out[996]), .A(rst), .Z(N1014) );
  ANDN U6039 ( .B(out[997]), .A(rst), .Z(N1015) );
  ANDN U6040 ( .B(out[998]), .A(rst), .Z(N1016) );
  ANDN U6041 ( .B(out[999]), .A(rst), .Z(N1017) );
  ANDN U6042 ( .B(out[1000]), .A(rst), .Z(N1018) );
  ANDN U6043 ( .B(out[1001]), .A(rst), .Z(N1019) );
  ANDN U6044 ( .B(out[84]), .A(rst), .Z(N102) );
  ANDN U6045 ( .B(out[1002]), .A(rst), .Z(N1020) );
  ANDN U6046 ( .B(out[1003]), .A(rst), .Z(N1021) );
  ANDN U6047 ( .B(out[1004]), .A(rst), .Z(N1022) );
  ANDN U6048 ( .B(out[1005]), .A(rst), .Z(N1023) );
  ANDN U6049 ( .B(out[1006]), .A(rst), .Z(N1024) );
  ANDN U6050 ( .B(out[1007]), .A(rst), .Z(N1025) );
  ANDN U6051 ( .B(out[1008]), .A(rst), .Z(N1026) );
  ANDN U6052 ( .B(out[1009]), .A(rst), .Z(N1027) );
  ANDN U6053 ( .B(out[1010]), .A(rst), .Z(N1028) );
  ANDN U6054 ( .B(out[1011]), .A(rst), .Z(N1029) );
  ANDN U6055 ( .B(out[85]), .A(rst), .Z(N103) );
  ANDN U6056 ( .B(out[1012]), .A(rst), .Z(N1030) );
  ANDN U6057 ( .B(out[1013]), .A(rst), .Z(N1031) );
  ANDN U6058 ( .B(out[1014]), .A(rst), .Z(N1032) );
  ANDN U6059 ( .B(out[1015]), .A(rst), .Z(N1033) );
  ANDN U6060 ( .B(out[1016]), .A(rst), .Z(N1034) );
  ANDN U6061 ( .B(out[1017]), .A(rst), .Z(N1035) );
  ANDN U6062 ( .B(out[1018]), .A(rst), .Z(N1036) );
  ANDN U6063 ( .B(out[1019]), .A(rst), .Z(N1037) );
  ANDN U6064 ( .B(out[1020]), .A(rst), .Z(N1038) );
  ANDN U6065 ( .B(out[1021]), .A(rst), .Z(N1039) );
  ANDN U6066 ( .B(out[86]), .A(rst), .Z(N104) );
  ANDN U6067 ( .B(out[1022]), .A(rst), .Z(N1040) );
  ANDN U6068 ( .B(out[1023]), .A(rst), .Z(N1041) );
  ANDN U6069 ( .B(out[1024]), .A(rst), .Z(N1042) );
  ANDN U6070 ( .B(out[1025]), .A(rst), .Z(N1043) );
  ANDN U6071 ( .B(out[1026]), .A(rst), .Z(N1044) );
  ANDN U6072 ( .B(out[1027]), .A(rst), .Z(N1045) );
  ANDN U6073 ( .B(out[1028]), .A(rst), .Z(N1046) );
  ANDN U6074 ( .B(out[1029]), .A(rst), .Z(N1047) );
  ANDN U6075 ( .B(out[1030]), .A(rst), .Z(N1048) );
  ANDN U6076 ( .B(out[1031]), .A(rst), .Z(N1049) );
  ANDN U6077 ( .B(out[87]), .A(rst), .Z(N105) );
  ANDN U6078 ( .B(out[1032]), .A(rst), .Z(N1050) );
  ANDN U6079 ( .B(out[1033]), .A(rst), .Z(N1051) );
  ANDN U6080 ( .B(out[1034]), .A(rst), .Z(N1052) );
  ANDN U6081 ( .B(out[1035]), .A(rst), .Z(N1053) );
  ANDN U6082 ( .B(out[1036]), .A(rst), .Z(N1054) );
  ANDN U6083 ( .B(out[1037]), .A(rst), .Z(N1055) );
  ANDN U6084 ( .B(out[1038]), .A(rst), .Z(N1056) );
  ANDN U6085 ( .B(out[1039]), .A(rst), .Z(N1057) );
  ANDN U6086 ( .B(out[1040]), .A(rst), .Z(N1058) );
  ANDN U6087 ( .B(out[1041]), .A(rst), .Z(N1059) );
  ANDN U6088 ( .B(out[88]), .A(rst), .Z(N106) );
  ANDN U6089 ( .B(out[1042]), .A(rst), .Z(N1060) );
  ANDN U6090 ( .B(out[1043]), .A(rst), .Z(N1061) );
  ANDN U6091 ( .B(out[1044]), .A(rst), .Z(N1062) );
  ANDN U6092 ( .B(out[1045]), .A(rst), .Z(N1063) );
  ANDN U6093 ( .B(out[1046]), .A(rst), .Z(N1064) );
  ANDN U6094 ( .B(out[1047]), .A(rst), .Z(N1065) );
  ANDN U6095 ( .B(out[1048]), .A(rst), .Z(N1066) );
  ANDN U6096 ( .B(out[1049]), .A(rst), .Z(N1067) );
  ANDN U6097 ( .B(out[1050]), .A(rst), .Z(N1068) );
  ANDN U6098 ( .B(out[1051]), .A(rst), .Z(N1069) );
  ANDN U6099 ( .B(out[89]), .A(rst), .Z(N107) );
  ANDN U6100 ( .B(out[1052]), .A(rst), .Z(N1070) );
  ANDN U6101 ( .B(out[1053]), .A(rst), .Z(N1071) );
  ANDN U6102 ( .B(out[1054]), .A(rst), .Z(N1072) );
  ANDN U6103 ( .B(out[1055]), .A(rst), .Z(N1073) );
  ANDN U6104 ( .B(out[1056]), .A(rst), .Z(N1074) );
  ANDN U6105 ( .B(out[1057]), .A(rst), .Z(N1075) );
  ANDN U6106 ( .B(out[1058]), .A(rst), .Z(N1076) );
  ANDN U6107 ( .B(out[1059]), .A(rst), .Z(N1077) );
  ANDN U6108 ( .B(out[1060]), .A(rst), .Z(N1078) );
  ANDN U6109 ( .B(out[1061]), .A(rst), .Z(N1079) );
  ANDN U6110 ( .B(out[90]), .A(rst), .Z(N108) );
  ANDN U6111 ( .B(out[1062]), .A(rst), .Z(N1080) );
  ANDN U6112 ( .B(out[1063]), .A(rst), .Z(N1081) );
  ANDN U6113 ( .B(out[1064]), .A(rst), .Z(N1082) );
  ANDN U6114 ( .B(out[1065]), .A(rst), .Z(N1083) );
  ANDN U6115 ( .B(out[1066]), .A(rst), .Z(N1084) );
  ANDN U6116 ( .B(out[1067]), .A(rst), .Z(N1085) );
  ANDN U6117 ( .B(out[1068]), .A(rst), .Z(N1086) );
  ANDN U6118 ( .B(out[1069]), .A(rst), .Z(N1087) );
  ANDN U6119 ( .B(out[1070]), .A(rst), .Z(N1088) );
  ANDN U6120 ( .B(out[1071]), .A(rst), .Z(N1089) );
  ANDN U6121 ( .B(out[91]), .A(rst), .Z(N109) );
  ANDN U6122 ( .B(out[1072]), .A(rst), .Z(N1090) );
  ANDN U6123 ( .B(out[1073]), .A(rst), .Z(N1091) );
  ANDN U6124 ( .B(out[1074]), .A(rst), .Z(N1092) );
  ANDN U6125 ( .B(out[1075]), .A(rst), .Z(N1093) );
  ANDN U6126 ( .B(out[1076]), .A(rst), .Z(N1094) );
  ANDN U6127 ( .B(out[1077]), .A(rst), .Z(N1095) );
  ANDN U6128 ( .B(out[1078]), .A(rst), .Z(N1096) );
  ANDN U6129 ( .B(out[1079]), .A(rst), .Z(N1097) );
  ANDN U6130 ( .B(out[1080]), .A(rst), .Z(N1098) );
  ANDN U6131 ( .B(out[1081]), .A(rst), .Z(N1099) );
  ANDN U6132 ( .B(rc_i[4]), .A(rst), .Z(N11) );
  ANDN U6133 ( .B(out[92]), .A(rst), .Z(N110) );
  ANDN U6134 ( .B(out[1082]), .A(rst), .Z(N1100) );
  ANDN U6135 ( .B(out[1083]), .A(rst), .Z(N1101) );
  ANDN U6136 ( .B(out[1084]), .A(rst), .Z(N1102) );
  ANDN U6137 ( .B(out[1085]), .A(rst), .Z(N1103) );
  ANDN U6138 ( .B(out[1086]), .A(rst), .Z(N1104) );
  ANDN U6139 ( .B(out[1087]), .A(rst), .Z(N1105) );
  ANDN U6140 ( .B(out[1088]), .A(rst), .Z(N1106) );
  ANDN U6141 ( .B(out[1089]), .A(rst), .Z(N1107) );
  ANDN U6142 ( .B(out[1090]), .A(rst), .Z(N1108) );
  ANDN U6143 ( .B(out[1091]), .A(rst), .Z(N1109) );
  ANDN U6144 ( .B(out[93]), .A(rst), .Z(N111) );
  ANDN U6145 ( .B(out[1092]), .A(rst), .Z(N1110) );
  ANDN U6146 ( .B(out[1093]), .A(rst), .Z(N1111) );
  ANDN U6147 ( .B(out[1094]), .A(rst), .Z(N1112) );
  ANDN U6148 ( .B(out[1095]), .A(rst), .Z(N1113) );
  ANDN U6149 ( .B(out[1096]), .A(rst), .Z(N1114) );
  ANDN U6150 ( .B(out[1097]), .A(rst), .Z(N1115) );
  ANDN U6151 ( .B(out[1098]), .A(rst), .Z(N1116) );
  ANDN U6152 ( .B(out[1099]), .A(rst), .Z(N1117) );
  ANDN U6153 ( .B(out[1100]), .A(rst), .Z(N1118) );
  ANDN U6154 ( .B(out[1101]), .A(rst), .Z(N1119) );
  ANDN U6155 ( .B(out[94]), .A(rst), .Z(N112) );
  ANDN U6156 ( .B(out[1102]), .A(rst), .Z(N1120) );
  ANDN U6157 ( .B(out[1103]), .A(rst), .Z(N1121) );
  ANDN U6158 ( .B(out[1104]), .A(rst), .Z(N1122) );
  ANDN U6159 ( .B(out[1105]), .A(rst), .Z(N1123) );
  ANDN U6160 ( .B(out[1106]), .A(rst), .Z(N1124) );
  ANDN U6161 ( .B(out[1107]), .A(rst), .Z(N1125) );
  ANDN U6162 ( .B(out[1108]), .A(rst), .Z(N1126) );
  ANDN U6163 ( .B(out[1109]), .A(rst), .Z(N1127) );
  ANDN U6164 ( .B(out[1110]), .A(rst), .Z(N1128) );
  ANDN U6165 ( .B(out[1111]), .A(rst), .Z(N1129) );
  ANDN U6166 ( .B(out[95]), .A(rst), .Z(N113) );
  ANDN U6167 ( .B(out[1112]), .A(rst), .Z(N1130) );
  ANDN U6168 ( .B(out[1113]), .A(rst), .Z(N1131) );
  ANDN U6169 ( .B(out[1114]), .A(rst), .Z(N1132) );
  ANDN U6170 ( .B(out[1115]), .A(rst), .Z(N1133) );
  ANDN U6171 ( .B(out[1116]), .A(rst), .Z(N1134) );
  ANDN U6172 ( .B(out[1117]), .A(rst), .Z(N1135) );
  ANDN U6173 ( .B(out[1118]), .A(rst), .Z(N1136) );
  ANDN U6174 ( .B(out[1119]), .A(rst), .Z(N1137) );
  ANDN U6175 ( .B(out[1120]), .A(rst), .Z(N1138) );
  ANDN U6176 ( .B(out[1121]), .A(rst), .Z(N1139) );
  ANDN U6177 ( .B(out[96]), .A(rst), .Z(N114) );
  ANDN U6178 ( .B(out[1122]), .A(rst), .Z(N1140) );
  ANDN U6179 ( .B(out[1123]), .A(rst), .Z(N1141) );
  ANDN U6180 ( .B(out[1124]), .A(rst), .Z(N1142) );
  ANDN U6181 ( .B(out[1125]), .A(rst), .Z(N1143) );
  ANDN U6182 ( .B(out[1126]), .A(rst), .Z(N1144) );
  ANDN U6183 ( .B(out[1127]), .A(rst), .Z(N1145) );
  ANDN U6184 ( .B(out[1128]), .A(rst), .Z(N1146) );
  ANDN U6185 ( .B(out[1129]), .A(rst), .Z(N1147) );
  ANDN U6186 ( .B(out[1130]), .A(rst), .Z(N1148) );
  ANDN U6187 ( .B(out[1131]), .A(rst), .Z(N1149) );
  ANDN U6188 ( .B(out[97]), .A(rst), .Z(N115) );
  ANDN U6189 ( .B(out[1132]), .A(rst), .Z(N1150) );
  ANDN U6190 ( .B(out[1133]), .A(rst), .Z(N1151) );
  ANDN U6191 ( .B(out[1134]), .A(rst), .Z(N1152) );
  ANDN U6192 ( .B(out[1135]), .A(rst), .Z(N1153) );
  ANDN U6193 ( .B(out[1136]), .A(rst), .Z(N1154) );
  ANDN U6194 ( .B(out[1137]), .A(rst), .Z(N1155) );
  ANDN U6195 ( .B(out[1138]), .A(rst), .Z(N1156) );
  ANDN U6196 ( .B(out[1139]), .A(rst), .Z(N1157) );
  ANDN U6197 ( .B(out[1140]), .A(rst), .Z(N1158) );
  ANDN U6198 ( .B(out[1141]), .A(rst), .Z(N1159) );
  ANDN U6199 ( .B(out[98]), .A(rst), .Z(N116) );
  ANDN U6200 ( .B(out[1142]), .A(rst), .Z(N1160) );
  ANDN U6201 ( .B(out[1143]), .A(rst), .Z(N1161) );
  ANDN U6202 ( .B(out[1144]), .A(rst), .Z(N1162) );
  ANDN U6203 ( .B(out[1145]), .A(rst), .Z(N1163) );
  ANDN U6204 ( .B(out[1146]), .A(rst), .Z(N1164) );
  ANDN U6205 ( .B(out[1147]), .A(rst), .Z(N1165) );
  ANDN U6206 ( .B(out[1148]), .A(rst), .Z(N1166) );
  ANDN U6207 ( .B(out[1149]), .A(rst), .Z(N1167) );
  ANDN U6208 ( .B(out[1150]), .A(rst), .Z(N1168) );
  ANDN U6209 ( .B(out[1151]), .A(rst), .Z(N1169) );
  ANDN U6210 ( .B(out[99]), .A(rst), .Z(N117) );
  ANDN U6211 ( .B(out[1152]), .A(rst), .Z(N1170) );
  ANDN U6212 ( .B(out[1153]), .A(rst), .Z(N1171) );
  ANDN U6213 ( .B(out[1154]), .A(rst), .Z(N1172) );
  ANDN U6214 ( .B(out[1155]), .A(rst), .Z(N1173) );
  ANDN U6215 ( .B(out[1156]), .A(rst), .Z(N1174) );
  ANDN U6216 ( .B(out[1157]), .A(rst), .Z(N1175) );
  ANDN U6217 ( .B(out[1158]), .A(rst), .Z(N1176) );
  ANDN U6218 ( .B(out[1159]), .A(rst), .Z(N1177) );
  ANDN U6219 ( .B(out[1160]), .A(rst), .Z(N1178) );
  ANDN U6220 ( .B(out[1161]), .A(rst), .Z(N1179) );
  ANDN U6221 ( .B(out[100]), .A(rst), .Z(N118) );
  ANDN U6222 ( .B(out[1162]), .A(rst), .Z(N1180) );
  ANDN U6223 ( .B(out[1163]), .A(rst), .Z(N1181) );
  ANDN U6224 ( .B(out[1164]), .A(rst), .Z(N1182) );
  ANDN U6225 ( .B(out[1165]), .A(rst), .Z(N1183) );
  ANDN U6226 ( .B(out[1166]), .A(rst), .Z(N1184) );
  ANDN U6227 ( .B(out[1167]), .A(rst), .Z(N1185) );
  ANDN U6228 ( .B(out[1168]), .A(rst), .Z(N1186) );
  ANDN U6229 ( .B(out[1169]), .A(rst), .Z(N1187) );
  ANDN U6230 ( .B(out[1170]), .A(rst), .Z(N1188) );
  ANDN U6231 ( .B(out[1171]), .A(rst), .Z(N1189) );
  ANDN U6232 ( .B(out[101]), .A(rst), .Z(N119) );
  ANDN U6233 ( .B(out[1172]), .A(rst), .Z(N1190) );
  ANDN U6234 ( .B(out[1173]), .A(rst), .Z(N1191) );
  ANDN U6235 ( .B(out[1174]), .A(rst), .Z(N1192) );
  ANDN U6236 ( .B(out[1175]), .A(rst), .Z(N1193) );
  ANDN U6237 ( .B(out[1176]), .A(rst), .Z(N1194) );
  ANDN U6238 ( .B(out[1177]), .A(rst), .Z(N1195) );
  ANDN U6239 ( .B(out[1178]), .A(rst), .Z(N1196) );
  ANDN U6240 ( .B(out[1179]), .A(rst), .Z(N1197) );
  ANDN U6241 ( .B(out[1180]), .A(rst), .Z(N1198) );
  ANDN U6242 ( .B(out[1181]), .A(rst), .Z(N1199) );
  ANDN U6243 ( .B(rc_i[5]), .A(rst), .Z(N12) );
  ANDN U6244 ( .B(out[102]), .A(rst), .Z(N120) );
  ANDN U6245 ( .B(out[1182]), .A(rst), .Z(N1200) );
  ANDN U6246 ( .B(out[1183]), .A(rst), .Z(N1201) );
  ANDN U6247 ( .B(out[1184]), .A(rst), .Z(N1202) );
  ANDN U6248 ( .B(out[1185]), .A(rst), .Z(N1203) );
  ANDN U6249 ( .B(out[1186]), .A(rst), .Z(N1204) );
  ANDN U6250 ( .B(out[1187]), .A(rst), .Z(N1205) );
  ANDN U6251 ( .B(out[1188]), .A(rst), .Z(N1206) );
  ANDN U6252 ( .B(out[1189]), .A(rst), .Z(N1207) );
  ANDN U6253 ( .B(out[1190]), .A(rst), .Z(N1208) );
  ANDN U6254 ( .B(out[1191]), .A(rst), .Z(N1209) );
  ANDN U6255 ( .B(out[103]), .A(rst), .Z(N121) );
  ANDN U6256 ( .B(out[1192]), .A(rst), .Z(N1210) );
  ANDN U6257 ( .B(out[1193]), .A(rst), .Z(N1211) );
  ANDN U6258 ( .B(out[1194]), .A(rst), .Z(N1212) );
  ANDN U6259 ( .B(out[1195]), .A(rst), .Z(N1213) );
  ANDN U6260 ( .B(out[1196]), .A(rst), .Z(N1214) );
  ANDN U6261 ( .B(out[1197]), .A(rst), .Z(N1215) );
  ANDN U6262 ( .B(out[1198]), .A(rst), .Z(N1216) );
  ANDN U6263 ( .B(out[1199]), .A(rst), .Z(N1217) );
  ANDN U6264 ( .B(out[1200]), .A(rst), .Z(N1218) );
  ANDN U6265 ( .B(out[1201]), .A(rst), .Z(N1219) );
  ANDN U6266 ( .B(out[104]), .A(rst), .Z(N122) );
  ANDN U6267 ( .B(out[1202]), .A(rst), .Z(N1220) );
  ANDN U6268 ( .B(out[1203]), .A(rst), .Z(N1221) );
  ANDN U6269 ( .B(out[1204]), .A(rst), .Z(N1222) );
  ANDN U6270 ( .B(out[1205]), .A(rst), .Z(N1223) );
  ANDN U6271 ( .B(out[1206]), .A(rst), .Z(N1224) );
  ANDN U6272 ( .B(out[1207]), .A(rst), .Z(N1225) );
  ANDN U6273 ( .B(out[1208]), .A(rst), .Z(N1226) );
  ANDN U6274 ( .B(out[1209]), .A(rst), .Z(N1227) );
  ANDN U6275 ( .B(out[1210]), .A(rst), .Z(N1228) );
  ANDN U6276 ( .B(out[1211]), .A(rst), .Z(N1229) );
  ANDN U6277 ( .B(out[105]), .A(rst), .Z(N123) );
  ANDN U6278 ( .B(out[1212]), .A(rst), .Z(N1230) );
  ANDN U6279 ( .B(out[1213]), .A(rst), .Z(N1231) );
  ANDN U6280 ( .B(out[1214]), .A(rst), .Z(N1232) );
  ANDN U6281 ( .B(out[1215]), .A(rst), .Z(N1233) );
  ANDN U6282 ( .B(out[1216]), .A(rst), .Z(N1234) );
  ANDN U6283 ( .B(out[1217]), .A(rst), .Z(N1235) );
  ANDN U6284 ( .B(out[1218]), .A(rst), .Z(N1236) );
  ANDN U6285 ( .B(out[1219]), .A(rst), .Z(N1237) );
  ANDN U6286 ( .B(out[1220]), .A(rst), .Z(N1238) );
  ANDN U6287 ( .B(out[1221]), .A(rst), .Z(N1239) );
  ANDN U6288 ( .B(out[106]), .A(rst), .Z(N124) );
  ANDN U6289 ( .B(out[1222]), .A(rst), .Z(N1240) );
  ANDN U6290 ( .B(out[1223]), .A(rst), .Z(N1241) );
  ANDN U6291 ( .B(out[1224]), .A(rst), .Z(N1242) );
  ANDN U6292 ( .B(out[1225]), .A(rst), .Z(N1243) );
  ANDN U6293 ( .B(out[1226]), .A(rst), .Z(N1244) );
  ANDN U6294 ( .B(out[1227]), .A(rst), .Z(N1245) );
  ANDN U6295 ( .B(out[1228]), .A(rst), .Z(N1246) );
  ANDN U6296 ( .B(out[1229]), .A(rst), .Z(N1247) );
  ANDN U6297 ( .B(out[1230]), .A(rst), .Z(N1248) );
  ANDN U6298 ( .B(out[1231]), .A(rst), .Z(N1249) );
  ANDN U6299 ( .B(out[107]), .A(rst), .Z(N125) );
  ANDN U6300 ( .B(out[1232]), .A(rst), .Z(N1250) );
  ANDN U6301 ( .B(out[1233]), .A(rst), .Z(N1251) );
  ANDN U6302 ( .B(out[1234]), .A(rst), .Z(N1252) );
  ANDN U6303 ( .B(out[1235]), .A(rst), .Z(N1253) );
  ANDN U6304 ( .B(out[1236]), .A(rst), .Z(N1254) );
  ANDN U6305 ( .B(out[1237]), .A(rst), .Z(N1255) );
  ANDN U6306 ( .B(out[1238]), .A(rst), .Z(N1256) );
  ANDN U6307 ( .B(out[1239]), .A(rst), .Z(N1257) );
  ANDN U6308 ( .B(out[1240]), .A(rst), .Z(N1258) );
  ANDN U6309 ( .B(out[1241]), .A(rst), .Z(N1259) );
  ANDN U6310 ( .B(out[108]), .A(rst), .Z(N126) );
  ANDN U6311 ( .B(out[1242]), .A(rst), .Z(N1260) );
  ANDN U6312 ( .B(out[1243]), .A(rst), .Z(N1261) );
  ANDN U6313 ( .B(out[1244]), .A(rst), .Z(N1262) );
  ANDN U6314 ( .B(out[1245]), .A(rst), .Z(N1263) );
  ANDN U6315 ( .B(out[1246]), .A(rst), .Z(N1264) );
  ANDN U6316 ( .B(out[1247]), .A(rst), .Z(N1265) );
  ANDN U6317 ( .B(out[1248]), .A(rst), .Z(N1266) );
  ANDN U6318 ( .B(out[1249]), .A(rst), .Z(N1267) );
  ANDN U6319 ( .B(out[1250]), .A(rst), .Z(N1268) );
  ANDN U6320 ( .B(out[1251]), .A(rst), .Z(N1269) );
  ANDN U6321 ( .B(out[109]), .A(rst), .Z(N127) );
  ANDN U6322 ( .B(out[1252]), .A(rst), .Z(N1270) );
  ANDN U6323 ( .B(out[1253]), .A(rst), .Z(N1271) );
  ANDN U6324 ( .B(out[1254]), .A(rst), .Z(N1272) );
  ANDN U6325 ( .B(out[1255]), .A(rst), .Z(N1273) );
  ANDN U6326 ( .B(out[1256]), .A(rst), .Z(N1274) );
  ANDN U6327 ( .B(out[1257]), .A(rst), .Z(N1275) );
  ANDN U6328 ( .B(out[1258]), .A(rst), .Z(N1276) );
  ANDN U6329 ( .B(out[1259]), .A(rst), .Z(N1277) );
  ANDN U6330 ( .B(out[1260]), .A(rst), .Z(N1278) );
  ANDN U6331 ( .B(out[1261]), .A(rst), .Z(N1279) );
  ANDN U6332 ( .B(out[110]), .A(rst), .Z(N128) );
  ANDN U6333 ( .B(out[1262]), .A(rst), .Z(N1280) );
  ANDN U6334 ( .B(out[1263]), .A(rst), .Z(N1281) );
  ANDN U6335 ( .B(out[1264]), .A(rst), .Z(N1282) );
  ANDN U6336 ( .B(out[1265]), .A(rst), .Z(N1283) );
  ANDN U6337 ( .B(out[1266]), .A(rst), .Z(N1284) );
  ANDN U6338 ( .B(out[1267]), .A(rst), .Z(N1285) );
  ANDN U6339 ( .B(out[1268]), .A(rst), .Z(N1286) );
  ANDN U6340 ( .B(out[1269]), .A(rst), .Z(N1287) );
  ANDN U6341 ( .B(out[1270]), .A(rst), .Z(N1288) );
  ANDN U6342 ( .B(out[1271]), .A(rst), .Z(N1289) );
  ANDN U6343 ( .B(out[111]), .A(rst), .Z(N129) );
  ANDN U6344 ( .B(out[1272]), .A(rst), .Z(N1290) );
  ANDN U6345 ( .B(out[1273]), .A(rst), .Z(N1291) );
  ANDN U6346 ( .B(out[1274]), .A(rst), .Z(N1292) );
  ANDN U6347 ( .B(out[1275]), .A(rst), .Z(N1293) );
  ANDN U6348 ( .B(out[1276]), .A(rst), .Z(N1294) );
  ANDN U6349 ( .B(out[1277]), .A(rst), .Z(N1295) );
  ANDN U6350 ( .B(out[1278]), .A(rst), .Z(N1296) );
  ANDN U6351 ( .B(out[1279]), .A(rst), .Z(N1297) );
  ANDN U6352 ( .B(out[1280]), .A(rst), .Z(N1298) );
  ANDN U6353 ( .B(out[1281]), .A(rst), .Z(N1299) );
  ANDN U6354 ( .B(rc_i[6]), .A(rst), .Z(N13) );
  ANDN U6355 ( .B(out[112]), .A(rst), .Z(N130) );
  ANDN U6356 ( .B(out[1282]), .A(rst), .Z(N1300) );
  ANDN U6357 ( .B(out[1283]), .A(rst), .Z(N1301) );
  ANDN U6358 ( .B(out[1284]), .A(rst), .Z(N1302) );
  ANDN U6359 ( .B(out[1285]), .A(rst), .Z(N1303) );
  ANDN U6360 ( .B(out[1286]), .A(rst), .Z(N1304) );
  ANDN U6361 ( .B(out[1287]), .A(rst), .Z(N1305) );
  ANDN U6362 ( .B(out[1288]), .A(rst), .Z(N1306) );
  ANDN U6363 ( .B(out[1289]), .A(rst), .Z(N1307) );
  ANDN U6364 ( .B(out[1290]), .A(rst), .Z(N1308) );
  ANDN U6365 ( .B(out[1291]), .A(rst), .Z(N1309) );
  ANDN U6366 ( .B(out[113]), .A(rst), .Z(N131) );
  ANDN U6367 ( .B(out[1292]), .A(rst), .Z(N1310) );
  ANDN U6368 ( .B(out[1293]), .A(rst), .Z(N1311) );
  ANDN U6369 ( .B(out[1294]), .A(rst), .Z(N1312) );
  ANDN U6370 ( .B(out[1295]), .A(rst), .Z(N1313) );
  ANDN U6371 ( .B(out[1296]), .A(rst), .Z(N1314) );
  ANDN U6372 ( .B(out[1297]), .A(rst), .Z(N1315) );
  ANDN U6373 ( .B(out[1298]), .A(rst), .Z(N1316) );
  ANDN U6374 ( .B(out[1299]), .A(rst), .Z(N1317) );
  ANDN U6375 ( .B(out[1300]), .A(rst), .Z(N1318) );
  ANDN U6376 ( .B(out[1301]), .A(rst), .Z(N1319) );
  ANDN U6377 ( .B(out[114]), .A(rst), .Z(N132) );
  ANDN U6378 ( .B(out[1302]), .A(rst), .Z(N1320) );
  ANDN U6379 ( .B(out[1303]), .A(rst), .Z(N1321) );
  ANDN U6380 ( .B(out[1304]), .A(rst), .Z(N1322) );
  ANDN U6381 ( .B(out[1305]), .A(rst), .Z(N1323) );
  ANDN U6382 ( .B(out[1306]), .A(rst), .Z(N1324) );
  ANDN U6383 ( .B(out[1307]), .A(rst), .Z(N1325) );
  ANDN U6384 ( .B(out[1308]), .A(rst), .Z(N1326) );
  ANDN U6385 ( .B(out[1309]), .A(rst), .Z(N1327) );
  ANDN U6386 ( .B(out[1310]), .A(rst), .Z(N1328) );
  ANDN U6387 ( .B(out[1311]), .A(rst), .Z(N1329) );
  ANDN U6388 ( .B(out[115]), .A(rst), .Z(N133) );
  ANDN U6389 ( .B(out[1312]), .A(rst), .Z(N1330) );
  ANDN U6390 ( .B(out[1313]), .A(rst), .Z(N1331) );
  ANDN U6391 ( .B(out[1314]), .A(rst), .Z(N1332) );
  ANDN U6392 ( .B(out[1315]), .A(rst), .Z(N1333) );
  ANDN U6393 ( .B(out[1316]), .A(rst), .Z(N1334) );
  ANDN U6394 ( .B(out[1317]), .A(rst), .Z(N1335) );
  ANDN U6395 ( .B(out[1318]), .A(rst), .Z(N1336) );
  ANDN U6396 ( .B(out[1319]), .A(rst), .Z(N1337) );
  ANDN U6397 ( .B(out[1320]), .A(rst), .Z(N1338) );
  ANDN U6398 ( .B(out[1321]), .A(rst), .Z(N1339) );
  ANDN U6399 ( .B(out[116]), .A(rst), .Z(N134) );
  ANDN U6400 ( .B(out[1322]), .A(rst), .Z(N1340) );
  ANDN U6401 ( .B(out[1323]), .A(rst), .Z(N1341) );
  ANDN U6402 ( .B(out[1324]), .A(rst), .Z(N1342) );
  ANDN U6403 ( .B(out[1325]), .A(rst), .Z(N1343) );
  ANDN U6404 ( .B(out[1326]), .A(rst), .Z(N1344) );
  ANDN U6405 ( .B(out[1327]), .A(rst), .Z(N1345) );
  ANDN U6406 ( .B(out[1328]), .A(rst), .Z(N1346) );
  ANDN U6407 ( .B(out[1329]), .A(rst), .Z(N1347) );
  ANDN U6408 ( .B(out[1330]), .A(rst), .Z(N1348) );
  ANDN U6409 ( .B(out[1331]), .A(rst), .Z(N1349) );
  ANDN U6410 ( .B(out[117]), .A(rst), .Z(N135) );
  ANDN U6411 ( .B(out[1332]), .A(rst), .Z(N1350) );
  ANDN U6412 ( .B(out[1333]), .A(rst), .Z(N1351) );
  ANDN U6413 ( .B(out[1334]), .A(rst), .Z(N1352) );
  ANDN U6414 ( .B(out[1335]), .A(rst), .Z(N1353) );
  ANDN U6415 ( .B(out[1336]), .A(rst), .Z(N1354) );
  ANDN U6416 ( .B(out[1337]), .A(rst), .Z(N1355) );
  ANDN U6417 ( .B(out[1338]), .A(rst), .Z(N1356) );
  ANDN U6418 ( .B(out[1339]), .A(rst), .Z(N1357) );
  ANDN U6419 ( .B(out[1340]), .A(rst), .Z(N1358) );
  ANDN U6420 ( .B(out[1341]), .A(rst), .Z(N1359) );
  ANDN U6421 ( .B(out[118]), .A(rst), .Z(N136) );
  ANDN U6422 ( .B(out[1342]), .A(rst), .Z(N1360) );
  ANDN U6423 ( .B(out[1343]), .A(rst), .Z(N1361) );
  ANDN U6424 ( .B(out[1344]), .A(rst), .Z(N1362) );
  ANDN U6425 ( .B(out[1345]), .A(rst), .Z(N1363) );
  ANDN U6426 ( .B(out[1346]), .A(rst), .Z(N1364) );
  ANDN U6427 ( .B(out[1347]), .A(rst), .Z(N1365) );
  ANDN U6428 ( .B(out[1348]), .A(rst), .Z(N1366) );
  ANDN U6429 ( .B(out[1349]), .A(rst), .Z(N1367) );
  ANDN U6430 ( .B(out[1350]), .A(rst), .Z(N1368) );
  ANDN U6431 ( .B(out[1351]), .A(rst), .Z(N1369) );
  ANDN U6432 ( .B(out[119]), .A(rst), .Z(N137) );
  ANDN U6433 ( .B(out[1352]), .A(rst), .Z(N1370) );
  ANDN U6434 ( .B(out[1353]), .A(rst), .Z(N1371) );
  ANDN U6435 ( .B(out[1354]), .A(rst), .Z(N1372) );
  ANDN U6436 ( .B(out[1355]), .A(rst), .Z(N1373) );
  ANDN U6437 ( .B(out[1356]), .A(rst), .Z(N1374) );
  ANDN U6438 ( .B(out[1357]), .A(rst), .Z(N1375) );
  ANDN U6439 ( .B(out[1358]), .A(rst), .Z(N1376) );
  ANDN U6440 ( .B(out[1359]), .A(rst), .Z(N1377) );
  ANDN U6441 ( .B(out[1360]), .A(rst), .Z(N1378) );
  ANDN U6442 ( .B(out[1361]), .A(rst), .Z(N1379) );
  ANDN U6443 ( .B(out[120]), .A(rst), .Z(N138) );
  ANDN U6444 ( .B(out[1362]), .A(rst), .Z(N1380) );
  ANDN U6445 ( .B(out[1363]), .A(rst), .Z(N1381) );
  ANDN U6446 ( .B(out[1364]), .A(rst), .Z(N1382) );
  ANDN U6447 ( .B(out[1365]), .A(rst), .Z(N1383) );
  ANDN U6448 ( .B(out[1366]), .A(rst), .Z(N1384) );
  ANDN U6449 ( .B(out[1367]), .A(rst), .Z(N1385) );
  ANDN U6450 ( .B(out[1368]), .A(rst), .Z(N1386) );
  ANDN U6451 ( .B(out[1369]), .A(rst), .Z(N1387) );
  ANDN U6452 ( .B(out[1370]), .A(rst), .Z(N1388) );
  ANDN U6453 ( .B(out[1371]), .A(rst), .Z(N1389) );
  ANDN U6454 ( .B(out[121]), .A(rst), .Z(N139) );
  ANDN U6455 ( .B(out[1372]), .A(rst), .Z(N1390) );
  ANDN U6456 ( .B(out[1373]), .A(rst), .Z(N1391) );
  ANDN U6457 ( .B(out[1374]), .A(rst), .Z(N1392) );
  ANDN U6458 ( .B(out[1375]), .A(rst), .Z(N1393) );
  ANDN U6459 ( .B(out[1376]), .A(rst), .Z(N1394) );
  ANDN U6460 ( .B(out[1377]), .A(rst), .Z(N1395) );
  ANDN U6461 ( .B(out[1378]), .A(rst), .Z(N1396) );
  ANDN U6462 ( .B(out[1379]), .A(rst), .Z(N1397) );
  ANDN U6463 ( .B(out[1380]), .A(rst), .Z(N1398) );
  ANDN U6464 ( .B(out[1381]), .A(rst), .Z(N1399) );
  ANDN U6465 ( .B(rc_i[7]), .A(rst), .Z(N14) );
  ANDN U6466 ( .B(out[122]), .A(rst), .Z(N140) );
  ANDN U6467 ( .B(out[1382]), .A(rst), .Z(N1400) );
  ANDN U6468 ( .B(out[1383]), .A(rst), .Z(N1401) );
  ANDN U6469 ( .B(out[1384]), .A(rst), .Z(N1402) );
  ANDN U6470 ( .B(out[1385]), .A(rst), .Z(N1403) );
  ANDN U6471 ( .B(out[1386]), .A(rst), .Z(N1404) );
  ANDN U6472 ( .B(out[1387]), .A(rst), .Z(N1405) );
  ANDN U6473 ( .B(out[1388]), .A(rst), .Z(N1406) );
  ANDN U6474 ( .B(out[1389]), .A(rst), .Z(N1407) );
  ANDN U6475 ( .B(out[1390]), .A(rst), .Z(N1408) );
  ANDN U6476 ( .B(out[1391]), .A(rst), .Z(N1409) );
  ANDN U6477 ( .B(out[123]), .A(rst), .Z(N141) );
  ANDN U6478 ( .B(out[1392]), .A(rst), .Z(N1410) );
  ANDN U6479 ( .B(out[1393]), .A(rst), .Z(N1411) );
  ANDN U6480 ( .B(out[1394]), .A(rst), .Z(N1412) );
  ANDN U6481 ( .B(out[1395]), .A(rst), .Z(N1413) );
  ANDN U6482 ( .B(out[1396]), .A(rst), .Z(N1414) );
  ANDN U6483 ( .B(out[1397]), .A(rst), .Z(N1415) );
  ANDN U6484 ( .B(out[1398]), .A(rst), .Z(N1416) );
  ANDN U6485 ( .B(out[1399]), .A(rst), .Z(N1417) );
  ANDN U6486 ( .B(out[1400]), .A(rst), .Z(N1418) );
  ANDN U6487 ( .B(out[1401]), .A(rst), .Z(N1419) );
  ANDN U6488 ( .B(out[124]), .A(rst), .Z(N142) );
  ANDN U6489 ( .B(out[1402]), .A(rst), .Z(N1420) );
  ANDN U6490 ( .B(out[1403]), .A(rst), .Z(N1421) );
  ANDN U6491 ( .B(out[1404]), .A(rst), .Z(N1422) );
  ANDN U6492 ( .B(out[1405]), .A(rst), .Z(N1423) );
  ANDN U6493 ( .B(out[1406]), .A(rst), .Z(N1424) );
  ANDN U6494 ( .B(out[1407]), .A(rst), .Z(N1425) );
  ANDN U6495 ( .B(out[1408]), .A(rst), .Z(N1426) );
  ANDN U6496 ( .B(out[1409]), .A(rst), .Z(N1427) );
  ANDN U6497 ( .B(out[1410]), .A(rst), .Z(N1428) );
  ANDN U6498 ( .B(out[1411]), .A(rst), .Z(N1429) );
  ANDN U6499 ( .B(out[125]), .A(rst), .Z(N143) );
  ANDN U6500 ( .B(out[1412]), .A(rst), .Z(N1430) );
  ANDN U6501 ( .B(out[1413]), .A(rst), .Z(N1431) );
  ANDN U6502 ( .B(out[1414]), .A(rst), .Z(N1432) );
  ANDN U6503 ( .B(out[1415]), .A(rst), .Z(N1433) );
  ANDN U6504 ( .B(out[1416]), .A(rst), .Z(N1434) );
  ANDN U6505 ( .B(out[1417]), .A(rst), .Z(N1435) );
  ANDN U6506 ( .B(out[1418]), .A(rst), .Z(N1436) );
  ANDN U6507 ( .B(out[1419]), .A(rst), .Z(N1437) );
  ANDN U6508 ( .B(out[1420]), .A(rst), .Z(N1438) );
  ANDN U6509 ( .B(out[1421]), .A(rst), .Z(N1439) );
  ANDN U6510 ( .B(out[126]), .A(rst), .Z(N144) );
  ANDN U6511 ( .B(out[1422]), .A(rst), .Z(N1440) );
  ANDN U6512 ( .B(out[1423]), .A(rst), .Z(N1441) );
  ANDN U6513 ( .B(out[1424]), .A(rst), .Z(N1442) );
  ANDN U6514 ( .B(out[1425]), .A(rst), .Z(N1443) );
  ANDN U6515 ( .B(out[1426]), .A(rst), .Z(N1444) );
  ANDN U6516 ( .B(out[1427]), .A(rst), .Z(N1445) );
  ANDN U6517 ( .B(out[1428]), .A(rst), .Z(N1446) );
  ANDN U6518 ( .B(out[1429]), .A(rst), .Z(N1447) );
  ANDN U6519 ( .B(out[1430]), .A(rst), .Z(N1448) );
  ANDN U6520 ( .B(out[1431]), .A(rst), .Z(N1449) );
  ANDN U6521 ( .B(out[127]), .A(rst), .Z(N145) );
  ANDN U6522 ( .B(out[1432]), .A(rst), .Z(N1450) );
  ANDN U6523 ( .B(out[1433]), .A(rst), .Z(N1451) );
  ANDN U6524 ( .B(out[1434]), .A(rst), .Z(N1452) );
  ANDN U6525 ( .B(out[1435]), .A(rst), .Z(N1453) );
  ANDN U6526 ( .B(out[1436]), .A(rst), .Z(N1454) );
  ANDN U6527 ( .B(out[1437]), .A(rst), .Z(N1455) );
  ANDN U6528 ( .B(out[1438]), .A(rst), .Z(N1456) );
  ANDN U6529 ( .B(out[1439]), .A(rst), .Z(N1457) );
  ANDN U6530 ( .B(out[1440]), .A(rst), .Z(N1458) );
  ANDN U6531 ( .B(out[1441]), .A(rst), .Z(N1459) );
  ANDN U6532 ( .B(out[128]), .A(rst), .Z(N146) );
  ANDN U6533 ( .B(out[1442]), .A(rst), .Z(N1460) );
  ANDN U6534 ( .B(out[1443]), .A(rst), .Z(N1461) );
  ANDN U6535 ( .B(out[1444]), .A(rst), .Z(N1462) );
  ANDN U6536 ( .B(out[1445]), .A(rst), .Z(N1463) );
  ANDN U6537 ( .B(out[1446]), .A(rst), .Z(N1464) );
  ANDN U6538 ( .B(out[1447]), .A(rst), .Z(N1465) );
  ANDN U6539 ( .B(out[1448]), .A(rst), .Z(N1466) );
  ANDN U6540 ( .B(out[1449]), .A(rst), .Z(N1467) );
  ANDN U6541 ( .B(out[1450]), .A(rst), .Z(N1468) );
  ANDN U6542 ( .B(out[1451]), .A(rst), .Z(N1469) );
  ANDN U6543 ( .B(out[129]), .A(rst), .Z(N147) );
  ANDN U6544 ( .B(out[1452]), .A(rst), .Z(N1470) );
  ANDN U6545 ( .B(out[1453]), .A(rst), .Z(N1471) );
  ANDN U6546 ( .B(out[1454]), .A(rst), .Z(N1472) );
  ANDN U6547 ( .B(out[1455]), .A(rst), .Z(N1473) );
  ANDN U6548 ( .B(out[1456]), .A(rst), .Z(N1474) );
  ANDN U6549 ( .B(out[1457]), .A(rst), .Z(N1475) );
  ANDN U6550 ( .B(out[1458]), .A(rst), .Z(N1476) );
  ANDN U6551 ( .B(out[1459]), .A(rst), .Z(N1477) );
  ANDN U6552 ( .B(out[1460]), .A(rst), .Z(N1478) );
  ANDN U6553 ( .B(out[1461]), .A(rst), .Z(N1479) );
  ANDN U6554 ( .B(out[130]), .A(rst), .Z(N148) );
  ANDN U6555 ( .B(out[1462]), .A(rst), .Z(N1480) );
  ANDN U6556 ( .B(out[1463]), .A(rst), .Z(N1481) );
  ANDN U6557 ( .B(out[1464]), .A(rst), .Z(N1482) );
  ANDN U6558 ( .B(out[1465]), .A(rst), .Z(N1483) );
  ANDN U6559 ( .B(out[1466]), .A(rst), .Z(N1484) );
  ANDN U6560 ( .B(out[1467]), .A(rst), .Z(N1485) );
  ANDN U6561 ( .B(out[1468]), .A(rst), .Z(N1486) );
  ANDN U6562 ( .B(out[1469]), .A(rst), .Z(N1487) );
  ANDN U6563 ( .B(out[1470]), .A(rst), .Z(N1488) );
  ANDN U6564 ( .B(out[1471]), .A(rst), .Z(N1489) );
  ANDN U6565 ( .B(out[131]), .A(rst), .Z(N149) );
  ANDN U6566 ( .B(out[1472]), .A(rst), .Z(N1490) );
  ANDN U6567 ( .B(out[1473]), .A(rst), .Z(N1491) );
  ANDN U6568 ( .B(out[1474]), .A(rst), .Z(N1492) );
  ANDN U6569 ( .B(out[1475]), .A(rst), .Z(N1493) );
  ANDN U6570 ( .B(out[1476]), .A(rst), .Z(N1494) );
  ANDN U6571 ( .B(out[1477]), .A(rst), .Z(N1495) );
  ANDN U6572 ( .B(out[1478]), .A(rst), .Z(N1496) );
  ANDN U6573 ( .B(out[1479]), .A(rst), .Z(N1497) );
  ANDN U6574 ( .B(out[1480]), .A(rst), .Z(N1498) );
  ANDN U6575 ( .B(out[1481]), .A(rst), .Z(N1499) );
  ANDN U6576 ( .B(rc_i[8]), .A(rst), .Z(N15) );
  ANDN U6577 ( .B(out[132]), .A(rst), .Z(N150) );
  ANDN U6578 ( .B(out[1482]), .A(rst), .Z(N1500) );
  ANDN U6579 ( .B(out[1483]), .A(rst), .Z(N1501) );
  ANDN U6580 ( .B(out[1484]), .A(rst), .Z(N1502) );
  ANDN U6581 ( .B(out[1485]), .A(rst), .Z(N1503) );
  ANDN U6582 ( .B(out[1486]), .A(rst), .Z(N1504) );
  ANDN U6583 ( .B(out[1487]), .A(rst), .Z(N1505) );
  ANDN U6584 ( .B(out[1488]), .A(rst), .Z(N1506) );
  ANDN U6585 ( .B(out[1489]), .A(rst), .Z(N1507) );
  ANDN U6586 ( .B(out[1490]), .A(rst), .Z(N1508) );
  ANDN U6587 ( .B(out[1491]), .A(rst), .Z(N1509) );
  ANDN U6588 ( .B(out[133]), .A(rst), .Z(N151) );
  ANDN U6589 ( .B(out[1492]), .A(rst), .Z(N1510) );
  ANDN U6590 ( .B(out[1493]), .A(rst), .Z(N1511) );
  ANDN U6591 ( .B(out[1494]), .A(rst), .Z(N1512) );
  ANDN U6592 ( .B(out[1495]), .A(rst), .Z(N1513) );
  ANDN U6593 ( .B(out[1496]), .A(rst), .Z(N1514) );
  ANDN U6594 ( .B(out[1497]), .A(rst), .Z(N1515) );
  ANDN U6595 ( .B(out[1498]), .A(rst), .Z(N1516) );
  ANDN U6596 ( .B(out[1499]), .A(rst), .Z(N1517) );
  ANDN U6597 ( .B(out[1500]), .A(rst), .Z(N1518) );
  ANDN U6598 ( .B(out[1501]), .A(rst), .Z(N1519) );
  ANDN U6599 ( .B(out[134]), .A(rst), .Z(N152) );
  ANDN U6600 ( .B(out[1502]), .A(rst), .Z(N1520) );
  ANDN U6601 ( .B(out[1503]), .A(rst), .Z(N1521) );
  ANDN U6602 ( .B(out[1504]), .A(rst), .Z(N1522) );
  ANDN U6603 ( .B(out[1505]), .A(rst), .Z(N1523) );
  ANDN U6604 ( .B(out[1506]), .A(rst), .Z(N1524) );
  ANDN U6605 ( .B(out[1507]), .A(rst), .Z(N1525) );
  ANDN U6606 ( .B(out[1508]), .A(rst), .Z(N1526) );
  ANDN U6607 ( .B(out[1509]), .A(rst), .Z(N1527) );
  ANDN U6608 ( .B(out[1510]), .A(rst), .Z(N1528) );
  ANDN U6609 ( .B(out[1511]), .A(rst), .Z(N1529) );
  ANDN U6610 ( .B(out[135]), .A(rst), .Z(N153) );
  ANDN U6611 ( .B(out[1512]), .A(rst), .Z(N1530) );
  ANDN U6612 ( .B(out[1513]), .A(rst), .Z(N1531) );
  ANDN U6613 ( .B(out[1514]), .A(rst), .Z(N1532) );
  ANDN U6614 ( .B(out[1515]), .A(rst), .Z(N1533) );
  ANDN U6615 ( .B(out[1516]), .A(rst), .Z(N1534) );
  ANDN U6616 ( .B(out[1517]), .A(rst), .Z(N1535) );
  ANDN U6617 ( .B(out[1518]), .A(rst), .Z(N1536) );
  ANDN U6618 ( .B(out[1519]), .A(rst), .Z(N1537) );
  ANDN U6619 ( .B(out[1520]), .A(rst), .Z(N1538) );
  ANDN U6620 ( .B(out[1521]), .A(rst), .Z(N1539) );
  ANDN U6621 ( .B(out[136]), .A(rst), .Z(N154) );
  ANDN U6622 ( .B(out[1522]), .A(rst), .Z(N1540) );
  ANDN U6623 ( .B(out[1523]), .A(rst), .Z(N1541) );
  ANDN U6624 ( .B(out[1524]), .A(rst), .Z(N1542) );
  ANDN U6625 ( .B(out[1525]), .A(rst), .Z(N1543) );
  ANDN U6626 ( .B(out[1526]), .A(rst), .Z(N1544) );
  ANDN U6627 ( .B(out[1527]), .A(rst), .Z(N1545) );
  ANDN U6628 ( .B(out[1528]), .A(rst), .Z(N1546) );
  ANDN U6629 ( .B(out[1529]), .A(rst), .Z(N1547) );
  ANDN U6630 ( .B(out[1530]), .A(rst), .Z(N1548) );
  ANDN U6631 ( .B(out[1531]), .A(rst), .Z(N1549) );
  ANDN U6632 ( .B(out[137]), .A(rst), .Z(N155) );
  ANDN U6633 ( .B(out[1532]), .A(rst), .Z(N1550) );
  ANDN U6634 ( .B(out[1533]), .A(rst), .Z(N1551) );
  ANDN U6635 ( .B(out[1534]), .A(rst), .Z(N1552) );
  ANDN U6636 ( .B(out[1535]), .A(rst), .Z(N1553) );
  ANDN U6637 ( .B(out[1536]), .A(rst), .Z(N1554) );
  ANDN U6638 ( .B(out[1537]), .A(rst), .Z(N1555) );
  ANDN U6639 ( .B(out[1538]), .A(rst), .Z(N1556) );
  ANDN U6640 ( .B(out[1539]), .A(rst), .Z(N1557) );
  ANDN U6641 ( .B(out[1540]), .A(rst), .Z(N1558) );
  ANDN U6642 ( .B(out[1541]), .A(rst), .Z(N1559) );
  ANDN U6643 ( .B(out[138]), .A(rst), .Z(N156) );
  ANDN U6644 ( .B(out[1542]), .A(rst), .Z(N1560) );
  ANDN U6645 ( .B(out[1543]), .A(rst), .Z(N1561) );
  ANDN U6646 ( .B(out[1544]), .A(rst), .Z(N1562) );
  ANDN U6647 ( .B(out[1545]), .A(rst), .Z(N1563) );
  ANDN U6648 ( .B(out[1546]), .A(rst), .Z(N1564) );
  ANDN U6649 ( .B(out[1547]), .A(rst), .Z(N1565) );
  ANDN U6650 ( .B(out[1548]), .A(rst), .Z(N1566) );
  ANDN U6651 ( .B(out[1549]), .A(rst), .Z(N1567) );
  ANDN U6652 ( .B(out[1550]), .A(rst), .Z(N1568) );
  ANDN U6653 ( .B(out[1551]), .A(rst), .Z(N1569) );
  ANDN U6654 ( .B(out[139]), .A(rst), .Z(N157) );
  ANDN U6655 ( .B(out[1552]), .A(rst), .Z(N1570) );
  ANDN U6656 ( .B(out[1553]), .A(rst), .Z(N1571) );
  ANDN U6657 ( .B(out[1554]), .A(rst), .Z(N1572) );
  ANDN U6658 ( .B(out[1555]), .A(rst), .Z(N1573) );
  ANDN U6659 ( .B(out[1556]), .A(rst), .Z(N1574) );
  ANDN U6660 ( .B(out[1557]), .A(rst), .Z(N1575) );
  ANDN U6661 ( .B(out[1558]), .A(rst), .Z(N1576) );
  ANDN U6662 ( .B(out[1559]), .A(rst), .Z(N1577) );
  ANDN U6663 ( .B(out[1560]), .A(rst), .Z(N1578) );
  ANDN U6664 ( .B(out[1561]), .A(rst), .Z(N1579) );
  ANDN U6665 ( .B(out[140]), .A(rst), .Z(N158) );
  ANDN U6666 ( .B(out[1562]), .A(rst), .Z(N1580) );
  ANDN U6667 ( .B(out[1563]), .A(rst), .Z(N1581) );
  ANDN U6668 ( .B(out[1564]), .A(rst), .Z(N1582) );
  ANDN U6669 ( .B(out[1565]), .A(rst), .Z(N1583) );
  ANDN U6670 ( .B(out[1566]), .A(rst), .Z(N1584) );
  ANDN U6671 ( .B(out[1567]), .A(rst), .Z(N1585) );
  ANDN U6672 ( .B(out[1568]), .A(rst), .Z(N1586) );
  ANDN U6673 ( .B(out[1569]), .A(rst), .Z(N1587) );
  ANDN U6674 ( .B(out[1570]), .A(rst), .Z(N1588) );
  ANDN U6675 ( .B(out[1571]), .A(rst), .Z(N1589) );
  ANDN U6676 ( .B(out[141]), .A(rst), .Z(N159) );
  ANDN U6677 ( .B(out[1572]), .A(rst), .Z(N1590) );
  ANDN U6678 ( .B(out[1573]), .A(rst), .Z(N1591) );
  ANDN U6679 ( .B(out[1574]), .A(rst), .Z(N1592) );
  ANDN U6680 ( .B(out[1575]), .A(rst), .Z(N1593) );
  ANDN U6681 ( .B(out[1576]), .A(rst), .Z(N1594) );
  ANDN U6682 ( .B(out[1577]), .A(rst), .Z(N1595) );
  ANDN U6683 ( .B(out[1578]), .A(rst), .Z(N1596) );
  ANDN U6684 ( .B(out[1579]), .A(rst), .Z(N1597) );
  ANDN U6685 ( .B(out[1580]), .A(rst), .Z(N1598) );
  ANDN U6686 ( .B(out[1581]), .A(rst), .Z(N1599) );
  ANDN U6687 ( .B(rc_i[9]), .A(rst), .Z(N16) );
  ANDN U6688 ( .B(out[142]), .A(rst), .Z(N160) );
  ANDN U6689 ( .B(out[1582]), .A(rst), .Z(N1600) );
  ANDN U6690 ( .B(out[1583]), .A(rst), .Z(N1601) );
  ANDN U6691 ( .B(out[1584]), .A(rst), .Z(N1602) );
  ANDN U6692 ( .B(out[1585]), .A(rst), .Z(N1603) );
  ANDN U6693 ( .B(out[1586]), .A(rst), .Z(N1604) );
  ANDN U6694 ( .B(out[1587]), .A(rst), .Z(N1605) );
  ANDN U6695 ( .B(out[1588]), .A(rst), .Z(N1606) );
  ANDN U6696 ( .B(out[1589]), .A(rst), .Z(N1607) );
  ANDN U6697 ( .B(out[1590]), .A(rst), .Z(N1608) );
  ANDN U6698 ( .B(out[1591]), .A(rst), .Z(N1609) );
  ANDN U6699 ( .B(out[143]), .A(rst), .Z(N161) );
  ANDN U6700 ( .B(out[1592]), .A(rst), .Z(N1610) );
  ANDN U6701 ( .B(out[1593]), .A(rst), .Z(N1611) );
  ANDN U6702 ( .B(out[1594]), .A(rst), .Z(N1612) );
  ANDN U6703 ( .B(out[1595]), .A(rst), .Z(N1613) );
  ANDN U6704 ( .B(out[1596]), .A(rst), .Z(N1614) );
  ANDN U6705 ( .B(out[1597]), .A(rst), .Z(N1615) );
  ANDN U6706 ( .B(out[1598]), .A(rst), .Z(N1616) );
  ANDN U6707 ( .B(out[1599]), .A(rst), .Z(N1617) );
  ANDN U6708 ( .B(out[144]), .A(rst), .Z(N162) );
  ANDN U6709 ( .B(out[145]), .A(rst), .Z(N163) );
  ANDN U6710 ( .B(out[146]), .A(rst), .Z(N164) );
  ANDN U6711 ( .B(out[147]), .A(rst), .Z(N165) );
  ANDN U6712 ( .B(out[148]), .A(rst), .Z(N166) );
  ANDN U6713 ( .B(out[149]), .A(rst), .Z(N167) );
  ANDN U6714 ( .B(out[150]), .A(rst), .Z(N168) );
  ANDN U6715 ( .B(out[151]), .A(rst), .Z(N169) );
  ANDN U6716 ( .B(rc_i[10]), .A(rst), .Z(N17) );
  ANDN U6717 ( .B(out[152]), .A(rst), .Z(N170) );
  ANDN U6718 ( .B(out[153]), .A(rst), .Z(N171) );
  ANDN U6719 ( .B(out[154]), .A(rst), .Z(N172) );
  ANDN U6720 ( .B(out[155]), .A(rst), .Z(N173) );
  ANDN U6721 ( .B(out[156]), .A(rst), .Z(N174) );
  ANDN U6722 ( .B(out[157]), .A(rst), .Z(N175) );
  ANDN U6723 ( .B(out[158]), .A(rst), .Z(N176) );
  ANDN U6724 ( .B(out[159]), .A(rst), .Z(N177) );
  ANDN U6725 ( .B(out[160]), .A(rst), .Z(N178) );
  ANDN U6726 ( .B(out[161]), .A(rst), .Z(N179) );
  ANDN U6727 ( .B(out[0]), .A(rst), .Z(N18) );
  ANDN U6728 ( .B(out[162]), .A(rst), .Z(N180) );
  ANDN U6729 ( .B(out[163]), .A(rst), .Z(N181) );
  ANDN U6730 ( .B(out[164]), .A(rst), .Z(N182) );
  ANDN U6731 ( .B(out[165]), .A(rst), .Z(N183) );
  ANDN U6732 ( .B(out[166]), .A(rst), .Z(N184) );
  ANDN U6733 ( .B(out[167]), .A(rst), .Z(N185) );
  ANDN U6734 ( .B(out[168]), .A(rst), .Z(N186) );
  ANDN U6735 ( .B(out[169]), .A(rst), .Z(N187) );
  ANDN U6736 ( .B(out[170]), .A(rst), .Z(N188) );
  ANDN U6737 ( .B(out[171]), .A(rst), .Z(N189) );
  ANDN U6738 ( .B(out[1]), .A(rst), .Z(N19) );
  ANDN U6739 ( .B(out[172]), .A(rst), .Z(N190) );
  ANDN U6740 ( .B(out[173]), .A(rst), .Z(N191) );
  ANDN U6741 ( .B(out[174]), .A(rst), .Z(N192) );
  ANDN U6742 ( .B(out[175]), .A(rst), .Z(N193) );
  ANDN U6743 ( .B(out[176]), .A(rst), .Z(N194) );
  ANDN U6744 ( .B(out[177]), .A(rst), .Z(N195) );
  ANDN U6745 ( .B(out[178]), .A(rst), .Z(N196) );
  ANDN U6746 ( .B(out[179]), .A(rst), .Z(N197) );
  ANDN U6747 ( .B(out[180]), .A(rst), .Z(N198) );
  ANDN U6748 ( .B(out[181]), .A(rst), .Z(N199) );
  ANDN U6749 ( .B(out[2]), .A(rst), .Z(N20) );
  ANDN U6750 ( .B(out[182]), .A(rst), .Z(N200) );
  ANDN U6751 ( .B(out[183]), .A(rst), .Z(N201) );
  ANDN U6752 ( .B(out[184]), .A(rst), .Z(N202) );
  ANDN U6753 ( .B(out[185]), .A(rst), .Z(N203) );
  ANDN U6754 ( .B(out[186]), .A(rst), .Z(N204) );
  ANDN U6755 ( .B(out[187]), .A(rst), .Z(N205) );
  ANDN U6756 ( .B(out[188]), .A(rst), .Z(N206) );
  ANDN U6757 ( .B(out[189]), .A(rst), .Z(N207) );
  ANDN U6758 ( .B(out[190]), .A(rst), .Z(N208) );
  ANDN U6759 ( .B(out[191]), .A(rst), .Z(N209) );
  ANDN U6760 ( .B(out[3]), .A(rst), .Z(N21) );
  ANDN U6761 ( .B(out[192]), .A(rst), .Z(N210) );
  ANDN U6762 ( .B(out[193]), .A(rst), .Z(N211) );
  ANDN U6763 ( .B(out[194]), .A(rst), .Z(N212) );
  ANDN U6764 ( .B(out[195]), .A(rst), .Z(N213) );
  ANDN U6765 ( .B(out[196]), .A(rst), .Z(N214) );
  ANDN U6766 ( .B(out[197]), .A(rst), .Z(N215) );
  ANDN U6767 ( .B(out[198]), .A(rst), .Z(N216) );
  ANDN U6768 ( .B(out[199]), .A(rst), .Z(N217) );
  ANDN U6769 ( .B(out[200]), .A(rst), .Z(N218) );
  ANDN U6770 ( .B(out[201]), .A(rst), .Z(N219) );
  ANDN U6771 ( .B(out[4]), .A(rst), .Z(N22) );
  ANDN U6772 ( .B(out[202]), .A(rst), .Z(N220) );
  ANDN U6773 ( .B(out[203]), .A(rst), .Z(N221) );
  ANDN U6774 ( .B(out[204]), .A(rst), .Z(N222) );
  ANDN U6775 ( .B(out[205]), .A(rst), .Z(N223) );
  ANDN U6776 ( .B(out[206]), .A(rst), .Z(N224) );
  ANDN U6777 ( .B(out[207]), .A(rst), .Z(N225) );
  ANDN U6778 ( .B(out[208]), .A(rst), .Z(N226) );
  ANDN U6779 ( .B(out[209]), .A(rst), .Z(N227) );
  ANDN U6780 ( .B(out[210]), .A(rst), .Z(N228) );
  ANDN U6781 ( .B(out[211]), .A(rst), .Z(N229) );
  ANDN U6782 ( .B(out[5]), .A(rst), .Z(N23) );
  ANDN U6783 ( .B(out[212]), .A(rst), .Z(N230) );
  ANDN U6784 ( .B(out[213]), .A(rst), .Z(N231) );
  ANDN U6785 ( .B(out[214]), .A(rst), .Z(N232) );
  ANDN U6786 ( .B(out[215]), .A(rst), .Z(N233) );
  ANDN U6787 ( .B(out[216]), .A(rst), .Z(N234) );
  ANDN U6788 ( .B(out[217]), .A(rst), .Z(N235) );
  ANDN U6789 ( .B(out[218]), .A(rst), .Z(N236) );
  ANDN U6790 ( .B(out[219]), .A(rst), .Z(N237) );
  ANDN U6791 ( .B(out[220]), .A(rst), .Z(N238) );
  ANDN U6792 ( .B(out[221]), .A(rst), .Z(N239) );
  ANDN U6793 ( .B(out[6]), .A(rst), .Z(N24) );
  ANDN U6794 ( .B(out[222]), .A(rst), .Z(N240) );
  ANDN U6795 ( .B(out[223]), .A(rst), .Z(N241) );
  ANDN U6796 ( .B(out[224]), .A(rst), .Z(N242) );
  ANDN U6797 ( .B(out[225]), .A(rst), .Z(N243) );
  ANDN U6798 ( .B(out[226]), .A(rst), .Z(N244) );
  ANDN U6799 ( .B(out[227]), .A(rst), .Z(N245) );
  ANDN U6800 ( .B(out[228]), .A(rst), .Z(N246) );
  ANDN U6801 ( .B(out[229]), .A(rst), .Z(N247) );
  ANDN U6802 ( .B(out[230]), .A(rst), .Z(N248) );
  ANDN U6803 ( .B(out[231]), .A(rst), .Z(N249) );
  ANDN U6804 ( .B(out[7]), .A(rst), .Z(N25) );
  ANDN U6805 ( .B(out[232]), .A(rst), .Z(N250) );
  ANDN U6806 ( .B(out[233]), .A(rst), .Z(N251) );
  ANDN U6807 ( .B(out[234]), .A(rst), .Z(N252) );
  ANDN U6808 ( .B(out[235]), .A(rst), .Z(N253) );
  ANDN U6809 ( .B(out[236]), .A(rst), .Z(N254) );
  ANDN U6810 ( .B(out[237]), .A(rst), .Z(N255) );
  ANDN U6811 ( .B(out[238]), .A(rst), .Z(N256) );
  ANDN U6812 ( .B(out[239]), .A(rst), .Z(N257) );
  ANDN U6813 ( .B(out[240]), .A(rst), .Z(N258) );
  ANDN U6814 ( .B(out[241]), .A(rst), .Z(N259) );
  ANDN U6815 ( .B(out[8]), .A(rst), .Z(N26) );
  ANDN U6816 ( .B(out[242]), .A(rst), .Z(N260) );
  ANDN U6817 ( .B(out[243]), .A(rst), .Z(N261) );
  ANDN U6818 ( .B(out[244]), .A(rst), .Z(N262) );
  ANDN U6819 ( .B(out[245]), .A(rst), .Z(N263) );
  ANDN U6820 ( .B(out[246]), .A(rst), .Z(N264) );
  ANDN U6821 ( .B(out[247]), .A(rst), .Z(N265) );
  ANDN U6822 ( .B(out[248]), .A(rst), .Z(N266) );
  ANDN U6823 ( .B(out[249]), .A(rst), .Z(N267) );
  ANDN U6824 ( .B(out[250]), .A(rst), .Z(N268) );
  ANDN U6825 ( .B(out[251]), .A(rst), .Z(N269) );
  ANDN U6826 ( .B(out[9]), .A(rst), .Z(N27) );
  ANDN U6827 ( .B(out[252]), .A(rst), .Z(N270) );
  ANDN U6828 ( .B(out[253]), .A(rst), .Z(N271) );
  ANDN U6829 ( .B(out[254]), .A(rst), .Z(N272) );
  ANDN U6830 ( .B(out[255]), .A(rst), .Z(N273) );
  ANDN U6831 ( .B(out[256]), .A(rst), .Z(N274) );
  ANDN U6832 ( .B(out[257]), .A(rst), .Z(N275) );
  ANDN U6833 ( .B(out[258]), .A(rst), .Z(N276) );
  ANDN U6834 ( .B(out[259]), .A(rst), .Z(N277) );
  ANDN U6835 ( .B(out[260]), .A(rst), .Z(N278) );
  ANDN U6836 ( .B(out[261]), .A(rst), .Z(N279) );
  ANDN U6837 ( .B(out[10]), .A(rst), .Z(N28) );
  ANDN U6838 ( .B(out[262]), .A(rst), .Z(N280) );
  ANDN U6839 ( .B(out[263]), .A(rst), .Z(N281) );
  ANDN U6840 ( .B(out[264]), .A(rst), .Z(N282) );
  ANDN U6841 ( .B(out[265]), .A(rst), .Z(N283) );
  ANDN U6842 ( .B(out[266]), .A(rst), .Z(N284) );
  ANDN U6843 ( .B(out[267]), .A(rst), .Z(N285) );
  ANDN U6844 ( .B(out[268]), .A(rst), .Z(N286) );
  ANDN U6845 ( .B(out[269]), .A(rst), .Z(N287) );
  ANDN U6846 ( .B(out[270]), .A(rst), .Z(N288) );
  ANDN U6847 ( .B(out[271]), .A(rst), .Z(N289) );
  ANDN U6848 ( .B(out[11]), .A(rst), .Z(N29) );
  ANDN U6849 ( .B(out[272]), .A(rst), .Z(N290) );
  ANDN U6850 ( .B(out[273]), .A(rst), .Z(N291) );
  ANDN U6851 ( .B(out[274]), .A(rst), .Z(N292) );
  ANDN U6852 ( .B(out[275]), .A(rst), .Z(N293) );
  ANDN U6853 ( .B(out[276]), .A(rst), .Z(N294) );
  ANDN U6854 ( .B(out[277]), .A(rst), .Z(N295) );
  ANDN U6855 ( .B(out[278]), .A(rst), .Z(N296) );
  ANDN U6856 ( .B(out[279]), .A(rst), .Z(N297) );
  ANDN U6857 ( .B(out[280]), .A(rst), .Z(N298) );
  ANDN U6858 ( .B(out[281]), .A(rst), .Z(N299) );
  ANDN U6859 ( .B(out[12]), .A(rst), .Z(N30) );
  ANDN U6860 ( .B(out[282]), .A(rst), .Z(N300) );
  ANDN U6861 ( .B(out[283]), .A(rst), .Z(N301) );
  ANDN U6862 ( .B(out[284]), .A(rst), .Z(N302) );
  ANDN U6863 ( .B(out[285]), .A(rst), .Z(N303) );
  ANDN U6864 ( .B(out[286]), .A(rst), .Z(N304) );
  ANDN U6865 ( .B(out[287]), .A(rst), .Z(N305) );
  ANDN U6866 ( .B(out[288]), .A(rst), .Z(N306) );
  ANDN U6867 ( .B(out[289]), .A(rst), .Z(N307) );
  ANDN U6868 ( .B(out[290]), .A(rst), .Z(N308) );
  ANDN U6869 ( .B(out[291]), .A(rst), .Z(N309) );
  ANDN U6870 ( .B(out[13]), .A(rst), .Z(N31) );
  ANDN U6871 ( .B(out[292]), .A(rst), .Z(N310) );
  ANDN U6872 ( .B(out[293]), .A(rst), .Z(N311) );
  ANDN U6873 ( .B(out[294]), .A(rst), .Z(N312) );
  ANDN U6874 ( .B(out[295]), .A(rst), .Z(N313) );
  ANDN U6875 ( .B(out[296]), .A(rst), .Z(N314) );
  ANDN U6876 ( .B(out[297]), .A(rst), .Z(N315) );
  ANDN U6877 ( .B(out[298]), .A(rst), .Z(N316) );
  ANDN U6878 ( .B(out[299]), .A(rst), .Z(N317) );
  ANDN U6879 ( .B(out[300]), .A(rst), .Z(N318) );
  ANDN U6880 ( .B(out[301]), .A(rst), .Z(N319) );
  ANDN U6881 ( .B(out[14]), .A(rst), .Z(N32) );
  ANDN U6882 ( .B(out[302]), .A(rst), .Z(N320) );
  ANDN U6883 ( .B(out[303]), .A(rst), .Z(N321) );
  ANDN U6884 ( .B(out[304]), .A(rst), .Z(N322) );
  ANDN U6885 ( .B(out[305]), .A(rst), .Z(N323) );
  ANDN U6886 ( .B(out[306]), .A(rst), .Z(N324) );
  ANDN U6887 ( .B(out[307]), .A(rst), .Z(N325) );
  ANDN U6888 ( .B(out[308]), .A(rst), .Z(N326) );
  ANDN U6889 ( .B(out[309]), .A(rst), .Z(N327) );
  ANDN U6890 ( .B(out[310]), .A(rst), .Z(N328) );
  ANDN U6891 ( .B(out[311]), .A(rst), .Z(N329) );
  ANDN U6892 ( .B(out[15]), .A(rst), .Z(N33) );
  ANDN U6893 ( .B(out[312]), .A(rst), .Z(N330) );
  ANDN U6894 ( .B(out[313]), .A(rst), .Z(N331) );
  ANDN U6895 ( .B(out[314]), .A(rst), .Z(N332) );
  ANDN U6896 ( .B(out[315]), .A(rst), .Z(N333) );
  ANDN U6897 ( .B(out[316]), .A(rst), .Z(N334) );
  ANDN U6898 ( .B(out[317]), .A(rst), .Z(N335) );
  ANDN U6899 ( .B(out[318]), .A(rst), .Z(N336) );
  ANDN U6900 ( .B(out[319]), .A(rst), .Z(N337) );
  ANDN U6901 ( .B(out[320]), .A(rst), .Z(N338) );
  ANDN U6902 ( .B(out[321]), .A(rst), .Z(N339) );
  ANDN U6903 ( .B(out[16]), .A(rst), .Z(N34) );
  ANDN U6904 ( .B(out[322]), .A(rst), .Z(N340) );
  ANDN U6905 ( .B(out[323]), .A(rst), .Z(N341) );
  ANDN U6906 ( .B(out[324]), .A(rst), .Z(N342) );
  ANDN U6907 ( .B(out[325]), .A(rst), .Z(N343) );
  ANDN U6908 ( .B(out[326]), .A(rst), .Z(N344) );
  ANDN U6909 ( .B(out[327]), .A(rst), .Z(N345) );
  ANDN U6910 ( .B(out[328]), .A(rst), .Z(N346) );
  ANDN U6911 ( .B(out[329]), .A(rst), .Z(N347) );
  ANDN U6912 ( .B(out[330]), .A(rst), .Z(N348) );
  ANDN U6913 ( .B(out[331]), .A(rst), .Z(N349) );
  ANDN U6914 ( .B(out[17]), .A(rst), .Z(N35) );
  ANDN U6915 ( .B(out[332]), .A(rst), .Z(N350) );
  ANDN U6916 ( .B(out[333]), .A(rst), .Z(N351) );
  ANDN U6917 ( .B(out[334]), .A(rst), .Z(N352) );
  ANDN U6918 ( .B(out[335]), .A(rst), .Z(N353) );
  ANDN U6919 ( .B(out[336]), .A(rst), .Z(N354) );
  ANDN U6920 ( .B(out[337]), .A(rst), .Z(N355) );
  ANDN U6921 ( .B(out[338]), .A(rst), .Z(N356) );
  ANDN U6922 ( .B(out[339]), .A(rst), .Z(N357) );
  ANDN U6923 ( .B(out[340]), .A(rst), .Z(N358) );
  ANDN U6924 ( .B(out[341]), .A(rst), .Z(N359) );
  ANDN U6925 ( .B(out[18]), .A(rst), .Z(N36) );
  ANDN U6926 ( .B(out[342]), .A(rst), .Z(N360) );
  ANDN U6927 ( .B(out[343]), .A(rst), .Z(N361) );
  ANDN U6928 ( .B(out[344]), .A(rst), .Z(N362) );
  ANDN U6929 ( .B(out[345]), .A(rst), .Z(N363) );
  ANDN U6930 ( .B(out[346]), .A(rst), .Z(N364) );
  ANDN U6931 ( .B(out[347]), .A(rst), .Z(N365) );
  ANDN U6932 ( .B(out[348]), .A(rst), .Z(N366) );
  ANDN U6933 ( .B(out[349]), .A(rst), .Z(N367) );
  ANDN U6934 ( .B(out[350]), .A(rst), .Z(N368) );
  ANDN U6935 ( .B(out[351]), .A(rst), .Z(N369) );
  ANDN U6936 ( .B(out[19]), .A(rst), .Z(N37) );
  ANDN U6937 ( .B(out[352]), .A(rst), .Z(N370) );
  ANDN U6938 ( .B(out[353]), .A(rst), .Z(N371) );
  ANDN U6939 ( .B(out[354]), .A(rst), .Z(N372) );
  ANDN U6940 ( .B(out[355]), .A(rst), .Z(N373) );
  ANDN U6941 ( .B(out[356]), .A(rst), .Z(N374) );
  ANDN U6942 ( .B(out[357]), .A(rst), .Z(N375) );
  ANDN U6943 ( .B(out[358]), .A(rst), .Z(N376) );
  ANDN U6944 ( .B(out[359]), .A(rst), .Z(N377) );
  ANDN U6945 ( .B(out[360]), .A(rst), .Z(N378) );
  ANDN U6946 ( .B(out[361]), .A(rst), .Z(N379) );
  ANDN U6947 ( .B(out[20]), .A(rst), .Z(N38) );
  ANDN U6948 ( .B(out[362]), .A(rst), .Z(N380) );
  ANDN U6949 ( .B(out[363]), .A(rst), .Z(N381) );
  ANDN U6950 ( .B(out[364]), .A(rst), .Z(N382) );
  ANDN U6951 ( .B(out[365]), .A(rst), .Z(N383) );
  ANDN U6952 ( .B(out[366]), .A(rst), .Z(N384) );
  ANDN U6953 ( .B(out[367]), .A(rst), .Z(N385) );
  ANDN U6954 ( .B(out[368]), .A(rst), .Z(N386) );
  ANDN U6955 ( .B(out[369]), .A(rst), .Z(N387) );
  ANDN U6956 ( .B(out[370]), .A(rst), .Z(N388) );
  ANDN U6957 ( .B(out[371]), .A(rst), .Z(N389) );
  ANDN U6958 ( .B(out[21]), .A(rst), .Z(N39) );
  ANDN U6959 ( .B(out[372]), .A(rst), .Z(N390) );
  ANDN U6960 ( .B(out[373]), .A(rst), .Z(N391) );
  ANDN U6961 ( .B(out[374]), .A(rst), .Z(N392) );
  ANDN U6962 ( .B(out[375]), .A(rst), .Z(N393) );
  ANDN U6963 ( .B(out[376]), .A(rst), .Z(N394) );
  ANDN U6964 ( .B(out[377]), .A(rst), .Z(N395) );
  ANDN U6965 ( .B(out[378]), .A(rst), .Z(N396) );
  ANDN U6966 ( .B(out[379]), .A(rst), .Z(N397) );
  ANDN U6967 ( .B(out[380]), .A(rst), .Z(N398) );
  ANDN U6968 ( .B(out[381]), .A(rst), .Z(N399) );
  ANDN U6969 ( .B(out[22]), .A(rst), .Z(N40) );
  ANDN U6970 ( .B(out[382]), .A(rst), .Z(N400) );
  ANDN U6971 ( .B(out[383]), .A(rst), .Z(N401) );
  ANDN U6972 ( .B(out[384]), .A(rst), .Z(N402) );
  ANDN U6973 ( .B(out[385]), .A(rst), .Z(N403) );
  ANDN U6974 ( .B(out[386]), .A(rst), .Z(N404) );
  ANDN U6975 ( .B(out[387]), .A(rst), .Z(N405) );
  ANDN U6976 ( .B(out[388]), .A(rst), .Z(N406) );
  ANDN U6977 ( .B(out[389]), .A(rst), .Z(N407) );
  ANDN U6978 ( .B(out[390]), .A(rst), .Z(N408) );
  ANDN U6979 ( .B(out[391]), .A(rst), .Z(N409) );
  ANDN U6980 ( .B(out[23]), .A(rst), .Z(N41) );
  ANDN U6981 ( .B(out[392]), .A(rst), .Z(N410) );
  ANDN U6982 ( .B(out[393]), .A(rst), .Z(N411) );
  ANDN U6983 ( .B(out[394]), .A(rst), .Z(N412) );
  ANDN U6984 ( .B(out[395]), .A(rst), .Z(N413) );
  ANDN U6985 ( .B(out[396]), .A(rst), .Z(N414) );
  ANDN U6986 ( .B(out[397]), .A(rst), .Z(N415) );
  ANDN U6987 ( .B(out[398]), .A(rst), .Z(N416) );
  ANDN U6988 ( .B(out[399]), .A(rst), .Z(N417) );
  ANDN U6989 ( .B(out[400]), .A(rst), .Z(N418) );
  ANDN U6990 ( .B(out[401]), .A(rst), .Z(N419) );
  ANDN U6991 ( .B(out[24]), .A(rst), .Z(N42) );
  ANDN U6992 ( .B(out[402]), .A(rst), .Z(N420) );
  ANDN U6993 ( .B(out[403]), .A(rst), .Z(N421) );
  ANDN U6994 ( .B(out[404]), .A(rst), .Z(N422) );
  ANDN U6995 ( .B(out[405]), .A(rst), .Z(N423) );
  ANDN U6996 ( .B(out[406]), .A(rst), .Z(N424) );
  ANDN U6997 ( .B(out[407]), .A(rst), .Z(N425) );
  ANDN U6998 ( .B(out[408]), .A(rst), .Z(N426) );
  ANDN U6999 ( .B(out[409]), .A(rst), .Z(N427) );
  ANDN U7000 ( .B(out[410]), .A(rst), .Z(N428) );
  ANDN U7001 ( .B(out[411]), .A(rst), .Z(N429) );
  ANDN U7002 ( .B(out[25]), .A(rst), .Z(N43) );
  ANDN U7003 ( .B(out[412]), .A(rst), .Z(N430) );
  ANDN U7004 ( .B(out[413]), .A(rst), .Z(N431) );
  ANDN U7005 ( .B(out[414]), .A(rst), .Z(N432) );
  ANDN U7006 ( .B(out[415]), .A(rst), .Z(N433) );
  ANDN U7007 ( .B(out[416]), .A(rst), .Z(N434) );
  ANDN U7008 ( .B(out[417]), .A(rst), .Z(N435) );
  ANDN U7009 ( .B(out[418]), .A(rst), .Z(N436) );
  ANDN U7010 ( .B(out[419]), .A(rst), .Z(N437) );
  ANDN U7011 ( .B(out[420]), .A(rst), .Z(N438) );
  ANDN U7012 ( .B(out[421]), .A(rst), .Z(N439) );
  ANDN U7013 ( .B(out[26]), .A(rst), .Z(N44) );
  ANDN U7014 ( .B(out[422]), .A(rst), .Z(N440) );
  ANDN U7015 ( .B(out[423]), .A(rst), .Z(N441) );
  ANDN U7016 ( .B(out[424]), .A(rst), .Z(N442) );
  ANDN U7017 ( .B(out[425]), .A(rst), .Z(N443) );
  ANDN U7018 ( .B(out[426]), .A(rst), .Z(N444) );
  ANDN U7019 ( .B(out[427]), .A(rst), .Z(N445) );
  ANDN U7020 ( .B(out[428]), .A(rst), .Z(N446) );
  ANDN U7021 ( .B(out[429]), .A(rst), .Z(N447) );
  ANDN U7022 ( .B(out[430]), .A(rst), .Z(N448) );
  ANDN U7023 ( .B(out[431]), .A(rst), .Z(N449) );
  ANDN U7024 ( .B(out[27]), .A(rst), .Z(N45) );
  ANDN U7025 ( .B(out[432]), .A(rst), .Z(N450) );
  ANDN U7026 ( .B(out[433]), .A(rst), .Z(N451) );
  ANDN U7027 ( .B(out[434]), .A(rst), .Z(N452) );
  ANDN U7028 ( .B(out[435]), .A(rst), .Z(N453) );
  ANDN U7029 ( .B(out[436]), .A(rst), .Z(N454) );
  ANDN U7030 ( .B(out[437]), .A(rst), .Z(N455) );
  ANDN U7031 ( .B(out[438]), .A(rst), .Z(N456) );
  ANDN U7032 ( .B(out[439]), .A(rst), .Z(N457) );
  ANDN U7033 ( .B(out[440]), .A(rst), .Z(N458) );
  ANDN U7034 ( .B(out[441]), .A(rst), .Z(N459) );
  ANDN U7035 ( .B(out[28]), .A(rst), .Z(N46) );
  ANDN U7036 ( .B(out[442]), .A(rst), .Z(N460) );
  ANDN U7037 ( .B(out[443]), .A(rst), .Z(N461) );
  ANDN U7038 ( .B(out[444]), .A(rst), .Z(N462) );
  ANDN U7039 ( .B(out[445]), .A(rst), .Z(N463) );
  ANDN U7040 ( .B(out[446]), .A(rst), .Z(N464) );
  ANDN U7041 ( .B(out[447]), .A(rst), .Z(N465) );
  ANDN U7042 ( .B(out[448]), .A(rst), .Z(N466) );
  ANDN U7043 ( .B(out[449]), .A(rst), .Z(N467) );
  ANDN U7044 ( .B(out[450]), .A(rst), .Z(N468) );
  ANDN U7045 ( .B(out[451]), .A(rst), .Z(N469) );
  ANDN U7046 ( .B(out[29]), .A(rst), .Z(N47) );
  ANDN U7047 ( .B(out[452]), .A(rst), .Z(N470) );
  ANDN U7048 ( .B(out[453]), .A(rst), .Z(N471) );
  ANDN U7049 ( .B(out[454]), .A(rst), .Z(N472) );
  ANDN U7050 ( .B(out[455]), .A(rst), .Z(N473) );
  ANDN U7051 ( .B(out[456]), .A(rst), .Z(N474) );
  ANDN U7052 ( .B(out[457]), .A(rst), .Z(N475) );
  ANDN U7053 ( .B(out[458]), .A(rst), .Z(N476) );
  ANDN U7054 ( .B(out[459]), .A(rst), .Z(N477) );
  ANDN U7055 ( .B(out[460]), .A(rst), .Z(N478) );
  ANDN U7056 ( .B(out[461]), .A(rst), .Z(N479) );
  ANDN U7057 ( .B(out[30]), .A(rst), .Z(N48) );
  ANDN U7058 ( .B(out[462]), .A(rst), .Z(N480) );
  ANDN U7059 ( .B(out[463]), .A(rst), .Z(N481) );
  ANDN U7060 ( .B(out[464]), .A(rst), .Z(N482) );
  ANDN U7061 ( .B(out[465]), .A(rst), .Z(N483) );
  ANDN U7062 ( .B(out[466]), .A(rst), .Z(N484) );
  ANDN U7063 ( .B(out[467]), .A(rst), .Z(N485) );
  ANDN U7064 ( .B(out[468]), .A(rst), .Z(N486) );
  ANDN U7065 ( .B(out[469]), .A(rst), .Z(N487) );
  ANDN U7066 ( .B(out[470]), .A(rst), .Z(N488) );
  ANDN U7067 ( .B(out[471]), .A(rst), .Z(N489) );
  ANDN U7068 ( .B(out[31]), .A(rst), .Z(N49) );
  ANDN U7069 ( .B(out[472]), .A(rst), .Z(N490) );
  ANDN U7070 ( .B(out[473]), .A(rst), .Z(N491) );
  ANDN U7071 ( .B(out[474]), .A(rst), .Z(N492) );
  ANDN U7072 ( .B(out[475]), .A(rst), .Z(N493) );
  ANDN U7073 ( .B(out[476]), .A(rst), .Z(N494) );
  ANDN U7074 ( .B(out[477]), .A(rst), .Z(N495) );
  ANDN U7075 ( .B(out[478]), .A(rst), .Z(N496) );
  ANDN U7076 ( .B(out[479]), .A(rst), .Z(N497) );
  ANDN U7077 ( .B(out[480]), .A(rst), .Z(N498) );
  ANDN U7078 ( .B(out[481]), .A(rst), .Z(N499) );
  ANDN U7079 ( .B(out[32]), .A(rst), .Z(N50) );
  ANDN U7080 ( .B(out[482]), .A(rst), .Z(N500) );
  ANDN U7081 ( .B(out[483]), .A(rst), .Z(N501) );
  ANDN U7082 ( .B(out[484]), .A(rst), .Z(N502) );
  ANDN U7083 ( .B(out[485]), .A(rst), .Z(N503) );
  ANDN U7084 ( .B(out[486]), .A(rst), .Z(N504) );
  ANDN U7085 ( .B(out[487]), .A(rst), .Z(N505) );
  ANDN U7086 ( .B(out[488]), .A(rst), .Z(N506) );
  ANDN U7087 ( .B(out[489]), .A(rst), .Z(N507) );
  ANDN U7088 ( .B(out[490]), .A(rst), .Z(N508) );
  ANDN U7089 ( .B(out[491]), .A(rst), .Z(N509) );
  ANDN U7090 ( .B(out[33]), .A(rst), .Z(N51) );
  ANDN U7091 ( .B(out[492]), .A(rst), .Z(N510) );
  ANDN U7092 ( .B(out[493]), .A(rst), .Z(N511) );
  ANDN U7093 ( .B(out[494]), .A(rst), .Z(N512) );
  ANDN U7094 ( .B(out[495]), .A(rst), .Z(N513) );
  ANDN U7095 ( .B(out[496]), .A(rst), .Z(N514) );
  ANDN U7096 ( .B(out[497]), .A(rst), .Z(N515) );
  ANDN U7097 ( .B(out[498]), .A(rst), .Z(N516) );
  ANDN U7098 ( .B(out[499]), .A(rst), .Z(N517) );
  ANDN U7099 ( .B(out[500]), .A(rst), .Z(N518) );
  ANDN U7100 ( .B(out[501]), .A(rst), .Z(N519) );
  ANDN U7101 ( .B(out[34]), .A(rst), .Z(N52) );
  ANDN U7102 ( .B(out[502]), .A(rst), .Z(N520) );
  ANDN U7103 ( .B(out[503]), .A(rst), .Z(N521) );
  ANDN U7104 ( .B(out[504]), .A(rst), .Z(N522) );
  ANDN U7105 ( .B(out[505]), .A(rst), .Z(N523) );
  ANDN U7106 ( .B(out[506]), .A(rst), .Z(N524) );
  ANDN U7107 ( .B(out[507]), .A(rst), .Z(N525) );
  ANDN U7108 ( .B(out[508]), .A(rst), .Z(N526) );
  ANDN U7109 ( .B(out[509]), .A(rst), .Z(N527) );
  ANDN U7110 ( .B(out[510]), .A(rst), .Z(N528) );
  ANDN U7111 ( .B(out[511]), .A(rst), .Z(N529) );
  ANDN U7112 ( .B(out[35]), .A(rst), .Z(N53) );
  ANDN U7113 ( .B(out[512]), .A(rst), .Z(N530) );
  ANDN U7114 ( .B(out[513]), .A(rst), .Z(N531) );
  ANDN U7115 ( .B(out[514]), .A(rst), .Z(N532) );
  ANDN U7116 ( .B(out[515]), .A(rst), .Z(N533) );
  ANDN U7117 ( .B(out[516]), .A(rst), .Z(N534) );
  ANDN U7118 ( .B(out[517]), .A(rst), .Z(N535) );
  ANDN U7119 ( .B(out[518]), .A(rst), .Z(N536) );
  ANDN U7120 ( .B(out[519]), .A(rst), .Z(N537) );
  ANDN U7121 ( .B(out[520]), .A(rst), .Z(N538) );
  ANDN U7122 ( .B(out[521]), .A(rst), .Z(N539) );
  ANDN U7123 ( .B(out[36]), .A(rst), .Z(N54) );
  ANDN U7124 ( .B(out[522]), .A(rst), .Z(N540) );
  ANDN U7125 ( .B(out[523]), .A(rst), .Z(N541) );
  ANDN U7126 ( .B(out[524]), .A(rst), .Z(N542) );
  ANDN U7127 ( .B(out[525]), .A(rst), .Z(N543) );
  ANDN U7128 ( .B(out[526]), .A(rst), .Z(N544) );
  ANDN U7129 ( .B(out[527]), .A(rst), .Z(N545) );
  ANDN U7130 ( .B(out[528]), .A(rst), .Z(N546) );
  ANDN U7131 ( .B(out[529]), .A(rst), .Z(N547) );
  ANDN U7132 ( .B(out[530]), .A(rst), .Z(N548) );
  ANDN U7133 ( .B(out[531]), .A(rst), .Z(N549) );
  ANDN U7134 ( .B(out[37]), .A(rst), .Z(N55) );
  ANDN U7135 ( .B(out[532]), .A(rst), .Z(N550) );
  ANDN U7136 ( .B(out[533]), .A(rst), .Z(N551) );
  ANDN U7137 ( .B(out[534]), .A(rst), .Z(N552) );
  ANDN U7138 ( .B(out[535]), .A(rst), .Z(N553) );
  ANDN U7139 ( .B(out[536]), .A(rst), .Z(N554) );
  ANDN U7140 ( .B(out[537]), .A(rst), .Z(N555) );
  ANDN U7141 ( .B(out[538]), .A(rst), .Z(N556) );
  ANDN U7142 ( .B(out[539]), .A(rst), .Z(N557) );
  ANDN U7143 ( .B(out[540]), .A(rst), .Z(N558) );
  ANDN U7144 ( .B(out[541]), .A(rst), .Z(N559) );
  ANDN U7145 ( .B(out[38]), .A(rst), .Z(N56) );
  ANDN U7146 ( .B(out[542]), .A(rst), .Z(N560) );
  ANDN U7147 ( .B(out[543]), .A(rst), .Z(N561) );
  ANDN U7148 ( .B(out[544]), .A(rst), .Z(N562) );
  ANDN U7149 ( .B(out[545]), .A(rst), .Z(N563) );
  ANDN U7150 ( .B(out[546]), .A(rst), .Z(N564) );
  ANDN U7151 ( .B(out[547]), .A(rst), .Z(N565) );
  ANDN U7152 ( .B(out[548]), .A(rst), .Z(N566) );
  ANDN U7153 ( .B(out[549]), .A(rst), .Z(N567) );
  ANDN U7154 ( .B(out[550]), .A(rst), .Z(N568) );
  ANDN U7155 ( .B(out[551]), .A(rst), .Z(N569) );
  ANDN U7156 ( .B(out[39]), .A(rst), .Z(N57) );
  ANDN U7157 ( .B(out[552]), .A(rst), .Z(N570) );
  ANDN U7158 ( .B(out[553]), .A(rst), .Z(N571) );
  ANDN U7159 ( .B(out[554]), .A(rst), .Z(N572) );
  ANDN U7160 ( .B(out[555]), .A(rst), .Z(N573) );
  ANDN U7161 ( .B(out[556]), .A(rst), .Z(N574) );
  ANDN U7162 ( .B(out[557]), .A(rst), .Z(N575) );
  ANDN U7163 ( .B(out[558]), .A(rst), .Z(N576) );
  ANDN U7164 ( .B(out[559]), .A(rst), .Z(N577) );
  ANDN U7165 ( .B(out[560]), .A(rst), .Z(N578) );
  ANDN U7166 ( .B(out[561]), .A(rst), .Z(N579) );
  ANDN U7167 ( .B(out[40]), .A(rst), .Z(N58) );
  ANDN U7168 ( .B(out[562]), .A(rst), .Z(N580) );
  ANDN U7169 ( .B(out[563]), .A(rst), .Z(N581) );
  ANDN U7170 ( .B(out[564]), .A(rst), .Z(N582) );
  ANDN U7171 ( .B(out[565]), .A(rst), .Z(N583) );
  ANDN U7172 ( .B(out[566]), .A(rst), .Z(N584) );
  ANDN U7173 ( .B(out[567]), .A(rst), .Z(N585) );
  ANDN U7174 ( .B(out[568]), .A(rst), .Z(N586) );
  ANDN U7175 ( .B(out[569]), .A(rst), .Z(N587) );
  ANDN U7176 ( .B(out[570]), .A(rst), .Z(N588) );
  ANDN U7177 ( .B(out[571]), .A(rst), .Z(N589) );
  ANDN U7178 ( .B(out[41]), .A(rst), .Z(N59) );
  ANDN U7179 ( .B(out[572]), .A(rst), .Z(N590) );
  ANDN U7180 ( .B(out[573]), .A(rst), .Z(N591) );
  ANDN U7181 ( .B(out[574]), .A(rst), .Z(N592) );
  ANDN U7182 ( .B(out[575]), .A(rst), .Z(N593) );
  ANDN U7183 ( .B(out[576]), .A(rst), .Z(N594) );
  ANDN U7184 ( .B(out[577]), .A(rst), .Z(N595) );
  ANDN U7185 ( .B(out[578]), .A(rst), .Z(N596) );
  ANDN U7186 ( .B(out[579]), .A(rst), .Z(N597) );
  ANDN U7187 ( .B(out[580]), .A(rst), .Z(N598) );
  ANDN U7188 ( .B(out[581]), .A(rst), .Z(N599) );
  NOR U7189 ( .A(rst), .B(init), .Z(N6) );
  ANDN U7190 ( .B(out[42]), .A(rst), .Z(N60) );
  ANDN U7191 ( .B(out[582]), .A(rst), .Z(N600) );
  ANDN U7192 ( .B(out[583]), .A(rst), .Z(N601) );
  ANDN U7193 ( .B(out[584]), .A(rst), .Z(N602) );
  ANDN U7194 ( .B(out[585]), .A(rst), .Z(N603) );
  ANDN U7195 ( .B(out[586]), .A(rst), .Z(N604) );
  ANDN U7196 ( .B(out[587]), .A(rst), .Z(N605) );
  ANDN U7197 ( .B(out[588]), .A(rst), .Z(N606) );
  ANDN U7198 ( .B(out[589]), .A(rst), .Z(N607) );
  ANDN U7199 ( .B(out[590]), .A(rst), .Z(N608) );
  ANDN U7200 ( .B(out[591]), .A(rst), .Z(N609) );
  ANDN U7201 ( .B(out[43]), .A(rst), .Z(N61) );
  ANDN U7202 ( .B(out[592]), .A(rst), .Z(N610) );
  ANDN U7203 ( .B(out[593]), .A(rst), .Z(N611) );
  ANDN U7204 ( .B(out[594]), .A(rst), .Z(N612) );
  ANDN U7205 ( .B(out[595]), .A(rst), .Z(N613) );
  ANDN U7206 ( .B(out[596]), .A(rst), .Z(N614) );
  ANDN U7207 ( .B(out[597]), .A(rst), .Z(N615) );
  ANDN U7208 ( .B(out[598]), .A(rst), .Z(N616) );
  ANDN U7209 ( .B(out[599]), .A(rst), .Z(N617) );
  ANDN U7210 ( .B(out[600]), .A(rst), .Z(N618) );
  ANDN U7211 ( .B(out[601]), .A(rst), .Z(N619) );
  ANDN U7212 ( .B(out[44]), .A(rst), .Z(N62) );
  ANDN U7213 ( .B(out[602]), .A(rst), .Z(N620) );
  ANDN U7214 ( .B(out[603]), .A(rst), .Z(N621) );
  ANDN U7215 ( .B(out[604]), .A(rst), .Z(N622) );
  ANDN U7216 ( .B(out[605]), .A(rst), .Z(N623) );
  ANDN U7217 ( .B(out[606]), .A(rst), .Z(N624) );
  ANDN U7218 ( .B(out[607]), .A(rst), .Z(N625) );
  ANDN U7219 ( .B(out[608]), .A(rst), .Z(N626) );
  ANDN U7220 ( .B(out[609]), .A(rst), .Z(N627) );
  ANDN U7221 ( .B(out[610]), .A(rst), .Z(N628) );
  ANDN U7222 ( .B(out[611]), .A(rst), .Z(N629) );
  ANDN U7223 ( .B(out[45]), .A(rst), .Z(N63) );
  ANDN U7224 ( .B(out[612]), .A(rst), .Z(N630) );
  ANDN U7225 ( .B(out[613]), .A(rst), .Z(N631) );
  ANDN U7226 ( .B(out[614]), .A(rst), .Z(N632) );
  ANDN U7227 ( .B(out[615]), .A(rst), .Z(N633) );
  ANDN U7228 ( .B(out[616]), .A(rst), .Z(N634) );
  ANDN U7229 ( .B(out[617]), .A(rst), .Z(N635) );
  ANDN U7230 ( .B(out[618]), .A(rst), .Z(N636) );
  ANDN U7231 ( .B(out[619]), .A(rst), .Z(N637) );
  ANDN U7232 ( .B(out[620]), .A(rst), .Z(N638) );
  ANDN U7233 ( .B(out[621]), .A(rst), .Z(N639) );
  ANDN U7234 ( .B(out[46]), .A(rst), .Z(N64) );
  ANDN U7235 ( .B(out[622]), .A(rst), .Z(N640) );
  ANDN U7236 ( .B(out[623]), .A(rst), .Z(N641) );
  ANDN U7237 ( .B(out[624]), .A(rst), .Z(N642) );
  ANDN U7238 ( .B(out[625]), .A(rst), .Z(N643) );
  ANDN U7239 ( .B(out[626]), .A(rst), .Z(N644) );
  ANDN U7240 ( .B(out[627]), .A(rst), .Z(N645) );
  ANDN U7241 ( .B(out[628]), .A(rst), .Z(N646) );
  ANDN U7242 ( .B(out[629]), .A(rst), .Z(N647) );
  ANDN U7243 ( .B(out[630]), .A(rst), .Z(N648) );
  ANDN U7244 ( .B(out[631]), .A(rst), .Z(N649) );
  ANDN U7245 ( .B(out[47]), .A(rst), .Z(N65) );
  ANDN U7246 ( .B(out[632]), .A(rst), .Z(N650) );
  ANDN U7247 ( .B(out[633]), .A(rst), .Z(N651) );
  ANDN U7248 ( .B(out[634]), .A(rst), .Z(N652) );
  ANDN U7249 ( .B(out[635]), .A(rst), .Z(N653) );
  ANDN U7250 ( .B(out[636]), .A(rst), .Z(N654) );
  ANDN U7251 ( .B(out[637]), .A(rst), .Z(N655) );
  ANDN U7252 ( .B(out[638]), .A(rst), .Z(N656) );
  ANDN U7253 ( .B(out[639]), .A(rst), .Z(N657) );
  ANDN U7254 ( .B(out[640]), .A(rst), .Z(N658) );
  ANDN U7255 ( .B(out[641]), .A(rst), .Z(N659) );
  ANDN U7256 ( .B(out[48]), .A(rst), .Z(N66) );
  ANDN U7257 ( .B(out[642]), .A(rst), .Z(N660) );
  ANDN U7258 ( .B(out[643]), .A(rst), .Z(N661) );
  ANDN U7259 ( .B(out[644]), .A(rst), .Z(N662) );
  ANDN U7260 ( .B(out[645]), .A(rst), .Z(N663) );
  ANDN U7261 ( .B(out[646]), .A(rst), .Z(N664) );
  ANDN U7262 ( .B(out[647]), .A(rst), .Z(N665) );
  ANDN U7263 ( .B(out[648]), .A(rst), .Z(N666) );
  ANDN U7264 ( .B(out[649]), .A(rst), .Z(N667) );
  ANDN U7265 ( .B(out[650]), .A(rst), .Z(N668) );
  ANDN U7266 ( .B(out[651]), .A(rst), .Z(N669) );
  ANDN U7267 ( .B(out[49]), .A(rst), .Z(N67) );
  ANDN U7268 ( .B(out[652]), .A(rst), .Z(N670) );
  ANDN U7269 ( .B(out[653]), .A(rst), .Z(N671) );
  ANDN U7270 ( .B(out[654]), .A(rst), .Z(N672) );
  ANDN U7271 ( .B(out[655]), .A(rst), .Z(N673) );
  ANDN U7272 ( .B(out[656]), .A(rst), .Z(N674) );
  ANDN U7273 ( .B(out[657]), .A(rst), .Z(N675) );
  ANDN U7274 ( .B(out[658]), .A(rst), .Z(N676) );
  ANDN U7275 ( .B(out[659]), .A(rst), .Z(N677) );
  ANDN U7276 ( .B(out[660]), .A(rst), .Z(N678) );
  ANDN U7277 ( .B(out[661]), .A(rst), .Z(N679) );
  ANDN U7278 ( .B(out[50]), .A(rst), .Z(N68) );
  ANDN U7279 ( .B(out[662]), .A(rst), .Z(N680) );
  ANDN U7280 ( .B(out[663]), .A(rst), .Z(N681) );
  ANDN U7281 ( .B(out[664]), .A(rst), .Z(N682) );
  ANDN U7282 ( .B(out[665]), .A(rst), .Z(N683) );
  ANDN U7283 ( .B(out[666]), .A(rst), .Z(N684) );
  ANDN U7284 ( .B(out[667]), .A(rst), .Z(N685) );
  ANDN U7285 ( .B(out[668]), .A(rst), .Z(N686) );
  ANDN U7286 ( .B(out[669]), .A(rst), .Z(N687) );
  ANDN U7287 ( .B(out[670]), .A(rst), .Z(N688) );
  ANDN U7288 ( .B(out[671]), .A(rst), .Z(N689) );
  ANDN U7289 ( .B(out[51]), .A(rst), .Z(N69) );
  ANDN U7290 ( .B(out[672]), .A(rst), .Z(N690) );
  ANDN U7291 ( .B(out[673]), .A(rst), .Z(N691) );
  ANDN U7292 ( .B(out[674]), .A(rst), .Z(N692) );
  ANDN U7293 ( .B(out[675]), .A(rst), .Z(N693) );
  ANDN U7294 ( .B(out[676]), .A(rst), .Z(N694) );
  ANDN U7295 ( .B(out[677]), .A(rst), .Z(N695) );
  ANDN U7296 ( .B(out[678]), .A(rst), .Z(N696) );
  ANDN U7297 ( .B(out[679]), .A(rst), .Z(N697) );
  ANDN U7298 ( .B(out[680]), .A(rst), .Z(N698) );
  ANDN U7299 ( .B(out[681]), .A(rst), .Z(N699) );
  ANDN U7300 ( .B(rc_i[0]), .A(rst), .Z(N7) );
  ANDN U7301 ( .B(out[52]), .A(rst), .Z(N70) );
  ANDN U7302 ( .B(out[682]), .A(rst), .Z(N700) );
  ANDN U7303 ( .B(out[683]), .A(rst), .Z(N701) );
  ANDN U7304 ( .B(out[684]), .A(rst), .Z(N702) );
  ANDN U7305 ( .B(out[685]), .A(rst), .Z(N703) );
  ANDN U7306 ( .B(out[686]), .A(rst), .Z(N704) );
  ANDN U7307 ( .B(out[687]), .A(rst), .Z(N705) );
  ANDN U7308 ( .B(out[688]), .A(rst), .Z(N706) );
  ANDN U7309 ( .B(out[689]), .A(rst), .Z(N707) );
  ANDN U7310 ( .B(out[690]), .A(rst), .Z(N708) );
  ANDN U7311 ( .B(out[691]), .A(rst), .Z(N709) );
  ANDN U7312 ( .B(out[53]), .A(rst), .Z(N71) );
  ANDN U7313 ( .B(out[692]), .A(rst), .Z(N710) );
  ANDN U7314 ( .B(out[693]), .A(rst), .Z(N711) );
  ANDN U7315 ( .B(out[694]), .A(rst), .Z(N712) );
  ANDN U7316 ( .B(out[695]), .A(rst), .Z(N713) );
  ANDN U7317 ( .B(out[696]), .A(rst), .Z(N714) );
  ANDN U7318 ( .B(out[697]), .A(rst), .Z(N715) );
  ANDN U7319 ( .B(out[698]), .A(rst), .Z(N716) );
  ANDN U7320 ( .B(out[699]), .A(rst), .Z(N717) );
  ANDN U7321 ( .B(out[700]), .A(rst), .Z(N718) );
  ANDN U7322 ( .B(out[701]), .A(rst), .Z(N719) );
  ANDN U7323 ( .B(out[54]), .A(rst), .Z(N72) );
  ANDN U7324 ( .B(out[702]), .A(rst), .Z(N720) );
  ANDN U7325 ( .B(out[703]), .A(rst), .Z(N721) );
  ANDN U7326 ( .B(out[704]), .A(rst), .Z(N722) );
  ANDN U7327 ( .B(out[705]), .A(rst), .Z(N723) );
  ANDN U7328 ( .B(out[706]), .A(rst), .Z(N724) );
  ANDN U7329 ( .B(out[707]), .A(rst), .Z(N725) );
  ANDN U7330 ( .B(out[708]), .A(rst), .Z(N726) );
  ANDN U7331 ( .B(out[709]), .A(rst), .Z(N727) );
  ANDN U7332 ( .B(out[710]), .A(rst), .Z(N728) );
  ANDN U7333 ( .B(out[711]), .A(rst), .Z(N729) );
  ANDN U7334 ( .B(out[55]), .A(rst), .Z(N73) );
  ANDN U7335 ( .B(out[712]), .A(rst), .Z(N730) );
  ANDN U7336 ( .B(out[713]), .A(rst), .Z(N731) );
  ANDN U7337 ( .B(out[714]), .A(rst), .Z(N732) );
  ANDN U7338 ( .B(out[715]), .A(rst), .Z(N733) );
  ANDN U7339 ( .B(out[716]), .A(rst), .Z(N734) );
  ANDN U7340 ( .B(out[717]), .A(rst), .Z(N735) );
  ANDN U7341 ( .B(out[718]), .A(rst), .Z(N736) );
  ANDN U7342 ( .B(out[719]), .A(rst), .Z(N737) );
  ANDN U7343 ( .B(out[720]), .A(rst), .Z(N738) );
  ANDN U7344 ( .B(out[721]), .A(rst), .Z(N739) );
  ANDN U7345 ( .B(out[56]), .A(rst), .Z(N74) );
  ANDN U7346 ( .B(out[722]), .A(rst), .Z(N740) );
  ANDN U7347 ( .B(out[723]), .A(rst), .Z(N741) );
  ANDN U7348 ( .B(out[724]), .A(rst), .Z(N742) );
  ANDN U7349 ( .B(out[725]), .A(rst), .Z(N743) );
  ANDN U7350 ( .B(out[726]), .A(rst), .Z(N744) );
  ANDN U7351 ( .B(out[727]), .A(rst), .Z(N745) );
  ANDN U7352 ( .B(out[728]), .A(rst), .Z(N746) );
  ANDN U7353 ( .B(out[729]), .A(rst), .Z(N747) );
  ANDN U7354 ( .B(out[730]), .A(rst), .Z(N748) );
  ANDN U7355 ( .B(out[731]), .A(rst), .Z(N749) );
  ANDN U7356 ( .B(out[57]), .A(rst), .Z(N75) );
  ANDN U7357 ( .B(out[732]), .A(rst), .Z(N750) );
  ANDN U7358 ( .B(out[733]), .A(rst), .Z(N751) );
  ANDN U7359 ( .B(out[734]), .A(rst), .Z(N752) );
  ANDN U7360 ( .B(out[735]), .A(rst), .Z(N753) );
  ANDN U7361 ( .B(out[736]), .A(rst), .Z(N754) );
  ANDN U7362 ( .B(out[737]), .A(rst), .Z(N755) );
  ANDN U7363 ( .B(out[738]), .A(rst), .Z(N756) );
  ANDN U7364 ( .B(out[739]), .A(rst), .Z(N757) );
  ANDN U7365 ( .B(out[740]), .A(rst), .Z(N758) );
  ANDN U7366 ( .B(out[741]), .A(rst), .Z(N759) );
  ANDN U7367 ( .B(out[58]), .A(rst), .Z(N76) );
  ANDN U7368 ( .B(out[742]), .A(rst), .Z(N760) );
  ANDN U7369 ( .B(out[743]), .A(rst), .Z(N761) );
  ANDN U7370 ( .B(out[744]), .A(rst), .Z(N762) );
  ANDN U7371 ( .B(out[745]), .A(rst), .Z(N763) );
  ANDN U7372 ( .B(out[746]), .A(rst), .Z(N764) );
  ANDN U7373 ( .B(out[747]), .A(rst), .Z(N765) );
  ANDN U7374 ( .B(out[748]), .A(rst), .Z(N766) );
  ANDN U7375 ( .B(out[749]), .A(rst), .Z(N767) );
  ANDN U7376 ( .B(out[750]), .A(rst), .Z(N768) );
  ANDN U7377 ( .B(out[751]), .A(rst), .Z(N769) );
  ANDN U7378 ( .B(out[59]), .A(rst), .Z(N77) );
  ANDN U7379 ( .B(out[752]), .A(rst), .Z(N770) );
  ANDN U7380 ( .B(out[753]), .A(rst), .Z(N771) );
  ANDN U7381 ( .B(out[754]), .A(rst), .Z(N772) );
  ANDN U7382 ( .B(out[755]), .A(rst), .Z(N773) );
  ANDN U7383 ( .B(out[756]), .A(rst), .Z(N774) );
  ANDN U7384 ( .B(out[757]), .A(rst), .Z(N775) );
  ANDN U7385 ( .B(out[758]), .A(rst), .Z(N776) );
  ANDN U7386 ( .B(out[759]), .A(rst), .Z(N777) );
  ANDN U7387 ( .B(out[760]), .A(rst), .Z(N778) );
  ANDN U7388 ( .B(out[761]), .A(rst), .Z(N779) );
  ANDN U7389 ( .B(out[60]), .A(rst), .Z(N78) );
  ANDN U7390 ( .B(out[762]), .A(rst), .Z(N780) );
  ANDN U7391 ( .B(out[763]), .A(rst), .Z(N781) );
  ANDN U7392 ( .B(out[764]), .A(rst), .Z(N782) );
  ANDN U7393 ( .B(out[765]), .A(rst), .Z(N783) );
  ANDN U7394 ( .B(out[766]), .A(rst), .Z(N784) );
  ANDN U7395 ( .B(out[767]), .A(rst), .Z(N785) );
  ANDN U7396 ( .B(out[768]), .A(rst), .Z(N786) );
  ANDN U7397 ( .B(out[769]), .A(rst), .Z(N787) );
  ANDN U7398 ( .B(out[770]), .A(rst), .Z(N788) );
  ANDN U7399 ( .B(out[771]), .A(rst), .Z(N789) );
  ANDN U7400 ( .B(out[61]), .A(rst), .Z(N79) );
  ANDN U7401 ( .B(out[772]), .A(rst), .Z(N790) );
  ANDN U7402 ( .B(out[773]), .A(rst), .Z(N791) );
  ANDN U7403 ( .B(out[774]), .A(rst), .Z(N792) );
  ANDN U7404 ( .B(out[775]), .A(rst), .Z(N793) );
  ANDN U7405 ( .B(out[776]), .A(rst), .Z(N794) );
  ANDN U7406 ( .B(out[777]), .A(rst), .Z(N795) );
  ANDN U7407 ( .B(out[778]), .A(rst), .Z(N796) );
  ANDN U7408 ( .B(out[779]), .A(rst), .Z(N797) );
  ANDN U7409 ( .B(out[780]), .A(rst), .Z(N798) );
  ANDN U7410 ( .B(out[781]), .A(rst), .Z(N799) );
  ANDN U7411 ( .B(rc_i[1]), .A(rst), .Z(N8) );
  ANDN U7412 ( .B(out[62]), .A(rst), .Z(N80) );
  ANDN U7413 ( .B(out[782]), .A(rst), .Z(N800) );
  ANDN U7414 ( .B(out[783]), .A(rst), .Z(N801) );
  ANDN U7415 ( .B(out[784]), .A(rst), .Z(N802) );
  ANDN U7416 ( .B(out[785]), .A(rst), .Z(N803) );
  ANDN U7417 ( .B(out[786]), .A(rst), .Z(N804) );
  ANDN U7418 ( .B(out[787]), .A(rst), .Z(N805) );
  ANDN U7419 ( .B(out[788]), .A(rst), .Z(N806) );
  ANDN U7420 ( .B(out[789]), .A(rst), .Z(N807) );
  ANDN U7421 ( .B(out[790]), .A(rst), .Z(N808) );
  ANDN U7422 ( .B(out[791]), .A(rst), .Z(N809) );
  ANDN U7423 ( .B(out[63]), .A(rst), .Z(N81) );
  ANDN U7424 ( .B(out[792]), .A(rst), .Z(N810) );
  ANDN U7425 ( .B(out[793]), .A(rst), .Z(N811) );
  ANDN U7426 ( .B(out[794]), .A(rst), .Z(N812) );
  ANDN U7427 ( .B(out[795]), .A(rst), .Z(N813) );
  ANDN U7428 ( .B(out[796]), .A(rst), .Z(N814) );
  ANDN U7429 ( .B(out[797]), .A(rst), .Z(N815) );
  ANDN U7430 ( .B(out[798]), .A(rst), .Z(N816) );
  ANDN U7431 ( .B(out[799]), .A(rst), .Z(N817) );
  ANDN U7432 ( .B(out[800]), .A(rst), .Z(N818) );
  ANDN U7433 ( .B(out[801]), .A(rst), .Z(N819) );
  ANDN U7434 ( .B(out[64]), .A(rst), .Z(N82) );
  ANDN U7435 ( .B(out[802]), .A(rst), .Z(N820) );
  ANDN U7436 ( .B(out[803]), .A(rst), .Z(N821) );
  ANDN U7437 ( .B(out[804]), .A(rst), .Z(N822) );
  ANDN U7438 ( .B(out[805]), .A(rst), .Z(N823) );
  ANDN U7439 ( .B(out[806]), .A(rst), .Z(N824) );
  ANDN U7440 ( .B(out[807]), .A(rst), .Z(N825) );
  ANDN U7441 ( .B(out[808]), .A(rst), .Z(N826) );
  ANDN U7442 ( .B(out[809]), .A(rst), .Z(N827) );
  ANDN U7443 ( .B(out[810]), .A(rst), .Z(N828) );
  ANDN U7444 ( .B(out[811]), .A(rst), .Z(N829) );
  ANDN U7445 ( .B(out[65]), .A(rst), .Z(N83) );
  ANDN U7446 ( .B(out[812]), .A(rst), .Z(N830) );
  ANDN U7447 ( .B(out[813]), .A(rst), .Z(N831) );
  ANDN U7448 ( .B(out[814]), .A(rst), .Z(N832) );
  ANDN U7449 ( .B(out[815]), .A(rst), .Z(N833) );
  ANDN U7450 ( .B(out[816]), .A(rst), .Z(N834) );
  ANDN U7451 ( .B(out[817]), .A(rst), .Z(N835) );
  ANDN U7452 ( .B(out[818]), .A(rst), .Z(N836) );
  ANDN U7453 ( .B(out[819]), .A(rst), .Z(N837) );
  ANDN U7454 ( .B(out[820]), .A(rst), .Z(N838) );
  ANDN U7455 ( .B(out[821]), .A(rst), .Z(N839) );
  ANDN U7456 ( .B(out[66]), .A(rst), .Z(N84) );
  ANDN U7457 ( .B(out[822]), .A(rst), .Z(N840) );
  ANDN U7458 ( .B(out[823]), .A(rst), .Z(N841) );
  ANDN U7459 ( .B(out[824]), .A(rst), .Z(N842) );
  ANDN U7460 ( .B(out[825]), .A(rst), .Z(N843) );
  ANDN U7461 ( .B(out[826]), .A(rst), .Z(N844) );
  ANDN U7462 ( .B(out[827]), .A(rst), .Z(N845) );
  ANDN U7463 ( .B(out[828]), .A(rst), .Z(N846) );
  ANDN U7464 ( .B(out[829]), .A(rst), .Z(N847) );
  ANDN U7465 ( .B(out[830]), .A(rst), .Z(N848) );
  ANDN U7466 ( .B(out[831]), .A(rst), .Z(N849) );
  ANDN U7467 ( .B(out[67]), .A(rst), .Z(N85) );
  ANDN U7468 ( .B(out[832]), .A(rst), .Z(N850) );
  ANDN U7469 ( .B(out[833]), .A(rst), .Z(N851) );
  ANDN U7470 ( .B(out[834]), .A(rst), .Z(N852) );
  ANDN U7471 ( .B(out[835]), .A(rst), .Z(N853) );
  ANDN U7472 ( .B(out[836]), .A(rst), .Z(N854) );
  ANDN U7473 ( .B(out[837]), .A(rst), .Z(N855) );
  ANDN U7474 ( .B(out[838]), .A(rst), .Z(N856) );
  ANDN U7475 ( .B(out[839]), .A(rst), .Z(N857) );
  ANDN U7476 ( .B(out[840]), .A(rst), .Z(N858) );
  ANDN U7477 ( .B(out[841]), .A(rst), .Z(N859) );
  ANDN U7478 ( .B(out[68]), .A(rst), .Z(N86) );
  ANDN U7479 ( .B(out[842]), .A(rst), .Z(N860) );
  ANDN U7480 ( .B(out[843]), .A(rst), .Z(N861) );
  ANDN U7481 ( .B(out[844]), .A(rst), .Z(N862) );
  ANDN U7482 ( .B(out[845]), .A(rst), .Z(N863) );
  ANDN U7483 ( .B(out[846]), .A(rst), .Z(N864) );
  ANDN U7484 ( .B(out[847]), .A(rst), .Z(N865) );
  ANDN U7485 ( .B(out[848]), .A(rst), .Z(N866) );
  ANDN U7486 ( .B(out[849]), .A(rst), .Z(N867) );
  ANDN U7487 ( .B(out[850]), .A(rst), .Z(N868) );
  ANDN U7488 ( .B(out[851]), .A(rst), .Z(N869) );
  ANDN U7489 ( .B(out[69]), .A(rst), .Z(N87) );
  ANDN U7490 ( .B(out[852]), .A(rst), .Z(N870) );
  ANDN U7491 ( .B(out[853]), .A(rst), .Z(N871) );
  ANDN U7492 ( .B(out[854]), .A(rst), .Z(N872) );
  ANDN U7493 ( .B(out[855]), .A(rst), .Z(N873) );
  ANDN U7494 ( .B(out[856]), .A(rst), .Z(N874) );
  ANDN U7495 ( .B(out[857]), .A(rst), .Z(N875) );
  ANDN U7496 ( .B(out[858]), .A(rst), .Z(N876) );
  ANDN U7497 ( .B(out[859]), .A(rst), .Z(N877) );
  ANDN U7498 ( .B(out[860]), .A(rst), .Z(N878) );
  ANDN U7499 ( .B(out[861]), .A(rst), .Z(N879) );
  ANDN U7500 ( .B(out[70]), .A(rst), .Z(N88) );
  ANDN U7501 ( .B(out[862]), .A(rst), .Z(N880) );
  ANDN U7502 ( .B(out[863]), .A(rst), .Z(N881) );
  ANDN U7503 ( .B(out[864]), .A(rst), .Z(N882) );
  ANDN U7504 ( .B(out[865]), .A(rst), .Z(N883) );
  ANDN U7505 ( .B(out[866]), .A(rst), .Z(N884) );
  ANDN U7506 ( .B(out[867]), .A(rst), .Z(N885) );
  ANDN U7507 ( .B(out[868]), .A(rst), .Z(N886) );
  ANDN U7508 ( .B(out[869]), .A(rst), .Z(N887) );
  ANDN U7509 ( .B(out[870]), .A(rst), .Z(N888) );
  ANDN U7510 ( .B(out[871]), .A(rst), .Z(N889) );
  ANDN U7511 ( .B(out[71]), .A(rst), .Z(N89) );
  ANDN U7512 ( .B(out[872]), .A(rst), .Z(N890) );
  ANDN U7513 ( .B(out[873]), .A(rst), .Z(N891) );
  ANDN U7514 ( .B(out[874]), .A(rst), .Z(N892) );
  ANDN U7515 ( .B(out[875]), .A(rst), .Z(N893) );
  ANDN U7516 ( .B(out[876]), .A(rst), .Z(N894) );
  ANDN U7517 ( .B(out[877]), .A(rst), .Z(N895) );
  ANDN U7518 ( .B(out[878]), .A(rst), .Z(N896) );
  ANDN U7519 ( .B(out[879]), .A(rst), .Z(N897) );
  ANDN U7520 ( .B(out[880]), .A(rst), .Z(N898) );
  ANDN U7521 ( .B(out[881]), .A(rst), .Z(N899) );
  ANDN U7522 ( .B(rc_i[2]), .A(rst), .Z(N9) );
  ANDN U7523 ( .B(out[72]), .A(rst), .Z(N90) );
  ANDN U7524 ( .B(out[882]), .A(rst), .Z(N900) );
  ANDN U7525 ( .B(out[883]), .A(rst), .Z(N901) );
  ANDN U7526 ( .B(out[884]), .A(rst), .Z(N902) );
  ANDN U7527 ( .B(out[885]), .A(rst), .Z(N903) );
  ANDN U7528 ( .B(out[886]), .A(rst), .Z(N904) );
  ANDN U7529 ( .B(out[887]), .A(rst), .Z(N905) );
  ANDN U7530 ( .B(out[888]), .A(rst), .Z(N906) );
  ANDN U7531 ( .B(out[889]), .A(rst), .Z(N907) );
  ANDN U7532 ( .B(out[890]), .A(rst), .Z(N908) );
  ANDN U7533 ( .B(out[891]), .A(rst), .Z(N909) );
  ANDN U7534 ( .B(out[73]), .A(rst), .Z(N91) );
  ANDN U7535 ( .B(out[892]), .A(rst), .Z(N910) );
  ANDN U7536 ( .B(out[893]), .A(rst), .Z(N911) );
  ANDN U7537 ( .B(out[894]), .A(rst), .Z(N912) );
  ANDN U7538 ( .B(out[895]), .A(rst), .Z(N913) );
  ANDN U7539 ( .B(out[896]), .A(rst), .Z(N914) );
  ANDN U7540 ( .B(out[897]), .A(rst), .Z(N915) );
  ANDN U7541 ( .B(out[898]), .A(rst), .Z(N916) );
  ANDN U7542 ( .B(out[899]), .A(rst), .Z(N917) );
  ANDN U7543 ( .B(out[900]), .A(rst), .Z(N918) );
  ANDN U7544 ( .B(out[901]), .A(rst), .Z(N919) );
  ANDN U7545 ( .B(out[74]), .A(rst), .Z(N92) );
  ANDN U7546 ( .B(out[902]), .A(rst), .Z(N920) );
  ANDN U7547 ( .B(out[903]), .A(rst), .Z(N921) );
  ANDN U7548 ( .B(out[904]), .A(rst), .Z(N922) );
  ANDN U7549 ( .B(out[905]), .A(rst), .Z(N923) );
  ANDN U7550 ( .B(out[906]), .A(rst), .Z(N924) );
  ANDN U7551 ( .B(out[907]), .A(rst), .Z(N925) );
  ANDN U7552 ( .B(out[908]), .A(rst), .Z(N926) );
  ANDN U7553 ( .B(out[909]), .A(rst), .Z(N927) );
  ANDN U7554 ( .B(out[910]), .A(rst), .Z(N928) );
  ANDN U7555 ( .B(out[911]), .A(rst), .Z(N929) );
  ANDN U7556 ( .B(out[75]), .A(rst), .Z(N93) );
  ANDN U7557 ( .B(out[912]), .A(rst), .Z(N930) );
  ANDN U7558 ( .B(out[913]), .A(rst), .Z(N931) );
  ANDN U7559 ( .B(out[914]), .A(rst), .Z(N932) );
  ANDN U7560 ( .B(out[915]), .A(rst), .Z(N933) );
  ANDN U7561 ( .B(out[916]), .A(rst), .Z(N934) );
  ANDN U7562 ( .B(out[917]), .A(rst), .Z(N935) );
  ANDN U7563 ( .B(out[918]), .A(rst), .Z(N936) );
  ANDN U7564 ( .B(out[919]), .A(rst), .Z(N937) );
  ANDN U7565 ( .B(out[920]), .A(rst), .Z(N938) );
  ANDN U7566 ( .B(out[921]), .A(rst), .Z(N939) );
  ANDN U7567 ( .B(out[76]), .A(rst), .Z(N94) );
  ANDN U7568 ( .B(out[922]), .A(rst), .Z(N940) );
  ANDN U7569 ( .B(out[923]), .A(rst), .Z(N941) );
  ANDN U7570 ( .B(out[924]), .A(rst), .Z(N942) );
  ANDN U7571 ( .B(out[925]), .A(rst), .Z(N943) );
  ANDN U7572 ( .B(out[926]), .A(rst), .Z(N944) );
  ANDN U7573 ( .B(out[927]), .A(rst), .Z(N945) );
  ANDN U7574 ( .B(out[928]), .A(rst), .Z(N946) );
  ANDN U7575 ( .B(out[929]), .A(rst), .Z(N947) );
  ANDN U7576 ( .B(out[930]), .A(rst), .Z(N948) );
  ANDN U7577 ( .B(out[931]), .A(rst), .Z(N949) );
  ANDN U7578 ( .B(out[77]), .A(rst), .Z(N95) );
  ANDN U7579 ( .B(out[932]), .A(rst), .Z(N950) );
  ANDN U7580 ( .B(out[933]), .A(rst), .Z(N951) );
  ANDN U7581 ( .B(out[934]), .A(rst), .Z(N952) );
  ANDN U7582 ( .B(out[935]), .A(rst), .Z(N953) );
  ANDN U7583 ( .B(out[936]), .A(rst), .Z(N954) );
  ANDN U7584 ( .B(out[937]), .A(rst), .Z(N955) );
  ANDN U7585 ( .B(out[938]), .A(rst), .Z(N956) );
  ANDN U7586 ( .B(out[939]), .A(rst), .Z(N957) );
  ANDN U7587 ( .B(out[940]), .A(rst), .Z(N958) );
  ANDN U7588 ( .B(out[941]), .A(rst), .Z(N959) );
  ANDN U7589 ( .B(out[78]), .A(rst), .Z(N96) );
  ANDN U7590 ( .B(out[942]), .A(rst), .Z(N960) );
  ANDN U7591 ( .B(out[943]), .A(rst), .Z(N961) );
  ANDN U7592 ( .B(out[944]), .A(rst), .Z(N962) );
  ANDN U7593 ( .B(out[945]), .A(rst), .Z(N963) );
  ANDN U7594 ( .B(out[946]), .A(rst), .Z(N964) );
  ANDN U7595 ( .B(out[947]), .A(rst), .Z(N965) );
  ANDN U7596 ( .B(out[948]), .A(rst), .Z(N966) );
  ANDN U7597 ( .B(out[949]), .A(rst), .Z(N967) );
  ANDN U7598 ( .B(out[950]), .A(rst), .Z(N968) );
  ANDN U7599 ( .B(out[951]), .A(rst), .Z(N969) );
  ANDN U7600 ( .B(out[79]), .A(rst), .Z(N97) );
  ANDN U7601 ( .B(out[952]), .A(rst), .Z(N970) );
  ANDN U7602 ( .B(out[953]), .A(rst), .Z(N971) );
  ANDN U7603 ( .B(out[954]), .A(rst), .Z(N972) );
  ANDN U7604 ( .B(out[955]), .A(rst), .Z(N973) );
  ANDN U7605 ( .B(out[956]), .A(rst), .Z(N974) );
  ANDN U7606 ( .B(out[957]), .A(rst), .Z(N975) );
  ANDN U7607 ( .B(out[958]), .A(rst), .Z(N976) );
  ANDN U7608 ( .B(out[959]), .A(rst), .Z(N977) );
  ANDN U7609 ( .B(out[960]), .A(rst), .Z(N978) );
  ANDN U7610 ( .B(out[961]), .A(rst), .Z(N979) );
  ANDN U7611 ( .B(out[80]), .A(rst), .Z(N98) );
  ANDN U7612 ( .B(out[962]), .A(rst), .Z(N980) );
  ANDN U7613 ( .B(out[963]), .A(rst), .Z(N981) );
  ANDN U7614 ( .B(out[964]), .A(rst), .Z(N982) );
  ANDN U7615 ( .B(out[965]), .A(rst), .Z(N983) );
  ANDN U7616 ( .B(out[966]), .A(rst), .Z(N984) );
  ANDN U7617 ( .B(out[967]), .A(rst), .Z(N985) );
  ANDN U7618 ( .B(out[968]), .A(rst), .Z(N986) );
  ANDN U7619 ( .B(out[969]), .A(rst), .Z(N987) );
  ANDN U7620 ( .B(out[970]), .A(rst), .Z(N988) );
  ANDN U7621 ( .B(out[971]), .A(rst), .Z(N989) );
  ANDN U7622 ( .B(out[81]), .A(rst), .Z(N99) );
  ANDN U7623 ( .B(out[972]), .A(rst), .Z(N990) );
  ANDN U7624 ( .B(out[973]), .A(rst), .Z(N991) );
  ANDN U7625 ( .B(out[974]), .A(rst), .Z(N992) );
  ANDN U7626 ( .B(out[975]), .A(rst), .Z(N993) );
  ANDN U7627 ( .B(out[976]), .A(rst), .Z(N994) );
  ANDN U7628 ( .B(out[977]), .A(rst), .Z(N995) );
  ANDN U7629 ( .B(out[978]), .A(rst), .Z(N996) );
  ANDN U7630 ( .B(out[979]), .A(rst), .Z(N997) );
  ANDN U7631 ( .B(out[980]), .A(rst), .Z(N998) );
  ANDN U7632 ( .B(out[981]), .A(rst), .Z(N999) );
  NOR U7633 ( .A(rc_i[6]), .B(rc_i[9]), .Z(n2794) );
  ANDN U7634 ( .B(n2794), .A(rc_i[8]), .Z(n2812) );
  NOR U7635 ( .A(rc_i[1]), .B(rc_i[4]), .Z(n2795) );
  AND U7636 ( .A(n2812), .B(n2795), .Z(n2793) );
  NANDN U7637 ( .A(rc_i[2]), .B(n2793), .Z(\RCONST[0].rconst_/N18 ) );
  ANDN U7638 ( .B(n2794), .A(rc_i[5]), .Z(n2809) );
  NOR U7639 ( .A(rc_i[2]), .B(rc_i[7]), .Z(n2796) );
  AND U7640 ( .A(n2795), .B(n2796), .Z(n2798) );
  NAND U7641 ( .A(n2809), .B(n2798), .Z(\RCONST[0].rconst_/N28 ) );
  NOR U7642 ( .A(rc_i[6]), .B(rc_i[3]), .Z(n2797) );
  NAND U7643 ( .A(n2797), .B(n2796), .Z(\RCONST[1].rconst_/N10 ) );
  ANDN U7644 ( .B(n2797), .A(rc_i[10]), .Z(n2802) );
  NAND U7645 ( .A(n2802), .B(n2798), .Z(\RCONST[0].rconst_/N37 ) );
  NOR U7646 ( .A(rc_i[7]), .B(rc_i[3]), .Z(n2799) );
  ANDN U7647 ( .B(n2799), .A(rc_i[1]), .Z(n2800) );
  ANDN U7648 ( .B(n2800), .A(rc_i[10]), .Z(n2804) );
  NANDN U7649 ( .A(rc_i[8]), .B(n2804), .Z(\RCONST[0].rconst_/N67 ) );
  NOR U7650 ( .A(rc_i[2]), .B(\RCONST[0].rconst_/N67 ), .Z(n2801) );
  NAND U7651 ( .A(n2809), .B(n2801), .Z(\RCONST[0].rconst_/N48 ) );
  NOR U7652 ( .A(rc_i[5]), .B(rc_i[11]), .Z(n2806) );
  NAND U7653 ( .A(n2806), .B(n2802), .Z(\RCONST[0].rconst_/N57 ) );
  NOR U7654 ( .A(rc_i[7]), .B(rc_i[0]), .Z(n2805) );
  ANDN U7655 ( .B(n2805), .A(\RCONST[0].rconst_/N57 ), .Z(n2803) );
  NANDN U7656 ( .A(rc_i[2]), .B(n2803), .Z(\rc[0][0] ) );
  ANDN U7657 ( .B(n2804), .A(rc_i[11]), .Z(n2813) );
  NANDN U7658 ( .A(rc_i[0]), .B(n2813), .Z(\rc[1][15] ) );
  NAND U7659 ( .A(n2809), .B(n2805), .Z(\rc[1][1] ) );
  ANDN U7660 ( .B(n2806), .A(rc_i[2]), .Z(n2807) );
  ANDN U7661 ( .B(n2807), .A(rc_i[1]), .Z(n2808) );
  NANDN U7662 ( .A(rc_i[9]), .B(n2808), .Z(\rc[1][31] ) );
  ANDN U7663 ( .B(n2809), .A(rc_i[3]), .Z(n2810) );
  ANDN U7664 ( .B(n2810), .A(rc_i[4]), .Z(n2811) );
  NANDN U7665 ( .A(rc_i[11]), .B(n2811), .Z(\rc[1][3] ) );
  NAND U7666 ( .A(n2813), .B(n2812), .Z(\rc[1][63] ) );
  NOR U7667 ( .A(rc_i[0]), .B(rc_i[4]), .Z(n2814) );
  ANDN U7668 ( .B(n2814), .A(rc_i[10]), .Z(n2815) );
  ANDN U7669 ( .B(n2815), .A(rc_i[8]), .Z(n2816) );
  NANDN U7670 ( .A(rc_i[6]), .B(n2816), .Z(\rc[1][7] ) );
  NAND U7671 ( .A(init), .B(round_reg[0]), .Z(n2818) );
  NANDN U7672 ( .A(init), .B(in[0]), .Z(n2817) );
  NAND U7673 ( .A(n2818), .B(n2817), .Z(\round_in[0][0] ) );
  AND U7674 ( .A(round_reg[1000]), .B(init), .Z(\round_in[0][1000] ) );
  AND U7675 ( .A(round_reg[1001]), .B(init), .Z(\round_in[0][1001] ) );
  AND U7676 ( .A(round_reg[1002]), .B(init), .Z(\round_in[0][1002] ) );
  AND U7677 ( .A(round_reg[1003]), .B(init), .Z(\round_in[0][1003] ) );
  AND U7678 ( .A(round_reg[1004]), .B(init), .Z(\round_in[0][1004] ) );
  AND U7679 ( .A(round_reg[1005]), .B(init), .Z(\round_in[0][1005] ) );
  AND U7680 ( .A(round_reg[1006]), .B(init), .Z(\round_in[0][1006] ) );
  AND U7681 ( .A(round_reg[1007]), .B(init), .Z(\round_in[0][1007] ) );
  AND U7682 ( .A(round_reg[1008]), .B(init), .Z(\round_in[0][1008] ) );
  AND U7683 ( .A(round_reg[1009]), .B(init), .Z(\round_in[0][1009] ) );
  NAND U7684 ( .A(init), .B(round_reg[100]), .Z(n2820) );
  NANDN U7685 ( .A(init), .B(in[100]), .Z(n2819) );
  NAND U7686 ( .A(n2820), .B(n2819), .Z(\round_in[0][100] ) );
  AND U7687 ( .A(round_reg[1010]), .B(init), .Z(\round_in[0][1010] ) );
  AND U7688 ( .A(round_reg[1011]), .B(init), .Z(\round_in[0][1011] ) );
  AND U7689 ( .A(round_reg[1012]), .B(init), .Z(\round_in[0][1012] ) );
  AND U7690 ( .A(round_reg[1013]), .B(init), .Z(\round_in[0][1013] ) );
  AND U7691 ( .A(round_reg[1014]), .B(init), .Z(\round_in[0][1014] ) );
  AND U7692 ( .A(round_reg[1015]), .B(init), .Z(\round_in[0][1015] ) );
  AND U7693 ( .A(round_reg[1016]), .B(init), .Z(\round_in[0][1016] ) );
  AND U7694 ( .A(round_reg[1017]), .B(init), .Z(\round_in[0][1017] ) );
  AND U7695 ( .A(round_reg[1018]), .B(init), .Z(\round_in[0][1018] ) );
  AND U7696 ( .A(round_reg[1019]), .B(init), .Z(\round_in[0][1019] ) );
  NAND U7697 ( .A(init), .B(round_reg[101]), .Z(n2822) );
  NANDN U7698 ( .A(init), .B(in[101]), .Z(n2821) );
  NAND U7699 ( .A(n2822), .B(n2821), .Z(\round_in[0][101] ) );
  AND U7700 ( .A(round_reg[1020]), .B(init), .Z(\round_in[0][1020] ) );
  AND U7701 ( .A(round_reg[1021]), .B(init), .Z(\round_in[0][1021] ) );
  AND U7702 ( .A(round_reg[1022]), .B(init), .Z(\round_in[0][1022] ) );
  AND U7703 ( .A(round_reg[1023]), .B(init), .Z(\round_in[0][1023] ) );
  AND U7704 ( .A(round_reg[1024]), .B(init), .Z(\round_in[0][1024] ) );
  AND U7705 ( .A(round_reg[1025]), .B(init), .Z(\round_in[0][1025] ) );
  AND U7706 ( .A(round_reg[1026]), .B(init), .Z(\round_in[0][1026] ) );
  AND U7707 ( .A(round_reg[1027]), .B(init), .Z(\round_in[0][1027] ) );
  AND U7708 ( .A(round_reg[1028]), .B(init), .Z(\round_in[0][1028] ) );
  AND U7709 ( .A(round_reg[1029]), .B(init), .Z(\round_in[0][1029] ) );
  NAND U7710 ( .A(init), .B(round_reg[102]), .Z(n2824) );
  NANDN U7711 ( .A(init), .B(in[102]), .Z(n2823) );
  NAND U7712 ( .A(n2824), .B(n2823), .Z(\round_in[0][102] ) );
  AND U7713 ( .A(round_reg[1030]), .B(init), .Z(\round_in[0][1030] ) );
  AND U7714 ( .A(round_reg[1031]), .B(init), .Z(\round_in[0][1031] ) );
  AND U7715 ( .A(round_reg[1032]), .B(init), .Z(\round_in[0][1032] ) );
  AND U7716 ( .A(round_reg[1033]), .B(init), .Z(\round_in[0][1033] ) );
  AND U7717 ( .A(round_reg[1034]), .B(init), .Z(\round_in[0][1034] ) );
  AND U7718 ( .A(round_reg[1035]), .B(init), .Z(\round_in[0][1035] ) );
  AND U7719 ( .A(round_reg[1036]), .B(init), .Z(\round_in[0][1036] ) );
  AND U7720 ( .A(round_reg[1037]), .B(init), .Z(\round_in[0][1037] ) );
  AND U7721 ( .A(round_reg[1038]), .B(init), .Z(\round_in[0][1038] ) );
  AND U7722 ( .A(round_reg[1039]), .B(init), .Z(\round_in[0][1039] ) );
  NAND U7723 ( .A(init), .B(round_reg[103]), .Z(n2826) );
  NANDN U7724 ( .A(init), .B(in[103]), .Z(n2825) );
  NAND U7725 ( .A(n2826), .B(n2825), .Z(\round_in[0][103] ) );
  AND U7726 ( .A(round_reg[1040]), .B(init), .Z(\round_in[0][1040] ) );
  AND U7727 ( .A(round_reg[1041]), .B(init), .Z(\round_in[0][1041] ) );
  AND U7728 ( .A(round_reg[1042]), .B(init), .Z(\round_in[0][1042] ) );
  AND U7729 ( .A(round_reg[1043]), .B(init), .Z(\round_in[0][1043] ) );
  AND U7730 ( .A(round_reg[1044]), .B(init), .Z(\round_in[0][1044] ) );
  AND U7731 ( .A(round_reg[1045]), .B(init), .Z(\round_in[0][1045] ) );
  AND U7732 ( .A(round_reg[1046]), .B(init), .Z(\round_in[0][1046] ) );
  AND U7733 ( .A(round_reg[1047]), .B(init), .Z(\round_in[0][1047] ) );
  AND U7734 ( .A(round_reg[1048]), .B(init), .Z(\round_in[0][1048] ) );
  AND U7735 ( .A(round_reg[1049]), .B(init), .Z(\round_in[0][1049] ) );
  NAND U7736 ( .A(init), .B(round_reg[104]), .Z(n2828) );
  NANDN U7737 ( .A(init), .B(in[104]), .Z(n2827) );
  NAND U7738 ( .A(n2828), .B(n2827), .Z(\round_in[0][104] ) );
  AND U7739 ( .A(round_reg[1050]), .B(init), .Z(\round_in[0][1050] ) );
  AND U7740 ( .A(round_reg[1051]), .B(init), .Z(\round_in[0][1051] ) );
  AND U7741 ( .A(round_reg[1052]), .B(init), .Z(\round_in[0][1052] ) );
  AND U7742 ( .A(round_reg[1053]), .B(init), .Z(\round_in[0][1053] ) );
  AND U7743 ( .A(round_reg[1054]), .B(init), .Z(\round_in[0][1054] ) );
  AND U7744 ( .A(round_reg[1055]), .B(init), .Z(\round_in[0][1055] ) );
  AND U7745 ( .A(round_reg[1056]), .B(init), .Z(\round_in[0][1056] ) );
  AND U7746 ( .A(round_reg[1057]), .B(init), .Z(\round_in[0][1057] ) );
  AND U7747 ( .A(round_reg[1058]), .B(init), .Z(\round_in[0][1058] ) );
  AND U7748 ( .A(round_reg[1059]), .B(init), .Z(\round_in[0][1059] ) );
  NAND U7749 ( .A(init), .B(round_reg[105]), .Z(n2830) );
  NANDN U7750 ( .A(init), .B(in[105]), .Z(n2829) );
  NAND U7751 ( .A(n2830), .B(n2829), .Z(\round_in[0][105] ) );
  AND U7752 ( .A(round_reg[1060]), .B(init), .Z(\round_in[0][1060] ) );
  AND U7753 ( .A(round_reg[1061]), .B(init), .Z(\round_in[0][1061] ) );
  AND U7754 ( .A(round_reg[1062]), .B(init), .Z(\round_in[0][1062] ) );
  AND U7755 ( .A(round_reg[1063]), .B(init), .Z(\round_in[0][1063] ) );
  AND U7756 ( .A(round_reg[1064]), .B(init), .Z(\round_in[0][1064] ) );
  AND U7757 ( .A(round_reg[1065]), .B(init), .Z(\round_in[0][1065] ) );
  AND U7758 ( .A(round_reg[1066]), .B(init), .Z(\round_in[0][1066] ) );
  AND U7759 ( .A(round_reg[1067]), .B(init), .Z(\round_in[0][1067] ) );
  AND U7760 ( .A(round_reg[1068]), .B(init), .Z(\round_in[0][1068] ) );
  AND U7761 ( .A(round_reg[1069]), .B(init), .Z(\round_in[0][1069] ) );
  NAND U7762 ( .A(init), .B(round_reg[106]), .Z(n2832) );
  NANDN U7763 ( .A(init), .B(in[106]), .Z(n2831) );
  NAND U7764 ( .A(n2832), .B(n2831), .Z(\round_in[0][106] ) );
  AND U7765 ( .A(round_reg[1070]), .B(init), .Z(\round_in[0][1070] ) );
  AND U7766 ( .A(round_reg[1071]), .B(init), .Z(\round_in[0][1071] ) );
  AND U7767 ( .A(round_reg[1072]), .B(init), .Z(\round_in[0][1072] ) );
  AND U7768 ( .A(round_reg[1073]), .B(init), .Z(\round_in[0][1073] ) );
  AND U7769 ( .A(round_reg[1074]), .B(init), .Z(\round_in[0][1074] ) );
  AND U7770 ( .A(round_reg[1075]), .B(init), .Z(\round_in[0][1075] ) );
  AND U7771 ( .A(round_reg[1076]), .B(init), .Z(\round_in[0][1076] ) );
  AND U7772 ( .A(round_reg[1077]), .B(init), .Z(\round_in[0][1077] ) );
  AND U7773 ( .A(round_reg[1078]), .B(init), .Z(\round_in[0][1078] ) );
  AND U7774 ( .A(round_reg[1079]), .B(init), .Z(\round_in[0][1079] ) );
  NAND U7775 ( .A(init), .B(round_reg[107]), .Z(n2834) );
  NANDN U7776 ( .A(init), .B(in[107]), .Z(n2833) );
  NAND U7777 ( .A(n2834), .B(n2833), .Z(\round_in[0][107] ) );
  AND U7778 ( .A(round_reg[1080]), .B(init), .Z(\round_in[0][1080] ) );
  AND U7779 ( .A(round_reg[1081]), .B(init), .Z(\round_in[0][1081] ) );
  AND U7780 ( .A(round_reg[1082]), .B(init), .Z(\round_in[0][1082] ) );
  AND U7781 ( .A(round_reg[1083]), .B(init), .Z(\round_in[0][1083] ) );
  AND U7782 ( .A(round_reg[1084]), .B(init), .Z(\round_in[0][1084] ) );
  AND U7783 ( .A(round_reg[1085]), .B(init), .Z(\round_in[0][1085] ) );
  AND U7784 ( .A(round_reg[1086]), .B(init), .Z(\round_in[0][1086] ) );
  AND U7785 ( .A(round_reg[1087]), .B(init), .Z(\round_in[0][1087] ) );
  AND U7786 ( .A(round_reg[1088]), .B(init), .Z(\round_in[0][1088] ) );
  AND U7787 ( .A(round_reg[1089]), .B(init), .Z(\round_in[0][1089] ) );
  NAND U7788 ( .A(init), .B(round_reg[108]), .Z(n2836) );
  NANDN U7789 ( .A(init), .B(in[108]), .Z(n2835) );
  NAND U7790 ( .A(n2836), .B(n2835), .Z(\round_in[0][108] ) );
  AND U7791 ( .A(round_reg[1090]), .B(init), .Z(\round_in[0][1090] ) );
  AND U7792 ( .A(round_reg[1091]), .B(init), .Z(\round_in[0][1091] ) );
  AND U7793 ( .A(round_reg[1092]), .B(init), .Z(\round_in[0][1092] ) );
  AND U7794 ( .A(round_reg[1093]), .B(init), .Z(\round_in[0][1093] ) );
  AND U7795 ( .A(round_reg[1094]), .B(init), .Z(\round_in[0][1094] ) );
  AND U7796 ( .A(round_reg[1095]), .B(init), .Z(\round_in[0][1095] ) );
  AND U7797 ( .A(round_reg[1096]), .B(init), .Z(\round_in[0][1096] ) );
  AND U7798 ( .A(round_reg[1097]), .B(init), .Z(\round_in[0][1097] ) );
  AND U7799 ( .A(round_reg[1098]), .B(init), .Z(\round_in[0][1098] ) );
  AND U7800 ( .A(round_reg[1099]), .B(init), .Z(\round_in[0][1099] ) );
  NAND U7801 ( .A(init), .B(round_reg[109]), .Z(n2838) );
  NANDN U7802 ( .A(init), .B(in[109]), .Z(n2837) );
  NAND U7803 ( .A(n2838), .B(n2837), .Z(\round_in[0][109] ) );
  NAND U7804 ( .A(init), .B(round_reg[10]), .Z(n2840) );
  NANDN U7805 ( .A(init), .B(in[10]), .Z(n2839) );
  NAND U7806 ( .A(n2840), .B(n2839), .Z(\round_in[0][10] ) );
  AND U7807 ( .A(round_reg[1100]), .B(init), .Z(\round_in[0][1100] ) );
  AND U7808 ( .A(round_reg[1101]), .B(init), .Z(\round_in[0][1101] ) );
  AND U7809 ( .A(round_reg[1102]), .B(init), .Z(\round_in[0][1102] ) );
  AND U7810 ( .A(round_reg[1103]), .B(init), .Z(\round_in[0][1103] ) );
  AND U7811 ( .A(round_reg[1104]), .B(init), .Z(\round_in[0][1104] ) );
  AND U7812 ( .A(round_reg[1105]), .B(init), .Z(\round_in[0][1105] ) );
  AND U7813 ( .A(round_reg[1106]), .B(init), .Z(\round_in[0][1106] ) );
  AND U7814 ( .A(round_reg[1107]), .B(init), .Z(\round_in[0][1107] ) );
  AND U7815 ( .A(round_reg[1108]), .B(init), .Z(\round_in[0][1108] ) );
  AND U7816 ( .A(round_reg[1109]), .B(init), .Z(\round_in[0][1109] ) );
  NAND U7817 ( .A(init), .B(round_reg[110]), .Z(n2842) );
  NANDN U7818 ( .A(init), .B(in[110]), .Z(n2841) );
  NAND U7819 ( .A(n2842), .B(n2841), .Z(\round_in[0][110] ) );
  AND U7820 ( .A(round_reg[1110]), .B(init), .Z(\round_in[0][1110] ) );
  AND U7821 ( .A(round_reg[1111]), .B(init), .Z(\round_in[0][1111] ) );
  AND U7822 ( .A(round_reg[1112]), .B(init), .Z(\round_in[0][1112] ) );
  AND U7823 ( .A(round_reg[1113]), .B(init), .Z(\round_in[0][1113] ) );
  AND U7824 ( .A(round_reg[1114]), .B(init), .Z(\round_in[0][1114] ) );
  AND U7825 ( .A(round_reg[1115]), .B(init), .Z(\round_in[0][1115] ) );
  AND U7826 ( .A(round_reg[1116]), .B(init), .Z(\round_in[0][1116] ) );
  AND U7827 ( .A(round_reg[1117]), .B(init), .Z(\round_in[0][1117] ) );
  AND U7828 ( .A(round_reg[1118]), .B(init), .Z(\round_in[0][1118] ) );
  AND U7829 ( .A(round_reg[1119]), .B(init), .Z(\round_in[0][1119] ) );
  NAND U7830 ( .A(init), .B(round_reg[111]), .Z(n2844) );
  NANDN U7831 ( .A(init), .B(in[111]), .Z(n2843) );
  NAND U7832 ( .A(n2844), .B(n2843), .Z(\round_in[0][111] ) );
  AND U7833 ( .A(round_reg[1120]), .B(init), .Z(\round_in[0][1120] ) );
  AND U7834 ( .A(round_reg[1121]), .B(init), .Z(\round_in[0][1121] ) );
  AND U7835 ( .A(round_reg[1122]), .B(init), .Z(\round_in[0][1122] ) );
  AND U7836 ( .A(round_reg[1123]), .B(init), .Z(\round_in[0][1123] ) );
  AND U7837 ( .A(round_reg[1124]), .B(init), .Z(\round_in[0][1124] ) );
  AND U7838 ( .A(round_reg[1125]), .B(init), .Z(\round_in[0][1125] ) );
  AND U7839 ( .A(round_reg[1126]), .B(init), .Z(\round_in[0][1126] ) );
  AND U7840 ( .A(round_reg[1127]), .B(init), .Z(\round_in[0][1127] ) );
  AND U7841 ( .A(round_reg[1128]), .B(init), .Z(\round_in[0][1128] ) );
  AND U7842 ( .A(round_reg[1129]), .B(init), .Z(\round_in[0][1129] ) );
  NAND U7843 ( .A(init), .B(round_reg[112]), .Z(n2846) );
  NANDN U7844 ( .A(init), .B(in[112]), .Z(n2845) );
  NAND U7845 ( .A(n2846), .B(n2845), .Z(\round_in[0][112] ) );
  AND U7846 ( .A(round_reg[1130]), .B(init), .Z(\round_in[0][1130] ) );
  AND U7847 ( .A(round_reg[1131]), .B(init), .Z(\round_in[0][1131] ) );
  AND U7848 ( .A(round_reg[1132]), .B(init), .Z(\round_in[0][1132] ) );
  AND U7849 ( .A(round_reg[1133]), .B(init), .Z(\round_in[0][1133] ) );
  AND U7850 ( .A(round_reg[1134]), .B(init), .Z(\round_in[0][1134] ) );
  AND U7851 ( .A(round_reg[1135]), .B(init), .Z(\round_in[0][1135] ) );
  AND U7852 ( .A(round_reg[1136]), .B(init), .Z(\round_in[0][1136] ) );
  AND U7853 ( .A(round_reg[1137]), .B(init), .Z(\round_in[0][1137] ) );
  AND U7854 ( .A(round_reg[1138]), .B(init), .Z(\round_in[0][1138] ) );
  AND U7855 ( .A(round_reg[1139]), .B(init), .Z(\round_in[0][1139] ) );
  NAND U7856 ( .A(init), .B(round_reg[113]), .Z(n2848) );
  NANDN U7857 ( .A(init), .B(in[113]), .Z(n2847) );
  NAND U7858 ( .A(n2848), .B(n2847), .Z(\round_in[0][113] ) );
  AND U7859 ( .A(round_reg[1140]), .B(init), .Z(\round_in[0][1140] ) );
  AND U7860 ( .A(round_reg[1141]), .B(init), .Z(\round_in[0][1141] ) );
  AND U7861 ( .A(round_reg[1142]), .B(init), .Z(\round_in[0][1142] ) );
  AND U7862 ( .A(round_reg[1143]), .B(init), .Z(\round_in[0][1143] ) );
  AND U7863 ( .A(round_reg[1144]), .B(init), .Z(\round_in[0][1144] ) );
  AND U7864 ( .A(round_reg[1145]), .B(init), .Z(\round_in[0][1145] ) );
  AND U7865 ( .A(round_reg[1146]), .B(init), .Z(\round_in[0][1146] ) );
  AND U7866 ( .A(round_reg[1147]), .B(init), .Z(\round_in[0][1147] ) );
  AND U7867 ( .A(round_reg[1148]), .B(init), .Z(\round_in[0][1148] ) );
  AND U7868 ( .A(round_reg[1149]), .B(init), .Z(\round_in[0][1149] ) );
  NAND U7869 ( .A(init), .B(round_reg[114]), .Z(n2850) );
  NANDN U7870 ( .A(init), .B(in[114]), .Z(n2849) );
  NAND U7871 ( .A(n2850), .B(n2849), .Z(\round_in[0][114] ) );
  AND U7872 ( .A(round_reg[1150]), .B(init), .Z(\round_in[0][1150] ) );
  AND U7873 ( .A(round_reg[1151]), .B(init), .Z(\round_in[0][1151] ) );
  AND U7874 ( .A(round_reg[1152]), .B(init), .Z(\round_in[0][1152] ) );
  AND U7875 ( .A(round_reg[1153]), .B(init), .Z(\round_in[0][1153] ) );
  AND U7876 ( .A(round_reg[1154]), .B(init), .Z(\round_in[0][1154] ) );
  AND U7877 ( .A(round_reg[1155]), .B(init), .Z(\round_in[0][1155] ) );
  AND U7878 ( .A(round_reg[1156]), .B(init), .Z(\round_in[0][1156] ) );
  AND U7879 ( .A(round_reg[1157]), .B(init), .Z(\round_in[0][1157] ) );
  AND U7880 ( .A(round_reg[1158]), .B(init), .Z(\round_in[0][1158] ) );
  AND U7881 ( .A(round_reg[1159]), .B(init), .Z(\round_in[0][1159] ) );
  NAND U7882 ( .A(init), .B(round_reg[115]), .Z(n2852) );
  NANDN U7883 ( .A(init), .B(in[115]), .Z(n2851) );
  NAND U7884 ( .A(n2852), .B(n2851), .Z(\round_in[0][115] ) );
  AND U7885 ( .A(round_reg[1160]), .B(init), .Z(\round_in[0][1160] ) );
  AND U7886 ( .A(round_reg[1161]), .B(init), .Z(\round_in[0][1161] ) );
  AND U7887 ( .A(round_reg[1162]), .B(init), .Z(\round_in[0][1162] ) );
  AND U7888 ( .A(round_reg[1163]), .B(init), .Z(\round_in[0][1163] ) );
  AND U7889 ( .A(round_reg[1164]), .B(init), .Z(\round_in[0][1164] ) );
  AND U7890 ( .A(round_reg[1165]), .B(init), .Z(\round_in[0][1165] ) );
  AND U7891 ( .A(round_reg[1166]), .B(init), .Z(\round_in[0][1166] ) );
  AND U7892 ( .A(round_reg[1167]), .B(init), .Z(\round_in[0][1167] ) );
  AND U7893 ( .A(round_reg[1168]), .B(init), .Z(\round_in[0][1168] ) );
  AND U7894 ( .A(round_reg[1169]), .B(init), .Z(\round_in[0][1169] ) );
  NAND U7895 ( .A(init), .B(round_reg[116]), .Z(n2854) );
  NANDN U7896 ( .A(init), .B(in[116]), .Z(n2853) );
  NAND U7897 ( .A(n2854), .B(n2853), .Z(\round_in[0][116] ) );
  AND U7898 ( .A(round_reg[1170]), .B(init), .Z(\round_in[0][1170] ) );
  AND U7899 ( .A(round_reg[1171]), .B(init), .Z(\round_in[0][1171] ) );
  AND U7900 ( .A(round_reg[1172]), .B(init), .Z(\round_in[0][1172] ) );
  AND U7901 ( .A(round_reg[1173]), .B(init), .Z(\round_in[0][1173] ) );
  AND U7902 ( .A(round_reg[1174]), .B(init), .Z(\round_in[0][1174] ) );
  AND U7903 ( .A(round_reg[1175]), .B(init), .Z(\round_in[0][1175] ) );
  AND U7904 ( .A(round_reg[1176]), .B(init), .Z(\round_in[0][1176] ) );
  AND U7905 ( .A(round_reg[1177]), .B(init), .Z(\round_in[0][1177] ) );
  AND U7906 ( .A(round_reg[1178]), .B(init), .Z(\round_in[0][1178] ) );
  AND U7907 ( .A(round_reg[1179]), .B(init), .Z(\round_in[0][1179] ) );
  NAND U7908 ( .A(init), .B(round_reg[117]), .Z(n2856) );
  NANDN U7909 ( .A(init), .B(in[117]), .Z(n2855) );
  NAND U7910 ( .A(n2856), .B(n2855), .Z(\round_in[0][117] ) );
  AND U7911 ( .A(round_reg[1180]), .B(init), .Z(\round_in[0][1180] ) );
  AND U7912 ( .A(round_reg[1181]), .B(init), .Z(\round_in[0][1181] ) );
  AND U7913 ( .A(round_reg[1182]), .B(init), .Z(\round_in[0][1182] ) );
  AND U7914 ( .A(round_reg[1183]), .B(init), .Z(\round_in[0][1183] ) );
  AND U7915 ( .A(round_reg[1184]), .B(init), .Z(\round_in[0][1184] ) );
  AND U7916 ( .A(round_reg[1185]), .B(init), .Z(\round_in[0][1185] ) );
  AND U7917 ( .A(round_reg[1186]), .B(init), .Z(\round_in[0][1186] ) );
  AND U7918 ( .A(round_reg[1187]), .B(init), .Z(\round_in[0][1187] ) );
  AND U7919 ( .A(round_reg[1188]), .B(init), .Z(\round_in[0][1188] ) );
  AND U7920 ( .A(round_reg[1189]), .B(init), .Z(\round_in[0][1189] ) );
  NAND U7921 ( .A(init), .B(round_reg[118]), .Z(n2858) );
  NANDN U7922 ( .A(init), .B(in[118]), .Z(n2857) );
  NAND U7923 ( .A(n2858), .B(n2857), .Z(\round_in[0][118] ) );
  AND U7924 ( .A(round_reg[1190]), .B(init), .Z(\round_in[0][1190] ) );
  AND U7925 ( .A(round_reg[1191]), .B(init), .Z(\round_in[0][1191] ) );
  AND U7926 ( .A(round_reg[1192]), .B(init), .Z(\round_in[0][1192] ) );
  AND U7927 ( .A(round_reg[1193]), .B(init), .Z(\round_in[0][1193] ) );
  AND U7928 ( .A(round_reg[1194]), .B(init), .Z(\round_in[0][1194] ) );
  AND U7929 ( .A(round_reg[1195]), .B(init), .Z(\round_in[0][1195] ) );
  AND U7930 ( .A(round_reg[1196]), .B(init), .Z(\round_in[0][1196] ) );
  AND U7931 ( .A(round_reg[1197]), .B(init), .Z(\round_in[0][1197] ) );
  AND U7932 ( .A(round_reg[1198]), .B(init), .Z(\round_in[0][1198] ) );
  AND U7933 ( .A(round_reg[1199]), .B(init), .Z(\round_in[0][1199] ) );
  NAND U7934 ( .A(init), .B(round_reg[119]), .Z(n2860) );
  NANDN U7935 ( .A(init), .B(in[119]), .Z(n2859) );
  NAND U7936 ( .A(n2860), .B(n2859), .Z(\round_in[0][119] ) );
  NAND U7937 ( .A(init), .B(round_reg[11]), .Z(n2862) );
  NANDN U7938 ( .A(init), .B(in[11]), .Z(n2861) );
  NAND U7939 ( .A(n2862), .B(n2861), .Z(\round_in[0][11] ) );
  AND U7940 ( .A(round_reg[1200]), .B(init), .Z(\round_in[0][1200] ) );
  AND U7941 ( .A(round_reg[1201]), .B(init), .Z(\round_in[0][1201] ) );
  AND U7942 ( .A(round_reg[1202]), .B(init), .Z(\round_in[0][1202] ) );
  AND U7943 ( .A(round_reg[1203]), .B(init), .Z(\round_in[0][1203] ) );
  AND U7944 ( .A(round_reg[1204]), .B(init), .Z(\round_in[0][1204] ) );
  AND U7945 ( .A(round_reg[1205]), .B(init), .Z(\round_in[0][1205] ) );
  AND U7946 ( .A(round_reg[1206]), .B(init), .Z(\round_in[0][1206] ) );
  AND U7947 ( .A(round_reg[1207]), .B(init), .Z(\round_in[0][1207] ) );
  AND U7948 ( .A(round_reg[1208]), .B(init), .Z(\round_in[0][1208] ) );
  AND U7949 ( .A(round_reg[1209]), .B(init), .Z(\round_in[0][1209] ) );
  NAND U7950 ( .A(init), .B(round_reg[120]), .Z(n2864) );
  NANDN U7951 ( .A(init), .B(in[120]), .Z(n2863) );
  NAND U7952 ( .A(n2864), .B(n2863), .Z(\round_in[0][120] ) );
  AND U7953 ( .A(round_reg[1210]), .B(init), .Z(\round_in[0][1210] ) );
  AND U7954 ( .A(round_reg[1211]), .B(init), .Z(\round_in[0][1211] ) );
  AND U7955 ( .A(round_reg[1212]), .B(init), .Z(\round_in[0][1212] ) );
  AND U7956 ( .A(round_reg[1213]), .B(init), .Z(\round_in[0][1213] ) );
  AND U7957 ( .A(round_reg[1214]), .B(init), .Z(\round_in[0][1214] ) );
  AND U7958 ( .A(round_reg[1215]), .B(init), .Z(\round_in[0][1215] ) );
  AND U7959 ( .A(round_reg[1216]), .B(init), .Z(\round_in[0][1216] ) );
  AND U7960 ( .A(round_reg[1217]), .B(init), .Z(\round_in[0][1217] ) );
  AND U7961 ( .A(round_reg[1218]), .B(init), .Z(\round_in[0][1218] ) );
  AND U7962 ( .A(round_reg[1219]), .B(init), .Z(\round_in[0][1219] ) );
  NAND U7963 ( .A(init), .B(round_reg[121]), .Z(n2866) );
  NANDN U7964 ( .A(init), .B(in[121]), .Z(n2865) );
  NAND U7965 ( .A(n2866), .B(n2865), .Z(\round_in[0][121] ) );
  AND U7966 ( .A(round_reg[1220]), .B(init), .Z(\round_in[0][1220] ) );
  AND U7967 ( .A(round_reg[1221]), .B(init), .Z(\round_in[0][1221] ) );
  AND U7968 ( .A(round_reg[1222]), .B(init), .Z(\round_in[0][1222] ) );
  AND U7969 ( .A(round_reg[1223]), .B(init), .Z(\round_in[0][1223] ) );
  AND U7970 ( .A(round_reg[1224]), .B(init), .Z(\round_in[0][1224] ) );
  AND U7971 ( .A(round_reg[1225]), .B(init), .Z(\round_in[0][1225] ) );
  AND U7972 ( .A(round_reg[1226]), .B(init), .Z(\round_in[0][1226] ) );
  AND U7973 ( .A(round_reg[1227]), .B(init), .Z(\round_in[0][1227] ) );
  AND U7974 ( .A(round_reg[1228]), .B(init), .Z(\round_in[0][1228] ) );
  AND U7975 ( .A(round_reg[1229]), .B(init), .Z(\round_in[0][1229] ) );
  NAND U7976 ( .A(init), .B(round_reg[122]), .Z(n2868) );
  NANDN U7977 ( .A(init), .B(in[122]), .Z(n2867) );
  NAND U7978 ( .A(n2868), .B(n2867), .Z(\round_in[0][122] ) );
  AND U7979 ( .A(round_reg[1230]), .B(init), .Z(\round_in[0][1230] ) );
  AND U7980 ( .A(round_reg[1231]), .B(init), .Z(\round_in[0][1231] ) );
  AND U7981 ( .A(round_reg[1232]), .B(init), .Z(\round_in[0][1232] ) );
  AND U7982 ( .A(round_reg[1233]), .B(init), .Z(\round_in[0][1233] ) );
  AND U7983 ( .A(round_reg[1234]), .B(init), .Z(\round_in[0][1234] ) );
  AND U7984 ( .A(round_reg[1235]), .B(init), .Z(\round_in[0][1235] ) );
  AND U7985 ( .A(round_reg[1236]), .B(init), .Z(\round_in[0][1236] ) );
  AND U7986 ( .A(round_reg[1237]), .B(init), .Z(\round_in[0][1237] ) );
  AND U7987 ( .A(round_reg[1238]), .B(init), .Z(\round_in[0][1238] ) );
  AND U7988 ( .A(round_reg[1239]), .B(init), .Z(\round_in[0][1239] ) );
  NAND U7989 ( .A(init), .B(round_reg[123]), .Z(n2870) );
  NANDN U7990 ( .A(init), .B(in[123]), .Z(n2869) );
  NAND U7991 ( .A(n2870), .B(n2869), .Z(\round_in[0][123] ) );
  AND U7992 ( .A(round_reg[1240]), .B(init), .Z(\round_in[0][1240] ) );
  AND U7993 ( .A(round_reg[1241]), .B(init), .Z(\round_in[0][1241] ) );
  AND U7994 ( .A(round_reg[1242]), .B(init), .Z(\round_in[0][1242] ) );
  AND U7995 ( .A(round_reg[1243]), .B(init), .Z(\round_in[0][1243] ) );
  AND U7996 ( .A(round_reg[1244]), .B(init), .Z(\round_in[0][1244] ) );
  AND U7997 ( .A(round_reg[1245]), .B(init), .Z(\round_in[0][1245] ) );
  AND U7998 ( .A(round_reg[1246]), .B(init), .Z(\round_in[0][1246] ) );
  AND U7999 ( .A(round_reg[1247]), .B(init), .Z(\round_in[0][1247] ) );
  AND U8000 ( .A(round_reg[1248]), .B(init), .Z(\round_in[0][1248] ) );
  AND U8001 ( .A(round_reg[1249]), .B(init), .Z(\round_in[0][1249] ) );
  NAND U8002 ( .A(init), .B(round_reg[124]), .Z(n2872) );
  NANDN U8003 ( .A(init), .B(in[124]), .Z(n2871) );
  NAND U8004 ( .A(n2872), .B(n2871), .Z(\round_in[0][124] ) );
  AND U8005 ( .A(round_reg[1250]), .B(init), .Z(\round_in[0][1250] ) );
  AND U8006 ( .A(round_reg[1251]), .B(init), .Z(\round_in[0][1251] ) );
  AND U8007 ( .A(round_reg[1252]), .B(init), .Z(\round_in[0][1252] ) );
  AND U8008 ( .A(round_reg[1253]), .B(init), .Z(\round_in[0][1253] ) );
  AND U8009 ( .A(round_reg[1254]), .B(init), .Z(\round_in[0][1254] ) );
  AND U8010 ( .A(round_reg[1255]), .B(init), .Z(\round_in[0][1255] ) );
  AND U8011 ( .A(round_reg[1256]), .B(init), .Z(\round_in[0][1256] ) );
  AND U8012 ( .A(round_reg[1257]), .B(init), .Z(\round_in[0][1257] ) );
  AND U8013 ( .A(round_reg[1258]), .B(init), .Z(\round_in[0][1258] ) );
  AND U8014 ( .A(round_reg[1259]), .B(init), .Z(\round_in[0][1259] ) );
  NAND U8015 ( .A(init), .B(round_reg[125]), .Z(n2874) );
  NANDN U8016 ( .A(init), .B(in[125]), .Z(n2873) );
  NAND U8017 ( .A(n2874), .B(n2873), .Z(\round_in[0][125] ) );
  AND U8018 ( .A(round_reg[1260]), .B(init), .Z(\round_in[0][1260] ) );
  AND U8019 ( .A(round_reg[1261]), .B(init), .Z(\round_in[0][1261] ) );
  AND U8020 ( .A(round_reg[1262]), .B(init), .Z(\round_in[0][1262] ) );
  AND U8021 ( .A(round_reg[1263]), .B(init), .Z(\round_in[0][1263] ) );
  AND U8022 ( .A(round_reg[1264]), .B(init), .Z(\round_in[0][1264] ) );
  AND U8023 ( .A(round_reg[1265]), .B(init), .Z(\round_in[0][1265] ) );
  AND U8024 ( .A(round_reg[1266]), .B(init), .Z(\round_in[0][1266] ) );
  AND U8025 ( .A(round_reg[1267]), .B(init), .Z(\round_in[0][1267] ) );
  AND U8026 ( .A(round_reg[1268]), .B(init), .Z(\round_in[0][1268] ) );
  AND U8027 ( .A(round_reg[1269]), .B(init), .Z(\round_in[0][1269] ) );
  NAND U8028 ( .A(init), .B(round_reg[126]), .Z(n2876) );
  NANDN U8029 ( .A(init), .B(in[126]), .Z(n2875) );
  NAND U8030 ( .A(n2876), .B(n2875), .Z(\round_in[0][126] ) );
  AND U8031 ( .A(round_reg[1270]), .B(init), .Z(\round_in[0][1270] ) );
  AND U8032 ( .A(round_reg[1271]), .B(init), .Z(\round_in[0][1271] ) );
  AND U8033 ( .A(round_reg[1272]), .B(init), .Z(\round_in[0][1272] ) );
  AND U8034 ( .A(round_reg[1273]), .B(init), .Z(\round_in[0][1273] ) );
  AND U8035 ( .A(round_reg[1274]), .B(init), .Z(\round_in[0][1274] ) );
  AND U8036 ( .A(round_reg[1275]), .B(init), .Z(\round_in[0][1275] ) );
  AND U8037 ( .A(round_reg[1276]), .B(init), .Z(\round_in[0][1276] ) );
  AND U8038 ( .A(round_reg[1277]), .B(init), .Z(\round_in[0][1277] ) );
  AND U8039 ( .A(round_reg[1278]), .B(init), .Z(\round_in[0][1278] ) );
  AND U8040 ( .A(round_reg[1279]), .B(init), .Z(\round_in[0][1279] ) );
  NAND U8041 ( .A(init), .B(round_reg[127]), .Z(n2878) );
  NANDN U8042 ( .A(init), .B(in[127]), .Z(n2877) );
  NAND U8043 ( .A(n2878), .B(n2877), .Z(\round_in[0][127] ) );
  AND U8044 ( .A(round_reg[1280]), .B(init), .Z(\round_in[0][1280] ) );
  AND U8045 ( .A(round_reg[1281]), .B(init), .Z(\round_in[0][1281] ) );
  AND U8046 ( .A(round_reg[1282]), .B(init), .Z(\round_in[0][1282] ) );
  AND U8047 ( .A(round_reg[1283]), .B(init), .Z(\round_in[0][1283] ) );
  AND U8048 ( .A(round_reg[1284]), .B(init), .Z(\round_in[0][1284] ) );
  AND U8049 ( .A(round_reg[1285]), .B(init), .Z(\round_in[0][1285] ) );
  AND U8050 ( .A(round_reg[1286]), .B(init), .Z(\round_in[0][1286] ) );
  AND U8051 ( .A(round_reg[1287]), .B(init), .Z(\round_in[0][1287] ) );
  AND U8052 ( .A(round_reg[1288]), .B(init), .Z(\round_in[0][1288] ) );
  AND U8053 ( .A(round_reg[1289]), .B(init), .Z(\round_in[0][1289] ) );
  NAND U8054 ( .A(init), .B(round_reg[128]), .Z(n2880) );
  NANDN U8055 ( .A(init), .B(in[128]), .Z(n2879) );
  NAND U8056 ( .A(n2880), .B(n2879), .Z(\round_in[0][128] ) );
  AND U8057 ( .A(round_reg[1290]), .B(init), .Z(\round_in[0][1290] ) );
  AND U8058 ( .A(round_reg[1291]), .B(init), .Z(\round_in[0][1291] ) );
  AND U8059 ( .A(round_reg[1292]), .B(init), .Z(\round_in[0][1292] ) );
  AND U8060 ( .A(round_reg[1293]), .B(init), .Z(\round_in[0][1293] ) );
  AND U8061 ( .A(round_reg[1294]), .B(init), .Z(\round_in[0][1294] ) );
  AND U8062 ( .A(round_reg[1295]), .B(init), .Z(\round_in[0][1295] ) );
  AND U8063 ( .A(round_reg[1296]), .B(init), .Z(\round_in[0][1296] ) );
  AND U8064 ( .A(round_reg[1297]), .B(init), .Z(\round_in[0][1297] ) );
  AND U8065 ( .A(round_reg[1298]), .B(init), .Z(\round_in[0][1298] ) );
  AND U8066 ( .A(round_reg[1299]), .B(init), .Z(\round_in[0][1299] ) );
  NAND U8067 ( .A(init), .B(round_reg[129]), .Z(n2882) );
  NANDN U8068 ( .A(init), .B(in[129]), .Z(n2881) );
  NAND U8069 ( .A(n2882), .B(n2881), .Z(\round_in[0][129] ) );
  NAND U8070 ( .A(init), .B(round_reg[12]), .Z(n2884) );
  NANDN U8071 ( .A(init), .B(in[12]), .Z(n2883) );
  NAND U8072 ( .A(n2884), .B(n2883), .Z(\round_in[0][12] ) );
  AND U8073 ( .A(round_reg[1300]), .B(init), .Z(\round_in[0][1300] ) );
  AND U8074 ( .A(round_reg[1301]), .B(init), .Z(\round_in[0][1301] ) );
  AND U8075 ( .A(round_reg[1302]), .B(init), .Z(\round_in[0][1302] ) );
  AND U8076 ( .A(round_reg[1303]), .B(init), .Z(\round_in[0][1303] ) );
  AND U8077 ( .A(round_reg[1304]), .B(init), .Z(\round_in[0][1304] ) );
  AND U8078 ( .A(round_reg[1305]), .B(init), .Z(\round_in[0][1305] ) );
  AND U8079 ( .A(round_reg[1306]), .B(init), .Z(\round_in[0][1306] ) );
  AND U8080 ( .A(round_reg[1307]), .B(init), .Z(\round_in[0][1307] ) );
  AND U8081 ( .A(round_reg[1308]), .B(init), .Z(\round_in[0][1308] ) );
  AND U8082 ( .A(round_reg[1309]), .B(init), .Z(\round_in[0][1309] ) );
  NAND U8083 ( .A(init), .B(round_reg[130]), .Z(n2886) );
  NANDN U8084 ( .A(init), .B(in[130]), .Z(n2885) );
  NAND U8085 ( .A(n2886), .B(n2885), .Z(\round_in[0][130] ) );
  AND U8086 ( .A(round_reg[1310]), .B(init), .Z(\round_in[0][1310] ) );
  AND U8087 ( .A(round_reg[1311]), .B(init), .Z(\round_in[0][1311] ) );
  AND U8088 ( .A(round_reg[1312]), .B(init), .Z(\round_in[0][1312] ) );
  AND U8089 ( .A(round_reg[1313]), .B(init), .Z(\round_in[0][1313] ) );
  AND U8090 ( .A(round_reg[1314]), .B(init), .Z(\round_in[0][1314] ) );
  AND U8091 ( .A(round_reg[1315]), .B(init), .Z(\round_in[0][1315] ) );
  AND U8092 ( .A(round_reg[1316]), .B(init), .Z(\round_in[0][1316] ) );
  AND U8093 ( .A(round_reg[1317]), .B(init), .Z(\round_in[0][1317] ) );
  AND U8094 ( .A(round_reg[1318]), .B(init), .Z(\round_in[0][1318] ) );
  AND U8095 ( .A(round_reg[1319]), .B(init), .Z(\round_in[0][1319] ) );
  NAND U8096 ( .A(init), .B(round_reg[131]), .Z(n2888) );
  NANDN U8097 ( .A(init), .B(in[131]), .Z(n2887) );
  NAND U8098 ( .A(n2888), .B(n2887), .Z(\round_in[0][131] ) );
  AND U8099 ( .A(round_reg[1320]), .B(init), .Z(\round_in[0][1320] ) );
  AND U8100 ( .A(round_reg[1321]), .B(init), .Z(\round_in[0][1321] ) );
  AND U8101 ( .A(round_reg[1322]), .B(init), .Z(\round_in[0][1322] ) );
  AND U8102 ( .A(round_reg[1323]), .B(init), .Z(\round_in[0][1323] ) );
  AND U8103 ( .A(round_reg[1324]), .B(init), .Z(\round_in[0][1324] ) );
  AND U8104 ( .A(round_reg[1325]), .B(init), .Z(\round_in[0][1325] ) );
  AND U8105 ( .A(round_reg[1326]), .B(init), .Z(\round_in[0][1326] ) );
  AND U8106 ( .A(round_reg[1327]), .B(init), .Z(\round_in[0][1327] ) );
  AND U8107 ( .A(round_reg[1328]), .B(init), .Z(\round_in[0][1328] ) );
  AND U8108 ( .A(round_reg[1329]), .B(init), .Z(\round_in[0][1329] ) );
  NAND U8109 ( .A(init), .B(round_reg[132]), .Z(n2890) );
  NANDN U8110 ( .A(init), .B(in[132]), .Z(n2889) );
  NAND U8111 ( .A(n2890), .B(n2889), .Z(\round_in[0][132] ) );
  AND U8112 ( .A(round_reg[1330]), .B(init), .Z(\round_in[0][1330] ) );
  AND U8113 ( .A(round_reg[1331]), .B(init), .Z(\round_in[0][1331] ) );
  AND U8114 ( .A(round_reg[1332]), .B(init), .Z(\round_in[0][1332] ) );
  AND U8115 ( .A(round_reg[1333]), .B(init), .Z(\round_in[0][1333] ) );
  AND U8116 ( .A(round_reg[1334]), .B(init), .Z(\round_in[0][1334] ) );
  AND U8117 ( .A(round_reg[1335]), .B(init), .Z(\round_in[0][1335] ) );
  AND U8118 ( .A(round_reg[1336]), .B(init), .Z(\round_in[0][1336] ) );
  AND U8119 ( .A(round_reg[1337]), .B(init), .Z(\round_in[0][1337] ) );
  AND U8120 ( .A(round_reg[1338]), .B(init), .Z(\round_in[0][1338] ) );
  AND U8121 ( .A(round_reg[1339]), .B(init), .Z(\round_in[0][1339] ) );
  NAND U8122 ( .A(init), .B(round_reg[133]), .Z(n2892) );
  NANDN U8123 ( .A(init), .B(in[133]), .Z(n2891) );
  NAND U8124 ( .A(n2892), .B(n2891), .Z(\round_in[0][133] ) );
  AND U8125 ( .A(round_reg[1340]), .B(init), .Z(\round_in[0][1340] ) );
  AND U8126 ( .A(round_reg[1341]), .B(init), .Z(\round_in[0][1341] ) );
  AND U8127 ( .A(round_reg[1342]), .B(init), .Z(\round_in[0][1342] ) );
  AND U8128 ( .A(round_reg[1343]), .B(init), .Z(\round_in[0][1343] ) );
  AND U8129 ( .A(round_reg[1344]), .B(init), .Z(\round_in[0][1344] ) );
  AND U8130 ( .A(round_reg[1345]), .B(init), .Z(\round_in[0][1345] ) );
  AND U8131 ( .A(round_reg[1346]), .B(init), .Z(\round_in[0][1346] ) );
  AND U8132 ( .A(round_reg[1347]), .B(init), .Z(\round_in[0][1347] ) );
  AND U8133 ( .A(round_reg[1348]), .B(init), .Z(\round_in[0][1348] ) );
  AND U8134 ( .A(round_reg[1349]), .B(init), .Z(\round_in[0][1349] ) );
  NAND U8135 ( .A(init), .B(round_reg[134]), .Z(n2894) );
  NANDN U8136 ( .A(init), .B(in[134]), .Z(n2893) );
  NAND U8137 ( .A(n2894), .B(n2893), .Z(\round_in[0][134] ) );
  AND U8138 ( .A(round_reg[1350]), .B(init), .Z(\round_in[0][1350] ) );
  AND U8139 ( .A(round_reg[1351]), .B(init), .Z(\round_in[0][1351] ) );
  AND U8140 ( .A(round_reg[1352]), .B(init), .Z(\round_in[0][1352] ) );
  AND U8141 ( .A(round_reg[1353]), .B(init), .Z(\round_in[0][1353] ) );
  AND U8142 ( .A(round_reg[1354]), .B(init), .Z(\round_in[0][1354] ) );
  AND U8143 ( .A(round_reg[1355]), .B(init), .Z(\round_in[0][1355] ) );
  AND U8144 ( .A(round_reg[1356]), .B(init), .Z(\round_in[0][1356] ) );
  AND U8145 ( .A(round_reg[1357]), .B(init), .Z(\round_in[0][1357] ) );
  AND U8146 ( .A(round_reg[1358]), .B(init), .Z(\round_in[0][1358] ) );
  AND U8147 ( .A(round_reg[1359]), .B(init), .Z(\round_in[0][1359] ) );
  NAND U8148 ( .A(init), .B(round_reg[135]), .Z(n2896) );
  NANDN U8149 ( .A(init), .B(in[135]), .Z(n2895) );
  NAND U8150 ( .A(n2896), .B(n2895), .Z(\round_in[0][135] ) );
  AND U8151 ( .A(round_reg[1360]), .B(init), .Z(\round_in[0][1360] ) );
  AND U8152 ( .A(round_reg[1361]), .B(init), .Z(\round_in[0][1361] ) );
  AND U8153 ( .A(round_reg[1362]), .B(init), .Z(\round_in[0][1362] ) );
  AND U8154 ( .A(round_reg[1363]), .B(init), .Z(\round_in[0][1363] ) );
  AND U8155 ( .A(round_reg[1364]), .B(init), .Z(\round_in[0][1364] ) );
  AND U8156 ( .A(round_reg[1365]), .B(init), .Z(\round_in[0][1365] ) );
  AND U8157 ( .A(round_reg[1366]), .B(init), .Z(\round_in[0][1366] ) );
  AND U8158 ( .A(round_reg[1367]), .B(init), .Z(\round_in[0][1367] ) );
  AND U8159 ( .A(round_reg[1368]), .B(init), .Z(\round_in[0][1368] ) );
  AND U8160 ( .A(round_reg[1369]), .B(init), .Z(\round_in[0][1369] ) );
  NAND U8161 ( .A(init), .B(round_reg[136]), .Z(n2898) );
  NANDN U8162 ( .A(init), .B(in[136]), .Z(n2897) );
  NAND U8163 ( .A(n2898), .B(n2897), .Z(\round_in[0][136] ) );
  AND U8164 ( .A(round_reg[1370]), .B(init), .Z(\round_in[0][1370] ) );
  AND U8165 ( .A(round_reg[1371]), .B(init), .Z(\round_in[0][1371] ) );
  AND U8166 ( .A(round_reg[1372]), .B(init), .Z(\round_in[0][1372] ) );
  AND U8167 ( .A(round_reg[1373]), .B(init), .Z(\round_in[0][1373] ) );
  AND U8168 ( .A(round_reg[1374]), .B(init), .Z(\round_in[0][1374] ) );
  AND U8169 ( .A(round_reg[1375]), .B(init), .Z(\round_in[0][1375] ) );
  AND U8170 ( .A(round_reg[1376]), .B(init), .Z(\round_in[0][1376] ) );
  AND U8171 ( .A(round_reg[1377]), .B(init), .Z(\round_in[0][1377] ) );
  AND U8172 ( .A(round_reg[1378]), .B(init), .Z(\round_in[0][1378] ) );
  AND U8173 ( .A(round_reg[1379]), .B(init), .Z(\round_in[0][1379] ) );
  NAND U8174 ( .A(init), .B(round_reg[137]), .Z(n2900) );
  NANDN U8175 ( .A(init), .B(in[137]), .Z(n2899) );
  NAND U8176 ( .A(n2900), .B(n2899), .Z(\round_in[0][137] ) );
  AND U8177 ( .A(round_reg[1380]), .B(init), .Z(\round_in[0][1380] ) );
  AND U8178 ( .A(round_reg[1381]), .B(init), .Z(\round_in[0][1381] ) );
  AND U8179 ( .A(round_reg[1382]), .B(init), .Z(\round_in[0][1382] ) );
  AND U8180 ( .A(round_reg[1383]), .B(init), .Z(\round_in[0][1383] ) );
  AND U8181 ( .A(round_reg[1384]), .B(init), .Z(\round_in[0][1384] ) );
  AND U8182 ( .A(round_reg[1385]), .B(init), .Z(\round_in[0][1385] ) );
  AND U8183 ( .A(round_reg[1386]), .B(init), .Z(\round_in[0][1386] ) );
  AND U8184 ( .A(round_reg[1387]), .B(init), .Z(\round_in[0][1387] ) );
  AND U8185 ( .A(round_reg[1388]), .B(init), .Z(\round_in[0][1388] ) );
  AND U8186 ( .A(round_reg[1389]), .B(init), .Z(\round_in[0][1389] ) );
  NAND U8187 ( .A(init), .B(round_reg[138]), .Z(n2902) );
  NANDN U8188 ( .A(init), .B(in[138]), .Z(n2901) );
  NAND U8189 ( .A(n2902), .B(n2901), .Z(\round_in[0][138] ) );
  AND U8190 ( .A(round_reg[1390]), .B(init), .Z(\round_in[0][1390] ) );
  AND U8191 ( .A(round_reg[1391]), .B(init), .Z(\round_in[0][1391] ) );
  AND U8192 ( .A(round_reg[1392]), .B(init), .Z(\round_in[0][1392] ) );
  AND U8193 ( .A(round_reg[1393]), .B(init), .Z(\round_in[0][1393] ) );
  AND U8194 ( .A(round_reg[1394]), .B(init), .Z(\round_in[0][1394] ) );
  AND U8195 ( .A(round_reg[1395]), .B(init), .Z(\round_in[0][1395] ) );
  AND U8196 ( .A(round_reg[1396]), .B(init), .Z(\round_in[0][1396] ) );
  AND U8197 ( .A(round_reg[1397]), .B(init), .Z(\round_in[0][1397] ) );
  AND U8198 ( .A(round_reg[1398]), .B(init), .Z(\round_in[0][1398] ) );
  AND U8199 ( .A(round_reg[1399]), .B(init), .Z(\round_in[0][1399] ) );
  NAND U8200 ( .A(init), .B(round_reg[139]), .Z(n2904) );
  NANDN U8201 ( .A(init), .B(in[139]), .Z(n2903) );
  NAND U8202 ( .A(n2904), .B(n2903), .Z(\round_in[0][139] ) );
  NAND U8203 ( .A(init), .B(round_reg[13]), .Z(n2906) );
  NANDN U8204 ( .A(init), .B(in[13]), .Z(n2905) );
  NAND U8205 ( .A(n2906), .B(n2905), .Z(\round_in[0][13] ) );
  AND U8206 ( .A(round_reg[1400]), .B(init), .Z(\round_in[0][1400] ) );
  AND U8207 ( .A(round_reg[1401]), .B(init), .Z(\round_in[0][1401] ) );
  AND U8208 ( .A(round_reg[1402]), .B(init), .Z(\round_in[0][1402] ) );
  AND U8209 ( .A(round_reg[1403]), .B(init), .Z(\round_in[0][1403] ) );
  AND U8210 ( .A(round_reg[1404]), .B(init), .Z(\round_in[0][1404] ) );
  AND U8211 ( .A(round_reg[1405]), .B(init), .Z(\round_in[0][1405] ) );
  AND U8212 ( .A(round_reg[1406]), .B(init), .Z(\round_in[0][1406] ) );
  AND U8213 ( .A(round_reg[1407]), .B(init), .Z(\round_in[0][1407] ) );
  AND U8214 ( .A(round_reg[1408]), .B(init), .Z(\round_in[0][1408] ) );
  AND U8215 ( .A(round_reg[1409]), .B(init), .Z(\round_in[0][1409] ) );
  NAND U8216 ( .A(init), .B(round_reg[140]), .Z(n2908) );
  NANDN U8217 ( .A(init), .B(in[140]), .Z(n2907) );
  NAND U8218 ( .A(n2908), .B(n2907), .Z(\round_in[0][140] ) );
  AND U8219 ( .A(round_reg[1410]), .B(init), .Z(\round_in[0][1410] ) );
  AND U8220 ( .A(round_reg[1411]), .B(init), .Z(\round_in[0][1411] ) );
  AND U8221 ( .A(round_reg[1412]), .B(init), .Z(\round_in[0][1412] ) );
  AND U8222 ( .A(round_reg[1413]), .B(init), .Z(\round_in[0][1413] ) );
  AND U8223 ( .A(round_reg[1414]), .B(init), .Z(\round_in[0][1414] ) );
  AND U8224 ( .A(round_reg[1415]), .B(init), .Z(\round_in[0][1415] ) );
  AND U8225 ( .A(round_reg[1416]), .B(init), .Z(\round_in[0][1416] ) );
  AND U8226 ( .A(round_reg[1417]), .B(init), .Z(\round_in[0][1417] ) );
  AND U8227 ( .A(round_reg[1418]), .B(init), .Z(\round_in[0][1418] ) );
  AND U8228 ( .A(round_reg[1419]), .B(init), .Z(\round_in[0][1419] ) );
  NAND U8229 ( .A(init), .B(round_reg[141]), .Z(n2910) );
  NANDN U8230 ( .A(init), .B(in[141]), .Z(n2909) );
  NAND U8231 ( .A(n2910), .B(n2909), .Z(\round_in[0][141] ) );
  AND U8232 ( .A(round_reg[1420]), .B(init), .Z(\round_in[0][1420] ) );
  AND U8233 ( .A(round_reg[1421]), .B(init), .Z(\round_in[0][1421] ) );
  AND U8234 ( .A(round_reg[1422]), .B(init), .Z(\round_in[0][1422] ) );
  AND U8235 ( .A(round_reg[1423]), .B(init), .Z(\round_in[0][1423] ) );
  AND U8236 ( .A(round_reg[1424]), .B(init), .Z(\round_in[0][1424] ) );
  AND U8237 ( .A(round_reg[1425]), .B(init), .Z(\round_in[0][1425] ) );
  AND U8238 ( .A(round_reg[1426]), .B(init), .Z(\round_in[0][1426] ) );
  AND U8239 ( .A(round_reg[1427]), .B(init), .Z(\round_in[0][1427] ) );
  AND U8240 ( .A(round_reg[1428]), .B(init), .Z(\round_in[0][1428] ) );
  AND U8241 ( .A(round_reg[1429]), .B(init), .Z(\round_in[0][1429] ) );
  NAND U8242 ( .A(init), .B(round_reg[142]), .Z(n2912) );
  NANDN U8243 ( .A(init), .B(in[142]), .Z(n2911) );
  NAND U8244 ( .A(n2912), .B(n2911), .Z(\round_in[0][142] ) );
  AND U8245 ( .A(round_reg[1430]), .B(init), .Z(\round_in[0][1430] ) );
  AND U8246 ( .A(round_reg[1431]), .B(init), .Z(\round_in[0][1431] ) );
  AND U8247 ( .A(round_reg[1432]), .B(init), .Z(\round_in[0][1432] ) );
  AND U8248 ( .A(round_reg[1433]), .B(init), .Z(\round_in[0][1433] ) );
  AND U8249 ( .A(round_reg[1434]), .B(init), .Z(\round_in[0][1434] ) );
  AND U8250 ( .A(round_reg[1435]), .B(init), .Z(\round_in[0][1435] ) );
  AND U8251 ( .A(round_reg[1436]), .B(init), .Z(\round_in[0][1436] ) );
  AND U8252 ( .A(round_reg[1437]), .B(init), .Z(\round_in[0][1437] ) );
  AND U8253 ( .A(round_reg[1438]), .B(init), .Z(\round_in[0][1438] ) );
  AND U8254 ( .A(round_reg[1439]), .B(init), .Z(\round_in[0][1439] ) );
  NAND U8255 ( .A(init), .B(round_reg[143]), .Z(n2914) );
  NANDN U8256 ( .A(init), .B(in[143]), .Z(n2913) );
  NAND U8257 ( .A(n2914), .B(n2913), .Z(\round_in[0][143] ) );
  AND U8258 ( .A(round_reg[1440]), .B(init), .Z(\round_in[0][1440] ) );
  AND U8259 ( .A(round_reg[1441]), .B(init), .Z(\round_in[0][1441] ) );
  AND U8260 ( .A(round_reg[1442]), .B(init), .Z(\round_in[0][1442] ) );
  AND U8261 ( .A(round_reg[1443]), .B(init), .Z(\round_in[0][1443] ) );
  AND U8262 ( .A(round_reg[1444]), .B(init), .Z(\round_in[0][1444] ) );
  AND U8263 ( .A(round_reg[1445]), .B(init), .Z(\round_in[0][1445] ) );
  AND U8264 ( .A(round_reg[1446]), .B(init), .Z(\round_in[0][1446] ) );
  AND U8265 ( .A(round_reg[1447]), .B(init), .Z(\round_in[0][1447] ) );
  AND U8266 ( .A(round_reg[1448]), .B(init), .Z(\round_in[0][1448] ) );
  AND U8267 ( .A(round_reg[1449]), .B(init), .Z(\round_in[0][1449] ) );
  NAND U8268 ( .A(init), .B(round_reg[144]), .Z(n2916) );
  NANDN U8269 ( .A(init), .B(in[144]), .Z(n2915) );
  NAND U8270 ( .A(n2916), .B(n2915), .Z(\round_in[0][144] ) );
  AND U8271 ( .A(round_reg[1450]), .B(init), .Z(\round_in[0][1450] ) );
  AND U8272 ( .A(round_reg[1451]), .B(init), .Z(\round_in[0][1451] ) );
  AND U8273 ( .A(round_reg[1452]), .B(init), .Z(\round_in[0][1452] ) );
  AND U8274 ( .A(round_reg[1453]), .B(init), .Z(\round_in[0][1453] ) );
  AND U8275 ( .A(round_reg[1454]), .B(init), .Z(\round_in[0][1454] ) );
  AND U8276 ( .A(round_reg[1455]), .B(init), .Z(\round_in[0][1455] ) );
  AND U8277 ( .A(round_reg[1456]), .B(init), .Z(\round_in[0][1456] ) );
  AND U8278 ( .A(round_reg[1457]), .B(init), .Z(\round_in[0][1457] ) );
  AND U8279 ( .A(round_reg[1458]), .B(init), .Z(\round_in[0][1458] ) );
  AND U8280 ( .A(round_reg[1459]), .B(init), .Z(\round_in[0][1459] ) );
  NAND U8281 ( .A(init), .B(round_reg[145]), .Z(n2918) );
  NANDN U8282 ( .A(init), .B(in[145]), .Z(n2917) );
  NAND U8283 ( .A(n2918), .B(n2917), .Z(\round_in[0][145] ) );
  AND U8284 ( .A(round_reg[1460]), .B(init), .Z(\round_in[0][1460] ) );
  AND U8285 ( .A(round_reg[1461]), .B(init), .Z(\round_in[0][1461] ) );
  AND U8286 ( .A(round_reg[1462]), .B(init), .Z(\round_in[0][1462] ) );
  AND U8287 ( .A(round_reg[1463]), .B(init), .Z(\round_in[0][1463] ) );
  AND U8288 ( .A(round_reg[1464]), .B(init), .Z(\round_in[0][1464] ) );
  AND U8289 ( .A(round_reg[1465]), .B(init), .Z(\round_in[0][1465] ) );
  AND U8290 ( .A(round_reg[1466]), .B(init), .Z(\round_in[0][1466] ) );
  AND U8291 ( .A(round_reg[1467]), .B(init), .Z(\round_in[0][1467] ) );
  AND U8292 ( .A(round_reg[1468]), .B(init), .Z(\round_in[0][1468] ) );
  AND U8293 ( .A(round_reg[1469]), .B(init), .Z(\round_in[0][1469] ) );
  NAND U8294 ( .A(init), .B(round_reg[146]), .Z(n2920) );
  NANDN U8295 ( .A(init), .B(in[146]), .Z(n2919) );
  NAND U8296 ( .A(n2920), .B(n2919), .Z(\round_in[0][146] ) );
  AND U8297 ( .A(round_reg[1470]), .B(init), .Z(\round_in[0][1470] ) );
  AND U8298 ( .A(round_reg[1471]), .B(init), .Z(\round_in[0][1471] ) );
  AND U8299 ( .A(round_reg[1472]), .B(init), .Z(\round_in[0][1472] ) );
  AND U8300 ( .A(round_reg[1473]), .B(init), .Z(\round_in[0][1473] ) );
  AND U8301 ( .A(round_reg[1474]), .B(init), .Z(\round_in[0][1474] ) );
  AND U8302 ( .A(round_reg[1475]), .B(init), .Z(\round_in[0][1475] ) );
  AND U8303 ( .A(round_reg[1476]), .B(init), .Z(\round_in[0][1476] ) );
  AND U8304 ( .A(round_reg[1477]), .B(init), .Z(\round_in[0][1477] ) );
  AND U8305 ( .A(round_reg[1478]), .B(init), .Z(\round_in[0][1478] ) );
  AND U8306 ( .A(round_reg[1479]), .B(init), .Z(\round_in[0][1479] ) );
  NAND U8307 ( .A(init), .B(round_reg[147]), .Z(n2922) );
  NANDN U8308 ( .A(init), .B(in[147]), .Z(n2921) );
  NAND U8309 ( .A(n2922), .B(n2921), .Z(\round_in[0][147] ) );
  AND U8310 ( .A(round_reg[1480]), .B(init), .Z(\round_in[0][1480] ) );
  AND U8311 ( .A(round_reg[1481]), .B(init), .Z(\round_in[0][1481] ) );
  AND U8312 ( .A(round_reg[1482]), .B(init), .Z(\round_in[0][1482] ) );
  AND U8313 ( .A(round_reg[1483]), .B(init), .Z(\round_in[0][1483] ) );
  AND U8314 ( .A(round_reg[1484]), .B(init), .Z(\round_in[0][1484] ) );
  AND U8315 ( .A(round_reg[1485]), .B(init), .Z(\round_in[0][1485] ) );
  AND U8316 ( .A(round_reg[1486]), .B(init), .Z(\round_in[0][1486] ) );
  AND U8317 ( .A(round_reg[1487]), .B(init), .Z(\round_in[0][1487] ) );
  AND U8318 ( .A(round_reg[1488]), .B(init), .Z(\round_in[0][1488] ) );
  AND U8319 ( .A(round_reg[1489]), .B(init), .Z(\round_in[0][1489] ) );
  NAND U8320 ( .A(init), .B(round_reg[148]), .Z(n2924) );
  NANDN U8321 ( .A(init), .B(in[148]), .Z(n2923) );
  NAND U8322 ( .A(n2924), .B(n2923), .Z(\round_in[0][148] ) );
  AND U8323 ( .A(round_reg[1490]), .B(init), .Z(\round_in[0][1490] ) );
  AND U8324 ( .A(round_reg[1491]), .B(init), .Z(\round_in[0][1491] ) );
  AND U8325 ( .A(round_reg[1492]), .B(init), .Z(\round_in[0][1492] ) );
  AND U8326 ( .A(round_reg[1493]), .B(init), .Z(\round_in[0][1493] ) );
  AND U8327 ( .A(round_reg[1494]), .B(init), .Z(\round_in[0][1494] ) );
  AND U8328 ( .A(round_reg[1495]), .B(init), .Z(\round_in[0][1495] ) );
  AND U8329 ( .A(round_reg[1496]), .B(init), .Z(\round_in[0][1496] ) );
  AND U8330 ( .A(round_reg[1497]), .B(init), .Z(\round_in[0][1497] ) );
  AND U8331 ( .A(round_reg[1498]), .B(init), .Z(\round_in[0][1498] ) );
  AND U8332 ( .A(round_reg[1499]), .B(init), .Z(\round_in[0][1499] ) );
  NAND U8333 ( .A(init), .B(round_reg[149]), .Z(n2926) );
  NANDN U8334 ( .A(init), .B(in[149]), .Z(n2925) );
  NAND U8335 ( .A(n2926), .B(n2925), .Z(\round_in[0][149] ) );
  NAND U8336 ( .A(init), .B(round_reg[14]), .Z(n2928) );
  NANDN U8337 ( .A(init), .B(in[14]), .Z(n2927) );
  NAND U8338 ( .A(n2928), .B(n2927), .Z(\round_in[0][14] ) );
  AND U8339 ( .A(round_reg[1500]), .B(init), .Z(\round_in[0][1500] ) );
  AND U8340 ( .A(round_reg[1501]), .B(init), .Z(\round_in[0][1501] ) );
  AND U8341 ( .A(round_reg[1502]), .B(init), .Z(\round_in[0][1502] ) );
  AND U8342 ( .A(round_reg[1503]), .B(init), .Z(\round_in[0][1503] ) );
  AND U8343 ( .A(round_reg[1504]), .B(init), .Z(\round_in[0][1504] ) );
  AND U8344 ( .A(round_reg[1505]), .B(init), .Z(\round_in[0][1505] ) );
  AND U8345 ( .A(round_reg[1506]), .B(init), .Z(\round_in[0][1506] ) );
  AND U8346 ( .A(round_reg[1507]), .B(init), .Z(\round_in[0][1507] ) );
  AND U8347 ( .A(round_reg[1508]), .B(init), .Z(\round_in[0][1508] ) );
  AND U8348 ( .A(round_reg[1509]), .B(init), .Z(\round_in[0][1509] ) );
  NAND U8349 ( .A(init), .B(round_reg[150]), .Z(n2930) );
  NANDN U8350 ( .A(init), .B(in[150]), .Z(n2929) );
  NAND U8351 ( .A(n2930), .B(n2929), .Z(\round_in[0][150] ) );
  AND U8352 ( .A(round_reg[1510]), .B(init), .Z(\round_in[0][1510] ) );
  AND U8353 ( .A(round_reg[1511]), .B(init), .Z(\round_in[0][1511] ) );
  AND U8354 ( .A(round_reg[1512]), .B(init), .Z(\round_in[0][1512] ) );
  AND U8355 ( .A(round_reg[1513]), .B(init), .Z(\round_in[0][1513] ) );
  AND U8356 ( .A(round_reg[1514]), .B(init), .Z(\round_in[0][1514] ) );
  AND U8357 ( .A(round_reg[1515]), .B(init), .Z(\round_in[0][1515] ) );
  AND U8358 ( .A(round_reg[1516]), .B(init), .Z(\round_in[0][1516] ) );
  AND U8359 ( .A(round_reg[1517]), .B(init), .Z(\round_in[0][1517] ) );
  AND U8360 ( .A(round_reg[1518]), .B(init), .Z(\round_in[0][1518] ) );
  AND U8361 ( .A(round_reg[1519]), .B(init), .Z(\round_in[0][1519] ) );
  NAND U8362 ( .A(init), .B(round_reg[151]), .Z(n2932) );
  NANDN U8363 ( .A(init), .B(in[151]), .Z(n2931) );
  NAND U8364 ( .A(n2932), .B(n2931), .Z(\round_in[0][151] ) );
  AND U8365 ( .A(round_reg[1520]), .B(init), .Z(\round_in[0][1520] ) );
  AND U8366 ( .A(round_reg[1521]), .B(init), .Z(\round_in[0][1521] ) );
  AND U8367 ( .A(round_reg[1522]), .B(init), .Z(\round_in[0][1522] ) );
  AND U8368 ( .A(round_reg[1523]), .B(init), .Z(\round_in[0][1523] ) );
  AND U8369 ( .A(round_reg[1524]), .B(init), .Z(\round_in[0][1524] ) );
  AND U8370 ( .A(round_reg[1525]), .B(init), .Z(\round_in[0][1525] ) );
  AND U8371 ( .A(round_reg[1526]), .B(init), .Z(\round_in[0][1526] ) );
  AND U8372 ( .A(round_reg[1527]), .B(init), .Z(\round_in[0][1527] ) );
  AND U8373 ( .A(round_reg[1528]), .B(init), .Z(\round_in[0][1528] ) );
  AND U8374 ( .A(round_reg[1529]), .B(init), .Z(\round_in[0][1529] ) );
  NAND U8375 ( .A(init), .B(round_reg[152]), .Z(n2934) );
  NANDN U8376 ( .A(init), .B(in[152]), .Z(n2933) );
  NAND U8377 ( .A(n2934), .B(n2933), .Z(\round_in[0][152] ) );
  AND U8378 ( .A(round_reg[1530]), .B(init), .Z(\round_in[0][1530] ) );
  AND U8379 ( .A(round_reg[1531]), .B(init), .Z(\round_in[0][1531] ) );
  AND U8380 ( .A(round_reg[1532]), .B(init), .Z(\round_in[0][1532] ) );
  AND U8381 ( .A(round_reg[1533]), .B(init), .Z(\round_in[0][1533] ) );
  AND U8382 ( .A(round_reg[1534]), .B(init), .Z(\round_in[0][1534] ) );
  AND U8383 ( .A(round_reg[1535]), .B(init), .Z(\round_in[0][1535] ) );
  AND U8384 ( .A(round_reg[1536]), .B(init), .Z(\round_in[0][1536] ) );
  AND U8385 ( .A(round_reg[1537]), .B(init), .Z(\round_in[0][1537] ) );
  AND U8386 ( .A(round_reg[1538]), .B(init), .Z(\round_in[0][1538] ) );
  AND U8387 ( .A(round_reg[1539]), .B(init), .Z(\round_in[0][1539] ) );
  NAND U8388 ( .A(init), .B(round_reg[153]), .Z(n2936) );
  NANDN U8389 ( .A(init), .B(in[153]), .Z(n2935) );
  NAND U8390 ( .A(n2936), .B(n2935), .Z(\round_in[0][153] ) );
  AND U8391 ( .A(round_reg[1540]), .B(init), .Z(\round_in[0][1540] ) );
  AND U8392 ( .A(round_reg[1541]), .B(init), .Z(\round_in[0][1541] ) );
  AND U8393 ( .A(round_reg[1542]), .B(init), .Z(\round_in[0][1542] ) );
  AND U8394 ( .A(round_reg[1543]), .B(init), .Z(\round_in[0][1543] ) );
  AND U8395 ( .A(round_reg[1544]), .B(init), .Z(\round_in[0][1544] ) );
  AND U8396 ( .A(round_reg[1545]), .B(init), .Z(\round_in[0][1545] ) );
  AND U8397 ( .A(round_reg[1546]), .B(init), .Z(\round_in[0][1546] ) );
  AND U8398 ( .A(round_reg[1547]), .B(init), .Z(\round_in[0][1547] ) );
  AND U8399 ( .A(round_reg[1548]), .B(init), .Z(\round_in[0][1548] ) );
  AND U8400 ( .A(round_reg[1549]), .B(init), .Z(\round_in[0][1549] ) );
  NAND U8401 ( .A(init), .B(round_reg[154]), .Z(n2938) );
  NANDN U8402 ( .A(init), .B(in[154]), .Z(n2937) );
  NAND U8403 ( .A(n2938), .B(n2937), .Z(\round_in[0][154] ) );
  AND U8404 ( .A(round_reg[1550]), .B(init), .Z(\round_in[0][1550] ) );
  AND U8405 ( .A(round_reg[1551]), .B(init), .Z(\round_in[0][1551] ) );
  AND U8406 ( .A(round_reg[1552]), .B(init), .Z(\round_in[0][1552] ) );
  AND U8407 ( .A(round_reg[1553]), .B(init), .Z(\round_in[0][1553] ) );
  AND U8408 ( .A(round_reg[1554]), .B(init), .Z(\round_in[0][1554] ) );
  AND U8409 ( .A(round_reg[1555]), .B(init), .Z(\round_in[0][1555] ) );
  AND U8410 ( .A(round_reg[1556]), .B(init), .Z(\round_in[0][1556] ) );
  AND U8411 ( .A(round_reg[1557]), .B(init), .Z(\round_in[0][1557] ) );
  AND U8412 ( .A(round_reg[1558]), .B(init), .Z(\round_in[0][1558] ) );
  AND U8413 ( .A(round_reg[1559]), .B(init), .Z(\round_in[0][1559] ) );
  NAND U8414 ( .A(init), .B(round_reg[155]), .Z(n2940) );
  NANDN U8415 ( .A(init), .B(in[155]), .Z(n2939) );
  NAND U8416 ( .A(n2940), .B(n2939), .Z(\round_in[0][155] ) );
  AND U8417 ( .A(round_reg[1560]), .B(init), .Z(\round_in[0][1560] ) );
  AND U8418 ( .A(round_reg[1561]), .B(init), .Z(\round_in[0][1561] ) );
  AND U8419 ( .A(round_reg[1562]), .B(init), .Z(\round_in[0][1562] ) );
  AND U8420 ( .A(round_reg[1563]), .B(init), .Z(\round_in[0][1563] ) );
  AND U8421 ( .A(round_reg[1564]), .B(init), .Z(\round_in[0][1564] ) );
  AND U8422 ( .A(round_reg[1565]), .B(init), .Z(\round_in[0][1565] ) );
  AND U8423 ( .A(round_reg[1566]), .B(init), .Z(\round_in[0][1566] ) );
  AND U8424 ( .A(round_reg[1567]), .B(init), .Z(\round_in[0][1567] ) );
  AND U8425 ( .A(round_reg[1568]), .B(init), .Z(\round_in[0][1568] ) );
  AND U8426 ( .A(round_reg[1569]), .B(init), .Z(\round_in[0][1569] ) );
  NAND U8427 ( .A(init), .B(round_reg[156]), .Z(n2942) );
  NANDN U8428 ( .A(init), .B(in[156]), .Z(n2941) );
  NAND U8429 ( .A(n2942), .B(n2941), .Z(\round_in[0][156] ) );
  AND U8430 ( .A(round_reg[1570]), .B(init), .Z(\round_in[0][1570] ) );
  AND U8431 ( .A(round_reg[1571]), .B(init), .Z(\round_in[0][1571] ) );
  AND U8432 ( .A(round_reg[1572]), .B(init), .Z(\round_in[0][1572] ) );
  AND U8433 ( .A(round_reg[1573]), .B(init), .Z(\round_in[0][1573] ) );
  AND U8434 ( .A(round_reg[1574]), .B(init), .Z(\round_in[0][1574] ) );
  AND U8435 ( .A(round_reg[1575]), .B(init), .Z(\round_in[0][1575] ) );
  AND U8436 ( .A(round_reg[1576]), .B(init), .Z(\round_in[0][1576] ) );
  AND U8437 ( .A(round_reg[1577]), .B(init), .Z(\round_in[0][1577] ) );
  AND U8438 ( .A(round_reg[1578]), .B(init), .Z(\round_in[0][1578] ) );
  AND U8439 ( .A(round_reg[1579]), .B(init), .Z(\round_in[0][1579] ) );
  NAND U8440 ( .A(init), .B(round_reg[157]), .Z(n2944) );
  NANDN U8441 ( .A(init), .B(in[157]), .Z(n2943) );
  NAND U8442 ( .A(n2944), .B(n2943), .Z(\round_in[0][157] ) );
  AND U8443 ( .A(round_reg[1580]), .B(init), .Z(\round_in[0][1580] ) );
  AND U8444 ( .A(round_reg[1581]), .B(init), .Z(\round_in[0][1581] ) );
  AND U8445 ( .A(round_reg[1582]), .B(init), .Z(\round_in[0][1582] ) );
  AND U8446 ( .A(round_reg[1583]), .B(init), .Z(\round_in[0][1583] ) );
  AND U8447 ( .A(round_reg[1584]), .B(init), .Z(\round_in[0][1584] ) );
  AND U8448 ( .A(round_reg[1585]), .B(init), .Z(\round_in[0][1585] ) );
  AND U8449 ( .A(round_reg[1586]), .B(init), .Z(\round_in[0][1586] ) );
  AND U8450 ( .A(round_reg[1587]), .B(init), .Z(\round_in[0][1587] ) );
  AND U8451 ( .A(round_reg[1588]), .B(init), .Z(\round_in[0][1588] ) );
  AND U8452 ( .A(round_reg[1589]), .B(init), .Z(\round_in[0][1589] ) );
  NAND U8453 ( .A(init), .B(round_reg[158]), .Z(n2946) );
  NANDN U8454 ( .A(init), .B(in[158]), .Z(n2945) );
  NAND U8455 ( .A(n2946), .B(n2945), .Z(\round_in[0][158] ) );
  AND U8456 ( .A(round_reg[1590]), .B(init), .Z(\round_in[0][1590] ) );
  AND U8457 ( .A(round_reg[1591]), .B(init), .Z(\round_in[0][1591] ) );
  AND U8458 ( .A(round_reg[1592]), .B(init), .Z(\round_in[0][1592] ) );
  AND U8459 ( .A(round_reg[1593]), .B(init), .Z(\round_in[0][1593] ) );
  AND U8460 ( .A(round_reg[1594]), .B(init), .Z(\round_in[0][1594] ) );
  AND U8461 ( .A(round_reg[1595]), .B(init), .Z(\round_in[0][1595] ) );
  AND U8462 ( .A(round_reg[1596]), .B(init), .Z(\round_in[0][1596] ) );
  AND U8463 ( .A(round_reg[1597]), .B(init), .Z(\round_in[0][1597] ) );
  AND U8464 ( .A(round_reg[1598]), .B(init), .Z(\round_in[0][1598] ) );
  AND U8465 ( .A(round_reg[1599]), .B(init), .Z(\round_in[0][1599] ) );
  NAND U8466 ( .A(init), .B(round_reg[159]), .Z(n2948) );
  NANDN U8467 ( .A(init), .B(in[159]), .Z(n2947) );
  NAND U8468 ( .A(n2948), .B(n2947), .Z(\round_in[0][159] ) );
  NAND U8469 ( .A(init), .B(round_reg[15]), .Z(n2950) );
  NANDN U8470 ( .A(init), .B(in[15]), .Z(n2949) );
  NAND U8471 ( .A(n2950), .B(n2949), .Z(\round_in[0][15] ) );
  NAND U8472 ( .A(init), .B(round_reg[160]), .Z(n2952) );
  NANDN U8473 ( .A(init), .B(in[160]), .Z(n2951) );
  NAND U8474 ( .A(n2952), .B(n2951), .Z(\round_in[0][160] ) );
  NAND U8475 ( .A(init), .B(round_reg[161]), .Z(n2954) );
  NANDN U8476 ( .A(init), .B(in[161]), .Z(n2953) );
  NAND U8477 ( .A(n2954), .B(n2953), .Z(\round_in[0][161] ) );
  NAND U8478 ( .A(init), .B(round_reg[162]), .Z(n2956) );
  NANDN U8479 ( .A(init), .B(in[162]), .Z(n2955) );
  NAND U8480 ( .A(n2956), .B(n2955), .Z(\round_in[0][162] ) );
  NAND U8481 ( .A(init), .B(round_reg[163]), .Z(n2958) );
  NANDN U8482 ( .A(init), .B(in[163]), .Z(n2957) );
  NAND U8483 ( .A(n2958), .B(n2957), .Z(\round_in[0][163] ) );
  NAND U8484 ( .A(init), .B(round_reg[164]), .Z(n2960) );
  NANDN U8485 ( .A(init), .B(in[164]), .Z(n2959) );
  NAND U8486 ( .A(n2960), .B(n2959), .Z(\round_in[0][164] ) );
  NAND U8487 ( .A(init), .B(round_reg[165]), .Z(n2962) );
  NANDN U8488 ( .A(init), .B(in[165]), .Z(n2961) );
  NAND U8489 ( .A(n2962), .B(n2961), .Z(\round_in[0][165] ) );
  NAND U8490 ( .A(init), .B(round_reg[166]), .Z(n2964) );
  NANDN U8491 ( .A(init), .B(in[166]), .Z(n2963) );
  NAND U8492 ( .A(n2964), .B(n2963), .Z(\round_in[0][166] ) );
  NAND U8493 ( .A(init), .B(round_reg[167]), .Z(n2966) );
  NANDN U8494 ( .A(init), .B(in[167]), .Z(n2965) );
  NAND U8495 ( .A(n2966), .B(n2965), .Z(\round_in[0][167] ) );
  NAND U8496 ( .A(init), .B(round_reg[168]), .Z(n2968) );
  NANDN U8497 ( .A(init), .B(in[168]), .Z(n2967) );
  NAND U8498 ( .A(n2968), .B(n2967), .Z(\round_in[0][168] ) );
  NAND U8499 ( .A(init), .B(round_reg[169]), .Z(n2970) );
  NANDN U8500 ( .A(init), .B(in[169]), .Z(n2969) );
  NAND U8501 ( .A(n2970), .B(n2969), .Z(\round_in[0][169] ) );
  NAND U8502 ( .A(init), .B(round_reg[16]), .Z(n2972) );
  NANDN U8503 ( .A(init), .B(in[16]), .Z(n2971) );
  NAND U8504 ( .A(n2972), .B(n2971), .Z(\round_in[0][16] ) );
  NAND U8505 ( .A(init), .B(round_reg[170]), .Z(n2974) );
  NANDN U8506 ( .A(init), .B(in[170]), .Z(n2973) );
  NAND U8507 ( .A(n2974), .B(n2973), .Z(\round_in[0][170] ) );
  NAND U8508 ( .A(init), .B(round_reg[171]), .Z(n2976) );
  NANDN U8509 ( .A(init), .B(in[171]), .Z(n2975) );
  NAND U8510 ( .A(n2976), .B(n2975), .Z(\round_in[0][171] ) );
  NAND U8511 ( .A(init), .B(round_reg[172]), .Z(n2978) );
  NANDN U8512 ( .A(init), .B(in[172]), .Z(n2977) );
  NAND U8513 ( .A(n2978), .B(n2977), .Z(\round_in[0][172] ) );
  NAND U8514 ( .A(init), .B(round_reg[173]), .Z(n2980) );
  NANDN U8515 ( .A(init), .B(in[173]), .Z(n2979) );
  NAND U8516 ( .A(n2980), .B(n2979), .Z(\round_in[0][173] ) );
  NAND U8517 ( .A(init), .B(round_reg[174]), .Z(n2982) );
  NANDN U8518 ( .A(init), .B(in[174]), .Z(n2981) );
  NAND U8519 ( .A(n2982), .B(n2981), .Z(\round_in[0][174] ) );
  NAND U8520 ( .A(init), .B(round_reg[175]), .Z(n2984) );
  NANDN U8521 ( .A(init), .B(in[175]), .Z(n2983) );
  NAND U8522 ( .A(n2984), .B(n2983), .Z(\round_in[0][175] ) );
  NAND U8523 ( .A(init), .B(round_reg[176]), .Z(n2986) );
  NANDN U8524 ( .A(init), .B(in[176]), .Z(n2985) );
  NAND U8525 ( .A(n2986), .B(n2985), .Z(\round_in[0][176] ) );
  NAND U8526 ( .A(init), .B(round_reg[177]), .Z(n2988) );
  NANDN U8527 ( .A(init), .B(in[177]), .Z(n2987) );
  NAND U8528 ( .A(n2988), .B(n2987), .Z(\round_in[0][177] ) );
  NAND U8529 ( .A(init), .B(round_reg[178]), .Z(n2990) );
  NANDN U8530 ( .A(init), .B(in[178]), .Z(n2989) );
  NAND U8531 ( .A(n2990), .B(n2989), .Z(\round_in[0][178] ) );
  NAND U8532 ( .A(init), .B(round_reg[179]), .Z(n2992) );
  NANDN U8533 ( .A(init), .B(in[179]), .Z(n2991) );
  NAND U8534 ( .A(n2992), .B(n2991), .Z(\round_in[0][179] ) );
  NAND U8535 ( .A(init), .B(round_reg[17]), .Z(n2994) );
  NANDN U8536 ( .A(init), .B(in[17]), .Z(n2993) );
  NAND U8537 ( .A(n2994), .B(n2993), .Z(\round_in[0][17] ) );
  NAND U8538 ( .A(init), .B(round_reg[180]), .Z(n2996) );
  NANDN U8539 ( .A(init), .B(in[180]), .Z(n2995) );
  NAND U8540 ( .A(n2996), .B(n2995), .Z(\round_in[0][180] ) );
  NAND U8541 ( .A(init), .B(round_reg[181]), .Z(n2998) );
  NANDN U8542 ( .A(init), .B(in[181]), .Z(n2997) );
  NAND U8543 ( .A(n2998), .B(n2997), .Z(\round_in[0][181] ) );
  NAND U8544 ( .A(init), .B(round_reg[182]), .Z(n3000) );
  NANDN U8545 ( .A(init), .B(in[182]), .Z(n2999) );
  NAND U8546 ( .A(n3000), .B(n2999), .Z(\round_in[0][182] ) );
  NAND U8547 ( .A(init), .B(round_reg[183]), .Z(n3002) );
  NANDN U8548 ( .A(init), .B(in[183]), .Z(n3001) );
  NAND U8549 ( .A(n3002), .B(n3001), .Z(\round_in[0][183] ) );
  NAND U8550 ( .A(init), .B(round_reg[184]), .Z(n3004) );
  NANDN U8551 ( .A(init), .B(in[184]), .Z(n3003) );
  NAND U8552 ( .A(n3004), .B(n3003), .Z(\round_in[0][184] ) );
  NAND U8553 ( .A(init), .B(round_reg[185]), .Z(n3006) );
  NANDN U8554 ( .A(init), .B(in[185]), .Z(n3005) );
  NAND U8555 ( .A(n3006), .B(n3005), .Z(\round_in[0][185] ) );
  NAND U8556 ( .A(init), .B(round_reg[186]), .Z(n3008) );
  NANDN U8557 ( .A(init), .B(in[186]), .Z(n3007) );
  NAND U8558 ( .A(n3008), .B(n3007), .Z(\round_in[0][186] ) );
  NAND U8559 ( .A(init), .B(round_reg[187]), .Z(n3010) );
  NANDN U8560 ( .A(init), .B(in[187]), .Z(n3009) );
  NAND U8561 ( .A(n3010), .B(n3009), .Z(\round_in[0][187] ) );
  NAND U8562 ( .A(init), .B(round_reg[188]), .Z(n3012) );
  NANDN U8563 ( .A(init), .B(in[188]), .Z(n3011) );
  NAND U8564 ( .A(n3012), .B(n3011), .Z(\round_in[0][188] ) );
  NAND U8565 ( .A(init), .B(round_reg[189]), .Z(n3014) );
  NANDN U8566 ( .A(init), .B(in[189]), .Z(n3013) );
  NAND U8567 ( .A(n3014), .B(n3013), .Z(\round_in[0][189] ) );
  NAND U8568 ( .A(init), .B(round_reg[18]), .Z(n3016) );
  NANDN U8569 ( .A(init), .B(in[18]), .Z(n3015) );
  NAND U8570 ( .A(n3016), .B(n3015), .Z(\round_in[0][18] ) );
  NAND U8571 ( .A(init), .B(round_reg[190]), .Z(n3018) );
  NANDN U8572 ( .A(init), .B(in[190]), .Z(n3017) );
  NAND U8573 ( .A(n3018), .B(n3017), .Z(\round_in[0][190] ) );
  NAND U8574 ( .A(init), .B(round_reg[191]), .Z(n3020) );
  NANDN U8575 ( .A(init), .B(in[191]), .Z(n3019) );
  NAND U8576 ( .A(n3020), .B(n3019), .Z(\round_in[0][191] ) );
  NAND U8577 ( .A(init), .B(round_reg[192]), .Z(n3022) );
  NANDN U8578 ( .A(init), .B(in[192]), .Z(n3021) );
  NAND U8579 ( .A(n3022), .B(n3021), .Z(\round_in[0][192] ) );
  NAND U8580 ( .A(init), .B(round_reg[193]), .Z(n3024) );
  NANDN U8581 ( .A(init), .B(in[193]), .Z(n3023) );
  NAND U8582 ( .A(n3024), .B(n3023), .Z(\round_in[0][193] ) );
  NAND U8583 ( .A(init), .B(round_reg[194]), .Z(n3026) );
  NANDN U8584 ( .A(init), .B(in[194]), .Z(n3025) );
  NAND U8585 ( .A(n3026), .B(n3025), .Z(\round_in[0][194] ) );
  NAND U8586 ( .A(init), .B(round_reg[195]), .Z(n3028) );
  NANDN U8587 ( .A(init), .B(in[195]), .Z(n3027) );
  NAND U8588 ( .A(n3028), .B(n3027), .Z(\round_in[0][195] ) );
  NAND U8589 ( .A(init), .B(round_reg[196]), .Z(n3030) );
  NANDN U8590 ( .A(init), .B(in[196]), .Z(n3029) );
  NAND U8591 ( .A(n3030), .B(n3029), .Z(\round_in[0][196] ) );
  NAND U8592 ( .A(init), .B(round_reg[197]), .Z(n3032) );
  NANDN U8593 ( .A(init), .B(in[197]), .Z(n3031) );
  NAND U8594 ( .A(n3032), .B(n3031), .Z(\round_in[0][197] ) );
  NAND U8595 ( .A(init), .B(round_reg[198]), .Z(n3034) );
  NANDN U8596 ( .A(init), .B(in[198]), .Z(n3033) );
  NAND U8597 ( .A(n3034), .B(n3033), .Z(\round_in[0][198] ) );
  NAND U8598 ( .A(init), .B(round_reg[199]), .Z(n3036) );
  NANDN U8599 ( .A(init), .B(in[199]), .Z(n3035) );
  NAND U8600 ( .A(n3036), .B(n3035), .Z(\round_in[0][199] ) );
  NAND U8601 ( .A(init), .B(round_reg[19]), .Z(n3038) );
  NANDN U8602 ( .A(init), .B(in[19]), .Z(n3037) );
  NAND U8603 ( .A(n3038), .B(n3037), .Z(\round_in[0][19] ) );
  NAND U8604 ( .A(init), .B(round_reg[1]), .Z(n3040) );
  NANDN U8605 ( .A(init), .B(in[1]), .Z(n3039) );
  NAND U8606 ( .A(n3040), .B(n3039), .Z(\round_in[0][1] ) );
  NAND U8607 ( .A(init), .B(round_reg[200]), .Z(n3042) );
  NANDN U8608 ( .A(init), .B(in[200]), .Z(n3041) );
  NAND U8609 ( .A(n3042), .B(n3041), .Z(\round_in[0][200] ) );
  NAND U8610 ( .A(init), .B(round_reg[201]), .Z(n3044) );
  NANDN U8611 ( .A(init), .B(in[201]), .Z(n3043) );
  NAND U8612 ( .A(n3044), .B(n3043), .Z(\round_in[0][201] ) );
  NAND U8613 ( .A(init), .B(round_reg[202]), .Z(n3046) );
  NANDN U8614 ( .A(init), .B(in[202]), .Z(n3045) );
  NAND U8615 ( .A(n3046), .B(n3045), .Z(\round_in[0][202] ) );
  NAND U8616 ( .A(init), .B(round_reg[203]), .Z(n3048) );
  NANDN U8617 ( .A(init), .B(in[203]), .Z(n3047) );
  NAND U8618 ( .A(n3048), .B(n3047), .Z(\round_in[0][203] ) );
  NAND U8619 ( .A(init), .B(round_reg[204]), .Z(n3050) );
  NANDN U8620 ( .A(init), .B(in[204]), .Z(n3049) );
  NAND U8621 ( .A(n3050), .B(n3049), .Z(\round_in[0][204] ) );
  NAND U8622 ( .A(init), .B(round_reg[205]), .Z(n3052) );
  NANDN U8623 ( .A(init), .B(in[205]), .Z(n3051) );
  NAND U8624 ( .A(n3052), .B(n3051), .Z(\round_in[0][205] ) );
  NAND U8625 ( .A(init), .B(round_reg[206]), .Z(n3054) );
  NANDN U8626 ( .A(init), .B(in[206]), .Z(n3053) );
  NAND U8627 ( .A(n3054), .B(n3053), .Z(\round_in[0][206] ) );
  NAND U8628 ( .A(init), .B(round_reg[207]), .Z(n3056) );
  NANDN U8629 ( .A(init), .B(in[207]), .Z(n3055) );
  NAND U8630 ( .A(n3056), .B(n3055), .Z(\round_in[0][207] ) );
  NAND U8631 ( .A(init), .B(round_reg[208]), .Z(n3058) );
  NANDN U8632 ( .A(init), .B(in[208]), .Z(n3057) );
  NAND U8633 ( .A(n3058), .B(n3057), .Z(\round_in[0][208] ) );
  NAND U8634 ( .A(init), .B(round_reg[209]), .Z(n3060) );
  NANDN U8635 ( .A(init), .B(in[209]), .Z(n3059) );
  NAND U8636 ( .A(n3060), .B(n3059), .Z(\round_in[0][209] ) );
  NAND U8637 ( .A(init), .B(round_reg[20]), .Z(n3062) );
  NANDN U8638 ( .A(init), .B(in[20]), .Z(n3061) );
  NAND U8639 ( .A(n3062), .B(n3061), .Z(\round_in[0][20] ) );
  NAND U8640 ( .A(init), .B(round_reg[210]), .Z(n3064) );
  NANDN U8641 ( .A(init), .B(in[210]), .Z(n3063) );
  NAND U8642 ( .A(n3064), .B(n3063), .Z(\round_in[0][210] ) );
  NAND U8643 ( .A(init), .B(round_reg[211]), .Z(n3066) );
  NANDN U8644 ( .A(init), .B(in[211]), .Z(n3065) );
  NAND U8645 ( .A(n3066), .B(n3065), .Z(\round_in[0][211] ) );
  NAND U8646 ( .A(init), .B(round_reg[212]), .Z(n3068) );
  NANDN U8647 ( .A(init), .B(in[212]), .Z(n3067) );
  NAND U8648 ( .A(n3068), .B(n3067), .Z(\round_in[0][212] ) );
  NAND U8649 ( .A(init), .B(round_reg[213]), .Z(n3070) );
  NANDN U8650 ( .A(init), .B(in[213]), .Z(n3069) );
  NAND U8651 ( .A(n3070), .B(n3069), .Z(\round_in[0][213] ) );
  NAND U8652 ( .A(init), .B(round_reg[214]), .Z(n3072) );
  NANDN U8653 ( .A(init), .B(in[214]), .Z(n3071) );
  NAND U8654 ( .A(n3072), .B(n3071), .Z(\round_in[0][214] ) );
  NAND U8655 ( .A(init), .B(round_reg[215]), .Z(n3074) );
  NANDN U8656 ( .A(init), .B(in[215]), .Z(n3073) );
  NAND U8657 ( .A(n3074), .B(n3073), .Z(\round_in[0][215] ) );
  NAND U8658 ( .A(init), .B(round_reg[216]), .Z(n3076) );
  NANDN U8659 ( .A(init), .B(in[216]), .Z(n3075) );
  NAND U8660 ( .A(n3076), .B(n3075), .Z(\round_in[0][216] ) );
  NAND U8661 ( .A(init), .B(round_reg[217]), .Z(n3078) );
  NANDN U8662 ( .A(init), .B(in[217]), .Z(n3077) );
  NAND U8663 ( .A(n3078), .B(n3077), .Z(\round_in[0][217] ) );
  NAND U8664 ( .A(init), .B(round_reg[218]), .Z(n3080) );
  NANDN U8665 ( .A(init), .B(in[218]), .Z(n3079) );
  NAND U8666 ( .A(n3080), .B(n3079), .Z(\round_in[0][218] ) );
  NAND U8667 ( .A(init), .B(round_reg[219]), .Z(n3082) );
  NANDN U8668 ( .A(init), .B(in[219]), .Z(n3081) );
  NAND U8669 ( .A(n3082), .B(n3081), .Z(\round_in[0][219] ) );
  NAND U8670 ( .A(init), .B(round_reg[21]), .Z(n3084) );
  NANDN U8671 ( .A(init), .B(in[21]), .Z(n3083) );
  NAND U8672 ( .A(n3084), .B(n3083), .Z(\round_in[0][21] ) );
  NAND U8673 ( .A(init), .B(round_reg[220]), .Z(n3086) );
  NANDN U8674 ( .A(init), .B(in[220]), .Z(n3085) );
  NAND U8675 ( .A(n3086), .B(n3085), .Z(\round_in[0][220] ) );
  NAND U8676 ( .A(init), .B(round_reg[221]), .Z(n3088) );
  NANDN U8677 ( .A(init), .B(in[221]), .Z(n3087) );
  NAND U8678 ( .A(n3088), .B(n3087), .Z(\round_in[0][221] ) );
  NAND U8679 ( .A(init), .B(round_reg[222]), .Z(n3090) );
  NANDN U8680 ( .A(init), .B(in[222]), .Z(n3089) );
  NAND U8681 ( .A(n3090), .B(n3089), .Z(\round_in[0][222] ) );
  NAND U8682 ( .A(init), .B(round_reg[223]), .Z(n3092) );
  NANDN U8683 ( .A(init), .B(in[223]), .Z(n3091) );
  NAND U8684 ( .A(n3092), .B(n3091), .Z(\round_in[0][223] ) );
  NAND U8685 ( .A(init), .B(round_reg[224]), .Z(n3094) );
  NANDN U8686 ( .A(init), .B(in[224]), .Z(n3093) );
  NAND U8687 ( .A(n3094), .B(n3093), .Z(\round_in[0][224] ) );
  NAND U8688 ( .A(init), .B(round_reg[225]), .Z(n3096) );
  NANDN U8689 ( .A(init), .B(in[225]), .Z(n3095) );
  NAND U8690 ( .A(n3096), .B(n3095), .Z(\round_in[0][225] ) );
  NAND U8691 ( .A(init), .B(round_reg[226]), .Z(n3098) );
  NANDN U8692 ( .A(init), .B(in[226]), .Z(n3097) );
  NAND U8693 ( .A(n3098), .B(n3097), .Z(\round_in[0][226] ) );
  NAND U8694 ( .A(init), .B(round_reg[227]), .Z(n3100) );
  NANDN U8695 ( .A(init), .B(in[227]), .Z(n3099) );
  NAND U8696 ( .A(n3100), .B(n3099), .Z(\round_in[0][227] ) );
  NAND U8697 ( .A(init), .B(round_reg[228]), .Z(n3102) );
  NANDN U8698 ( .A(init), .B(in[228]), .Z(n3101) );
  NAND U8699 ( .A(n3102), .B(n3101), .Z(\round_in[0][228] ) );
  NAND U8700 ( .A(init), .B(round_reg[229]), .Z(n3104) );
  NANDN U8701 ( .A(init), .B(in[229]), .Z(n3103) );
  NAND U8702 ( .A(n3104), .B(n3103), .Z(\round_in[0][229] ) );
  NAND U8703 ( .A(init), .B(round_reg[22]), .Z(n3106) );
  NANDN U8704 ( .A(init), .B(in[22]), .Z(n3105) );
  NAND U8705 ( .A(n3106), .B(n3105), .Z(\round_in[0][22] ) );
  NAND U8706 ( .A(init), .B(round_reg[230]), .Z(n3108) );
  NANDN U8707 ( .A(init), .B(in[230]), .Z(n3107) );
  NAND U8708 ( .A(n3108), .B(n3107), .Z(\round_in[0][230] ) );
  NAND U8709 ( .A(init), .B(round_reg[231]), .Z(n3110) );
  NANDN U8710 ( .A(init), .B(in[231]), .Z(n3109) );
  NAND U8711 ( .A(n3110), .B(n3109), .Z(\round_in[0][231] ) );
  NAND U8712 ( .A(init), .B(round_reg[232]), .Z(n3112) );
  NANDN U8713 ( .A(init), .B(in[232]), .Z(n3111) );
  NAND U8714 ( .A(n3112), .B(n3111), .Z(\round_in[0][232] ) );
  NAND U8715 ( .A(init), .B(round_reg[233]), .Z(n3114) );
  NANDN U8716 ( .A(init), .B(in[233]), .Z(n3113) );
  NAND U8717 ( .A(n3114), .B(n3113), .Z(\round_in[0][233] ) );
  NAND U8718 ( .A(init), .B(round_reg[234]), .Z(n3116) );
  NANDN U8719 ( .A(init), .B(in[234]), .Z(n3115) );
  NAND U8720 ( .A(n3116), .B(n3115), .Z(\round_in[0][234] ) );
  NAND U8721 ( .A(init), .B(round_reg[235]), .Z(n3118) );
  NANDN U8722 ( .A(init), .B(in[235]), .Z(n3117) );
  NAND U8723 ( .A(n3118), .B(n3117), .Z(\round_in[0][235] ) );
  NAND U8724 ( .A(init), .B(round_reg[236]), .Z(n3120) );
  NANDN U8725 ( .A(init), .B(in[236]), .Z(n3119) );
  NAND U8726 ( .A(n3120), .B(n3119), .Z(\round_in[0][236] ) );
  NAND U8727 ( .A(init), .B(round_reg[237]), .Z(n3122) );
  NANDN U8728 ( .A(init), .B(in[237]), .Z(n3121) );
  NAND U8729 ( .A(n3122), .B(n3121), .Z(\round_in[0][237] ) );
  NAND U8730 ( .A(init), .B(round_reg[238]), .Z(n3124) );
  NANDN U8731 ( .A(init), .B(in[238]), .Z(n3123) );
  NAND U8732 ( .A(n3124), .B(n3123), .Z(\round_in[0][238] ) );
  NAND U8733 ( .A(init), .B(round_reg[239]), .Z(n3126) );
  NANDN U8734 ( .A(init), .B(in[239]), .Z(n3125) );
  NAND U8735 ( .A(n3126), .B(n3125), .Z(\round_in[0][239] ) );
  NAND U8736 ( .A(init), .B(round_reg[23]), .Z(n3128) );
  NANDN U8737 ( .A(init), .B(in[23]), .Z(n3127) );
  NAND U8738 ( .A(n3128), .B(n3127), .Z(\round_in[0][23] ) );
  NAND U8739 ( .A(init), .B(round_reg[240]), .Z(n3130) );
  NANDN U8740 ( .A(init), .B(in[240]), .Z(n3129) );
  NAND U8741 ( .A(n3130), .B(n3129), .Z(\round_in[0][240] ) );
  NAND U8742 ( .A(init), .B(round_reg[241]), .Z(n3132) );
  NANDN U8743 ( .A(init), .B(in[241]), .Z(n3131) );
  NAND U8744 ( .A(n3132), .B(n3131), .Z(\round_in[0][241] ) );
  NAND U8745 ( .A(init), .B(round_reg[242]), .Z(n3134) );
  NANDN U8746 ( .A(init), .B(in[242]), .Z(n3133) );
  NAND U8747 ( .A(n3134), .B(n3133), .Z(\round_in[0][242] ) );
  NAND U8748 ( .A(init), .B(round_reg[243]), .Z(n3136) );
  NANDN U8749 ( .A(init), .B(in[243]), .Z(n3135) );
  NAND U8750 ( .A(n3136), .B(n3135), .Z(\round_in[0][243] ) );
  NAND U8751 ( .A(init), .B(round_reg[244]), .Z(n3138) );
  NANDN U8752 ( .A(init), .B(in[244]), .Z(n3137) );
  NAND U8753 ( .A(n3138), .B(n3137), .Z(\round_in[0][244] ) );
  NAND U8754 ( .A(init), .B(round_reg[245]), .Z(n3140) );
  NANDN U8755 ( .A(init), .B(in[245]), .Z(n3139) );
  NAND U8756 ( .A(n3140), .B(n3139), .Z(\round_in[0][245] ) );
  NAND U8757 ( .A(init), .B(round_reg[246]), .Z(n3142) );
  NANDN U8758 ( .A(init), .B(in[246]), .Z(n3141) );
  NAND U8759 ( .A(n3142), .B(n3141), .Z(\round_in[0][246] ) );
  NAND U8760 ( .A(init), .B(round_reg[247]), .Z(n3144) );
  NANDN U8761 ( .A(init), .B(in[247]), .Z(n3143) );
  NAND U8762 ( .A(n3144), .B(n3143), .Z(\round_in[0][247] ) );
  NAND U8763 ( .A(init), .B(round_reg[248]), .Z(n3146) );
  NANDN U8764 ( .A(init), .B(in[248]), .Z(n3145) );
  NAND U8765 ( .A(n3146), .B(n3145), .Z(\round_in[0][248] ) );
  NAND U8766 ( .A(init), .B(round_reg[249]), .Z(n3148) );
  NANDN U8767 ( .A(init), .B(in[249]), .Z(n3147) );
  NAND U8768 ( .A(n3148), .B(n3147), .Z(\round_in[0][249] ) );
  NAND U8769 ( .A(init), .B(round_reg[24]), .Z(n3150) );
  NANDN U8770 ( .A(init), .B(in[24]), .Z(n3149) );
  NAND U8771 ( .A(n3150), .B(n3149), .Z(\round_in[0][24] ) );
  NAND U8772 ( .A(init), .B(round_reg[250]), .Z(n3152) );
  NANDN U8773 ( .A(init), .B(in[250]), .Z(n3151) );
  NAND U8774 ( .A(n3152), .B(n3151), .Z(\round_in[0][250] ) );
  NAND U8775 ( .A(init), .B(round_reg[251]), .Z(n3154) );
  NANDN U8776 ( .A(init), .B(in[251]), .Z(n3153) );
  NAND U8777 ( .A(n3154), .B(n3153), .Z(\round_in[0][251] ) );
  NAND U8778 ( .A(init), .B(round_reg[252]), .Z(n3156) );
  NANDN U8779 ( .A(init), .B(in[252]), .Z(n3155) );
  NAND U8780 ( .A(n3156), .B(n3155), .Z(\round_in[0][252] ) );
  NAND U8781 ( .A(init), .B(round_reg[253]), .Z(n3158) );
  NANDN U8782 ( .A(init), .B(in[253]), .Z(n3157) );
  NAND U8783 ( .A(n3158), .B(n3157), .Z(\round_in[0][253] ) );
  NAND U8784 ( .A(init), .B(round_reg[254]), .Z(n3160) );
  NANDN U8785 ( .A(init), .B(in[254]), .Z(n3159) );
  NAND U8786 ( .A(n3160), .B(n3159), .Z(\round_in[0][254] ) );
  NAND U8787 ( .A(init), .B(round_reg[255]), .Z(n3162) );
  NANDN U8788 ( .A(init), .B(in[255]), .Z(n3161) );
  NAND U8789 ( .A(n3162), .B(n3161), .Z(\round_in[0][255] ) );
  NAND U8790 ( .A(init), .B(round_reg[256]), .Z(n3164) );
  NANDN U8791 ( .A(init), .B(in[256]), .Z(n3163) );
  NAND U8792 ( .A(n3164), .B(n3163), .Z(\round_in[0][256] ) );
  NAND U8793 ( .A(init), .B(round_reg[257]), .Z(n3166) );
  NANDN U8794 ( .A(init), .B(in[257]), .Z(n3165) );
  NAND U8795 ( .A(n3166), .B(n3165), .Z(\round_in[0][257] ) );
  NAND U8796 ( .A(init), .B(round_reg[258]), .Z(n3168) );
  NANDN U8797 ( .A(init), .B(in[258]), .Z(n3167) );
  NAND U8798 ( .A(n3168), .B(n3167), .Z(\round_in[0][258] ) );
  NAND U8799 ( .A(init), .B(round_reg[259]), .Z(n3170) );
  NANDN U8800 ( .A(init), .B(in[259]), .Z(n3169) );
  NAND U8801 ( .A(n3170), .B(n3169), .Z(\round_in[0][259] ) );
  NAND U8802 ( .A(init), .B(round_reg[25]), .Z(n3172) );
  NANDN U8803 ( .A(init), .B(in[25]), .Z(n3171) );
  NAND U8804 ( .A(n3172), .B(n3171), .Z(\round_in[0][25] ) );
  NAND U8805 ( .A(init), .B(round_reg[260]), .Z(n3174) );
  NANDN U8806 ( .A(init), .B(in[260]), .Z(n3173) );
  NAND U8807 ( .A(n3174), .B(n3173), .Z(\round_in[0][260] ) );
  NAND U8808 ( .A(init), .B(round_reg[261]), .Z(n3176) );
  NANDN U8809 ( .A(init), .B(in[261]), .Z(n3175) );
  NAND U8810 ( .A(n3176), .B(n3175), .Z(\round_in[0][261] ) );
  NAND U8811 ( .A(init), .B(round_reg[262]), .Z(n3178) );
  NANDN U8812 ( .A(init), .B(in[262]), .Z(n3177) );
  NAND U8813 ( .A(n3178), .B(n3177), .Z(\round_in[0][262] ) );
  NAND U8814 ( .A(init), .B(round_reg[263]), .Z(n3180) );
  NANDN U8815 ( .A(init), .B(in[263]), .Z(n3179) );
  NAND U8816 ( .A(n3180), .B(n3179), .Z(\round_in[0][263] ) );
  NAND U8817 ( .A(init), .B(round_reg[264]), .Z(n3182) );
  NANDN U8818 ( .A(init), .B(in[264]), .Z(n3181) );
  NAND U8819 ( .A(n3182), .B(n3181), .Z(\round_in[0][264] ) );
  NAND U8820 ( .A(init), .B(round_reg[265]), .Z(n3184) );
  NANDN U8821 ( .A(init), .B(in[265]), .Z(n3183) );
  NAND U8822 ( .A(n3184), .B(n3183), .Z(\round_in[0][265] ) );
  NAND U8823 ( .A(init), .B(round_reg[266]), .Z(n3186) );
  NANDN U8824 ( .A(init), .B(in[266]), .Z(n3185) );
  NAND U8825 ( .A(n3186), .B(n3185), .Z(\round_in[0][266] ) );
  NAND U8826 ( .A(init), .B(round_reg[267]), .Z(n3188) );
  NANDN U8827 ( .A(init), .B(in[267]), .Z(n3187) );
  NAND U8828 ( .A(n3188), .B(n3187), .Z(\round_in[0][267] ) );
  NAND U8829 ( .A(init), .B(round_reg[268]), .Z(n3190) );
  NANDN U8830 ( .A(init), .B(in[268]), .Z(n3189) );
  NAND U8831 ( .A(n3190), .B(n3189), .Z(\round_in[0][268] ) );
  NAND U8832 ( .A(init), .B(round_reg[269]), .Z(n3192) );
  NANDN U8833 ( .A(init), .B(in[269]), .Z(n3191) );
  NAND U8834 ( .A(n3192), .B(n3191), .Z(\round_in[0][269] ) );
  NAND U8835 ( .A(init), .B(round_reg[26]), .Z(n3194) );
  NANDN U8836 ( .A(init), .B(in[26]), .Z(n3193) );
  NAND U8837 ( .A(n3194), .B(n3193), .Z(\round_in[0][26] ) );
  NAND U8838 ( .A(init), .B(round_reg[270]), .Z(n3196) );
  NANDN U8839 ( .A(init), .B(in[270]), .Z(n3195) );
  NAND U8840 ( .A(n3196), .B(n3195), .Z(\round_in[0][270] ) );
  NAND U8841 ( .A(init), .B(round_reg[271]), .Z(n3198) );
  NANDN U8842 ( .A(init), .B(in[271]), .Z(n3197) );
  NAND U8843 ( .A(n3198), .B(n3197), .Z(\round_in[0][271] ) );
  NAND U8844 ( .A(init), .B(round_reg[272]), .Z(n3200) );
  NANDN U8845 ( .A(init), .B(in[272]), .Z(n3199) );
  NAND U8846 ( .A(n3200), .B(n3199), .Z(\round_in[0][272] ) );
  NAND U8847 ( .A(init), .B(round_reg[273]), .Z(n3202) );
  NANDN U8848 ( .A(init), .B(in[273]), .Z(n3201) );
  NAND U8849 ( .A(n3202), .B(n3201), .Z(\round_in[0][273] ) );
  NAND U8850 ( .A(init), .B(round_reg[274]), .Z(n3204) );
  NANDN U8851 ( .A(init), .B(in[274]), .Z(n3203) );
  NAND U8852 ( .A(n3204), .B(n3203), .Z(\round_in[0][274] ) );
  NAND U8853 ( .A(init), .B(round_reg[275]), .Z(n3206) );
  NANDN U8854 ( .A(init), .B(in[275]), .Z(n3205) );
  NAND U8855 ( .A(n3206), .B(n3205), .Z(\round_in[0][275] ) );
  NAND U8856 ( .A(init), .B(round_reg[276]), .Z(n3208) );
  NANDN U8857 ( .A(init), .B(in[276]), .Z(n3207) );
  NAND U8858 ( .A(n3208), .B(n3207), .Z(\round_in[0][276] ) );
  NAND U8859 ( .A(init), .B(round_reg[277]), .Z(n3210) );
  NANDN U8860 ( .A(init), .B(in[277]), .Z(n3209) );
  NAND U8861 ( .A(n3210), .B(n3209), .Z(\round_in[0][277] ) );
  NAND U8862 ( .A(init), .B(round_reg[278]), .Z(n3212) );
  NANDN U8863 ( .A(init), .B(in[278]), .Z(n3211) );
  NAND U8864 ( .A(n3212), .B(n3211), .Z(\round_in[0][278] ) );
  NAND U8865 ( .A(init), .B(round_reg[279]), .Z(n3214) );
  NANDN U8866 ( .A(init), .B(in[279]), .Z(n3213) );
  NAND U8867 ( .A(n3214), .B(n3213), .Z(\round_in[0][279] ) );
  NAND U8868 ( .A(init), .B(round_reg[27]), .Z(n3216) );
  NANDN U8869 ( .A(init), .B(in[27]), .Z(n3215) );
  NAND U8870 ( .A(n3216), .B(n3215), .Z(\round_in[0][27] ) );
  NAND U8871 ( .A(init), .B(round_reg[280]), .Z(n3218) );
  NANDN U8872 ( .A(init), .B(in[280]), .Z(n3217) );
  NAND U8873 ( .A(n3218), .B(n3217), .Z(\round_in[0][280] ) );
  NAND U8874 ( .A(init), .B(round_reg[281]), .Z(n3220) );
  NANDN U8875 ( .A(init), .B(in[281]), .Z(n3219) );
  NAND U8876 ( .A(n3220), .B(n3219), .Z(\round_in[0][281] ) );
  NAND U8877 ( .A(init), .B(round_reg[282]), .Z(n3222) );
  NANDN U8878 ( .A(init), .B(in[282]), .Z(n3221) );
  NAND U8879 ( .A(n3222), .B(n3221), .Z(\round_in[0][282] ) );
  NAND U8880 ( .A(init), .B(round_reg[283]), .Z(n3224) );
  NANDN U8881 ( .A(init), .B(in[283]), .Z(n3223) );
  NAND U8882 ( .A(n3224), .B(n3223), .Z(\round_in[0][283] ) );
  NAND U8883 ( .A(init), .B(round_reg[284]), .Z(n3226) );
  NANDN U8884 ( .A(init), .B(in[284]), .Z(n3225) );
  NAND U8885 ( .A(n3226), .B(n3225), .Z(\round_in[0][284] ) );
  NAND U8886 ( .A(init), .B(round_reg[285]), .Z(n3228) );
  NANDN U8887 ( .A(init), .B(in[285]), .Z(n3227) );
  NAND U8888 ( .A(n3228), .B(n3227), .Z(\round_in[0][285] ) );
  NAND U8889 ( .A(init), .B(round_reg[286]), .Z(n3230) );
  NANDN U8890 ( .A(init), .B(in[286]), .Z(n3229) );
  NAND U8891 ( .A(n3230), .B(n3229), .Z(\round_in[0][286] ) );
  NAND U8892 ( .A(init), .B(round_reg[287]), .Z(n3232) );
  NANDN U8893 ( .A(init), .B(in[287]), .Z(n3231) );
  NAND U8894 ( .A(n3232), .B(n3231), .Z(\round_in[0][287] ) );
  NAND U8895 ( .A(init), .B(round_reg[288]), .Z(n3234) );
  NANDN U8896 ( .A(init), .B(in[288]), .Z(n3233) );
  NAND U8897 ( .A(n3234), .B(n3233), .Z(\round_in[0][288] ) );
  NAND U8898 ( .A(init), .B(round_reg[289]), .Z(n3236) );
  NANDN U8899 ( .A(init), .B(in[289]), .Z(n3235) );
  NAND U8900 ( .A(n3236), .B(n3235), .Z(\round_in[0][289] ) );
  NAND U8901 ( .A(init), .B(round_reg[28]), .Z(n3238) );
  NANDN U8902 ( .A(init), .B(in[28]), .Z(n3237) );
  NAND U8903 ( .A(n3238), .B(n3237), .Z(\round_in[0][28] ) );
  NAND U8904 ( .A(init), .B(round_reg[290]), .Z(n3240) );
  NANDN U8905 ( .A(init), .B(in[290]), .Z(n3239) );
  NAND U8906 ( .A(n3240), .B(n3239), .Z(\round_in[0][290] ) );
  NAND U8907 ( .A(init), .B(round_reg[291]), .Z(n3242) );
  NANDN U8908 ( .A(init), .B(in[291]), .Z(n3241) );
  NAND U8909 ( .A(n3242), .B(n3241), .Z(\round_in[0][291] ) );
  NAND U8910 ( .A(init), .B(round_reg[292]), .Z(n3244) );
  NANDN U8911 ( .A(init), .B(in[292]), .Z(n3243) );
  NAND U8912 ( .A(n3244), .B(n3243), .Z(\round_in[0][292] ) );
  NAND U8913 ( .A(init), .B(round_reg[293]), .Z(n3246) );
  NANDN U8914 ( .A(init), .B(in[293]), .Z(n3245) );
  NAND U8915 ( .A(n3246), .B(n3245), .Z(\round_in[0][293] ) );
  NAND U8916 ( .A(init), .B(round_reg[294]), .Z(n3248) );
  NANDN U8917 ( .A(init), .B(in[294]), .Z(n3247) );
  NAND U8918 ( .A(n3248), .B(n3247), .Z(\round_in[0][294] ) );
  NAND U8919 ( .A(init), .B(round_reg[295]), .Z(n3250) );
  NANDN U8920 ( .A(init), .B(in[295]), .Z(n3249) );
  NAND U8921 ( .A(n3250), .B(n3249), .Z(\round_in[0][295] ) );
  NAND U8922 ( .A(init), .B(round_reg[296]), .Z(n3252) );
  NANDN U8923 ( .A(init), .B(in[296]), .Z(n3251) );
  NAND U8924 ( .A(n3252), .B(n3251), .Z(\round_in[0][296] ) );
  NAND U8925 ( .A(init), .B(round_reg[297]), .Z(n3254) );
  NANDN U8926 ( .A(init), .B(in[297]), .Z(n3253) );
  NAND U8927 ( .A(n3254), .B(n3253), .Z(\round_in[0][297] ) );
  NAND U8928 ( .A(init), .B(round_reg[298]), .Z(n3256) );
  NANDN U8929 ( .A(init), .B(in[298]), .Z(n3255) );
  NAND U8930 ( .A(n3256), .B(n3255), .Z(\round_in[0][298] ) );
  NAND U8931 ( .A(init), .B(round_reg[299]), .Z(n3258) );
  NANDN U8932 ( .A(init), .B(in[299]), .Z(n3257) );
  NAND U8933 ( .A(n3258), .B(n3257), .Z(\round_in[0][299] ) );
  NAND U8934 ( .A(init), .B(round_reg[29]), .Z(n3260) );
  NANDN U8935 ( .A(init), .B(in[29]), .Z(n3259) );
  NAND U8936 ( .A(n3260), .B(n3259), .Z(\round_in[0][29] ) );
  NAND U8937 ( .A(init), .B(round_reg[2]), .Z(n3262) );
  NANDN U8938 ( .A(init), .B(in[2]), .Z(n3261) );
  NAND U8939 ( .A(n3262), .B(n3261), .Z(\round_in[0][2] ) );
  NAND U8940 ( .A(init), .B(round_reg[300]), .Z(n3264) );
  NANDN U8941 ( .A(init), .B(in[300]), .Z(n3263) );
  NAND U8942 ( .A(n3264), .B(n3263), .Z(\round_in[0][300] ) );
  NAND U8943 ( .A(init), .B(round_reg[301]), .Z(n3266) );
  NANDN U8944 ( .A(init), .B(in[301]), .Z(n3265) );
  NAND U8945 ( .A(n3266), .B(n3265), .Z(\round_in[0][301] ) );
  NAND U8946 ( .A(init), .B(round_reg[302]), .Z(n3268) );
  NANDN U8947 ( .A(init), .B(in[302]), .Z(n3267) );
  NAND U8948 ( .A(n3268), .B(n3267), .Z(\round_in[0][302] ) );
  NAND U8949 ( .A(init), .B(round_reg[303]), .Z(n3270) );
  NANDN U8950 ( .A(init), .B(in[303]), .Z(n3269) );
  NAND U8951 ( .A(n3270), .B(n3269), .Z(\round_in[0][303] ) );
  NAND U8952 ( .A(init), .B(round_reg[304]), .Z(n3272) );
  NANDN U8953 ( .A(init), .B(in[304]), .Z(n3271) );
  NAND U8954 ( .A(n3272), .B(n3271), .Z(\round_in[0][304] ) );
  NAND U8955 ( .A(init), .B(round_reg[305]), .Z(n3274) );
  NANDN U8956 ( .A(init), .B(in[305]), .Z(n3273) );
  NAND U8957 ( .A(n3274), .B(n3273), .Z(\round_in[0][305] ) );
  NAND U8958 ( .A(init), .B(round_reg[306]), .Z(n3276) );
  NANDN U8959 ( .A(init), .B(in[306]), .Z(n3275) );
  NAND U8960 ( .A(n3276), .B(n3275), .Z(\round_in[0][306] ) );
  NAND U8961 ( .A(init), .B(round_reg[307]), .Z(n3278) );
  NANDN U8962 ( .A(init), .B(in[307]), .Z(n3277) );
  NAND U8963 ( .A(n3278), .B(n3277), .Z(\round_in[0][307] ) );
  NAND U8964 ( .A(init), .B(round_reg[308]), .Z(n3280) );
  NANDN U8965 ( .A(init), .B(in[308]), .Z(n3279) );
  NAND U8966 ( .A(n3280), .B(n3279), .Z(\round_in[0][308] ) );
  NAND U8967 ( .A(init), .B(round_reg[309]), .Z(n3282) );
  NANDN U8968 ( .A(init), .B(in[309]), .Z(n3281) );
  NAND U8969 ( .A(n3282), .B(n3281), .Z(\round_in[0][309] ) );
  NAND U8970 ( .A(init), .B(round_reg[30]), .Z(n3284) );
  NANDN U8971 ( .A(init), .B(in[30]), .Z(n3283) );
  NAND U8972 ( .A(n3284), .B(n3283), .Z(\round_in[0][30] ) );
  NAND U8973 ( .A(init), .B(round_reg[310]), .Z(n3286) );
  NANDN U8974 ( .A(init), .B(in[310]), .Z(n3285) );
  NAND U8975 ( .A(n3286), .B(n3285), .Z(\round_in[0][310] ) );
  NAND U8976 ( .A(init), .B(round_reg[311]), .Z(n3288) );
  NANDN U8977 ( .A(init), .B(in[311]), .Z(n3287) );
  NAND U8978 ( .A(n3288), .B(n3287), .Z(\round_in[0][311] ) );
  NAND U8979 ( .A(init), .B(round_reg[312]), .Z(n3290) );
  NANDN U8980 ( .A(init), .B(in[312]), .Z(n3289) );
  NAND U8981 ( .A(n3290), .B(n3289), .Z(\round_in[0][312] ) );
  NAND U8982 ( .A(init), .B(round_reg[313]), .Z(n3292) );
  NANDN U8983 ( .A(init), .B(in[313]), .Z(n3291) );
  NAND U8984 ( .A(n3292), .B(n3291), .Z(\round_in[0][313] ) );
  NAND U8985 ( .A(init), .B(round_reg[314]), .Z(n3294) );
  NANDN U8986 ( .A(init), .B(in[314]), .Z(n3293) );
  NAND U8987 ( .A(n3294), .B(n3293), .Z(\round_in[0][314] ) );
  NAND U8988 ( .A(init), .B(round_reg[315]), .Z(n3296) );
  NANDN U8989 ( .A(init), .B(in[315]), .Z(n3295) );
  NAND U8990 ( .A(n3296), .B(n3295), .Z(\round_in[0][315] ) );
  NAND U8991 ( .A(init), .B(round_reg[316]), .Z(n3298) );
  NANDN U8992 ( .A(init), .B(in[316]), .Z(n3297) );
  NAND U8993 ( .A(n3298), .B(n3297), .Z(\round_in[0][316] ) );
  NAND U8994 ( .A(init), .B(round_reg[317]), .Z(n3300) );
  NANDN U8995 ( .A(init), .B(in[317]), .Z(n3299) );
  NAND U8996 ( .A(n3300), .B(n3299), .Z(\round_in[0][317] ) );
  NAND U8997 ( .A(init), .B(round_reg[318]), .Z(n3302) );
  NANDN U8998 ( .A(init), .B(in[318]), .Z(n3301) );
  NAND U8999 ( .A(n3302), .B(n3301), .Z(\round_in[0][318] ) );
  NAND U9000 ( .A(init), .B(round_reg[319]), .Z(n3304) );
  NANDN U9001 ( .A(init), .B(in[319]), .Z(n3303) );
  NAND U9002 ( .A(n3304), .B(n3303), .Z(\round_in[0][319] ) );
  NAND U9003 ( .A(init), .B(round_reg[31]), .Z(n3306) );
  NANDN U9004 ( .A(init), .B(in[31]), .Z(n3305) );
  NAND U9005 ( .A(n3306), .B(n3305), .Z(\round_in[0][31] ) );
  NAND U9006 ( .A(init), .B(round_reg[320]), .Z(n3308) );
  NANDN U9007 ( .A(init), .B(in[320]), .Z(n3307) );
  NAND U9008 ( .A(n3308), .B(n3307), .Z(\round_in[0][320] ) );
  NAND U9009 ( .A(init), .B(round_reg[321]), .Z(n3310) );
  NANDN U9010 ( .A(init), .B(in[321]), .Z(n3309) );
  NAND U9011 ( .A(n3310), .B(n3309), .Z(\round_in[0][321] ) );
  NAND U9012 ( .A(init), .B(round_reg[322]), .Z(n3312) );
  NANDN U9013 ( .A(init), .B(in[322]), .Z(n3311) );
  NAND U9014 ( .A(n3312), .B(n3311), .Z(\round_in[0][322] ) );
  NAND U9015 ( .A(init), .B(round_reg[323]), .Z(n3314) );
  NANDN U9016 ( .A(init), .B(in[323]), .Z(n3313) );
  NAND U9017 ( .A(n3314), .B(n3313), .Z(\round_in[0][323] ) );
  NAND U9018 ( .A(init), .B(round_reg[324]), .Z(n3316) );
  NANDN U9019 ( .A(init), .B(in[324]), .Z(n3315) );
  NAND U9020 ( .A(n3316), .B(n3315), .Z(\round_in[0][324] ) );
  NAND U9021 ( .A(init), .B(round_reg[325]), .Z(n3318) );
  NANDN U9022 ( .A(init), .B(in[325]), .Z(n3317) );
  NAND U9023 ( .A(n3318), .B(n3317), .Z(\round_in[0][325] ) );
  NAND U9024 ( .A(init), .B(round_reg[326]), .Z(n3320) );
  NANDN U9025 ( .A(init), .B(in[326]), .Z(n3319) );
  NAND U9026 ( .A(n3320), .B(n3319), .Z(\round_in[0][326] ) );
  NAND U9027 ( .A(init), .B(round_reg[327]), .Z(n3322) );
  NANDN U9028 ( .A(init), .B(in[327]), .Z(n3321) );
  NAND U9029 ( .A(n3322), .B(n3321), .Z(\round_in[0][327] ) );
  NAND U9030 ( .A(init), .B(round_reg[328]), .Z(n3324) );
  NANDN U9031 ( .A(init), .B(in[328]), .Z(n3323) );
  NAND U9032 ( .A(n3324), .B(n3323), .Z(\round_in[0][328] ) );
  NAND U9033 ( .A(init), .B(round_reg[329]), .Z(n3326) );
  NANDN U9034 ( .A(init), .B(in[329]), .Z(n3325) );
  NAND U9035 ( .A(n3326), .B(n3325), .Z(\round_in[0][329] ) );
  NAND U9036 ( .A(init), .B(round_reg[32]), .Z(n3328) );
  NANDN U9037 ( .A(init), .B(in[32]), .Z(n3327) );
  NAND U9038 ( .A(n3328), .B(n3327), .Z(\round_in[0][32] ) );
  NAND U9039 ( .A(init), .B(round_reg[330]), .Z(n3330) );
  NANDN U9040 ( .A(init), .B(in[330]), .Z(n3329) );
  NAND U9041 ( .A(n3330), .B(n3329), .Z(\round_in[0][330] ) );
  NAND U9042 ( .A(init), .B(round_reg[331]), .Z(n3332) );
  NANDN U9043 ( .A(init), .B(in[331]), .Z(n3331) );
  NAND U9044 ( .A(n3332), .B(n3331), .Z(\round_in[0][331] ) );
  NAND U9045 ( .A(init), .B(round_reg[332]), .Z(n3334) );
  NANDN U9046 ( .A(init), .B(in[332]), .Z(n3333) );
  NAND U9047 ( .A(n3334), .B(n3333), .Z(\round_in[0][332] ) );
  NAND U9048 ( .A(init), .B(round_reg[333]), .Z(n3336) );
  NANDN U9049 ( .A(init), .B(in[333]), .Z(n3335) );
  NAND U9050 ( .A(n3336), .B(n3335), .Z(\round_in[0][333] ) );
  NAND U9051 ( .A(init), .B(round_reg[334]), .Z(n3338) );
  NANDN U9052 ( .A(init), .B(in[334]), .Z(n3337) );
  NAND U9053 ( .A(n3338), .B(n3337), .Z(\round_in[0][334] ) );
  NAND U9054 ( .A(init), .B(round_reg[335]), .Z(n3340) );
  NANDN U9055 ( .A(init), .B(in[335]), .Z(n3339) );
  NAND U9056 ( .A(n3340), .B(n3339), .Z(\round_in[0][335] ) );
  NAND U9057 ( .A(init), .B(round_reg[336]), .Z(n3342) );
  NANDN U9058 ( .A(init), .B(in[336]), .Z(n3341) );
  NAND U9059 ( .A(n3342), .B(n3341), .Z(\round_in[0][336] ) );
  NAND U9060 ( .A(init), .B(round_reg[337]), .Z(n3344) );
  NANDN U9061 ( .A(init), .B(in[337]), .Z(n3343) );
  NAND U9062 ( .A(n3344), .B(n3343), .Z(\round_in[0][337] ) );
  NAND U9063 ( .A(init), .B(round_reg[338]), .Z(n3346) );
  NANDN U9064 ( .A(init), .B(in[338]), .Z(n3345) );
  NAND U9065 ( .A(n3346), .B(n3345), .Z(\round_in[0][338] ) );
  NAND U9066 ( .A(init), .B(round_reg[339]), .Z(n3348) );
  NANDN U9067 ( .A(init), .B(in[339]), .Z(n3347) );
  NAND U9068 ( .A(n3348), .B(n3347), .Z(\round_in[0][339] ) );
  NAND U9069 ( .A(init), .B(round_reg[33]), .Z(n3350) );
  NANDN U9070 ( .A(init), .B(in[33]), .Z(n3349) );
  NAND U9071 ( .A(n3350), .B(n3349), .Z(\round_in[0][33] ) );
  NAND U9072 ( .A(init), .B(round_reg[340]), .Z(n3352) );
  NANDN U9073 ( .A(init), .B(in[340]), .Z(n3351) );
  NAND U9074 ( .A(n3352), .B(n3351), .Z(\round_in[0][340] ) );
  NAND U9075 ( .A(init), .B(round_reg[341]), .Z(n3354) );
  NANDN U9076 ( .A(init), .B(in[341]), .Z(n3353) );
  NAND U9077 ( .A(n3354), .B(n3353), .Z(\round_in[0][341] ) );
  NAND U9078 ( .A(init), .B(round_reg[342]), .Z(n3356) );
  NANDN U9079 ( .A(init), .B(in[342]), .Z(n3355) );
  NAND U9080 ( .A(n3356), .B(n3355), .Z(\round_in[0][342] ) );
  NAND U9081 ( .A(init), .B(round_reg[343]), .Z(n3358) );
  NANDN U9082 ( .A(init), .B(in[343]), .Z(n3357) );
  NAND U9083 ( .A(n3358), .B(n3357), .Z(\round_in[0][343] ) );
  NAND U9084 ( .A(init), .B(round_reg[344]), .Z(n3360) );
  NANDN U9085 ( .A(init), .B(in[344]), .Z(n3359) );
  NAND U9086 ( .A(n3360), .B(n3359), .Z(\round_in[0][344] ) );
  NAND U9087 ( .A(init), .B(round_reg[345]), .Z(n3362) );
  NANDN U9088 ( .A(init), .B(in[345]), .Z(n3361) );
  NAND U9089 ( .A(n3362), .B(n3361), .Z(\round_in[0][345] ) );
  NAND U9090 ( .A(init), .B(round_reg[346]), .Z(n3364) );
  NANDN U9091 ( .A(init), .B(in[346]), .Z(n3363) );
  NAND U9092 ( .A(n3364), .B(n3363), .Z(\round_in[0][346] ) );
  NAND U9093 ( .A(init), .B(round_reg[347]), .Z(n3366) );
  NANDN U9094 ( .A(init), .B(in[347]), .Z(n3365) );
  NAND U9095 ( .A(n3366), .B(n3365), .Z(\round_in[0][347] ) );
  NAND U9096 ( .A(init), .B(round_reg[348]), .Z(n3368) );
  NANDN U9097 ( .A(init), .B(in[348]), .Z(n3367) );
  NAND U9098 ( .A(n3368), .B(n3367), .Z(\round_in[0][348] ) );
  NAND U9099 ( .A(init), .B(round_reg[349]), .Z(n3370) );
  NANDN U9100 ( .A(init), .B(in[349]), .Z(n3369) );
  NAND U9101 ( .A(n3370), .B(n3369), .Z(\round_in[0][349] ) );
  NAND U9102 ( .A(init), .B(round_reg[34]), .Z(n3372) );
  NANDN U9103 ( .A(init), .B(in[34]), .Z(n3371) );
  NAND U9104 ( .A(n3372), .B(n3371), .Z(\round_in[0][34] ) );
  NAND U9105 ( .A(init), .B(round_reg[350]), .Z(n3374) );
  NANDN U9106 ( .A(init), .B(in[350]), .Z(n3373) );
  NAND U9107 ( .A(n3374), .B(n3373), .Z(\round_in[0][350] ) );
  NAND U9108 ( .A(init), .B(round_reg[351]), .Z(n3376) );
  NANDN U9109 ( .A(init), .B(in[351]), .Z(n3375) );
  NAND U9110 ( .A(n3376), .B(n3375), .Z(\round_in[0][351] ) );
  NAND U9111 ( .A(init), .B(round_reg[352]), .Z(n3378) );
  NANDN U9112 ( .A(init), .B(in[352]), .Z(n3377) );
  NAND U9113 ( .A(n3378), .B(n3377), .Z(\round_in[0][352] ) );
  NAND U9114 ( .A(init), .B(round_reg[353]), .Z(n3380) );
  NANDN U9115 ( .A(init), .B(in[353]), .Z(n3379) );
  NAND U9116 ( .A(n3380), .B(n3379), .Z(\round_in[0][353] ) );
  NAND U9117 ( .A(init), .B(round_reg[354]), .Z(n3382) );
  NANDN U9118 ( .A(init), .B(in[354]), .Z(n3381) );
  NAND U9119 ( .A(n3382), .B(n3381), .Z(\round_in[0][354] ) );
  NAND U9120 ( .A(init), .B(round_reg[355]), .Z(n3384) );
  NANDN U9121 ( .A(init), .B(in[355]), .Z(n3383) );
  NAND U9122 ( .A(n3384), .B(n3383), .Z(\round_in[0][355] ) );
  NAND U9123 ( .A(init), .B(round_reg[356]), .Z(n3386) );
  NANDN U9124 ( .A(init), .B(in[356]), .Z(n3385) );
  NAND U9125 ( .A(n3386), .B(n3385), .Z(\round_in[0][356] ) );
  NAND U9126 ( .A(init), .B(round_reg[357]), .Z(n3388) );
  NANDN U9127 ( .A(init), .B(in[357]), .Z(n3387) );
  NAND U9128 ( .A(n3388), .B(n3387), .Z(\round_in[0][357] ) );
  NAND U9129 ( .A(init), .B(round_reg[358]), .Z(n3390) );
  NANDN U9130 ( .A(init), .B(in[358]), .Z(n3389) );
  NAND U9131 ( .A(n3390), .B(n3389), .Z(\round_in[0][358] ) );
  NAND U9132 ( .A(init), .B(round_reg[359]), .Z(n3392) );
  NANDN U9133 ( .A(init), .B(in[359]), .Z(n3391) );
  NAND U9134 ( .A(n3392), .B(n3391), .Z(\round_in[0][359] ) );
  NAND U9135 ( .A(init), .B(round_reg[35]), .Z(n3394) );
  NANDN U9136 ( .A(init), .B(in[35]), .Z(n3393) );
  NAND U9137 ( .A(n3394), .B(n3393), .Z(\round_in[0][35] ) );
  NAND U9138 ( .A(init), .B(round_reg[360]), .Z(n3396) );
  NANDN U9139 ( .A(init), .B(in[360]), .Z(n3395) );
  NAND U9140 ( .A(n3396), .B(n3395), .Z(\round_in[0][360] ) );
  NAND U9141 ( .A(init), .B(round_reg[361]), .Z(n3398) );
  NANDN U9142 ( .A(init), .B(in[361]), .Z(n3397) );
  NAND U9143 ( .A(n3398), .B(n3397), .Z(\round_in[0][361] ) );
  NAND U9144 ( .A(init), .B(round_reg[362]), .Z(n3400) );
  NANDN U9145 ( .A(init), .B(in[362]), .Z(n3399) );
  NAND U9146 ( .A(n3400), .B(n3399), .Z(\round_in[0][362] ) );
  NAND U9147 ( .A(init), .B(round_reg[363]), .Z(n3402) );
  NANDN U9148 ( .A(init), .B(in[363]), .Z(n3401) );
  NAND U9149 ( .A(n3402), .B(n3401), .Z(\round_in[0][363] ) );
  NAND U9150 ( .A(init), .B(round_reg[364]), .Z(n3404) );
  NANDN U9151 ( .A(init), .B(in[364]), .Z(n3403) );
  NAND U9152 ( .A(n3404), .B(n3403), .Z(\round_in[0][364] ) );
  NAND U9153 ( .A(init), .B(round_reg[365]), .Z(n3406) );
  NANDN U9154 ( .A(init), .B(in[365]), .Z(n3405) );
  NAND U9155 ( .A(n3406), .B(n3405), .Z(\round_in[0][365] ) );
  NAND U9156 ( .A(init), .B(round_reg[366]), .Z(n3408) );
  NANDN U9157 ( .A(init), .B(in[366]), .Z(n3407) );
  NAND U9158 ( .A(n3408), .B(n3407), .Z(\round_in[0][366] ) );
  NAND U9159 ( .A(init), .B(round_reg[367]), .Z(n3410) );
  NANDN U9160 ( .A(init), .B(in[367]), .Z(n3409) );
  NAND U9161 ( .A(n3410), .B(n3409), .Z(\round_in[0][367] ) );
  NAND U9162 ( .A(init), .B(round_reg[368]), .Z(n3412) );
  NANDN U9163 ( .A(init), .B(in[368]), .Z(n3411) );
  NAND U9164 ( .A(n3412), .B(n3411), .Z(\round_in[0][368] ) );
  NAND U9165 ( .A(init), .B(round_reg[369]), .Z(n3414) );
  NANDN U9166 ( .A(init), .B(in[369]), .Z(n3413) );
  NAND U9167 ( .A(n3414), .B(n3413), .Z(\round_in[0][369] ) );
  NAND U9168 ( .A(init), .B(round_reg[36]), .Z(n3416) );
  NANDN U9169 ( .A(init), .B(in[36]), .Z(n3415) );
  NAND U9170 ( .A(n3416), .B(n3415), .Z(\round_in[0][36] ) );
  NAND U9171 ( .A(init), .B(round_reg[370]), .Z(n3418) );
  NANDN U9172 ( .A(init), .B(in[370]), .Z(n3417) );
  NAND U9173 ( .A(n3418), .B(n3417), .Z(\round_in[0][370] ) );
  NAND U9174 ( .A(init), .B(round_reg[371]), .Z(n3420) );
  NANDN U9175 ( .A(init), .B(in[371]), .Z(n3419) );
  NAND U9176 ( .A(n3420), .B(n3419), .Z(\round_in[0][371] ) );
  NAND U9177 ( .A(init), .B(round_reg[372]), .Z(n3422) );
  NANDN U9178 ( .A(init), .B(in[372]), .Z(n3421) );
  NAND U9179 ( .A(n3422), .B(n3421), .Z(\round_in[0][372] ) );
  NAND U9180 ( .A(init), .B(round_reg[373]), .Z(n3424) );
  NANDN U9181 ( .A(init), .B(in[373]), .Z(n3423) );
  NAND U9182 ( .A(n3424), .B(n3423), .Z(\round_in[0][373] ) );
  NAND U9183 ( .A(init), .B(round_reg[374]), .Z(n3426) );
  NANDN U9184 ( .A(init), .B(in[374]), .Z(n3425) );
  NAND U9185 ( .A(n3426), .B(n3425), .Z(\round_in[0][374] ) );
  NAND U9186 ( .A(init), .B(round_reg[375]), .Z(n3428) );
  NANDN U9187 ( .A(init), .B(in[375]), .Z(n3427) );
  NAND U9188 ( .A(n3428), .B(n3427), .Z(\round_in[0][375] ) );
  NAND U9189 ( .A(init), .B(round_reg[376]), .Z(n3430) );
  NANDN U9190 ( .A(init), .B(in[376]), .Z(n3429) );
  NAND U9191 ( .A(n3430), .B(n3429), .Z(\round_in[0][376] ) );
  NAND U9192 ( .A(init), .B(round_reg[377]), .Z(n3432) );
  NANDN U9193 ( .A(init), .B(in[377]), .Z(n3431) );
  NAND U9194 ( .A(n3432), .B(n3431), .Z(\round_in[0][377] ) );
  NAND U9195 ( .A(init), .B(round_reg[378]), .Z(n3434) );
  NANDN U9196 ( .A(init), .B(in[378]), .Z(n3433) );
  NAND U9197 ( .A(n3434), .B(n3433), .Z(\round_in[0][378] ) );
  NAND U9198 ( .A(init), .B(round_reg[379]), .Z(n3436) );
  NANDN U9199 ( .A(init), .B(in[379]), .Z(n3435) );
  NAND U9200 ( .A(n3436), .B(n3435), .Z(\round_in[0][379] ) );
  NAND U9201 ( .A(init), .B(round_reg[37]), .Z(n3438) );
  NANDN U9202 ( .A(init), .B(in[37]), .Z(n3437) );
  NAND U9203 ( .A(n3438), .B(n3437), .Z(\round_in[0][37] ) );
  NAND U9204 ( .A(init), .B(round_reg[380]), .Z(n3440) );
  NANDN U9205 ( .A(init), .B(in[380]), .Z(n3439) );
  NAND U9206 ( .A(n3440), .B(n3439), .Z(\round_in[0][380] ) );
  NAND U9207 ( .A(init), .B(round_reg[381]), .Z(n3442) );
  NANDN U9208 ( .A(init), .B(in[381]), .Z(n3441) );
  NAND U9209 ( .A(n3442), .B(n3441), .Z(\round_in[0][381] ) );
  NAND U9210 ( .A(init), .B(round_reg[382]), .Z(n3444) );
  NANDN U9211 ( .A(init), .B(in[382]), .Z(n3443) );
  NAND U9212 ( .A(n3444), .B(n3443), .Z(\round_in[0][382] ) );
  NAND U9213 ( .A(init), .B(round_reg[383]), .Z(n3446) );
  NANDN U9214 ( .A(init), .B(in[383]), .Z(n3445) );
  NAND U9215 ( .A(n3446), .B(n3445), .Z(\round_in[0][383] ) );
  NAND U9216 ( .A(init), .B(round_reg[384]), .Z(n3448) );
  NANDN U9217 ( .A(init), .B(in[384]), .Z(n3447) );
  NAND U9218 ( .A(n3448), .B(n3447), .Z(\round_in[0][384] ) );
  NAND U9219 ( .A(init), .B(round_reg[385]), .Z(n3450) );
  NANDN U9220 ( .A(init), .B(in[385]), .Z(n3449) );
  NAND U9221 ( .A(n3450), .B(n3449), .Z(\round_in[0][385] ) );
  NAND U9222 ( .A(init), .B(round_reg[386]), .Z(n3452) );
  NANDN U9223 ( .A(init), .B(in[386]), .Z(n3451) );
  NAND U9224 ( .A(n3452), .B(n3451), .Z(\round_in[0][386] ) );
  NAND U9225 ( .A(init), .B(round_reg[387]), .Z(n3454) );
  NANDN U9226 ( .A(init), .B(in[387]), .Z(n3453) );
  NAND U9227 ( .A(n3454), .B(n3453), .Z(\round_in[0][387] ) );
  NAND U9228 ( .A(init), .B(round_reg[388]), .Z(n3456) );
  NANDN U9229 ( .A(init), .B(in[388]), .Z(n3455) );
  NAND U9230 ( .A(n3456), .B(n3455), .Z(\round_in[0][388] ) );
  NAND U9231 ( .A(init), .B(round_reg[389]), .Z(n3458) );
  NANDN U9232 ( .A(init), .B(in[389]), .Z(n3457) );
  NAND U9233 ( .A(n3458), .B(n3457), .Z(\round_in[0][389] ) );
  NAND U9234 ( .A(init), .B(round_reg[38]), .Z(n3460) );
  NANDN U9235 ( .A(init), .B(in[38]), .Z(n3459) );
  NAND U9236 ( .A(n3460), .B(n3459), .Z(\round_in[0][38] ) );
  NAND U9237 ( .A(init), .B(round_reg[390]), .Z(n3462) );
  NANDN U9238 ( .A(init), .B(in[390]), .Z(n3461) );
  NAND U9239 ( .A(n3462), .B(n3461), .Z(\round_in[0][390] ) );
  NAND U9240 ( .A(init), .B(round_reg[391]), .Z(n3464) );
  NANDN U9241 ( .A(init), .B(in[391]), .Z(n3463) );
  NAND U9242 ( .A(n3464), .B(n3463), .Z(\round_in[0][391] ) );
  NAND U9243 ( .A(init), .B(round_reg[392]), .Z(n3466) );
  NANDN U9244 ( .A(init), .B(in[392]), .Z(n3465) );
  NAND U9245 ( .A(n3466), .B(n3465), .Z(\round_in[0][392] ) );
  NAND U9246 ( .A(init), .B(round_reg[393]), .Z(n3468) );
  NANDN U9247 ( .A(init), .B(in[393]), .Z(n3467) );
  NAND U9248 ( .A(n3468), .B(n3467), .Z(\round_in[0][393] ) );
  NAND U9249 ( .A(init), .B(round_reg[394]), .Z(n3470) );
  NANDN U9250 ( .A(init), .B(in[394]), .Z(n3469) );
  NAND U9251 ( .A(n3470), .B(n3469), .Z(\round_in[0][394] ) );
  NAND U9252 ( .A(init), .B(round_reg[395]), .Z(n3472) );
  NANDN U9253 ( .A(init), .B(in[395]), .Z(n3471) );
  NAND U9254 ( .A(n3472), .B(n3471), .Z(\round_in[0][395] ) );
  NAND U9255 ( .A(init), .B(round_reg[396]), .Z(n3474) );
  NANDN U9256 ( .A(init), .B(in[396]), .Z(n3473) );
  NAND U9257 ( .A(n3474), .B(n3473), .Z(\round_in[0][396] ) );
  NAND U9258 ( .A(init), .B(round_reg[397]), .Z(n3476) );
  NANDN U9259 ( .A(init), .B(in[397]), .Z(n3475) );
  NAND U9260 ( .A(n3476), .B(n3475), .Z(\round_in[0][397] ) );
  NAND U9261 ( .A(init), .B(round_reg[398]), .Z(n3478) );
  NANDN U9262 ( .A(init), .B(in[398]), .Z(n3477) );
  NAND U9263 ( .A(n3478), .B(n3477), .Z(\round_in[0][398] ) );
  NAND U9264 ( .A(init), .B(round_reg[399]), .Z(n3480) );
  NANDN U9265 ( .A(init), .B(in[399]), .Z(n3479) );
  NAND U9266 ( .A(n3480), .B(n3479), .Z(\round_in[0][399] ) );
  NAND U9267 ( .A(init), .B(round_reg[39]), .Z(n3482) );
  NANDN U9268 ( .A(init), .B(in[39]), .Z(n3481) );
  NAND U9269 ( .A(n3482), .B(n3481), .Z(\round_in[0][39] ) );
  NAND U9270 ( .A(init), .B(round_reg[3]), .Z(n3484) );
  NANDN U9271 ( .A(init), .B(in[3]), .Z(n3483) );
  NAND U9272 ( .A(n3484), .B(n3483), .Z(\round_in[0][3] ) );
  NAND U9273 ( .A(init), .B(round_reg[400]), .Z(n3486) );
  NANDN U9274 ( .A(init), .B(in[400]), .Z(n3485) );
  NAND U9275 ( .A(n3486), .B(n3485), .Z(\round_in[0][400] ) );
  NAND U9276 ( .A(init), .B(round_reg[401]), .Z(n3488) );
  NANDN U9277 ( .A(init), .B(in[401]), .Z(n3487) );
  NAND U9278 ( .A(n3488), .B(n3487), .Z(\round_in[0][401] ) );
  NAND U9279 ( .A(init), .B(round_reg[402]), .Z(n3490) );
  NANDN U9280 ( .A(init), .B(in[402]), .Z(n3489) );
  NAND U9281 ( .A(n3490), .B(n3489), .Z(\round_in[0][402] ) );
  NAND U9282 ( .A(init), .B(round_reg[403]), .Z(n3492) );
  NANDN U9283 ( .A(init), .B(in[403]), .Z(n3491) );
  NAND U9284 ( .A(n3492), .B(n3491), .Z(\round_in[0][403] ) );
  NAND U9285 ( .A(init), .B(round_reg[404]), .Z(n3494) );
  NANDN U9286 ( .A(init), .B(in[404]), .Z(n3493) );
  NAND U9287 ( .A(n3494), .B(n3493), .Z(\round_in[0][404] ) );
  NAND U9288 ( .A(init), .B(round_reg[405]), .Z(n3496) );
  NANDN U9289 ( .A(init), .B(in[405]), .Z(n3495) );
  NAND U9290 ( .A(n3496), .B(n3495), .Z(\round_in[0][405] ) );
  NAND U9291 ( .A(init), .B(round_reg[406]), .Z(n3498) );
  NANDN U9292 ( .A(init), .B(in[406]), .Z(n3497) );
  NAND U9293 ( .A(n3498), .B(n3497), .Z(\round_in[0][406] ) );
  NAND U9294 ( .A(init), .B(round_reg[407]), .Z(n3500) );
  NANDN U9295 ( .A(init), .B(in[407]), .Z(n3499) );
  NAND U9296 ( .A(n3500), .B(n3499), .Z(\round_in[0][407] ) );
  NAND U9297 ( .A(init), .B(round_reg[408]), .Z(n3502) );
  NANDN U9298 ( .A(init), .B(in[408]), .Z(n3501) );
  NAND U9299 ( .A(n3502), .B(n3501), .Z(\round_in[0][408] ) );
  NAND U9300 ( .A(init), .B(round_reg[409]), .Z(n3504) );
  NANDN U9301 ( .A(init), .B(in[409]), .Z(n3503) );
  NAND U9302 ( .A(n3504), .B(n3503), .Z(\round_in[0][409] ) );
  NAND U9303 ( .A(init), .B(round_reg[40]), .Z(n3506) );
  NANDN U9304 ( .A(init), .B(in[40]), .Z(n3505) );
  NAND U9305 ( .A(n3506), .B(n3505), .Z(\round_in[0][40] ) );
  NAND U9306 ( .A(init), .B(round_reg[410]), .Z(n3508) );
  NANDN U9307 ( .A(init), .B(in[410]), .Z(n3507) );
  NAND U9308 ( .A(n3508), .B(n3507), .Z(\round_in[0][410] ) );
  NAND U9309 ( .A(init), .B(round_reg[411]), .Z(n3510) );
  NANDN U9310 ( .A(init), .B(in[411]), .Z(n3509) );
  NAND U9311 ( .A(n3510), .B(n3509), .Z(\round_in[0][411] ) );
  NAND U9312 ( .A(init), .B(round_reg[412]), .Z(n3512) );
  NANDN U9313 ( .A(init), .B(in[412]), .Z(n3511) );
  NAND U9314 ( .A(n3512), .B(n3511), .Z(\round_in[0][412] ) );
  NAND U9315 ( .A(init), .B(round_reg[413]), .Z(n3514) );
  NANDN U9316 ( .A(init), .B(in[413]), .Z(n3513) );
  NAND U9317 ( .A(n3514), .B(n3513), .Z(\round_in[0][413] ) );
  NAND U9318 ( .A(init), .B(round_reg[414]), .Z(n3516) );
  NANDN U9319 ( .A(init), .B(in[414]), .Z(n3515) );
  NAND U9320 ( .A(n3516), .B(n3515), .Z(\round_in[0][414] ) );
  NAND U9321 ( .A(init), .B(round_reg[415]), .Z(n3518) );
  NANDN U9322 ( .A(init), .B(in[415]), .Z(n3517) );
  NAND U9323 ( .A(n3518), .B(n3517), .Z(\round_in[0][415] ) );
  NAND U9324 ( .A(init), .B(round_reg[416]), .Z(n3520) );
  NANDN U9325 ( .A(init), .B(in[416]), .Z(n3519) );
  NAND U9326 ( .A(n3520), .B(n3519), .Z(\round_in[0][416] ) );
  NAND U9327 ( .A(init), .B(round_reg[417]), .Z(n3522) );
  NANDN U9328 ( .A(init), .B(in[417]), .Z(n3521) );
  NAND U9329 ( .A(n3522), .B(n3521), .Z(\round_in[0][417] ) );
  NAND U9330 ( .A(init), .B(round_reg[418]), .Z(n3524) );
  NANDN U9331 ( .A(init), .B(in[418]), .Z(n3523) );
  NAND U9332 ( .A(n3524), .B(n3523), .Z(\round_in[0][418] ) );
  NAND U9333 ( .A(init), .B(round_reg[419]), .Z(n3526) );
  NANDN U9334 ( .A(init), .B(in[419]), .Z(n3525) );
  NAND U9335 ( .A(n3526), .B(n3525), .Z(\round_in[0][419] ) );
  NAND U9336 ( .A(init), .B(round_reg[41]), .Z(n3528) );
  NANDN U9337 ( .A(init), .B(in[41]), .Z(n3527) );
  NAND U9338 ( .A(n3528), .B(n3527), .Z(\round_in[0][41] ) );
  NAND U9339 ( .A(init), .B(round_reg[420]), .Z(n3530) );
  NANDN U9340 ( .A(init), .B(in[420]), .Z(n3529) );
  NAND U9341 ( .A(n3530), .B(n3529), .Z(\round_in[0][420] ) );
  NAND U9342 ( .A(init), .B(round_reg[421]), .Z(n3532) );
  NANDN U9343 ( .A(init), .B(in[421]), .Z(n3531) );
  NAND U9344 ( .A(n3532), .B(n3531), .Z(\round_in[0][421] ) );
  NAND U9345 ( .A(init), .B(round_reg[422]), .Z(n3534) );
  NANDN U9346 ( .A(init), .B(in[422]), .Z(n3533) );
  NAND U9347 ( .A(n3534), .B(n3533), .Z(\round_in[0][422] ) );
  NAND U9348 ( .A(init), .B(round_reg[423]), .Z(n3536) );
  NANDN U9349 ( .A(init), .B(in[423]), .Z(n3535) );
  NAND U9350 ( .A(n3536), .B(n3535), .Z(\round_in[0][423] ) );
  NAND U9351 ( .A(init), .B(round_reg[424]), .Z(n3538) );
  NANDN U9352 ( .A(init), .B(in[424]), .Z(n3537) );
  NAND U9353 ( .A(n3538), .B(n3537), .Z(\round_in[0][424] ) );
  NAND U9354 ( .A(init), .B(round_reg[425]), .Z(n3540) );
  NANDN U9355 ( .A(init), .B(in[425]), .Z(n3539) );
  NAND U9356 ( .A(n3540), .B(n3539), .Z(\round_in[0][425] ) );
  NAND U9357 ( .A(init), .B(round_reg[426]), .Z(n3542) );
  NANDN U9358 ( .A(init), .B(in[426]), .Z(n3541) );
  NAND U9359 ( .A(n3542), .B(n3541), .Z(\round_in[0][426] ) );
  NAND U9360 ( .A(init), .B(round_reg[427]), .Z(n3544) );
  NANDN U9361 ( .A(init), .B(in[427]), .Z(n3543) );
  NAND U9362 ( .A(n3544), .B(n3543), .Z(\round_in[0][427] ) );
  NAND U9363 ( .A(init), .B(round_reg[428]), .Z(n3546) );
  NANDN U9364 ( .A(init), .B(in[428]), .Z(n3545) );
  NAND U9365 ( .A(n3546), .B(n3545), .Z(\round_in[0][428] ) );
  NAND U9366 ( .A(init), .B(round_reg[429]), .Z(n3548) );
  NANDN U9367 ( .A(init), .B(in[429]), .Z(n3547) );
  NAND U9368 ( .A(n3548), .B(n3547), .Z(\round_in[0][429] ) );
  NAND U9369 ( .A(init), .B(round_reg[42]), .Z(n3550) );
  NANDN U9370 ( .A(init), .B(in[42]), .Z(n3549) );
  NAND U9371 ( .A(n3550), .B(n3549), .Z(\round_in[0][42] ) );
  NAND U9372 ( .A(init), .B(round_reg[430]), .Z(n3552) );
  NANDN U9373 ( .A(init), .B(in[430]), .Z(n3551) );
  NAND U9374 ( .A(n3552), .B(n3551), .Z(\round_in[0][430] ) );
  NAND U9375 ( .A(init), .B(round_reg[431]), .Z(n3554) );
  NANDN U9376 ( .A(init), .B(in[431]), .Z(n3553) );
  NAND U9377 ( .A(n3554), .B(n3553), .Z(\round_in[0][431] ) );
  NAND U9378 ( .A(init), .B(round_reg[432]), .Z(n3556) );
  NANDN U9379 ( .A(init), .B(in[432]), .Z(n3555) );
  NAND U9380 ( .A(n3556), .B(n3555), .Z(\round_in[0][432] ) );
  NAND U9381 ( .A(init), .B(round_reg[433]), .Z(n3558) );
  NANDN U9382 ( .A(init), .B(in[433]), .Z(n3557) );
  NAND U9383 ( .A(n3558), .B(n3557), .Z(\round_in[0][433] ) );
  NAND U9384 ( .A(init), .B(round_reg[434]), .Z(n3560) );
  NANDN U9385 ( .A(init), .B(in[434]), .Z(n3559) );
  NAND U9386 ( .A(n3560), .B(n3559), .Z(\round_in[0][434] ) );
  NAND U9387 ( .A(init), .B(round_reg[435]), .Z(n3562) );
  NANDN U9388 ( .A(init), .B(in[435]), .Z(n3561) );
  NAND U9389 ( .A(n3562), .B(n3561), .Z(\round_in[0][435] ) );
  NAND U9390 ( .A(init), .B(round_reg[436]), .Z(n3564) );
  NANDN U9391 ( .A(init), .B(in[436]), .Z(n3563) );
  NAND U9392 ( .A(n3564), .B(n3563), .Z(\round_in[0][436] ) );
  NAND U9393 ( .A(init), .B(round_reg[437]), .Z(n3566) );
  NANDN U9394 ( .A(init), .B(in[437]), .Z(n3565) );
  NAND U9395 ( .A(n3566), .B(n3565), .Z(\round_in[0][437] ) );
  NAND U9396 ( .A(init), .B(round_reg[438]), .Z(n3568) );
  NANDN U9397 ( .A(init), .B(in[438]), .Z(n3567) );
  NAND U9398 ( .A(n3568), .B(n3567), .Z(\round_in[0][438] ) );
  NAND U9399 ( .A(init), .B(round_reg[439]), .Z(n3570) );
  NANDN U9400 ( .A(init), .B(in[439]), .Z(n3569) );
  NAND U9401 ( .A(n3570), .B(n3569), .Z(\round_in[0][439] ) );
  NAND U9402 ( .A(init), .B(round_reg[43]), .Z(n3572) );
  NANDN U9403 ( .A(init), .B(in[43]), .Z(n3571) );
  NAND U9404 ( .A(n3572), .B(n3571), .Z(\round_in[0][43] ) );
  NAND U9405 ( .A(init), .B(round_reg[440]), .Z(n3574) );
  NANDN U9406 ( .A(init), .B(in[440]), .Z(n3573) );
  NAND U9407 ( .A(n3574), .B(n3573), .Z(\round_in[0][440] ) );
  NAND U9408 ( .A(init), .B(round_reg[441]), .Z(n3576) );
  NANDN U9409 ( .A(init), .B(in[441]), .Z(n3575) );
  NAND U9410 ( .A(n3576), .B(n3575), .Z(\round_in[0][441] ) );
  NAND U9411 ( .A(init), .B(round_reg[442]), .Z(n3578) );
  NANDN U9412 ( .A(init), .B(in[442]), .Z(n3577) );
  NAND U9413 ( .A(n3578), .B(n3577), .Z(\round_in[0][442] ) );
  NAND U9414 ( .A(init), .B(round_reg[443]), .Z(n3580) );
  NANDN U9415 ( .A(init), .B(in[443]), .Z(n3579) );
  NAND U9416 ( .A(n3580), .B(n3579), .Z(\round_in[0][443] ) );
  NAND U9417 ( .A(init), .B(round_reg[444]), .Z(n3582) );
  NANDN U9418 ( .A(init), .B(in[444]), .Z(n3581) );
  NAND U9419 ( .A(n3582), .B(n3581), .Z(\round_in[0][444] ) );
  NAND U9420 ( .A(init), .B(round_reg[445]), .Z(n3584) );
  NANDN U9421 ( .A(init), .B(in[445]), .Z(n3583) );
  NAND U9422 ( .A(n3584), .B(n3583), .Z(\round_in[0][445] ) );
  NAND U9423 ( .A(init), .B(round_reg[446]), .Z(n3586) );
  NANDN U9424 ( .A(init), .B(in[446]), .Z(n3585) );
  NAND U9425 ( .A(n3586), .B(n3585), .Z(\round_in[0][446] ) );
  NAND U9426 ( .A(init), .B(round_reg[447]), .Z(n3588) );
  NANDN U9427 ( .A(init), .B(in[447]), .Z(n3587) );
  NAND U9428 ( .A(n3588), .B(n3587), .Z(\round_in[0][447] ) );
  NAND U9429 ( .A(init), .B(round_reg[448]), .Z(n3590) );
  NANDN U9430 ( .A(init), .B(in[448]), .Z(n3589) );
  NAND U9431 ( .A(n3590), .B(n3589), .Z(\round_in[0][448] ) );
  NAND U9432 ( .A(init), .B(round_reg[449]), .Z(n3592) );
  NANDN U9433 ( .A(init), .B(in[449]), .Z(n3591) );
  NAND U9434 ( .A(n3592), .B(n3591), .Z(\round_in[0][449] ) );
  NAND U9435 ( .A(init), .B(round_reg[44]), .Z(n3594) );
  NANDN U9436 ( .A(init), .B(in[44]), .Z(n3593) );
  NAND U9437 ( .A(n3594), .B(n3593), .Z(\round_in[0][44] ) );
  NAND U9438 ( .A(init), .B(round_reg[450]), .Z(n3596) );
  NANDN U9439 ( .A(init), .B(in[450]), .Z(n3595) );
  NAND U9440 ( .A(n3596), .B(n3595), .Z(\round_in[0][450] ) );
  NAND U9441 ( .A(init), .B(round_reg[451]), .Z(n3598) );
  NANDN U9442 ( .A(init), .B(in[451]), .Z(n3597) );
  NAND U9443 ( .A(n3598), .B(n3597), .Z(\round_in[0][451] ) );
  NAND U9444 ( .A(init), .B(round_reg[452]), .Z(n3600) );
  NANDN U9445 ( .A(init), .B(in[452]), .Z(n3599) );
  NAND U9446 ( .A(n3600), .B(n3599), .Z(\round_in[0][452] ) );
  NAND U9447 ( .A(init), .B(round_reg[453]), .Z(n3602) );
  NANDN U9448 ( .A(init), .B(in[453]), .Z(n3601) );
  NAND U9449 ( .A(n3602), .B(n3601), .Z(\round_in[0][453] ) );
  NAND U9450 ( .A(init), .B(round_reg[454]), .Z(n3604) );
  NANDN U9451 ( .A(init), .B(in[454]), .Z(n3603) );
  NAND U9452 ( .A(n3604), .B(n3603), .Z(\round_in[0][454] ) );
  NAND U9453 ( .A(init), .B(round_reg[455]), .Z(n3606) );
  NANDN U9454 ( .A(init), .B(in[455]), .Z(n3605) );
  NAND U9455 ( .A(n3606), .B(n3605), .Z(\round_in[0][455] ) );
  NAND U9456 ( .A(init), .B(round_reg[456]), .Z(n3608) );
  NANDN U9457 ( .A(init), .B(in[456]), .Z(n3607) );
  NAND U9458 ( .A(n3608), .B(n3607), .Z(\round_in[0][456] ) );
  NAND U9459 ( .A(init), .B(round_reg[457]), .Z(n3610) );
  NANDN U9460 ( .A(init), .B(in[457]), .Z(n3609) );
  NAND U9461 ( .A(n3610), .B(n3609), .Z(\round_in[0][457] ) );
  NAND U9462 ( .A(init), .B(round_reg[458]), .Z(n3612) );
  NANDN U9463 ( .A(init), .B(in[458]), .Z(n3611) );
  NAND U9464 ( .A(n3612), .B(n3611), .Z(\round_in[0][458] ) );
  NAND U9465 ( .A(init), .B(round_reg[459]), .Z(n3614) );
  NANDN U9466 ( .A(init), .B(in[459]), .Z(n3613) );
  NAND U9467 ( .A(n3614), .B(n3613), .Z(\round_in[0][459] ) );
  NAND U9468 ( .A(init), .B(round_reg[45]), .Z(n3616) );
  NANDN U9469 ( .A(init), .B(in[45]), .Z(n3615) );
  NAND U9470 ( .A(n3616), .B(n3615), .Z(\round_in[0][45] ) );
  NAND U9471 ( .A(init), .B(round_reg[460]), .Z(n3618) );
  NANDN U9472 ( .A(init), .B(in[460]), .Z(n3617) );
  NAND U9473 ( .A(n3618), .B(n3617), .Z(\round_in[0][460] ) );
  NAND U9474 ( .A(init), .B(round_reg[461]), .Z(n3620) );
  NANDN U9475 ( .A(init), .B(in[461]), .Z(n3619) );
  NAND U9476 ( .A(n3620), .B(n3619), .Z(\round_in[0][461] ) );
  NAND U9477 ( .A(init), .B(round_reg[462]), .Z(n3622) );
  NANDN U9478 ( .A(init), .B(in[462]), .Z(n3621) );
  NAND U9479 ( .A(n3622), .B(n3621), .Z(\round_in[0][462] ) );
  NAND U9480 ( .A(init), .B(round_reg[463]), .Z(n3624) );
  NANDN U9481 ( .A(init), .B(in[463]), .Z(n3623) );
  NAND U9482 ( .A(n3624), .B(n3623), .Z(\round_in[0][463] ) );
  NAND U9483 ( .A(init), .B(round_reg[464]), .Z(n3626) );
  NANDN U9484 ( .A(init), .B(in[464]), .Z(n3625) );
  NAND U9485 ( .A(n3626), .B(n3625), .Z(\round_in[0][464] ) );
  NAND U9486 ( .A(init), .B(round_reg[465]), .Z(n3628) );
  NANDN U9487 ( .A(init), .B(in[465]), .Z(n3627) );
  NAND U9488 ( .A(n3628), .B(n3627), .Z(\round_in[0][465] ) );
  NAND U9489 ( .A(init), .B(round_reg[466]), .Z(n3630) );
  NANDN U9490 ( .A(init), .B(in[466]), .Z(n3629) );
  NAND U9491 ( .A(n3630), .B(n3629), .Z(\round_in[0][466] ) );
  NAND U9492 ( .A(init), .B(round_reg[467]), .Z(n3632) );
  NANDN U9493 ( .A(init), .B(in[467]), .Z(n3631) );
  NAND U9494 ( .A(n3632), .B(n3631), .Z(\round_in[0][467] ) );
  NAND U9495 ( .A(init), .B(round_reg[468]), .Z(n3634) );
  NANDN U9496 ( .A(init), .B(in[468]), .Z(n3633) );
  NAND U9497 ( .A(n3634), .B(n3633), .Z(\round_in[0][468] ) );
  NAND U9498 ( .A(init), .B(round_reg[469]), .Z(n3636) );
  NANDN U9499 ( .A(init), .B(in[469]), .Z(n3635) );
  NAND U9500 ( .A(n3636), .B(n3635), .Z(\round_in[0][469] ) );
  NAND U9501 ( .A(init), .B(round_reg[46]), .Z(n3638) );
  NANDN U9502 ( .A(init), .B(in[46]), .Z(n3637) );
  NAND U9503 ( .A(n3638), .B(n3637), .Z(\round_in[0][46] ) );
  NAND U9504 ( .A(init), .B(round_reg[470]), .Z(n3640) );
  NANDN U9505 ( .A(init), .B(in[470]), .Z(n3639) );
  NAND U9506 ( .A(n3640), .B(n3639), .Z(\round_in[0][470] ) );
  NAND U9507 ( .A(init), .B(round_reg[471]), .Z(n3642) );
  NANDN U9508 ( .A(init), .B(in[471]), .Z(n3641) );
  NAND U9509 ( .A(n3642), .B(n3641), .Z(\round_in[0][471] ) );
  NAND U9510 ( .A(init), .B(round_reg[472]), .Z(n3644) );
  NANDN U9511 ( .A(init), .B(in[472]), .Z(n3643) );
  NAND U9512 ( .A(n3644), .B(n3643), .Z(\round_in[0][472] ) );
  NAND U9513 ( .A(init), .B(round_reg[473]), .Z(n3646) );
  NANDN U9514 ( .A(init), .B(in[473]), .Z(n3645) );
  NAND U9515 ( .A(n3646), .B(n3645), .Z(\round_in[0][473] ) );
  NAND U9516 ( .A(init), .B(round_reg[474]), .Z(n3648) );
  NANDN U9517 ( .A(init), .B(in[474]), .Z(n3647) );
  NAND U9518 ( .A(n3648), .B(n3647), .Z(\round_in[0][474] ) );
  NAND U9519 ( .A(init), .B(round_reg[475]), .Z(n3650) );
  NANDN U9520 ( .A(init), .B(in[475]), .Z(n3649) );
  NAND U9521 ( .A(n3650), .B(n3649), .Z(\round_in[0][475] ) );
  NAND U9522 ( .A(init), .B(round_reg[476]), .Z(n3652) );
  NANDN U9523 ( .A(init), .B(in[476]), .Z(n3651) );
  NAND U9524 ( .A(n3652), .B(n3651), .Z(\round_in[0][476] ) );
  NAND U9525 ( .A(init), .B(round_reg[477]), .Z(n3654) );
  NANDN U9526 ( .A(init), .B(in[477]), .Z(n3653) );
  NAND U9527 ( .A(n3654), .B(n3653), .Z(\round_in[0][477] ) );
  NAND U9528 ( .A(init), .B(round_reg[478]), .Z(n3656) );
  NANDN U9529 ( .A(init), .B(in[478]), .Z(n3655) );
  NAND U9530 ( .A(n3656), .B(n3655), .Z(\round_in[0][478] ) );
  NAND U9531 ( .A(init), .B(round_reg[479]), .Z(n3658) );
  NANDN U9532 ( .A(init), .B(in[479]), .Z(n3657) );
  NAND U9533 ( .A(n3658), .B(n3657), .Z(\round_in[0][479] ) );
  NAND U9534 ( .A(init), .B(round_reg[47]), .Z(n3660) );
  NANDN U9535 ( .A(init), .B(in[47]), .Z(n3659) );
  NAND U9536 ( .A(n3660), .B(n3659), .Z(\round_in[0][47] ) );
  NAND U9537 ( .A(init), .B(round_reg[480]), .Z(n3662) );
  NANDN U9538 ( .A(init), .B(in[480]), .Z(n3661) );
  NAND U9539 ( .A(n3662), .B(n3661), .Z(\round_in[0][480] ) );
  NAND U9540 ( .A(init), .B(round_reg[481]), .Z(n3664) );
  NANDN U9541 ( .A(init), .B(in[481]), .Z(n3663) );
  NAND U9542 ( .A(n3664), .B(n3663), .Z(\round_in[0][481] ) );
  NAND U9543 ( .A(init), .B(round_reg[482]), .Z(n3666) );
  NANDN U9544 ( .A(init), .B(in[482]), .Z(n3665) );
  NAND U9545 ( .A(n3666), .B(n3665), .Z(\round_in[0][482] ) );
  NAND U9546 ( .A(init), .B(round_reg[483]), .Z(n3668) );
  NANDN U9547 ( .A(init), .B(in[483]), .Z(n3667) );
  NAND U9548 ( .A(n3668), .B(n3667), .Z(\round_in[0][483] ) );
  NAND U9549 ( .A(init), .B(round_reg[484]), .Z(n3670) );
  NANDN U9550 ( .A(init), .B(in[484]), .Z(n3669) );
  NAND U9551 ( .A(n3670), .B(n3669), .Z(\round_in[0][484] ) );
  NAND U9552 ( .A(init), .B(round_reg[485]), .Z(n3672) );
  NANDN U9553 ( .A(init), .B(in[485]), .Z(n3671) );
  NAND U9554 ( .A(n3672), .B(n3671), .Z(\round_in[0][485] ) );
  NAND U9555 ( .A(init), .B(round_reg[486]), .Z(n3674) );
  NANDN U9556 ( .A(init), .B(in[486]), .Z(n3673) );
  NAND U9557 ( .A(n3674), .B(n3673), .Z(\round_in[0][486] ) );
  NAND U9558 ( .A(init), .B(round_reg[487]), .Z(n3676) );
  NANDN U9559 ( .A(init), .B(in[487]), .Z(n3675) );
  NAND U9560 ( .A(n3676), .B(n3675), .Z(\round_in[0][487] ) );
  NAND U9561 ( .A(init), .B(round_reg[488]), .Z(n3678) );
  NANDN U9562 ( .A(init), .B(in[488]), .Z(n3677) );
  NAND U9563 ( .A(n3678), .B(n3677), .Z(\round_in[0][488] ) );
  NAND U9564 ( .A(init), .B(round_reg[489]), .Z(n3680) );
  NANDN U9565 ( .A(init), .B(in[489]), .Z(n3679) );
  NAND U9566 ( .A(n3680), .B(n3679), .Z(\round_in[0][489] ) );
  NAND U9567 ( .A(init), .B(round_reg[48]), .Z(n3682) );
  NANDN U9568 ( .A(init), .B(in[48]), .Z(n3681) );
  NAND U9569 ( .A(n3682), .B(n3681), .Z(\round_in[0][48] ) );
  NAND U9570 ( .A(init), .B(round_reg[490]), .Z(n3684) );
  NANDN U9571 ( .A(init), .B(in[490]), .Z(n3683) );
  NAND U9572 ( .A(n3684), .B(n3683), .Z(\round_in[0][490] ) );
  NAND U9573 ( .A(init), .B(round_reg[491]), .Z(n3686) );
  NANDN U9574 ( .A(init), .B(in[491]), .Z(n3685) );
  NAND U9575 ( .A(n3686), .B(n3685), .Z(\round_in[0][491] ) );
  NAND U9576 ( .A(init), .B(round_reg[492]), .Z(n3688) );
  NANDN U9577 ( .A(init), .B(in[492]), .Z(n3687) );
  NAND U9578 ( .A(n3688), .B(n3687), .Z(\round_in[0][492] ) );
  NAND U9579 ( .A(init), .B(round_reg[493]), .Z(n3690) );
  NANDN U9580 ( .A(init), .B(in[493]), .Z(n3689) );
  NAND U9581 ( .A(n3690), .B(n3689), .Z(\round_in[0][493] ) );
  NAND U9582 ( .A(init), .B(round_reg[494]), .Z(n3692) );
  NANDN U9583 ( .A(init), .B(in[494]), .Z(n3691) );
  NAND U9584 ( .A(n3692), .B(n3691), .Z(\round_in[0][494] ) );
  NAND U9585 ( .A(init), .B(round_reg[495]), .Z(n3694) );
  NANDN U9586 ( .A(init), .B(in[495]), .Z(n3693) );
  NAND U9587 ( .A(n3694), .B(n3693), .Z(\round_in[0][495] ) );
  NAND U9588 ( .A(init), .B(round_reg[496]), .Z(n3696) );
  NANDN U9589 ( .A(init), .B(in[496]), .Z(n3695) );
  NAND U9590 ( .A(n3696), .B(n3695), .Z(\round_in[0][496] ) );
  NAND U9591 ( .A(init), .B(round_reg[497]), .Z(n3698) );
  NANDN U9592 ( .A(init), .B(in[497]), .Z(n3697) );
  NAND U9593 ( .A(n3698), .B(n3697), .Z(\round_in[0][497] ) );
  NAND U9594 ( .A(init), .B(round_reg[498]), .Z(n3700) );
  NANDN U9595 ( .A(init), .B(in[498]), .Z(n3699) );
  NAND U9596 ( .A(n3700), .B(n3699), .Z(\round_in[0][498] ) );
  NAND U9597 ( .A(init), .B(round_reg[499]), .Z(n3702) );
  NANDN U9598 ( .A(init), .B(in[499]), .Z(n3701) );
  NAND U9599 ( .A(n3702), .B(n3701), .Z(\round_in[0][499] ) );
  NAND U9600 ( .A(init), .B(round_reg[49]), .Z(n3704) );
  NANDN U9601 ( .A(init), .B(in[49]), .Z(n3703) );
  NAND U9602 ( .A(n3704), .B(n3703), .Z(\round_in[0][49] ) );
  NAND U9603 ( .A(init), .B(round_reg[4]), .Z(n3706) );
  NANDN U9604 ( .A(init), .B(in[4]), .Z(n3705) );
  NAND U9605 ( .A(n3706), .B(n3705), .Z(\round_in[0][4] ) );
  NAND U9606 ( .A(init), .B(round_reg[500]), .Z(n3708) );
  NANDN U9607 ( .A(init), .B(in[500]), .Z(n3707) );
  NAND U9608 ( .A(n3708), .B(n3707), .Z(\round_in[0][500] ) );
  NAND U9609 ( .A(init), .B(round_reg[501]), .Z(n3710) );
  NANDN U9610 ( .A(init), .B(in[501]), .Z(n3709) );
  NAND U9611 ( .A(n3710), .B(n3709), .Z(\round_in[0][501] ) );
  NAND U9612 ( .A(init), .B(round_reg[502]), .Z(n3712) );
  NANDN U9613 ( .A(init), .B(in[502]), .Z(n3711) );
  NAND U9614 ( .A(n3712), .B(n3711), .Z(\round_in[0][502] ) );
  NAND U9615 ( .A(init), .B(round_reg[503]), .Z(n3714) );
  NANDN U9616 ( .A(init), .B(in[503]), .Z(n3713) );
  NAND U9617 ( .A(n3714), .B(n3713), .Z(\round_in[0][503] ) );
  NAND U9618 ( .A(init), .B(round_reg[504]), .Z(n3716) );
  NANDN U9619 ( .A(init), .B(in[504]), .Z(n3715) );
  NAND U9620 ( .A(n3716), .B(n3715), .Z(\round_in[0][504] ) );
  NAND U9621 ( .A(init), .B(round_reg[505]), .Z(n3718) );
  NANDN U9622 ( .A(init), .B(in[505]), .Z(n3717) );
  NAND U9623 ( .A(n3718), .B(n3717), .Z(\round_in[0][505] ) );
  NAND U9624 ( .A(init), .B(round_reg[506]), .Z(n3720) );
  NANDN U9625 ( .A(init), .B(in[506]), .Z(n3719) );
  NAND U9626 ( .A(n3720), .B(n3719), .Z(\round_in[0][506] ) );
  NAND U9627 ( .A(init), .B(round_reg[507]), .Z(n3722) );
  NANDN U9628 ( .A(init), .B(in[507]), .Z(n3721) );
  NAND U9629 ( .A(n3722), .B(n3721), .Z(\round_in[0][507] ) );
  NAND U9630 ( .A(init), .B(round_reg[508]), .Z(n3724) );
  NANDN U9631 ( .A(init), .B(in[508]), .Z(n3723) );
  NAND U9632 ( .A(n3724), .B(n3723), .Z(\round_in[0][508] ) );
  NAND U9633 ( .A(init), .B(round_reg[509]), .Z(n3726) );
  NANDN U9634 ( .A(init), .B(in[509]), .Z(n3725) );
  NAND U9635 ( .A(n3726), .B(n3725), .Z(\round_in[0][509] ) );
  NAND U9636 ( .A(init), .B(round_reg[50]), .Z(n3728) );
  NANDN U9637 ( .A(init), .B(in[50]), .Z(n3727) );
  NAND U9638 ( .A(n3728), .B(n3727), .Z(\round_in[0][50] ) );
  NAND U9639 ( .A(init), .B(round_reg[510]), .Z(n3730) );
  NANDN U9640 ( .A(init), .B(in[510]), .Z(n3729) );
  NAND U9641 ( .A(n3730), .B(n3729), .Z(\round_in[0][510] ) );
  NAND U9642 ( .A(init), .B(round_reg[511]), .Z(n3732) );
  NANDN U9643 ( .A(init), .B(in[511]), .Z(n3731) );
  NAND U9644 ( .A(n3732), .B(n3731), .Z(\round_in[0][511] ) );
  NAND U9645 ( .A(init), .B(round_reg[512]), .Z(n3734) );
  NANDN U9646 ( .A(init), .B(in[512]), .Z(n3733) );
  NAND U9647 ( .A(n3734), .B(n3733), .Z(\round_in[0][512] ) );
  NAND U9648 ( .A(init), .B(round_reg[513]), .Z(n3736) );
  NANDN U9649 ( .A(init), .B(in[513]), .Z(n3735) );
  NAND U9650 ( .A(n3736), .B(n3735), .Z(\round_in[0][513] ) );
  NAND U9651 ( .A(init), .B(round_reg[514]), .Z(n3738) );
  NANDN U9652 ( .A(init), .B(in[514]), .Z(n3737) );
  NAND U9653 ( .A(n3738), .B(n3737), .Z(\round_in[0][514] ) );
  NAND U9654 ( .A(init), .B(round_reg[515]), .Z(n3740) );
  NANDN U9655 ( .A(init), .B(in[515]), .Z(n3739) );
  NAND U9656 ( .A(n3740), .B(n3739), .Z(\round_in[0][515] ) );
  NAND U9657 ( .A(init), .B(round_reg[516]), .Z(n3742) );
  NANDN U9658 ( .A(init), .B(in[516]), .Z(n3741) );
  NAND U9659 ( .A(n3742), .B(n3741), .Z(\round_in[0][516] ) );
  NAND U9660 ( .A(init), .B(round_reg[517]), .Z(n3744) );
  NANDN U9661 ( .A(init), .B(in[517]), .Z(n3743) );
  NAND U9662 ( .A(n3744), .B(n3743), .Z(\round_in[0][517] ) );
  NAND U9663 ( .A(init), .B(round_reg[518]), .Z(n3746) );
  NANDN U9664 ( .A(init), .B(in[518]), .Z(n3745) );
  NAND U9665 ( .A(n3746), .B(n3745), .Z(\round_in[0][518] ) );
  NAND U9666 ( .A(init), .B(round_reg[519]), .Z(n3748) );
  NANDN U9667 ( .A(init), .B(in[519]), .Z(n3747) );
  NAND U9668 ( .A(n3748), .B(n3747), .Z(\round_in[0][519] ) );
  NAND U9669 ( .A(init), .B(round_reg[51]), .Z(n3750) );
  NANDN U9670 ( .A(init), .B(in[51]), .Z(n3749) );
  NAND U9671 ( .A(n3750), .B(n3749), .Z(\round_in[0][51] ) );
  NAND U9672 ( .A(init), .B(round_reg[520]), .Z(n3752) );
  NANDN U9673 ( .A(init), .B(in[520]), .Z(n3751) );
  NAND U9674 ( .A(n3752), .B(n3751), .Z(\round_in[0][520] ) );
  NAND U9675 ( .A(init), .B(round_reg[521]), .Z(n3754) );
  NANDN U9676 ( .A(init), .B(in[521]), .Z(n3753) );
  NAND U9677 ( .A(n3754), .B(n3753), .Z(\round_in[0][521] ) );
  NAND U9678 ( .A(init), .B(round_reg[522]), .Z(n3756) );
  NANDN U9679 ( .A(init), .B(in[522]), .Z(n3755) );
  NAND U9680 ( .A(n3756), .B(n3755), .Z(\round_in[0][522] ) );
  NAND U9681 ( .A(init), .B(round_reg[523]), .Z(n3758) );
  NANDN U9682 ( .A(init), .B(in[523]), .Z(n3757) );
  NAND U9683 ( .A(n3758), .B(n3757), .Z(\round_in[0][523] ) );
  NAND U9684 ( .A(init), .B(round_reg[524]), .Z(n3760) );
  NANDN U9685 ( .A(init), .B(in[524]), .Z(n3759) );
  NAND U9686 ( .A(n3760), .B(n3759), .Z(\round_in[0][524] ) );
  NAND U9687 ( .A(init), .B(round_reg[525]), .Z(n3762) );
  NANDN U9688 ( .A(init), .B(in[525]), .Z(n3761) );
  NAND U9689 ( .A(n3762), .B(n3761), .Z(\round_in[0][525] ) );
  NAND U9690 ( .A(init), .B(round_reg[526]), .Z(n3764) );
  NANDN U9691 ( .A(init), .B(in[526]), .Z(n3763) );
  NAND U9692 ( .A(n3764), .B(n3763), .Z(\round_in[0][526] ) );
  NAND U9693 ( .A(init), .B(round_reg[527]), .Z(n3766) );
  NANDN U9694 ( .A(init), .B(in[527]), .Z(n3765) );
  NAND U9695 ( .A(n3766), .B(n3765), .Z(\round_in[0][527] ) );
  NAND U9696 ( .A(init), .B(round_reg[528]), .Z(n3768) );
  NANDN U9697 ( .A(init), .B(in[528]), .Z(n3767) );
  NAND U9698 ( .A(n3768), .B(n3767), .Z(\round_in[0][528] ) );
  NAND U9699 ( .A(init), .B(round_reg[529]), .Z(n3770) );
  NANDN U9700 ( .A(init), .B(in[529]), .Z(n3769) );
  NAND U9701 ( .A(n3770), .B(n3769), .Z(\round_in[0][529] ) );
  NAND U9702 ( .A(init), .B(round_reg[52]), .Z(n3772) );
  NANDN U9703 ( .A(init), .B(in[52]), .Z(n3771) );
  NAND U9704 ( .A(n3772), .B(n3771), .Z(\round_in[0][52] ) );
  NAND U9705 ( .A(init), .B(round_reg[530]), .Z(n3774) );
  NANDN U9706 ( .A(init), .B(in[530]), .Z(n3773) );
  NAND U9707 ( .A(n3774), .B(n3773), .Z(\round_in[0][530] ) );
  NAND U9708 ( .A(init), .B(round_reg[531]), .Z(n3776) );
  NANDN U9709 ( .A(init), .B(in[531]), .Z(n3775) );
  NAND U9710 ( .A(n3776), .B(n3775), .Z(\round_in[0][531] ) );
  NAND U9711 ( .A(init), .B(round_reg[532]), .Z(n3778) );
  NANDN U9712 ( .A(init), .B(in[532]), .Z(n3777) );
  NAND U9713 ( .A(n3778), .B(n3777), .Z(\round_in[0][532] ) );
  NAND U9714 ( .A(init), .B(round_reg[533]), .Z(n3780) );
  NANDN U9715 ( .A(init), .B(in[533]), .Z(n3779) );
  NAND U9716 ( .A(n3780), .B(n3779), .Z(\round_in[0][533] ) );
  NAND U9717 ( .A(init), .B(round_reg[534]), .Z(n3782) );
  NANDN U9718 ( .A(init), .B(in[534]), .Z(n3781) );
  NAND U9719 ( .A(n3782), .B(n3781), .Z(\round_in[0][534] ) );
  NAND U9720 ( .A(init), .B(round_reg[535]), .Z(n3784) );
  NANDN U9721 ( .A(init), .B(in[535]), .Z(n3783) );
  NAND U9722 ( .A(n3784), .B(n3783), .Z(\round_in[0][535] ) );
  NAND U9723 ( .A(init), .B(round_reg[536]), .Z(n3786) );
  NANDN U9724 ( .A(init), .B(in[536]), .Z(n3785) );
  NAND U9725 ( .A(n3786), .B(n3785), .Z(\round_in[0][536] ) );
  NAND U9726 ( .A(init), .B(round_reg[537]), .Z(n3788) );
  NANDN U9727 ( .A(init), .B(in[537]), .Z(n3787) );
  NAND U9728 ( .A(n3788), .B(n3787), .Z(\round_in[0][537] ) );
  NAND U9729 ( .A(init), .B(round_reg[538]), .Z(n3790) );
  NANDN U9730 ( .A(init), .B(in[538]), .Z(n3789) );
  NAND U9731 ( .A(n3790), .B(n3789), .Z(\round_in[0][538] ) );
  NAND U9732 ( .A(init), .B(round_reg[539]), .Z(n3792) );
  NANDN U9733 ( .A(init), .B(in[539]), .Z(n3791) );
  NAND U9734 ( .A(n3792), .B(n3791), .Z(\round_in[0][539] ) );
  NAND U9735 ( .A(init), .B(round_reg[53]), .Z(n3794) );
  NANDN U9736 ( .A(init), .B(in[53]), .Z(n3793) );
  NAND U9737 ( .A(n3794), .B(n3793), .Z(\round_in[0][53] ) );
  NAND U9738 ( .A(init), .B(round_reg[540]), .Z(n3796) );
  NANDN U9739 ( .A(init), .B(in[540]), .Z(n3795) );
  NAND U9740 ( .A(n3796), .B(n3795), .Z(\round_in[0][540] ) );
  NAND U9741 ( .A(init), .B(round_reg[541]), .Z(n3798) );
  NANDN U9742 ( .A(init), .B(in[541]), .Z(n3797) );
  NAND U9743 ( .A(n3798), .B(n3797), .Z(\round_in[0][541] ) );
  NAND U9744 ( .A(init), .B(round_reg[542]), .Z(n3800) );
  NANDN U9745 ( .A(init), .B(in[542]), .Z(n3799) );
  NAND U9746 ( .A(n3800), .B(n3799), .Z(\round_in[0][542] ) );
  NAND U9747 ( .A(init), .B(round_reg[543]), .Z(n3802) );
  NANDN U9748 ( .A(init), .B(in[543]), .Z(n3801) );
  NAND U9749 ( .A(n3802), .B(n3801), .Z(\round_in[0][543] ) );
  NAND U9750 ( .A(init), .B(round_reg[544]), .Z(n3804) );
  NANDN U9751 ( .A(init), .B(in[544]), .Z(n3803) );
  NAND U9752 ( .A(n3804), .B(n3803), .Z(\round_in[0][544] ) );
  NAND U9753 ( .A(init), .B(round_reg[545]), .Z(n3806) );
  NANDN U9754 ( .A(init), .B(in[545]), .Z(n3805) );
  NAND U9755 ( .A(n3806), .B(n3805), .Z(\round_in[0][545] ) );
  NAND U9756 ( .A(init), .B(round_reg[546]), .Z(n3808) );
  NANDN U9757 ( .A(init), .B(in[546]), .Z(n3807) );
  NAND U9758 ( .A(n3808), .B(n3807), .Z(\round_in[0][546] ) );
  NAND U9759 ( .A(init), .B(round_reg[547]), .Z(n3810) );
  NANDN U9760 ( .A(init), .B(in[547]), .Z(n3809) );
  NAND U9761 ( .A(n3810), .B(n3809), .Z(\round_in[0][547] ) );
  NAND U9762 ( .A(init), .B(round_reg[548]), .Z(n3812) );
  NANDN U9763 ( .A(init), .B(in[548]), .Z(n3811) );
  NAND U9764 ( .A(n3812), .B(n3811), .Z(\round_in[0][548] ) );
  NAND U9765 ( .A(init), .B(round_reg[549]), .Z(n3814) );
  NANDN U9766 ( .A(init), .B(in[549]), .Z(n3813) );
  NAND U9767 ( .A(n3814), .B(n3813), .Z(\round_in[0][549] ) );
  NAND U9768 ( .A(init), .B(round_reg[54]), .Z(n3816) );
  NANDN U9769 ( .A(init), .B(in[54]), .Z(n3815) );
  NAND U9770 ( .A(n3816), .B(n3815), .Z(\round_in[0][54] ) );
  NAND U9771 ( .A(init), .B(round_reg[550]), .Z(n3818) );
  NANDN U9772 ( .A(init), .B(in[550]), .Z(n3817) );
  NAND U9773 ( .A(n3818), .B(n3817), .Z(\round_in[0][550] ) );
  NAND U9774 ( .A(init), .B(round_reg[551]), .Z(n3820) );
  NANDN U9775 ( .A(init), .B(in[551]), .Z(n3819) );
  NAND U9776 ( .A(n3820), .B(n3819), .Z(\round_in[0][551] ) );
  NAND U9777 ( .A(init), .B(round_reg[552]), .Z(n3822) );
  NANDN U9778 ( .A(init), .B(in[552]), .Z(n3821) );
  NAND U9779 ( .A(n3822), .B(n3821), .Z(\round_in[0][552] ) );
  NAND U9780 ( .A(init), .B(round_reg[553]), .Z(n3824) );
  NANDN U9781 ( .A(init), .B(in[553]), .Z(n3823) );
  NAND U9782 ( .A(n3824), .B(n3823), .Z(\round_in[0][553] ) );
  NAND U9783 ( .A(init), .B(round_reg[554]), .Z(n3826) );
  NANDN U9784 ( .A(init), .B(in[554]), .Z(n3825) );
  NAND U9785 ( .A(n3826), .B(n3825), .Z(\round_in[0][554] ) );
  NAND U9786 ( .A(init), .B(round_reg[555]), .Z(n3828) );
  NANDN U9787 ( .A(init), .B(in[555]), .Z(n3827) );
  NAND U9788 ( .A(n3828), .B(n3827), .Z(\round_in[0][555] ) );
  NAND U9789 ( .A(init), .B(round_reg[556]), .Z(n3830) );
  NANDN U9790 ( .A(init), .B(in[556]), .Z(n3829) );
  NAND U9791 ( .A(n3830), .B(n3829), .Z(\round_in[0][556] ) );
  NAND U9792 ( .A(init), .B(round_reg[557]), .Z(n3832) );
  NANDN U9793 ( .A(init), .B(in[557]), .Z(n3831) );
  NAND U9794 ( .A(n3832), .B(n3831), .Z(\round_in[0][557] ) );
  NAND U9795 ( .A(init), .B(round_reg[558]), .Z(n3834) );
  NANDN U9796 ( .A(init), .B(in[558]), .Z(n3833) );
  NAND U9797 ( .A(n3834), .B(n3833), .Z(\round_in[0][558] ) );
  NAND U9798 ( .A(init), .B(round_reg[559]), .Z(n3836) );
  NANDN U9799 ( .A(init), .B(in[559]), .Z(n3835) );
  NAND U9800 ( .A(n3836), .B(n3835), .Z(\round_in[0][559] ) );
  NAND U9801 ( .A(init), .B(round_reg[55]), .Z(n3838) );
  NANDN U9802 ( .A(init), .B(in[55]), .Z(n3837) );
  NAND U9803 ( .A(n3838), .B(n3837), .Z(\round_in[0][55] ) );
  NAND U9804 ( .A(init), .B(round_reg[560]), .Z(n3840) );
  NANDN U9805 ( .A(init), .B(in[560]), .Z(n3839) );
  NAND U9806 ( .A(n3840), .B(n3839), .Z(\round_in[0][560] ) );
  NAND U9807 ( .A(init), .B(round_reg[561]), .Z(n3842) );
  NANDN U9808 ( .A(init), .B(in[561]), .Z(n3841) );
  NAND U9809 ( .A(n3842), .B(n3841), .Z(\round_in[0][561] ) );
  NAND U9810 ( .A(init), .B(round_reg[562]), .Z(n3844) );
  NANDN U9811 ( .A(init), .B(in[562]), .Z(n3843) );
  NAND U9812 ( .A(n3844), .B(n3843), .Z(\round_in[0][562] ) );
  NAND U9813 ( .A(init), .B(round_reg[563]), .Z(n3846) );
  NANDN U9814 ( .A(init), .B(in[563]), .Z(n3845) );
  NAND U9815 ( .A(n3846), .B(n3845), .Z(\round_in[0][563] ) );
  NAND U9816 ( .A(init), .B(round_reg[564]), .Z(n3848) );
  NANDN U9817 ( .A(init), .B(in[564]), .Z(n3847) );
  NAND U9818 ( .A(n3848), .B(n3847), .Z(\round_in[0][564] ) );
  NAND U9819 ( .A(init), .B(round_reg[565]), .Z(n3850) );
  NANDN U9820 ( .A(init), .B(in[565]), .Z(n3849) );
  NAND U9821 ( .A(n3850), .B(n3849), .Z(\round_in[0][565] ) );
  NAND U9822 ( .A(init), .B(round_reg[566]), .Z(n3852) );
  NANDN U9823 ( .A(init), .B(in[566]), .Z(n3851) );
  NAND U9824 ( .A(n3852), .B(n3851), .Z(\round_in[0][566] ) );
  NAND U9825 ( .A(init), .B(round_reg[567]), .Z(n3854) );
  NANDN U9826 ( .A(init), .B(in[567]), .Z(n3853) );
  NAND U9827 ( .A(n3854), .B(n3853), .Z(\round_in[0][567] ) );
  NAND U9828 ( .A(init), .B(round_reg[568]), .Z(n3856) );
  NANDN U9829 ( .A(init), .B(in[568]), .Z(n3855) );
  NAND U9830 ( .A(n3856), .B(n3855), .Z(\round_in[0][568] ) );
  NAND U9831 ( .A(init), .B(round_reg[569]), .Z(n3858) );
  NANDN U9832 ( .A(init), .B(in[569]), .Z(n3857) );
  NAND U9833 ( .A(n3858), .B(n3857), .Z(\round_in[0][569] ) );
  NAND U9834 ( .A(init), .B(round_reg[56]), .Z(n3860) );
  NANDN U9835 ( .A(init), .B(in[56]), .Z(n3859) );
  NAND U9836 ( .A(n3860), .B(n3859), .Z(\round_in[0][56] ) );
  NAND U9837 ( .A(init), .B(round_reg[570]), .Z(n3862) );
  NANDN U9838 ( .A(init), .B(in[570]), .Z(n3861) );
  NAND U9839 ( .A(n3862), .B(n3861), .Z(\round_in[0][570] ) );
  NAND U9840 ( .A(init), .B(round_reg[571]), .Z(n3864) );
  NANDN U9841 ( .A(init), .B(in[571]), .Z(n3863) );
  NAND U9842 ( .A(n3864), .B(n3863), .Z(\round_in[0][571] ) );
  NAND U9843 ( .A(init), .B(round_reg[572]), .Z(n3866) );
  NANDN U9844 ( .A(init), .B(in[572]), .Z(n3865) );
  NAND U9845 ( .A(n3866), .B(n3865), .Z(\round_in[0][572] ) );
  NAND U9846 ( .A(init), .B(round_reg[573]), .Z(n3868) );
  NANDN U9847 ( .A(init), .B(in[573]), .Z(n3867) );
  NAND U9848 ( .A(n3868), .B(n3867), .Z(\round_in[0][573] ) );
  NAND U9849 ( .A(init), .B(round_reg[574]), .Z(n3870) );
  NANDN U9850 ( .A(init), .B(in[574]), .Z(n3869) );
  NAND U9851 ( .A(n3870), .B(n3869), .Z(\round_in[0][574] ) );
  NAND U9852 ( .A(init), .B(round_reg[575]), .Z(n3872) );
  NANDN U9853 ( .A(init), .B(in[575]), .Z(n3871) );
  NAND U9854 ( .A(n3872), .B(n3871), .Z(\round_in[0][575] ) );
  AND U9855 ( .A(round_reg[576]), .B(init), .Z(\round_in[0][576] ) );
  AND U9856 ( .A(round_reg[577]), .B(init), .Z(\round_in[0][577] ) );
  AND U9857 ( .A(round_reg[578]), .B(init), .Z(\round_in[0][578] ) );
  AND U9858 ( .A(round_reg[579]), .B(init), .Z(\round_in[0][579] ) );
  NAND U9859 ( .A(init), .B(round_reg[57]), .Z(n3874) );
  NANDN U9860 ( .A(init), .B(in[57]), .Z(n3873) );
  NAND U9861 ( .A(n3874), .B(n3873), .Z(\round_in[0][57] ) );
  AND U9862 ( .A(round_reg[580]), .B(init), .Z(\round_in[0][580] ) );
  AND U9863 ( .A(round_reg[581]), .B(init), .Z(\round_in[0][581] ) );
  AND U9864 ( .A(round_reg[582]), .B(init), .Z(\round_in[0][582] ) );
  AND U9865 ( .A(round_reg[583]), .B(init), .Z(\round_in[0][583] ) );
  AND U9866 ( .A(round_reg[584]), .B(init), .Z(\round_in[0][584] ) );
  AND U9867 ( .A(round_reg[585]), .B(init), .Z(\round_in[0][585] ) );
  AND U9868 ( .A(round_reg[586]), .B(init), .Z(\round_in[0][586] ) );
  AND U9869 ( .A(round_reg[587]), .B(init), .Z(\round_in[0][587] ) );
  AND U9870 ( .A(round_reg[588]), .B(init), .Z(\round_in[0][588] ) );
  AND U9871 ( .A(round_reg[589]), .B(init), .Z(\round_in[0][589] ) );
  NAND U9872 ( .A(init), .B(round_reg[58]), .Z(n3876) );
  NANDN U9873 ( .A(init), .B(in[58]), .Z(n3875) );
  NAND U9874 ( .A(n3876), .B(n3875), .Z(\round_in[0][58] ) );
  AND U9875 ( .A(round_reg[590]), .B(init), .Z(\round_in[0][590] ) );
  AND U9876 ( .A(round_reg[591]), .B(init), .Z(\round_in[0][591] ) );
  AND U9877 ( .A(round_reg[592]), .B(init), .Z(\round_in[0][592] ) );
  AND U9878 ( .A(round_reg[593]), .B(init), .Z(\round_in[0][593] ) );
  AND U9879 ( .A(round_reg[594]), .B(init), .Z(\round_in[0][594] ) );
  AND U9880 ( .A(round_reg[595]), .B(init), .Z(\round_in[0][595] ) );
  AND U9881 ( .A(round_reg[596]), .B(init), .Z(\round_in[0][596] ) );
  AND U9882 ( .A(round_reg[597]), .B(init), .Z(\round_in[0][597] ) );
  AND U9883 ( .A(round_reg[598]), .B(init), .Z(\round_in[0][598] ) );
  AND U9884 ( .A(round_reg[599]), .B(init), .Z(\round_in[0][599] ) );
  NAND U9885 ( .A(init), .B(round_reg[59]), .Z(n3878) );
  NANDN U9886 ( .A(init), .B(in[59]), .Z(n3877) );
  NAND U9887 ( .A(n3878), .B(n3877), .Z(\round_in[0][59] ) );
  NAND U9888 ( .A(init), .B(round_reg[5]), .Z(n3880) );
  NANDN U9889 ( .A(init), .B(in[5]), .Z(n3879) );
  NAND U9890 ( .A(n3880), .B(n3879), .Z(\round_in[0][5] ) );
  AND U9891 ( .A(round_reg[600]), .B(init), .Z(\round_in[0][600] ) );
  AND U9892 ( .A(round_reg[601]), .B(init), .Z(\round_in[0][601] ) );
  AND U9893 ( .A(round_reg[602]), .B(init), .Z(\round_in[0][602] ) );
  AND U9894 ( .A(round_reg[603]), .B(init), .Z(\round_in[0][603] ) );
  AND U9895 ( .A(round_reg[604]), .B(init), .Z(\round_in[0][604] ) );
  AND U9896 ( .A(round_reg[605]), .B(init), .Z(\round_in[0][605] ) );
  AND U9897 ( .A(round_reg[606]), .B(init), .Z(\round_in[0][606] ) );
  AND U9898 ( .A(round_reg[607]), .B(init), .Z(\round_in[0][607] ) );
  AND U9899 ( .A(round_reg[608]), .B(init), .Z(\round_in[0][608] ) );
  AND U9900 ( .A(round_reg[609]), .B(init), .Z(\round_in[0][609] ) );
  NAND U9901 ( .A(init), .B(round_reg[60]), .Z(n3882) );
  NANDN U9902 ( .A(init), .B(in[60]), .Z(n3881) );
  NAND U9903 ( .A(n3882), .B(n3881), .Z(\round_in[0][60] ) );
  AND U9904 ( .A(round_reg[610]), .B(init), .Z(\round_in[0][610] ) );
  AND U9905 ( .A(round_reg[611]), .B(init), .Z(\round_in[0][611] ) );
  AND U9906 ( .A(round_reg[612]), .B(init), .Z(\round_in[0][612] ) );
  AND U9907 ( .A(round_reg[613]), .B(init), .Z(\round_in[0][613] ) );
  AND U9908 ( .A(round_reg[614]), .B(init), .Z(\round_in[0][614] ) );
  AND U9909 ( .A(round_reg[615]), .B(init), .Z(\round_in[0][615] ) );
  AND U9910 ( .A(round_reg[616]), .B(init), .Z(\round_in[0][616] ) );
  AND U9911 ( .A(round_reg[617]), .B(init), .Z(\round_in[0][617] ) );
  AND U9912 ( .A(round_reg[618]), .B(init), .Z(\round_in[0][618] ) );
  AND U9913 ( .A(round_reg[619]), .B(init), .Z(\round_in[0][619] ) );
  NAND U9914 ( .A(init), .B(round_reg[61]), .Z(n3884) );
  NANDN U9915 ( .A(init), .B(in[61]), .Z(n3883) );
  NAND U9916 ( .A(n3884), .B(n3883), .Z(\round_in[0][61] ) );
  AND U9917 ( .A(round_reg[620]), .B(init), .Z(\round_in[0][620] ) );
  AND U9918 ( .A(round_reg[621]), .B(init), .Z(\round_in[0][621] ) );
  AND U9919 ( .A(round_reg[622]), .B(init), .Z(\round_in[0][622] ) );
  AND U9920 ( .A(round_reg[623]), .B(init), .Z(\round_in[0][623] ) );
  AND U9921 ( .A(round_reg[624]), .B(init), .Z(\round_in[0][624] ) );
  AND U9922 ( .A(round_reg[625]), .B(init), .Z(\round_in[0][625] ) );
  AND U9923 ( .A(round_reg[626]), .B(init), .Z(\round_in[0][626] ) );
  AND U9924 ( .A(round_reg[627]), .B(init), .Z(\round_in[0][627] ) );
  AND U9925 ( .A(round_reg[628]), .B(init), .Z(\round_in[0][628] ) );
  AND U9926 ( .A(round_reg[629]), .B(init), .Z(\round_in[0][629] ) );
  NAND U9927 ( .A(init), .B(round_reg[62]), .Z(n3886) );
  NANDN U9928 ( .A(init), .B(in[62]), .Z(n3885) );
  NAND U9929 ( .A(n3886), .B(n3885), .Z(\round_in[0][62] ) );
  AND U9930 ( .A(round_reg[630]), .B(init), .Z(\round_in[0][630] ) );
  AND U9931 ( .A(round_reg[631]), .B(init), .Z(\round_in[0][631] ) );
  AND U9932 ( .A(round_reg[632]), .B(init), .Z(\round_in[0][632] ) );
  AND U9933 ( .A(round_reg[633]), .B(init), .Z(\round_in[0][633] ) );
  AND U9934 ( .A(round_reg[634]), .B(init), .Z(\round_in[0][634] ) );
  AND U9935 ( .A(round_reg[635]), .B(init), .Z(\round_in[0][635] ) );
  AND U9936 ( .A(round_reg[636]), .B(init), .Z(\round_in[0][636] ) );
  AND U9937 ( .A(round_reg[637]), .B(init), .Z(\round_in[0][637] ) );
  AND U9938 ( .A(round_reg[638]), .B(init), .Z(\round_in[0][638] ) );
  AND U9939 ( .A(round_reg[639]), .B(init), .Z(\round_in[0][639] ) );
  NAND U9940 ( .A(init), .B(round_reg[63]), .Z(n3888) );
  NANDN U9941 ( .A(init), .B(in[63]), .Z(n3887) );
  NAND U9942 ( .A(n3888), .B(n3887), .Z(\round_in[0][63] ) );
  AND U9943 ( .A(round_reg[640]), .B(init), .Z(\round_in[0][640] ) );
  AND U9944 ( .A(round_reg[641]), .B(init), .Z(\round_in[0][641] ) );
  AND U9945 ( .A(round_reg[642]), .B(init), .Z(\round_in[0][642] ) );
  AND U9946 ( .A(round_reg[643]), .B(init), .Z(\round_in[0][643] ) );
  AND U9947 ( .A(round_reg[644]), .B(init), .Z(\round_in[0][644] ) );
  AND U9948 ( .A(round_reg[645]), .B(init), .Z(\round_in[0][645] ) );
  AND U9949 ( .A(round_reg[646]), .B(init), .Z(\round_in[0][646] ) );
  AND U9950 ( .A(round_reg[647]), .B(init), .Z(\round_in[0][647] ) );
  AND U9951 ( .A(round_reg[648]), .B(init), .Z(\round_in[0][648] ) );
  AND U9952 ( .A(round_reg[649]), .B(init), .Z(\round_in[0][649] ) );
  NAND U9953 ( .A(init), .B(round_reg[64]), .Z(n3890) );
  NANDN U9954 ( .A(init), .B(in[64]), .Z(n3889) );
  NAND U9955 ( .A(n3890), .B(n3889), .Z(\round_in[0][64] ) );
  AND U9956 ( .A(round_reg[650]), .B(init), .Z(\round_in[0][650] ) );
  AND U9957 ( .A(round_reg[651]), .B(init), .Z(\round_in[0][651] ) );
  AND U9958 ( .A(round_reg[652]), .B(init), .Z(\round_in[0][652] ) );
  AND U9959 ( .A(round_reg[653]), .B(init), .Z(\round_in[0][653] ) );
  AND U9960 ( .A(round_reg[654]), .B(init), .Z(\round_in[0][654] ) );
  AND U9961 ( .A(round_reg[655]), .B(init), .Z(\round_in[0][655] ) );
  AND U9962 ( .A(round_reg[656]), .B(init), .Z(\round_in[0][656] ) );
  AND U9963 ( .A(round_reg[657]), .B(init), .Z(\round_in[0][657] ) );
  AND U9964 ( .A(round_reg[658]), .B(init), .Z(\round_in[0][658] ) );
  AND U9965 ( .A(round_reg[659]), .B(init), .Z(\round_in[0][659] ) );
  NAND U9966 ( .A(init), .B(round_reg[65]), .Z(n3892) );
  NANDN U9967 ( .A(init), .B(in[65]), .Z(n3891) );
  NAND U9968 ( .A(n3892), .B(n3891), .Z(\round_in[0][65] ) );
  AND U9969 ( .A(round_reg[660]), .B(init), .Z(\round_in[0][660] ) );
  AND U9970 ( .A(round_reg[661]), .B(init), .Z(\round_in[0][661] ) );
  AND U9971 ( .A(round_reg[662]), .B(init), .Z(\round_in[0][662] ) );
  AND U9972 ( .A(round_reg[663]), .B(init), .Z(\round_in[0][663] ) );
  AND U9973 ( .A(round_reg[664]), .B(init), .Z(\round_in[0][664] ) );
  AND U9974 ( .A(round_reg[665]), .B(init), .Z(\round_in[0][665] ) );
  AND U9975 ( .A(round_reg[666]), .B(init), .Z(\round_in[0][666] ) );
  AND U9976 ( .A(round_reg[667]), .B(init), .Z(\round_in[0][667] ) );
  AND U9977 ( .A(round_reg[668]), .B(init), .Z(\round_in[0][668] ) );
  AND U9978 ( .A(round_reg[669]), .B(init), .Z(\round_in[0][669] ) );
  NAND U9979 ( .A(init), .B(round_reg[66]), .Z(n3894) );
  NANDN U9980 ( .A(init), .B(in[66]), .Z(n3893) );
  NAND U9981 ( .A(n3894), .B(n3893), .Z(\round_in[0][66] ) );
  AND U9982 ( .A(round_reg[670]), .B(init), .Z(\round_in[0][670] ) );
  AND U9983 ( .A(round_reg[671]), .B(init), .Z(\round_in[0][671] ) );
  AND U9984 ( .A(round_reg[672]), .B(init), .Z(\round_in[0][672] ) );
  AND U9985 ( .A(round_reg[673]), .B(init), .Z(\round_in[0][673] ) );
  AND U9986 ( .A(round_reg[674]), .B(init), .Z(\round_in[0][674] ) );
  AND U9987 ( .A(round_reg[675]), .B(init), .Z(\round_in[0][675] ) );
  AND U9988 ( .A(round_reg[676]), .B(init), .Z(\round_in[0][676] ) );
  AND U9989 ( .A(round_reg[677]), .B(init), .Z(\round_in[0][677] ) );
  AND U9990 ( .A(round_reg[678]), .B(init), .Z(\round_in[0][678] ) );
  AND U9991 ( .A(round_reg[679]), .B(init), .Z(\round_in[0][679] ) );
  NAND U9992 ( .A(init), .B(round_reg[67]), .Z(n3896) );
  NANDN U9993 ( .A(init), .B(in[67]), .Z(n3895) );
  NAND U9994 ( .A(n3896), .B(n3895), .Z(\round_in[0][67] ) );
  AND U9995 ( .A(round_reg[680]), .B(init), .Z(\round_in[0][680] ) );
  AND U9996 ( .A(round_reg[681]), .B(init), .Z(\round_in[0][681] ) );
  AND U9997 ( .A(round_reg[682]), .B(init), .Z(\round_in[0][682] ) );
  AND U9998 ( .A(round_reg[683]), .B(init), .Z(\round_in[0][683] ) );
  AND U9999 ( .A(round_reg[684]), .B(init), .Z(\round_in[0][684] ) );
  AND U10000 ( .A(round_reg[685]), .B(init), .Z(\round_in[0][685] ) );
  AND U10001 ( .A(round_reg[686]), .B(init), .Z(\round_in[0][686] ) );
  AND U10002 ( .A(round_reg[687]), .B(init), .Z(\round_in[0][687] ) );
  AND U10003 ( .A(round_reg[688]), .B(init), .Z(\round_in[0][688] ) );
  AND U10004 ( .A(round_reg[689]), .B(init), .Z(\round_in[0][689] ) );
  NAND U10005 ( .A(init), .B(round_reg[68]), .Z(n3898) );
  NANDN U10006 ( .A(init), .B(in[68]), .Z(n3897) );
  NAND U10007 ( .A(n3898), .B(n3897), .Z(\round_in[0][68] ) );
  AND U10008 ( .A(round_reg[690]), .B(init), .Z(\round_in[0][690] ) );
  AND U10009 ( .A(round_reg[691]), .B(init), .Z(\round_in[0][691] ) );
  AND U10010 ( .A(round_reg[692]), .B(init), .Z(\round_in[0][692] ) );
  AND U10011 ( .A(round_reg[693]), .B(init), .Z(\round_in[0][693] ) );
  AND U10012 ( .A(round_reg[694]), .B(init), .Z(\round_in[0][694] ) );
  AND U10013 ( .A(round_reg[695]), .B(init), .Z(\round_in[0][695] ) );
  AND U10014 ( .A(round_reg[696]), .B(init), .Z(\round_in[0][696] ) );
  AND U10015 ( .A(round_reg[697]), .B(init), .Z(\round_in[0][697] ) );
  AND U10016 ( .A(round_reg[698]), .B(init), .Z(\round_in[0][698] ) );
  AND U10017 ( .A(round_reg[699]), .B(init), .Z(\round_in[0][699] ) );
  NAND U10018 ( .A(init), .B(round_reg[69]), .Z(n3900) );
  NANDN U10019 ( .A(init), .B(in[69]), .Z(n3899) );
  NAND U10020 ( .A(n3900), .B(n3899), .Z(\round_in[0][69] ) );
  NAND U10021 ( .A(init), .B(round_reg[6]), .Z(n3902) );
  NANDN U10022 ( .A(init), .B(in[6]), .Z(n3901) );
  NAND U10023 ( .A(n3902), .B(n3901), .Z(\round_in[0][6] ) );
  AND U10024 ( .A(round_reg[700]), .B(init), .Z(\round_in[0][700] ) );
  AND U10025 ( .A(round_reg[701]), .B(init), .Z(\round_in[0][701] ) );
  AND U10026 ( .A(round_reg[702]), .B(init), .Z(\round_in[0][702] ) );
  AND U10027 ( .A(round_reg[703]), .B(init), .Z(\round_in[0][703] ) );
  AND U10028 ( .A(round_reg[704]), .B(init), .Z(\round_in[0][704] ) );
  AND U10029 ( .A(round_reg[705]), .B(init), .Z(\round_in[0][705] ) );
  AND U10030 ( .A(round_reg[706]), .B(init), .Z(\round_in[0][706] ) );
  AND U10031 ( .A(round_reg[707]), .B(init), .Z(\round_in[0][707] ) );
  AND U10032 ( .A(round_reg[708]), .B(init), .Z(\round_in[0][708] ) );
  AND U10033 ( .A(round_reg[709]), .B(init), .Z(\round_in[0][709] ) );
  NAND U10034 ( .A(init), .B(round_reg[70]), .Z(n3904) );
  NANDN U10035 ( .A(init), .B(in[70]), .Z(n3903) );
  NAND U10036 ( .A(n3904), .B(n3903), .Z(\round_in[0][70] ) );
  AND U10037 ( .A(round_reg[710]), .B(init), .Z(\round_in[0][710] ) );
  AND U10038 ( .A(round_reg[711]), .B(init), .Z(\round_in[0][711] ) );
  AND U10039 ( .A(round_reg[712]), .B(init), .Z(\round_in[0][712] ) );
  AND U10040 ( .A(round_reg[713]), .B(init), .Z(\round_in[0][713] ) );
  AND U10041 ( .A(round_reg[714]), .B(init), .Z(\round_in[0][714] ) );
  AND U10042 ( .A(round_reg[715]), .B(init), .Z(\round_in[0][715] ) );
  AND U10043 ( .A(round_reg[716]), .B(init), .Z(\round_in[0][716] ) );
  AND U10044 ( .A(round_reg[717]), .B(init), .Z(\round_in[0][717] ) );
  AND U10045 ( .A(round_reg[718]), .B(init), .Z(\round_in[0][718] ) );
  AND U10046 ( .A(round_reg[719]), .B(init), .Z(\round_in[0][719] ) );
  NAND U10047 ( .A(init), .B(round_reg[71]), .Z(n3906) );
  NANDN U10048 ( .A(init), .B(in[71]), .Z(n3905) );
  NAND U10049 ( .A(n3906), .B(n3905), .Z(\round_in[0][71] ) );
  AND U10050 ( .A(round_reg[720]), .B(init), .Z(\round_in[0][720] ) );
  AND U10051 ( .A(round_reg[721]), .B(init), .Z(\round_in[0][721] ) );
  AND U10052 ( .A(round_reg[722]), .B(init), .Z(\round_in[0][722] ) );
  AND U10053 ( .A(round_reg[723]), .B(init), .Z(\round_in[0][723] ) );
  AND U10054 ( .A(round_reg[724]), .B(init), .Z(\round_in[0][724] ) );
  AND U10055 ( .A(round_reg[725]), .B(init), .Z(\round_in[0][725] ) );
  AND U10056 ( .A(round_reg[726]), .B(init), .Z(\round_in[0][726] ) );
  AND U10057 ( .A(round_reg[727]), .B(init), .Z(\round_in[0][727] ) );
  AND U10058 ( .A(round_reg[728]), .B(init), .Z(\round_in[0][728] ) );
  AND U10059 ( .A(round_reg[729]), .B(init), .Z(\round_in[0][729] ) );
  NAND U10060 ( .A(init), .B(round_reg[72]), .Z(n3908) );
  NANDN U10061 ( .A(init), .B(in[72]), .Z(n3907) );
  NAND U10062 ( .A(n3908), .B(n3907), .Z(\round_in[0][72] ) );
  AND U10063 ( .A(round_reg[730]), .B(init), .Z(\round_in[0][730] ) );
  AND U10064 ( .A(round_reg[731]), .B(init), .Z(\round_in[0][731] ) );
  AND U10065 ( .A(round_reg[732]), .B(init), .Z(\round_in[0][732] ) );
  AND U10066 ( .A(round_reg[733]), .B(init), .Z(\round_in[0][733] ) );
  AND U10067 ( .A(round_reg[734]), .B(init), .Z(\round_in[0][734] ) );
  AND U10068 ( .A(round_reg[735]), .B(init), .Z(\round_in[0][735] ) );
  AND U10069 ( .A(round_reg[736]), .B(init), .Z(\round_in[0][736] ) );
  AND U10070 ( .A(round_reg[737]), .B(init), .Z(\round_in[0][737] ) );
  AND U10071 ( .A(round_reg[738]), .B(init), .Z(\round_in[0][738] ) );
  AND U10072 ( .A(round_reg[739]), .B(init), .Z(\round_in[0][739] ) );
  NAND U10073 ( .A(init), .B(round_reg[73]), .Z(n3910) );
  NANDN U10074 ( .A(init), .B(in[73]), .Z(n3909) );
  NAND U10075 ( .A(n3910), .B(n3909), .Z(\round_in[0][73] ) );
  AND U10076 ( .A(round_reg[740]), .B(init), .Z(\round_in[0][740] ) );
  AND U10077 ( .A(round_reg[741]), .B(init), .Z(\round_in[0][741] ) );
  AND U10078 ( .A(round_reg[742]), .B(init), .Z(\round_in[0][742] ) );
  AND U10079 ( .A(round_reg[743]), .B(init), .Z(\round_in[0][743] ) );
  AND U10080 ( .A(round_reg[744]), .B(init), .Z(\round_in[0][744] ) );
  AND U10081 ( .A(round_reg[745]), .B(init), .Z(\round_in[0][745] ) );
  AND U10082 ( .A(round_reg[746]), .B(init), .Z(\round_in[0][746] ) );
  AND U10083 ( .A(round_reg[747]), .B(init), .Z(\round_in[0][747] ) );
  AND U10084 ( .A(round_reg[748]), .B(init), .Z(\round_in[0][748] ) );
  AND U10085 ( .A(round_reg[749]), .B(init), .Z(\round_in[0][749] ) );
  NAND U10086 ( .A(init), .B(round_reg[74]), .Z(n3912) );
  NANDN U10087 ( .A(init), .B(in[74]), .Z(n3911) );
  NAND U10088 ( .A(n3912), .B(n3911), .Z(\round_in[0][74] ) );
  AND U10089 ( .A(round_reg[750]), .B(init), .Z(\round_in[0][750] ) );
  AND U10090 ( .A(round_reg[751]), .B(init), .Z(\round_in[0][751] ) );
  AND U10091 ( .A(round_reg[752]), .B(init), .Z(\round_in[0][752] ) );
  AND U10092 ( .A(round_reg[753]), .B(init), .Z(\round_in[0][753] ) );
  AND U10093 ( .A(round_reg[754]), .B(init), .Z(\round_in[0][754] ) );
  AND U10094 ( .A(round_reg[755]), .B(init), .Z(\round_in[0][755] ) );
  AND U10095 ( .A(round_reg[756]), .B(init), .Z(\round_in[0][756] ) );
  AND U10096 ( .A(round_reg[757]), .B(init), .Z(\round_in[0][757] ) );
  AND U10097 ( .A(round_reg[758]), .B(init), .Z(\round_in[0][758] ) );
  AND U10098 ( .A(round_reg[759]), .B(init), .Z(\round_in[0][759] ) );
  NAND U10099 ( .A(init), .B(round_reg[75]), .Z(n3914) );
  NANDN U10100 ( .A(init), .B(in[75]), .Z(n3913) );
  NAND U10101 ( .A(n3914), .B(n3913), .Z(\round_in[0][75] ) );
  AND U10102 ( .A(round_reg[760]), .B(init), .Z(\round_in[0][760] ) );
  AND U10103 ( .A(round_reg[761]), .B(init), .Z(\round_in[0][761] ) );
  AND U10104 ( .A(round_reg[762]), .B(init), .Z(\round_in[0][762] ) );
  AND U10105 ( .A(round_reg[763]), .B(init), .Z(\round_in[0][763] ) );
  AND U10106 ( .A(round_reg[764]), .B(init), .Z(\round_in[0][764] ) );
  AND U10107 ( .A(round_reg[765]), .B(init), .Z(\round_in[0][765] ) );
  AND U10108 ( .A(round_reg[766]), .B(init), .Z(\round_in[0][766] ) );
  AND U10109 ( .A(round_reg[767]), .B(init), .Z(\round_in[0][767] ) );
  AND U10110 ( .A(round_reg[768]), .B(init), .Z(\round_in[0][768] ) );
  AND U10111 ( .A(round_reg[769]), .B(init), .Z(\round_in[0][769] ) );
  NAND U10112 ( .A(init), .B(round_reg[76]), .Z(n3916) );
  NANDN U10113 ( .A(init), .B(in[76]), .Z(n3915) );
  NAND U10114 ( .A(n3916), .B(n3915), .Z(\round_in[0][76] ) );
  AND U10115 ( .A(round_reg[770]), .B(init), .Z(\round_in[0][770] ) );
  AND U10116 ( .A(round_reg[771]), .B(init), .Z(\round_in[0][771] ) );
  AND U10117 ( .A(round_reg[772]), .B(init), .Z(\round_in[0][772] ) );
  AND U10118 ( .A(round_reg[773]), .B(init), .Z(\round_in[0][773] ) );
  AND U10119 ( .A(round_reg[774]), .B(init), .Z(\round_in[0][774] ) );
  AND U10120 ( .A(round_reg[775]), .B(init), .Z(\round_in[0][775] ) );
  AND U10121 ( .A(round_reg[776]), .B(init), .Z(\round_in[0][776] ) );
  AND U10122 ( .A(round_reg[777]), .B(init), .Z(\round_in[0][777] ) );
  AND U10123 ( .A(round_reg[778]), .B(init), .Z(\round_in[0][778] ) );
  AND U10124 ( .A(round_reg[779]), .B(init), .Z(\round_in[0][779] ) );
  NAND U10125 ( .A(init), .B(round_reg[77]), .Z(n3918) );
  NANDN U10126 ( .A(init), .B(in[77]), .Z(n3917) );
  NAND U10127 ( .A(n3918), .B(n3917), .Z(\round_in[0][77] ) );
  AND U10128 ( .A(round_reg[780]), .B(init), .Z(\round_in[0][780] ) );
  AND U10129 ( .A(round_reg[781]), .B(init), .Z(\round_in[0][781] ) );
  AND U10130 ( .A(round_reg[782]), .B(init), .Z(\round_in[0][782] ) );
  AND U10131 ( .A(round_reg[783]), .B(init), .Z(\round_in[0][783] ) );
  AND U10132 ( .A(round_reg[784]), .B(init), .Z(\round_in[0][784] ) );
  AND U10133 ( .A(round_reg[785]), .B(init), .Z(\round_in[0][785] ) );
  AND U10134 ( .A(round_reg[786]), .B(init), .Z(\round_in[0][786] ) );
  AND U10135 ( .A(round_reg[787]), .B(init), .Z(\round_in[0][787] ) );
  AND U10136 ( .A(round_reg[788]), .B(init), .Z(\round_in[0][788] ) );
  AND U10137 ( .A(round_reg[789]), .B(init), .Z(\round_in[0][789] ) );
  NAND U10138 ( .A(init), .B(round_reg[78]), .Z(n3920) );
  NANDN U10139 ( .A(init), .B(in[78]), .Z(n3919) );
  NAND U10140 ( .A(n3920), .B(n3919), .Z(\round_in[0][78] ) );
  AND U10141 ( .A(round_reg[790]), .B(init), .Z(\round_in[0][790] ) );
  AND U10142 ( .A(round_reg[791]), .B(init), .Z(\round_in[0][791] ) );
  AND U10143 ( .A(round_reg[792]), .B(init), .Z(\round_in[0][792] ) );
  AND U10144 ( .A(round_reg[793]), .B(init), .Z(\round_in[0][793] ) );
  AND U10145 ( .A(round_reg[794]), .B(init), .Z(\round_in[0][794] ) );
  AND U10146 ( .A(round_reg[795]), .B(init), .Z(\round_in[0][795] ) );
  AND U10147 ( .A(round_reg[796]), .B(init), .Z(\round_in[0][796] ) );
  AND U10148 ( .A(round_reg[797]), .B(init), .Z(\round_in[0][797] ) );
  AND U10149 ( .A(round_reg[798]), .B(init), .Z(\round_in[0][798] ) );
  AND U10150 ( .A(round_reg[799]), .B(init), .Z(\round_in[0][799] ) );
  NAND U10151 ( .A(init), .B(round_reg[79]), .Z(n3922) );
  NANDN U10152 ( .A(init), .B(in[79]), .Z(n3921) );
  NAND U10153 ( .A(n3922), .B(n3921), .Z(\round_in[0][79] ) );
  NAND U10154 ( .A(init), .B(round_reg[7]), .Z(n3924) );
  NANDN U10155 ( .A(init), .B(in[7]), .Z(n3923) );
  NAND U10156 ( .A(n3924), .B(n3923), .Z(\round_in[0][7] ) );
  AND U10157 ( .A(round_reg[800]), .B(init), .Z(\round_in[0][800] ) );
  AND U10158 ( .A(round_reg[801]), .B(init), .Z(\round_in[0][801] ) );
  AND U10159 ( .A(round_reg[802]), .B(init), .Z(\round_in[0][802] ) );
  AND U10160 ( .A(round_reg[803]), .B(init), .Z(\round_in[0][803] ) );
  AND U10161 ( .A(round_reg[804]), .B(init), .Z(\round_in[0][804] ) );
  AND U10162 ( .A(round_reg[805]), .B(init), .Z(\round_in[0][805] ) );
  AND U10163 ( .A(round_reg[806]), .B(init), .Z(\round_in[0][806] ) );
  AND U10164 ( .A(round_reg[807]), .B(init), .Z(\round_in[0][807] ) );
  AND U10165 ( .A(round_reg[808]), .B(init), .Z(\round_in[0][808] ) );
  AND U10166 ( .A(round_reg[809]), .B(init), .Z(\round_in[0][809] ) );
  NAND U10167 ( .A(init), .B(round_reg[80]), .Z(n3926) );
  NANDN U10168 ( .A(init), .B(in[80]), .Z(n3925) );
  NAND U10169 ( .A(n3926), .B(n3925), .Z(\round_in[0][80] ) );
  AND U10170 ( .A(round_reg[810]), .B(init), .Z(\round_in[0][810] ) );
  AND U10171 ( .A(round_reg[811]), .B(init), .Z(\round_in[0][811] ) );
  AND U10172 ( .A(round_reg[812]), .B(init), .Z(\round_in[0][812] ) );
  AND U10173 ( .A(round_reg[813]), .B(init), .Z(\round_in[0][813] ) );
  AND U10174 ( .A(round_reg[814]), .B(init), .Z(\round_in[0][814] ) );
  AND U10175 ( .A(round_reg[815]), .B(init), .Z(\round_in[0][815] ) );
  AND U10176 ( .A(round_reg[816]), .B(init), .Z(\round_in[0][816] ) );
  AND U10177 ( .A(round_reg[817]), .B(init), .Z(\round_in[0][817] ) );
  AND U10178 ( .A(round_reg[818]), .B(init), .Z(\round_in[0][818] ) );
  AND U10179 ( .A(round_reg[819]), .B(init), .Z(\round_in[0][819] ) );
  NAND U10180 ( .A(init), .B(round_reg[81]), .Z(n3928) );
  NANDN U10181 ( .A(init), .B(in[81]), .Z(n3927) );
  NAND U10182 ( .A(n3928), .B(n3927), .Z(\round_in[0][81] ) );
  AND U10183 ( .A(round_reg[820]), .B(init), .Z(\round_in[0][820] ) );
  AND U10184 ( .A(round_reg[821]), .B(init), .Z(\round_in[0][821] ) );
  AND U10185 ( .A(round_reg[822]), .B(init), .Z(\round_in[0][822] ) );
  AND U10186 ( .A(round_reg[823]), .B(init), .Z(\round_in[0][823] ) );
  AND U10187 ( .A(round_reg[824]), .B(init), .Z(\round_in[0][824] ) );
  AND U10188 ( .A(round_reg[825]), .B(init), .Z(\round_in[0][825] ) );
  AND U10189 ( .A(round_reg[826]), .B(init), .Z(\round_in[0][826] ) );
  AND U10190 ( .A(round_reg[827]), .B(init), .Z(\round_in[0][827] ) );
  AND U10191 ( .A(round_reg[828]), .B(init), .Z(\round_in[0][828] ) );
  AND U10192 ( .A(round_reg[829]), .B(init), .Z(\round_in[0][829] ) );
  NAND U10193 ( .A(init), .B(round_reg[82]), .Z(n3930) );
  NANDN U10194 ( .A(init), .B(in[82]), .Z(n3929) );
  NAND U10195 ( .A(n3930), .B(n3929), .Z(\round_in[0][82] ) );
  AND U10196 ( .A(round_reg[830]), .B(init), .Z(\round_in[0][830] ) );
  AND U10197 ( .A(round_reg[831]), .B(init), .Z(\round_in[0][831] ) );
  AND U10198 ( .A(round_reg[832]), .B(init), .Z(\round_in[0][832] ) );
  AND U10199 ( .A(round_reg[833]), .B(init), .Z(\round_in[0][833] ) );
  AND U10200 ( .A(round_reg[834]), .B(init), .Z(\round_in[0][834] ) );
  AND U10201 ( .A(round_reg[835]), .B(init), .Z(\round_in[0][835] ) );
  AND U10202 ( .A(round_reg[836]), .B(init), .Z(\round_in[0][836] ) );
  AND U10203 ( .A(round_reg[837]), .B(init), .Z(\round_in[0][837] ) );
  AND U10204 ( .A(round_reg[838]), .B(init), .Z(\round_in[0][838] ) );
  AND U10205 ( .A(round_reg[839]), .B(init), .Z(\round_in[0][839] ) );
  NAND U10206 ( .A(init), .B(round_reg[83]), .Z(n3932) );
  NANDN U10207 ( .A(init), .B(in[83]), .Z(n3931) );
  NAND U10208 ( .A(n3932), .B(n3931), .Z(\round_in[0][83] ) );
  AND U10209 ( .A(round_reg[840]), .B(init), .Z(\round_in[0][840] ) );
  AND U10210 ( .A(round_reg[841]), .B(init), .Z(\round_in[0][841] ) );
  AND U10211 ( .A(round_reg[842]), .B(init), .Z(\round_in[0][842] ) );
  AND U10212 ( .A(round_reg[843]), .B(init), .Z(\round_in[0][843] ) );
  AND U10213 ( .A(round_reg[844]), .B(init), .Z(\round_in[0][844] ) );
  AND U10214 ( .A(round_reg[845]), .B(init), .Z(\round_in[0][845] ) );
  AND U10215 ( .A(round_reg[846]), .B(init), .Z(\round_in[0][846] ) );
  AND U10216 ( .A(round_reg[847]), .B(init), .Z(\round_in[0][847] ) );
  AND U10217 ( .A(round_reg[848]), .B(init), .Z(\round_in[0][848] ) );
  AND U10218 ( .A(round_reg[849]), .B(init), .Z(\round_in[0][849] ) );
  NAND U10219 ( .A(init), .B(round_reg[84]), .Z(n3934) );
  NANDN U10220 ( .A(init), .B(in[84]), .Z(n3933) );
  NAND U10221 ( .A(n3934), .B(n3933), .Z(\round_in[0][84] ) );
  AND U10222 ( .A(round_reg[850]), .B(init), .Z(\round_in[0][850] ) );
  AND U10223 ( .A(round_reg[851]), .B(init), .Z(\round_in[0][851] ) );
  AND U10224 ( .A(round_reg[852]), .B(init), .Z(\round_in[0][852] ) );
  AND U10225 ( .A(round_reg[853]), .B(init), .Z(\round_in[0][853] ) );
  AND U10226 ( .A(round_reg[854]), .B(init), .Z(\round_in[0][854] ) );
  AND U10227 ( .A(round_reg[855]), .B(init), .Z(\round_in[0][855] ) );
  AND U10228 ( .A(round_reg[856]), .B(init), .Z(\round_in[0][856] ) );
  AND U10229 ( .A(round_reg[857]), .B(init), .Z(\round_in[0][857] ) );
  AND U10230 ( .A(round_reg[858]), .B(init), .Z(\round_in[0][858] ) );
  AND U10231 ( .A(round_reg[859]), .B(init), .Z(\round_in[0][859] ) );
  NAND U10232 ( .A(init), .B(round_reg[85]), .Z(n3936) );
  NANDN U10233 ( .A(init), .B(in[85]), .Z(n3935) );
  NAND U10234 ( .A(n3936), .B(n3935), .Z(\round_in[0][85] ) );
  AND U10235 ( .A(round_reg[860]), .B(init), .Z(\round_in[0][860] ) );
  AND U10236 ( .A(round_reg[861]), .B(init), .Z(\round_in[0][861] ) );
  AND U10237 ( .A(round_reg[862]), .B(init), .Z(\round_in[0][862] ) );
  AND U10238 ( .A(round_reg[863]), .B(init), .Z(\round_in[0][863] ) );
  AND U10239 ( .A(round_reg[864]), .B(init), .Z(\round_in[0][864] ) );
  AND U10240 ( .A(round_reg[865]), .B(init), .Z(\round_in[0][865] ) );
  AND U10241 ( .A(round_reg[866]), .B(init), .Z(\round_in[0][866] ) );
  AND U10242 ( .A(round_reg[867]), .B(init), .Z(\round_in[0][867] ) );
  AND U10243 ( .A(round_reg[868]), .B(init), .Z(\round_in[0][868] ) );
  AND U10244 ( .A(round_reg[869]), .B(init), .Z(\round_in[0][869] ) );
  NAND U10245 ( .A(init), .B(round_reg[86]), .Z(n3938) );
  NANDN U10246 ( .A(init), .B(in[86]), .Z(n3937) );
  NAND U10247 ( .A(n3938), .B(n3937), .Z(\round_in[0][86] ) );
  AND U10248 ( .A(round_reg[870]), .B(init), .Z(\round_in[0][870] ) );
  AND U10249 ( .A(round_reg[871]), .B(init), .Z(\round_in[0][871] ) );
  AND U10250 ( .A(round_reg[872]), .B(init), .Z(\round_in[0][872] ) );
  AND U10251 ( .A(round_reg[873]), .B(init), .Z(\round_in[0][873] ) );
  AND U10252 ( .A(round_reg[874]), .B(init), .Z(\round_in[0][874] ) );
  AND U10253 ( .A(round_reg[875]), .B(init), .Z(\round_in[0][875] ) );
  AND U10254 ( .A(round_reg[876]), .B(init), .Z(\round_in[0][876] ) );
  AND U10255 ( .A(round_reg[877]), .B(init), .Z(\round_in[0][877] ) );
  AND U10256 ( .A(round_reg[878]), .B(init), .Z(\round_in[0][878] ) );
  AND U10257 ( .A(round_reg[879]), .B(init), .Z(\round_in[0][879] ) );
  NAND U10258 ( .A(init), .B(round_reg[87]), .Z(n3940) );
  NANDN U10259 ( .A(init), .B(in[87]), .Z(n3939) );
  NAND U10260 ( .A(n3940), .B(n3939), .Z(\round_in[0][87] ) );
  AND U10261 ( .A(round_reg[880]), .B(init), .Z(\round_in[0][880] ) );
  AND U10262 ( .A(round_reg[881]), .B(init), .Z(\round_in[0][881] ) );
  AND U10263 ( .A(round_reg[882]), .B(init), .Z(\round_in[0][882] ) );
  AND U10264 ( .A(round_reg[883]), .B(init), .Z(\round_in[0][883] ) );
  AND U10265 ( .A(round_reg[884]), .B(init), .Z(\round_in[0][884] ) );
  AND U10266 ( .A(round_reg[885]), .B(init), .Z(\round_in[0][885] ) );
  AND U10267 ( .A(round_reg[886]), .B(init), .Z(\round_in[0][886] ) );
  AND U10268 ( .A(round_reg[887]), .B(init), .Z(\round_in[0][887] ) );
  AND U10269 ( .A(round_reg[888]), .B(init), .Z(\round_in[0][888] ) );
  AND U10270 ( .A(round_reg[889]), .B(init), .Z(\round_in[0][889] ) );
  NAND U10271 ( .A(init), .B(round_reg[88]), .Z(n3942) );
  NANDN U10272 ( .A(init), .B(in[88]), .Z(n3941) );
  NAND U10273 ( .A(n3942), .B(n3941), .Z(\round_in[0][88] ) );
  AND U10274 ( .A(round_reg[890]), .B(init), .Z(\round_in[0][890] ) );
  AND U10275 ( .A(round_reg[891]), .B(init), .Z(\round_in[0][891] ) );
  AND U10276 ( .A(round_reg[892]), .B(init), .Z(\round_in[0][892] ) );
  AND U10277 ( .A(round_reg[893]), .B(init), .Z(\round_in[0][893] ) );
  AND U10278 ( .A(round_reg[894]), .B(init), .Z(\round_in[0][894] ) );
  AND U10279 ( .A(round_reg[895]), .B(init), .Z(\round_in[0][895] ) );
  AND U10280 ( .A(round_reg[896]), .B(init), .Z(\round_in[0][896] ) );
  AND U10281 ( .A(round_reg[897]), .B(init), .Z(\round_in[0][897] ) );
  AND U10282 ( .A(round_reg[898]), .B(init), .Z(\round_in[0][898] ) );
  AND U10283 ( .A(round_reg[899]), .B(init), .Z(\round_in[0][899] ) );
  NAND U10284 ( .A(init), .B(round_reg[89]), .Z(n3944) );
  NANDN U10285 ( .A(init), .B(in[89]), .Z(n3943) );
  NAND U10286 ( .A(n3944), .B(n3943), .Z(\round_in[0][89] ) );
  NAND U10287 ( .A(init), .B(round_reg[8]), .Z(n3946) );
  NANDN U10288 ( .A(init), .B(in[8]), .Z(n3945) );
  NAND U10289 ( .A(n3946), .B(n3945), .Z(\round_in[0][8] ) );
  AND U10290 ( .A(round_reg[900]), .B(init), .Z(\round_in[0][900] ) );
  AND U10291 ( .A(round_reg[901]), .B(init), .Z(\round_in[0][901] ) );
  AND U10292 ( .A(round_reg[902]), .B(init), .Z(\round_in[0][902] ) );
  AND U10293 ( .A(round_reg[903]), .B(init), .Z(\round_in[0][903] ) );
  AND U10294 ( .A(round_reg[904]), .B(init), .Z(\round_in[0][904] ) );
  AND U10295 ( .A(round_reg[905]), .B(init), .Z(\round_in[0][905] ) );
  AND U10296 ( .A(round_reg[906]), .B(init), .Z(\round_in[0][906] ) );
  AND U10297 ( .A(round_reg[907]), .B(init), .Z(\round_in[0][907] ) );
  AND U10298 ( .A(round_reg[908]), .B(init), .Z(\round_in[0][908] ) );
  AND U10299 ( .A(round_reg[909]), .B(init), .Z(\round_in[0][909] ) );
  NAND U10300 ( .A(init), .B(round_reg[90]), .Z(n3948) );
  NANDN U10301 ( .A(init), .B(in[90]), .Z(n3947) );
  NAND U10302 ( .A(n3948), .B(n3947), .Z(\round_in[0][90] ) );
  AND U10303 ( .A(round_reg[910]), .B(init), .Z(\round_in[0][910] ) );
  AND U10304 ( .A(round_reg[911]), .B(init), .Z(\round_in[0][911] ) );
  AND U10305 ( .A(round_reg[912]), .B(init), .Z(\round_in[0][912] ) );
  AND U10306 ( .A(round_reg[913]), .B(init), .Z(\round_in[0][913] ) );
  AND U10307 ( .A(round_reg[914]), .B(init), .Z(\round_in[0][914] ) );
  AND U10308 ( .A(round_reg[915]), .B(init), .Z(\round_in[0][915] ) );
  AND U10309 ( .A(round_reg[916]), .B(init), .Z(\round_in[0][916] ) );
  AND U10310 ( .A(round_reg[917]), .B(init), .Z(\round_in[0][917] ) );
  AND U10311 ( .A(round_reg[918]), .B(init), .Z(\round_in[0][918] ) );
  AND U10312 ( .A(round_reg[919]), .B(init), .Z(\round_in[0][919] ) );
  NAND U10313 ( .A(init), .B(round_reg[91]), .Z(n3950) );
  NANDN U10314 ( .A(init), .B(in[91]), .Z(n3949) );
  NAND U10315 ( .A(n3950), .B(n3949), .Z(\round_in[0][91] ) );
  AND U10316 ( .A(round_reg[920]), .B(init), .Z(\round_in[0][920] ) );
  AND U10317 ( .A(round_reg[921]), .B(init), .Z(\round_in[0][921] ) );
  AND U10318 ( .A(round_reg[922]), .B(init), .Z(\round_in[0][922] ) );
  AND U10319 ( .A(round_reg[923]), .B(init), .Z(\round_in[0][923] ) );
  AND U10320 ( .A(round_reg[924]), .B(init), .Z(\round_in[0][924] ) );
  AND U10321 ( .A(round_reg[925]), .B(init), .Z(\round_in[0][925] ) );
  AND U10322 ( .A(round_reg[926]), .B(init), .Z(\round_in[0][926] ) );
  AND U10323 ( .A(round_reg[927]), .B(init), .Z(\round_in[0][927] ) );
  AND U10324 ( .A(round_reg[928]), .B(init), .Z(\round_in[0][928] ) );
  AND U10325 ( .A(round_reg[929]), .B(init), .Z(\round_in[0][929] ) );
  NAND U10326 ( .A(init), .B(round_reg[92]), .Z(n3952) );
  NANDN U10327 ( .A(init), .B(in[92]), .Z(n3951) );
  NAND U10328 ( .A(n3952), .B(n3951), .Z(\round_in[0][92] ) );
  AND U10329 ( .A(round_reg[930]), .B(init), .Z(\round_in[0][930] ) );
  AND U10330 ( .A(round_reg[931]), .B(init), .Z(\round_in[0][931] ) );
  AND U10331 ( .A(round_reg[932]), .B(init), .Z(\round_in[0][932] ) );
  AND U10332 ( .A(round_reg[933]), .B(init), .Z(\round_in[0][933] ) );
  AND U10333 ( .A(round_reg[934]), .B(init), .Z(\round_in[0][934] ) );
  AND U10334 ( .A(round_reg[935]), .B(init), .Z(\round_in[0][935] ) );
  AND U10335 ( .A(round_reg[936]), .B(init), .Z(\round_in[0][936] ) );
  AND U10336 ( .A(round_reg[937]), .B(init), .Z(\round_in[0][937] ) );
  AND U10337 ( .A(round_reg[938]), .B(init), .Z(\round_in[0][938] ) );
  AND U10338 ( .A(round_reg[939]), .B(init), .Z(\round_in[0][939] ) );
  NAND U10339 ( .A(init), .B(round_reg[93]), .Z(n3954) );
  NANDN U10340 ( .A(init), .B(in[93]), .Z(n3953) );
  NAND U10341 ( .A(n3954), .B(n3953), .Z(\round_in[0][93] ) );
  AND U10342 ( .A(round_reg[940]), .B(init), .Z(\round_in[0][940] ) );
  AND U10343 ( .A(round_reg[941]), .B(init), .Z(\round_in[0][941] ) );
  AND U10344 ( .A(round_reg[942]), .B(init), .Z(\round_in[0][942] ) );
  AND U10345 ( .A(round_reg[943]), .B(init), .Z(\round_in[0][943] ) );
  AND U10346 ( .A(round_reg[944]), .B(init), .Z(\round_in[0][944] ) );
  AND U10347 ( .A(round_reg[945]), .B(init), .Z(\round_in[0][945] ) );
  AND U10348 ( .A(round_reg[946]), .B(init), .Z(\round_in[0][946] ) );
  AND U10349 ( .A(round_reg[947]), .B(init), .Z(\round_in[0][947] ) );
  AND U10350 ( .A(round_reg[948]), .B(init), .Z(\round_in[0][948] ) );
  AND U10351 ( .A(round_reg[949]), .B(init), .Z(\round_in[0][949] ) );
  NAND U10352 ( .A(init), .B(round_reg[94]), .Z(n3956) );
  NANDN U10353 ( .A(init), .B(in[94]), .Z(n3955) );
  NAND U10354 ( .A(n3956), .B(n3955), .Z(\round_in[0][94] ) );
  AND U10355 ( .A(round_reg[950]), .B(init), .Z(\round_in[0][950] ) );
  AND U10356 ( .A(round_reg[951]), .B(init), .Z(\round_in[0][951] ) );
  AND U10357 ( .A(round_reg[952]), .B(init), .Z(\round_in[0][952] ) );
  AND U10358 ( .A(round_reg[953]), .B(init), .Z(\round_in[0][953] ) );
  AND U10359 ( .A(round_reg[954]), .B(init), .Z(\round_in[0][954] ) );
  AND U10360 ( .A(round_reg[955]), .B(init), .Z(\round_in[0][955] ) );
  AND U10361 ( .A(round_reg[956]), .B(init), .Z(\round_in[0][956] ) );
  AND U10362 ( .A(round_reg[957]), .B(init), .Z(\round_in[0][957] ) );
  AND U10363 ( .A(round_reg[958]), .B(init), .Z(\round_in[0][958] ) );
  AND U10364 ( .A(round_reg[959]), .B(init), .Z(\round_in[0][959] ) );
  NAND U10365 ( .A(init), .B(round_reg[95]), .Z(n3958) );
  NANDN U10366 ( .A(init), .B(in[95]), .Z(n3957) );
  NAND U10367 ( .A(n3958), .B(n3957), .Z(\round_in[0][95] ) );
  AND U10368 ( .A(round_reg[960]), .B(init), .Z(\round_in[0][960] ) );
  AND U10369 ( .A(round_reg[961]), .B(init), .Z(\round_in[0][961] ) );
  AND U10370 ( .A(round_reg[962]), .B(init), .Z(\round_in[0][962] ) );
  AND U10371 ( .A(round_reg[963]), .B(init), .Z(\round_in[0][963] ) );
  AND U10372 ( .A(round_reg[964]), .B(init), .Z(\round_in[0][964] ) );
  AND U10373 ( .A(round_reg[965]), .B(init), .Z(\round_in[0][965] ) );
  AND U10374 ( .A(round_reg[966]), .B(init), .Z(\round_in[0][966] ) );
  AND U10375 ( .A(round_reg[967]), .B(init), .Z(\round_in[0][967] ) );
  AND U10376 ( .A(round_reg[968]), .B(init), .Z(\round_in[0][968] ) );
  AND U10377 ( .A(round_reg[969]), .B(init), .Z(\round_in[0][969] ) );
  NAND U10378 ( .A(init), .B(round_reg[96]), .Z(n3960) );
  NANDN U10379 ( .A(init), .B(in[96]), .Z(n3959) );
  NAND U10380 ( .A(n3960), .B(n3959), .Z(\round_in[0][96] ) );
  AND U10381 ( .A(round_reg[970]), .B(init), .Z(\round_in[0][970] ) );
  AND U10382 ( .A(round_reg[971]), .B(init), .Z(\round_in[0][971] ) );
  AND U10383 ( .A(round_reg[972]), .B(init), .Z(\round_in[0][972] ) );
  AND U10384 ( .A(round_reg[973]), .B(init), .Z(\round_in[0][973] ) );
  AND U10385 ( .A(round_reg[974]), .B(init), .Z(\round_in[0][974] ) );
  AND U10386 ( .A(round_reg[975]), .B(init), .Z(\round_in[0][975] ) );
  AND U10387 ( .A(round_reg[976]), .B(init), .Z(\round_in[0][976] ) );
  AND U10388 ( .A(round_reg[977]), .B(init), .Z(\round_in[0][977] ) );
  AND U10389 ( .A(round_reg[978]), .B(init), .Z(\round_in[0][978] ) );
  AND U10390 ( .A(round_reg[979]), .B(init), .Z(\round_in[0][979] ) );
  NAND U10391 ( .A(init), .B(round_reg[97]), .Z(n3962) );
  NANDN U10392 ( .A(init), .B(in[97]), .Z(n3961) );
  NAND U10393 ( .A(n3962), .B(n3961), .Z(\round_in[0][97] ) );
  AND U10394 ( .A(round_reg[980]), .B(init), .Z(\round_in[0][980] ) );
  AND U10395 ( .A(round_reg[981]), .B(init), .Z(\round_in[0][981] ) );
  AND U10396 ( .A(round_reg[982]), .B(init), .Z(\round_in[0][982] ) );
  AND U10397 ( .A(round_reg[983]), .B(init), .Z(\round_in[0][983] ) );
  AND U10398 ( .A(round_reg[984]), .B(init), .Z(\round_in[0][984] ) );
  AND U10399 ( .A(round_reg[985]), .B(init), .Z(\round_in[0][985] ) );
  AND U10400 ( .A(round_reg[986]), .B(init), .Z(\round_in[0][986] ) );
  AND U10401 ( .A(round_reg[987]), .B(init), .Z(\round_in[0][987] ) );
  AND U10402 ( .A(round_reg[988]), .B(init), .Z(\round_in[0][988] ) );
  AND U10403 ( .A(round_reg[989]), .B(init), .Z(\round_in[0][989] ) );
  NAND U10404 ( .A(init), .B(round_reg[98]), .Z(n3964) );
  NANDN U10405 ( .A(init), .B(in[98]), .Z(n3963) );
  NAND U10406 ( .A(n3964), .B(n3963), .Z(\round_in[0][98] ) );
  AND U10407 ( .A(round_reg[990]), .B(init), .Z(\round_in[0][990] ) );
  AND U10408 ( .A(round_reg[991]), .B(init), .Z(\round_in[0][991] ) );
  AND U10409 ( .A(round_reg[992]), .B(init), .Z(\round_in[0][992] ) );
  AND U10410 ( .A(round_reg[993]), .B(init), .Z(\round_in[0][993] ) );
  AND U10411 ( .A(round_reg[994]), .B(init), .Z(\round_in[0][994] ) );
  AND U10412 ( .A(round_reg[995]), .B(init), .Z(\round_in[0][995] ) );
  AND U10413 ( .A(round_reg[996]), .B(init), .Z(\round_in[0][996] ) );
  AND U10414 ( .A(round_reg[997]), .B(init), .Z(\round_in[0][997] ) );
  AND U10415 ( .A(round_reg[998]), .B(init), .Z(\round_in[0][998] ) );
  AND U10416 ( .A(round_reg[999]), .B(init), .Z(\round_in[0][999] ) );
  NAND U10417 ( .A(init), .B(round_reg[99]), .Z(n3966) );
  NANDN U10418 ( .A(init), .B(in[99]), .Z(n3965) );
  NAND U10419 ( .A(n3966), .B(n3965), .Z(\round_in[0][99] ) );
  NAND U10420 ( .A(init), .B(round_reg[9]), .Z(n3968) );
  NANDN U10421 ( .A(init), .B(in[9]), .Z(n3967) );
  NAND U10422 ( .A(n3968), .B(n3967), .Z(\round_in[0][9] ) );
endmodule

