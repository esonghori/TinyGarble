
module modexp_2N_NN_N4_CC8 ( clk, rst, m, e, n, c );
  input [3:0] m;
  input [3:0] e;
  input [3:0] n;
  output [3:0] c;
  input clk, rst;
  wire   init, mul_pow, first_one, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594;
  wire   [3:0] ereg;
  wire   [3:0] creg;

  DFF init_reg ( .D(1'b1), .CLK(clk), .RST(rst), .Q(init) );
  DFF mul_pow_reg ( .D(n43), .CLK(clk), .RST(rst), .Q(mul_pow) );
  DFF \ereg_reg[0]  ( .D(n42), .CLK(clk), .RST(rst), .Q(ereg[0]) );
  DFF \ereg_reg[1]  ( .D(n41), .CLK(clk), .RST(rst), .Q(ereg[1]) );
  DFF \ereg_reg[2]  ( .D(n40), .CLK(clk), .RST(rst), .Q(ereg[2]) );
  DFF \ereg_reg[3]  ( .D(n39), .CLK(clk), .RST(rst), .Q(ereg[3]) );
  DFF first_one_reg ( .D(n38), .CLK(clk), .RST(rst), .Q(first_one) );
  DFF \creg_reg[3]  ( .D(n37), .CLK(clk), .RST(rst), .Q(creg[3]) );
  DFF \creg_reg[2]  ( .D(n36), .CLK(clk), .RST(rst), .Q(creg[2]) );
  DFF \creg_reg[1]  ( .D(n35), .CLK(clk), .RST(rst), .Q(creg[1]) );
  DFF \creg_reg[0]  ( .D(n34), .CLK(clk), .RST(rst), .Q(creg[0]) );
  NAND U209 ( .A(n259), .B(n[1]), .Z(n152) );
  XOR U210 ( .A(n259), .B(n[1]), .Z(n153) );
  NANDN U211 ( .A(n262), .B(n153), .Z(n154) );
  NAND U212 ( .A(n152), .B(n154), .Z(n251) );
  ANDN U213 ( .B(n364), .A(n363), .Z(n155) );
  AND U214 ( .A(n[0]), .B(n155), .Z(n156) );
  NAND U215 ( .A(n357), .B(n[1]), .Z(n157) );
  XOR U216 ( .A(n357), .B(n[1]), .Z(n158) );
  NAND U217 ( .A(n158), .B(n156), .Z(n159) );
  NAND U218 ( .A(n157), .B(n159), .Z(n160) );
  XOR U219 ( .A(n[2]), .B(n378), .Z(n161) );
  NAND U220 ( .A(n161), .B(n160), .Z(n162) );
  NAND U221 ( .A(n[2]), .B(n378), .Z(n163) );
  AND U222 ( .A(n162), .B(n163), .Z(n164) );
  NANDN U223 ( .A(n394), .B(n346), .Z(n165) );
  NAND U224 ( .A(n388), .B(n522), .Z(n166) );
  ANDN U225 ( .B(n166), .A(n165), .Z(n167) );
  XOR U226 ( .A(n388), .B(n522), .Z(n168) );
  NAND U227 ( .A(n168), .B(n164), .Z(n169) );
  NAND U228 ( .A(n167), .B(n169), .Z(n384) );
  NAND U229 ( .A(n512), .B(n[1]), .Z(n170) );
  XOR U230 ( .A(n512), .B(n[1]), .Z(n171) );
  NAND U231 ( .A(n171), .B(n509), .Z(n172) );
  NAND U232 ( .A(n170), .B(n172), .Z(n516) );
  XOR U233 ( .A(n481), .B(n482), .Z(n520) );
  XOR U234 ( .A(n263), .B(n265), .Z(n173) );
  AND U235 ( .A(n[0]), .B(n173), .Z(n174) );
  NAND U236 ( .A(n174), .B(n[1]), .Z(n175) );
  XOR U237 ( .A(n174), .B(n[1]), .Z(n176) );
  NANDN U238 ( .A(n281), .B(n176), .Z(n177) );
  NAND U239 ( .A(n175), .B(n177), .Z(n178) );
  NAND U240 ( .A(n296), .B(n[2]), .Z(n179) );
  XOR U241 ( .A(n296), .B(n[2]), .Z(n180) );
  NAND U242 ( .A(n180), .B(n178), .Z(n181) );
  NAND U243 ( .A(n179), .B(n181), .Z(n302) );
  XOR U244 ( .A(n360), .B(n361), .Z(n401) );
  NAND U245 ( .A(n439), .B(n[1]), .Z(n182) );
  XOR U246 ( .A(n439), .B(n[1]), .Z(n183) );
  NAND U247 ( .A(n183), .B(n435), .Z(n184) );
  NAND U248 ( .A(n182), .B(n184), .Z(n431) );
  XOR U249 ( .A(n391), .B(n392), .Z(n429) );
  AND U250 ( .A(n[0]), .B(n530), .Z(n185) );
  NAND U251 ( .A(n537), .B(n[1]), .Z(n186) );
  XOR U252 ( .A(n537), .B(n[1]), .Z(n187) );
  NAND U253 ( .A(n187), .B(n185), .Z(n188) );
  NAND U254 ( .A(n186), .B(n188), .Z(n189) );
  XOR U255 ( .A(n[2]), .B(n542), .Z(n190) );
  NAND U256 ( .A(n190), .B(n189), .Z(n191) );
  NAND U257 ( .A(n[2]), .B(n542), .Z(n192) );
  AND U258 ( .A(n191), .B(n192), .Z(n193) );
  AND U259 ( .A(n[3]), .B(n525), .Z(n194) );
  NANDN U260 ( .A(n523), .B(n527), .Z(n195) );
  AND U261 ( .A(n194), .B(n195), .Z(n196) );
  XNOR U262 ( .A(n520), .B(n196), .Z(n197) );
  NANDN U263 ( .A(n521), .B(n197), .Z(n198) );
  NAND U264 ( .A(n550), .B(n522), .Z(n199) );
  ANDN U265 ( .B(n199), .A(n198), .Z(n200) );
  XOR U266 ( .A(n550), .B(n522), .Z(n201) );
  NAND U267 ( .A(n201), .B(n193), .Z(n202) );
  NAND U268 ( .A(n200), .B(n202), .Z(n546) );
  ANDN U269 ( .B(n274), .A(n272), .Z(n284) );
  NAND U270 ( .A(n350), .B(n[1]), .Z(n203) );
  XOR U271 ( .A(n350), .B(n[1]), .Z(n204) );
  NAND U272 ( .A(n204), .B(n347), .Z(n205) );
  NAND U273 ( .A(n203), .B(n205), .Z(n333) );
  XOR U274 ( .A(n307), .B(n305), .Z(n206) );
  XNOR U275 ( .A(n306), .B(n206), .Z(n345) );
  ANDN U276 ( .B(n443), .A(n442), .Z(n207) );
  AND U277 ( .A(n[0]), .B(n207), .Z(n208) );
  NAND U278 ( .A(n451), .B(n[1]), .Z(n209) );
  XOR U279 ( .A(n451), .B(n[1]), .Z(n210) );
  NAND U280 ( .A(n210), .B(n208), .Z(n211) );
  NAND U281 ( .A(n209), .B(n211), .Z(n212) );
  XOR U282 ( .A(n[2]), .B(n468), .Z(n213) );
  NAND U283 ( .A(n213), .B(n212), .Z(n214) );
  NAND U284 ( .A(n[2]), .B(n468), .Z(n215) );
  AND U285 ( .A(n214), .B(n215), .Z(n216) );
  OR U286 ( .A(n484), .B(n430), .Z(n217) );
  NAND U287 ( .A(n478), .B(n522), .Z(n218) );
  ANDN U288 ( .B(n218), .A(n217), .Z(n219) );
  XOR U289 ( .A(n478), .B(n522), .Z(n220) );
  NAND U290 ( .A(n220), .B(n216), .Z(n221) );
  NAND U291 ( .A(n219), .B(n221), .Z(n474) );
  XOR U292 ( .A(n537), .B(n535), .Z(n222) );
  NANDN U293 ( .A(n536), .B(n222), .Z(n223) );
  NAND U294 ( .A(n537), .B(n535), .Z(n224) );
  AND U295 ( .A(n223), .B(n224), .Z(n543) );
  IV U296 ( .A(n[2]), .Z(n225) );
  NANDN U297 ( .A(init), .B(e[3]), .Z(n581) );
  NAND U298 ( .A(ereg[3]), .B(init), .Z(n226) );
  AND U299 ( .A(n581), .B(n226), .Z(n551) );
  NAND U300 ( .A(creg[0]), .B(n551), .Z(n529) );
  IV U301 ( .A(n[3]), .Z(n522) );
  IV U302 ( .A(mul_pow), .Z(n43) );
  AND U303 ( .A(init), .B(n43), .Z(n592) );
  NAND U304 ( .A(creg[0]), .B(n592), .Z(n228) );
  NANDN U305 ( .A(n592), .B(m[0]), .Z(n227) );
  NAND U306 ( .A(n228), .B(n227), .Z(n505) );
  NANDN U307 ( .A(init), .B(m[1]), .Z(n564) );
  NAND U308 ( .A(creg[1]), .B(init), .Z(n229) );
  AND U309 ( .A(n564), .B(n229), .Z(n399) );
  ANDN U310 ( .B(n505), .A(n399), .Z(n416) );
  NANDN U311 ( .A(init), .B(m[3]), .Z(n576) );
  NAND U312 ( .A(init), .B(creg[3]), .Z(n230) );
  AND U313 ( .A(n576), .B(n230), .Z(n244) );
  NANDN U314 ( .A(n244), .B(n505), .Z(n263) );
  NOR U315 ( .A(n263), .B(n[0]), .Z(n273) );
  NANDN U316 ( .A(n273), .B(n[1]), .Z(n235) );
  NAND U317 ( .A(creg[1]), .B(n592), .Z(n232) );
  NANDN U318 ( .A(n592), .B(m[1]), .Z(n231) );
  NAND U319 ( .A(n232), .B(n231), .Z(n446) );
  ANDN U320 ( .B(n446), .A(n244), .Z(n262) );
  XNOR U321 ( .A(n273), .B(n[1]), .Z(n233) );
  NANDN U322 ( .A(n262), .B(n233), .Z(n234) );
  NAND U323 ( .A(n235), .B(n234), .Z(n238) );
  NAND U324 ( .A(n[2]), .B(n238), .Z(n241) );
  NAND U325 ( .A(creg[2]), .B(n592), .Z(n237) );
  NANDN U326 ( .A(n592), .B(m[2]), .Z(n236) );
  NAND U327 ( .A(n237), .B(n236), .Z(n459) );
  ANDN U328 ( .B(n459), .A(n244), .Z(n267) );
  IV U329 ( .A(n267), .Z(n252) );
  XOR U330 ( .A(n238), .B(n[2]), .Z(n239) );
  NAND U331 ( .A(n252), .B(n239), .Z(n240) );
  NAND U332 ( .A(n241), .B(n240), .Z(n246) );
  XOR U333 ( .A(n[3]), .B(n246), .Z(n245) );
  NAND U334 ( .A(creg[3]), .B(n592), .Z(n243) );
  NANDN U335 ( .A(n592), .B(m[3]), .Z(n242) );
  NAND U336 ( .A(n243), .B(n242), .Z(n456) );
  NANDN U337 ( .A(n244), .B(n456), .Z(n257) );
  NAND U338 ( .A(n245), .B(n257), .Z(n248) );
  NAND U339 ( .A(n[3]), .B(n246), .Z(n247) );
  AND U340 ( .A(n248), .B(n247), .Z(n265) );
  XNOR U341 ( .A(n263), .B(n265), .Z(n250) );
  NANDN U342 ( .A(n[0]), .B(n263), .Z(n249) );
  NAND U343 ( .A(n250), .B(n249), .Z(n274) );
  AND U344 ( .A(n[0]), .B(n263), .Z(n259) );
  NAND U345 ( .A(n[2]), .B(n251), .Z(n254) );
  XOR U346 ( .A(n251), .B(n[2]), .Z(n264) );
  NAND U347 ( .A(n252), .B(n264), .Z(n253) );
  NAND U348 ( .A(n254), .B(n253), .Z(n255) );
  OR U349 ( .A(n255), .B(n[3]), .Z(n256) );
  NAND U350 ( .A(n265), .B(n256), .Z(n258) );
  ANDN U351 ( .B(n258), .A(n257), .Z(n304) );
  XOR U352 ( .A(n[1]), .B(n259), .Z(n260) );
  NAND U353 ( .A(n265), .B(n260), .Z(n261) );
  XNOR U354 ( .A(n262), .B(n261), .Z(n281) );
  AND U355 ( .A(n265), .B(n264), .Z(n266) );
  XOR U356 ( .A(n267), .B(n266), .Z(n280) );
  IV U357 ( .A(n280), .Z(n296) );
  XOR U358 ( .A(n[3]), .B(n302), .Z(n268) );
  NANDN U359 ( .A(n304), .B(n268), .Z(n270) );
  NAND U360 ( .A(n[3]), .B(n302), .Z(n269) );
  AND U361 ( .A(n270), .B(n269), .Z(n279) );
  NAND U362 ( .A(n[0]), .B(n279), .Z(n272) );
  AND U363 ( .A(n[1]), .B(n279), .Z(n282) );
  XNOR U364 ( .A(n281), .B(n282), .Z(n283) );
  XNOR U365 ( .A(n284), .B(n283), .Z(n287) );
  NANDN U366 ( .A(init), .B(m[2]), .Z(n569) );
  NAND U367 ( .A(init), .B(creg[2]), .Z(n271) );
  AND U368 ( .A(n569), .B(n271), .Z(n310) );
  XNOR U369 ( .A(n274), .B(n272), .Z(n276) );
  NAND U370 ( .A(n274), .B(n273), .Z(n275) );
  NAND U371 ( .A(n276), .B(n275), .Z(n319) );
  AND U372 ( .A(n319), .B(n446), .Z(n288) );
  XOR U373 ( .A(n459), .B(n288), .Z(n277) );
  NANDN U374 ( .A(n310), .B(n277), .Z(n278) );
  XNOR U375 ( .A(n287), .B(n278), .Z(n331) );
  AND U376 ( .A(n279), .B(n[2]), .Z(n297) );
  XNOR U377 ( .A(n280), .B(n297), .Z(n299) );
  NANDN U378 ( .A(n282), .B(n281), .Z(n286) );
  NANDN U379 ( .A(n284), .B(n283), .Z(n285) );
  NAND U380 ( .A(n286), .B(n285), .Z(n298) );
  XOR U381 ( .A(n299), .B(n298), .Z(n314) );
  AND U382 ( .A(n314), .B(n456), .Z(n294) );
  IV U383 ( .A(n456), .Z(n496) );
  XNOR U384 ( .A(n496), .B(n314), .Z(n292) );
  NAND U385 ( .A(n459), .B(n287), .Z(n291) );
  IV U386 ( .A(n459), .Z(n457) );
  XNOR U387 ( .A(n457), .B(n287), .Z(n289) );
  NAND U388 ( .A(n289), .B(n288), .Z(n290) );
  AND U389 ( .A(n291), .B(n290), .Z(n311) );
  ANDN U390 ( .B(n292), .A(n311), .Z(n293) );
  OR U391 ( .A(n294), .B(n293), .Z(n295) );
  ANDN U392 ( .B(n295), .A(n310), .Z(n307) );
  OR U393 ( .A(n297), .B(n296), .Z(n301) );
  NAND U394 ( .A(n299), .B(n298), .Z(n300) );
  NAND U395 ( .A(n301), .B(n300), .Z(n305) );
  NANDN U396 ( .A(n302), .B(n[3]), .Z(n303) );
  AND U397 ( .A(n304), .B(n303), .Z(n306) );
  XNOR U398 ( .A(n305), .B(n307), .Z(n309) );
  XNOR U399 ( .A(n307), .B(n306), .Z(n308) );
  NAND U400 ( .A(n309), .B(n308), .Z(n346) );
  IV U401 ( .A(n310), .Z(n317) );
  XOR U402 ( .A(n496), .B(n311), .Z(n312) );
  NAND U403 ( .A(n317), .B(n312), .Z(n313) );
  XNOR U404 ( .A(n314), .B(n313), .Z(n338) );
  ANDN U405 ( .B(n338), .A(n[3]), .Z(n340) );
  ANDN U406 ( .B(n346), .A(n340), .Z(n327) );
  AND U407 ( .A(n505), .B(n317), .Z(n352) );
  ANDN U408 ( .B(n352), .A(n[0]), .Z(n363) );
  NANDN U409 ( .A(n[1]), .B(n363), .Z(n316) );
  ANDN U410 ( .B(n331), .A(n[2]), .Z(n315) );
  ANDN U411 ( .B(n316), .A(n315), .Z(n322) );
  IV U412 ( .A(n446), .Z(n487) );
  ANDN U413 ( .B(n317), .A(n487), .Z(n318) );
  XNOR U414 ( .A(n319), .B(n318), .Z(n350) );
  XNOR U415 ( .A(n363), .B(n[1]), .Z(n320) );
  NANDN U416 ( .A(n350), .B(n320), .Z(n321) );
  NAND U417 ( .A(n322), .B(n321), .Z(n325) );
  ANDN U418 ( .B(n522), .A(n[2]), .Z(n492) );
  ANDN U419 ( .B(n[3]), .A(n338), .Z(n342) );
  NANDN U420 ( .A(n342), .B(n331), .Z(n323) );
  NANDN U421 ( .A(n492), .B(n323), .Z(n324) );
  AND U422 ( .A(n325), .B(n324), .Z(n326) );
  ANDN U423 ( .B(n327), .A(n326), .Z(n328) );
  NANDN U424 ( .A(n345), .B(n328), .Z(n351) );
  ANDN U425 ( .B(n[0]), .A(n352), .Z(n347) );
  XOR U426 ( .A(n[2]), .B(n333), .Z(n329) );
  NAND U427 ( .A(n351), .B(n329), .Z(n330) );
  XNOR U428 ( .A(n331), .B(n330), .Z(n355) );
  NAND U429 ( .A(n225), .B(n331), .Z(n335) );
  XOR U430 ( .A(n225), .B(n331), .Z(n332) );
  NANDN U431 ( .A(n333), .B(n332), .Z(n334) );
  AND U432 ( .A(n335), .B(n334), .Z(n339) );
  XNOR U433 ( .A(n522), .B(n339), .Z(n336) );
  NAND U434 ( .A(n351), .B(n336), .Z(n337) );
  XNOR U435 ( .A(n338), .B(n337), .Z(n388) );
  NANDN U436 ( .A(n340), .B(n339), .Z(n341) );
  NANDN U437 ( .A(n342), .B(n341), .Z(n343) );
  AND U438 ( .A(n351), .B(n343), .Z(n344) );
  XOR U439 ( .A(n345), .B(n344), .Z(n394) );
  IV U440 ( .A(n355), .Z(n378) );
  XOR U441 ( .A(n[1]), .B(n347), .Z(n348) );
  NAND U442 ( .A(n351), .B(n348), .Z(n349) );
  XNOR U443 ( .A(n350), .B(n349), .Z(n357) );
  XOR U444 ( .A(n352), .B(n351), .Z(n354) );
  OR U445 ( .A(n[0]), .B(n352), .Z(n353) );
  NAND U446 ( .A(n354), .B(n353), .Z(n364) );
  AND U447 ( .A(n384), .B(n[2]), .Z(n379) );
  XNOR U448 ( .A(n355), .B(n379), .Z(n381) );
  NAND U449 ( .A(n[1]), .B(n384), .Z(n356) );
  NANDN U450 ( .A(n357), .B(n356), .Z(n359) );
  NAND U451 ( .A(n[0]), .B(n384), .Z(n362) );
  NANDN U452 ( .A(n362), .B(n364), .Z(n360) );
  XNOR U453 ( .A(n357), .B(n356), .Z(n361) );
  NAND U454 ( .A(n360), .B(n361), .Z(n358) );
  NAND U455 ( .A(n359), .B(n358), .Z(n380) );
  XOR U456 ( .A(n381), .B(n380), .Z(n372) );
  NAND U457 ( .A(n459), .B(n401), .Z(n369) );
  XNOR U458 ( .A(n457), .B(n401), .Z(n367) );
  XNOR U459 ( .A(n364), .B(n362), .Z(n366) );
  NAND U460 ( .A(n364), .B(n363), .Z(n365) );
  NAND U461 ( .A(n366), .B(n365), .Z(n405) );
  AND U462 ( .A(n405), .B(n446), .Z(n397) );
  NAND U463 ( .A(n367), .B(n397), .Z(n368) );
  AND U464 ( .A(n369), .B(n368), .Z(n373) );
  XOR U465 ( .A(n496), .B(n373), .Z(n370) );
  NANDN U466 ( .A(n399), .B(n370), .Z(n371) );
  XNOR U467 ( .A(n372), .B(n371), .Z(n422) );
  ANDN U468 ( .B(n422), .A(n[3]), .Z(n424) );
  AND U469 ( .A(n372), .B(n456), .Z(n376) );
  XNOR U470 ( .A(n496), .B(n372), .Z(n374) );
  ANDN U471 ( .B(n374), .A(n373), .Z(n375) );
  OR U472 ( .A(n376), .B(n375), .Z(n377) );
  IV U473 ( .A(n399), .Z(n403) );
  AND U474 ( .A(n377), .B(n403), .Z(n392) );
  OR U475 ( .A(n379), .B(n378), .Z(n383) );
  NAND U476 ( .A(n381), .B(n380), .Z(n382) );
  NAND U477 ( .A(n383), .B(n382), .Z(n385) );
  NAND U478 ( .A(n[3]), .B(n384), .Z(n387) );
  XOR U479 ( .A(n388), .B(n387), .Z(n386) );
  XOR U480 ( .A(n385), .B(n386), .Z(n391) );
  NAND U481 ( .A(n386), .B(n385), .Z(n390) );
  NAND U482 ( .A(n388), .B(n387), .Z(n389) );
  AND U483 ( .A(n390), .B(n389), .Z(n396) );
  AND U484 ( .A(n392), .B(n391), .Z(n393) );
  XNOR U485 ( .A(n394), .B(n393), .Z(n395) );
  XNOR U486 ( .A(n396), .B(n395), .Z(n430) );
  NOR U487 ( .A(n429), .B(n430), .Z(n412) );
  XOR U488 ( .A(n459), .B(n397), .Z(n398) );
  NANDN U489 ( .A(n399), .B(n398), .Z(n400) );
  XOR U490 ( .A(n401), .B(n400), .Z(n434) );
  ANDN U491 ( .B(n[3]), .A(n422), .Z(n426) );
  OR U492 ( .A(n434), .B(n426), .Z(n402) );
  NANDN U493 ( .A(n492), .B(n402), .Z(n410) );
  OR U494 ( .A(n434), .B(n[2]), .Z(n408) );
  ANDN U495 ( .B(n403), .A(n487), .Z(n404) );
  XNOR U496 ( .A(n405), .B(n404), .Z(n439) );
  ANDN U497 ( .B(n416), .A(n[0]), .Z(n442) );
  NANDN U498 ( .A(n442), .B(n[1]), .Z(n406) );
  NANDN U499 ( .A(n439), .B(n406), .Z(n407) );
  AND U500 ( .A(n408), .B(n407), .Z(n409) );
  ANDN U501 ( .B(n410), .A(n409), .Z(n411) );
  ANDN U502 ( .B(n412), .A(n411), .Z(n413) );
  NANDN U503 ( .A(n424), .B(n413), .Z(n437) );
  XOR U504 ( .A(n416), .B(n437), .Z(n415) );
  OR U505 ( .A(n[0]), .B(n416), .Z(n414) );
  NAND U506 ( .A(n415), .B(n414), .Z(n443) );
  NAND U507 ( .A(n[2]), .B(n434), .Z(n419) );
  XOR U508 ( .A(n434), .B(n[2]), .Z(n417) );
  ANDN U509 ( .B(n[0]), .A(n416), .Z(n435) );
  NAND U510 ( .A(n417), .B(n431), .Z(n418) );
  NAND U511 ( .A(n419), .B(n418), .Z(n423) );
  XOR U512 ( .A(n[3]), .B(n423), .Z(n420) );
  NAND U513 ( .A(n437), .B(n420), .Z(n421) );
  XNOR U514 ( .A(n422), .B(n421), .Z(n478) );
  NANDN U515 ( .A(n424), .B(n423), .Z(n425) );
  NANDN U516 ( .A(n426), .B(n425), .Z(n427) );
  AND U517 ( .A(n437), .B(n427), .Z(n428) );
  XOR U518 ( .A(n429), .B(n428), .Z(n484) );
  XOR U519 ( .A(n[2]), .B(n431), .Z(n432) );
  NAND U520 ( .A(n437), .B(n432), .Z(n433) );
  XNOR U521 ( .A(n434), .B(n433), .Z(n468) );
  XOR U522 ( .A(n[1]), .B(n435), .Z(n436) );
  NAND U523 ( .A(n437), .B(n436), .Z(n438) );
  XNOR U524 ( .A(n439), .B(n438), .Z(n451) );
  AND U525 ( .A(n[0]), .B(n474), .Z(n441) );
  AND U526 ( .A(n443), .B(n441), .Z(n453) );
  AND U527 ( .A(n[1]), .B(n474), .Z(n450) );
  XOR U528 ( .A(n451), .B(n450), .Z(n452) );
  XOR U529 ( .A(n453), .B(n452), .Z(n458) );
  NANDN U530 ( .A(init), .B(m[0]), .Z(n559) );
  NAND U531 ( .A(creg[0]), .B(init), .Z(n440) );
  AND U532 ( .A(n559), .B(n440), .Z(n506) );
  XOR U533 ( .A(n443), .B(n441), .Z(n445) );
  NAND U534 ( .A(n443), .B(n442), .Z(n444) );
  NAND U535 ( .A(n445), .B(n444), .Z(n489) );
  AND U536 ( .A(n489), .B(n446), .Z(n461) );
  XOR U537 ( .A(n459), .B(n461), .Z(n447) );
  NANDN U538 ( .A(n506), .B(n447), .Z(n448) );
  XNOR U539 ( .A(n458), .B(n448), .Z(n515) );
  NAND U540 ( .A(n[2]), .B(n474), .Z(n449) );
  XNOR U541 ( .A(n468), .B(n449), .Z(n471) );
  OR U542 ( .A(n451), .B(n450), .Z(n455) );
  NANDN U543 ( .A(n453), .B(n452), .Z(n454) );
  NAND U544 ( .A(n455), .B(n454), .Z(n470) );
  XOR U545 ( .A(n471), .B(n470), .Z(n499) );
  AND U546 ( .A(n499), .B(n456), .Z(n466) );
  XNOR U547 ( .A(n496), .B(n499), .Z(n464) );
  OR U548 ( .A(n458), .B(n457), .Z(n463) );
  XNOR U549 ( .A(n459), .B(n458), .Z(n460) );
  NAND U550 ( .A(n461), .B(n460), .Z(n462) );
  AND U551 ( .A(n463), .B(n462), .Z(n495) );
  ANDN U552 ( .B(n464), .A(n495), .Z(n465) );
  OR U553 ( .A(n466), .B(n465), .Z(n467) );
  ANDN U554 ( .B(n467), .A(n506), .Z(n482) );
  NANDN U555 ( .A(n225), .B(n474), .Z(n469) );
  ANDN U556 ( .B(n469), .A(n468), .Z(n473) );
  NAND U557 ( .A(n471), .B(n470), .Z(n472) );
  NANDN U558 ( .A(n473), .B(n472), .Z(n475) );
  NAND U559 ( .A(n[3]), .B(n474), .Z(n477) );
  XOR U560 ( .A(n478), .B(n477), .Z(n476) );
  XOR U561 ( .A(n475), .B(n476), .Z(n481) );
  NAND U562 ( .A(n476), .B(n475), .Z(n480) );
  NAND U563 ( .A(n478), .B(n477), .Z(n479) );
  AND U564 ( .A(n480), .B(n479), .Z(n486) );
  AND U565 ( .A(n482), .B(n481), .Z(n483) );
  XNOR U566 ( .A(n484), .B(n483), .Z(n485) );
  XNOR U567 ( .A(n486), .B(n485), .Z(n521) );
  NOR U568 ( .A(n520), .B(n521), .Z(n494) );
  OR U569 ( .A(n515), .B(n[2]), .Z(n491) );
  NOR U570 ( .A(n487), .B(n506), .Z(n488) );
  XNOR U571 ( .A(n489), .B(n488), .Z(n512) );
  OR U572 ( .A(n[1]), .B(n512), .Z(n490) );
  AND U573 ( .A(n491), .B(n490), .Z(n500) );
  NANDN U574 ( .A(n500), .B(n492), .Z(n493) );
  AND U575 ( .A(n494), .B(n493), .Z(n504) );
  XOR U576 ( .A(n496), .B(n495), .Z(n497) );
  NANDN U577 ( .A(n506), .B(n497), .Z(n498) );
  XNOR U578 ( .A(n499), .B(n498), .Z(n527) );
  OR U579 ( .A(n515), .B(n500), .Z(n501) );
  NAND U580 ( .A(n[3]), .B(n501), .Z(n502) );
  NAND U581 ( .A(n527), .B(n502), .Z(n503) );
  NAND U582 ( .A(n504), .B(n503), .Z(n525) );
  NANDN U583 ( .A(n506), .B(n505), .Z(n514) );
  AND U584 ( .A(n[0]), .B(n514), .Z(n509) );
  XOR U585 ( .A(n[2]), .B(n516), .Z(n507) );
  NAND U586 ( .A(n525), .B(n507), .Z(n508) );
  XNOR U587 ( .A(n515), .B(n508), .Z(n542) );
  XOR U588 ( .A(n[1]), .B(n509), .Z(n510) );
  NAND U589 ( .A(n525), .B(n510), .Z(n511) );
  XNOR U590 ( .A(n512), .B(n511), .Z(n537) );
  NAND U591 ( .A(n525), .B(n[0]), .Z(n513) );
  XNOR U592 ( .A(n514), .B(n513), .Z(n530) );
  NAND U593 ( .A(n[2]), .B(n515), .Z(n519) );
  XOR U594 ( .A(n515), .B(n[2]), .Z(n517) );
  NAND U595 ( .A(n517), .B(n516), .Z(n518) );
  NAND U596 ( .A(n519), .B(n518), .Z(n523) );
  XOR U597 ( .A(n[3]), .B(n523), .Z(n524) );
  NAND U598 ( .A(n525), .B(n524), .Z(n526) );
  XNOR U599 ( .A(n527), .B(n526), .Z(n550) );
  AND U600 ( .A(n[0]), .B(n546), .Z(n531) );
  XNOR U601 ( .A(n531), .B(n530), .Z(n556) );
  NANDN U602 ( .A(n551), .B(n556), .Z(n528) );
  NAND U603 ( .A(n529), .B(n528), .Z(c[0]) );
  NAND U604 ( .A(creg[1]), .B(n551), .Z(n534) );
  AND U605 ( .A(n[1]), .B(n546), .Z(n535) );
  NAND U606 ( .A(n531), .B(n530), .Z(n536) );
  XOR U607 ( .A(n537), .B(n536), .Z(n532) );
  XOR U608 ( .A(n535), .B(n532), .Z(n561) );
  NANDN U609 ( .A(n551), .B(n561), .Z(n533) );
  NAND U610 ( .A(n534), .B(n533), .Z(c[1]) );
  NAND U611 ( .A(creg[2]), .B(n551), .Z(n539) );
  XNOR U612 ( .A(n542), .B(n543), .Z(n541) );
  AND U613 ( .A(n546), .B(n[2]), .Z(n540) );
  XNOR U614 ( .A(n541), .B(n540), .Z(n566) );
  NANDN U615 ( .A(n551), .B(n566), .Z(n538) );
  NAND U616 ( .A(n539), .B(n538), .Z(c[2]) );
  NAND U617 ( .A(creg[3]), .B(n551), .Z(n553) );
  NAND U618 ( .A(n541), .B(n540), .Z(n545) );
  NANDN U619 ( .A(n543), .B(n542), .Z(n544) );
  AND U620 ( .A(n545), .B(n544), .Z(n548) );
  NAND U621 ( .A(n[3]), .B(n546), .Z(n547) );
  XNOR U622 ( .A(n548), .B(n547), .Z(n549) );
  XNOR U623 ( .A(n550), .B(n549), .Z(n572) );
  NANDN U624 ( .A(n551), .B(n572), .Z(n552) );
  NAND U625 ( .A(n553), .B(n552), .Z(c[3]) );
  OR U626 ( .A(ereg[3]), .B(n43), .Z(n554) );
  AND U627 ( .A(first_one), .B(n554), .Z(n555) );
  ANDN U628 ( .B(init), .A(n555), .Z(n571) );
  NAND U629 ( .A(creg[0]), .B(n571), .Z(n558) );
  AND U630 ( .A(init), .B(n555), .Z(n573) );
  NAND U631 ( .A(n573), .B(n556), .Z(n557) );
  AND U632 ( .A(n558), .B(n557), .Z(n560) );
  NAND U633 ( .A(n560), .B(n559), .Z(n34) );
  NAND U634 ( .A(creg[1]), .B(n571), .Z(n563) );
  NAND U635 ( .A(n573), .B(n561), .Z(n562) );
  AND U636 ( .A(n563), .B(n562), .Z(n565) );
  NAND U637 ( .A(n565), .B(n564), .Z(n35) );
  NAND U638 ( .A(creg[2]), .B(n571), .Z(n568) );
  NAND U639 ( .A(n573), .B(n566), .Z(n567) );
  AND U640 ( .A(n568), .B(n567), .Z(n570) );
  NAND U641 ( .A(n570), .B(n569), .Z(n36) );
  NAND U642 ( .A(creg[3]), .B(n571), .Z(n575) );
  NAND U643 ( .A(n573), .B(n572), .Z(n574) );
  AND U644 ( .A(n575), .B(n574), .Z(n577) );
  NAND U645 ( .A(n577), .B(n576), .Z(n37) );
  AND U646 ( .A(init), .B(mul_pow), .Z(n587) );
  NAND U647 ( .A(ereg[3]), .B(n587), .Z(n578) );
  NANDN U648 ( .A(first_one), .B(n578), .Z(n38) );
  NAND U649 ( .A(ereg[2]), .B(n587), .Z(n580) );
  NAND U650 ( .A(ereg[3]), .B(n592), .Z(n579) );
  AND U651 ( .A(n580), .B(n579), .Z(n582) );
  NAND U652 ( .A(n582), .B(n581), .Z(n39) );
  NAND U653 ( .A(ereg[1]), .B(n587), .Z(n584) );
  NAND U654 ( .A(ereg[2]), .B(n592), .Z(n583) );
  AND U655 ( .A(n584), .B(n583), .Z(n586) );
  NANDN U656 ( .A(init), .B(e[2]), .Z(n585) );
  NAND U657 ( .A(n586), .B(n585), .Z(n40) );
  NAND U658 ( .A(ereg[0]), .B(n587), .Z(n589) );
  NAND U659 ( .A(ereg[1]), .B(n592), .Z(n588) );
  AND U660 ( .A(n589), .B(n588), .Z(n591) );
  NANDN U661 ( .A(init), .B(e[1]), .Z(n590) );
  NAND U662 ( .A(n591), .B(n590), .Z(n41) );
  NAND U663 ( .A(ereg[0]), .B(n592), .Z(n594) );
  NANDN U664 ( .A(init), .B(e[0]), .Z(n593) );
  NAND U665 ( .A(n594), .B(n593), .Z(n42) );
endmodule

