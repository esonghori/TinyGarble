
module sum_N128_CC1 ( clk, rst, a, b, c );
  input [127:0] a;
  input [127:0] b;
  output [127:0] c;
  input clk, rst;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508;

  NANDN U2 ( .A(n314), .B(b[126]), .Z(n2) );
  XNOR U3 ( .A(n314), .B(b[126]), .Z(n3) );
  NAND U4 ( .A(n3), .B(a[126]), .Z(n4) );
  NAND U5 ( .A(n2), .B(n4), .Z(n5) );
  XNOR U6 ( .A(a[127]), .B(n5), .Z(n6) );
  XNOR U7 ( .A(b[127]), .B(n6), .Z(c[127]) );
  XOR U8 ( .A(a[0]), .B(b[0]), .Z(c[0]) );
  XOR U9 ( .A(a[100]), .B(b[100]), .Z(n205) );
  NAND U10 ( .A(b[99]), .B(a[99]), .Z(n204) );
  XNOR U11 ( .A(b[99]), .B(a[99]), .Z(n506) );
  NAND U12 ( .A(b[98]), .B(a[98]), .Z(n202) );
  NAND U13 ( .A(b[97]), .B(a[97]), .Z(n200) );
  NAND U14 ( .A(b[96]), .B(a[96]), .Z(n198) );
  NAND U15 ( .A(b[95]), .B(a[95]), .Z(n196) );
  NAND U16 ( .A(b[94]), .B(a[94]), .Z(n194) );
  NAND U17 ( .A(b[93]), .B(a[93]), .Z(n192) );
  NAND U18 ( .A(b[92]), .B(a[92]), .Z(n190) );
  NAND U19 ( .A(b[91]), .B(a[91]), .Z(n188) );
  NAND U20 ( .A(b[90]), .B(a[90]), .Z(n186) );
  NAND U21 ( .A(b[89]), .B(a[89]), .Z(n184) );
  NAND U22 ( .A(b[88]), .B(a[88]), .Z(n182) );
  NAND U23 ( .A(b[87]), .B(a[87]), .Z(n180) );
  NAND U24 ( .A(b[86]), .B(a[86]), .Z(n178) );
  NAND U25 ( .A(b[85]), .B(a[85]), .Z(n176) );
  NAND U26 ( .A(b[84]), .B(a[84]), .Z(n174) );
  NAND U27 ( .A(b[83]), .B(a[83]), .Z(n172) );
  NAND U28 ( .A(b[82]), .B(a[82]), .Z(n170) );
  NAND U29 ( .A(b[81]), .B(a[81]), .Z(n168) );
  NAND U30 ( .A(b[80]), .B(a[80]), .Z(n166) );
  NAND U31 ( .A(b[79]), .B(a[79]), .Z(n164) );
  NAND U32 ( .A(b[78]), .B(a[78]), .Z(n162) );
  NAND U33 ( .A(b[77]), .B(a[77]), .Z(n160) );
  NAND U34 ( .A(b[76]), .B(a[76]), .Z(n158) );
  NAND U35 ( .A(b[75]), .B(a[75]), .Z(n156) );
  NAND U36 ( .A(b[74]), .B(a[74]), .Z(n154) );
  NAND U37 ( .A(b[73]), .B(a[73]), .Z(n152) );
  NAND U38 ( .A(b[72]), .B(a[72]), .Z(n150) );
  NAND U39 ( .A(b[71]), .B(a[71]), .Z(n148) );
  NAND U40 ( .A(b[70]), .B(a[70]), .Z(n146) );
  NAND U41 ( .A(b[69]), .B(a[69]), .Z(n144) );
  NAND U42 ( .A(b[68]), .B(a[68]), .Z(n142) );
  NAND U43 ( .A(b[67]), .B(a[67]), .Z(n140) );
  NAND U44 ( .A(b[66]), .B(a[66]), .Z(n138) );
  NAND U45 ( .A(b[65]), .B(a[65]), .Z(n136) );
  NAND U46 ( .A(b[64]), .B(a[64]), .Z(n134) );
  NAND U47 ( .A(b[63]), .B(a[63]), .Z(n132) );
  NAND U48 ( .A(b[62]), .B(a[62]), .Z(n130) );
  NAND U49 ( .A(b[61]), .B(a[61]), .Z(n128) );
  NAND U50 ( .A(b[60]), .B(a[60]), .Z(n126) );
  NAND U51 ( .A(b[59]), .B(a[59]), .Z(n124) );
  NAND U52 ( .A(b[58]), .B(a[58]), .Z(n122) );
  NAND U53 ( .A(b[57]), .B(a[57]), .Z(n120) );
  NAND U54 ( .A(b[56]), .B(a[56]), .Z(n118) );
  NAND U55 ( .A(b[55]), .B(a[55]), .Z(n116) );
  NAND U56 ( .A(b[54]), .B(a[54]), .Z(n114) );
  NAND U57 ( .A(b[53]), .B(a[53]), .Z(n112) );
  NAND U58 ( .A(b[52]), .B(a[52]), .Z(n110) );
  NAND U59 ( .A(b[51]), .B(a[51]), .Z(n108) );
  NAND U60 ( .A(b[50]), .B(a[50]), .Z(n106) );
  NAND U61 ( .A(b[49]), .B(a[49]), .Z(n104) );
  NAND U62 ( .A(b[48]), .B(a[48]), .Z(n102) );
  NAND U63 ( .A(b[47]), .B(a[47]), .Z(n100) );
  NAND U64 ( .A(b[46]), .B(a[46]), .Z(n98) );
  NAND U65 ( .A(b[45]), .B(a[45]), .Z(n96) );
  NAND U66 ( .A(b[44]), .B(a[44]), .Z(n94) );
  NAND U67 ( .A(b[43]), .B(a[43]), .Z(n92) );
  NAND U68 ( .A(b[42]), .B(a[42]), .Z(n90) );
  NAND U69 ( .A(b[41]), .B(a[41]), .Z(n88) );
  NAND U70 ( .A(b[40]), .B(a[40]), .Z(n86) );
  NAND U71 ( .A(b[39]), .B(a[39]), .Z(n84) );
  NAND U72 ( .A(b[38]), .B(a[38]), .Z(n82) );
  NAND U73 ( .A(b[37]), .B(a[37]), .Z(n80) );
  NAND U74 ( .A(b[36]), .B(a[36]), .Z(n78) );
  NAND U75 ( .A(b[35]), .B(a[35]), .Z(n76) );
  NAND U76 ( .A(b[34]), .B(a[34]), .Z(n74) );
  NAND U77 ( .A(b[33]), .B(a[33]), .Z(n72) );
  NAND U78 ( .A(b[32]), .B(a[32]), .Z(n70) );
  NAND U79 ( .A(b[31]), .B(a[31]), .Z(n68) );
  NAND U80 ( .A(b[30]), .B(a[30]), .Z(n66) );
  NAND U81 ( .A(b[29]), .B(a[29]), .Z(n64) );
  NAND U82 ( .A(b[28]), .B(a[28]), .Z(n62) );
  NAND U83 ( .A(b[27]), .B(a[27]), .Z(n60) );
  NAND U84 ( .A(b[26]), .B(a[26]), .Z(n58) );
  NAND U85 ( .A(b[25]), .B(a[25]), .Z(n56) );
  NAND U86 ( .A(b[24]), .B(a[24]), .Z(n54) );
  NAND U87 ( .A(b[23]), .B(a[23]), .Z(n52) );
  NAND U88 ( .A(b[22]), .B(a[22]), .Z(n50) );
  NAND U89 ( .A(b[21]), .B(a[21]), .Z(n48) );
  NAND U90 ( .A(b[20]), .B(a[20]), .Z(n46) );
  NAND U91 ( .A(b[19]), .B(a[19]), .Z(n44) );
  NAND U92 ( .A(b[18]), .B(a[18]), .Z(n42) );
  NAND U93 ( .A(b[17]), .B(a[17]), .Z(n40) );
  NAND U94 ( .A(b[16]), .B(a[16]), .Z(n38) );
  NAND U95 ( .A(b[15]), .B(a[15]), .Z(n36) );
  NAND U96 ( .A(b[14]), .B(a[14]), .Z(n34) );
  NAND U97 ( .A(b[13]), .B(a[13]), .Z(n32) );
  NAND U98 ( .A(b[12]), .B(a[12]), .Z(n30) );
  NAND U99 ( .A(b[11]), .B(a[11]), .Z(n28) );
  NAND U100 ( .A(b[10]), .B(a[10]), .Z(n26) );
  NAND U101 ( .A(b[9]), .B(a[9]), .Z(n24) );
  XNOR U102 ( .A(b[9]), .B(a[9]), .Z(n508) );
  NAND U103 ( .A(b[8]), .B(a[8]), .Z(n22) );
  NAND U104 ( .A(b[7]), .B(a[7]), .Z(n20) );
  NAND U105 ( .A(b[6]), .B(a[6]), .Z(n18) );
  NAND U106 ( .A(b[5]), .B(a[5]), .Z(n16) );
  NAND U107 ( .A(b[4]), .B(a[4]), .Z(n14) );
  NAND U108 ( .A(b[3]), .B(a[3]), .Z(n12) );
  NAND U109 ( .A(b[2]), .B(a[2]), .Z(n10) );
  NAND U110 ( .A(b[1]), .B(a[1]), .Z(n8) );
  NAND U111 ( .A(a[0]), .B(b[0]), .Z(n331) );
  XOR U112 ( .A(a[1]), .B(b[1]), .Z(n332) );
  NANDN U113 ( .A(n331), .B(n332), .Z(n7) );
  AND U114 ( .A(n8), .B(n7), .Z(n353) );
  XOR U115 ( .A(a[2]), .B(b[2]), .Z(n354) );
  NANDN U116 ( .A(n353), .B(n354), .Z(n9) );
  AND U117 ( .A(n10), .B(n9), .Z(n375) );
  XOR U118 ( .A(a[3]), .B(b[3]), .Z(n376) );
  NANDN U119 ( .A(n375), .B(n376), .Z(n11) );
  AND U120 ( .A(n12), .B(n11), .Z(n397) );
  XOR U121 ( .A(a[4]), .B(b[4]), .Z(n398) );
  NANDN U122 ( .A(n397), .B(n398), .Z(n13) );
  AND U123 ( .A(n14), .B(n13), .Z(n419) );
  XOR U124 ( .A(a[5]), .B(b[5]), .Z(n420) );
  NANDN U125 ( .A(n419), .B(n420), .Z(n15) );
  AND U126 ( .A(n16), .B(n15), .Z(n441) );
  XOR U127 ( .A(a[6]), .B(b[6]), .Z(n442) );
  NANDN U128 ( .A(n441), .B(n442), .Z(n17) );
  AND U129 ( .A(n18), .B(n17), .Z(n463) );
  XOR U130 ( .A(a[7]), .B(b[7]), .Z(n464) );
  NANDN U131 ( .A(n463), .B(n464), .Z(n19) );
  AND U132 ( .A(n20), .B(n19), .Z(n485) );
  XOR U133 ( .A(a[8]), .B(b[8]), .Z(n486) );
  NANDN U134 ( .A(n485), .B(n486), .Z(n21) );
  AND U135 ( .A(n22), .B(n21), .Z(n507) );
  OR U136 ( .A(n508), .B(n507), .Z(n23) );
  AND U137 ( .A(n24), .B(n23), .Z(n241) );
  XOR U138 ( .A(a[10]), .B(b[10]), .Z(n242) );
  NANDN U139 ( .A(n241), .B(n242), .Z(n25) );
  AND U140 ( .A(n26), .B(n25), .Z(n283) );
  XOR U141 ( .A(a[11]), .B(b[11]), .Z(n284) );
  NANDN U142 ( .A(n283), .B(n284), .Z(n27) );
  AND U143 ( .A(n28), .B(n27), .Z(n315) );
  XOR U144 ( .A(a[12]), .B(b[12]), .Z(n316) );
  NANDN U145 ( .A(n315), .B(n316), .Z(n29) );
  AND U146 ( .A(n30), .B(n29), .Z(n317) );
  XOR U147 ( .A(a[13]), .B(b[13]), .Z(n318) );
  NANDN U148 ( .A(n317), .B(n318), .Z(n31) );
  AND U149 ( .A(n32), .B(n31), .Z(n319) );
  XOR U150 ( .A(a[14]), .B(b[14]), .Z(n320) );
  NANDN U151 ( .A(n319), .B(n320), .Z(n33) );
  AND U152 ( .A(n34), .B(n33), .Z(n321) );
  XOR U153 ( .A(a[15]), .B(b[15]), .Z(n322) );
  NANDN U154 ( .A(n321), .B(n322), .Z(n35) );
  AND U155 ( .A(n36), .B(n35), .Z(n323) );
  XOR U156 ( .A(a[16]), .B(b[16]), .Z(n324) );
  NANDN U157 ( .A(n323), .B(n324), .Z(n37) );
  AND U158 ( .A(n38), .B(n37), .Z(n325) );
  XOR U159 ( .A(a[17]), .B(b[17]), .Z(n326) );
  NANDN U160 ( .A(n325), .B(n326), .Z(n39) );
  AND U161 ( .A(n40), .B(n39), .Z(n327) );
  XOR U162 ( .A(a[18]), .B(b[18]), .Z(n328) );
  NANDN U163 ( .A(n327), .B(n328), .Z(n41) );
  AND U164 ( .A(n42), .B(n41), .Z(n329) );
  XOR U165 ( .A(a[19]), .B(b[19]), .Z(n330) );
  NANDN U166 ( .A(n329), .B(n330), .Z(n43) );
  AND U167 ( .A(n44), .B(n43), .Z(n333) );
  XOR U168 ( .A(a[20]), .B(b[20]), .Z(n334) );
  NANDN U169 ( .A(n333), .B(n334), .Z(n45) );
  AND U170 ( .A(n46), .B(n45), .Z(n335) );
  XOR U171 ( .A(a[21]), .B(b[21]), .Z(n336) );
  NANDN U172 ( .A(n335), .B(n336), .Z(n47) );
  AND U173 ( .A(n48), .B(n47), .Z(n337) );
  XOR U174 ( .A(a[22]), .B(b[22]), .Z(n338) );
  NANDN U175 ( .A(n337), .B(n338), .Z(n49) );
  AND U176 ( .A(n50), .B(n49), .Z(n339) );
  XOR U177 ( .A(a[23]), .B(b[23]), .Z(n340) );
  NANDN U178 ( .A(n339), .B(n340), .Z(n51) );
  AND U179 ( .A(n52), .B(n51), .Z(n341) );
  XOR U180 ( .A(a[24]), .B(b[24]), .Z(n342) );
  NANDN U181 ( .A(n341), .B(n342), .Z(n53) );
  AND U182 ( .A(n54), .B(n53), .Z(n343) );
  XOR U183 ( .A(a[25]), .B(b[25]), .Z(n344) );
  NANDN U184 ( .A(n343), .B(n344), .Z(n55) );
  AND U185 ( .A(n56), .B(n55), .Z(n345) );
  XOR U186 ( .A(a[26]), .B(b[26]), .Z(n346) );
  NANDN U187 ( .A(n345), .B(n346), .Z(n57) );
  AND U188 ( .A(n58), .B(n57), .Z(n347) );
  XOR U189 ( .A(a[27]), .B(b[27]), .Z(n348) );
  NANDN U190 ( .A(n347), .B(n348), .Z(n59) );
  AND U191 ( .A(n60), .B(n59), .Z(n349) );
  XOR U192 ( .A(a[28]), .B(b[28]), .Z(n350) );
  NANDN U193 ( .A(n349), .B(n350), .Z(n61) );
  AND U194 ( .A(n62), .B(n61), .Z(n351) );
  XOR U195 ( .A(a[29]), .B(b[29]), .Z(n352) );
  NANDN U196 ( .A(n351), .B(n352), .Z(n63) );
  AND U197 ( .A(n64), .B(n63), .Z(n355) );
  XOR U198 ( .A(a[30]), .B(b[30]), .Z(n356) );
  NANDN U199 ( .A(n355), .B(n356), .Z(n65) );
  AND U200 ( .A(n66), .B(n65), .Z(n357) );
  XOR U201 ( .A(a[31]), .B(b[31]), .Z(n358) );
  NANDN U202 ( .A(n357), .B(n358), .Z(n67) );
  AND U203 ( .A(n68), .B(n67), .Z(n359) );
  XOR U204 ( .A(a[32]), .B(b[32]), .Z(n360) );
  NANDN U205 ( .A(n359), .B(n360), .Z(n69) );
  AND U206 ( .A(n70), .B(n69), .Z(n361) );
  XOR U207 ( .A(a[33]), .B(b[33]), .Z(n362) );
  NANDN U208 ( .A(n361), .B(n362), .Z(n71) );
  AND U209 ( .A(n72), .B(n71), .Z(n363) );
  XOR U210 ( .A(a[34]), .B(b[34]), .Z(n364) );
  NANDN U211 ( .A(n363), .B(n364), .Z(n73) );
  AND U212 ( .A(n74), .B(n73), .Z(n365) );
  XOR U213 ( .A(a[35]), .B(b[35]), .Z(n366) );
  NANDN U214 ( .A(n365), .B(n366), .Z(n75) );
  AND U215 ( .A(n76), .B(n75), .Z(n367) );
  XOR U216 ( .A(a[36]), .B(b[36]), .Z(n368) );
  NANDN U217 ( .A(n367), .B(n368), .Z(n77) );
  AND U218 ( .A(n78), .B(n77), .Z(n369) );
  XOR U219 ( .A(a[37]), .B(b[37]), .Z(n370) );
  NANDN U220 ( .A(n369), .B(n370), .Z(n79) );
  AND U221 ( .A(n80), .B(n79), .Z(n371) );
  XOR U222 ( .A(a[38]), .B(b[38]), .Z(n372) );
  NANDN U223 ( .A(n371), .B(n372), .Z(n81) );
  AND U224 ( .A(n82), .B(n81), .Z(n373) );
  XOR U225 ( .A(a[39]), .B(b[39]), .Z(n374) );
  NANDN U226 ( .A(n373), .B(n374), .Z(n83) );
  AND U227 ( .A(n84), .B(n83), .Z(n377) );
  XOR U228 ( .A(a[40]), .B(b[40]), .Z(n378) );
  NANDN U229 ( .A(n377), .B(n378), .Z(n85) );
  AND U230 ( .A(n86), .B(n85), .Z(n379) );
  XOR U231 ( .A(a[41]), .B(b[41]), .Z(n380) );
  NANDN U232 ( .A(n379), .B(n380), .Z(n87) );
  AND U233 ( .A(n88), .B(n87), .Z(n381) );
  XOR U234 ( .A(a[42]), .B(b[42]), .Z(n382) );
  NANDN U235 ( .A(n381), .B(n382), .Z(n89) );
  AND U236 ( .A(n90), .B(n89), .Z(n383) );
  XOR U237 ( .A(a[43]), .B(b[43]), .Z(n384) );
  NANDN U238 ( .A(n383), .B(n384), .Z(n91) );
  AND U239 ( .A(n92), .B(n91), .Z(n385) );
  XOR U240 ( .A(a[44]), .B(b[44]), .Z(n386) );
  NANDN U241 ( .A(n385), .B(n386), .Z(n93) );
  AND U242 ( .A(n94), .B(n93), .Z(n387) );
  XOR U243 ( .A(a[45]), .B(b[45]), .Z(n388) );
  NANDN U244 ( .A(n387), .B(n388), .Z(n95) );
  AND U245 ( .A(n96), .B(n95), .Z(n389) );
  XOR U246 ( .A(a[46]), .B(b[46]), .Z(n390) );
  NANDN U247 ( .A(n389), .B(n390), .Z(n97) );
  AND U248 ( .A(n98), .B(n97), .Z(n391) );
  XOR U249 ( .A(a[47]), .B(b[47]), .Z(n392) );
  NANDN U250 ( .A(n391), .B(n392), .Z(n99) );
  AND U251 ( .A(n100), .B(n99), .Z(n393) );
  XOR U252 ( .A(a[48]), .B(b[48]), .Z(n394) );
  NANDN U253 ( .A(n393), .B(n394), .Z(n101) );
  AND U254 ( .A(n102), .B(n101), .Z(n395) );
  XOR U255 ( .A(a[49]), .B(b[49]), .Z(n396) );
  NANDN U256 ( .A(n395), .B(n396), .Z(n103) );
  AND U257 ( .A(n104), .B(n103), .Z(n399) );
  XOR U258 ( .A(a[50]), .B(b[50]), .Z(n400) );
  NANDN U259 ( .A(n399), .B(n400), .Z(n105) );
  AND U260 ( .A(n106), .B(n105), .Z(n401) );
  XOR U261 ( .A(a[51]), .B(b[51]), .Z(n402) );
  NANDN U262 ( .A(n401), .B(n402), .Z(n107) );
  AND U263 ( .A(n108), .B(n107), .Z(n403) );
  XOR U264 ( .A(a[52]), .B(b[52]), .Z(n404) );
  NANDN U265 ( .A(n403), .B(n404), .Z(n109) );
  AND U266 ( .A(n110), .B(n109), .Z(n405) );
  XOR U267 ( .A(a[53]), .B(b[53]), .Z(n406) );
  NANDN U268 ( .A(n405), .B(n406), .Z(n111) );
  AND U269 ( .A(n112), .B(n111), .Z(n407) );
  XOR U270 ( .A(a[54]), .B(b[54]), .Z(n408) );
  NANDN U271 ( .A(n407), .B(n408), .Z(n113) );
  AND U272 ( .A(n114), .B(n113), .Z(n409) );
  XOR U273 ( .A(a[55]), .B(b[55]), .Z(n410) );
  NANDN U274 ( .A(n409), .B(n410), .Z(n115) );
  AND U275 ( .A(n116), .B(n115), .Z(n411) );
  XOR U276 ( .A(a[56]), .B(b[56]), .Z(n412) );
  NANDN U277 ( .A(n411), .B(n412), .Z(n117) );
  AND U278 ( .A(n118), .B(n117), .Z(n413) );
  XOR U279 ( .A(a[57]), .B(b[57]), .Z(n414) );
  NANDN U280 ( .A(n413), .B(n414), .Z(n119) );
  AND U281 ( .A(n120), .B(n119), .Z(n415) );
  XOR U282 ( .A(a[58]), .B(b[58]), .Z(n416) );
  NANDN U283 ( .A(n415), .B(n416), .Z(n121) );
  AND U284 ( .A(n122), .B(n121), .Z(n417) );
  XOR U285 ( .A(a[59]), .B(b[59]), .Z(n418) );
  NANDN U286 ( .A(n417), .B(n418), .Z(n123) );
  AND U287 ( .A(n124), .B(n123), .Z(n421) );
  XOR U288 ( .A(a[60]), .B(b[60]), .Z(n422) );
  NANDN U289 ( .A(n421), .B(n422), .Z(n125) );
  AND U290 ( .A(n126), .B(n125), .Z(n423) );
  XOR U291 ( .A(a[61]), .B(b[61]), .Z(n424) );
  NANDN U292 ( .A(n423), .B(n424), .Z(n127) );
  AND U293 ( .A(n128), .B(n127), .Z(n425) );
  XOR U294 ( .A(a[62]), .B(b[62]), .Z(n426) );
  NANDN U295 ( .A(n425), .B(n426), .Z(n129) );
  AND U296 ( .A(n130), .B(n129), .Z(n427) );
  XOR U297 ( .A(a[63]), .B(b[63]), .Z(n428) );
  NANDN U298 ( .A(n427), .B(n428), .Z(n131) );
  AND U299 ( .A(n132), .B(n131), .Z(n429) );
  XOR U300 ( .A(a[64]), .B(b[64]), .Z(n430) );
  NANDN U301 ( .A(n429), .B(n430), .Z(n133) );
  AND U302 ( .A(n134), .B(n133), .Z(n431) );
  XOR U303 ( .A(a[65]), .B(b[65]), .Z(n432) );
  NANDN U304 ( .A(n431), .B(n432), .Z(n135) );
  AND U305 ( .A(n136), .B(n135), .Z(n433) );
  XOR U306 ( .A(a[66]), .B(b[66]), .Z(n434) );
  NANDN U307 ( .A(n433), .B(n434), .Z(n137) );
  AND U308 ( .A(n138), .B(n137), .Z(n435) );
  XOR U309 ( .A(a[67]), .B(b[67]), .Z(n436) );
  NANDN U310 ( .A(n435), .B(n436), .Z(n139) );
  AND U311 ( .A(n140), .B(n139), .Z(n437) );
  XOR U312 ( .A(a[68]), .B(b[68]), .Z(n438) );
  NANDN U313 ( .A(n437), .B(n438), .Z(n141) );
  AND U314 ( .A(n142), .B(n141), .Z(n439) );
  XOR U315 ( .A(a[69]), .B(b[69]), .Z(n440) );
  NANDN U316 ( .A(n439), .B(n440), .Z(n143) );
  AND U317 ( .A(n144), .B(n143), .Z(n443) );
  XOR U318 ( .A(a[70]), .B(b[70]), .Z(n444) );
  NANDN U319 ( .A(n443), .B(n444), .Z(n145) );
  AND U320 ( .A(n146), .B(n145), .Z(n445) );
  XOR U321 ( .A(a[71]), .B(b[71]), .Z(n446) );
  NANDN U322 ( .A(n445), .B(n446), .Z(n147) );
  AND U323 ( .A(n148), .B(n147), .Z(n447) );
  XOR U324 ( .A(a[72]), .B(b[72]), .Z(n448) );
  NANDN U325 ( .A(n447), .B(n448), .Z(n149) );
  AND U326 ( .A(n150), .B(n149), .Z(n449) );
  XOR U327 ( .A(a[73]), .B(b[73]), .Z(n450) );
  NANDN U328 ( .A(n449), .B(n450), .Z(n151) );
  AND U329 ( .A(n152), .B(n151), .Z(n451) );
  XOR U330 ( .A(a[74]), .B(b[74]), .Z(n452) );
  NANDN U331 ( .A(n451), .B(n452), .Z(n153) );
  AND U332 ( .A(n154), .B(n153), .Z(n453) );
  XOR U333 ( .A(a[75]), .B(b[75]), .Z(n454) );
  NANDN U334 ( .A(n453), .B(n454), .Z(n155) );
  AND U335 ( .A(n156), .B(n155), .Z(n455) );
  XOR U336 ( .A(a[76]), .B(b[76]), .Z(n456) );
  NANDN U337 ( .A(n455), .B(n456), .Z(n157) );
  AND U338 ( .A(n158), .B(n157), .Z(n457) );
  XOR U339 ( .A(a[77]), .B(b[77]), .Z(n458) );
  NANDN U340 ( .A(n457), .B(n458), .Z(n159) );
  AND U341 ( .A(n160), .B(n159), .Z(n459) );
  XOR U342 ( .A(a[78]), .B(b[78]), .Z(n460) );
  NANDN U343 ( .A(n459), .B(n460), .Z(n161) );
  AND U344 ( .A(n162), .B(n161), .Z(n461) );
  XOR U345 ( .A(a[79]), .B(b[79]), .Z(n462) );
  NANDN U346 ( .A(n461), .B(n462), .Z(n163) );
  AND U347 ( .A(n164), .B(n163), .Z(n465) );
  XOR U348 ( .A(a[80]), .B(b[80]), .Z(n466) );
  NANDN U349 ( .A(n465), .B(n466), .Z(n165) );
  AND U350 ( .A(n166), .B(n165), .Z(n467) );
  XOR U351 ( .A(a[81]), .B(b[81]), .Z(n468) );
  NANDN U352 ( .A(n467), .B(n468), .Z(n167) );
  AND U353 ( .A(n168), .B(n167), .Z(n469) );
  XOR U354 ( .A(a[82]), .B(b[82]), .Z(n470) );
  NANDN U355 ( .A(n469), .B(n470), .Z(n169) );
  AND U356 ( .A(n170), .B(n169), .Z(n471) );
  XOR U357 ( .A(a[83]), .B(b[83]), .Z(n472) );
  NANDN U358 ( .A(n471), .B(n472), .Z(n171) );
  AND U359 ( .A(n172), .B(n171), .Z(n473) );
  XOR U360 ( .A(a[84]), .B(b[84]), .Z(n474) );
  NANDN U361 ( .A(n473), .B(n474), .Z(n173) );
  AND U362 ( .A(n174), .B(n173), .Z(n475) );
  XOR U363 ( .A(a[85]), .B(b[85]), .Z(n476) );
  NANDN U364 ( .A(n475), .B(n476), .Z(n175) );
  AND U365 ( .A(n176), .B(n175), .Z(n477) );
  XOR U366 ( .A(a[86]), .B(b[86]), .Z(n478) );
  NANDN U367 ( .A(n477), .B(n478), .Z(n177) );
  AND U368 ( .A(n178), .B(n177), .Z(n479) );
  XOR U369 ( .A(a[87]), .B(b[87]), .Z(n480) );
  NANDN U370 ( .A(n479), .B(n480), .Z(n179) );
  AND U371 ( .A(n180), .B(n179), .Z(n481) );
  XOR U372 ( .A(a[88]), .B(b[88]), .Z(n482) );
  NANDN U373 ( .A(n481), .B(n482), .Z(n181) );
  AND U374 ( .A(n182), .B(n181), .Z(n483) );
  XOR U375 ( .A(a[89]), .B(b[89]), .Z(n484) );
  NANDN U376 ( .A(n483), .B(n484), .Z(n183) );
  AND U377 ( .A(n184), .B(n183), .Z(n487) );
  XOR U378 ( .A(a[90]), .B(b[90]), .Z(n488) );
  NANDN U379 ( .A(n487), .B(n488), .Z(n185) );
  AND U380 ( .A(n186), .B(n185), .Z(n489) );
  XOR U381 ( .A(a[91]), .B(b[91]), .Z(n490) );
  NANDN U382 ( .A(n489), .B(n490), .Z(n187) );
  AND U383 ( .A(n188), .B(n187), .Z(n491) );
  XOR U384 ( .A(a[92]), .B(b[92]), .Z(n492) );
  NANDN U385 ( .A(n491), .B(n492), .Z(n189) );
  AND U386 ( .A(n190), .B(n189), .Z(n493) );
  XOR U387 ( .A(a[93]), .B(b[93]), .Z(n494) );
  NANDN U388 ( .A(n493), .B(n494), .Z(n191) );
  AND U389 ( .A(n192), .B(n191), .Z(n495) );
  XOR U390 ( .A(a[94]), .B(b[94]), .Z(n496) );
  NANDN U391 ( .A(n495), .B(n496), .Z(n193) );
  AND U392 ( .A(n194), .B(n193), .Z(n497) );
  XOR U393 ( .A(a[95]), .B(b[95]), .Z(n498) );
  NANDN U394 ( .A(n497), .B(n498), .Z(n195) );
  AND U395 ( .A(n196), .B(n195), .Z(n499) );
  XOR U396 ( .A(a[96]), .B(b[96]), .Z(n500) );
  NANDN U397 ( .A(n499), .B(n500), .Z(n197) );
  AND U398 ( .A(n198), .B(n197), .Z(n501) );
  XOR U399 ( .A(a[97]), .B(b[97]), .Z(n502) );
  NANDN U400 ( .A(n501), .B(n502), .Z(n199) );
  AND U401 ( .A(n200), .B(n199), .Z(n503) );
  XOR U402 ( .A(a[98]), .B(b[98]), .Z(n504) );
  NANDN U403 ( .A(n503), .B(n504), .Z(n201) );
  AND U404 ( .A(n202), .B(n201), .Z(n505) );
  OR U405 ( .A(n506), .B(n505), .Z(n203) );
  AND U406 ( .A(n204), .B(n203), .Z(n206) );
  XNOR U407 ( .A(n205), .B(n206), .Z(c[100]) );
  XOR U408 ( .A(a[101]), .B(b[101]), .Z(n209) );
  NAND U409 ( .A(b[100]), .B(a[100]), .Z(n208) );
  NANDN U410 ( .A(n206), .B(n205), .Z(n207) );
  AND U411 ( .A(n208), .B(n207), .Z(n210) );
  XNOR U412 ( .A(n209), .B(n210), .Z(c[101]) );
  XOR U413 ( .A(a[102]), .B(b[102]), .Z(n213) );
  NAND U414 ( .A(b[101]), .B(a[101]), .Z(n212) );
  NANDN U415 ( .A(n210), .B(n209), .Z(n211) );
  AND U416 ( .A(n212), .B(n211), .Z(n214) );
  XNOR U417 ( .A(n213), .B(n214), .Z(c[102]) );
  XOR U418 ( .A(a[103]), .B(b[103]), .Z(n217) );
  NAND U419 ( .A(b[102]), .B(a[102]), .Z(n216) );
  NANDN U420 ( .A(n214), .B(n213), .Z(n215) );
  AND U421 ( .A(n216), .B(n215), .Z(n218) );
  XNOR U422 ( .A(n217), .B(n218), .Z(c[103]) );
  XOR U423 ( .A(a[104]), .B(b[104]), .Z(n221) );
  NAND U424 ( .A(b[103]), .B(a[103]), .Z(n220) );
  NANDN U425 ( .A(n218), .B(n217), .Z(n219) );
  AND U426 ( .A(n220), .B(n219), .Z(n222) );
  XNOR U427 ( .A(n221), .B(n222), .Z(c[104]) );
  XOR U428 ( .A(a[105]), .B(b[105]), .Z(n225) );
  NAND U429 ( .A(b[104]), .B(a[104]), .Z(n224) );
  NANDN U430 ( .A(n222), .B(n221), .Z(n223) );
  AND U431 ( .A(n224), .B(n223), .Z(n226) );
  XNOR U432 ( .A(n225), .B(n226), .Z(c[105]) );
  XOR U433 ( .A(a[106]), .B(b[106]), .Z(n229) );
  NAND U434 ( .A(b[105]), .B(a[105]), .Z(n228) );
  NANDN U435 ( .A(n226), .B(n225), .Z(n227) );
  AND U436 ( .A(n228), .B(n227), .Z(n230) );
  XNOR U437 ( .A(n229), .B(n230), .Z(c[106]) );
  XOR U438 ( .A(a[107]), .B(b[107]), .Z(n233) );
  NAND U439 ( .A(b[106]), .B(a[106]), .Z(n232) );
  NANDN U440 ( .A(n230), .B(n229), .Z(n231) );
  AND U441 ( .A(n232), .B(n231), .Z(n234) );
  XNOR U442 ( .A(n233), .B(n234), .Z(c[107]) );
  XOR U443 ( .A(a[108]), .B(b[108]), .Z(n237) );
  NAND U444 ( .A(b[107]), .B(a[107]), .Z(n236) );
  NANDN U445 ( .A(n234), .B(n233), .Z(n235) );
  AND U446 ( .A(n236), .B(n235), .Z(n238) );
  XNOR U447 ( .A(n237), .B(n238), .Z(c[108]) );
  XOR U448 ( .A(a[109]), .B(b[109]), .Z(n243) );
  NAND U449 ( .A(b[108]), .B(a[108]), .Z(n240) );
  NANDN U450 ( .A(n238), .B(n237), .Z(n239) );
  AND U451 ( .A(n240), .B(n239), .Z(n244) );
  XNOR U452 ( .A(n243), .B(n244), .Z(c[109]) );
  XNOR U453 ( .A(n242), .B(n241), .Z(c[10]) );
  XOR U454 ( .A(a[110]), .B(b[110]), .Z(n247) );
  NAND U455 ( .A(b[109]), .B(a[109]), .Z(n246) );
  NANDN U456 ( .A(n244), .B(n243), .Z(n245) );
  AND U457 ( .A(n246), .B(n245), .Z(n248) );
  XNOR U458 ( .A(n247), .B(n248), .Z(c[110]) );
  XOR U459 ( .A(a[111]), .B(b[111]), .Z(n251) );
  NAND U460 ( .A(b[110]), .B(a[110]), .Z(n250) );
  NANDN U461 ( .A(n248), .B(n247), .Z(n249) );
  AND U462 ( .A(n250), .B(n249), .Z(n252) );
  XNOR U463 ( .A(n251), .B(n252), .Z(c[111]) );
  XOR U464 ( .A(a[112]), .B(b[112]), .Z(n255) );
  NAND U465 ( .A(b[111]), .B(a[111]), .Z(n254) );
  NANDN U466 ( .A(n252), .B(n251), .Z(n253) );
  AND U467 ( .A(n254), .B(n253), .Z(n256) );
  XNOR U468 ( .A(n255), .B(n256), .Z(c[112]) );
  XOR U469 ( .A(a[113]), .B(b[113]), .Z(n259) );
  NAND U470 ( .A(b[112]), .B(a[112]), .Z(n258) );
  NANDN U471 ( .A(n256), .B(n255), .Z(n257) );
  AND U472 ( .A(n258), .B(n257), .Z(n260) );
  XNOR U473 ( .A(n259), .B(n260), .Z(c[113]) );
  XOR U474 ( .A(a[114]), .B(b[114]), .Z(n263) );
  NAND U475 ( .A(b[113]), .B(a[113]), .Z(n262) );
  NANDN U476 ( .A(n260), .B(n259), .Z(n261) );
  AND U477 ( .A(n262), .B(n261), .Z(n264) );
  XNOR U478 ( .A(n263), .B(n264), .Z(c[114]) );
  XOR U479 ( .A(a[115]), .B(b[115]), .Z(n267) );
  NAND U480 ( .A(b[114]), .B(a[114]), .Z(n266) );
  NANDN U481 ( .A(n264), .B(n263), .Z(n265) );
  AND U482 ( .A(n266), .B(n265), .Z(n268) );
  XNOR U483 ( .A(n267), .B(n268), .Z(c[115]) );
  XOR U484 ( .A(a[116]), .B(b[116]), .Z(n271) );
  NAND U485 ( .A(b[115]), .B(a[115]), .Z(n270) );
  NANDN U486 ( .A(n268), .B(n267), .Z(n269) );
  AND U487 ( .A(n270), .B(n269), .Z(n272) );
  XNOR U488 ( .A(n271), .B(n272), .Z(c[116]) );
  XOR U489 ( .A(a[117]), .B(b[117]), .Z(n275) );
  NAND U490 ( .A(b[116]), .B(a[116]), .Z(n274) );
  NANDN U491 ( .A(n272), .B(n271), .Z(n273) );
  AND U492 ( .A(n274), .B(n273), .Z(n276) );
  XNOR U493 ( .A(n275), .B(n276), .Z(c[117]) );
  XOR U494 ( .A(a[118]), .B(b[118]), .Z(n279) );
  NAND U495 ( .A(b[117]), .B(a[117]), .Z(n278) );
  NANDN U496 ( .A(n276), .B(n275), .Z(n277) );
  AND U497 ( .A(n278), .B(n277), .Z(n280) );
  XNOR U498 ( .A(n279), .B(n280), .Z(c[118]) );
  XOR U499 ( .A(a[119]), .B(b[119]), .Z(n285) );
  NAND U500 ( .A(b[118]), .B(a[118]), .Z(n282) );
  NANDN U501 ( .A(n280), .B(n279), .Z(n281) );
  AND U502 ( .A(n282), .B(n281), .Z(n286) );
  XNOR U503 ( .A(n285), .B(n286), .Z(c[119]) );
  XNOR U504 ( .A(n284), .B(n283), .Z(c[11]) );
  XOR U505 ( .A(a[120]), .B(b[120]), .Z(n289) );
  NAND U506 ( .A(b[119]), .B(a[119]), .Z(n288) );
  NANDN U507 ( .A(n286), .B(n285), .Z(n287) );
  AND U508 ( .A(n288), .B(n287), .Z(n290) );
  XNOR U509 ( .A(n289), .B(n290), .Z(c[120]) );
  XOR U510 ( .A(a[121]), .B(b[121]), .Z(n293) );
  NAND U511 ( .A(b[120]), .B(a[120]), .Z(n292) );
  NANDN U512 ( .A(n290), .B(n289), .Z(n291) );
  AND U513 ( .A(n292), .B(n291), .Z(n294) );
  XNOR U514 ( .A(n293), .B(n294), .Z(c[121]) );
  XOR U515 ( .A(a[122]), .B(b[122]), .Z(n297) );
  NAND U516 ( .A(b[121]), .B(a[121]), .Z(n296) );
  NANDN U517 ( .A(n294), .B(n293), .Z(n295) );
  AND U518 ( .A(n296), .B(n295), .Z(n298) );
  XNOR U519 ( .A(n297), .B(n298), .Z(c[122]) );
  XOR U520 ( .A(a[123]), .B(b[123]), .Z(n301) );
  NAND U521 ( .A(b[122]), .B(a[122]), .Z(n300) );
  NANDN U522 ( .A(n298), .B(n297), .Z(n299) );
  AND U523 ( .A(n300), .B(n299), .Z(n302) );
  XNOR U524 ( .A(n301), .B(n302), .Z(c[123]) );
  XOR U525 ( .A(a[124]), .B(b[124]), .Z(n305) );
  NAND U526 ( .A(b[123]), .B(a[123]), .Z(n304) );
  NANDN U527 ( .A(n302), .B(n301), .Z(n303) );
  AND U528 ( .A(n304), .B(n303), .Z(n306) );
  XNOR U529 ( .A(n305), .B(n306), .Z(c[124]) );
  XOR U530 ( .A(a[125]), .B(b[125]), .Z(n309) );
  NAND U531 ( .A(b[124]), .B(a[124]), .Z(n308) );
  NANDN U532 ( .A(n306), .B(n305), .Z(n307) );
  AND U533 ( .A(n308), .B(n307), .Z(n310) );
  XNOR U534 ( .A(n309), .B(n310), .Z(c[125]) );
  NAND U535 ( .A(b[125]), .B(a[125]), .Z(n312) );
  NANDN U536 ( .A(n310), .B(n309), .Z(n311) );
  AND U537 ( .A(n312), .B(n311), .Z(n314) );
  XOR U538 ( .A(a[126]), .B(n314), .Z(n313) );
  XNOR U539 ( .A(b[126]), .B(n313), .Z(c[126]) );
  XNOR U540 ( .A(n316), .B(n315), .Z(c[12]) );
  XNOR U541 ( .A(n318), .B(n317), .Z(c[13]) );
  XNOR U542 ( .A(n320), .B(n319), .Z(c[14]) );
  XNOR U543 ( .A(n322), .B(n321), .Z(c[15]) );
  XNOR U544 ( .A(n324), .B(n323), .Z(c[16]) );
  XNOR U545 ( .A(n326), .B(n325), .Z(c[17]) );
  XNOR U546 ( .A(n328), .B(n327), .Z(c[18]) );
  XNOR U547 ( .A(n330), .B(n329), .Z(c[19]) );
  XNOR U548 ( .A(n332), .B(n331), .Z(c[1]) );
  XNOR U549 ( .A(n334), .B(n333), .Z(c[20]) );
  XNOR U550 ( .A(n336), .B(n335), .Z(c[21]) );
  XNOR U551 ( .A(n338), .B(n337), .Z(c[22]) );
  XNOR U552 ( .A(n340), .B(n339), .Z(c[23]) );
  XNOR U553 ( .A(n342), .B(n341), .Z(c[24]) );
  XNOR U554 ( .A(n344), .B(n343), .Z(c[25]) );
  XNOR U555 ( .A(n346), .B(n345), .Z(c[26]) );
  XNOR U556 ( .A(n348), .B(n347), .Z(c[27]) );
  XNOR U557 ( .A(n350), .B(n349), .Z(c[28]) );
  XNOR U558 ( .A(n352), .B(n351), .Z(c[29]) );
  XNOR U559 ( .A(n354), .B(n353), .Z(c[2]) );
  XNOR U560 ( .A(n356), .B(n355), .Z(c[30]) );
  XNOR U561 ( .A(n358), .B(n357), .Z(c[31]) );
  XNOR U562 ( .A(n360), .B(n359), .Z(c[32]) );
  XNOR U563 ( .A(n362), .B(n361), .Z(c[33]) );
  XNOR U564 ( .A(n364), .B(n363), .Z(c[34]) );
  XNOR U565 ( .A(n366), .B(n365), .Z(c[35]) );
  XNOR U566 ( .A(n368), .B(n367), .Z(c[36]) );
  XNOR U567 ( .A(n370), .B(n369), .Z(c[37]) );
  XNOR U568 ( .A(n372), .B(n371), .Z(c[38]) );
  XNOR U569 ( .A(n374), .B(n373), .Z(c[39]) );
  XNOR U570 ( .A(n376), .B(n375), .Z(c[3]) );
  XNOR U571 ( .A(n378), .B(n377), .Z(c[40]) );
  XNOR U572 ( .A(n380), .B(n379), .Z(c[41]) );
  XNOR U573 ( .A(n382), .B(n381), .Z(c[42]) );
  XNOR U574 ( .A(n384), .B(n383), .Z(c[43]) );
  XNOR U575 ( .A(n386), .B(n385), .Z(c[44]) );
  XNOR U576 ( .A(n388), .B(n387), .Z(c[45]) );
  XNOR U577 ( .A(n390), .B(n389), .Z(c[46]) );
  XNOR U578 ( .A(n392), .B(n391), .Z(c[47]) );
  XNOR U579 ( .A(n394), .B(n393), .Z(c[48]) );
  XNOR U580 ( .A(n396), .B(n395), .Z(c[49]) );
  XNOR U581 ( .A(n398), .B(n397), .Z(c[4]) );
  XNOR U582 ( .A(n400), .B(n399), .Z(c[50]) );
  XNOR U583 ( .A(n402), .B(n401), .Z(c[51]) );
  XNOR U584 ( .A(n404), .B(n403), .Z(c[52]) );
  XNOR U585 ( .A(n406), .B(n405), .Z(c[53]) );
  XNOR U586 ( .A(n408), .B(n407), .Z(c[54]) );
  XNOR U587 ( .A(n410), .B(n409), .Z(c[55]) );
  XNOR U588 ( .A(n412), .B(n411), .Z(c[56]) );
  XNOR U589 ( .A(n414), .B(n413), .Z(c[57]) );
  XNOR U590 ( .A(n416), .B(n415), .Z(c[58]) );
  XNOR U591 ( .A(n418), .B(n417), .Z(c[59]) );
  XNOR U592 ( .A(n420), .B(n419), .Z(c[5]) );
  XNOR U593 ( .A(n422), .B(n421), .Z(c[60]) );
  XNOR U594 ( .A(n424), .B(n423), .Z(c[61]) );
  XNOR U595 ( .A(n426), .B(n425), .Z(c[62]) );
  XNOR U596 ( .A(n428), .B(n427), .Z(c[63]) );
  XNOR U597 ( .A(n430), .B(n429), .Z(c[64]) );
  XNOR U598 ( .A(n432), .B(n431), .Z(c[65]) );
  XNOR U599 ( .A(n434), .B(n433), .Z(c[66]) );
  XNOR U600 ( .A(n436), .B(n435), .Z(c[67]) );
  XNOR U601 ( .A(n438), .B(n437), .Z(c[68]) );
  XNOR U602 ( .A(n440), .B(n439), .Z(c[69]) );
  XNOR U603 ( .A(n442), .B(n441), .Z(c[6]) );
  XNOR U604 ( .A(n444), .B(n443), .Z(c[70]) );
  XNOR U605 ( .A(n446), .B(n445), .Z(c[71]) );
  XNOR U606 ( .A(n448), .B(n447), .Z(c[72]) );
  XNOR U607 ( .A(n450), .B(n449), .Z(c[73]) );
  XNOR U608 ( .A(n452), .B(n451), .Z(c[74]) );
  XNOR U609 ( .A(n454), .B(n453), .Z(c[75]) );
  XNOR U610 ( .A(n456), .B(n455), .Z(c[76]) );
  XNOR U611 ( .A(n458), .B(n457), .Z(c[77]) );
  XNOR U612 ( .A(n460), .B(n459), .Z(c[78]) );
  XNOR U613 ( .A(n462), .B(n461), .Z(c[79]) );
  XNOR U614 ( .A(n464), .B(n463), .Z(c[7]) );
  XNOR U615 ( .A(n466), .B(n465), .Z(c[80]) );
  XNOR U616 ( .A(n468), .B(n467), .Z(c[81]) );
  XNOR U617 ( .A(n470), .B(n469), .Z(c[82]) );
  XNOR U618 ( .A(n472), .B(n471), .Z(c[83]) );
  XNOR U619 ( .A(n474), .B(n473), .Z(c[84]) );
  XNOR U620 ( .A(n476), .B(n475), .Z(c[85]) );
  XNOR U621 ( .A(n478), .B(n477), .Z(c[86]) );
  XNOR U622 ( .A(n480), .B(n479), .Z(c[87]) );
  XNOR U623 ( .A(n482), .B(n481), .Z(c[88]) );
  XNOR U624 ( .A(n484), .B(n483), .Z(c[89]) );
  XNOR U625 ( .A(n486), .B(n485), .Z(c[8]) );
  XNOR U626 ( .A(n488), .B(n487), .Z(c[90]) );
  XNOR U627 ( .A(n490), .B(n489), .Z(c[91]) );
  XNOR U628 ( .A(n492), .B(n491), .Z(c[92]) );
  XNOR U629 ( .A(n494), .B(n493), .Z(c[93]) );
  XNOR U630 ( .A(n496), .B(n495), .Z(c[94]) );
  XNOR U631 ( .A(n498), .B(n497), .Z(c[95]) );
  XNOR U632 ( .A(n500), .B(n499), .Z(c[96]) );
  XNOR U633 ( .A(n502), .B(n501), .Z(c[97]) );
  XNOR U634 ( .A(n504), .B(n503), .Z(c[98]) );
  XOR U635 ( .A(n506), .B(n505), .Z(c[99]) );
  XOR U636 ( .A(n508), .B(n507), .Z(c[9]) );
endmodule

