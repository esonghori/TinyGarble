`include "../defined.vh"

module Control 
( 
	opcode,
	rs_index,
	rt_index,
	rd_index,
	imm_out,
	alu_func,
	shift_func,
	mult_func,
	branch_func,
	a_source_out,
	b_source_out,
	c_source_out,
	pc_source_out,
	mem_source_out
);

	input 	[31:0]	opcode;
	output	[4:0]	rs_index;
	output	[4:0]	rt_index;
	output	[4:0]	rd_index;
	output	[15:0]	imm_out;
	output	[3:0]	alu_func;
	output	[1:0]	shift_func;
	output	[3:0]	mult_func;
	output	[2:0]	branch_func;
	output	[1:0]	a_source_out;
	output	[1:0]	b_source_out;
	output	[2:0]	c_source_out;
	output	[1:0]	pc_source_out;
	output	[3:0]	mem_source_out;


	reg	[4:0]	rs_index;
	reg	[4:0]	rt_index;
	reg	[4:0]	rd_index;
	reg	[3:0]	alu_func;
	reg	[1:0]	shift_func;
	reg	[3:0]	mult_func;
	reg	[2:0]	branch_func;
	reg	[1:0]	a_source_out;
	reg	[1:0]	b_source_out;
	reg	[2:0]	c_source_out;
	reg	[1:0]	pc_source_out;
	reg	[3:0]	mem_source_out;

	
	wire	[5:0]	op,func;
	wire	[4:0]	r1,r2,r3,sham;
	
	
	assign op=opcode[31:26];
	assign func=opcode[5:0];
	assign r1=opcode[25:21];
	assign r2=opcode[20:16];
	assign r3=opcode[15:11];
	assign sham=opcode[10:6];

	assign imm_out=opcode[15:0];
	
	always@(*)
	begin
		rs_index<=r1;
		rt_index<=r2;
		rd_index<=5'b0;
		alu_func<=`ALU_NOTHING;
		shift_func<=`SHIFT_NOTHING;
		mult_func<=`MULT_NOTHING;
		branch_func<=`BRANCH_NO;
		a_source_out<=`A_FROM_REG_SOURCE;
		b_source_out<=`B_FROM_REG_TARGET;
		c_source_out<=`C_FROM_ALU;//`C_FROM_SHIFT,`C_FROM_MULT
		pc_source_out<=`FROM_INC4;
		mem_source_out<=`MEM_FETCH;
		//////
		case(opcode[31:29])
		3'b000:
			case(opcode[28:26])
			3'b000://SPECIAL
				begin
					rs_index<=r1;
					rt_index<=r2;
					case(func[5:3])
					3'b000:
						case(func[2:0])
						3'b000://SLL
							begin
								if(r2==0 && r3==0)
									$display("NOP");
								else
									$display("SLL");
								shift_func<=`SHIFT_LEFT_UNSIGNED;
								a_source_out<=`A_FROM_IMM10_6;//shift amount
								b_source_out<=`B_FROM_REG_TARGET;
								rt_index<=r2;
								rd_index<=r3;
							end
						3'b001://-
							;
						3'b010://SRL
							begin
								$display("SLR");
								shift_func<=`SHIFT_RIGHT_UNSIGNED;
								a_source_out<=`A_FROM_IMM10_6;//shift amount
								b_source_out<=`B_FROM_REG_TARGET;
								rt_index<=r2;
								rd_index<=r3;
							end
						3'b011://SRA
							begin
								$display("SRA");
								shift_func<=`SHIFT_RIGHT_SIGNED;
								a_source_out<=`A_FROM_IMM10_6;//shift amount
								b_source_out<=`B_FROM_REG_TARGET;
								rt_index<=r2;
								rd_index<=r3;
							end
						3'b100://SLLV
							begin
								$display("SLLV");
								shift_func<=`SHIFT_LEFT_UNSIGNED;
								a_source_out<=`A_FROM_REG_SOURCE;
								b_source_out<=`B_FROM_REG_TARGET;
								rs_index<=r1;
								rt_index<=r2;
								rd_index<=r3;
							end
						3'b101://-
							;
						3'b110://SRLV
							begin
								$display("SRLV");
								shift_func<=`SHIFT_RIGHT_UNSIGNED;
								a_source_out<=`A_FROM_REG_SOURCE;
								b_source_out<=`B_FROM_REG_TARGET;
								rs_index<=r1;
								rt_index<=r2;
								rd_index<=r3;
							end
						3'b111://SRAV
							begin
								$display("SRAV");
								shift_func<=`SHIFT_RIGHT_SIGNED;
								a_source_out<=`A_FROM_REG_SOURCE;
								b_source_out<=`B_FROM_REG_TARGET;
								rs_index<=r1;
								rt_index<=r2;
								rd_index<=r3;
							end
						endcase
					3'b001:
						case(func[2:0])
						3'b000://JR
							begin
								$display("JR");
								rs_index<=r1;
								rt_index<=0;
								rd_index<=0;
								branch_func<=`BRANCH_YES;
								pc_source_out<=`FROM_LBRANCH;
								alu_func<=`ALU_OR;
							end
						3'b001://JALR
							begin
								$display("JALR");
								rs_index<=r1;
								rt_index<=0;
								rd_index<=r3;
								branch_func<=`BRANCH_YES;
								pc_source_out<=`FROM_LBRANCH;
								c_source_out<=`C_FROM_PC_PLUS4;
								alu_func<=`ALU_OR;
							end
						3'b010://--
							;
						3'b011://--
							;
						3'b100://SYSCALL
						begin
							$display("SYSCALL");
							rs_index<=63;//ISR
							rt_index<=0;
							rd_index<=46;//EPC
							branch_func<=`BRANCH_YES;
							pc_source_out<=`FROM_LBRANCH;
							c_source_out<=`C_FROM_PC_PLUS4;
							alu_func<=`ALU_OR;
						end
						3'b101://BREAK
						begin
							$display("BREAK");
							rs_index<=63;//ISR
							rt_index<=0;
							rd_index<=46;//EPC
							branch_func<=`BRANCH_YES;
							pc_source_out<=`FROM_LBRANCH;
							c_source_out<=`C_FROM_PC_PLUS4;
							alu_func<=`ALU_OR;
						end
						3'b110://--
							;
						3'b111://SYNC
							$display("SYNC");
						endcase
					3'b010:
						case(func[2:0])
						3'b000://MFHI
						begin
							$display("MFHI");
							mult_func<=`MULT_READ_HI;
							rd_index<=r3;
						end
						3'b001://MTHI
						begin
							$display("MTHI");
							mult_func<=`MULT_WRITE_HI;
						end
						3'b010://MFLO
						begin
							$display("MFLO");
							mult_func<=`MULT_READ_LO;
							rd_index<=r3;
						end
						3'b011://MTLO
						begin
							$display("MTLO");
							mult_func<=`MULT_WRITE_LO;
						end
						3'b100://-
							;
						3'b101://-
							;
						3'b110://-
							;
						3'b111://-
							;
						endcase
					3'b011:
						case(func[2:0])
						3'b000://MULT
						begin
							$display("MULT");
							mult_func<=`MULT_SIGNED_MULT;
						end
						3'b001://MULTU
						begin
							$display("MULTU");
							mult_func<=`MULT_MULT;
						end
						3'b010://DIV
						begin
							$display("DIV");
							mult_func<=`MULT_SIGNED_DIVIDE;
						end
						3'b011://DIVU
						begin
							$display("DIVU");
							mult_func<=`MULT_DIVIDE;
						end
						3'b100://--
							;
						3'b101://-
							;
						3'b110://-
							;
						3'b111://-
							;
						endcase
					3'b100:
					begin
						rd_index<=r3;
						case(func[2:0])
						3'b000://ADD
						begin
							$display("ADD");
							alu_func<=`ALU_ADD;
						end
						3'b001://ADDU
						begin
							$display("ADDU");
							alu_func<=`ALU_ADD;
						end
						3'b010://SUB
						begin
							$display("SUB");
							alu_func<=`ALU_SUBTRACT;
						end
						3'b011://SUBU
						begin
							$display("SUBU");
							alu_func<=`ALU_SUBTRACT;
						end
						3'b100://AND
						begin
							$display("AND");
							alu_func<=`ALU_AND;
						end
						3'b101://OR
						begin
							$display("OR");
							alu_func<=`ALU_OR;
						end
						3'b110://XOR
						begin
							$display("XOR");
							alu_func<=`ALU_XOR;
						end
						3'b111://NOR
						begin
							$display("NOR");
							alu_func<=`ALU_NOR;
						end
						endcase
					end
					3'b101:
						case(func[2:0])
						3'b000://-
							;
						3'b001://-
							;
						3'b010://SLT
						begin
							$display("SLT");
							rd_index<=r3;
							alu_func<=`ALU_LESS_THAN_SIGNED;
						end
						3'b011://SLTU
						begin
							$display("SLTU");
							rd_index<=r3;
							alu_func<=`ALU_LESS_THAN;
						end
						3'b100://-
							;
						3'b101://-
							;
						3'b110://-
							;
						3'b111://-
							;
						endcase
					3'b110:
						case(func[2:0])
						3'b000://TGE
							;
						3'b001://TGEU
							;
						3'b010://TLT
							;
						3'b011://TLTU
							;
						3'b100://TEQ
							;
						3'b101://-
							;
						3'b110://TNE
							;
						3'b111://-
							;
						endcase
					3'b111:
						case(func[2:0])
						3'b000://-
							;
						3'b001://-
							;
						3'b010://-
							;
						3'b011://-
							;
						3'b100://-
							;
						3'b101://-
							;
						3'b110://-
							;
						3'b111://-
							;
						endcase
					endcase
				end
			3'b001://REGIMM
				begin
					case(opcode[20:19])
					2'b00:
						case(opcode[18:16])
						3'b000://BLTZ
						begin	
							$display("BLTZ");
							rs_index<=r1;
							rt_index<=0;
							alu_func<=`ALU_OR;
							branch_func<=`BRANCH_LTZ;
							pc_source_out<=`FROM_BRANCH;
						end
						3'b001://BGEZ
						begin	
							$display("BGEZ");
							rs_index<=r1;
							rt_index<=0;
							alu_func<=`ALU_OR;
							branch_func<=`BRANCH_GEZ;
							pc_source_out<=`FROM_BRANCH;
						end
						3'b010://BLTZL
							;
						3'b011://BGEZL
							;
						3'b100://-
							;
						3'b101://-
							;
						3'b110://-
							;
						3'b111://-
							;
						endcase
					2'b01:
						case(opcode[18:16])
						3'b000://TGEI
							;
						3'b001://TGEI
							;
						3'b010://TLTI
							;
						3'b011://TLTIU
							;
						3'b100://TEQI
							;
						3'b101://-
							;
						3'b110://TNEI
							;
						3'b111://-
							;
						endcase
					2'b10:
						case(opcode[18:16])
						3'b000://BLTZAL
						begin	
							$display("BLTZAL");
							rs_index<=r1;
							rt_index<=0;
							rd_index<=31;
							alu_func<=`ALU_OR;
							branch_func<=`BRANCH_LTZ;
							pc_source_out<=`FROM_BRANCH;
							c_source_out<=`C_FROM_PC_PLUS4;
						end
						3'b001://BGEZAL
						begin	
							$display("BGEZAL");
							rs_index<=r1;
							rt_index<=0;
							rd_index<=31;
							alu_func<=`ALU_OR;
							branch_func<=`BRANCH_GEZ;
							pc_source_out<=`FROM_BRANCH;
							c_source_out<=`C_FROM_PC_PLUS4;
						end
						3'b010://BLTZALL
							;
						3'b011://BGEZALL
							;
						3'b100://
							;
						3'b101://
							;
						3'b110://
							;
						3'b111://
							;
						endcase
					2'b11:
						case(opcode[18:16])
						3'b000://-
							;
						3'b001://-
							;
						3'b010://-
							;
						3'b011://-
							;
						3'b100://-
							;
						3'b101://-
							;
						3'b110://-
							;
						3'b111://-
							;
						endcase
					endcase
				end
			3'b010://J
			begin
				$display("J");
				branch_func<=`BRANCH_YES;
				pc_source_out<=`FROM_OPCODE25_0;
			end
			3'b011://JAL
			begin
				$display("JAL");
				rd_index<=31;
				c_source_out<=`C_FROM_PC_PLUS4;
				branch_func<=`BRANCH_YES;
				pc_source_out<=`FROM_OPCODE25_0;
			end
			3'b100://BEQ
			begin
				$display("BEQ");
				rs_index<=r1;
				rt_index<=r2;
				alu_func<=`ALU_XOR;
				branch_func<=`BRANCH_EQ;
				pc_source_out<=`FROM_BRANCH;
			end
			3'b101://BNE
			begin
				$display("BNE");
				rs_index<=r1;
				rt_index<=r2;
				alu_func<=`ALU_XOR;
				branch_func<=`BRANCH_NE;
				pc_source_out<=`FROM_BRANCH;
			end
			3'b110://BLEZ
			begin
				$display("BLEZ");
				rs_index<=r1;
				rt_index<=0;
				alu_func<=`ALU_OR;
				branch_func<=`BRANCH_LEZ;
				pc_source_out<=`FROM_BRANCH;
			end
			3'b111://BGTZ
			begin
				$display("BGTZ");
				rs_index<=r1;
				rt_index<=0;
				alu_func<=`ALU_OR;
				branch_func<=`BRANCH_GTZ;
				pc_source_out<=`FROM_BRANCH;
			end
			endcase
		3'b001:
			case(opcode[28:26])
			3'b000://ADDI
			begin
				$display("ADDI");
				rs_index<=r1;
				rd_index<=r2;
				b_source_out<=`B_FROM_SIGNED_IMM;
				alu_func<=`ALU_ADD;
			end
			3'b001://ADDIU
			begin
				$display("ADDIU");
				rs_index<=r1;
				rd_index<=r2;
				b_source_out<=`B_FROM_SIGNED_IMM;
				alu_func<=`ALU_ADD;
			end
			3'b010://SLTI
			begin
				$display("SLTI");
				rs_index<=r1;
				rd_index<=r2;
				b_source_out<=`B_FROM_SIGNED_IMM;
				alu_func<=`ALU_LESS_THAN_SIGNED;
			end
			3'b011://SLTIU
			begin
				$display("SLTIU");
				rs_index<=r1;
				rd_index<=r2;
				b_source_out<=`B_FROM_IMM;
				alu_func<=`ALU_LESS_THAN;
			end
			3'b100://ANDI
			begin
				$display("ANDI");
				rs_index<=r1;
				rd_index<=r2;
				b_source_out<=`B_FROM_IMM;
				alu_func<=`ALU_AND;
			end
			3'b101://ORI
			begin
				$display("ORI");
				rs_index<=r1;
				rd_index<=r2;
				b_source_out<=`B_FROM_IMM;
				alu_func<=`ALU_OR;
			end
			3'b110://XORI
			begin
				$display("XORI");
				rs_index<=r1;
				rd_index<=r2;
				b_source_out<=`B_FROM_IMM;
				alu_func<=`ALU_XOR;
			end
			3'b111://LUI
			begin
				$display("LUI");
				rd_index<=r2;
				c_source_out<=`C_FROM_IMM_SHIFT16;
			end
			endcase
		3'b010:
			case(opcode[28:26])
			3'b000://COP0
			begin
				case(opcode[25:21])
				5'b00000://MFC0
				begin
					$display("MFC0");
					rs_index<={1'b1,r3};
					rt_index<=6'b0;
					rd_index<=r2;
					alu_func<=`ALU_OR;
				end
				5'b00100://MTC0
				begin
					$display("MTC0");
					rs_index<=r2;
					rt_index<=6'b0;
					rd_index<={1'b1,r3};
					alu_func<=`ALU_OR;
				end
				default:
					;
				endcase
			end
			3'b001://COP1
				;
			3'b010://COP2
				;
			3'b011://COP3
				;
			3'b100://BEQL
				;
			3'b101://BNEL
				;
			3'b110://BLEZL
				;
			3'b111://BGTZL
				;
			endcase
		3'b011:
			case(opcode[28:26])
			3'b000://-
				;
			3'b001://-
				;
			3'b010://-
				;
			3'b011://-
				;
			3'b100://-
				;
			3'b101://-
				;
			3'b110://-
				;
			3'b111://-
				;
			endcase
		3'b100:
			case(opcode[28:26])
			3'b000://LB
			begin
				$display("LB");
				rs_index<=r1;
				rd_index<=r2;
				b_source_out<=`B_FROM_SIGNED_IMM;
				alu_func<=`ALU_ADD;
				c_source_out<=`C_FROM_MEMORY;
				mem_source_out<=`MEM_READ8S;
			end
			3'b001://LH
			begin
				$display("LH");
				rs_index<=r1;
				rd_index<=r2;
				b_source_out<=`B_FROM_SIGNED_IMM;
				alu_func<=`ALU_ADD;
				c_source_out<=`C_FROM_MEMORY;
				mem_source_out<=`MEM_READ16S;
			end
			3'b010://LWL
			begin
				$display("LWL");
				rs_index<=r1;
				rd_index<=r2;
				b_source_out<=`B_FROM_SIGNED_IMM;
				alu_func<=`ALU_ADD;
				c_source_out<=`C_FROM_MEMORY;
				mem_source_out<=`MEM_READ32; //TODO: fix it
			end
			3'b011://LW
			begin
				$display("LW");
				rs_index<=r1;
				rd_index<=r2;
				b_source_out<=`B_FROM_SIGNED_IMM;
				alu_func<=`ALU_ADD;
				c_source_out<=`C_FROM_MEMORY;
				mem_source_out<=`MEM_READ32;
			end
			3'b100://LBU
			begin
				$display("LBU");
				rs_index<=r1;
				rd_index<=r2;
				b_source_out<=`B_FROM_SIGNED_IMM;
				alu_func<=`ALU_ADD;
				c_source_out<=`C_FROM_MEMORY;
				mem_source_out<=`MEM_READ8;
			end
			3'b101://LHU
			begin
				$display("LHU");
				rs_index<=r1;
				rd_index<=r2;
				b_source_out<=`B_FROM_SIGNED_IMM;
				alu_func<=`ALU_ADD;
				c_source_out<=`C_FROM_MEMORY;
				mem_source_out<=`MEM_READ16;
			end
			3'b110://LWR
			begin
				$display("LWR");
				rs_index<=r1;
				rd_index<=r2;
				b_source_out<=`B_FROM_SIGNED_IMM;
				alu_func<=`ALU_ADD;
				c_source_out<=`C_FROM_MEMORY;
				mem_source_out<=`MEM_READ32; //TODO: fix it
			end
			3'b111://-
				;
			endcase
		3'b101:
			case(opcode[28:26])
			3'b000://SB
			begin
				$display("SB");
				rs_index<=r1;
				rt_index<=r2;
				b_source_out<=`B_FROM_SIGNED_IMM;
				alu_func<=`ALU_ADD;
				mem_source_out<=`MEM_WRITE8;
			end
			3'b001://SH
			begin
				$display("SH");
				rs_index<=r1;
				rt_index<=r2;
				b_source_out<=`B_FROM_SIGNED_IMM;
				alu_func<=`ALU_ADD;
				mem_source_out<=`MEM_WRITE16;
			end
			3'b010://SWL
			begin
				$display("SWL");
				rs_index<=r1;
				rt_index<=r2;
				b_source_out<=`B_FROM_SIGNED_IMM;
				alu_func<=`ALU_ADD;
				mem_source_out<=`MEM_WRITE32;
			end
			3'b011://SW
			begin
				$display("SW");
				rs_index<=r1;
				rt_index<=r2;
				b_source_out<=`B_FROM_SIGNED_IMM;
				alu_func<=`ALU_ADD;
				mem_source_out<=`MEM_WRITE32;
			end
			3'b100://-
				;
			3'b101://-
				;
			3'b110://SWR
				;
			3'b111://ro
				;
			endcase
		3'b110:
			case(opcode[28:26])
			3'b000://LL
				;
			3'b001://LWC1
				;
			3'b010://LWC1
				;
			3'b011://LWC3
				;
			3'b100://-
				;
			3'b101://LDC1
				;
			3'b110://LDC2
				;
			3'b111://LDC3
				;
			endcase
		3'b111:
			case(opcode[28:26])
			3'b000://SC
				;
			3'b001://SWC1
				;
			3'b010://SWC2
				;
			3'b011://SWC3
				;
			3'b100://-
				;
			3'b101://SDC1
				;
			3'b110://SDC2
				;
			3'b111://SDC3
				;
			endcase
		endcase
	end
endmodule
