
module mult_N128_CC8 ( clk, rst, a, b, c );
  input [127:0] a;
  input [15:0] b;
  output [127:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294;
  wire   [127:16] swire;
  wire   [255:128] sreg;

  DFF \sreg_reg[128]  ( .D(swire[16]), .CLK(clk), .RST(rst), .Q(sreg[128]) );
  DFF \sreg_reg[129]  ( .D(swire[17]), .CLK(clk), .RST(rst), .Q(sreg[129]) );
  DFF \sreg_reg[130]  ( .D(swire[18]), .CLK(clk), .RST(rst), .Q(sreg[130]) );
  DFF \sreg_reg[131]  ( .D(swire[19]), .CLK(clk), .RST(rst), .Q(sreg[131]) );
  DFF \sreg_reg[132]  ( .D(swire[20]), .CLK(clk), .RST(rst), .Q(sreg[132]) );
  DFF \sreg_reg[133]  ( .D(swire[21]), .CLK(clk), .RST(rst), .Q(sreg[133]) );
  DFF \sreg_reg[134]  ( .D(swire[22]), .CLK(clk), .RST(rst), .Q(sreg[134]) );
  DFF \sreg_reg[135]  ( .D(swire[23]), .CLK(clk), .RST(rst), .Q(sreg[135]) );
  DFF \sreg_reg[136]  ( .D(swire[24]), .CLK(clk), .RST(rst), .Q(sreg[136]) );
  DFF \sreg_reg[137]  ( .D(swire[25]), .CLK(clk), .RST(rst), .Q(sreg[137]) );
  DFF \sreg_reg[138]  ( .D(swire[26]), .CLK(clk), .RST(rst), .Q(sreg[138]) );
  DFF \sreg_reg[139]  ( .D(swire[27]), .CLK(clk), .RST(rst), .Q(sreg[139]) );
  DFF \sreg_reg[140]  ( .D(swire[28]), .CLK(clk), .RST(rst), .Q(sreg[140]) );
  DFF \sreg_reg[141]  ( .D(swire[29]), .CLK(clk), .RST(rst), .Q(sreg[141]) );
  DFF \sreg_reg[142]  ( .D(swire[30]), .CLK(clk), .RST(rst), .Q(sreg[142]) );
  DFF \sreg_reg[143]  ( .D(swire[31]), .CLK(clk), .RST(rst), .Q(sreg[143]) );
  DFF \sreg_reg[144]  ( .D(swire[32]), .CLK(clk), .RST(rst), .Q(sreg[144]) );
  DFF \sreg_reg[145]  ( .D(swire[33]), .CLK(clk), .RST(rst), .Q(sreg[145]) );
  DFF \sreg_reg[146]  ( .D(swire[34]), .CLK(clk), .RST(rst), .Q(sreg[146]) );
  DFF \sreg_reg[147]  ( .D(swire[35]), .CLK(clk), .RST(rst), .Q(sreg[147]) );
  DFF \sreg_reg[148]  ( .D(swire[36]), .CLK(clk), .RST(rst), .Q(sreg[148]) );
  DFF \sreg_reg[149]  ( .D(swire[37]), .CLK(clk), .RST(rst), .Q(sreg[149]) );
  DFF \sreg_reg[150]  ( .D(swire[38]), .CLK(clk), .RST(rst), .Q(sreg[150]) );
  DFF \sreg_reg[151]  ( .D(swire[39]), .CLK(clk), .RST(rst), .Q(sreg[151]) );
  DFF \sreg_reg[152]  ( .D(swire[40]), .CLK(clk), .RST(rst), .Q(sreg[152]) );
  DFF \sreg_reg[153]  ( .D(swire[41]), .CLK(clk), .RST(rst), .Q(sreg[153]) );
  DFF \sreg_reg[154]  ( .D(swire[42]), .CLK(clk), .RST(rst), .Q(sreg[154]) );
  DFF \sreg_reg[155]  ( .D(swire[43]), .CLK(clk), .RST(rst), .Q(sreg[155]) );
  DFF \sreg_reg[156]  ( .D(swire[44]), .CLK(clk), .RST(rst), .Q(sreg[156]) );
  DFF \sreg_reg[157]  ( .D(swire[45]), .CLK(clk), .RST(rst), .Q(sreg[157]) );
  DFF \sreg_reg[158]  ( .D(swire[46]), .CLK(clk), .RST(rst), .Q(sreg[158]) );
  DFF \sreg_reg[159]  ( .D(swire[47]), .CLK(clk), .RST(rst), .Q(sreg[159]) );
  DFF \sreg_reg[160]  ( .D(swire[48]), .CLK(clk), .RST(rst), .Q(sreg[160]) );
  DFF \sreg_reg[161]  ( .D(swire[49]), .CLK(clk), .RST(rst), .Q(sreg[161]) );
  DFF \sreg_reg[162]  ( .D(swire[50]), .CLK(clk), .RST(rst), .Q(sreg[162]) );
  DFF \sreg_reg[163]  ( .D(swire[51]), .CLK(clk), .RST(rst), .Q(sreg[163]) );
  DFF \sreg_reg[164]  ( .D(swire[52]), .CLK(clk), .RST(rst), .Q(sreg[164]) );
  DFF \sreg_reg[165]  ( .D(swire[53]), .CLK(clk), .RST(rst), .Q(sreg[165]) );
  DFF \sreg_reg[166]  ( .D(swire[54]), .CLK(clk), .RST(rst), .Q(sreg[166]) );
  DFF \sreg_reg[167]  ( .D(swire[55]), .CLK(clk), .RST(rst), .Q(sreg[167]) );
  DFF \sreg_reg[168]  ( .D(swire[56]), .CLK(clk), .RST(rst), .Q(sreg[168]) );
  DFF \sreg_reg[169]  ( .D(swire[57]), .CLK(clk), .RST(rst), .Q(sreg[169]) );
  DFF \sreg_reg[170]  ( .D(swire[58]), .CLK(clk), .RST(rst), .Q(sreg[170]) );
  DFF \sreg_reg[171]  ( .D(swire[59]), .CLK(clk), .RST(rst), .Q(sreg[171]) );
  DFF \sreg_reg[172]  ( .D(swire[60]), .CLK(clk), .RST(rst), .Q(sreg[172]) );
  DFF \sreg_reg[173]  ( .D(swire[61]), .CLK(clk), .RST(rst), .Q(sreg[173]) );
  DFF \sreg_reg[174]  ( .D(swire[62]), .CLK(clk), .RST(rst), .Q(sreg[174]) );
  DFF \sreg_reg[175]  ( .D(swire[63]), .CLK(clk), .RST(rst), .Q(sreg[175]) );
  DFF \sreg_reg[176]  ( .D(swire[64]), .CLK(clk), .RST(rst), .Q(sreg[176]) );
  DFF \sreg_reg[177]  ( .D(swire[65]), .CLK(clk), .RST(rst), .Q(sreg[177]) );
  DFF \sreg_reg[178]  ( .D(swire[66]), .CLK(clk), .RST(rst), .Q(sreg[178]) );
  DFF \sreg_reg[179]  ( .D(swire[67]), .CLK(clk), .RST(rst), .Q(sreg[179]) );
  DFF \sreg_reg[180]  ( .D(swire[68]), .CLK(clk), .RST(rst), .Q(sreg[180]) );
  DFF \sreg_reg[181]  ( .D(swire[69]), .CLK(clk), .RST(rst), .Q(sreg[181]) );
  DFF \sreg_reg[182]  ( .D(swire[70]), .CLK(clk), .RST(rst), .Q(sreg[182]) );
  DFF \sreg_reg[183]  ( .D(swire[71]), .CLK(clk), .RST(rst), .Q(sreg[183]) );
  DFF \sreg_reg[184]  ( .D(swire[72]), .CLK(clk), .RST(rst), .Q(sreg[184]) );
  DFF \sreg_reg[185]  ( .D(swire[73]), .CLK(clk), .RST(rst), .Q(sreg[185]) );
  DFF \sreg_reg[186]  ( .D(swire[74]), .CLK(clk), .RST(rst), .Q(sreg[186]) );
  DFF \sreg_reg[187]  ( .D(swire[75]), .CLK(clk), .RST(rst), .Q(sreg[187]) );
  DFF \sreg_reg[188]  ( .D(swire[76]), .CLK(clk), .RST(rst), .Q(sreg[188]) );
  DFF \sreg_reg[189]  ( .D(swire[77]), .CLK(clk), .RST(rst), .Q(sreg[189]) );
  DFF \sreg_reg[190]  ( .D(swire[78]), .CLK(clk), .RST(rst), .Q(sreg[190]) );
  DFF \sreg_reg[191]  ( .D(swire[79]), .CLK(clk), .RST(rst), .Q(sreg[191]) );
  DFF \sreg_reg[192]  ( .D(swire[80]), .CLK(clk), .RST(rst), .Q(sreg[192]) );
  DFF \sreg_reg[193]  ( .D(swire[81]), .CLK(clk), .RST(rst), .Q(sreg[193]) );
  DFF \sreg_reg[194]  ( .D(swire[82]), .CLK(clk), .RST(rst), .Q(sreg[194]) );
  DFF \sreg_reg[195]  ( .D(swire[83]), .CLK(clk), .RST(rst), .Q(sreg[195]) );
  DFF \sreg_reg[196]  ( .D(swire[84]), .CLK(clk), .RST(rst), .Q(sreg[196]) );
  DFF \sreg_reg[197]  ( .D(swire[85]), .CLK(clk), .RST(rst), .Q(sreg[197]) );
  DFF \sreg_reg[198]  ( .D(swire[86]), .CLK(clk), .RST(rst), .Q(sreg[198]) );
  DFF \sreg_reg[199]  ( .D(swire[87]), .CLK(clk), .RST(rst), .Q(sreg[199]) );
  DFF \sreg_reg[200]  ( .D(swire[88]), .CLK(clk), .RST(rst), .Q(sreg[200]) );
  DFF \sreg_reg[201]  ( .D(swire[89]), .CLK(clk), .RST(rst), .Q(sreg[201]) );
  DFF \sreg_reg[202]  ( .D(swire[90]), .CLK(clk), .RST(rst), .Q(sreg[202]) );
  DFF \sreg_reg[203]  ( .D(swire[91]), .CLK(clk), .RST(rst), .Q(sreg[203]) );
  DFF \sreg_reg[204]  ( .D(swire[92]), .CLK(clk), .RST(rst), .Q(sreg[204]) );
  DFF \sreg_reg[205]  ( .D(swire[93]), .CLK(clk), .RST(rst), .Q(sreg[205]) );
  DFF \sreg_reg[206]  ( .D(swire[94]), .CLK(clk), .RST(rst), .Q(sreg[206]) );
  DFF \sreg_reg[207]  ( .D(swire[95]), .CLK(clk), .RST(rst), .Q(sreg[207]) );
  DFF \sreg_reg[208]  ( .D(swire[96]), .CLK(clk), .RST(rst), .Q(sreg[208]) );
  DFF \sreg_reg[209]  ( .D(swire[97]), .CLK(clk), .RST(rst), .Q(sreg[209]) );
  DFF \sreg_reg[210]  ( .D(swire[98]), .CLK(clk), .RST(rst), .Q(sreg[210]) );
  DFF \sreg_reg[211]  ( .D(swire[99]), .CLK(clk), .RST(rst), .Q(sreg[211]) );
  DFF \sreg_reg[212]  ( .D(swire[100]), .CLK(clk), .RST(rst), .Q(sreg[212]) );
  DFF \sreg_reg[213]  ( .D(swire[101]), .CLK(clk), .RST(rst), .Q(sreg[213]) );
  DFF \sreg_reg[214]  ( .D(swire[102]), .CLK(clk), .RST(rst), .Q(sreg[214]) );
  DFF \sreg_reg[215]  ( .D(swire[103]), .CLK(clk), .RST(rst), .Q(sreg[215]) );
  DFF \sreg_reg[216]  ( .D(swire[104]), .CLK(clk), .RST(rst), .Q(sreg[216]) );
  DFF \sreg_reg[217]  ( .D(swire[105]), .CLK(clk), .RST(rst), .Q(sreg[217]) );
  DFF \sreg_reg[218]  ( .D(swire[106]), .CLK(clk), .RST(rst), .Q(sreg[218]) );
  DFF \sreg_reg[219]  ( .D(swire[107]), .CLK(clk), .RST(rst), .Q(sreg[219]) );
  DFF \sreg_reg[220]  ( .D(swire[108]), .CLK(clk), .RST(rst), .Q(sreg[220]) );
  DFF \sreg_reg[221]  ( .D(swire[109]), .CLK(clk), .RST(rst), .Q(sreg[221]) );
  DFF \sreg_reg[222]  ( .D(swire[110]), .CLK(clk), .RST(rst), .Q(sreg[222]) );
  DFF \sreg_reg[223]  ( .D(swire[111]), .CLK(clk), .RST(rst), .Q(sreg[223]) );
  DFF \sreg_reg[224]  ( .D(swire[112]), .CLK(clk), .RST(rst), .Q(sreg[224]) );
  DFF \sreg_reg[225]  ( .D(swire[113]), .CLK(clk), .RST(rst), .Q(sreg[225]) );
  DFF \sreg_reg[226]  ( .D(swire[114]), .CLK(clk), .RST(rst), .Q(sreg[226]) );
  DFF \sreg_reg[227]  ( .D(swire[115]), .CLK(clk), .RST(rst), .Q(sreg[227]) );
  DFF \sreg_reg[228]  ( .D(swire[116]), .CLK(clk), .RST(rst), .Q(sreg[228]) );
  DFF \sreg_reg[229]  ( .D(swire[117]), .CLK(clk), .RST(rst), .Q(sreg[229]) );
  DFF \sreg_reg[230]  ( .D(swire[118]), .CLK(clk), .RST(rst), .Q(sreg[230]) );
  DFF \sreg_reg[231]  ( .D(swire[119]), .CLK(clk), .RST(rst), .Q(sreg[231]) );
  DFF \sreg_reg[232]  ( .D(swire[120]), .CLK(clk), .RST(rst), .Q(sreg[232]) );
  DFF \sreg_reg[233]  ( .D(swire[121]), .CLK(clk), .RST(rst), .Q(sreg[233]) );
  DFF \sreg_reg[234]  ( .D(swire[122]), .CLK(clk), .RST(rst), .Q(sreg[234]) );
  DFF \sreg_reg[235]  ( .D(swire[123]), .CLK(clk), .RST(rst), .Q(sreg[235]) );
  DFF \sreg_reg[236]  ( .D(swire[124]), .CLK(clk), .RST(rst), .Q(sreg[236]) );
  DFF \sreg_reg[237]  ( .D(swire[125]), .CLK(clk), .RST(rst), .Q(sreg[237]) );
  DFF \sreg_reg[238]  ( .D(swire[126]), .CLK(clk), .RST(rst), .Q(sreg[238]) );
  DFF \sreg_reg[239]  ( .D(swire[127]), .CLK(clk), .RST(rst), .Q(sreg[239]) );
  DFF \sreg_reg[127]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[126]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[125]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[124]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[123]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[122]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[121]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[120]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[119]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[118]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[117]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[116]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[115]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[114]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[113]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[112]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[111]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[110]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[109]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[108]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[107]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[106]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[105]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[104]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[103]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[102]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[101]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[100]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[99]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[98]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[97]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[96]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[95]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[94]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[93]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[92]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[91]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[90]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[89]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[88]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[87]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[86]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[85]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[84]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[83]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[82]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[81]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[80]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[79]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[78]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[77]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[76]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[75]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[74]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[73]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[72]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[71]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[70]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[69]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[68]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[67]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[66]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[65]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[64]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[63]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[62]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[61]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[60]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[59]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[58]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[57]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[56]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[55]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[54]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[53]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[52]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[51]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[50]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[49]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[48]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[47]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[46]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[45]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[44]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[43]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[42]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[41]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[40]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[39]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[38]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[37]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[36]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[35]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[34]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[33]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[32]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[31]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[30]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[29]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[28]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[27]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[26]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[25]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[24]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[23]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[22]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[21]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[20]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[19]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[18]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[17]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[16]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[0]) );
  XOR U19 ( .A(n9235), .B(n9293), .Z(n9240) );
  XOR U20 ( .A(n2981), .B(n3006), .Z(n2985) );
  XOR U21 ( .A(n3141), .B(n3166), .Z(n3145) );
  XOR U22 ( .A(n3110), .B(n3172), .Z(n3115) );
  XOR U23 ( .A(n4164), .B(n4225), .Z(n4168) );
  XOR U24 ( .A(n4323), .B(n4385), .Z(n4328) );
  XOR U25 ( .A(n5383), .B(n5444), .Z(n5387) );
  XOR U26 ( .A(n5542), .B(n5604), .Z(n5547) );
  XOR U27 ( .A(n6608), .B(n6669), .Z(n6612) );
  XOR U28 ( .A(n6767), .B(n6829), .Z(n6772) );
  XOR U29 ( .A(n7839), .B(n7900), .Z(n7843) );
  XOR U30 ( .A(n7998), .B(n8060), .Z(n8003) );
  XNOR U31 ( .A(n9242), .B(n9159), .Z(n9161) );
  XNOR U32 ( .A(n9317), .B(n9239), .Z(n9241) );
  XNOR U33 ( .A(n9386), .B(n9314), .Z(n9316) );
  XOR U34 ( .A(n2966), .B(n3009), .Z(n2970) );
  XOR U35 ( .A(n3061), .B(n3086), .Z(n3065) );
  XOR U36 ( .A(n3220), .B(n3245), .Z(n3224) );
  XOR U37 ( .A(n3457), .B(n3482), .Z(n3461) );
  XOR U38 ( .A(n3615), .B(n3640), .Z(n3619) );
  XOR U39 ( .A(n4194), .B(n4219), .Z(n4198) );
  XOR U40 ( .A(n4354), .B(n4379), .Z(n4358) );
  XOR U41 ( .A(n4512), .B(n4537), .Z(n4516) );
  XOR U42 ( .A(n4670), .B(n4695), .Z(n4674) );
  XOR U43 ( .A(n4828), .B(n4853), .Z(n4832) );
  XOR U44 ( .A(n5413), .B(n5418), .Z(n5336) );
  XOR U45 ( .A(n5573), .B(n5578), .Z(n5503) );
  XOR U46 ( .A(n5731), .B(n5736), .Z(n5662) );
  XOR U47 ( .A(n5889), .B(n5894), .Z(n5820) );
  XOR U48 ( .A(n6047), .B(n6052), .Z(n5978) );
  XOR U49 ( .A(n6578), .B(n6556), .Z(n6530) );
  XOR U50 ( .A(n6744), .B(n6722), .Z(n6648) );
  XOR U51 ( .A(n6903), .B(n6881), .Z(n6808) );
  XOR U52 ( .A(n7061), .B(n7039), .Z(n6966) );
  XOR U53 ( .A(n7219), .B(n7197), .Z(n7124) );
  XOR U54 ( .A(n7772), .B(n7750), .Z(n7676) );
  XOR U55 ( .A(n7895), .B(n7873), .Z(n7794) );
  XOR U56 ( .A(n8055), .B(n8033), .Z(n7959) );
  XOR U57 ( .A(n8213), .B(n8191), .Z(n8118) );
  XOR U58 ( .A(n8371), .B(n8349), .Z(n8276) );
  XOR U59 ( .A(n9004), .B(n8982), .Z(n8908) );
  XOR U60 ( .A(n9132), .B(n9110), .Z(n9032) );
  XOR U61 ( .A(n9288), .B(n9270), .Z(n9196) );
  XOR U62 ( .A(n1739), .B(n1814), .Z(n1744) );
  XOR U63 ( .A(n3264), .B(n3332), .Z(n3273) );
  XOR U64 ( .A(n4477), .B(n4545), .Z(n4486) );
  XOR U65 ( .A(n5696), .B(n5764), .Z(n5705) );
  XOR U66 ( .A(n6921), .B(n6989), .Z(n6930) );
  XOR U67 ( .A(n2261), .B(n2329), .Z(n2265) );
  XOR U68 ( .A(n9156), .B(n9217), .Z(n9160) );
  XNOR U69 ( .A(n3122), .B(n3039), .Z(n3041) );
  XOR U70 ( .A(n3512), .B(n3567), .Z(n3516) );
  XOR U71 ( .A(n3907), .B(n3962), .Z(n3911) );
  XOR U72 ( .A(n4725), .B(n4780), .Z(n4729) );
  XOR U73 ( .A(n5120), .B(n5175), .Z(n5124) );
  XOR U74 ( .A(n5944), .B(n5999), .Z(n5948) );
  XOR U75 ( .A(n6339), .B(n6395), .Z(n6343) );
  XOR U76 ( .A(n7169), .B(n7224), .Z(n7173) );
  XOR U77 ( .A(n7565), .B(n7621), .Z(n7569) );
  XOR U78 ( .A(n8797), .B(n8853), .Z(n8801) );
  XOR U79 ( .A(n388), .B(n448), .Z(n392) );
  XOR U80 ( .A(n2013), .B(n2069), .Z(n2017) );
  XNOR U81 ( .A(n3285), .B(n3203), .Z(n3205) );
  XNOR U82 ( .A(n3364), .B(n3282), .Z(n3284) );
  XNOR U83 ( .A(n3443), .B(n3361), .Z(n3363) );
  XNOR U84 ( .A(n4260), .B(n4177), .Z(n4179) );
  XNOR U85 ( .A(n4340), .B(n4257), .Z(n4259) );
  XNOR U86 ( .A(n4419), .B(n4337), .Z(n4339) );
  XNOR U87 ( .A(n4498), .B(n4416), .Z(n4418) );
  XNOR U88 ( .A(n4577), .B(n4495), .Z(n4497) );
  XNOR U89 ( .A(n4656), .B(n4574), .Z(n4576) );
  XNOR U90 ( .A(n5479), .B(n5396), .Z(n5398) );
  XNOR U91 ( .A(n5559), .B(n5476), .Z(n5478) );
  XNOR U92 ( .A(n5638), .B(n5556), .Z(n5558) );
  XNOR U93 ( .A(n5717), .B(n5635), .Z(n5637) );
  XNOR U94 ( .A(n5796), .B(n5714), .Z(n5716) );
  XNOR U95 ( .A(n5875), .B(n5793), .Z(n5795) );
  XNOR U96 ( .A(n6704), .B(n6621), .Z(n6623) );
  XNOR U97 ( .A(n6784), .B(n6701), .Z(n6703) );
  XNOR U98 ( .A(n6863), .B(n6781), .Z(n6783) );
  XNOR U99 ( .A(n6942), .B(n6860), .Z(n6862) );
  XNOR U100 ( .A(n7021), .B(n6939), .Z(n6941) );
  XNOR U101 ( .A(n7100), .B(n7018), .Z(n7020) );
  XNOR U102 ( .A(n7935), .B(n7852), .Z(n7854) );
  XNOR U103 ( .A(n8015), .B(n7932), .Z(n7934) );
  XNOR U104 ( .A(n8094), .B(n8012), .Z(n8014) );
  XNOR U105 ( .A(n8173), .B(n8091), .Z(n8093) );
  XNOR U106 ( .A(n8252), .B(n8170), .Z(n8172) );
  XOR U107 ( .A(n8241), .B(n8295), .Z(n8250) );
  XNOR U108 ( .A(n9172), .B(n9089), .Z(n9091) );
  XNOR U109 ( .A(n9252), .B(n9169), .Z(n9171) );
  XNOR U110 ( .A(n9327), .B(n9249), .Z(n9251) );
  XOR U111 ( .A(n9390), .B(n9423), .Z(n9394) );
  XNOR U112 ( .A(n3132), .B(n3049), .Z(n3051) );
  XNOR U113 ( .A(n8414), .B(n8453), .Z(n8409) );
  XOR U114 ( .A(n2971), .B(n3008), .Z(n2975) );
  XNOR U115 ( .A(n9403), .B(n9402), .Z(n9358) );
  XOR U116 ( .A(n328), .B(n364), .Z(n332) );
  XOR U117 ( .A(n488), .B(n525), .Z(n492) );
  XOR U118 ( .A(n2883), .B(n2918), .Z(n2887) );
  XNOR U119 ( .A(n3384), .B(n3302), .Z(n3304) );
  XOR U120 ( .A(n3378), .B(n3403), .Z(n3382) );
  XOR U121 ( .A(n3536), .B(n3561), .Z(n3540) );
  XOR U122 ( .A(n3689), .B(n3719), .Z(n3698) );
  XOR U123 ( .A(n4274), .B(n4299), .Z(n4278) );
  XOR U124 ( .A(n4433), .B(n4458), .Z(n4437) );
  XOR U125 ( .A(n4591), .B(n4616), .Z(n4595) );
  XOR U126 ( .A(n4749), .B(n4774), .Z(n4753) );
  XOR U127 ( .A(n4902), .B(n4932), .Z(n4911) );
  XOR U128 ( .A(n5493), .B(n5498), .Z(n5423) );
  XOR U129 ( .A(n5652), .B(n5657), .Z(n5583) );
  XOR U130 ( .A(n5810), .B(n5815), .Z(n5741) );
  XOR U131 ( .A(n5968), .B(n5973), .Z(n5899) );
  XOR U132 ( .A(n6121), .B(n6131), .Z(n6057) );
  XOR U133 ( .A(n6664), .B(n6642), .Z(n6562) );
  XOR U134 ( .A(n6824), .B(n6802), .Z(n6728) );
  XOR U135 ( .A(n6982), .B(n6960), .Z(n6887) );
  XOR U136 ( .A(n7140), .B(n7118), .Z(n7045) );
  XOR U137 ( .A(n7298), .B(n7276), .Z(n7203) );
  XOR U138 ( .A(n7810), .B(n7788), .Z(n7756) );
  XOR U139 ( .A(n7975), .B(n7953), .Z(n7879) );
  XOR U140 ( .A(n8134), .B(n8112), .Z(n8039) );
  XOR U141 ( .A(n8292), .B(n8270), .Z(n8197) );
  XOR U142 ( .A(n8450), .B(n8428), .Z(n8355) );
  XOR U143 ( .A(n8924), .B(n8902), .Z(n8828) );
  XOR U144 ( .A(n9048), .B(n9026), .Z(n8988) );
  XNOR U145 ( .A(n9189), .B(n9188), .Z(n9131) );
  XNOR U146 ( .A(n9269), .B(n9268), .Z(n9211) );
  XNOR U147 ( .A(n9344), .B(n9343), .Z(n9287) );
  XOR U148 ( .A(n3066), .B(n3085), .Z(n3070) );
  XOR U149 ( .A(n3225), .B(n3244), .Z(n3229) );
  XOR U150 ( .A(n9732), .B(n9806), .Z(n9736) );
  XOR U151 ( .A(n9591), .B(n9636), .Z(n9596) );
  XNOR U152 ( .A(n3032), .B(n2949), .Z(n2951) );
  XOR U153 ( .A(n3659), .B(n3727), .Z(n3664) );
  XOR U154 ( .A(n3896), .B(n3964), .Z(n3901) );
  XOR U155 ( .A(n4872), .B(n4940), .Z(n4877) );
  XOR U156 ( .A(n5109), .B(n5177), .Z(n5114) );
  XOR U157 ( .A(n6091), .B(n6159), .Z(n6096) );
  XOR U158 ( .A(n6328), .B(n6397), .Z(n6333) );
  XOR U159 ( .A(n7316), .B(n7384), .Z(n7321) );
  XOR U160 ( .A(n7554), .B(n7623), .Z(n7559) );
  XOR U161 ( .A(n8152), .B(n8220), .Z(n8161) );
  XOR U162 ( .A(n8786), .B(n8855), .Z(n8791) );
  XOR U163 ( .A(n9438), .B(n9484), .Z(n9443) );
  XOR U164 ( .A(n720), .B(n787), .Z(n724) );
  XOR U165 ( .A(n890), .B(n956), .Z(n894) );
  XOR U166 ( .A(n1059), .B(n1125), .Z(n1063) );
  XOR U167 ( .A(n1228), .B(n1294), .Z(n1232) );
  XOR U168 ( .A(n1397), .B(n1469), .Z(n1401) );
  XOR U169 ( .A(n1573), .B(n1641), .Z(n1577) );
  XOR U170 ( .A(n1745), .B(n1813), .Z(n1749) );
  XOR U171 ( .A(n2003), .B(n2071), .Z(n2007) );
  XNOR U172 ( .A(n3275), .B(n3193), .Z(n3195) );
  XOR U173 ( .A(n3823), .B(n3884), .Z(n3827) );
  XOR U174 ( .A(n4244), .B(n4305), .Z(n4248) );
  XNOR U175 ( .A(n4488), .B(n4406), .Z(n4408) );
  XOR U176 ( .A(n5036), .B(n5097), .Z(n5040) );
  XOR U177 ( .A(n5463), .B(n5524), .Z(n5467) );
  XNOR U178 ( .A(n5707), .B(n5625), .Z(n5627) );
  XOR U179 ( .A(n6255), .B(n6316), .Z(n6259) );
  XOR U180 ( .A(n6688), .B(n6749), .Z(n6692) );
  XNOR U181 ( .A(n6932), .B(n6850), .Z(n6852) );
  XOR U182 ( .A(n7480), .B(n7542), .Z(n7484) );
  XOR U183 ( .A(n7919), .B(n7980), .Z(n7923) );
  XOR U184 ( .A(n8073), .B(n8139), .Z(n8082) );
  XOR U185 ( .A(n8395), .B(n8456), .Z(n8399) );
  XOR U186 ( .A(n8553), .B(n8614), .Z(n8557) );
  XOR U187 ( .A(n8712), .B(n8774), .Z(n8716) );
  XNOR U188 ( .A(n9162), .B(n9079), .Z(n9081) );
  XOR U189 ( .A(n3433), .B(n3488), .Z(n3441) );
  XOR U190 ( .A(n3591), .B(n3646), .Z(n3595) );
  XOR U191 ( .A(n4646), .B(n4701), .Z(n4654) );
  XOR U192 ( .A(n4804), .B(n4859), .Z(n4808) );
  XOR U193 ( .A(n5865), .B(n5920), .Z(n5873) );
  XOR U194 ( .A(n6023), .B(n6078), .Z(n6027) );
  XOR U195 ( .A(n7090), .B(n7145), .Z(n7098) );
  XOR U196 ( .A(n7248), .B(n7303), .Z(n7252) );
  XOR U197 ( .A(n9380), .B(n9424), .Z(n9389) );
  XOR U198 ( .A(n9954), .B(n10010), .Z(n9958) );
  XOR U199 ( .A(n9822), .B(n9878), .Z(n9826) );
  XOR U200 ( .A(n9663), .B(n9719), .Z(n9667) );
  XOR U201 ( .A(n561), .B(n615), .Z(n565) );
  XOR U202 ( .A(n2271), .B(n2327), .Z(n2275) );
  XOR U203 ( .A(n9321), .B(n9360), .Z(n9325) );
  XOR U204 ( .A(n9562), .B(n9577), .Z(n9566) );
  XOR U205 ( .A(n478), .B(n527), .Z(n482) );
  XOR U206 ( .A(n820), .B(n869), .Z(n824) );
  XOR U207 ( .A(n989), .B(n1038), .Z(n993) );
  XOR U208 ( .A(n1158), .B(n1207), .Z(n1162) );
  XOR U209 ( .A(n1327), .B(n1376), .Z(n1331) );
  XOR U210 ( .A(n1502), .B(n1552), .Z(n1506) );
  XOR U211 ( .A(n1674), .B(n1724), .Z(n1678) );
  XOR U212 ( .A(n1846), .B(n1896), .Z(n1850) );
  XOR U213 ( .A(n2018), .B(n2068), .Z(n2022) );
  XOR U214 ( .A(n2868), .B(n2924), .Z(n2872) );
  XNOR U215 ( .A(n3211), .B(n3129), .Z(n3131) );
  XNOR U216 ( .A(n3290), .B(n3208), .Z(n3210) );
  XNOR U217 ( .A(n3369), .B(n3287), .Z(n3289) );
  XNOR U218 ( .A(n3448), .B(n3366), .Z(n3368) );
  XNOR U219 ( .A(n3527), .B(n3445), .Z(n3447) );
  XOR U220 ( .A(n3917), .B(n3960), .Z(n3921) );
  XNOR U221 ( .A(n4265), .B(n4182), .Z(n4184) );
  XNOR U222 ( .A(n4345), .B(n4262), .Z(n4264) );
  XNOR U223 ( .A(n4424), .B(n4342), .Z(n4344) );
  XNOR U224 ( .A(n4503), .B(n4421), .Z(n4423) );
  XNOR U225 ( .A(n4582), .B(n4500), .Z(n4502) );
  XNOR U226 ( .A(n4661), .B(n4579), .Z(n4581) );
  XNOR U227 ( .A(n4740), .B(n4658), .Z(n4660) );
  XOR U228 ( .A(n5130), .B(n5173), .Z(n5134) );
  XNOR U229 ( .A(n5484), .B(n5401), .Z(n5403) );
  XNOR U230 ( .A(n5564), .B(n5481), .Z(n5483) );
  XNOR U231 ( .A(n5643), .B(n5561), .Z(n5563) );
  XNOR U232 ( .A(n5722), .B(n5640), .Z(n5642) );
  XNOR U233 ( .A(n5801), .B(n5719), .Z(n5721) );
  XNOR U234 ( .A(n5880), .B(n5798), .Z(n5800) );
  XNOR U235 ( .A(n5959), .B(n5877), .Z(n5879) );
  XOR U236 ( .A(n6349), .B(n6393), .Z(n6353) );
  XNOR U237 ( .A(n6709), .B(n6626), .Z(n6628) );
  XNOR U238 ( .A(n6789), .B(n6706), .Z(n6708) );
  XNOR U239 ( .A(n6868), .B(n6786), .Z(n6788) );
  XNOR U240 ( .A(n6947), .B(n6865), .Z(n6867) );
  XNOR U241 ( .A(n7026), .B(n6944), .Z(n6946) );
  XNOR U242 ( .A(n7105), .B(n7023), .Z(n7025) );
  XNOR U243 ( .A(n7184), .B(n7102), .Z(n7104) );
  XOR U244 ( .A(n7575), .B(n7619), .Z(n7579) );
  XNOR U245 ( .A(n7940), .B(n7857), .Z(n7859) );
  XNOR U246 ( .A(n8020), .B(n7937), .Z(n7939) );
  XNOR U247 ( .A(n8099), .B(n8017), .Z(n8019) );
  XNOR U248 ( .A(n8178), .B(n8096), .Z(n8098) );
  XNOR U249 ( .A(n8257), .B(n8175), .Z(n8177) );
  XNOR U250 ( .A(n8336), .B(n8254), .Z(n8256) );
  XNOR U251 ( .A(n8415), .B(n8333), .Z(n8335) );
  XOR U252 ( .A(n8489), .B(n8532), .Z(n8493) );
  XOR U253 ( .A(n8647), .B(n8691), .Z(n8652) );
  XOR U254 ( .A(n8807), .B(n8851), .Z(n8812) );
  XNOR U255 ( .A(n9095), .B(n9094), .Z(n9050) );
  XNOR U256 ( .A(n9175), .B(n9174), .Z(n9134) );
  XNOR U257 ( .A(n9255), .B(n9254), .Z(n9214) );
  XNOR U258 ( .A(n9330), .B(n9329), .Z(n9290) );
  XNOR U259 ( .A(n9462), .B(n9461), .Z(n9422) );
  XOR U260 ( .A(n3051), .B(n3088), .Z(n3055) );
  XOR U261 ( .A(n3843), .B(n3880), .Z(n3847) );
  XOR U262 ( .A(n5056), .B(n5093), .Z(n5060) );
  XOR U263 ( .A(n6275), .B(n6312), .Z(n6279) );
  XOR U264 ( .A(n7500), .B(n7538), .Z(n7505) );
  XOR U265 ( .A(n10122), .B(n10160), .Z(n10126) );
  XOR U266 ( .A(n10026), .B(n10064), .Z(n10030) );
  XOR U267 ( .A(n9906), .B(n9944), .Z(n9910) );
  XOR U268 ( .A(n9762), .B(n9800), .Z(n9766) );
  XOR U269 ( .A(n9572), .B(n9630), .Z(n9528) );
  XOR U270 ( .A(n2286), .B(n2324), .Z(n2290) );
  XOR U271 ( .A(n333), .B(n363), .Z(n337) );
  XOR U272 ( .A(n493), .B(n524), .Z(n497) );
  XOR U273 ( .A(n665), .B(n696), .Z(n669) );
  XOR U274 ( .A(n835), .B(n866), .Z(n839) );
  XOR U275 ( .A(n1004), .B(n1035), .Z(n1008) );
  XOR U276 ( .A(n1173), .B(n1204), .Z(n1177) );
  XOR U277 ( .A(n1342), .B(n1373), .Z(n1346) );
  XOR U278 ( .A(n1517), .B(n1549), .Z(n1521) );
  XOR U279 ( .A(n1689), .B(n1721), .Z(n1693) );
  XOR U280 ( .A(n1861), .B(n1893), .Z(n1865) );
  XOR U281 ( .A(n2033), .B(n2065), .Z(n2037) );
  XOR U282 ( .A(n2205), .B(n2237), .Z(n2209) );
  XNOR U283 ( .A(n3463), .B(n3381), .Z(n3383) );
  XNOR U284 ( .A(n3542), .B(n3460), .Z(n3462) );
  XNOR U285 ( .A(n3621), .B(n3539), .Z(n3541) );
  XNOR U286 ( .A(n3700), .B(n3618), .Z(n3620) );
  XNOR U287 ( .A(n3779), .B(n3697), .Z(n3699) );
  XNOR U288 ( .A(n3778), .B(n3799), .Z(n3773) );
  XOR U289 ( .A(n4090), .B(n4131), .Z(n4094) );
  XNOR U290 ( .A(n4280), .B(n4197), .Z(n4199) );
  XNOR U291 ( .A(n4360), .B(n4277), .Z(n4279) );
  XNOR U292 ( .A(n4439), .B(n4357), .Z(n4359) );
  XNOR U293 ( .A(n4518), .B(n4436), .Z(n4438) );
  XNOR U294 ( .A(n4597), .B(n4515), .Z(n4517) );
  XNOR U295 ( .A(n4676), .B(n4594), .Z(n4596) );
  XNOR U296 ( .A(n4755), .B(n4673), .Z(n4675) );
  XNOR U297 ( .A(n4834), .B(n4752), .Z(n4754) );
  XNOR U298 ( .A(n4913), .B(n4831), .Z(n4833) );
  XNOR U299 ( .A(n4992), .B(n4910), .Z(n4912) );
  XNOR U300 ( .A(n4991), .B(n5012), .Z(n4986) );
  XOR U301 ( .A(n5304), .B(n5331), .Z(n5310) );
  XNOR U302 ( .A(n5417), .B(n5416), .Z(n5351) );
  XNOR U303 ( .A(n5497), .B(n5496), .Z(n5438) );
  XNOR U304 ( .A(n5577), .B(n5576), .Z(n5518) );
  XNOR U305 ( .A(n5656), .B(n5655), .Z(n5598) );
  XNOR U306 ( .A(n5735), .B(n5734), .Z(n5677) );
  XNOR U307 ( .A(n5814), .B(n5813), .Z(n5756) );
  XNOR U308 ( .A(n5893), .B(n5892), .Z(n5835) );
  XNOR U309 ( .A(n5972), .B(n5971), .Z(n5914) );
  XNOR U310 ( .A(n6051), .B(n6050), .Z(n5993) );
  XNOR U311 ( .A(n6130), .B(n6129), .Z(n6072) );
  XNOR U312 ( .A(n6206), .B(n6204), .Z(n6151) );
  XOR U313 ( .A(n6546), .B(n6524), .Z(n6450) );
  XNOR U314 ( .A(n6555), .B(n6554), .Z(n6545) );
  XNOR U315 ( .A(n6641), .B(n6640), .Z(n6577) );
  XNOR U316 ( .A(n6721), .B(n6720), .Z(n6663) );
  XNOR U317 ( .A(n6801), .B(n6800), .Z(n6743) );
  XNOR U318 ( .A(n6880), .B(n6879), .Z(n6823) );
  XNOR U319 ( .A(n6959), .B(n6958), .Z(n6902) );
  XNOR U320 ( .A(n7038), .B(n7037), .Z(n6981) );
  XNOR U321 ( .A(n7117), .B(n7116), .Z(n7060) );
  XNOR U322 ( .A(n7196), .B(n7195), .Z(n7139) );
  XNOR U323 ( .A(n7275), .B(n7274), .Z(n7218) );
  XNOR U324 ( .A(n7353), .B(n7351), .Z(n7297) );
  XOR U325 ( .A(n7692), .B(n7670), .Z(n7596) );
  XNOR U326 ( .A(n7749), .B(n7748), .Z(n7691) );
  XNOR U327 ( .A(n7787), .B(n7786), .Z(n7771) );
  XNOR U328 ( .A(n7872), .B(n7871), .Z(n7809) );
  XNOR U329 ( .A(n7952), .B(n7951), .Z(n7894) );
  XNOR U330 ( .A(n8032), .B(n8031), .Z(n7974) );
  XNOR U331 ( .A(n8111), .B(n8110), .Z(n8054) );
  XNOR U332 ( .A(n8190), .B(n8189), .Z(n8133) );
  XNOR U333 ( .A(n8269), .B(n8268), .Z(n8212) );
  XNOR U334 ( .A(n8348), .B(n8347), .Z(n8291) );
  XNOR U335 ( .A(n8427), .B(n8426), .Z(n8370) );
  XNOR U336 ( .A(n8506), .B(n8504), .Z(n8449) );
  XOR U337 ( .A(n8684), .B(n8661), .Z(n8588) );
  XOR U338 ( .A(n8844), .B(n8822), .Z(n8748) );
  XNOR U339 ( .A(n8901), .B(n8900), .Z(n8843) );
  XNOR U340 ( .A(n8981), .B(n8980), .Z(n8923) );
  XNOR U341 ( .A(n9025), .B(n9024), .Z(n9003) );
  XNOR U342 ( .A(n9109), .B(n9108), .Z(n9047) );
  XOR U343 ( .A(n9212), .B(n9190), .Z(n9116) );
  XOR U344 ( .A(n9357), .B(n9345), .Z(n9276) );
  XOR U345 ( .A(n2986), .B(n3005), .Z(n2990) );
  XOR U346 ( .A(n3146), .B(n3165), .Z(n3150) );
  XOR U347 ( .A(n3304), .B(n3323), .Z(n3308) );
  XOR U348 ( .A(n3937), .B(n3956), .Z(n3942) );
  XOR U349 ( .A(n5165), .B(n5149), .Z(n5077) );
  XOR U350 ( .A(n6305), .B(n6289), .Z(n6218) );
  XOR U351 ( .A(n7451), .B(n7435), .Z(n7365) );
  XNOR U352 ( .A(n9274), .B(n9273), .Z(n9210) );
  XNOR U353 ( .A(n10236), .B(n10256), .Z(n10244) );
  XNOR U354 ( .A(n10176), .B(n10196), .Z(n10184) );
  XNOR U355 ( .A(n10092), .B(n10112), .Z(n10100) );
  XNOR U356 ( .A(n9984), .B(n10004), .Z(n9992) );
  XNOR U357 ( .A(n9852), .B(n9872), .Z(n9860) );
  XNOR U358 ( .A(n9693), .B(n9713), .Z(n9701) );
  XOR U359 ( .A(n9647), .B(n9722), .Z(n9652) );
  XOR U360 ( .A(n1911), .B(n1986), .Z(n1916) );
  XOR U361 ( .A(n2083), .B(n2158), .Z(n2088) );
  XOR U362 ( .A(n2255), .B(n2330), .Z(n2260) );
  XOR U363 ( .A(n8389), .B(n8457), .Z(n8394) );
  XNOR U364 ( .A(n9310), .B(n9364), .Z(n9306) );
  XOR U365 ( .A(n9546), .B(n9580), .Z(n9551) );
  XOR U366 ( .A(n462), .B(n530), .Z(n467) );
  XOR U367 ( .A(n635), .B(n702), .Z(n639) );
  XOR U368 ( .A(n805), .B(n872), .Z(n809) );
  XOR U369 ( .A(n974), .B(n1041), .Z(n978) );
  XOR U370 ( .A(n1143), .B(n1210), .Z(n1147) );
  XOR U371 ( .A(n1312), .B(n1379), .Z(n1316) );
  XOR U372 ( .A(n1487), .B(n1555), .Z(n1491) );
  XOR U373 ( .A(n1659), .B(n1727), .Z(n1663) );
  XOR U374 ( .A(n1831), .B(n1899), .Z(n1835) );
  XOR U375 ( .A(n2853), .B(n2930), .Z(n2857) );
  XNOR U376 ( .A(n3037), .B(n2954), .Z(n2956) );
  XNOR U377 ( .A(n3117), .B(n3034), .Z(n3036) );
  XNOR U378 ( .A(n3196), .B(n3114), .Z(n3116) );
  XOR U379 ( .A(n3185), .B(n3251), .Z(n3194) );
  XOR U380 ( .A(n3349), .B(n3410), .Z(n3357) );
  XOR U381 ( .A(n3665), .B(n3726), .Z(n3669) );
  XOR U382 ( .A(n3902), .B(n3963), .Z(n3906) );
  XOR U383 ( .A(n4060), .B(n4143), .Z(n4064) );
  XNOR U384 ( .A(n4250), .B(n4167), .Z(n4169) );
  XNOR U385 ( .A(n4330), .B(n4247), .Z(n4249) );
  XNOR U386 ( .A(n4409), .B(n4327), .Z(n4329) );
  XOR U387 ( .A(n4398), .B(n4464), .Z(n4407) );
  XOR U388 ( .A(n4562), .B(n4623), .Z(n4570) );
  XOR U389 ( .A(n4878), .B(n4939), .Z(n4882) );
  XOR U390 ( .A(n5115), .B(n5176), .Z(n5119) );
  XOR U391 ( .A(n5274), .B(n5362), .Z(n5278) );
  XNOR U392 ( .A(n5469), .B(n5386), .Z(n5388) );
  XNOR U393 ( .A(n5549), .B(n5466), .Z(n5468) );
  XNOR U394 ( .A(n5628), .B(n5546), .Z(n5548) );
  XOR U395 ( .A(n5617), .B(n5683), .Z(n5626) );
  XOR U396 ( .A(n5781), .B(n5842), .Z(n5789) );
  XOR U397 ( .A(n6097), .B(n6158), .Z(n6101) );
  XOR U398 ( .A(n6334), .B(n6396), .Z(n6338) );
  XOR U399 ( .A(n6494), .B(n6587), .Z(n6498) );
  XNOR U400 ( .A(n6694), .B(n6611), .Z(n6613) );
  XNOR U401 ( .A(n6774), .B(n6691), .Z(n6693) );
  XNOR U402 ( .A(n6853), .B(n6771), .Z(n6773) );
  XOR U403 ( .A(n6842), .B(n6908), .Z(n6851) );
  XOR U404 ( .A(n7006), .B(n7067), .Z(n7014) );
  XOR U405 ( .A(n7322), .B(n7383), .Z(n7326) );
  XOR U406 ( .A(n7560), .B(n7622), .Z(n7564) );
  XOR U407 ( .A(n7720), .B(n7818), .Z(n7724) );
  XNOR U408 ( .A(n7925), .B(n7842), .Z(n7844) );
  XNOR U409 ( .A(n8005), .B(n7922), .Z(n7924) );
  XNOR U410 ( .A(n8084), .B(n8002), .Z(n8004) );
  XNOR U411 ( .A(n8163), .B(n8081), .Z(n8083) );
  XNOR U412 ( .A(n8162), .B(n8219), .Z(n8157) );
  XOR U413 ( .A(n8792), .B(n8854), .Z(n8796) );
  XOR U414 ( .A(n8952), .B(n9055), .Z(n8956) );
  XOR U415 ( .A(n9076), .B(n9137), .Z(n9080) );
  XOR U416 ( .A(n8321), .B(n8376), .Z(n8329) );
  XOR U417 ( .A(n8637), .B(n8693), .Z(n8641) );
  XOR U418 ( .A(n9506), .B(n9533), .Z(n9514) );
  XOR U419 ( .A(n9891), .B(n9947), .Z(n9895) );
  XOR U420 ( .A(n9747), .B(n9803), .Z(n9751) );
  XOR U421 ( .A(n9607), .B(n9633), .Z(n9615) );
  XOR U422 ( .A(n2185), .B(n2241), .Z(n2189) );
  XOR U423 ( .A(n2357), .B(n2833), .Z(n2361) );
  XOR U424 ( .A(n8563), .B(n8612), .Z(n8567) );
  XNOR U425 ( .A(n9396), .B(n9324), .Z(n9326) );
  XNOR U426 ( .A(n9459), .B(n9393), .Z(n9395) );
  XOR U427 ( .A(n9448), .B(n9480), .Z(n9457) );
  XOR U428 ( .A(n393), .B(n447), .Z(n397) );
  XOR U429 ( .A(n566), .B(n614), .Z(n570) );
  XOR U430 ( .A(n735), .B(n784), .Z(n739) );
  XOR U431 ( .A(n905), .B(n953), .Z(n909) );
  XOR U432 ( .A(n1074), .B(n1122), .Z(n1078) );
  XOR U433 ( .A(n1243), .B(n1291), .Z(n1247) );
  XOR U434 ( .A(n1412), .B(n1466), .Z(n1416) );
  XOR U435 ( .A(n1588), .B(n1638), .Z(n1592) );
  XOR U436 ( .A(n1760), .B(n1810), .Z(n1764) );
  XOR U437 ( .A(n1932), .B(n1982), .Z(n1936) );
  XOR U438 ( .A(n2104), .B(n2154), .Z(n2108) );
  XOR U439 ( .A(n3126), .B(n3169), .Z(n3130) );
  XNOR U440 ( .A(n3526), .B(n3565), .Z(n3521) );
  XOR U441 ( .A(n3759), .B(n3802), .Z(n3763) );
  XOR U442 ( .A(n3996), .B(n4039), .Z(n4000) );
  XNOR U443 ( .A(n4739), .B(n4778), .Z(n4734) );
  XOR U444 ( .A(n4972), .B(n5015), .Z(n4976) );
  XOR U445 ( .A(n5209), .B(n5253), .Z(n5213) );
  XNOR U446 ( .A(n5958), .B(n5997), .Z(n5953) );
  XOR U447 ( .A(n6191), .B(n6234), .Z(n6195) );
  XOR U448 ( .A(n6429), .B(n6473), .Z(n6433) );
  XNOR U449 ( .A(n7183), .B(n7222), .Z(n7178) );
  XOR U450 ( .A(n7416), .B(n7459), .Z(n7420) );
  XOR U451 ( .A(n7655), .B(n7699), .Z(n7659) );
  XOR U452 ( .A(n8887), .B(n8931), .Z(n8892) );
  XNOR U453 ( .A(n3216), .B(n3134), .Z(n3136) );
  XNOR U454 ( .A(n3374), .B(n3292), .Z(n3294) );
  XNOR U455 ( .A(n3453), .B(n3371), .Z(n3373) );
  XNOR U456 ( .A(n3532), .B(n3450), .Z(n3452) );
  XNOR U457 ( .A(n3611), .B(n3529), .Z(n3531) );
  XOR U458 ( .A(n3685), .B(n3722), .Z(n3693) );
  XOR U459 ( .A(n3922), .B(n3959), .Z(n3926) );
  XNOR U460 ( .A(n4270), .B(n4187), .Z(n4189) );
  XNOR U461 ( .A(n4350), .B(n4267), .Z(n4269) );
  XNOR U462 ( .A(n4429), .B(n4347), .Z(n4349) );
  XNOR U463 ( .A(n4508), .B(n4426), .Z(n4428) );
  XNOR U464 ( .A(n4587), .B(n4505), .Z(n4507) );
  XNOR U465 ( .A(n4666), .B(n4584), .Z(n4586) );
  XNOR U466 ( .A(n4745), .B(n4663), .Z(n4665) );
  XNOR U467 ( .A(n4824), .B(n4742), .Z(n4744) );
  XOR U468 ( .A(n4898), .B(n4935), .Z(n4906) );
  XOR U469 ( .A(n5135), .B(n5172), .Z(n5139) );
  XNOR U470 ( .A(n5489), .B(n5406), .Z(n5408) );
  XNOR U471 ( .A(n5569), .B(n5486), .Z(n5488) );
  XNOR U472 ( .A(n5648), .B(n5566), .Z(n5568) );
  XNOR U473 ( .A(n5727), .B(n5645), .Z(n5647) );
  XNOR U474 ( .A(n5806), .B(n5724), .Z(n5726) );
  XNOR U475 ( .A(n5885), .B(n5803), .Z(n5805) );
  XNOR U476 ( .A(n5964), .B(n5882), .Z(n5884) );
  XNOR U477 ( .A(n6043), .B(n5961), .Z(n5963) );
  XOR U478 ( .A(n6117), .B(n6154), .Z(n6125) );
  XOR U479 ( .A(n6354), .B(n6392), .Z(n6358) );
  XNOR U480 ( .A(n6714), .B(n6631), .Z(n6633) );
  XNOR U481 ( .A(n6794), .B(n6711), .Z(n6713) );
  XNOR U482 ( .A(n6873), .B(n6791), .Z(n6793) );
  XNOR U483 ( .A(n6952), .B(n6870), .Z(n6872) );
  XNOR U484 ( .A(n7031), .B(n6949), .Z(n6951) );
  XNOR U485 ( .A(n7110), .B(n7028), .Z(n7030) );
  XNOR U486 ( .A(n7189), .B(n7107), .Z(n7109) );
  XNOR U487 ( .A(n7268), .B(n7186), .Z(n7188) );
  XOR U488 ( .A(n7342), .B(n7379), .Z(n7346) );
  XOR U489 ( .A(n7580), .B(n7618), .Z(n7585) );
  XNOR U490 ( .A(n7863), .B(n7862), .Z(n7811) );
  XNOR U491 ( .A(n7943), .B(n7942), .Z(n7896) );
  XNOR U492 ( .A(n8023), .B(n8022), .Z(n7976) );
  XNOR U493 ( .A(n8102), .B(n8101), .Z(n8056) );
  XNOR U494 ( .A(n8181), .B(n8180), .Z(n8135) );
  XNOR U495 ( .A(n8260), .B(n8259), .Z(n8214) );
  XNOR U496 ( .A(n8339), .B(n8338), .Z(n8293) );
  XOR U497 ( .A(n8409), .B(n8419), .Z(n8345) );
  XOR U498 ( .A(n8846), .B(n8811), .Z(n8737) );
  XNOR U499 ( .A(n9015), .B(n9014), .Z(n9005) );
  XNOR U500 ( .A(n9099), .B(n9098), .Z(n9049) );
  XNOR U501 ( .A(n9179), .B(n9178), .Z(n9133) );
  XNOR U502 ( .A(n9259), .B(n9258), .Z(n9213) );
  XNOR U503 ( .A(n9334), .B(n9333), .Z(n9289) );
  XOR U504 ( .A(n10077), .B(n10115), .Z(n10081) );
  XOR U505 ( .A(n9969), .B(n10007), .Z(n9973) );
  XOR U506 ( .A(n9837), .B(n9875), .Z(n9841) );
  XOR U507 ( .A(n9678), .B(n9716), .Z(n9682) );
  XOR U508 ( .A(n2372), .B(n2830), .Z(n2376) );
  XOR U509 ( .A(n3056), .B(n3087), .Z(n3060) );
  XOR U510 ( .A(n8605), .B(n8577), .Z(n8505) );
  XNOR U511 ( .A(n9408), .B(n9407), .Z(n9357) );
  XOR U512 ( .A(n9478), .B(n9472), .Z(n9415) );
  XOR U513 ( .A(n413), .B(n443), .Z(n417) );
  XOR U514 ( .A(n581), .B(n611), .Z(n585) );
  XOR U515 ( .A(n750), .B(n781), .Z(n754) );
  XOR U516 ( .A(n920), .B(n950), .Z(n924) );
  XOR U517 ( .A(n1089), .B(n1119), .Z(n1093) );
  XOR U518 ( .A(n1258), .B(n1288), .Z(n1262) );
  XOR U519 ( .A(n1427), .B(n1463), .Z(n1431) );
  XOR U520 ( .A(n1603), .B(n1635), .Z(n1607) );
  XOR U521 ( .A(n1775), .B(n1807), .Z(n1779) );
  XOR U522 ( .A(n1947), .B(n1979), .Z(n1951) );
  XOR U523 ( .A(n2119), .B(n2151), .Z(n2123) );
  XOR U524 ( .A(n2291), .B(n2323), .Z(n2295) );
  XNOR U525 ( .A(n3468), .B(n3386), .Z(n3388) );
  XNOR U526 ( .A(n3547), .B(n3465), .Z(n3467) );
  XNOR U527 ( .A(n3626), .B(n3544), .Z(n3546) );
  XNOR U528 ( .A(n3705), .B(n3623), .Z(n3625) );
  XNOR U529 ( .A(n3784), .B(n3702), .Z(n3704) );
  XNOR U530 ( .A(n3863), .B(n3781), .Z(n3783) );
  XOR U531 ( .A(n4016), .B(n4035), .Z(n4021) );
  XNOR U532 ( .A(n4203), .B(n4202), .Z(n4130) );
  XNOR U533 ( .A(n4283), .B(n4282), .Z(n4218) );
  XNOR U534 ( .A(n4363), .B(n4362), .Z(n4298) );
  XNOR U535 ( .A(n4442), .B(n4441), .Z(n4378) );
  XNOR U536 ( .A(n4521), .B(n4520), .Z(n4457) );
  XNOR U537 ( .A(n4600), .B(n4599), .Z(n4536) );
  XNOR U538 ( .A(n4679), .B(n4678), .Z(n4615) );
  XNOR U539 ( .A(n4758), .B(n4757), .Z(n4694) );
  XNOR U540 ( .A(n4837), .B(n4836), .Z(n4773) );
  XNOR U541 ( .A(n4916), .B(n4915), .Z(n4852) );
  XNOR U542 ( .A(n4995), .B(n4994), .Z(n4931) );
  XOR U543 ( .A(n5245), .B(n5228), .Z(n5155) );
  XNOR U544 ( .A(n5334), .B(n5333), .Z(n5324) );
  XNOR U545 ( .A(n5421), .B(n5420), .Z(n5350) );
  XNOR U546 ( .A(n5501), .B(n5500), .Z(n5437) );
  XNOR U547 ( .A(n5581), .B(n5580), .Z(n5517) );
  XNOR U548 ( .A(n5660), .B(n5659), .Z(n5597) );
  XNOR U549 ( .A(n5739), .B(n5738), .Z(n5676) );
  XNOR U550 ( .A(n5818), .B(n5817), .Z(n5755) );
  XNOR U551 ( .A(n5897), .B(n5896), .Z(n5834) );
  XNOR U552 ( .A(n5976), .B(n5975), .Z(n5913) );
  XNOR U553 ( .A(n6055), .B(n6054), .Z(n5992) );
  XNOR U554 ( .A(n6134), .B(n6133), .Z(n6071) );
  XOR U555 ( .A(n6385), .B(n6368), .Z(n6295) );
  XNOR U556 ( .A(n6528), .B(n6527), .Z(n6464) );
  XNOR U557 ( .A(n6560), .B(n6559), .Z(n6544) );
  XNOR U558 ( .A(n6646), .B(n6645), .Z(n6576) );
  XNOR U559 ( .A(n6726), .B(n6725), .Z(n6662) );
  XNOR U560 ( .A(n6806), .B(n6805), .Z(n6742) );
  XNOR U561 ( .A(n6885), .B(n6884), .Z(n6822) );
  XNOR U562 ( .A(n6964), .B(n6963), .Z(n6901) );
  XNOR U563 ( .A(n7043), .B(n7042), .Z(n6980) );
  XNOR U564 ( .A(n7122), .B(n7121), .Z(n7059) );
  XNOR U565 ( .A(n7201), .B(n7200), .Z(n7138) );
  XNOR U566 ( .A(n7280), .B(n7279), .Z(n7217) );
  XOR U567 ( .A(n7531), .B(n7514), .Z(n7441) );
  XNOR U568 ( .A(n7674), .B(n7673), .Z(n7610) );
  XNOR U569 ( .A(n7754), .B(n7753), .Z(n7690) );
  XNOR U570 ( .A(n7792), .B(n7791), .Z(n7770) );
  XNOR U571 ( .A(n7877), .B(n7876), .Z(n7808) );
  XNOR U572 ( .A(n7957), .B(n7956), .Z(n7893) );
  XNOR U573 ( .A(n8037), .B(n8036), .Z(n7973) );
  XNOR U574 ( .A(n8116), .B(n8115), .Z(n8053) );
  XNOR U575 ( .A(n8195), .B(n8194), .Z(n8132) );
  XNOR U576 ( .A(n8274), .B(n8273), .Z(n8211) );
  XNOR U577 ( .A(n8353), .B(n8352), .Z(n8290) );
  XNOR U578 ( .A(n8432), .B(n8431), .Z(n8369) );
  XOR U579 ( .A(n8683), .B(n8666), .Z(n8593) );
  XNOR U580 ( .A(n8826), .B(n8825), .Z(n8762) );
  XNOR U581 ( .A(n8906), .B(n8905), .Z(n8842) );
  XNOR U582 ( .A(n8986), .B(n8985), .Z(n8922) );
  XNOR U583 ( .A(n9030), .B(n9029), .Z(n9002) );
  XNOR U584 ( .A(n9114), .B(n9113), .Z(n9046) );
  XNOR U585 ( .A(n9194), .B(n9193), .Z(n9130) );
  XNOR U586 ( .A(n10209), .B(n10229), .Z(n10217) );
  XNOR U587 ( .A(n10137), .B(n10157), .Z(n10145) );
  XNOR U588 ( .A(n10041), .B(n10061), .Z(n10049) );
  XNOR U589 ( .A(n9921), .B(n9941), .Z(n9929) );
  XNOR U590 ( .A(n9777), .B(n9797), .Z(n9785) );
  XNOR U591 ( .A(n9419), .B(n9627), .Z(n9354) );
  XOR U592 ( .A(n2991), .B(n2996), .Z(n2912) );
  XOR U593 ( .A(n3151), .B(n3156), .Z(n3081) );
  XOR U594 ( .A(n3309), .B(n3314), .Z(n3240) );
  XNOR U595 ( .A(n3951), .B(n3941), .Z(n3873) );
  XNOR U596 ( .A(n5086), .B(n5076), .Z(n5007) );
  XNOR U597 ( .A(n6227), .B(n6217), .Z(n6147) );
  XNOR U598 ( .A(n7374), .B(n7364), .Z(n7293) );
  XNOR U599 ( .A(n8527), .B(n8517), .Z(n8445) );
  XNOR U600 ( .A(n9279), .B(n9278), .Z(n9207) );
  XOR U601 ( .A(n2169), .B(n2244), .Z(n2174) );
  XOR U602 ( .A(n3738), .B(n3806), .Z(n3743) );
  XOR U603 ( .A(n4951), .B(n5019), .Z(n4956) );
  XOR U604 ( .A(n6170), .B(n6238), .Z(n6175) );
  XOR U605 ( .A(n7395), .B(n7463), .Z(n7400) );
  XOR U606 ( .A(n8547), .B(n8615), .Z(n8552) );
  XOR U607 ( .A(n9375), .B(n9427), .Z(n9384) );
  XOR U608 ( .A(n9495), .B(n9535), .Z(n9500) );
  XOR U609 ( .A(n9737), .B(n9805), .Z(n9741) );
  XOR U610 ( .A(n9597), .B(n9635), .Z(n9601) );
  XOR U611 ( .A(n551), .B(n617), .Z(n555) );
  XOR U612 ( .A(n1917), .B(n1985), .Z(n1921) );
  XOR U613 ( .A(n2089), .B(n2157), .Z(n2093) );
  XOR U614 ( .A(n2347), .B(n2835), .Z(n2351) );
  XOR U615 ( .A(n3507), .B(n3568), .Z(n3511) );
  XOR U616 ( .A(n4720), .B(n4781), .Z(n4724) );
  XOR U617 ( .A(n5939), .B(n6000), .Z(n5943) );
  XOR U618 ( .A(n7164), .B(n7225), .Z(n7168) );
  XOR U619 ( .A(n8316), .B(n8377), .Z(n8320) );
  XOR U620 ( .A(n382), .B(n449), .Z(n387) );
  XOR U621 ( .A(n725), .B(n786), .Z(n729) );
  XOR U622 ( .A(n895), .B(n955), .Z(n899) );
  XOR U623 ( .A(n1064), .B(n1124), .Z(n1068) );
  XOR U624 ( .A(n1233), .B(n1293), .Z(n1237) );
  XOR U625 ( .A(n1402), .B(n1468), .Z(n1406) );
  XOR U626 ( .A(n1578), .B(n1640), .Z(n1582) );
  XOR U627 ( .A(n1750), .B(n1812), .Z(n1754) );
  XNOR U628 ( .A(n3042), .B(n2959), .Z(n2961) );
  XOR U629 ( .A(n3036), .B(n3091), .Z(n3040) );
  XNOR U630 ( .A(n3201), .B(n3119), .Z(n3121) );
  XNOR U631 ( .A(n3280), .B(n3198), .Z(n3200) );
  XNOR U632 ( .A(n3359), .B(n3277), .Z(n3279) );
  XNOR U633 ( .A(n3358), .B(n3409), .Z(n3353) );
  XOR U634 ( .A(n3670), .B(n3725), .Z(n3674) );
  XOR U635 ( .A(n3986), .B(n4041), .Z(n3990) );
  XNOR U636 ( .A(n4255), .B(n4172), .Z(n4174) );
  XNOR U637 ( .A(n4335), .B(n4252), .Z(n4254) );
  XNOR U638 ( .A(n4414), .B(n4332), .Z(n4334) );
  XNOR U639 ( .A(n4493), .B(n4411), .Z(n4413) );
  XNOR U640 ( .A(n4572), .B(n4490), .Z(n4492) );
  XNOR U641 ( .A(n4571), .B(n4622), .Z(n4566) );
  XOR U642 ( .A(n4883), .B(n4938), .Z(n4887) );
  XOR U643 ( .A(n5199), .B(n5255), .Z(n5203) );
  XNOR U644 ( .A(n5474), .B(n5391), .Z(n5393) );
  XNOR U645 ( .A(n5554), .B(n5471), .Z(n5473) );
  XNOR U646 ( .A(n5633), .B(n5551), .Z(n5553) );
  XNOR U647 ( .A(n5712), .B(n5630), .Z(n5632) );
  XNOR U648 ( .A(n5791), .B(n5709), .Z(n5711) );
  XNOR U649 ( .A(n5790), .B(n5841), .Z(n5785) );
  XOR U650 ( .A(n6102), .B(n6157), .Z(n6106) );
  XOR U651 ( .A(n6419), .B(n6475), .Z(n6423) );
  XNOR U652 ( .A(n6699), .B(n6616), .Z(n6618) );
  XNOR U653 ( .A(n6779), .B(n6696), .Z(n6698) );
  XNOR U654 ( .A(n6858), .B(n6776), .Z(n6778) );
  XNOR U655 ( .A(n6937), .B(n6855), .Z(n6857) );
  XNOR U656 ( .A(n7016), .B(n6934), .Z(n6936) );
  XNOR U657 ( .A(n7015), .B(n7066), .Z(n7010) );
  XOR U658 ( .A(n7327), .B(n7382), .Z(n7331) );
  XOR U659 ( .A(n7645), .B(n7701), .Z(n7649) );
  XNOR U660 ( .A(n7930), .B(n7847), .Z(n7849) );
  XNOR U661 ( .A(n8010), .B(n7927), .Z(n7929) );
  XNOR U662 ( .A(n8089), .B(n8007), .Z(n8009) );
  XNOR U663 ( .A(n8168), .B(n8086), .Z(n8088) );
  XNOR U664 ( .A(n8247), .B(n8165), .Z(n8167) );
  XNOR U665 ( .A(n8246), .B(n8297), .Z(n8241) );
  XOR U666 ( .A(n8479), .B(n8534), .Z(n8483) );
  XOR U667 ( .A(n8877), .B(n8933), .Z(n8881) );
  XNOR U668 ( .A(n9167), .B(n9084), .Z(n9086) );
  XNOR U669 ( .A(n9247), .B(n9164), .Z(n9166) );
  XNOR U670 ( .A(n9322), .B(n9244), .Z(n9246) );
  XNOR U671 ( .A(n9391), .B(n9319), .Z(n9321) );
  XNOR U672 ( .A(n3047), .B(n2964), .Z(n2966) );
  XOR U673 ( .A(n3833), .B(n3882), .Z(n3837) );
  XOR U674 ( .A(n5046), .B(n5095), .Z(n5050) );
  XOR U675 ( .A(n6265), .B(n6314), .Z(n6269) );
  XOR U676 ( .A(n7490), .B(n7540), .Z(n7494) );
  XOR U677 ( .A(n8722), .B(n8772), .Z(n8726) );
  XNOR U678 ( .A(n9516), .B(n9456), .Z(n9458) );
  XNOR U679 ( .A(n9515), .B(n9532), .Z(n9510) );
  XOR U680 ( .A(n10016), .B(n10066), .Z(n10020) );
  XOR U681 ( .A(n9896), .B(n9946), .Z(n9900) );
  XOR U682 ( .A(n9752), .B(n9802), .Z(n9756) );
  XOR U683 ( .A(n9616), .B(n9632), .Z(n9610) );
  XOR U684 ( .A(n650), .B(n699), .Z(n654) );
  XOR U685 ( .A(n2190), .B(n2240), .Z(n2194) );
  XOR U686 ( .A(n2362), .B(n2832), .Z(n2366) );
  XOR U687 ( .A(n3601), .B(n3644), .Z(n3609) );
  XOR U688 ( .A(n4814), .B(n4857), .Z(n4822) );
  XOR U689 ( .A(n6033), .B(n6076), .Z(n6041) );
  XOR U690 ( .A(n7258), .B(n7301), .Z(n7266) );
  XOR U691 ( .A(n398), .B(n446), .Z(n402) );
  XOR U692 ( .A(n323), .B(n365), .Z(n327) );
  XOR U693 ( .A(n571), .B(n613), .Z(n575) );
  XOR U694 ( .A(n825), .B(n868), .Z(n829) );
  XOR U695 ( .A(n994), .B(n1037), .Z(n998) );
  XOR U696 ( .A(n1163), .B(n1206), .Z(n1167) );
  XOR U697 ( .A(n1332), .B(n1375), .Z(n1336) );
  XOR U698 ( .A(n1507), .B(n1551), .Z(n1511) );
  XOR U699 ( .A(n1679), .B(n1723), .Z(n1683) );
  XOR U700 ( .A(n1851), .B(n1895), .Z(n1855) );
  XOR U701 ( .A(n2023), .B(n2067), .Z(n2027) );
  XNOR U702 ( .A(n3295), .B(n3213), .Z(n3215) );
  XOR U703 ( .A(n3289), .B(n3326), .Z(n3293) );
  XOR U704 ( .A(n3368), .B(n3405), .Z(n3372) );
  XOR U705 ( .A(n3447), .B(n3484), .Z(n3451) );
  XOR U706 ( .A(n3521), .B(n3563), .Z(n3530) );
  XOR U707 ( .A(n3764), .B(n3801), .Z(n3768) );
  XOR U708 ( .A(n4080), .B(n4135), .Z(n4084) );
  XOR U709 ( .A(n4184), .B(n4221), .Z(n4188) );
  XOR U710 ( .A(n4264), .B(n4301), .Z(n4268) );
  XOR U711 ( .A(n4344), .B(n4381), .Z(n4348) );
  XOR U712 ( .A(n4423), .B(n4460), .Z(n4427) );
  XOR U713 ( .A(n4502), .B(n4539), .Z(n4506) );
  XOR U714 ( .A(n4581), .B(n4618), .Z(n4585) );
  XOR U715 ( .A(n4660), .B(n4697), .Z(n4664) );
  XOR U716 ( .A(n4734), .B(n4776), .Z(n4743) );
  XOR U717 ( .A(n4977), .B(n5014), .Z(n4981) );
  XOR U718 ( .A(n5294), .B(n5354), .Z(n5298) );
  XOR U719 ( .A(n5403), .B(n5440), .Z(n5407) );
  XOR U720 ( .A(n5483), .B(n5520), .Z(n5487) );
  XOR U721 ( .A(n5563), .B(n5600), .Z(n5567) );
  XOR U722 ( .A(n5642), .B(n5679), .Z(n5646) );
  XOR U723 ( .A(n5721), .B(n5758), .Z(n5725) );
  XOR U724 ( .A(n5800), .B(n5837), .Z(n5804) );
  XOR U725 ( .A(n5879), .B(n5916), .Z(n5883) );
  XOR U726 ( .A(n5953), .B(n5995), .Z(n5962) );
  XOR U727 ( .A(n6196), .B(n6233), .Z(n6200) );
  XOR U728 ( .A(n6514), .B(n6579), .Z(n6518) );
  XOR U729 ( .A(n6628), .B(n6665), .Z(n6632) );
  XOR U730 ( .A(n6708), .B(n6745), .Z(n6712) );
  XOR U731 ( .A(n6788), .B(n6825), .Z(n6792) );
  XOR U732 ( .A(n6867), .B(n6904), .Z(n6871) );
  XOR U733 ( .A(n6946), .B(n6983), .Z(n6950) );
  XOR U734 ( .A(n7025), .B(n7062), .Z(n7029) );
  XOR U735 ( .A(n7104), .B(n7141), .Z(n7108) );
  XOR U736 ( .A(n7178), .B(n7220), .Z(n7187) );
  XOR U737 ( .A(n7421), .B(n7458), .Z(n7426) );
  XOR U738 ( .A(n7740), .B(n7779), .Z(n7746) );
  XOR U739 ( .A(n7859), .B(n7864), .Z(n7784) );
  XOR U740 ( .A(n7939), .B(n7944), .Z(n7869) );
  XOR U741 ( .A(n8019), .B(n8024), .Z(n7949) );
  XOR U742 ( .A(n8098), .B(n8103), .Z(n8029) );
  XOR U743 ( .A(n8177), .B(n8182), .Z(n8108) );
  XOR U744 ( .A(n8256), .B(n8261), .Z(n8187) );
  XOR U745 ( .A(n8335), .B(n8340), .Z(n8266) );
  XNOR U746 ( .A(n8418), .B(n8417), .Z(n8372) );
  XNOR U747 ( .A(n8494), .B(n8492), .Z(n8451) );
  XOR U748 ( .A(n8686), .B(n8651), .Z(n8578) );
  XOR U749 ( .A(n9006), .B(n8972), .Z(n8898) );
  XOR U750 ( .A(n9050), .B(n9016), .Z(n8978) );
  XOR U751 ( .A(n9134), .B(n9100), .Z(n9022) );
  XOR U752 ( .A(n9214), .B(n9180), .Z(n9106) );
  XOR U753 ( .A(n9290), .B(n9260), .Z(n9186) );
  XOR U754 ( .A(n9359), .B(n9335), .Z(n9266) );
  XOR U755 ( .A(n2976), .B(n3007), .Z(n2980) );
  XOR U756 ( .A(n3136), .B(n3167), .Z(n3140) );
  XNOR U757 ( .A(n3300), .B(n3218), .Z(n3220) );
  XOR U758 ( .A(n3927), .B(n3958), .Z(n3931) );
  XOR U759 ( .A(n5140), .B(n5171), .Z(n5144) );
  XOR U760 ( .A(n6359), .B(n6391), .Z(n6364) );
  XOR U761 ( .A(n7613), .B(n7584), .Z(n7510) );
  XOR U762 ( .A(n8765), .B(n8736), .Z(n8662) );
  XOR U763 ( .A(n9421), .B(n9409), .Z(n9346) );
  XOR U764 ( .A(n10127), .B(n10159), .Z(n10131) );
  XOR U765 ( .A(n10031), .B(n10063), .Z(n10035) );
  XOR U766 ( .A(n9911), .B(n9943), .Z(n9915) );
  XOR U767 ( .A(n9767), .B(n9799), .Z(n9771) );
  XOR U768 ( .A(n9529), .B(n9629), .Z(n9476) );
  XOR U769 ( .A(n338), .B(n362), .Z(n342) );
  XOR U770 ( .A(n498), .B(n523), .Z(n502) );
  XOR U771 ( .A(n670), .B(n695), .Z(n674) );
  XOR U772 ( .A(n840), .B(n865), .Z(n844) );
  XOR U773 ( .A(n1009), .B(n1034), .Z(n1013) );
  XOR U774 ( .A(n1178), .B(n1203), .Z(n1182) );
  XOR U775 ( .A(n1347), .B(n1372), .Z(n1351) );
  XOR U776 ( .A(n1522), .B(n1548), .Z(n1526) );
  XOR U777 ( .A(n1694), .B(n1720), .Z(n1698) );
  XOR U778 ( .A(n1866), .B(n1892), .Z(n1870) );
  XOR U779 ( .A(n2038), .B(n2064), .Z(n2042) );
  XOR U780 ( .A(n2210), .B(n2236), .Z(n2214) );
  XOR U781 ( .A(n2382), .B(n2828), .Z(n2386) );
  XNOR U782 ( .A(n3862), .B(n3877), .Z(n3857) );
  XNOR U783 ( .A(n5071), .B(n5069), .Z(n5010) );
  XNOR U784 ( .A(n6212), .B(n6210), .Z(n6150) );
  XNOR U785 ( .A(n7359), .B(n7357), .Z(n7296) );
  XNOR U786 ( .A(n8512), .B(n8510), .Z(n8448) );
  XOR U787 ( .A(n3071), .B(n3076), .Z(n3001) );
  XOR U788 ( .A(n3230), .B(n3235), .Z(n3161) );
  XOR U789 ( .A(n3388), .B(n3393), .Z(n3319) );
  XNOR U790 ( .A(n3471), .B(n3470), .Z(n3399) );
  XNOR U791 ( .A(n3550), .B(n3549), .Z(n3478) );
  XNOR U792 ( .A(n3629), .B(n3628), .Z(n3557) );
  XNOR U793 ( .A(n3708), .B(n3707), .Z(n3636) );
  XNOR U794 ( .A(n3787), .B(n3786), .Z(n3715) );
  XNOR U795 ( .A(n3866), .B(n3865), .Z(n3794) );
  XNOR U796 ( .A(n4030), .B(n4020), .Z(n3947) );
  XNOR U797 ( .A(n4119), .B(n4118), .Z(n4107) );
  XNOR U798 ( .A(n4207), .B(n4206), .Z(n4127) );
  XNOR U799 ( .A(n4287), .B(n4286), .Z(n4215) );
  XNOR U800 ( .A(n4367), .B(n4366), .Z(n4295) );
  XNOR U801 ( .A(n4446), .B(n4445), .Z(n4375) );
  XNOR U802 ( .A(n4525), .B(n4524), .Z(n4454) );
  XNOR U803 ( .A(n4604), .B(n4603), .Z(n4533) );
  XNOR U804 ( .A(n4683), .B(n4682), .Z(n4612) );
  XNOR U805 ( .A(n4762), .B(n4761), .Z(n4691) );
  XNOR U806 ( .A(n4841), .B(n4840), .Z(n4770) );
  XNOR U807 ( .A(n4920), .B(n4919), .Z(n4849) );
  XNOR U808 ( .A(n4999), .B(n4998), .Z(n4928) );
  XNOR U809 ( .A(n5164), .B(n5154), .Z(n5082) );
  XNOR U810 ( .A(n5313), .B(n5312), .Z(n5241) );
  XNOR U811 ( .A(n5339), .B(n5338), .Z(n5321) );
  XNOR U812 ( .A(n5426), .B(n5425), .Z(n5347) );
  XNOR U813 ( .A(n5506), .B(n5505), .Z(n5434) );
  XNOR U814 ( .A(n5586), .B(n5585), .Z(n5514) );
  XNOR U815 ( .A(n5665), .B(n5664), .Z(n5594) );
  XNOR U816 ( .A(n5744), .B(n5743), .Z(n5673) );
  XNOR U817 ( .A(n5823), .B(n5822), .Z(n5752) );
  XNOR U818 ( .A(n5902), .B(n5901), .Z(n5831) );
  XNOR U819 ( .A(n5981), .B(n5980), .Z(n5910) );
  XNOR U820 ( .A(n6060), .B(n6059), .Z(n5989) );
  XNOR U821 ( .A(n6139), .B(n6138), .Z(n6068) );
  XNOR U822 ( .A(n6304), .B(n6294), .Z(n6223) );
  XNOR U823 ( .A(n6453), .B(n6452), .Z(n6381) );
  XNOR U824 ( .A(n6533), .B(n6532), .Z(n6461) );
  XNOR U825 ( .A(n6565), .B(n6564), .Z(n6541) );
  XNOR U826 ( .A(n6651), .B(n6650), .Z(n6573) );
  XNOR U827 ( .A(n6731), .B(n6730), .Z(n6659) );
  XNOR U828 ( .A(n6811), .B(n6810), .Z(n6739) );
  XNOR U829 ( .A(n6890), .B(n6889), .Z(n6819) );
  XNOR U830 ( .A(n6969), .B(n6968), .Z(n6898) );
  XNOR U831 ( .A(n7048), .B(n7047), .Z(n6977) );
  XNOR U832 ( .A(n7127), .B(n7126), .Z(n7056) );
  XNOR U833 ( .A(n7206), .B(n7205), .Z(n7135) );
  XNOR U834 ( .A(n7285), .B(n7284), .Z(n7214) );
  XNOR U835 ( .A(n7450), .B(n7440), .Z(n7370) );
  XNOR U836 ( .A(n7599), .B(n7598), .Z(n7527) );
  XNOR U837 ( .A(n7679), .B(n7678), .Z(n7607) );
  XNOR U838 ( .A(n7759), .B(n7758), .Z(n7687) );
  XNOR U839 ( .A(n7797), .B(n7796), .Z(n7767) );
  XNOR U840 ( .A(n7882), .B(n7881), .Z(n7805) );
  XNOR U841 ( .A(n7962), .B(n7961), .Z(n7890) );
  XNOR U842 ( .A(n8042), .B(n8041), .Z(n7970) );
  XNOR U843 ( .A(n8121), .B(n8120), .Z(n8050) );
  XNOR U844 ( .A(n8200), .B(n8199), .Z(n8129) );
  XNOR U845 ( .A(n8279), .B(n8278), .Z(n8208) );
  XNOR U846 ( .A(n8358), .B(n8357), .Z(n8287) );
  XNOR U847 ( .A(n8437), .B(n8436), .Z(n8366) );
  XNOR U848 ( .A(n8602), .B(n8592), .Z(n8523) );
  XNOR U849 ( .A(n8751), .B(n8750), .Z(n8679) );
  XNOR U850 ( .A(n8831), .B(n8830), .Z(n8759) );
  XNOR U851 ( .A(n8911), .B(n8910), .Z(n8839) );
  XNOR U852 ( .A(n8991), .B(n8990), .Z(n8919) );
  XNOR U853 ( .A(n9035), .B(n9034), .Z(n8999) );
  XNOR U854 ( .A(n9119), .B(n9118), .Z(n9043) );
  XNOR U855 ( .A(n9199), .B(n9198), .Z(n9127) );
  XOR U856 ( .A(n9286), .B(n9280), .Z(n9206) );
  XNOR U857 ( .A(n10279), .B(n10289), .Z(n10282) );
  XNOR U858 ( .A(n10244), .B(n10252), .Z(n10240) );
  XNOR U859 ( .A(n10184), .B(n10192), .Z(n10180) );
  XNOR U860 ( .A(n10100), .B(n10108), .Z(n10096) );
  XNOR U861 ( .A(n9992), .B(n10000), .Z(n9988) );
  XNOR U862 ( .A(n9860), .B(n9868), .Z(n9856) );
  XNOR U863 ( .A(n9701), .B(n9709), .Z(n9697) );
  AND U864 ( .A(n434), .B(n433), .Z(n353) );
  AND U865 ( .A(n771), .B(n770), .Z(n685) );
  AND U866 ( .A(n1110), .B(n1109), .Z(n1024) );
  XOR U867 ( .A(n2341), .B(n2836), .Z(n2346) );
  XOR U868 ( .A(n2945), .B(n3013), .Z(n2950) );
  XNOR U869 ( .A(n3112), .B(n3029), .Z(n3031) );
  XNOR U870 ( .A(n3189), .B(n3253), .Z(n3185) );
  XOR U871 ( .A(n3343), .B(n3411), .Z(n3348) );
  XOR U872 ( .A(n3501), .B(n3569), .Z(n3506) );
  XOR U873 ( .A(n3975), .B(n4043), .Z(n3980) );
  XOR U874 ( .A(n4158), .B(n4226), .Z(n4163) );
  XOR U875 ( .A(n4238), .B(n4306), .Z(n4243) );
  XNOR U876 ( .A(n4402), .B(n4466), .Z(n4398) );
  XOR U877 ( .A(n4556), .B(n4624), .Z(n4561) );
  XOR U878 ( .A(n4714), .B(n4782), .Z(n4719) );
  XOR U879 ( .A(n5188), .B(n5257), .Z(n5193) );
  XOR U880 ( .A(n5377), .B(n5445), .Z(n5382) );
  XOR U881 ( .A(n5457), .B(n5525), .Z(n5462) );
  XNOR U882 ( .A(n5621), .B(n5685), .Z(n5617) );
  XOR U883 ( .A(n5775), .B(n5843), .Z(n5780) );
  XOR U884 ( .A(n5933), .B(n6001), .Z(n5938) );
  XOR U885 ( .A(n6408), .B(n6477), .Z(n6413) );
  XOR U886 ( .A(n6602), .B(n6670), .Z(n6607) );
  XOR U887 ( .A(n6682), .B(n6750), .Z(n6687) );
  XNOR U888 ( .A(n6846), .B(n6910), .Z(n6842) );
  XOR U889 ( .A(n7000), .B(n7068), .Z(n7005) );
  XOR U890 ( .A(n7158), .B(n7226), .Z(n7163) );
  XOR U891 ( .A(n7634), .B(n7703), .Z(n7639) );
  XOR U892 ( .A(n7833), .B(n7901), .Z(n7838) );
  XOR U893 ( .A(n7913), .B(n7981), .Z(n7918) );
  XNOR U894 ( .A(n8077), .B(n8141), .Z(n8073) );
  XOR U895 ( .A(n8231), .B(n8299), .Z(n8236) );
  XOR U896 ( .A(n8468), .B(n8536), .Z(n8473) );
  XOR U897 ( .A(n8626), .B(n8695), .Z(n8631) );
  XOR U898 ( .A(n8866), .B(n8935), .Z(n8871) );
  XOR U899 ( .A(n9070), .B(n9138), .Z(n9075) );
  XOR U900 ( .A(n9150), .B(n9218), .Z(n9155) );
  XOR U901 ( .A(n9812), .B(n9880), .Z(n9816) );
  XOR U902 ( .A(n9653), .B(n9721), .Z(n9657) );
  XOR U903 ( .A(n9306), .B(n9362), .Z(n9315) );
  XOR U904 ( .A(n9444), .B(n9483), .Z(n9452) );
  XOR U905 ( .A(n9552), .B(n9579), .Z(n9556) );
  XOR U906 ( .A(n468), .B(n529), .Z(n472) );
  XOR U907 ( .A(n640), .B(n701), .Z(n644) );
  XOR U908 ( .A(n810), .B(n871), .Z(n814) );
  XOR U909 ( .A(n979), .B(n1040), .Z(n983) );
  XOR U910 ( .A(n1148), .B(n1209), .Z(n1152) );
  XOR U911 ( .A(n1317), .B(n1378), .Z(n1321) );
  XOR U912 ( .A(n1492), .B(n1554), .Z(n1496) );
  XOR U913 ( .A(n1664), .B(n1726), .Z(n1668) );
  XOR U914 ( .A(n1836), .B(n1898), .Z(n1840) );
  XOR U915 ( .A(n2008), .B(n2070), .Z(n2012) );
  XOR U916 ( .A(n2180), .B(n2242), .Z(n2184) );
  XOR U917 ( .A(n3749), .B(n3804), .Z(n3753) );
  XOR U918 ( .A(n4962), .B(n5017), .Z(n4966) );
  XOR U919 ( .A(n6181), .B(n6236), .Z(n6185) );
  XOR U920 ( .A(n7406), .B(n7461), .Z(n7410) );
  XOR U921 ( .A(n2863), .B(n2926), .Z(n2867) );
  XOR U922 ( .A(n2961), .B(n3010), .Z(n2965) );
  XNOR U923 ( .A(n3127), .B(n3044), .Z(n3046) );
  XNOR U924 ( .A(n3206), .B(n3124), .Z(n3126) );
  XOR U925 ( .A(n3200), .B(n3249), .Z(n3204) );
  XOR U926 ( .A(n3279), .B(n3328), .Z(n3283) );
  XOR U927 ( .A(n3353), .B(n3407), .Z(n3362) );
  XOR U928 ( .A(n3517), .B(n3566), .Z(n3525) );
  XOR U929 ( .A(n3675), .B(n3724), .Z(n3679) );
  XOR U930 ( .A(n3912), .B(n3961), .Z(n3916) );
  XOR U931 ( .A(n4070), .B(n4139), .Z(n4074) );
  XOR U932 ( .A(n4174), .B(n4223), .Z(n4178) );
  XOR U933 ( .A(n4254), .B(n4303), .Z(n4258) );
  XOR U934 ( .A(n4334), .B(n4383), .Z(n4338) );
  XOR U935 ( .A(n4413), .B(n4462), .Z(n4417) );
  XOR U936 ( .A(n4492), .B(n4541), .Z(n4496) );
  XOR U937 ( .A(n4566), .B(n4620), .Z(n4575) );
  XOR U938 ( .A(n4730), .B(n4779), .Z(n4738) );
  XOR U939 ( .A(n4888), .B(n4937), .Z(n4892) );
  XOR U940 ( .A(n5125), .B(n5174), .Z(n5129) );
  XOR U941 ( .A(n5284), .B(n5358), .Z(n5288) );
  XOR U942 ( .A(n5393), .B(n5442), .Z(n5397) );
  XOR U943 ( .A(n5473), .B(n5522), .Z(n5477) );
  XOR U944 ( .A(n5553), .B(n5602), .Z(n5557) );
  XOR U945 ( .A(n5632), .B(n5681), .Z(n5636) );
  XOR U946 ( .A(n5711), .B(n5760), .Z(n5715) );
  XOR U947 ( .A(n5785), .B(n5839), .Z(n5794) );
  XOR U948 ( .A(n5949), .B(n5998), .Z(n5957) );
  XOR U949 ( .A(n6107), .B(n6156), .Z(n6111) );
  XOR U950 ( .A(n6344), .B(n6394), .Z(n6348) );
  XOR U951 ( .A(n6504), .B(n6583), .Z(n6508) );
  XOR U952 ( .A(n6618), .B(n6667), .Z(n6622) );
  XOR U953 ( .A(n6698), .B(n6747), .Z(n6702) );
  XOR U954 ( .A(n6778), .B(n6827), .Z(n6782) );
  XOR U955 ( .A(n6857), .B(n6906), .Z(n6861) );
  XOR U956 ( .A(n6936), .B(n6985), .Z(n6940) );
  XOR U957 ( .A(n7010), .B(n7064), .Z(n7019) );
  XOR U958 ( .A(n7174), .B(n7223), .Z(n7182) );
  XOR U959 ( .A(n7332), .B(n7381), .Z(n7336) );
  XOR U960 ( .A(n7570), .B(n7620), .Z(n7574) );
  XOR U961 ( .A(n7730), .B(n7814), .Z(n7734) );
  XOR U962 ( .A(n7849), .B(n7898), .Z(n7853) );
  XOR U963 ( .A(n7929), .B(n7978), .Z(n7933) );
  XOR U964 ( .A(n8009), .B(n8058), .Z(n8013) );
  XOR U965 ( .A(n8088), .B(n8137), .Z(n8092) );
  XOR U966 ( .A(n8167), .B(n8216), .Z(n8171) );
  XNOR U967 ( .A(n8331), .B(n8249), .Z(n8251) );
  XNOR U968 ( .A(n8330), .B(n8375), .Z(n8325) );
  XOR U969 ( .A(n8484), .B(n8533), .Z(n8488) );
  XOR U970 ( .A(n8642), .B(n8692), .Z(n8646) );
  XOR U971 ( .A(n8802), .B(n8852), .Z(n8806) );
  XOR U972 ( .A(n8962), .B(n9051), .Z(n8966) );
  XOR U973 ( .A(n9086), .B(n9135), .Z(n9090) );
  XOR U974 ( .A(n9166), .B(n9215), .Z(n9170) );
  XOR U975 ( .A(n9246), .B(n9291), .Z(n9250) );
  XOR U976 ( .A(n9959), .B(n10009), .Z(n9963) );
  XOR U977 ( .A(n9827), .B(n9877), .Z(n9831) );
  XOR U978 ( .A(n9668), .B(n9718), .Z(n9672) );
  XNOR U979 ( .A(n9399), .B(n9398), .Z(n9359) );
  XOR U980 ( .A(n9458), .B(n9463), .Z(n9405) );
  XNOR U981 ( .A(n9519), .B(n9518), .Z(n9479) );
  XNOR U982 ( .A(n9567), .B(n9565), .Z(n9530) );
  XOR U983 ( .A(n308), .B(n368), .Z(n312) );
  XOR U984 ( .A(n740), .B(n783), .Z(n744) );
  XOR U985 ( .A(n910), .B(n952), .Z(n914) );
  XOR U986 ( .A(n1079), .B(n1121), .Z(n1083) );
  XOR U987 ( .A(n1248), .B(n1290), .Z(n1252) );
  XOR U988 ( .A(n1417), .B(n1465), .Z(n1421) );
  XOR U989 ( .A(n1593), .B(n1637), .Z(n1597) );
  XOR U990 ( .A(n1765), .B(n1809), .Z(n1769) );
  XOR U991 ( .A(n1937), .B(n1981), .Z(n1941) );
  XOR U992 ( .A(n2109), .B(n2153), .Z(n2113) );
  XOR U993 ( .A(n2281), .B(n2325), .Z(n2285) );
  XOR U994 ( .A(n403), .B(n445), .Z(n407) );
  XOR U995 ( .A(n660), .B(n697), .Z(n664) );
  XOR U996 ( .A(n2878), .B(n2920), .Z(n2882) );
  XNOR U997 ( .A(n3062), .B(n2979), .Z(n2981) );
  XNOR U998 ( .A(n3142), .B(n3059), .Z(n3061) );
  XNOR U999 ( .A(n3221), .B(n3139), .Z(n3141) );
  XOR U1000 ( .A(n3215), .B(n3246), .Z(n3219) );
  XNOR U1001 ( .A(n3379), .B(n3297), .Z(n3299) );
  XNOR U1002 ( .A(n3458), .B(n3376), .Z(n3378) );
  XNOR U1003 ( .A(n3537), .B(n3455), .Z(n3457) );
  XNOR U1004 ( .A(n3616), .B(n3534), .Z(n3536) );
  XNOR U1005 ( .A(n3695), .B(n3613), .Z(n3615) );
  XNOR U1006 ( .A(n3694), .B(n3721), .Z(n3689) );
  XOR U1007 ( .A(n3848), .B(n3879), .Z(n3852) );
  XOR U1008 ( .A(n4006), .B(n4037), .Z(n4010) );
  XNOR U1009 ( .A(n4275), .B(n4192), .Z(n4194) );
  XNOR U1010 ( .A(n4355), .B(n4272), .Z(n4274) );
  XNOR U1011 ( .A(n4434), .B(n4352), .Z(n4354) );
  XNOR U1012 ( .A(n4513), .B(n4431), .Z(n4433) );
  XNOR U1013 ( .A(n4592), .B(n4510), .Z(n4512) );
  XNOR U1014 ( .A(n4671), .B(n4589), .Z(n4591) );
  XNOR U1015 ( .A(n4750), .B(n4668), .Z(n4670) );
  XNOR U1016 ( .A(n4829), .B(n4747), .Z(n4749) );
  XNOR U1017 ( .A(n4908), .B(n4826), .Z(n4828) );
  XNOR U1018 ( .A(n4907), .B(n4934), .Z(n4902) );
  XOR U1019 ( .A(n5061), .B(n5092), .Z(n5065) );
  XOR U1020 ( .A(n5219), .B(n5251), .Z(n5223) );
  XNOR U1021 ( .A(n5494), .B(n5411), .Z(n5413) );
  XNOR U1022 ( .A(n5574), .B(n5491), .Z(n5493) );
  XNOR U1023 ( .A(n5653), .B(n5571), .Z(n5573) );
  XNOR U1024 ( .A(n5732), .B(n5650), .Z(n5652) );
  XNOR U1025 ( .A(n5811), .B(n5729), .Z(n5731) );
  XNOR U1026 ( .A(n5890), .B(n5808), .Z(n5810) );
  XNOR U1027 ( .A(n5969), .B(n5887), .Z(n5889) );
  XNOR U1028 ( .A(n6048), .B(n5966), .Z(n5968) );
  XNOR U1029 ( .A(n6127), .B(n6045), .Z(n6047) );
  XNOR U1030 ( .A(n6126), .B(n6153), .Z(n6121) );
  XOR U1031 ( .A(n6280), .B(n6311), .Z(n6285) );
  XOR U1032 ( .A(n6439), .B(n6471), .Z(n6444) );
  XNOR U1033 ( .A(n6637), .B(n6636), .Z(n6578) );
  XNOR U1034 ( .A(n6717), .B(n6716), .Z(n6664) );
  XNOR U1035 ( .A(n6797), .B(n6796), .Z(n6744) );
  XNOR U1036 ( .A(n6876), .B(n6875), .Z(n6824) );
  XNOR U1037 ( .A(n6955), .B(n6954), .Z(n6903) );
  XNOR U1038 ( .A(n7034), .B(n7033), .Z(n6982) );
  XNOR U1039 ( .A(n7113), .B(n7112), .Z(n7061) );
  XNOR U1040 ( .A(n7192), .B(n7191), .Z(n7140) );
  XNOR U1041 ( .A(n7271), .B(n7270), .Z(n7219) );
  XNOR U1042 ( .A(n7347), .B(n7345), .Z(n7298) );
  XOR U1043 ( .A(n7533), .B(n7504), .Z(n7431) );
  XOR U1044 ( .A(n7693), .B(n7664), .Z(n7590) );
  XNOR U1045 ( .A(n7782), .B(n7781), .Z(n7772) );
  XNOR U1046 ( .A(n7867), .B(n7866), .Z(n7810) );
  XNOR U1047 ( .A(n7947), .B(n7946), .Z(n7895) );
  XNOR U1048 ( .A(n8027), .B(n8026), .Z(n7975) );
  XNOR U1049 ( .A(n8106), .B(n8105), .Z(n8055) );
  XNOR U1050 ( .A(n8185), .B(n8184), .Z(n8134) );
  XNOR U1051 ( .A(n8264), .B(n8263), .Z(n8213) );
  XNOR U1052 ( .A(n8343), .B(n8342), .Z(n8292) );
  XNOR U1053 ( .A(n8422), .B(n8421), .Z(n8371) );
  XNOR U1054 ( .A(n8500), .B(n8498), .Z(n8450) );
  XOR U1055 ( .A(n8685), .B(n8656), .Z(n8583) );
  XOR U1056 ( .A(n8845), .B(n8816), .Z(n8742) );
  XNOR U1057 ( .A(n8976), .B(n8975), .Z(n8924) );
  XNOR U1058 ( .A(n9020), .B(n9019), .Z(n9004) );
  XNOR U1059 ( .A(n9104), .B(n9103), .Z(n9048) );
  XNOR U1060 ( .A(n9184), .B(n9183), .Z(n9132) );
  XNOR U1061 ( .A(n9264), .B(n9263), .Z(n9212) );
  XNOR U1062 ( .A(n9339), .B(n9338), .Z(n9288) );
  XOR U1063 ( .A(n10166), .B(n10198), .Z(n10170) );
  XOR U1064 ( .A(n10082), .B(n10114), .Z(n10086) );
  XOR U1065 ( .A(n9974), .B(n10006), .Z(n9978) );
  XOR U1066 ( .A(n9842), .B(n9874), .Z(n9846) );
  XOR U1067 ( .A(n9683), .B(n9715), .Z(n9687) );
  XOR U1068 ( .A(n9420), .B(n9414), .Z(n9351) );
  XOR U1069 ( .A(n418), .B(n442), .Z(n422) );
  XOR U1070 ( .A(n586), .B(n610), .Z(n590) );
  XOR U1071 ( .A(n925), .B(n949), .Z(n929) );
  XOR U1072 ( .A(n1094), .B(n1118), .Z(n1098) );
  XOR U1073 ( .A(n1263), .B(n1287), .Z(n1267) );
  XOR U1074 ( .A(n1432), .B(n1462), .Z(n1436) );
  XOR U1075 ( .A(n1608), .B(n1634), .Z(n1612) );
  XOR U1076 ( .A(n1780), .B(n1806), .Z(n1784) );
  XOR U1077 ( .A(n1952), .B(n1978), .Z(n1956) );
  XOR U1078 ( .A(n2124), .B(n2150), .Z(n2128) );
  XOR U1079 ( .A(n2296), .B(n2322), .Z(n2300) );
  XNOR U1080 ( .A(n760), .B(n779), .Z(n768) );
  XOR U1081 ( .A(n2893), .B(n2907), .Z(n2898) );
  XNOR U1082 ( .A(n2995), .B(n2994), .Z(n2913) );
  XNOR U1083 ( .A(n3075), .B(n3074), .Z(n3002) );
  XNOR U1084 ( .A(n3155), .B(n3154), .Z(n3082) );
  XNOR U1085 ( .A(n3234), .B(n3233), .Z(n3162) );
  XNOR U1086 ( .A(n3313), .B(n3312), .Z(n3241) );
  XNOR U1087 ( .A(n3392), .B(n3391), .Z(n3320) );
  XOR U1088 ( .A(n3467), .B(n3472), .Z(n3398) );
  XOR U1089 ( .A(n3546), .B(n3551), .Z(n3477) );
  XOR U1090 ( .A(n3625), .B(n3630), .Z(n3556) );
  XOR U1091 ( .A(n3704), .B(n3709), .Z(n3635) );
  XOR U1092 ( .A(n3783), .B(n3788), .Z(n3714) );
  XOR U1093 ( .A(n4110), .B(n4100), .Z(n4026) );
  XOR U1094 ( .A(n4130), .B(n4120), .Z(n4106) );
  XOR U1095 ( .A(n4218), .B(n4208), .Z(n4126) );
  XOR U1096 ( .A(n4298), .B(n4288), .Z(n4214) );
  XOR U1097 ( .A(n4378), .B(n4368), .Z(n4294) );
  XOR U1098 ( .A(n4457), .B(n4447), .Z(n4374) );
  XOR U1099 ( .A(n4536), .B(n4526), .Z(n4453) );
  XOR U1100 ( .A(n4615), .B(n4605), .Z(n4532) );
  XOR U1101 ( .A(n4694), .B(n4684), .Z(n4611) );
  XOR U1102 ( .A(n4773), .B(n4763), .Z(n4690) );
  XOR U1103 ( .A(n4852), .B(n4842), .Z(n4769) );
  XOR U1104 ( .A(n4931), .B(n4921), .Z(n4848) );
  XOR U1105 ( .A(n5244), .B(n5234), .Z(n5160) );
  XOR U1106 ( .A(n5324), .B(n5314), .Z(n5240) );
  XOR U1107 ( .A(n5350), .B(n5340), .Z(n5320) );
  XOR U1108 ( .A(n5437), .B(n5427), .Z(n5346) );
  XOR U1109 ( .A(n5517), .B(n5507), .Z(n5433) );
  XOR U1110 ( .A(n5597), .B(n5587), .Z(n5513) );
  XOR U1111 ( .A(n5676), .B(n5666), .Z(n5593) );
  XOR U1112 ( .A(n5755), .B(n5745), .Z(n5672) );
  XOR U1113 ( .A(n5834), .B(n5824), .Z(n5751) );
  XOR U1114 ( .A(n5913), .B(n5903), .Z(n5830) );
  XOR U1115 ( .A(n5992), .B(n5982), .Z(n5909) );
  XOR U1116 ( .A(n6071), .B(n6061), .Z(n5988) );
  XOR U1117 ( .A(n6384), .B(n6374), .Z(n6300) );
  XOR U1118 ( .A(n6464), .B(n6454), .Z(n6380) );
  XOR U1119 ( .A(n6544), .B(n6534), .Z(n6460) );
  XOR U1120 ( .A(n6576), .B(n6566), .Z(n6540) );
  XOR U1121 ( .A(n6662), .B(n6652), .Z(n6572) );
  XOR U1122 ( .A(n6742), .B(n6732), .Z(n6658) );
  XOR U1123 ( .A(n6822), .B(n6812), .Z(n6738) );
  XOR U1124 ( .A(n6901), .B(n6891), .Z(n6818) );
  XOR U1125 ( .A(n6980), .B(n6970), .Z(n6897) );
  XOR U1126 ( .A(n7059), .B(n7049), .Z(n6976) );
  XOR U1127 ( .A(n7138), .B(n7128), .Z(n7055) );
  XOR U1128 ( .A(n7217), .B(n7207), .Z(n7134) );
  XOR U1129 ( .A(n7530), .B(n7520), .Z(n7446) );
  XOR U1130 ( .A(n7610), .B(n7600), .Z(n7526) );
  XOR U1131 ( .A(n7690), .B(n7680), .Z(n7606) );
  XOR U1132 ( .A(n7770), .B(n7760), .Z(n7686) );
  XOR U1133 ( .A(n7808), .B(n7798), .Z(n7766) );
  XOR U1134 ( .A(n7893), .B(n7883), .Z(n7804) );
  XOR U1135 ( .A(n7973), .B(n7963), .Z(n7889) );
  XOR U1136 ( .A(n8053), .B(n8043), .Z(n7969) );
  XOR U1137 ( .A(n8132), .B(n8122), .Z(n8049) );
  XOR U1138 ( .A(n8211), .B(n8201), .Z(n8128) );
  XOR U1139 ( .A(n8290), .B(n8280), .Z(n8207) );
  XOR U1140 ( .A(n8369), .B(n8359), .Z(n8286) );
  XOR U1141 ( .A(n8448), .B(n8438), .Z(n8365) );
  XOR U1142 ( .A(n8682), .B(n8672), .Z(n8598) );
  XOR U1143 ( .A(n8762), .B(n8752), .Z(n8678) );
  XOR U1144 ( .A(n8842), .B(n8832), .Z(n8758) );
  XOR U1145 ( .A(n8922), .B(n8912), .Z(n8838) );
  XOR U1146 ( .A(n9002), .B(n8992), .Z(n8918) );
  XOR U1147 ( .A(n9046), .B(n9036), .Z(n8998) );
  XOR U1148 ( .A(n9130), .B(n9120), .Z(n9042) );
  XOR U1149 ( .A(n9210), .B(n9200), .Z(n9126) );
  XNOR U1150 ( .A(n10265), .B(n10273), .Z(n10261) );
  XNOR U1151 ( .A(n10217), .B(n10225), .Z(n10213) );
  XNOR U1152 ( .A(n10145), .B(n10153), .Z(n10141) );
  XNOR U1153 ( .A(n10049), .B(n10057), .Z(n10045) );
  XNOR U1154 ( .A(n9929), .B(n9937), .Z(n9925) );
  XNOR U1155 ( .A(n9785), .B(n9793), .Z(n9781) );
  XNOR U1156 ( .A(n9354), .B(n9623), .Z(n9285) );
  XNOR U1157 ( .A(n3873), .B(n3871), .Z(n3796) );
  XNOR U1158 ( .A(n5007), .B(n5005), .Z(n4930) );
  XNOR U1159 ( .A(n6147), .B(n6145), .Z(n6070) );
  XNOR U1160 ( .A(n7293), .B(n7291), .Z(n7216) );
  XNOR U1161 ( .A(n8523), .B(n8521), .Z(n8447) );
  AND U1162 ( .A(n514), .B(n513), .Z(n433) );
  AND U1163 ( .A(n856), .B(n855), .Z(n770) );
  AND U1164 ( .A(n1194), .B(n1193), .Z(n1109) );
  XOR U1165 ( .A(n545), .B(n618), .Z(n550) );
  XOR U1166 ( .A(n714), .B(n788), .Z(n719) );
  XOR U1167 ( .A(n884), .B(n957), .Z(n889) );
  XOR U1168 ( .A(n1053), .B(n1126), .Z(n1058) );
  XOR U1169 ( .A(n1222), .B(n1295), .Z(n1227) );
  XOR U1170 ( .A(n1391), .B(n1470), .Z(n1396) );
  XOR U1171 ( .A(n1567), .B(n1642), .Z(n1572) );
  XOR U1172 ( .A(n3025), .B(n3093), .Z(n3030) );
  XOR U1173 ( .A(n3422), .B(n3490), .Z(n3427) );
  XOR U1174 ( .A(n3580), .B(n3648), .Z(n3585) );
  XOR U1175 ( .A(n4054), .B(n4145), .Z(n4059) );
  XNOR U1176 ( .A(n4325), .B(n4242), .Z(n4244) );
  XOR U1177 ( .A(n4635), .B(n4703), .Z(n4640) );
  XOR U1178 ( .A(n4793), .B(n4861), .Z(n4798) );
  XOR U1179 ( .A(n5268), .B(n5364), .Z(n5273) );
  XNOR U1180 ( .A(n5544), .B(n5461), .Z(n5463) );
  XOR U1181 ( .A(n5854), .B(n5922), .Z(n5859) );
  XOR U1182 ( .A(n6012), .B(n6080), .Z(n6017) );
  XOR U1183 ( .A(n6488), .B(n6589), .Z(n6493) );
  XNOR U1184 ( .A(n6769), .B(n6686), .Z(n6688) );
  XOR U1185 ( .A(n7079), .B(n7147), .Z(n7084) );
  XOR U1186 ( .A(n7237), .B(n7305), .Z(n7242) );
  XOR U1187 ( .A(n7714), .B(n7820), .Z(n7719) );
  XNOR U1188 ( .A(n8000), .B(n7917), .Z(n7919) );
  XOR U1189 ( .A(n8310), .B(n8378), .Z(n8315) );
  XOR U1190 ( .A(n8706), .B(n8775), .Z(n8711) );
  XNOR U1191 ( .A(n9157), .B(n9074), .Z(n9076) );
  XNOR U1192 ( .A(n9312), .B(n9234), .Z(n9235) );
  XOR U1193 ( .A(n2951), .B(n3012), .Z(n2955) );
  XOR U1194 ( .A(n3981), .B(n4042), .Z(n3985) );
  XOR U1195 ( .A(n5194), .B(n5256), .Z(n5198) );
  XOR U1196 ( .A(n6414), .B(n6476), .Z(n6418) );
  XOR U1197 ( .A(n7640), .B(n7702), .Z(n7644) );
  XOR U1198 ( .A(n8474), .B(n8535), .Z(n8478) );
  XOR U1199 ( .A(n8632), .B(n8694), .Z(n8636) );
  XNOR U1200 ( .A(n9385), .B(n9426), .Z(n9380) );
  XOR U1201 ( .A(n9501), .B(n9534), .Z(n9505) );
  XOR U1202 ( .A(n9886), .B(n9948), .Z(n9890) );
  XOR U1203 ( .A(n9742), .B(n9804), .Z(n9746) );
  XOR U1204 ( .A(n9602), .B(n9634), .Z(n9606) );
  XOR U1205 ( .A(n1922), .B(n1984), .Z(n1926) );
  XOR U1206 ( .A(n2094), .B(n2156), .Z(n2098) );
  XOR U1207 ( .A(n2266), .B(n2328), .Z(n2270) );
  XOR U1208 ( .A(n2858), .B(n2928), .Z(n2862) );
  XOR U1209 ( .A(n3116), .B(n3171), .Z(n3120) );
  XOR U1210 ( .A(n3269), .B(n3329), .Z(n3278) );
  XOR U1211 ( .A(n3828), .B(n3883), .Z(n3832) );
  XOR U1212 ( .A(n4169), .B(n4224), .Z(n4173) );
  XOR U1213 ( .A(n4329), .B(n4384), .Z(n4333) );
  XOR U1214 ( .A(n4482), .B(n4542), .Z(n4491) );
  XOR U1215 ( .A(n5041), .B(n5096), .Z(n5045) );
  XOR U1216 ( .A(n5388), .B(n5443), .Z(n5392) );
  XOR U1217 ( .A(n5548), .B(n5603), .Z(n5552) );
  XOR U1218 ( .A(n5701), .B(n5761), .Z(n5710) );
  XOR U1219 ( .A(n6260), .B(n6315), .Z(n6264) );
  XOR U1220 ( .A(n6613), .B(n6668), .Z(n6617) );
  XOR U1221 ( .A(n6773), .B(n6828), .Z(n6777) );
  XOR U1222 ( .A(n6926), .B(n6986), .Z(n6935) );
  XOR U1223 ( .A(n7485), .B(n7541), .Z(n7489) );
  XOR U1224 ( .A(n7844), .B(n7899), .Z(n7848) );
  XOR U1225 ( .A(n8004), .B(n8059), .Z(n8008) );
  XOR U1226 ( .A(n8157), .B(n8217), .Z(n8166) );
  XOR U1227 ( .A(n8957), .B(n9053), .Z(n8961) );
  XOR U1228 ( .A(n9161), .B(n9216), .Z(n9165) );
  XOR U1229 ( .A(n9316), .B(n9361), .Z(n9320) );
  XOR U1230 ( .A(n473), .B(n528), .Z(n477) );
  XOR U1231 ( .A(n645), .B(n700), .Z(n649) );
  XOR U1232 ( .A(n815), .B(n870), .Z(n819) );
  XOR U1233 ( .A(n984), .B(n1039), .Z(n988) );
  XOR U1234 ( .A(n1153), .B(n1208), .Z(n1157) );
  XOR U1235 ( .A(n1322), .B(n1377), .Z(n1326) );
  XOR U1236 ( .A(n1497), .B(n1553), .Z(n1501) );
  XOR U1237 ( .A(n1669), .B(n1725), .Z(n1673) );
  XOR U1238 ( .A(n1841), .B(n1897), .Z(n1845) );
  XOR U1239 ( .A(n3041), .B(n3090), .Z(n3045) );
  XNOR U1240 ( .A(n3442), .B(n3487), .Z(n3437) );
  XOR U1241 ( .A(n3596), .B(n3645), .Z(n3600) );
  XOR U1242 ( .A(n3754), .B(n3803), .Z(n3758) );
  XNOR U1243 ( .A(n4655), .B(n4700), .Z(n4650) );
  XOR U1244 ( .A(n4809), .B(n4858), .Z(n4813) );
  XOR U1245 ( .A(n4967), .B(n5016), .Z(n4971) );
  XNOR U1246 ( .A(n5874), .B(n5919), .Z(n5869) );
  XOR U1247 ( .A(n6028), .B(n6077), .Z(n6032) );
  XOR U1248 ( .A(n6186), .B(n6235), .Z(n6190) );
  XNOR U1249 ( .A(n7099), .B(n7144), .Z(n7094) );
  XOR U1250 ( .A(n7253), .B(n7302), .Z(n7257) );
  XOR U1251 ( .A(n7411), .B(n7460), .Z(n7415) );
  XOR U1252 ( .A(n8405), .B(n8454), .Z(n8413) );
  XOR U1253 ( .A(n8882), .B(n8932), .Z(n8886) );
  XNOR U1254 ( .A(n3052), .B(n2969), .Z(n2971) );
  XOR U1255 ( .A(n3205), .B(n3248), .Z(n3209) );
  XOR U1256 ( .A(n3363), .B(n3406), .Z(n3367) );
  XOR U1257 ( .A(n4075), .B(n4137), .Z(n4079) );
  XOR U1258 ( .A(n4259), .B(n4302), .Z(n4263) );
  XOR U1259 ( .A(n4418), .B(n4461), .Z(n4422) );
  XOR U1260 ( .A(n4576), .B(n4619), .Z(n4580) );
  XOR U1261 ( .A(n5289), .B(n5356), .Z(n5293) );
  XOR U1262 ( .A(n5478), .B(n5521), .Z(n5482) );
  XOR U1263 ( .A(n5637), .B(n5680), .Z(n5641) );
  XOR U1264 ( .A(n5795), .B(n5838), .Z(n5799) );
  XOR U1265 ( .A(n6509), .B(n6581), .Z(n6513) );
  XOR U1266 ( .A(n6703), .B(n6746), .Z(n6707) );
  XOR U1267 ( .A(n6862), .B(n6905), .Z(n6866) );
  XOR U1268 ( .A(n7020), .B(n7063), .Z(n7024) );
  XOR U1269 ( .A(n7735), .B(n7812), .Z(n7739) );
  XOR U1270 ( .A(n7934), .B(n7977), .Z(n7938) );
  XOR U1271 ( .A(n8093), .B(n8136), .Z(n8097) );
  XOR U1272 ( .A(n8251), .B(n8294), .Z(n8255) );
  XOR U1273 ( .A(n8568), .B(n8611), .Z(n8573) );
  XOR U1274 ( .A(n8727), .B(n8771), .Z(n8732) );
  XOR U1275 ( .A(n9091), .B(n9096), .Z(n9017) );
  XOR U1276 ( .A(n9251), .B(n9256), .Z(n9181) );
  XOR U1277 ( .A(n9395), .B(n9400), .Z(n9336) );
  XOR U1278 ( .A(n9510), .B(n9520), .Z(n9468) );
  XOR U1279 ( .A(n10021), .B(n10065), .Z(n10025) );
  XOR U1280 ( .A(n9901), .B(n9945), .Z(n9905) );
  XOR U1281 ( .A(n9757), .B(n9801), .Z(n9761) );
  XOR U1282 ( .A(n9611), .B(n9631), .Z(n9571) );
  XOR U1283 ( .A(n2195), .B(n2239), .Z(n2199) );
  XOR U1284 ( .A(n2367), .B(n2831), .Z(n2371) );
  XNOR U1285 ( .A(n3057), .B(n2974), .Z(n2976) );
  XOR U1286 ( .A(n3131), .B(n3168), .Z(n3135) );
  XOR U1287 ( .A(n4001), .B(n4038), .Z(n4005) );
  XOR U1288 ( .A(n5214), .B(n5252), .Z(n5218) );
  XOR U1289 ( .A(n6434), .B(n6472), .Z(n6438) );
  XOR U1290 ( .A(n7660), .B(n7698), .Z(n7665) );
  XNOR U1291 ( .A(n9466), .B(n9465), .Z(n9421) );
  XOR U1292 ( .A(n313), .B(n367), .Z(n317) );
  XOR U1293 ( .A(n408), .B(n444), .Z(n412) );
  XOR U1294 ( .A(n576), .B(n612), .Z(n580) );
  XOR U1295 ( .A(n745), .B(n782), .Z(n749) );
  XOR U1296 ( .A(n915), .B(n951), .Z(n919) );
  XOR U1297 ( .A(n1084), .B(n1120), .Z(n1088) );
  XOR U1298 ( .A(n1253), .B(n1289), .Z(n1257) );
  XOR U1299 ( .A(n1422), .B(n1464), .Z(n1426) );
  XOR U1300 ( .A(n1598), .B(n1636), .Z(n1602) );
  XOR U1301 ( .A(n1770), .B(n1808), .Z(n1774) );
  XOR U1302 ( .A(n1942), .B(n1980), .Z(n1946) );
  XOR U1303 ( .A(n2114), .B(n2152), .Z(n2118) );
  XOR U1304 ( .A(n3294), .B(n3325), .Z(n3298) );
  XOR U1305 ( .A(n3452), .B(n3483), .Z(n3456) );
  XOR U1306 ( .A(n3605), .B(n3641), .Z(n3614) );
  XOR U1307 ( .A(n3769), .B(n3800), .Z(n3777) );
  XOR U1308 ( .A(n4189), .B(n4220), .Z(n4193) );
  XOR U1309 ( .A(n4349), .B(n4380), .Z(n4353) );
  XOR U1310 ( .A(n4507), .B(n4538), .Z(n4511) );
  XOR U1311 ( .A(n4665), .B(n4696), .Z(n4669) );
  XOR U1312 ( .A(n4818), .B(n4854), .Z(n4827) );
  XOR U1313 ( .A(n4982), .B(n5013), .Z(n4990) );
  XOR U1314 ( .A(n5408), .B(n5439), .Z(n5412) );
  XOR U1315 ( .A(n5568), .B(n5599), .Z(n5572) );
  XOR U1316 ( .A(n5726), .B(n5757), .Z(n5730) );
  XOR U1317 ( .A(n5884), .B(n5915), .Z(n5888) );
  XOR U1318 ( .A(n6037), .B(n6073), .Z(n6046) );
  XOR U1319 ( .A(n6201), .B(n6232), .Z(n6205) );
  XOR U1320 ( .A(n6633), .B(n6638), .Z(n6557) );
  XOR U1321 ( .A(n6793), .B(n6798), .Z(n6723) );
  XOR U1322 ( .A(n6951), .B(n6956), .Z(n6882) );
  XOR U1323 ( .A(n7109), .B(n7114), .Z(n7040) );
  XOR U1324 ( .A(n7262), .B(n7272), .Z(n7198) );
  XOR U1325 ( .A(n7453), .B(n7425), .Z(n7352) );
  XOR U1326 ( .A(n7811), .B(n7783), .Z(n7751) );
  XOR U1327 ( .A(n7976), .B(n7948), .Z(n7874) );
  XOR U1328 ( .A(n8135), .B(n8107), .Z(n8034) );
  XOR U1329 ( .A(n8293), .B(n8265), .Z(n8192) );
  XOR U1330 ( .A(n8451), .B(n8423), .Z(n8350) );
  XOR U1331 ( .A(n8925), .B(n8897), .Z(n8823) );
  XOR U1332 ( .A(n9049), .B(n9021), .Z(n8983) );
  XOR U1333 ( .A(n9213), .B(n9185), .Z(n9111) );
  XOR U1334 ( .A(n9358), .B(n9340), .Z(n9271) );
  XNOR U1335 ( .A(n3147), .B(n3064), .Z(n3066) );
  XNOR U1336 ( .A(n3305), .B(n3223), .Z(n3225) );
  XOR U1337 ( .A(n3932), .B(n3957), .Z(n3936) );
  XOR U1338 ( .A(n5145), .B(n5170), .Z(n5150) );
  XOR U1339 ( .A(n6386), .B(n6363), .Z(n6290) );
  XOR U1340 ( .A(n7532), .B(n7509), .Z(n7436) );
  XOR U1341 ( .A(n8604), .B(n8582), .Z(n8511) );
  XOR U1342 ( .A(n8764), .B(n8741), .Z(n8667) );
  XOR U1343 ( .A(n10204), .B(n10230), .Z(n10208) );
  XOR U1344 ( .A(n10132), .B(n10158), .Z(n10136) );
  XOR U1345 ( .A(n10036), .B(n10062), .Z(n10040) );
  XOR U1346 ( .A(n9916), .B(n9942), .Z(n9920) );
  XOR U1347 ( .A(n9772), .B(n9798), .Z(n9776) );
  XOR U1348 ( .A(n9477), .B(n9628), .Z(n9418) );
  XOR U1349 ( .A(n2888), .B(n2916), .Z(n2892) );
  XNOR U1350 ( .A(n3152), .B(n3069), .Z(n3071) );
  XNOR U1351 ( .A(n3310), .B(n3228), .Z(n3230) );
  XOR U1352 ( .A(n3383), .B(n3402), .Z(n3387) );
  XOR U1353 ( .A(n3541), .B(n3560), .Z(n3545) );
  XOR U1354 ( .A(n3699), .B(n3718), .Z(n3703) );
  XOR U1355 ( .A(n4095), .B(n4116), .Z(n4101) );
  XOR U1356 ( .A(n4279), .B(n4284), .Z(n4209) );
  XOR U1357 ( .A(n4438), .B(n4443), .Z(n4369) );
  XOR U1358 ( .A(n4596), .B(n4601), .Z(n4527) );
  XOR U1359 ( .A(n4754), .B(n4759), .Z(n4685) );
  XOR U1360 ( .A(n4912), .B(n4917), .Z(n4843) );
  XOR U1361 ( .A(n5325), .B(n5309), .Z(n5235) );
  XOR U1362 ( .A(n5438), .B(n5422), .Z(n5341) );
  XOR U1363 ( .A(n5598), .B(n5582), .Z(n5508) );
  XOR U1364 ( .A(n5756), .B(n5740), .Z(n5667) );
  XOR U1365 ( .A(n5914), .B(n5898), .Z(n5825) );
  XOR U1366 ( .A(n6072), .B(n6056), .Z(n5983) );
  XOR U1367 ( .A(n6465), .B(n6449), .Z(n6375) );
  XOR U1368 ( .A(n6577), .B(n6561), .Z(n6535) );
  XOR U1369 ( .A(n6743), .B(n6727), .Z(n6653) );
  XOR U1370 ( .A(n6902), .B(n6886), .Z(n6813) );
  XOR U1371 ( .A(n7060), .B(n7044), .Z(n6971) );
  XOR U1372 ( .A(n7218), .B(n7202), .Z(n7129) );
  XOR U1373 ( .A(n7611), .B(n7595), .Z(n7521) );
  XOR U1374 ( .A(n7771), .B(n7755), .Z(n7681) );
  XOR U1375 ( .A(n7894), .B(n7878), .Z(n7799) );
  XOR U1376 ( .A(n8054), .B(n8038), .Z(n7964) );
  XOR U1377 ( .A(n8212), .B(n8196), .Z(n8123) );
  XOR U1378 ( .A(n8370), .B(n8354), .Z(n8281) );
  XOR U1379 ( .A(n8843), .B(n8827), .Z(n8753) );
  XOR U1380 ( .A(n9003), .B(n8987), .Z(n8913) );
  XOR U1381 ( .A(n9131), .B(n9115), .Z(n9037) );
  XOR U1382 ( .A(n9287), .B(n9275), .Z(n9201) );
  XOR U1383 ( .A(n423), .B(n441), .Z(n432) );
  XOR U1384 ( .A(n591), .B(n609), .Z(n600) );
  XOR U1385 ( .A(n845), .B(n864), .Z(n854) );
  XOR U1386 ( .A(n1014), .B(n1033), .Z(n1023) );
  XOR U1387 ( .A(n1183), .B(n1202), .Z(n1192) );
  XOR U1388 ( .A(n1352), .B(n1371), .Z(n1361) );
  XOR U1389 ( .A(n1527), .B(n1547), .Z(n1536) );
  XOR U1390 ( .A(n1699), .B(n1719), .Z(n1708) );
  XOR U1391 ( .A(n1871), .B(n1891), .Z(n1880) );
  XOR U1392 ( .A(n2043), .B(n2063), .Z(n2052) );
  XOR U1393 ( .A(n2215), .B(n2235), .Z(n2224) );
  XOR U1394 ( .A(n2387), .B(n2827), .Z(n2396) );
  XOR U1395 ( .A(n3857), .B(n3867), .Z(n3793) );
  XOR U1396 ( .A(n5010), .B(n5000), .Z(n4927) );
  XOR U1397 ( .A(n6150), .B(n6140), .Z(n6067) );
  XOR U1398 ( .A(n7296), .B(n7286), .Z(n7213) );
  XOR U1399 ( .A(n768), .B(n775), .Z(n764) );
  XNOR U1400 ( .A(n2913), .B(n2911), .Z(n2901) );
  XNOR U1401 ( .A(n3082), .B(n3080), .Z(n3004) );
  XNOR U1402 ( .A(n3241), .B(n3239), .Z(n3164) );
  XNOR U1403 ( .A(n3399), .B(n3397), .Z(n3322) );
  XNOR U1404 ( .A(n3557), .B(n3555), .Z(n3480) );
  XNOR U1405 ( .A(n3715), .B(n3713), .Z(n3638) );
  XNOR U1406 ( .A(n3947), .B(n3945), .Z(n3875) );
  XNOR U1407 ( .A(n4107), .B(n4105), .Z(n4029) );
  XNOR U1408 ( .A(n4215), .B(n4213), .Z(n4129) );
  XNOR U1409 ( .A(n4375), .B(n4373), .Z(n4297) );
  XNOR U1410 ( .A(n4533), .B(n4531), .Z(n4456) );
  XNOR U1411 ( .A(n4691), .B(n4689), .Z(n4614) );
  XNOR U1412 ( .A(n4849), .B(n4847), .Z(n4772) );
  XNOR U1413 ( .A(n5082), .B(n5080), .Z(n5009) );
  XNOR U1414 ( .A(n5241), .B(n5239), .Z(n5163) );
  XNOR U1415 ( .A(n5347), .B(n5345), .Z(n5323) );
  XNOR U1416 ( .A(n5514), .B(n5512), .Z(n5436) );
  XNOR U1417 ( .A(n5673), .B(n5671), .Z(n5596) );
  XNOR U1418 ( .A(n5831), .B(n5829), .Z(n5754) );
  XNOR U1419 ( .A(n5989), .B(n5987), .Z(n5912) );
  XNOR U1420 ( .A(n6223), .B(n6221), .Z(n6149) );
  XNOR U1421 ( .A(n6381), .B(n6379), .Z(n6303) );
  XNOR U1422 ( .A(n6541), .B(n6539), .Z(n6463) );
  XNOR U1423 ( .A(n6659), .B(n6657), .Z(n6575) );
  XNOR U1424 ( .A(n6819), .B(n6817), .Z(n6741) );
  XNOR U1425 ( .A(n6977), .B(n6975), .Z(n6900) );
  XNOR U1426 ( .A(n7135), .B(n7133), .Z(n7058) );
  XNOR U1427 ( .A(n7370), .B(n7368), .Z(n7295) );
  XNOR U1428 ( .A(n7527), .B(n7525), .Z(n7449) );
  XNOR U1429 ( .A(n7687), .B(n7685), .Z(n7609) );
  XNOR U1430 ( .A(n7805), .B(n7803), .Z(n7769) );
  XNOR U1431 ( .A(n7970), .B(n7968), .Z(n7892) );
  XNOR U1432 ( .A(n8129), .B(n8127), .Z(n8052) );
  XNOR U1433 ( .A(n8287), .B(n8285), .Z(n8210) );
  XNOR U1434 ( .A(n8445), .B(n8443), .Z(n8368) );
  XNOR U1435 ( .A(n8599), .B(n8597), .Z(n8526) );
  XNOR U1436 ( .A(n8759), .B(n8757), .Z(n8681) );
  XNOR U1437 ( .A(n8919), .B(n8917), .Z(n8841) );
  XNOR U1438 ( .A(n9043), .B(n9041), .Z(n9001) );
  XNOR U1439 ( .A(n9207), .B(n9205), .Z(n9129) );
  XNOR U1440 ( .A(n10281), .B(n10282), .Z(n10276) );
  XNOR U1441 ( .A(n10240), .B(n10239), .Z(n10228) );
  XNOR U1442 ( .A(n10180), .B(n10179), .Z(n10156) );
  XNOR U1443 ( .A(n10096), .B(n10095), .Z(n10060) );
  XNOR U1444 ( .A(n9988), .B(n9987), .Z(n9940) );
  XNOR U1445 ( .A(n9856), .B(n9855), .Z(n9796) );
  XNOR U1446 ( .A(n9697), .B(n9696), .Z(n9626) );
  AND U1447 ( .A(n602), .B(n601), .Z(n513) );
  AND U1448 ( .A(n941), .B(n940), .Z(n855) );
  AND U1449 ( .A(n1279), .B(n1278), .Z(n1193) );
  XOR U1450 ( .A(n629), .B(n703), .Z(n634) );
  XOR U1451 ( .A(n799), .B(n873), .Z(n804) );
  XOR U1452 ( .A(n968), .B(n1042), .Z(n973) );
  XOR U1453 ( .A(n1137), .B(n1211), .Z(n1142) );
  XOR U1454 ( .A(n1306), .B(n1380), .Z(n1311) );
  XOR U1455 ( .A(n1481), .B(n1556), .Z(n1486) );
  XOR U1456 ( .A(n1653), .B(n1728), .Z(n1658) );
  XOR U1457 ( .A(n1825), .B(n1900), .Z(n1830) );
  XOR U1458 ( .A(n1997), .B(n2072), .Z(n2002) );
  XOR U1459 ( .A(n2847), .B(n2932), .Z(n2852) );
  XNOR U1460 ( .A(n3191), .B(n3109), .Z(n3110) );
  XOR U1461 ( .A(n3817), .B(n3885), .Z(n3822) );
  XNOR U1462 ( .A(n4245), .B(n4162), .Z(n4164) );
  XNOR U1463 ( .A(n4404), .B(n4322), .Z(n4323) );
  XOR U1464 ( .A(n5030), .B(n5098), .Z(n5035) );
  XNOR U1465 ( .A(n5464), .B(n5381), .Z(n5383) );
  XNOR U1466 ( .A(n5623), .B(n5541), .Z(n5542) );
  XOR U1467 ( .A(n6249), .B(n6317), .Z(n6254) );
  XNOR U1468 ( .A(n6689), .B(n6606), .Z(n6608) );
  XNOR U1469 ( .A(n6848), .B(n6766), .Z(n6767) );
  XOR U1470 ( .A(n7474), .B(n7543), .Z(n7479) );
  XNOR U1471 ( .A(n7920), .B(n7837), .Z(n7839) );
  XNOR U1472 ( .A(n8079), .B(n7997), .Z(n7998) );
  XOR U1473 ( .A(n8946), .B(n9057), .Z(n8951) );
  XNOR U1474 ( .A(n9237), .B(n9154), .Z(n9156) );
  XOR U1475 ( .A(n2175), .B(n2243), .Z(n2179) );
  XOR U1476 ( .A(n3031), .B(n3092), .Z(n3035) );
  XNOR U1477 ( .A(n3274), .B(n3331), .Z(n3269) );
  XOR U1478 ( .A(n3428), .B(n3489), .Z(n3432) );
  XOR U1479 ( .A(n3586), .B(n3647), .Z(n3590) );
  XOR U1480 ( .A(n3744), .B(n3805), .Z(n3748) );
  XNOR U1481 ( .A(n4487), .B(n4544), .Z(n4482) );
  XOR U1482 ( .A(n4641), .B(n4702), .Z(n4645) );
  XOR U1483 ( .A(n4799), .B(n4860), .Z(n4803) );
  XOR U1484 ( .A(n4957), .B(n5018), .Z(n4961) );
  XNOR U1485 ( .A(n5706), .B(n5763), .Z(n5701) );
  XOR U1486 ( .A(n5860), .B(n5921), .Z(n5864) );
  XOR U1487 ( .A(n6018), .B(n6079), .Z(n6022) );
  XOR U1488 ( .A(n6176), .B(n6237), .Z(n6180) );
  XNOR U1489 ( .A(n6931), .B(n6988), .Z(n6926) );
  XOR U1490 ( .A(n7085), .B(n7146), .Z(n7089) );
  XOR U1491 ( .A(n7243), .B(n7304), .Z(n7247) );
  XOR U1492 ( .A(n7401), .B(n7462), .Z(n7405) );
  XOR U1493 ( .A(n8237), .B(n8298), .Z(n8245) );
  XOR U1494 ( .A(n8872), .B(n8934), .Z(n8876) );
  XOR U1495 ( .A(n9817), .B(n9879), .Z(n9821) );
  XOR U1496 ( .A(n9658), .B(n9720), .Z(n9662) );
  XOR U1497 ( .A(n556), .B(n616), .Z(n560) );
  XOR U1498 ( .A(n2352), .B(n2834), .Z(n2356) );
  XOR U1499 ( .A(n2956), .B(n3011), .Z(n2960) );
  XOR U1500 ( .A(n3195), .B(n3250), .Z(n3199) );
  XOR U1501 ( .A(n4065), .B(n4141), .Z(n4069) );
  XOR U1502 ( .A(n4249), .B(n4304), .Z(n4253) );
  XOR U1503 ( .A(n4408), .B(n4463), .Z(n4412) );
  XOR U1504 ( .A(n5279), .B(n5360), .Z(n5283) );
  XOR U1505 ( .A(n5468), .B(n5523), .Z(n5472) );
  XOR U1506 ( .A(n5627), .B(n5682), .Z(n5631) );
  XOR U1507 ( .A(n6499), .B(n6585), .Z(n6503) );
  XOR U1508 ( .A(n6693), .B(n6748), .Z(n6697) );
  XOR U1509 ( .A(n6852), .B(n6907), .Z(n6856) );
  XOR U1510 ( .A(n7725), .B(n7816), .Z(n7729) );
  XOR U1511 ( .A(n7924), .B(n7979), .Z(n7928) );
  XOR U1512 ( .A(n8083), .B(n8138), .Z(n8087) );
  XOR U1513 ( .A(n8400), .B(n8455), .Z(n8404) );
  XOR U1514 ( .A(n8558), .B(n8613), .Z(n8562) );
  XOR U1515 ( .A(n8717), .B(n8773), .Z(n8721) );
  XOR U1516 ( .A(n9081), .B(n9136), .Z(n9085) );
  XOR U1517 ( .A(n9241), .B(n9292), .Z(n9245) );
  XNOR U1518 ( .A(n9454), .B(n9388), .Z(n9390) );
  XNOR U1519 ( .A(n9453), .B(n9482), .Z(n9448) );
  XOR U1520 ( .A(n9557), .B(n9578), .Z(n9561) );
  XOR U1521 ( .A(n730), .B(n785), .Z(n734) );
  XOR U1522 ( .A(n900), .B(n954), .Z(n904) );
  XOR U1523 ( .A(n1069), .B(n1123), .Z(n1073) );
  XOR U1524 ( .A(n1238), .B(n1292), .Z(n1242) );
  XOR U1525 ( .A(n1407), .B(n1467), .Z(n1411) );
  XOR U1526 ( .A(n1583), .B(n1639), .Z(n1587) );
  XOR U1527 ( .A(n1755), .B(n1811), .Z(n1759) );
  XOR U1528 ( .A(n1927), .B(n1983), .Z(n1931) );
  XOR U1529 ( .A(n2099), .B(n2155), .Z(n2103) );
  XOR U1530 ( .A(n3121), .B(n3170), .Z(n3125) );
  XOR U1531 ( .A(n3991), .B(n4040), .Z(n3995) );
  XOR U1532 ( .A(n5204), .B(n5254), .Z(n5208) );
  XOR U1533 ( .A(n6424), .B(n6474), .Z(n6428) );
  XOR U1534 ( .A(n7650), .B(n7700), .Z(n7654) );
  XOR U1535 ( .A(n302), .B(n369), .Z(n307) );
  XOR U1536 ( .A(n2276), .B(n2326), .Z(n2280) );
  XOR U1537 ( .A(n3046), .B(n3089), .Z(n3050) );
  XOR U1538 ( .A(n3284), .B(n3327), .Z(n3288) );
  XOR U1539 ( .A(n3437), .B(n3485), .Z(n3446) );
  XOR U1540 ( .A(n3680), .B(n3723), .Z(n3684) );
  XOR U1541 ( .A(n3838), .B(n3881), .Z(n3842) );
  XOR U1542 ( .A(n4179), .B(n4222), .Z(n4183) );
  XOR U1543 ( .A(n4339), .B(n4382), .Z(n4343) );
  XOR U1544 ( .A(n4497), .B(n4540), .Z(n4501) );
  XOR U1545 ( .A(n4650), .B(n4698), .Z(n4659) );
  XOR U1546 ( .A(n4893), .B(n4936), .Z(n4897) );
  XOR U1547 ( .A(n5051), .B(n5094), .Z(n5055) );
  XOR U1548 ( .A(n5398), .B(n5441), .Z(n5402) );
  XOR U1549 ( .A(n5558), .B(n5601), .Z(n5562) );
  XOR U1550 ( .A(n5716), .B(n5759), .Z(n5720) );
  XOR U1551 ( .A(n5869), .B(n5917), .Z(n5878) );
  XOR U1552 ( .A(n6112), .B(n6155), .Z(n6116) );
  XOR U1553 ( .A(n6270), .B(n6313), .Z(n6274) );
  XOR U1554 ( .A(n6623), .B(n6666), .Z(n6627) );
  XOR U1555 ( .A(n6783), .B(n6826), .Z(n6787) );
  XOR U1556 ( .A(n6941), .B(n6984), .Z(n6945) );
  XOR U1557 ( .A(n7094), .B(n7142), .Z(n7103) );
  XOR U1558 ( .A(n7337), .B(n7380), .Z(n7341) );
  XOR U1559 ( .A(n7495), .B(n7539), .Z(n7499) );
  XOR U1560 ( .A(n7854), .B(n7897), .Z(n7858) );
  XOR U1561 ( .A(n8014), .B(n8057), .Z(n8018) );
  XOR U1562 ( .A(n8172), .B(n8215), .Z(n8176) );
  XOR U1563 ( .A(n8325), .B(n8373), .Z(n8334) );
  XOR U1564 ( .A(n8967), .B(n9012), .Z(n8973) );
  XOR U1565 ( .A(n9171), .B(n9176), .Z(n9101) );
  XOR U1566 ( .A(n9326), .B(n9331), .Z(n9261) );
  XOR U1567 ( .A(n10072), .B(n10116), .Z(n10076) );
  XOR U1568 ( .A(n9964), .B(n10008), .Z(n9968) );
  XOR U1569 ( .A(n9832), .B(n9876), .Z(n9836) );
  XOR U1570 ( .A(n9673), .B(n9717), .Z(n9677) );
  XOR U1571 ( .A(n483), .B(n526), .Z(n487) );
  XOR U1572 ( .A(n655), .B(n698), .Z(n659) );
  XOR U1573 ( .A(n2873), .B(n2922), .Z(n2877) );
  XNOR U1574 ( .A(n3137), .B(n3054), .Z(n3056) );
  XOR U1575 ( .A(n3210), .B(n3247), .Z(n3214) );
  XNOR U1576 ( .A(n3610), .B(n3643), .Z(n3605) );
  XNOR U1577 ( .A(n4823), .B(n4856), .Z(n4818) );
  XNOR U1578 ( .A(n6042), .B(n6075), .Z(n6037) );
  XNOR U1579 ( .A(n7267), .B(n7300), .Z(n7262) );
  XOR U1580 ( .A(n8606), .B(n8572), .Z(n8499) );
  XOR U1581 ( .A(n8766), .B(n8731), .Z(n8657) );
  XOR U1582 ( .A(n8926), .B(n8891), .Z(n8817) );
  XOR U1583 ( .A(n9422), .B(n9404), .Z(n9341) );
  XOR U1584 ( .A(n9479), .B(n9467), .Z(n9410) );
  XOR U1585 ( .A(n9530), .B(n9524), .Z(n9473) );
  XOR U1586 ( .A(n830), .B(n867), .Z(n834) );
  XOR U1587 ( .A(n999), .B(n1036), .Z(n1003) );
  XOR U1588 ( .A(n1168), .B(n1205), .Z(n1172) );
  XOR U1589 ( .A(n1337), .B(n1374), .Z(n1341) );
  XOR U1590 ( .A(n1512), .B(n1550), .Z(n1516) );
  XOR U1591 ( .A(n1684), .B(n1722), .Z(n1688) );
  XOR U1592 ( .A(n1856), .B(n1894), .Z(n1860) );
  XOR U1593 ( .A(n2028), .B(n2066), .Z(n2032) );
  XOR U1594 ( .A(n2200), .B(n2238), .Z(n2204) );
  XOR U1595 ( .A(n3373), .B(n3404), .Z(n3377) );
  XOR U1596 ( .A(n3531), .B(n3562), .Z(n3535) );
  XOR U1597 ( .A(n4085), .B(n4133), .Z(n4089) );
  XOR U1598 ( .A(n4269), .B(n4300), .Z(n4273) );
  XOR U1599 ( .A(n4428), .B(n4459), .Z(n4432) );
  XOR U1600 ( .A(n4586), .B(n4617), .Z(n4590) );
  XOR U1601 ( .A(n4744), .B(n4775), .Z(n4748) );
  XOR U1602 ( .A(n5299), .B(n5352), .Z(n5303) );
  XOR U1603 ( .A(n5488), .B(n5519), .Z(n5492) );
  XOR U1604 ( .A(n5647), .B(n5678), .Z(n5651) );
  XOR U1605 ( .A(n5805), .B(n5836), .Z(n5809) );
  XOR U1606 ( .A(n5963), .B(n5994), .Z(n5967) );
  XOR U1607 ( .A(n6519), .B(n6552), .Z(n6525) );
  XOR U1608 ( .A(n6713), .B(n6718), .Z(n6643) );
  XOR U1609 ( .A(n6872), .B(n6877), .Z(n6803) );
  XOR U1610 ( .A(n7030), .B(n7035), .Z(n6961) );
  XOR U1611 ( .A(n7188), .B(n7193), .Z(n7119) );
  XOR U1612 ( .A(n7773), .B(n7745), .Z(n7671) );
  XOR U1613 ( .A(n7896), .B(n7868), .Z(n7789) );
  XOR U1614 ( .A(n8056), .B(n8028), .Z(n7954) );
  XOR U1615 ( .A(n8214), .B(n8186), .Z(n8113) );
  XOR U1616 ( .A(n8372), .B(n8344), .Z(n8271) );
  XOR U1617 ( .A(n9005), .B(n8977), .Z(n8903) );
  XOR U1618 ( .A(n9133), .B(n9105), .Z(n9027) );
  XOR U1619 ( .A(n9289), .B(n9265), .Z(n9191) );
  XOR U1620 ( .A(n318), .B(n366), .Z(n322) );
  XOR U1621 ( .A(n2377), .B(n2829), .Z(n2381) );
  XNOR U1622 ( .A(n3067), .B(n2984), .Z(n2986) );
  XNOR U1623 ( .A(n3226), .B(n3144), .Z(n3146) );
  XOR U1624 ( .A(n3299), .B(n3324), .Z(n3303) );
  XOR U1625 ( .A(n3853), .B(n3878), .Z(n3861) );
  XOR U1626 ( .A(n4011), .B(n4036), .Z(n4015) );
  XOR U1627 ( .A(n5066), .B(n5091), .Z(n5070) );
  XOR U1628 ( .A(n5224), .B(n5250), .Z(n5229) );
  XOR U1629 ( .A(n6306), .B(n6284), .Z(n6211) );
  XOR U1630 ( .A(n6466), .B(n6443), .Z(n6369) );
  XOR U1631 ( .A(n7452), .B(n7430), .Z(n7358) );
  XOR U1632 ( .A(n7612), .B(n7589), .Z(n7515) );
  XOR U1633 ( .A(n10171), .B(n10197), .Z(n10175) );
  XOR U1634 ( .A(n10087), .B(n10113), .Z(n10091) );
  XOR U1635 ( .A(n9979), .B(n10005), .Z(n9983) );
  XOR U1636 ( .A(n9847), .B(n9873), .Z(n9851) );
  XOR U1637 ( .A(n9688), .B(n9714), .Z(n9692) );
  XOR U1638 ( .A(n755), .B(n780), .Z(n759) );
  XNOR U1639 ( .A(n3072), .B(n2989), .Z(n2991) );
  XNOR U1640 ( .A(n3231), .B(n3149), .Z(n3151) );
  XNOR U1641 ( .A(n3389), .B(n3307), .Z(n3309) );
  XOR U1642 ( .A(n3462), .B(n3481), .Z(n3466) );
  XOR U1643 ( .A(n3620), .B(n3639), .Z(n3624) );
  XOR U1644 ( .A(n3773), .B(n3797), .Z(n3782) );
  XOR U1645 ( .A(n4199), .B(n4204), .Z(n4121) );
  XOR U1646 ( .A(n4359), .B(n4364), .Z(n4289) );
  XOR U1647 ( .A(n4517), .B(n4522), .Z(n4448) );
  XOR U1648 ( .A(n4675), .B(n4680), .Z(n4606) );
  XOR U1649 ( .A(n4833), .B(n4838), .Z(n4764) );
  XOR U1650 ( .A(n4986), .B(n4996), .Z(n4922) );
  XOR U1651 ( .A(n5351), .B(n5335), .Z(n5315) );
  XOR U1652 ( .A(n5518), .B(n5502), .Z(n5428) );
  XOR U1653 ( .A(n5677), .B(n5661), .Z(n5588) );
  XOR U1654 ( .A(n5835), .B(n5819), .Z(n5746) );
  XOR U1655 ( .A(n5993), .B(n5977), .Z(n5904) );
  XOR U1656 ( .A(n6151), .B(n6135), .Z(n6062) );
  XOR U1657 ( .A(n6545), .B(n6529), .Z(n6455) );
  XOR U1658 ( .A(n6663), .B(n6647), .Z(n6567) );
  XOR U1659 ( .A(n6823), .B(n6807), .Z(n6733) );
  XOR U1660 ( .A(n6981), .B(n6965), .Z(n6892) );
  XOR U1661 ( .A(n7139), .B(n7123), .Z(n7050) );
  XOR U1662 ( .A(n7297), .B(n7281), .Z(n7208) );
  XOR U1663 ( .A(n7691), .B(n7675), .Z(n7601) );
  XOR U1664 ( .A(n7809), .B(n7793), .Z(n7761) );
  XOR U1665 ( .A(n7974), .B(n7958), .Z(n7884) );
  XOR U1666 ( .A(n8133), .B(n8117), .Z(n8044) );
  XOR U1667 ( .A(n8291), .B(n8275), .Z(n8202) );
  XOR U1668 ( .A(n8449), .B(n8433), .Z(n8360) );
  XOR U1669 ( .A(n8603), .B(n8587), .Z(n8518) );
  XOR U1670 ( .A(n8763), .B(n8747), .Z(n8673) );
  XOR U1671 ( .A(n8923), .B(n8907), .Z(n8833) );
  XOR U1672 ( .A(n9047), .B(n9031), .Z(n8993) );
  XOR U1673 ( .A(n9211), .B(n9195), .Z(n9121) );
  XOR U1674 ( .A(n9356), .B(n9350), .Z(n9281) );
  XOR U1675 ( .A(n343), .B(n361), .Z(n352) );
  XOR U1676 ( .A(n503), .B(n522), .Z(n512) );
  XOR U1677 ( .A(n675), .B(n694), .Z(n683) );
  XOR U1678 ( .A(n930), .B(n948), .Z(n939) );
  XOR U1679 ( .A(n1099), .B(n1117), .Z(n1108) );
  XOR U1680 ( .A(n1268), .B(n1286), .Z(n1277) );
  XOR U1681 ( .A(n1437), .B(n1461), .Z(n1446) );
  XOR U1682 ( .A(n1613), .B(n1633), .Z(n1622) );
  XOR U1683 ( .A(n1785), .B(n1805), .Z(n1794) );
  XOR U1684 ( .A(n1957), .B(n1977), .Z(n1966) );
  XOR U1685 ( .A(n2129), .B(n2149), .Z(n2138) );
  XOR U1686 ( .A(n2301), .B(n2321), .Z(n2310) );
  XNOR U1687 ( .A(n2899), .B(n2897), .Z(n2826) );
  XNOR U1688 ( .A(n3002), .B(n3000), .Z(n2915) );
  XNOR U1689 ( .A(n3162), .B(n3160), .Z(n3084) );
  XNOR U1690 ( .A(n3320), .B(n3318), .Z(n3243) );
  XNOR U1691 ( .A(n3478), .B(n3476), .Z(n3401) );
  XNOR U1692 ( .A(n3636), .B(n3634), .Z(n3559) );
  XNOR U1693 ( .A(n3794), .B(n3792), .Z(n3717) );
  XNOR U1694 ( .A(n4027), .B(n4025), .Z(n3950) );
  XNOR U1695 ( .A(n4127), .B(n4125), .Z(n4109) );
  XNOR U1696 ( .A(n4295), .B(n4293), .Z(n4217) );
  XNOR U1697 ( .A(n4454), .B(n4452), .Z(n4377) );
  XNOR U1698 ( .A(n4612), .B(n4610), .Z(n4535) );
  XNOR U1699 ( .A(n4770), .B(n4768), .Z(n4693) );
  XNOR U1700 ( .A(n4928), .B(n4926), .Z(n4851) );
  XNOR U1701 ( .A(n5161), .B(n5159), .Z(n5085) );
  XNOR U1702 ( .A(n5321), .B(n5319), .Z(n5243) );
  XNOR U1703 ( .A(n5434), .B(n5432), .Z(n5349) );
  XNOR U1704 ( .A(n5594), .B(n5592), .Z(n5516) );
  XNOR U1705 ( .A(n5752), .B(n5750), .Z(n5675) );
  XNOR U1706 ( .A(n5910), .B(n5908), .Z(n5833) );
  XNOR U1707 ( .A(n6068), .B(n6066), .Z(n5991) );
  XNOR U1708 ( .A(n6301), .B(n6299), .Z(n6226) );
  XNOR U1709 ( .A(n6461), .B(n6459), .Z(n6383) );
  XNOR U1710 ( .A(n6573), .B(n6571), .Z(n6543) );
  XNOR U1711 ( .A(n6739), .B(n6737), .Z(n6661) );
  XNOR U1712 ( .A(n6898), .B(n6896), .Z(n6821) );
  XNOR U1713 ( .A(n7056), .B(n7054), .Z(n6979) );
  XNOR U1714 ( .A(n7214), .B(n7212), .Z(n7137) );
  XNOR U1715 ( .A(n7447), .B(n7445), .Z(n7373) );
  XNOR U1716 ( .A(n7607), .B(n7605), .Z(n7529) );
  XNOR U1717 ( .A(n7767), .B(n7765), .Z(n7689) );
  XNOR U1718 ( .A(n7890), .B(n7888), .Z(n7807) );
  XNOR U1719 ( .A(n8050), .B(n8048), .Z(n7972) );
  XNOR U1720 ( .A(n8208), .B(n8206), .Z(n8131) );
  XNOR U1721 ( .A(n8366), .B(n8364), .Z(n8289) );
  XNOR U1722 ( .A(n8679), .B(n8677), .Z(n8601) );
  XNOR U1723 ( .A(n8839), .B(n8837), .Z(n8761) );
  XNOR U1724 ( .A(n8999), .B(n8997), .Z(n8921) );
  XNOR U1725 ( .A(n9127), .B(n9125), .Z(n9045) );
  XNOR U1726 ( .A(n10261), .B(n10260), .Z(n10255) );
  XNOR U1727 ( .A(n10213), .B(n10212), .Z(n10195) );
  XNOR U1728 ( .A(n10141), .B(n10140), .Z(n10111) );
  XNOR U1729 ( .A(n10045), .B(n10044), .Z(n10003) );
  XNOR U1730 ( .A(n9925), .B(n9924), .Z(n9871) );
  XNOR U1731 ( .A(n9781), .B(n9780), .Z(n9712) );
  XNOR U1732 ( .A(n9285), .B(n9284), .Z(n9209) );
  XNOR U1733 ( .A(n764), .B(n763), .Z(n693) );
  XNOR U1734 ( .A(n3875), .B(n3874), .Z(n2470) );
  XNOR U1735 ( .A(n5009), .B(n5008), .Z(n2545) );
  XNOR U1736 ( .A(n6149), .B(n6148), .Z(n2620) );
  XNOR U1737 ( .A(n7295), .B(n7294), .Z(n2695) );
  XNOR U1738 ( .A(n8447), .B(n8446), .Z(n2770) );
  XOR U1739 ( .A(n10276), .B(n10283), .Z(n10270) );
  NANDN U1740 ( .A(n354), .B(n353), .Z(n244) );
  AND U1741 ( .A(n686), .B(n685), .Z(n601) );
  AND U1742 ( .A(n1025), .B(n1024), .Z(n940) );
  AND U1743 ( .A(n1363), .B(n1362), .Z(n1278) );
  XNOR U1744 ( .A(n1), .B(n2), .Z(swire[99]) );
  XNOR U1745 ( .A(n3), .B(n4), .Z(swire[98]) );
  XNOR U1746 ( .A(n5), .B(n6), .Z(swire[97]) );
  XNOR U1747 ( .A(n7), .B(n8), .Z(swire[96]) );
  XNOR U1748 ( .A(n9), .B(n10), .Z(swire[95]) );
  XNOR U1749 ( .A(n11), .B(n12), .Z(swire[94]) );
  XNOR U1750 ( .A(n13), .B(n14), .Z(swire[93]) );
  XNOR U1751 ( .A(n15), .B(n16), .Z(swire[92]) );
  XNOR U1752 ( .A(n17), .B(n18), .Z(swire[91]) );
  XNOR U1753 ( .A(n19), .B(n20), .Z(swire[90]) );
  XNOR U1754 ( .A(n21), .B(n22), .Z(swire[89]) );
  XNOR U1755 ( .A(n23), .B(n24), .Z(swire[88]) );
  XNOR U1756 ( .A(n25), .B(n26), .Z(swire[87]) );
  XNOR U1757 ( .A(n27), .B(n28), .Z(swire[86]) );
  XNOR U1758 ( .A(n29), .B(n30), .Z(swire[85]) );
  XNOR U1759 ( .A(n31), .B(n32), .Z(swire[84]) );
  XNOR U1760 ( .A(n33), .B(n34), .Z(swire[83]) );
  XNOR U1761 ( .A(n35), .B(n36), .Z(swire[82]) );
  XNOR U1762 ( .A(n37), .B(n38), .Z(swire[81]) );
  XNOR U1763 ( .A(n39), .B(n40), .Z(swire[80]) );
  XNOR U1764 ( .A(n41), .B(n42), .Z(swire[79]) );
  XNOR U1765 ( .A(n43), .B(n44), .Z(swire[78]) );
  XNOR U1766 ( .A(n45), .B(n46), .Z(swire[77]) );
  XNOR U1767 ( .A(n47), .B(n48), .Z(swire[76]) );
  XNOR U1768 ( .A(n49), .B(n50), .Z(swire[75]) );
  XNOR U1769 ( .A(n51), .B(n52), .Z(swire[74]) );
  XNOR U1770 ( .A(n53), .B(n54), .Z(swire[73]) );
  XNOR U1771 ( .A(n55), .B(n56), .Z(swire[72]) );
  XNOR U1772 ( .A(n57), .B(n58), .Z(swire[71]) );
  XNOR U1773 ( .A(n59), .B(n60), .Z(swire[70]) );
  XNOR U1774 ( .A(n61), .B(n62), .Z(swire[69]) );
  XNOR U1775 ( .A(n63), .B(n64), .Z(swire[68]) );
  XNOR U1776 ( .A(n65), .B(n66), .Z(swire[67]) );
  XNOR U1777 ( .A(n67), .B(n68), .Z(swire[66]) );
  XNOR U1778 ( .A(n69), .B(n70), .Z(swire[65]) );
  XNOR U1779 ( .A(n71), .B(n72), .Z(swire[64]) );
  XNOR U1780 ( .A(n73), .B(n74), .Z(swire[63]) );
  XNOR U1781 ( .A(n75), .B(n76), .Z(swire[62]) );
  XNOR U1782 ( .A(n77), .B(n78), .Z(swire[61]) );
  XNOR U1783 ( .A(n79), .B(n80), .Z(swire[60]) );
  XNOR U1784 ( .A(n81), .B(n82), .Z(swire[59]) );
  XNOR U1785 ( .A(n83), .B(n84), .Z(swire[58]) );
  XNOR U1786 ( .A(n85), .B(n86), .Z(swire[57]) );
  XNOR U1787 ( .A(n87), .B(n88), .Z(swire[56]) );
  XNOR U1788 ( .A(n89), .B(n90), .Z(swire[55]) );
  XNOR U1789 ( .A(n91), .B(n92), .Z(swire[54]) );
  XNOR U1790 ( .A(n93), .B(n94), .Z(swire[53]) );
  XNOR U1791 ( .A(n95), .B(n96), .Z(swire[52]) );
  XNOR U1792 ( .A(n97), .B(n98), .Z(swire[51]) );
  XNOR U1793 ( .A(n99), .B(n100), .Z(swire[50]) );
  XNOR U1794 ( .A(n101), .B(n102), .Z(swire[49]) );
  XNOR U1795 ( .A(n103), .B(n104), .Z(swire[48]) );
  XNOR U1796 ( .A(n105), .B(n106), .Z(swire[47]) );
  XNOR U1797 ( .A(n107), .B(n108), .Z(swire[46]) );
  XNOR U1798 ( .A(n109), .B(n110), .Z(swire[45]) );
  XNOR U1799 ( .A(n111), .B(n112), .Z(swire[44]) );
  XNOR U1800 ( .A(n113), .B(n114), .Z(swire[43]) );
  XNOR U1801 ( .A(n115), .B(n116), .Z(swire[42]) );
  XNOR U1802 ( .A(n117), .B(n118), .Z(swire[41]) );
  XNOR U1803 ( .A(n119), .B(n120), .Z(swire[40]) );
  XNOR U1804 ( .A(n121), .B(n122), .Z(swire[39]) );
  XNOR U1805 ( .A(n123), .B(n124), .Z(swire[38]) );
  XNOR U1806 ( .A(n125), .B(n126), .Z(swire[37]) );
  XNOR U1807 ( .A(n127), .B(n128), .Z(swire[36]) );
  XNOR U1808 ( .A(n129), .B(n130), .Z(swire[35]) );
  XNOR U1809 ( .A(n131), .B(n132), .Z(swire[34]) );
  XNOR U1810 ( .A(n133), .B(n134), .Z(swire[33]) );
  XNOR U1811 ( .A(n135), .B(n136), .Z(swire[32]) );
  XNOR U1812 ( .A(n137), .B(n138), .Z(swire[31]) );
  XNOR U1813 ( .A(n139), .B(n140), .Z(swire[30]) );
  XNOR U1814 ( .A(n141), .B(n142), .Z(swire[29]) );
  XNOR U1815 ( .A(n143), .B(n144), .Z(swire[28]) );
  XNOR U1816 ( .A(n145), .B(n146), .Z(swire[27]) );
  XNOR U1817 ( .A(n147), .B(n148), .Z(swire[26]) );
  XNOR U1818 ( .A(n149), .B(n150), .Z(swire[25]) );
  XNOR U1819 ( .A(n151), .B(n152), .Z(swire[24]) );
  XNOR U1820 ( .A(n153), .B(n154), .Z(swire[23]) );
  XNOR U1821 ( .A(n155), .B(n156), .Z(swire[22]) );
  XNOR U1822 ( .A(n157), .B(n158), .Z(swire[21]) );
  XNOR U1823 ( .A(n159), .B(n160), .Z(swire[20]) );
  XNOR U1824 ( .A(n161), .B(n162), .Z(swire[19]) );
  XNOR U1825 ( .A(n163), .B(n164), .Z(swire[18]) );
  XNOR U1826 ( .A(n165), .B(n166), .Z(swire[17]) );
  XNOR U1827 ( .A(n167), .B(n168), .Z(swire[16]) );
  XOR U1828 ( .A(n169), .B(n170), .Z(swire[127]) );
  XOR U1829 ( .A(n171), .B(n172), .Z(n170) );
  AND U1830 ( .A(b[1]), .B(a[126]), .Z(n172) );
  AND U1831 ( .A(b[2]), .B(a[125]), .Z(n171) );
  XOR U1832 ( .A(n173), .B(n174), .Z(n169) );
  XOR U1833 ( .A(n175), .B(n176), .Z(n174) );
  XOR U1834 ( .A(n177), .B(n178), .Z(n176) );
  ANDN U1835 ( .B(a[127]), .A(n179), .Z(n178) );
  AND U1836 ( .A(b[3]), .B(a[124]), .Z(n177) );
  XOR U1837 ( .A(n180), .B(n181), .Z(n175) );
  XOR U1838 ( .A(n182), .B(n183), .Z(n181) );
  XOR U1839 ( .A(n184), .B(n185), .Z(n183) );
  AND U1840 ( .A(b[4]), .B(a[123]), .Z(n185) );
  AND U1841 ( .A(b[9]), .B(a[118]), .Z(n184) );
  XOR U1842 ( .A(n186), .B(n187), .Z(n182) );
  AND U1843 ( .A(b[10]), .B(a[117]), .Z(n187) );
  AND U1844 ( .A(b[11]), .B(a[116]), .Z(n186) );
  XOR U1845 ( .A(n188), .B(n189), .Z(n180) );
  XOR U1846 ( .A(n190), .B(n191), .Z(n189) );
  AND U1847 ( .A(b[12]), .B(a[115]), .Z(n191) );
  AND U1848 ( .A(b[13]), .B(a[114]), .Z(n190) );
  XOR U1849 ( .A(n192), .B(n193), .Z(n188) );
  AND U1850 ( .A(b[14]), .B(a[113]), .Z(n193) );
  AND U1851 ( .A(b[15]), .B(a[112]), .Z(n192) );
  XOR U1852 ( .A(n194), .B(n195), .Z(n173) );
  XOR U1853 ( .A(n196), .B(n197), .Z(n195) );
  AND U1854 ( .A(b[5]), .B(a[122]), .Z(n197) );
  AND U1855 ( .A(b[6]), .B(a[121]), .Z(n196) );
  XOR U1856 ( .A(n198), .B(n199), .Z(n194) );
  AND U1857 ( .A(b[7]), .B(a[120]), .Z(n199) );
  AND U1858 ( .A(b[8]), .B(a[119]), .Z(n198) );
  XOR U1859 ( .A(n200), .B(n201), .Z(swire[126]) );
  XOR U1860 ( .A(n202), .B(n203), .Z(n201) );
  XOR U1861 ( .A(n204), .B(n205), .Z(n203) );
  XOR U1862 ( .A(n206), .B(n207), .Z(n205) );
  XOR U1863 ( .A(n208), .B(n209), .Z(n207) );
  XOR U1864 ( .A(n210), .B(n211), .Z(n209) );
  AND U1865 ( .A(b[3]), .B(a[123]), .Z(n210) );
  XOR U1866 ( .A(n212), .B(n213), .Z(n208) );
  XOR U1867 ( .A(n214), .B(n215), .Z(n213) );
  XOR U1868 ( .A(n216), .B(n217), .Z(n215) );
  XOR U1869 ( .A(n218), .B(n216), .Z(n217) );
  AND U1870 ( .A(b[9]), .B(a[117]), .Z(n218) );
  XOR U1871 ( .A(n219), .B(n220), .Z(n216) );
  ANDN U1872 ( .B(n221), .A(n222), .Z(n219) );
  XOR U1873 ( .A(n223), .B(n224), .Z(n214) );
  AND U1874 ( .A(b[10]), .B(a[116]), .Z(n224) );
  AND U1875 ( .A(b[11]), .B(a[115]), .Z(n223) );
  XOR U1876 ( .A(n225), .B(n226), .Z(n212) );
  XOR U1877 ( .A(n227), .B(n228), .Z(n226) );
  AND U1878 ( .A(b[12]), .B(a[114]), .Z(n228) );
  AND U1879 ( .A(b[13]), .B(a[113]), .Z(n227) );
  XOR U1880 ( .A(n229), .B(n230), .Z(n225) );
  AND U1881 ( .A(b[14]), .B(a[112]), .Z(n230) );
  AND U1882 ( .A(b[15]), .B(a[111]), .Z(n229) );
  XOR U1883 ( .A(n231), .B(n211), .Z(n206) );
  XNOR U1884 ( .A(n232), .B(n233), .Z(n211) );
  ANDN U1885 ( .B(n234), .A(n235), .Z(n232) );
  AND U1886 ( .A(b[4]), .B(a[122]), .Z(n231) );
  XOR U1887 ( .A(n236), .B(n237), .Z(n204) );
  XOR U1888 ( .A(n238), .B(n239), .Z(n237) );
  AND U1889 ( .A(b[5]), .B(a[121]), .Z(n239) );
  AND U1890 ( .A(b[6]), .B(a[120]), .Z(n238) );
  XOR U1891 ( .A(n240), .B(n241), .Z(n236) );
  AND U1892 ( .A(b[7]), .B(a[119]), .Z(n241) );
  AND U1893 ( .A(b[8]), .B(a[118]), .Z(n240) );
  ANDN U1894 ( .B(a[126]), .A(n179), .Z(n202) );
  XOR U1895 ( .A(n242), .B(n243), .Z(n200) );
  AND U1896 ( .A(b[1]), .B(a[125]), .Z(n243) );
  AND U1897 ( .A(b[2]), .B(a[124]), .Z(n242) );
  XNOR U1898 ( .A(n244), .B(n245), .Z(swire[125]) );
  XOR U1899 ( .A(n246), .B(n247), .Z(n245) );
  XNOR U1900 ( .A(n248), .B(n244), .Z(n247) );
  ANDN U1901 ( .B(a[125]), .A(n179), .Z(n248) );
  XOR U1902 ( .A(n249), .B(n250), .Z(n246) );
  XNOR U1903 ( .A(n251), .B(n252), .Z(n250) );
  AND U1904 ( .A(b[1]), .B(a[124]), .Z(n252) );
  XNOR U1905 ( .A(n235), .B(n253), .Z(n249) );
  XNOR U1906 ( .A(n251), .B(n234), .Z(n253) );
  XNOR U1907 ( .A(n254), .B(n233), .Z(n234) );
  AND U1908 ( .A(b[2]), .B(a[123]), .Z(n254) );
  OR U1909 ( .A(n255), .B(n256), .Z(n251) );
  XOR U1910 ( .A(n257), .B(n258), .Z(n235) );
  XNOR U1911 ( .A(n233), .B(n259), .Z(n258) );
  XOR U1912 ( .A(n260), .B(n261), .Z(n259) );
  XOR U1913 ( .A(n262), .B(n263), .Z(n261) );
  XOR U1914 ( .A(n264), .B(n265), .Z(n263) );
  XOR U1915 ( .A(n266), .B(n267), .Z(n265) );
  XOR U1916 ( .A(n268), .B(n269), .Z(n267) );
  XOR U1917 ( .A(n270), .B(n271), .Z(n269) );
  XOR U1918 ( .A(n272), .B(n273), .Z(n271) );
  XOR U1919 ( .A(n274), .B(n275), .Z(n273) );
  XOR U1920 ( .A(n221), .B(n276), .Z(n275) );
  XOR U1921 ( .A(n277), .B(n222), .Z(n276) );
  XOR U1922 ( .A(n278), .B(n279), .Z(n222) );
  XOR U1923 ( .A(n220), .B(n280), .Z(n279) );
  XOR U1924 ( .A(n281), .B(n282), .Z(n280) );
  XOR U1925 ( .A(n283), .B(n284), .Z(n282) );
  XOR U1926 ( .A(n285), .B(n286), .Z(n284) );
  XOR U1927 ( .A(n287), .B(n288), .Z(n286) );
  XOR U1928 ( .A(n289), .B(n290), .Z(n288) );
  XOR U1929 ( .A(n291), .B(n292), .Z(n290) );
  XOR U1930 ( .A(n293), .B(n294), .Z(n292) );
  XNOR U1931 ( .A(n295), .B(n296), .Z(n294) );
  AND U1932 ( .A(b[13]), .B(a[112]), .Z(n295) );
  XOR U1933 ( .A(n297), .B(n298), .Z(n293) );
  AND U1934 ( .A(b[14]), .B(a[111]), .Z(n298) );
  AND U1935 ( .A(b[15]), .B(a[110]), .Z(n297) );
  XOR U1936 ( .A(n299), .B(n296), .Z(n289) );
  XOR U1937 ( .A(n300), .B(n301), .Z(n296) );
  NOR U1938 ( .A(n302), .B(n303), .Z(n300) );
  AND U1939 ( .A(b[12]), .B(a[113]), .Z(n299) );
  XOR U1940 ( .A(n304), .B(n291), .Z(n285) );
  XOR U1941 ( .A(n305), .B(n306), .Z(n291) );
  ANDN U1942 ( .B(n307), .A(n308), .Z(n305) );
  AND U1943 ( .A(b[11]), .B(a[114]), .Z(n304) );
  XOR U1944 ( .A(n309), .B(n287), .Z(n281) );
  XOR U1945 ( .A(n310), .B(n311), .Z(n287) );
  ANDN U1946 ( .B(n312), .A(n313), .Z(n310) );
  AND U1947 ( .A(b[10]), .B(a[115]), .Z(n309) );
  XOR U1948 ( .A(n314), .B(n283), .Z(n278) );
  XOR U1949 ( .A(n315), .B(n316), .Z(n283) );
  ANDN U1950 ( .B(n317), .A(n318), .Z(n315) );
  AND U1951 ( .A(b[9]), .B(a[116]), .Z(n314) );
  XOR U1952 ( .A(n319), .B(n220), .Z(n221) );
  XOR U1953 ( .A(n320), .B(n321), .Z(n220) );
  ANDN U1954 ( .B(n322), .A(n323), .Z(n320) );
  AND U1955 ( .A(b[8]), .B(a[117]), .Z(n319) );
  XOR U1956 ( .A(n324), .B(n277), .Z(n272) );
  XOR U1957 ( .A(n325), .B(n326), .Z(n277) );
  ANDN U1958 ( .B(n327), .A(n328), .Z(n325) );
  AND U1959 ( .A(b[7]), .B(a[118]), .Z(n324) );
  XOR U1960 ( .A(n329), .B(n274), .Z(n268) );
  XOR U1961 ( .A(n330), .B(n331), .Z(n274) );
  ANDN U1962 ( .B(n332), .A(n333), .Z(n330) );
  AND U1963 ( .A(b[6]), .B(a[119]), .Z(n329) );
  XOR U1964 ( .A(n334), .B(n270), .Z(n264) );
  XOR U1965 ( .A(n335), .B(n336), .Z(n270) );
  ANDN U1966 ( .B(n337), .A(n338), .Z(n335) );
  AND U1967 ( .A(b[5]), .B(a[120]), .Z(n334) );
  XOR U1968 ( .A(n339), .B(n266), .Z(n260) );
  XOR U1969 ( .A(n340), .B(n341), .Z(n266) );
  ANDN U1970 ( .B(n342), .A(n343), .Z(n340) );
  AND U1971 ( .A(b[4]), .B(a[121]), .Z(n339) );
  XNOR U1972 ( .A(n344), .B(n345), .Z(n233) );
  NANDN U1973 ( .A(n346), .B(n347), .Z(n345) );
  XOR U1974 ( .A(n348), .B(n262), .Z(n257) );
  XNOR U1975 ( .A(n349), .B(n350), .Z(n262) );
  AND U1976 ( .A(n351), .B(n352), .Z(n349) );
  AND U1977 ( .A(b[3]), .B(a[122]), .Z(n348) );
  XOR U1978 ( .A(n353), .B(n354), .Z(swire[124]) );
  XOR U1979 ( .A(n256), .B(n355), .Z(n354) );
  XOR U1980 ( .A(n255), .B(n353), .Z(n355) );
  NANDN U1981 ( .A(n179), .B(a[124]), .Z(n255) );
  XOR U1982 ( .A(n346), .B(n347), .Z(n256) );
  XOR U1983 ( .A(n344), .B(n356), .Z(n347) );
  NAND U1984 ( .A(b[1]), .B(a[123]), .Z(n356) );
  XOR U1985 ( .A(n352), .B(n357), .Z(n346) );
  XOR U1986 ( .A(n344), .B(n351), .Z(n357) );
  XNOR U1987 ( .A(n358), .B(n350), .Z(n351) );
  AND U1988 ( .A(b[2]), .B(a[122]), .Z(n358) );
  NANDN U1989 ( .A(n359), .B(n360), .Z(n344) );
  XOR U1990 ( .A(n350), .B(n342), .Z(n361) );
  XNOR U1991 ( .A(n341), .B(n337), .Z(n362) );
  XNOR U1992 ( .A(n336), .B(n332), .Z(n363) );
  XNOR U1993 ( .A(n331), .B(n327), .Z(n364) );
  XNOR U1994 ( .A(n326), .B(n322), .Z(n365) );
  XNOR U1995 ( .A(n321), .B(n317), .Z(n366) );
  XNOR U1996 ( .A(n316), .B(n312), .Z(n367) );
  XNOR U1997 ( .A(n311), .B(n307), .Z(n368) );
  XOR U1998 ( .A(n306), .B(n303), .Z(n369) );
  XOR U1999 ( .A(n370), .B(n371), .Z(n303) );
  XOR U2000 ( .A(n301), .B(n372), .Z(n371) );
  XOR U2001 ( .A(n373), .B(n374), .Z(n372) );
  XNOR U2002 ( .A(n375), .B(n376), .Z(n374) );
  AND U2003 ( .A(b[13]), .B(a[111]), .Z(n375) );
  XOR U2004 ( .A(n377), .B(n378), .Z(n373) );
  AND U2005 ( .A(b[14]), .B(a[110]), .Z(n378) );
  AND U2006 ( .A(b[15]), .B(a[109]), .Z(n377) );
  XOR U2007 ( .A(n379), .B(n376), .Z(n370) );
  XOR U2008 ( .A(n380), .B(n381), .Z(n376) );
  NOR U2009 ( .A(n382), .B(n383), .Z(n380) );
  AND U2010 ( .A(b[12]), .B(a[112]), .Z(n379) );
  XNOR U2011 ( .A(n384), .B(n301), .Z(n302) );
  XOR U2012 ( .A(n385), .B(n386), .Z(n301) );
  ANDN U2013 ( .B(n387), .A(n388), .Z(n385) );
  AND U2014 ( .A(b[11]), .B(a[113]), .Z(n384) );
  XNOR U2015 ( .A(n389), .B(n306), .Z(n308) );
  XOR U2016 ( .A(n390), .B(n391), .Z(n306) );
  ANDN U2017 ( .B(n392), .A(n393), .Z(n390) );
  AND U2018 ( .A(b[10]), .B(a[114]), .Z(n389) );
  XNOR U2019 ( .A(n394), .B(n311), .Z(n313) );
  XOR U2020 ( .A(n395), .B(n396), .Z(n311) );
  ANDN U2021 ( .B(n397), .A(n398), .Z(n395) );
  AND U2022 ( .A(b[9]), .B(a[115]), .Z(n394) );
  XNOR U2023 ( .A(n399), .B(n316), .Z(n318) );
  XOR U2024 ( .A(n400), .B(n401), .Z(n316) );
  ANDN U2025 ( .B(n402), .A(n403), .Z(n400) );
  AND U2026 ( .A(b[8]), .B(a[116]), .Z(n399) );
  XNOR U2027 ( .A(n404), .B(n321), .Z(n323) );
  XOR U2028 ( .A(n405), .B(n406), .Z(n321) );
  ANDN U2029 ( .B(n407), .A(n408), .Z(n405) );
  AND U2030 ( .A(b[7]), .B(a[117]), .Z(n404) );
  XNOR U2031 ( .A(n409), .B(n326), .Z(n328) );
  XOR U2032 ( .A(n410), .B(n411), .Z(n326) );
  ANDN U2033 ( .B(n412), .A(n413), .Z(n410) );
  AND U2034 ( .A(b[6]), .B(a[118]), .Z(n409) );
  XNOR U2035 ( .A(n414), .B(n331), .Z(n333) );
  XOR U2036 ( .A(n415), .B(n416), .Z(n331) );
  ANDN U2037 ( .B(n417), .A(n418), .Z(n415) );
  AND U2038 ( .A(b[5]), .B(a[119]), .Z(n414) );
  XNOR U2039 ( .A(n419), .B(n336), .Z(n338) );
  XOR U2040 ( .A(n420), .B(n421), .Z(n336) );
  ANDN U2041 ( .B(n422), .A(n423), .Z(n420) );
  AND U2042 ( .A(b[4]), .B(a[120]), .Z(n419) );
  XNOR U2043 ( .A(n424), .B(n425), .Z(n350) );
  NANDN U2044 ( .A(n426), .B(n427), .Z(n425) );
  XNOR U2045 ( .A(n428), .B(n341), .Z(n343) );
  XNOR U2046 ( .A(n429), .B(n430), .Z(n341) );
  AND U2047 ( .A(n431), .B(n432), .Z(n429) );
  AND U2048 ( .A(b[3]), .B(a[121]), .Z(n428) );
  XNOR U2049 ( .A(n433), .B(n434), .Z(swire[123]) );
  XOR U2050 ( .A(n360), .B(n435), .Z(n434) );
  XOR U2051 ( .A(n359), .B(n433), .Z(n435) );
  NANDN U2052 ( .A(n179), .B(a[123]), .Z(n359) );
  XNOR U2053 ( .A(n426), .B(n427), .Z(n360) );
  XOR U2054 ( .A(n424), .B(n436), .Z(n427) );
  NAND U2055 ( .A(b[1]), .B(a[122]), .Z(n436) );
  XOR U2056 ( .A(n432), .B(n437), .Z(n426) );
  XOR U2057 ( .A(n424), .B(n431), .Z(n437) );
  XNOR U2058 ( .A(n438), .B(n430), .Z(n431) );
  AND U2059 ( .A(b[2]), .B(a[121]), .Z(n438) );
  NANDN U2060 ( .A(n439), .B(n440), .Z(n424) );
  XOR U2061 ( .A(n430), .B(n422), .Z(n441) );
  XNOR U2062 ( .A(n421), .B(n417), .Z(n442) );
  XNOR U2063 ( .A(n416), .B(n412), .Z(n443) );
  XNOR U2064 ( .A(n411), .B(n407), .Z(n444) );
  XNOR U2065 ( .A(n406), .B(n402), .Z(n445) );
  XNOR U2066 ( .A(n401), .B(n397), .Z(n446) );
  XNOR U2067 ( .A(n396), .B(n392), .Z(n447) );
  XNOR U2068 ( .A(n391), .B(n387), .Z(n448) );
  XOR U2069 ( .A(n386), .B(n383), .Z(n449) );
  XOR U2070 ( .A(n450), .B(n451), .Z(n383) );
  XOR U2071 ( .A(n381), .B(n452), .Z(n451) );
  XOR U2072 ( .A(n453), .B(n454), .Z(n452) );
  XNOR U2073 ( .A(n455), .B(n456), .Z(n454) );
  AND U2074 ( .A(b[13]), .B(a[110]), .Z(n455) );
  XOR U2075 ( .A(n457), .B(n458), .Z(n453) );
  AND U2076 ( .A(b[14]), .B(a[109]), .Z(n458) );
  AND U2077 ( .A(b[15]), .B(a[108]), .Z(n457) );
  XOR U2078 ( .A(n459), .B(n456), .Z(n450) );
  XOR U2079 ( .A(n460), .B(n461), .Z(n456) );
  NOR U2080 ( .A(n462), .B(n463), .Z(n460) );
  AND U2081 ( .A(b[12]), .B(a[111]), .Z(n459) );
  XNOR U2082 ( .A(n464), .B(n381), .Z(n382) );
  XOR U2083 ( .A(n465), .B(n466), .Z(n381) );
  ANDN U2084 ( .B(n467), .A(n468), .Z(n465) );
  AND U2085 ( .A(b[11]), .B(a[112]), .Z(n464) );
  XNOR U2086 ( .A(n469), .B(n386), .Z(n388) );
  XOR U2087 ( .A(n470), .B(n471), .Z(n386) );
  ANDN U2088 ( .B(n472), .A(n473), .Z(n470) );
  AND U2089 ( .A(b[10]), .B(a[113]), .Z(n469) );
  XNOR U2090 ( .A(n474), .B(n391), .Z(n393) );
  XOR U2091 ( .A(n475), .B(n476), .Z(n391) );
  ANDN U2092 ( .B(n477), .A(n478), .Z(n475) );
  AND U2093 ( .A(b[9]), .B(a[114]), .Z(n474) );
  XNOR U2094 ( .A(n479), .B(n396), .Z(n398) );
  XOR U2095 ( .A(n480), .B(n481), .Z(n396) );
  ANDN U2096 ( .B(n482), .A(n483), .Z(n480) );
  AND U2097 ( .A(b[8]), .B(a[115]), .Z(n479) );
  XNOR U2098 ( .A(n484), .B(n401), .Z(n403) );
  XOR U2099 ( .A(n485), .B(n486), .Z(n401) );
  ANDN U2100 ( .B(n487), .A(n488), .Z(n485) );
  AND U2101 ( .A(b[7]), .B(a[116]), .Z(n484) );
  XNOR U2102 ( .A(n489), .B(n406), .Z(n408) );
  XOR U2103 ( .A(n490), .B(n491), .Z(n406) );
  ANDN U2104 ( .B(n492), .A(n493), .Z(n490) );
  AND U2105 ( .A(b[6]), .B(a[117]), .Z(n489) );
  XNOR U2106 ( .A(n494), .B(n411), .Z(n413) );
  XOR U2107 ( .A(n495), .B(n496), .Z(n411) );
  ANDN U2108 ( .B(n497), .A(n498), .Z(n495) );
  AND U2109 ( .A(b[5]), .B(a[118]), .Z(n494) );
  XNOR U2110 ( .A(n499), .B(n416), .Z(n418) );
  XOR U2111 ( .A(n500), .B(n501), .Z(n416) );
  ANDN U2112 ( .B(n502), .A(n503), .Z(n500) );
  AND U2113 ( .A(b[4]), .B(a[119]), .Z(n499) );
  XNOR U2114 ( .A(n504), .B(n505), .Z(n430) );
  NANDN U2115 ( .A(n506), .B(n507), .Z(n505) );
  XNOR U2116 ( .A(n508), .B(n421), .Z(n423) );
  XNOR U2117 ( .A(n509), .B(n510), .Z(n421) );
  AND U2118 ( .A(n511), .B(n512), .Z(n509) );
  AND U2119 ( .A(b[3]), .B(a[120]), .Z(n508) );
  XNOR U2120 ( .A(n513), .B(n514), .Z(swire[122]) );
  XOR U2121 ( .A(n440), .B(n516), .Z(n514) );
  XNOR U2122 ( .A(n439), .B(n515), .Z(n516) );
  IV U2123 ( .A(n513), .Z(n515) );
  NANDN U2124 ( .A(n179), .B(a[122]), .Z(n439) );
  XNOR U2125 ( .A(n506), .B(n507), .Z(n440) );
  XOR U2126 ( .A(n504), .B(n517), .Z(n507) );
  NAND U2127 ( .A(b[1]), .B(a[121]), .Z(n517) );
  XOR U2128 ( .A(n512), .B(n518), .Z(n506) );
  XOR U2129 ( .A(n504), .B(n511), .Z(n518) );
  XNOR U2130 ( .A(n519), .B(n510), .Z(n511) );
  AND U2131 ( .A(b[2]), .B(a[120]), .Z(n519) );
  NANDN U2132 ( .A(n520), .B(n521), .Z(n504) );
  XOR U2133 ( .A(n510), .B(n502), .Z(n522) );
  XNOR U2134 ( .A(n501), .B(n497), .Z(n523) );
  XNOR U2135 ( .A(n496), .B(n492), .Z(n524) );
  XNOR U2136 ( .A(n491), .B(n487), .Z(n525) );
  XNOR U2137 ( .A(n486), .B(n482), .Z(n526) );
  XNOR U2138 ( .A(n481), .B(n477), .Z(n527) );
  XNOR U2139 ( .A(n476), .B(n472), .Z(n528) );
  XNOR U2140 ( .A(n471), .B(n467), .Z(n529) );
  XOR U2141 ( .A(n466), .B(n463), .Z(n530) );
  XOR U2142 ( .A(n531), .B(n532), .Z(n463) );
  XOR U2143 ( .A(n461), .B(n533), .Z(n532) );
  XOR U2144 ( .A(n534), .B(n535), .Z(n533) );
  XOR U2145 ( .A(n536), .B(n537), .Z(n535) );
  XOR U2146 ( .A(n538), .B(n539), .Z(n537) );
  XOR U2147 ( .A(n540), .B(n541), .Z(n539) );
  NAND U2148 ( .A(b[14]), .B(a[108]), .Z(n541) );
  AND U2149 ( .A(b[15]), .B(a[107]), .Z(n540) );
  XOR U2150 ( .A(n542), .B(n538), .Z(n534) );
  XOR U2151 ( .A(n543), .B(n544), .Z(n538) );
  NOR U2152 ( .A(n545), .B(n546), .Z(n543) );
  AND U2153 ( .A(b[13]), .B(a[109]), .Z(n542) );
  XOR U2154 ( .A(n547), .B(n536), .Z(n531) );
  XOR U2155 ( .A(n548), .B(n549), .Z(n536) );
  ANDN U2156 ( .B(n550), .A(n551), .Z(n548) );
  AND U2157 ( .A(b[12]), .B(a[110]), .Z(n547) );
  XNOR U2158 ( .A(n552), .B(n461), .Z(n462) );
  XOR U2159 ( .A(n553), .B(n554), .Z(n461) );
  ANDN U2160 ( .B(n555), .A(n556), .Z(n553) );
  AND U2161 ( .A(b[11]), .B(a[111]), .Z(n552) );
  XNOR U2162 ( .A(n557), .B(n466), .Z(n468) );
  XOR U2163 ( .A(n558), .B(n559), .Z(n466) );
  ANDN U2164 ( .B(n560), .A(n561), .Z(n558) );
  AND U2165 ( .A(b[10]), .B(a[112]), .Z(n557) );
  XNOR U2166 ( .A(n562), .B(n471), .Z(n473) );
  XOR U2167 ( .A(n563), .B(n564), .Z(n471) );
  ANDN U2168 ( .B(n565), .A(n566), .Z(n563) );
  AND U2169 ( .A(b[9]), .B(a[113]), .Z(n562) );
  XNOR U2170 ( .A(n567), .B(n476), .Z(n478) );
  XOR U2171 ( .A(n568), .B(n569), .Z(n476) );
  ANDN U2172 ( .B(n570), .A(n571), .Z(n568) );
  AND U2173 ( .A(b[8]), .B(a[114]), .Z(n567) );
  XNOR U2174 ( .A(n572), .B(n481), .Z(n483) );
  XOR U2175 ( .A(n573), .B(n574), .Z(n481) );
  ANDN U2176 ( .B(n575), .A(n576), .Z(n573) );
  AND U2177 ( .A(b[7]), .B(a[115]), .Z(n572) );
  XNOR U2178 ( .A(n577), .B(n486), .Z(n488) );
  XOR U2179 ( .A(n578), .B(n579), .Z(n486) );
  ANDN U2180 ( .B(n580), .A(n581), .Z(n578) );
  AND U2181 ( .A(b[6]), .B(a[116]), .Z(n577) );
  XNOR U2182 ( .A(n582), .B(n491), .Z(n493) );
  XOR U2183 ( .A(n583), .B(n584), .Z(n491) );
  ANDN U2184 ( .B(n585), .A(n586), .Z(n583) );
  AND U2185 ( .A(b[5]), .B(a[117]), .Z(n582) );
  XNOR U2186 ( .A(n587), .B(n496), .Z(n498) );
  XOR U2187 ( .A(n588), .B(n589), .Z(n496) );
  ANDN U2188 ( .B(n590), .A(n591), .Z(n588) );
  AND U2189 ( .A(b[4]), .B(a[118]), .Z(n587) );
  XNOR U2190 ( .A(n592), .B(n593), .Z(n510) );
  NANDN U2191 ( .A(n594), .B(n595), .Z(n593) );
  XNOR U2192 ( .A(n596), .B(n501), .Z(n503) );
  XNOR U2193 ( .A(n597), .B(n598), .Z(n501) );
  AND U2194 ( .A(n599), .B(n600), .Z(n597) );
  AND U2195 ( .A(b[3]), .B(a[119]), .Z(n596) );
  XNOR U2196 ( .A(n601), .B(n602), .Z(swire[121]) );
  XOR U2197 ( .A(n521), .B(n603), .Z(n602) );
  XOR U2198 ( .A(n520), .B(n601), .Z(n603) );
  NANDN U2199 ( .A(n179), .B(a[121]), .Z(n520) );
  XNOR U2200 ( .A(n594), .B(n595), .Z(n521) );
  XOR U2201 ( .A(n592), .B(n604), .Z(n595) );
  NAND U2202 ( .A(b[1]), .B(a[120]), .Z(n604) );
  XOR U2203 ( .A(n600), .B(n605), .Z(n594) );
  XOR U2204 ( .A(n592), .B(n599), .Z(n605) );
  XNOR U2205 ( .A(n606), .B(n598), .Z(n599) );
  AND U2206 ( .A(b[2]), .B(a[119]), .Z(n606) );
  NANDN U2207 ( .A(n607), .B(n608), .Z(n592) );
  XOR U2208 ( .A(n598), .B(n590), .Z(n609) );
  XNOR U2209 ( .A(n589), .B(n585), .Z(n610) );
  XNOR U2210 ( .A(n584), .B(n580), .Z(n611) );
  XNOR U2211 ( .A(n579), .B(n575), .Z(n612) );
  XNOR U2212 ( .A(n574), .B(n570), .Z(n613) );
  XNOR U2213 ( .A(n569), .B(n565), .Z(n614) );
  XNOR U2214 ( .A(n564), .B(n560), .Z(n615) );
  XNOR U2215 ( .A(n559), .B(n555), .Z(n616) );
  XNOR U2216 ( .A(n554), .B(n550), .Z(n617) );
  XOR U2217 ( .A(n549), .B(n546), .Z(n618) );
  XOR U2218 ( .A(n619), .B(n620), .Z(n546) );
  XOR U2219 ( .A(n544), .B(n621), .Z(n620) );
  XOR U2220 ( .A(n622), .B(n623), .Z(n621) );
  XOR U2221 ( .A(n624), .B(n625), .Z(n623) );
  NAND U2222 ( .A(b[14]), .B(a[107]), .Z(n625) );
  AND U2223 ( .A(b[15]), .B(a[106]), .Z(n624) );
  XOR U2224 ( .A(n626), .B(n622), .Z(n619) );
  XOR U2225 ( .A(n627), .B(n628), .Z(n622) );
  NOR U2226 ( .A(n629), .B(n630), .Z(n627) );
  AND U2227 ( .A(b[13]), .B(a[108]), .Z(n626) );
  XNOR U2228 ( .A(n631), .B(n544), .Z(n545) );
  XOR U2229 ( .A(n632), .B(n633), .Z(n544) );
  ANDN U2230 ( .B(n634), .A(n635), .Z(n632) );
  AND U2231 ( .A(b[12]), .B(a[109]), .Z(n631) );
  XNOR U2232 ( .A(n636), .B(n549), .Z(n551) );
  XOR U2233 ( .A(n637), .B(n638), .Z(n549) );
  ANDN U2234 ( .B(n639), .A(n640), .Z(n637) );
  AND U2235 ( .A(b[11]), .B(a[110]), .Z(n636) );
  XNOR U2236 ( .A(n641), .B(n554), .Z(n556) );
  XOR U2237 ( .A(n642), .B(n643), .Z(n554) );
  ANDN U2238 ( .B(n644), .A(n645), .Z(n642) );
  AND U2239 ( .A(b[10]), .B(a[111]), .Z(n641) );
  XNOR U2240 ( .A(n646), .B(n559), .Z(n561) );
  XOR U2241 ( .A(n647), .B(n648), .Z(n559) );
  ANDN U2242 ( .B(n649), .A(n650), .Z(n647) );
  AND U2243 ( .A(b[9]), .B(a[112]), .Z(n646) );
  XNOR U2244 ( .A(n651), .B(n564), .Z(n566) );
  XOR U2245 ( .A(n652), .B(n653), .Z(n564) );
  ANDN U2246 ( .B(n654), .A(n655), .Z(n652) );
  AND U2247 ( .A(b[8]), .B(a[113]), .Z(n651) );
  XNOR U2248 ( .A(n656), .B(n569), .Z(n571) );
  XOR U2249 ( .A(n657), .B(n658), .Z(n569) );
  ANDN U2250 ( .B(n659), .A(n660), .Z(n657) );
  AND U2251 ( .A(b[7]), .B(a[114]), .Z(n656) );
  XNOR U2252 ( .A(n661), .B(n574), .Z(n576) );
  XOR U2253 ( .A(n662), .B(n663), .Z(n574) );
  ANDN U2254 ( .B(n664), .A(n665), .Z(n662) );
  AND U2255 ( .A(b[6]), .B(a[115]), .Z(n661) );
  XNOR U2256 ( .A(n666), .B(n579), .Z(n581) );
  XOR U2257 ( .A(n667), .B(n668), .Z(n579) );
  ANDN U2258 ( .B(n669), .A(n670), .Z(n667) );
  AND U2259 ( .A(b[5]), .B(a[116]), .Z(n666) );
  XNOR U2260 ( .A(n671), .B(n584), .Z(n586) );
  XOR U2261 ( .A(n672), .B(n673), .Z(n584) );
  ANDN U2262 ( .B(n674), .A(n675), .Z(n672) );
  AND U2263 ( .A(b[4]), .B(a[117]), .Z(n671) );
  XNOR U2264 ( .A(n676), .B(n677), .Z(n598) );
  NANDN U2265 ( .A(n678), .B(n679), .Z(n677) );
  XNOR U2266 ( .A(n680), .B(n589), .Z(n591) );
  XNOR U2267 ( .A(n681), .B(n682), .Z(n589) );
  AND U2268 ( .A(n683), .B(n684), .Z(n681) );
  AND U2269 ( .A(b[3]), .B(a[118]), .Z(n680) );
  XNOR U2270 ( .A(n685), .B(n686), .Z(swire[120]) );
  XOR U2271 ( .A(n608), .B(n688), .Z(n686) );
  XNOR U2272 ( .A(n607), .B(n687), .Z(n688) );
  IV U2273 ( .A(n685), .Z(n687) );
  NANDN U2274 ( .A(n179), .B(a[120]), .Z(n607) );
  XNOR U2275 ( .A(n678), .B(n679), .Z(n608) );
  XOR U2276 ( .A(n676), .B(n689), .Z(n679) );
  NAND U2277 ( .A(b[1]), .B(a[119]), .Z(n689) );
  XOR U2278 ( .A(n683), .B(n690), .Z(n678) );
  XOR U2279 ( .A(n676), .B(n684), .Z(n690) );
  XNOR U2280 ( .A(n691), .B(n682), .Z(n684) );
  AND U2281 ( .A(b[2]), .B(a[118]), .Z(n691) );
  NANDN U2282 ( .A(n692), .B(n693), .Z(n676) );
  XOR U2283 ( .A(n682), .B(n674), .Z(n694) );
  XNOR U2284 ( .A(n673), .B(n669), .Z(n695) );
  XNOR U2285 ( .A(n668), .B(n664), .Z(n696) );
  XNOR U2286 ( .A(n663), .B(n659), .Z(n697) );
  XNOR U2287 ( .A(n658), .B(n654), .Z(n698) );
  XNOR U2288 ( .A(n653), .B(n649), .Z(n699) );
  XNOR U2289 ( .A(n648), .B(n644), .Z(n700) );
  XNOR U2290 ( .A(n643), .B(n639), .Z(n701) );
  XNOR U2291 ( .A(n638), .B(n634), .Z(n702) );
  XOR U2292 ( .A(n633), .B(n630), .Z(n703) );
  XOR U2293 ( .A(n704), .B(n705), .Z(n630) );
  XOR U2294 ( .A(n628), .B(n706), .Z(n705) );
  XOR U2295 ( .A(n707), .B(n708), .Z(n706) );
  XOR U2296 ( .A(n709), .B(n710), .Z(n708) );
  NAND U2297 ( .A(b[14]), .B(a[106]), .Z(n710) );
  AND U2298 ( .A(b[15]), .B(a[105]), .Z(n709) );
  XOR U2299 ( .A(n711), .B(n707), .Z(n704) );
  XOR U2300 ( .A(n712), .B(n713), .Z(n707) );
  NOR U2301 ( .A(n714), .B(n715), .Z(n712) );
  AND U2302 ( .A(b[13]), .B(a[107]), .Z(n711) );
  XNOR U2303 ( .A(n716), .B(n628), .Z(n629) );
  XOR U2304 ( .A(n717), .B(n718), .Z(n628) );
  ANDN U2305 ( .B(n719), .A(n720), .Z(n717) );
  AND U2306 ( .A(b[12]), .B(a[108]), .Z(n716) );
  XNOR U2307 ( .A(n721), .B(n633), .Z(n635) );
  XOR U2308 ( .A(n722), .B(n723), .Z(n633) );
  ANDN U2309 ( .B(n724), .A(n725), .Z(n722) );
  AND U2310 ( .A(b[11]), .B(a[109]), .Z(n721) );
  XNOR U2311 ( .A(n726), .B(n638), .Z(n640) );
  XOR U2312 ( .A(n727), .B(n728), .Z(n638) );
  ANDN U2313 ( .B(n729), .A(n730), .Z(n727) );
  AND U2314 ( .A(b[10]), .B(a[110]), .Z(n726) );
  XNOR U2315 ( .A(n731), .B(n643), .Z(n645) );
  XOR U2316 ( .A(n732), .B(n733), .Z(n643) );
  ANDN U2317 ( .B(n734), .A(n735), .Z(n732) );
  AND U2318 ( .A(b[9]), .B(a[111]), .Z(n731) );
  XNOR U2319 ( .A(n736), .B(n648), .Z(n650) );
  XOR U2320 ( .A(n737), .B(n738), .Z(n648) );
  ANDN U2321 ( .B(n739), .A(n740), .Z(n737) );
  AND U2322 ( .A(b[8]), .B(a[112]), .Z(n736) );
  XNOR U2323 ( .A(n741), .B(n653), .Z(n655) );
  XOR U2324 ( .A(n742), .B(n743), .Z(n653) );
  ANDN U2325 ( .B(n744), .A(n745), .Z(n742) );
  AND U2326 ( .A(b[7]), .B(a[113]), .Z(n741) );
  XNOR U2327 ( .A(n746), .B(n658), .Z(n660) );
  XOR U2328 ( .A(n747), .B(n748), .Z(n658) );
  ANDN U2329 ( .B(n749), .A(n750), .Z(n747) );
  AND U2330 ( .A(b[6]), .B(a[114]), .Z(n746) );
  XNOR U2331 ( .A(n751), .B(n663), .Z(n665) );
  XOR U2332 ( .A(n752), .B(n753), .Z(n663) );
  ANDN U2333 ( .B(n754), .A(n755), .Z(n752) );
  AND U2334 ( .A(b[5]), .B(a[115]), .Z(n751) );
  XNOR U2335 ( .A(n756), .B(n668), .Z(n670) );
  XOR U2336 ( .A(n757), .B(n758), .Z(n668) );
  ANDN U2337 ( .B(n759), .A(n760), .Z(n757) );
  AND U2338 ( .A(b[4]), .B(a[116]), .Z(n756) );
  XNOR U2339 ( .A(n761), .B(n762), .Z(n682) );
  NANDN U2340 ( .A(n763), .B(n764), .Z(n762) );
  XNOR U2341 ( .A(n765), .B(n673), .Z(n675) );
  XNOR U2342 ( .A(n766), .B(n767), .Z(n673) );
  NOR U2343 ( .A(n768), .B(n769), .Z(n766) );
  AND U2344 ( .A(b[3]), .B(a[117]), .Z(n765) );
  XNOR U2345 ( .A(n770), .B(n771), .Z(swire[119]) );
  XOR U2346 ( .A(n693), .B(n772), .Z(n771) );
  XOR U2347 ( .A(n692), .B(n770), .Z(n772) );
  NANDN U2348 ( .A(n179), .B(a[119]), .Z(n692) );
  XOR U2349 ( .A(n773), .B(n774), .Z(n763) );
  NAND U2350 ( .A(b[1]), .B(a[118]), .Z(n774) );
  XOR U2351 ( .A(n773), .B(n769), .Z(n775) );
  XOR U2352 ( .A(n776), .B(n767), .Z(n769) );
  AND U2353 ( .A(b[2]), .B(a[117]), .Z(n776) );
  IV U2354 ( .A(n761), .Z(n773) );
  NANDN U2355 ( .A(n777), .B(n778), .Z(n761) );
  XOR U2356 ( .A(n767), .B(n759), .Z(n779) );
  XNOR U2357 ( .A(n758), .B(n754), .Z(n780) );
  XNOR U2358 ( .A(n753), .B(n749), .Z(n781) );
  XNOR U2359 ( .A(n748), .B(n744), .Z(n782) );
  XNOR U2360 ( .A(n743), .B(n739), .Z(n783) );
  XNOR U2361 ( .A(n738), .B(n734), .Z(n784) );
  XNOR U2362 ( .A(n733), .B(n729), .Z(n785) );
  XNOR U2363 ( .A(n728), .B(n724), .Z(n786) );
  XNOR U2364 ( .A(n723), .B(n719), .Z(n787) );
  XOR U2365 ( .A(n718), .B(n715), .Z(n788) );
  XOR U2366 ( .A(n789), .B(n790), .Z(n715) );
  XOR U2367 ( .A(n713), .B(n791), .Z(n790) );
  XOR U2368 ( .A(n792), .B(n793), .Z(n791) );
  XOR U2369 ( .A(n794), .B(n795), .Z(n793) );
  NAND U2370 ( .A(b[14]), .B(a[105]), .Z(n795) );
  AND U2371 ( .A(b[15]), .B(a[104]), .Z(n794) );
  XOR U2372 ( .A(n796), .B(n792), .Z(n789) );
  XOR U2373 ( .A(n797), .B(n798), .Z(n792) );
  NOR U2374 ( .A(n799), .B(n800), .Z(n797) );
  AND U2375 ( .A(b[13]), .B(a[106]), .Z(n796) );
  XNOR U2376 ( .A(n801), .B(n713), .Z(n714) );
  XOR U2377 ( .A(n802), .B(n803), .Z(n713) );
  ANDN U2378 ( .B(n804), .A(n805), .Z(n802) );
  AND U2379 ( .A(b[12]), .B(a[107]), .Z(n801) );
  XNOR U2380 ( .A(n806), .B(n718), .Z(n720) );
  XOR U2381 ( .A(n807), .B(n808), .Z(n718) );
  ANDN U2382 ( .B(n809), .A(n810), .Z(n807) );
  AND U2383 ( .A(b[11]), .B(a[108]), .Z(n806) );
  XNOR U2384 ( .A(n811), .B(n723), .Z(n725) );
  XOR U2385 ( .A(n812), .B(n813), .Z(n723) );
  ANDN U2386 ( .B(n814), .A(n815), .Z(n812) );
  AND U2387 ( .A(b[10]), .B(a[109]), .Z(n811) );
  XNOR U2388 ( .A(n816), .B(n728), .Z(n730) );
  XOR U2389 ( .A(n817), .B(n818), .Z(n728) );
  ANDN U2390 ( .B(n819), .A(n820), .Z(n817) );
  AND U2391 ( .A(b[9]), .B(a[110]), .Z(n816) );
  XNOR U2392 ( .A(n821), .B(n733), .Z(n735) );
  XOR U2393 ( .A(n822), .B(n823), .Z(n733) );
  ANDN U2394 ( .B(n824), .A(n825), .Z(n822) );
  AND U2395 ( .A(b[8]), .B(a[111]), .Z(n821) );
  XNOR U2396 ( .A(n826), .B(n738), .Z(n740) );
  XOR U2397 ( .A(n827), .B(n828), .Z(n738) );
  ANDN U2398 ( .B(n829), .A(n830), .Z(n827) );
  AND U2399 ( .A(b[7]), .B(a[112]), .Z(n826) );
  XNOR U2400 ( .A(n831), .B(n743), .Z(n745) );
  XOR U2401 ( .A(n832), .B(n833), .Z(n743) );
  ANDN U2402 ( .B(n834), .A(n835), .Z(n832) );
  AND U2403 ( .A(b[6]), .B(a[113]), .Z(n831) );
  XNOR U2404 ( .A(n836), .B(n748), .Z(n750) );
  XOR U2405 ( .A(n837), .B(n838), .Z(n748) );
  ANDN U2406 ( .B(n839), .A(n840), .Z(n837) );
  AND U2407 ( .A(b[5]), .B(a[114]), .Z(n836) );
  XNOR U2408 ( .A(n841), .B(n753), .Z(n755) );
  XOR U2409 ( .A(n842), .B(n843), .Z(n753) );
  ANDN U2410 ( .B(n844), .A(n845), .Z(n842) );
  AND U2411 ( .A(b[4]), .B(a[115]), .Z(n841) );
  XOR U2412 ( .A(n846), .B(n847), .Z(n767) );
  NANDN U2413 ( .A(n848), .B(n849), .Z(n847) );
  XNOR U2414 ( .A(n850), .B(n758), .Z(n760) );
  XNOR U2415 ( .A(n851), .B(n852), .Z(n758) );
  AND U2416 ( .A(n853), .B(n854), .Z(n851) );
  AND U2417 ( .A(b[3]), .B(a[116]), .Z(n850) );
  XNOR U2418 ( .A(n855), .B(n856), .Z(swire[118]) );
  XOR U2419 ( .A(n778), .B(n858), .Z(n856) );
  XNOR U2420 ( .A(n777), .B(n857), .Z(n858) );
  IV U2421 ( .A(n855), .Z(n857) );
  NANDN U2422 ( .A(n179), .B(a[118]), .Z(n777) );
  XNOR U2423 ( .A(n849), .B(n848), .Z(n778) );
  XOR U2424 ( .A(n846), .B(n859), .Z(n848) );
  NAND U2425 ( .A(b[1]), .B(a[117]), .Z(n859) );
  XNOR U2426 ( .A(n854), .B(n860), .Z(n849) );
  XNOR U2427 ( .A(n846), .B(n853), .Z(n860) );
  XNOR U2428 ( .A(n861), .B(n852), .Z(n853) );
  AND U2429 ( .A(b[2]), .B(a[116]), .Z(n861) );
  ANDN U2430 ( .B(n862), .A(n863), .Z(n846) );
  XOR U2431 ( .A(n852), .B(n844), .Z(n864) );
  XNOR U2432 ( .A(n843), .B(n839), .Z(n865) );
  XNOR U2433 ( .A(n838), .B(n834), .Z(n866) );
  XNOR U2434 ( .A(n833), .B(n829), .Z(n867) );
  XNOR U2435 ( .A(n828), .B(n824), .Z(n868) );
  XNOR U2436 ( .A(n823), .B(n819), .Z(n869) );
  XNOR U2437 ( .A(n818), .B(n814), .Z(n870) );
  XNOR U2438 ( .A(n813), .B(n809), .Z(n871) );
  XNOR U2439 ( .A(n808), .B(n804), .Z(n872) );
  XOR U2440 ( .A(n803), .B(n800), .Z(n873) );
  XOR U2441 ( .A(n874), .B(n875), .Z(n800) );
  XOR U2442 ( .A(n798), .B(n876), .Z(n875) );
  XOR U2443 ( .A(n877), .B(n878), .Z(n876) );
  XOR U2444 ( .A(n879), .B(n880), .Z(n878) );
  NAND U2445 ( .A(b[14]), .B(a[104]), .Z(n880) );
  AND U2446 ( .A(b[15]), .B(a[103]), .Z(n879) );
  XOR U2447 ( .A(n881), .B(n877), .Z(n874) );
  XOR U2448 ( .A(n882), .B(n883), .Z(n877) );
  NOR U2449 ( .A(n884), .B(n885), .Z(n882) );
  AND U2450 ( .A(b[13]), .B(a[105]), .Z(n881) );
  XNOR U2451 ( .A(n886), .B(n798), .Z(n799) );
  XOR U2452 ( .A(n887), .B(n888), .Z(n798) );
  ANDN U2453 ( .B(n889), .A(n890), .Z(n887) );
  AND U2454 ( .A(b[12]), .B(a[106]), .Z(n886) );
  XNOR U2455 ( .A(n891), .B(n803), .Z(n805) );
  XOR U2456 ( .A(n892), .B(n893), .Z(n803) );
  ANDN U2457 ( .B(n894), .A(n895), .Z(n892) );
  AND U2458 ( .A(b[11]), .B(a[107]), .Z(n891) );
  XNOR U2459 ( .A(n896), .B(n808), .Z(n810) );
  XOR U2460 ( .A(n897), .B(n898), .Z(n808) );
  ANDN U2461 ( .B(n899), .A(n900), .Z(n897) );
  AND U2462 ( .A(b[10]), .B(a[108]), .Z(n896) );
  XNOR U2463 ( .A(n901), .B(n813), .Z(n815) );
  XOR U2464 ( .A(n902), .B(n903), .Z(n813) );
  ANDN U2465 ( .B(n904), .A(n905), .Z(n902) );
  AND U2466 ( .A(b[9]), .B(a[109]), .Z(n901) );
  XNOR U2467 ( .A(n906), .B(n818), .Z(n820) );
  XOR U2468 ( .A(n907), .B(n908), .Z(n818) );
  ANDN U2469 ( .B(n909), .A(n910), .Z(n907) );
  AND U2470 ( .A(b[8]), .B(a[110]), .Z(n906) );
  XNOR U2471 ( .A(n911), .B(n823), .Z(n825) );
  XOR U2472 ( .A(n912), .B(n913), .Z(n823) );
  ANDN U2473 ( .B(n914), .A(n915), .Z(n912) );
  AND U2474 ( .A(b[7]), .B(a[111]), .Z(n911) );
  XNOR U2475 ( .A(n916), .B(n828), .Z(n830) );
  XOR U2476 ( .A(n917), .B(n918), .Z(n828) );
  ANDN U2477 ( .B(n919), .A(n920), .Z(n917) );
  AND U2478 ( .A(b[6]), .B(a[112]), .Z(n916) );
  XNOR U2479 ( .A(n921), .B(n833), .Z(n835) );
  XOR U2480 ( .A(n922), .B(n923), .Z(n833) );
  ANDN U2481 ( .B(n924), .A(n925), .Z(n922) );
  AND U2482 ( .A(b[5]), .B(a[113]), .Z(n921) );
  XNOR U2483 ( .A(n926), .B(n838), .Z(n840) );
  XOR U2484 ( .A(n927), .B(n928), .Z(n838) );
  ANDN U2485 ( .B(n929), .A(n930), .Z(n927) );
  AND U2486 ( .A(b[4]), .B(a[114]), .Z(n926) );
  XNOR U2487 ( .A(n931), .B(n932), .Z(n852) );
  NANDN U2488 ( .A(n933), .B(n934), .Z(n932) );
  XNOR U2489 ( .A(n935), .B(n843), .Z(n845) );
  XNOR U2490 ( .A(n936), .B(n937), .Z(n843) );
  AND U2491 ( .A(n938), .B(n939), .Z(n936) );
  AND U2492 ( .A(b[3]), .B(a[115]), .Z(n935) );
  XNOR U2493 ( .A(n940), .B(n941), .Z(swire[117]) );
  XOR U2494 ( .A(n862), .B(n942), .Z(n941) );
  XOR U2495 ( .A(n863), .B(n940), .Z(n942) );
  NANDN U2496 ( .A(n179), .B(a[117]), .Z(n863) );
  XNOR U2497 ( .A(n933), .B(n934), .Z(n862) );
  XOR U2498 ( .A(n931), .B(n943), .Z(n934) );
  NAND U2499 ( .A(b[1]), .B(a[116]), .Z(n943) );
  XOR U2500 ( .A(n939), .B(n944), .Z(n933) );
  XOR U2501 ( .A(n931), .B(n938), .Z(n944) );
  XNOR U2502 ( .A(n945), .B(n937), .Z(n938) );
  AND U2503 ( .A(b[2]), .B(a[115]), .Z(n945) );
  NANDN U2504 ( .A(n946), .B(n947), .Z(n931) );
  XOR U2505 ( .A(n937), .B(n929), .Z(n948) );
  XNOR U2506 ( .A(n928), .B(n924), .Z(n949) );
  XNOR U2507 ( .A(n923), .B(n919), .Z(n950) );
  XNOR U2508 ( .A(n918), .B(n914), .Z(n951) );
  XNOR U2509 ( .A(n913), .B(n909), .Z(n952) );
  XNOR U2510 ( .A(n908), .B(n904), .Z(n953) );
  XNOR U2511 ( .A(n903), .B(n899), .Z(n954) );
  XNOR U2512 ( .A(n898), .B(n894), .Z(n955) );
  XNOR U2513 ( .A(n893), .B(n889), .Z(n956) );
  XOR U2514 ( .A(n888), .B(n885), .Z(n957) );
  XOR U2515 ( .A(n958), .B(n959), .Z(n885) );
  XOR U2516 ( .A(n883), .B(n960), .Z(n959) );
  XOR U2517 ( .A(n961), .B(n962), .Z(n960) );
  XOR U2518 ( .A(n963), .B(n964), .Z(n962) );
  NAND U2519 ( .A(b[14]), .B(a[103]), .Z(n964) );
  AND U2520 ( .A(b[15]), .B(a[102]), .Z(n963) );
  XOR U2521 ( .A(n965), .B(n961), .Z(n958) );
  XOR U2522 ( .A(n966), .B(n967), .Z(n961) );
  NOR U2523 ( .A(n968), .B(n969), .Z(n966) );
  AND U2524 ( .A(b[13]), .B(a[104]), .Z(n965) );
  XNOR U2525 ( .A(n970), .B(n883), .Z(n884) );
  XOR U2526 ( .A(n971), .B(n972), .Z(n883) );
  ANDN U2527 ( .B(n973), .A(n974), .Z(n971) );
  AND U2528 ( .A(b[12]), .B(a[105]), .Z(n970) );
  XNOR U2529 ( .A(n975), .B(n888), .Z(n890) );
  XOR U2530 ( .A(n976), .B(n977), .Z(n888) );
  ANDN U2531 ( .B(n978), .A(n979), .Z(n976) );
  AND U2532 ( .A(b[11]), .B(a[106]), .Z(n975) );
  XNOR U2533 ( .A(n980), .B(n893), .Z(n895) );
  XOR U2534 ( .A(n981), .B(n982), .Z(n893) );
  ANDN U2535 ( .B(n983), .A(n984), .Z(n981) );
  AND U2536 ( .A(b[10]), .B(a[107]), .Z(n980) );
  XNOR U2537 ( .A(n985), .B(n898), .Z(n900) );
  XOR U2538 ( .A(n986), .B(n987), .Z(n898) );
  ANDN U2539 ( .B(n988), .A(n989), .Z(n986) );
  AND U2540 ( .A(b[9]), .B(a[108]), .Z(n985) );
  XNOR U2541 ( .A(n990), .B(n903), .Z(n905) );
  XOR U2542 ( .A(n991), .B(n992), .Z(n903) );
  ANDN U2543 ( .B(n993), .A(n994), .Z(n991) );
  AND U2544 ( .A(b[8]), .B(a[109]), .Z(n990) );
  XNOR U2545 ( .A(n995), .B(n908), .Z(n910) );
  XOR U2546 ( .A(n996), .B(n997), .Z(n908) );
  ANDN U2547 ( .B(n998), .A(n999), .Z(n996) );
  AND U2548 ( .A(b[7]), .B(a[110]), .Z(n995) );
  XNOR U2549 ( .A(n1000), .B(n913), .Z(n915) );
  XOR U2550 ( .A(n1001), .B(n1002), .Z(n913) );
  ANDN U2551 ( .B(n1003), .A(n1004), .Z(n1001) );
  AND U2552 ( .A(b[6]), .B(a[111]), .Z(n1000) );
  XNOR U2553 ( .A(n1005), .B(n918), .Z(n920) );
  XOR U2554 ( .A(n1006), .B(n1007), .Z(n918) );
  ANDN U2555 ( .B(n1008), .A(n1009), .Z(n1006) );
  AND U2556 ( .A(b[5]), .B(a[112]), .Z(n1005) );
  XNOR U2557 ( .A(n1010), .B(n923), .Z(n925) );
  XOR U2558 ( .A(n1011), .B(n1012), .Z(n923) );
  ANDN U2559 ( .B(n1013), .A(n1014), .Z(n1011) );
  AND U2560 ( .A(b[4]), .B(a[113]), .Z(n1010) );
  XNOR U2561 ( .A(n1015), .B(n1016), .Z(n937) );
  NANDN U2562 ( .A(n1017), .B(n1018), .Z(n1016) );
  XNOR U2563 ( .A(n1019), .B(n928), .Z(n930) );
  XNOR U2564 ( .A(n1020), .B(n1021), .Z(n928) );
  AND U2565 ( .A(n1022), .B(n1023), .Z(n1020) );
  AND U2566 ( .A(b[3]), .B(a[114]), .Z(n1019) );
  XNOR U2567 ( .A(n1024), .B(n1025), .Z(swire[116]) );
  XOR U2568 ( .A(n947), .B(n1027), .Z(n1025) );
  XNOR U2569 ( .A(n946), .B(n1026), .Z(n1027) );
  IV U2570 ( .A(n1024), .Z(n1026) );
  NANDN U2571 ( .A(n179), .B(a[116]), .Z(n946) );
  XNOR U2572 ( .A(n1017), .B(n1018), .Z(n947) );
  XOR U2573 ( .A(n1015), .B(n1028), .Z(n1018) );
  NAND U2574 ( .A(b[1]), .B(a[115]), .Z(n1028) );
  XOR U2575 ( .A(n1023), .B(n1029), .Z(n1017) );
  XOR U2576 ( .A(n1015), .B(n1022), .Z(n1029) );
  XNOR U2577 ( .A(n1030), .B(n1021), .Z(n1022) );
  AND U2578 ( .A(b[2]), .B(a[114]), .Z(n1030) );
  NANDN U2579 ( .A(n1031), .B(n1032), .Z(n1015) );
  XOR U2580 ( .A(n1021), .B(n1013), .Z(n1033) );
  XNOR U2581 ( .A(n1012), .B(n1008), .Z(n1034) );
  XNOR U2582 ( .A(n1007), .B(n1003), .Z(n1035) );
  XNOR U2583 ( .A(n1002), .B(n998), .Z(n1036) );
  XNOR U2584 ( .A(n997), .B(n993), .Z(n1037) );
  XNOR U2585 ( .A(n992), .B(n988), .Z(n1038) );
  XNOR U2586 ( .A(n987), .B(n983), .Z(n1039) );
  XNOR U2587 ( .A(n982), .B(n978), .Z(n1040) );
  XNOR U2588 ( .A(n977), .B(n973), .Z(n1041) );
  XOR U2589 ( .A(n972), .B(n969), .Z(n1042) );
  XOR U2590 ( .A(n1043), .B(n1044), .Z(n969) );
  XOR U2591 ( .A(n967), .B(n1045), .Z(n1044) );
  XOR U2592 ( .A(n1046), .B(n1047), .Z(n1045) );
  XOR U2593 ( .A(n1048), .B(n1049), .Z(n1047) );
  NAND U2594 ( .A(b[14]), .B(a[102]), .Z(n1049) );
  AND U2595 ( .A(b[15]), .B(a[101]), .Z(n1048) );
  XOR U2596 ( .A(n1050), .B(n1046), .Z(n1043) );
  XOR U2597 ( .A(n1051), .B(n1052), .Z(n1046) );
  NOR U2598 ( .A(n1053), .B(n1054), .Z(n1051) );
  AND U2599 ( .A(b[13]), .B(a[103]), .Z(n1050) );
  XNOR U2600 ( .A(n1055), .B(n967), .Z(n968) );
  XOR U2601 ( .A(n1056), .B(n1057), .Z(n967) );
  ANDN U2602 ( .B(n1058), .A(n1059), .Z(n1056) );
  AND U2603 ( .A(b[12]), .B(a[104]), .Z(n1055) );
  XNOR U2604 ( .A(n1060), .B(n972), .Z(n974) );
  XOR U2605 ( .A(n1061), .B(n1062), .Z(n972) );
  ANDN U2606 ( .B(n1063), .A(n1064), .Z(n1061) );
  AND U2607 ( .A(b[11]), .B(a[105]), .Z(n1060) );
  XNOR U2608 ( .A(n1065), .B(n977), .Z(n979) );
  XOR U2609 ( .A(n1066), .B(n1067), .Z(n977) );
  ANDN U2610 ( .B(n1068), .A(n1069), .Z(n1066) );
  AND U2611 ( .A(b[10]), .B(a[106]), .Z(n1065) );
  XNOR U2612 ( .A(n1070), .B(n982), .Z(n984) );
  XOR U2613 ( .A(n1071), .B(n1072), .Z(n982) );
  ANDN U2614 ( .B(n1073), .A(n1074), .Z(n1071) );
  AND U2615 ( .A(b[9]), .B(a[107]), .Z(n1070) );
  XNOR U2616 ( .A(n1075), .B(n987), .Z(n989) );
  XOR U2617 ( .A(n1076), .B(n1077), .Z(n987) );
  ANDN U2618 ( .B(n1078), .A(n1079), .Z(n1076) );
  AND U2619 ( .A(b[8]), .B(a[108]), .Z(n1075) );
  XNOR U2620 ( .A(n1080), .B(n992), .Z(n994) );
  XOR U2621 ( .A(n1081), .B(n1082), .Z(n992) );
  ANDN U2622 ( .B(n1083), .A(n1084), .Z(n1081) );
  AND U2623 ( .A(b[7]), .B(a[109]), .Z(n1080) );
  XNOR U2624 ( .A(n1085), .B(n997), .Z(n999) );
  XOR U2625 ( .A(n1086), .B(n1087), .Z(n997) );
  ANDN U2626 ( .B(n1088), .A(n1089), .Z(n1086) );
  AND U2627 ( .A(b[6]), .B(a[110]), .Z(n1085) );
  XNOR U2628 ( .A(n1090), .B(n1002), .Z(n1004) );
  XOR U2629 ( .A(n1091), .B(n1092), .Z(n1002) );
  ANDN U2630 ( .B(n1093), .A(n1094), .Z(n1091) );
  AND U2631 ( .A(b[5]), .B(a[111]), .Z(n1090) );
  XNOR U2632 ( .A(n1095), .B(n1007), .Z(n1009) );
  XOR U2633 ( .A(n1096), .B(n1097), .Z(n1007) );
  ANDN U2634 ( .B(n1098), .A(n1099), .Z(n1096) );
  AND U2635 ( .A(b[4]), .B(a[112]), .Z(n1095) );
  XNOR U2636 ( .A(n1100), .B(n1101), .Z(n1021) );
  NANDN U2637 ( .A(n1102), .B(n1103), .Z(n1101) );
  XNOR U2638 ( .A(n1104), .B(n1012), .Z(n1014) );
  XNOR U2639 ( .A(n1105), .B(n1106), .Z(n1012) );
  AND U2640 ( .A(n1107), .B(n1108), .Z(n1105) );
  AND U2641 ( .A(b[3]), .B(a[113]), .Z(n1104) );
  XNOR U2642 ( .A(n1109), .B(n1110), .Z(swire[115]) );
  XOR U2643 ( .A(n1032), .B(n1111), .Z(n1110) );
  XOR U2644 ( .A(n1031), .B(n1109), .Z(n1111) );
  NANDN U2645 ( .A(n179), .B(a[115]), .Z(n1031) );
  XNOR U2646 ( .A(n1102), .B(n1103), .Z(n1032) );
  XOR U2647 ( .A(n1100), .B(n1112), .Z(n1103) );
  NAND U2648 ( .A(b[1]), .B(a[114]), .Z(n1112) );
  XOR U2649 ( .A(n1108), .B(n1113), .Z(n1102) );
  XOR U2650 ( .A(n1100), .B(n1107), .Z(n1113) );
  XNOR U2651 ( .A(n1114), .B(n1106), .Z(n1107) );
  AND U2652 ( .A(b[2]), .B(a[113]), .Z(n1114) );
  NANDN U2653 ( .A(n1115), .B(n1116), .Z(n1100) );
  XOR U2654 ( .A(n1106), .B(n1098), .Z(n1117) );
  XNOR U2655 ( .A(n1097), .B(n1093), .Z(n1118) );
  XNOR U2656 ( .A(n1092), .B(n1088), .Z(n1119) );
  XNOR U2657 ( .A(n1087), .B(n1083), .Z(n1120) );
  XNOR U2658 ( .A(n1082), .B(n1078), .Z(n1121) );
  XNOR U2659 ( .A(n1077), .B(n1073), .Z(n1122) );
  XNOR U2660 ( .A(n1072), .B(n1068), .Z(n1123) );
  XNOR U2661 ( .A(n1067), .B(n1063), .Z(n1124) );
  XNOR U2662 ( .A(n1062), .B(n1058), .Z(n1125) );
  XOR U2663 ( .A(n1057), .B(n1054), .Z(n1126) );
  XOR U2664 ( .A(n1127), .B(n1128), .Z(n1054) );
  XOR U2665 ( .A(n1052), .B(n1129), .Z(n1128) );
  XOR U2666 ( .A(n1130), .B(n1131), .Z(n1129) );
  XOR U2667 ( .A(n1132), .B(n1133), .Z(n1131) );
  NAND U2668 ( .A(b[14]), .B(a[101]), .Z(n1133) );
  AND U2669 ( .A(b[15]), .B(a[100]), .Z(n1132) );
  XOR U2670 ( .A(n1134), .B(n1130), .Z(n1127) );
  XOR U2671 ( .A(n1135), .B(n1136), .Z(n1130) );
  NOR U2672 ( .A(n1137), .B(n1138), .Z(n1135) );
  AND U2673 ( .A(b[13]), .B(a[102]), .Z(n1134) );
  XNOR U2674 ( .A(n1139), .B(n1052), .Z(n1053) );
  XOR U2675 ( .A(n1140), .B(n1141), .Z(n1052) );
  ANDN U2676 ( .B(n1142), .A(n1143), .Z(n1140) );
  AND U2677 ( .A(b[12]), .B(a[103]), .Z(n1139) );
  XNOR U2678 ( .A(n1144), .B(n1057), .Z(n1059) );
  XOR U2679 ( .A(n1145), .B(n1146), .Z(n1057) );
  ANDN U2680 ( .B(n1147), .A(n1148), .Z(n1145) );
  AND U2681 ( .A(b[11]), .B(a[104]), .Z(n1144) );
  XNOR U2682 ( .A(n1149), .B(n1062), .Z(n1064) );
  XOR U2683 ( .A(n1150), .B(n1151), .Z(n1062) );
  ANDN U2684 ( .B(n1152), .A(n1153), .Z(n1150) );
  AND U2685 ( .A(b[10]), .B(a[105]), .Z(n1149) );
  XNOR U2686 ( .A(n1154), .B(n1067), .Z(n1069) );
  XOR U2687 ( .A(n1155), .B(n1156), .Z(n1067) );
  ANDN U2688 ( .B(n1157), .A(n1158), .Z(n1155) );
  AND U2689 ( .A(b[9]), .B(a[106]), .Z(n1154) );
  XNOR U2690 ( .A(n1159), .B(n1072), .Z(n1074) );
  XOR U2691 ( .A(n1160), .B(n1161), .Z(n1072) );
  ANDN U2692 ( .B(n1162), .A(n1163), .Z(n1160) );
  AND U2693 ( .A(b[8]), .B(a[107]), .Z(n1159) );
  XNOR U2694 ( .A(n1164), .B(n1077), .Z(n1079) );
  XOR U2695 ( .A(n1165), .B(n1166), .Z(n1077) );
  ANDN U2696 ( .B(n1167), .A(n1168), .Z(n1165) );
  AND U2697 ( .A(b[7]), .B(a[108]), .Z(n1164) );
  XNOR U2698 ( .A(n1169), .B(n1082), .Z(n1084) );
  XOR U2699 ( .A(n1170), .B(n1171), .Z(n1082) );
  ANDN U2700 ( .B(n1172), .A(n1173), .Z(n1170) );
  AND U2701 ( .A(b[6]), .B(a[109]), .Z(n1169) );
  XNOR U2702 ( .A(n1174), .B(n1087), .Z(n1089) );
  XOR U2703 ( .A(n1175), .B(n1176), .Z(n1087) );
  ANDN U2704 ( .B(n1177), .A(n1178), .Z(n1175) );
  AND U2705 ( .A(b[5]), .B(a[110]), .Z(n1174) );
  XNOR U2706 ( .A(n1179), .B(n1092), .Z(n1094) );
  XOR U2707 ( .A(n1180), .B(n1181), .Z(n1092) );
  ANDN U2708 ( .B(n1182), .A(n1183), .Z(n1180) );
  AND U2709 ( .A(b[4]), .B(a[111]), .Z(n1179) );
  XNOR U2710 ( .A(n1184), .B(n1185), .Z(n1106) );
  NANDN U2711 ( .A(n1186), .B(n1187), .Z(n1185) );
  XNOR U2712 ( .A(n1188), .B(n1097), .Z(n1099) );
  XNOR U2713 ( .A(n1189), .B(n1190), .Z(n1097) );
  AND U2714 ( .A(n1191), .B(n1192), .Z(n1189) );
  AND U2715 ( .A(b[3]), .B(a[112]), .Z(n1188) );
  XNOR U2716 ( .A(n1193), .B(n1194), .Z(swire[114]) );
  XOR U2717 ( .A(n1116), .B(n1196), .Z(n1194) );
  XNOR U2718 ( .A(n1115), .B(n1195), .Z(n1196) );
  IV U2719 ( .A(n1193), .Z(n1195) );
  NANDN U2720 ( .A(n179), .B(a[114]), .Z(n1115) );
  XNOR U2721 ( .A(n1186), .B(n1187), .Z(n1116) );
  XOR U2722 ( .A(n1184), .B(n1197), .Z(n1187) );
  NAND U2723 ( .A(b[1]), .B(a[113]), .Z(n1197) );
  XOR U2724 ( .A(n1192), .B(n1198), .Z(n1186) );
  XOR U2725 ( .A(n1184), .B(n1191), .Z(n1198) );
  XNOR U2726 ( .A(n1199), .B(n1190), .Z(n1191) );
  AND U2727 ( .A(b[2]), .B(a[112]), .Z(n1199) );
  NANDN U2728 ( .A(n1200), .B(n1201), .Z(n1184) );
  XOR U2729 ( .A(n1190), .B(n1182), .Z(n1202) );
  XNOR U2730 ( .A(n1181), .B(n1177), .Z(n1203) );
  XNOR U2731 ( .A(n1176), .B(n1172), .Z(n1204) );
  XNOR U2732 ( .A(n1171), .B(n1167), .Z(n1205) );
  XNOR U2733 ( .A(n1166), .B(n1162), .Z(n1206) );
  XNOR U2734 ( .A(n1161), .B(n1157), .Z(n1207) );
  XNOR U2735 ( .A(n1156), .B(n1152), .Z(n1208) );
  XNOR U2736 ( .A(n1151), .B(n1147), .Z(n1209) );
  XNOR U2737 ( .A(n1146), .B(n1142), .Z(n1210) );
  XOR U2738 ( .A(n1141), .B(n1138), .Z(n1211) );
  XOR U2739 ( .A(n1212), .B(n1213), .Z(n1138) );
  XOR U2740 ( .A(n1136), .B(n1214), .Z(n1213) );
  XOR U2741 ( .A(n1215), .B(n1216), .Z(n1214) );
  XOR U2742 ( .A(n1217), .B(n1218), .Z(n1216) );
  NAND U2743 ( .A(b[14]), .B(a[100]), .Z(n1218) );
  AND U2744 ( .A(b[15]), .B(a[99]), .Z(n1217) );
  XOR U2745 ( .A(n1219), .B(n1215), .Z(n1212) );
  XOR U2746 ( .A(n1220), .B(n1221), .Z(n1215) );
  NOR U2747 ( .A(n1222), .B(n1223), .Z(n1220) );
  AND U2748 ( .A(b[13]), .B(a[101]), .Z(n1219) );
  XNOR U2749 ( .A(n1224), .B(n1136), .Z(n1137) );
  XOR U2750 ( .A(n1225), .B(n1226), .Z(n1136) );
  ANDN U2751 ( .B(n1227), .A(n1228), .Z(n1225) );
  AND U2752 ( .A(b[12]), .B(a[102]), .Z(n1224) );
  XNOR U2753 ( .A(n1229), .B(n1141), .Z(n1143) );
  XOR U2754 ( .A(n1230), .B(n1231), .Z(n1141) );
  ANDN U2755 ( .B(n1232), .A(n1233), .Z(n1230) );
  AND U2756 ( .A(b[11]), .B(a[103]), .Z(n1229) );
  XNOR U2757 ( .A(n1234), .B(n1146), .Z(n1148) );
  XOR U2758 ( .A(n1235), .B(n1236), .Z(n1146) );
  ANDN U2759 ( .B(n1237), .A(n1238), .Z(n1235) );
  AND U2760 ( .A(b[10]), .B(a[104]), .Z(n1234) );
  XNOR U2761 ( .A(n1239), .B(n1151), .Z(n1153) );
  XOR U2762 ( .A(n1240), .B(n1241), .Z(n1151) );
  ANDN U2763 ( .B(n1242), .A(n1243), .Z(n1240) );
  AND U2764 ( .A(b[9]), .B(a[105]), .Z(n1239) );
  XNOR U2765 ( .A(n1244), .B(n1156), .Z(n1158) );
  XOR U2766 ( .A(n1245), .B(n1246), .Z(n1156) );
  ANDN U2767 ( .B(n1247), .A(n1248), .Z(n1245) );
  AND U2768 ( .A(b[8]), .B(a[106]), .Z(n1244) );
  XNOR U2769 ( .A(n1249), .B(n1161), .Z(n1163) );
  XOR U2770 ( .A(n1250), .B(n1251), .Z(n1161) );
  ANDN U2771 ( .B(n1252), .A(n1253), .Z(n1250) );
  AND U2772 ( .A(b[7]), .B(a[107]), .Z(n1249) );
  XNOR U2773 ( .A(n1254), .B(n1166), .Z(n1168) );
  XOR U2774 ( .A(n1255), .B(n1256), .Z(n1166) );
  ANDN U2775 ( .B(n1257), .A(n1258), .Z(n1255) );
  AND U2776 ( .A(b[6]), .B(a[108]), .Z(n1254) );
  XNOR U2777 ( .A(n1259), .B(n1171), .Z(n1173) );
  XOR U2778 ( .A(n1260), .B(n1261), .Z(n1171) );
  ANDN U2779 ( .B(n1262), .A(n1263), .Z(n1260) );
  AND U2780 ( .A(b[5]), .B(a[109]), .Z(n1259) );
  XNOR U2781 ( .A(n1264), .B(n1176), .Z(n1178) );
  XOR U2782 ( .A(n1265), .B(n1266), .Z(n1176) );
  ANDN U2783 ( .B(n1267), .A(n1268), .Z(n1265) );
  AND U2784 ( .A(b[4]), .B(a[110]), .Z(n1264) );
  XNOR U2785 ( .A(n1269), .B(n1270), .Z(n1190) );
  NANDN U2786 ( .A(n1271), .B(n1272), .Z(n1270) );
  XNOR U2787 ( .A(n1273), .B(n1181), .Z(n1183) );
  XNOR U2788 ( .A(n1274), .B(n1275), .Z(n1181) );
  AND U2789 ( .A(n1276), .B(n1277), .Z(n1274) );
  AND U2790 ( .A(b[3]), .B(a[111]), .Z(n1273) );
  XNOR U2791 ( .A(n1278), .B(n1279), .Z(swire[113]) );
  XOR U2792 ( .A(n1201), .B(n1280), .Z(n1279) );
  XOR U2793 ( .A(n1200), .B(n1278), .Z(n1280) );
  NANDN U2794 ( .A(n179), .B(a[113]), .Z(n1200) );
  XNOR U2795 ( .A(n1271), .B(n1272), .Z(n1201) );
  XOR U2796 ( .A(n1269), .B(n1281), .Z(n1272) );
  NAND U2797 ( .A(b[1]), .B(a[112]), .Z(n1281) );
  XOR U2798 ( .A(n1277), .B(n1282), .Z(n1271) );
  XOR U2799 ( .A(n1269), .B(n1276), .Z(n1282) );
  XNOR U2800 ( .A(n1283), .B(n1275), .Z(n1276) );
  AND U2801 ( .A(b[2]), .B(a[111]), .Z(n1283) );
  NANDN U2802 ( .A(n1284), .B(n1285), .Z(n1269) );
  XOR U2803 ( .A(n1275), .B(n1267), .Z(n1286) );
  XNOR U2804 ( .A(n1266), .B(n1262), .Z(n1287) );
  XNOR U2805 ( .A(n1261), .B(n1257), .Z(n1288) );
  XNOR U2806 ( .A(n1256), .B(n1252), .Z(n1289) );
  XNOR U2807 ( .A(n1251), .B(n1247), .Z(n1290) );
  XNOR U2808 ( .A(n1246), .B(n1242), .Z(n1291) );
  XNOR U2809 ( .A(n1241), .B(n1237), .Z(n1292) );
  XNOR U2810 ( .A(n1236), .B(n1232), .Z(n1293) );
  XNOR U2811 ( .A(n1231), .B(n1227), .Z(n1294) );
  XOR U2812 ( .A(n1226), .B(n1223), .Z(n1295) );
  XOR U2813 ( .A(n1296), .B(n1297), .Z(n1223) );
  XOR U2814 ( .A(n1221), .B(n1298), .Z(n1297) );
  XOR U2815 ( .A(n1299), .B(n1300), .Z(n1298) );
  XOR U2816 ( .A(n1301), .B(n1302), .Z(n1300) );
  NAND U2817 ( .A(b[14]), .B(a[99]), .Z(n1302) );
  AND U2818 ( .A(b[15]), .B(a[98]), .Z(n1301) );
  XOR U2819 ( .A(n1303), .B(n1299), .Z(n1296) );
  XOR U2820 ( .A(n1304), .B(n1305), .Z(n1299) );
  NOR U2821 ( .A(n1306), .B(n1307), .Z(n1304) );
  AND U2822 ( .A(b[13]), .B(a[100]), .Z(n1303) );
  XNOR U2823 ( .A(n1308), .B(n1221), .Z(n1222) );
  XOR U2824 ( .A(n1309), .B(n1310), .Z(n1221) );
  ANDN U2825 ( .B(n1311), .A(n1312), .Z(n1309) );
  AND U2826 ( .A(b[12]), .B(a[101]), .Z(n1308) );
  XNOR U2827 ( .A(n1313), .B(n1226), .Z(n1228) );
  XOR U2828 ( .A(n1314), .B(n1315), .Z(n1226) );
  ANDN U2829 ( .B(n1316), .A(n1317), .Z(n1314) );
  AND U2830 ( .A(b[11]), .B(a[102]), .Z(n1313) );
  XNOR U2831 ( .A(n1318), .B(n1231), .Z(n1233) );
  XOR U2832 ( .A(n1319), .B(n1320), .Z(n1231) );
  ANDN U2833 ( .B(n1321), .A(n1322), .Z(n1319) );
  AND U2834 ( .A(b[10]), .B(a[103]), .Z(n1318) );
  XNOR U2835 ( .A(n1323), .B(n1236), .Z(n1238) );
  XOR U2836 ( .A(n1324), .B(n1325), .Z(n1236) );
  ANDN U2837 ( .B(n1326), .A(n1327), .Z(n1324) );
  AND U2838 ( .A(b[9]), .B(a[104]), .Z(n1323) );
  XNOR U2839 ( .A(n1328), .B(n1241), .Z(n1243) );
  XOR U2840 ( .A(n1329), .B(n1330), .Z(n1241) );
  ANDN U2841 ( .B(n1331), .A(n1332), .Z(n1329) );
  AND U2842 ( .A(b[8]), .B(a[105]), .Z(n1328) );
  XNOR U2843 ( .A(n1333), .B(n1246), .Z(n1248) );
  XOR U2844 ( .A(n1334), .B(n1335), .Z(n1246) );
  ANDN U2845 ( .B(n1336), .A(n1337), .Z(n1334) );
  AND U2846 ( .A(b[7]), .B(a[106]), .Z(n1333) );
  XNOR U2847 ( .A(n1338), .B(n1251), .Z(n1253) );
  XOR U2848 ( .A(n1339), .B(n1340), .Z(n1251) );
  ANDN U2849 ( .B(n1341), .A(n1342), .Z(n1339) );
  AND U2850 ( .A(b[6]), .B(a[107]), .Z(n1338) );
  XNOR U2851 ( .A(n1343), .B(n1256), .Z(n1258) );
  XOR U2852 ( .A(n1344), .B(n1345), .Z(n1256) );
  ANDN U2853 ( .B(n1346), .A(n1347), .Z(n1344) );
  AND U2854 ( .A(b[5]), .B(a[108]), .Z(n1343) );
  XNOR U2855 ( .A(n1348), .B(n1261), .Z(n1263) );
  XOR U2856 ( .A(n1349), .B(n1350), .Z(n1261) );
  ANDN U2857 ( .B(n1351), .A(n1352), .Z(n1349) );
  AND U2858 ( .A(b[4]), .B(a[109]), .Z(n1348) );
  XNOR U2859 ( .A(n1353), .B(n1354), .Z(n1275) );
  NANDN U2860 ( .A(n1355), .B(n1356), .Z(n1354) );
  XNOR U2861 ( .A(n1357), .B(n1266), .Z(n1268) );
  XNOR U2862 ( .A(n1358), .B(n1359), .Z(n1266) );
  AND U2863 ( .A(n1360), .B(n1361), .Z(n1358) );
  AND U2864 ( .A(b[3]), .B(a[110]), .Z(n1357) );
  XNOR U2865 ( .A(n1362), .B(n1363), .Z(swire[112]) );
  XOR U2866 ( .A(n1285), .B(n1365), .Z(n1363) );
  XNOR U2867 ( .A(n1284), .B(n1364), .Z(n1365) );
  IV U2868 ( .A(n1362), .Z(n1364) );
  NANDN U2869 ( .A(n179), .B(a[112]), .Z(n1284) );
  XNOR U2870 ( .A(n1355), .B(n1356), .Z(n1285) );
  XOR U2871 ( .A(n1353), .B(n1366), .Z(n1356) );
  NAND U2872 ( .A(b[1]), .B(a[111]), .Z(n1366) );
  XOR U2873 ( .A(n1361), .B(n1367), .Z(n1355) );
  XOR U2874 ( .A(n1353), .B(n1360), .Z(n1367) );
  XNOR U2875 ( .A(n1368), .B(n1359), .Z(n1360) );
  AND U2876 ( .A(b[2]), .B(a[110]), .Z(n1368) );
  NANDN U2877 ( .A(n1369), .B(n1370), .Z(n1353) );
  XOR U2878 ( .A(n1359), .B(n1351), .Z(n1371) );
  XNOR U2879 ( .A(n1350), .B(n1346), .Z(n1372) );
  XNOR U2880 ( .A(n1345), .B(n1341), .Z(n1373) );
  XNOR U2881 ( .A(n1340), .B(n1336), .Z(n1374) );
  XNOR U2882 ( .A(n1335), .B(n1331), .Z(n1375) );
  XNOR U2883 ( .A(n1330), .B(n1326), .Z(n1376) );
  XNOR U2884 ( .A(n1325), .B(n1321), .Z(n1377) );
  XNOR U2885 ( .A(n1320), .B(n1316), .Z(n1378) );
  XNOR U2886 ( .A(n1315), .B(n1311), .Z(n1379) );
  XOR U2887 ( .A(n1310), .B(n1307), .Z(n1380) );
  XOR U2888 ( .A(n1381), .B(n1382), .Z(n1307) );
  XOR U2889 ( .A(n1305), .B(n1383), .Z(n1382) );
  XOR U2890 ( .A(n1384), .B(n1385), .Z(n1383) );
  XOR U2891 ( .A(n1386), .B(n1387), .Z(n1385) );
  NAND U2892 ( .A(b[14]), .B(a[98]), .Z(n1387) );
  AND U2893 ( .A(a[97]), .B(b[15]), .Z(n1386) );
  XOR U2894 ( .A(n1388), .B(n1384), .Z(n1381) );
  XOR U2895 ( .A(n1389), .B(n1390), .Z(n1384) );
  NOR U2896 ( .A(n1391), .B(n1392), .Z(n1389) );
  AND U2897 ( .A(b[13]), .B(a[99]), .Z(n1388) );
  XNOR U2898 ( .A(n1393), .B(n1305), .Z(n1306) );
  XOR U2899 ( .A(n1394), .B(n1395), .Z(n1305) );
  ANDN U2900 ( .B(n1396), .A(n1397), .Z(n1394) );
  AND U2901 ( .A(b[12]), .B(a[100]), .Z(n1393) );
  XNOR U2902 ( .A(n1398), .B(n1310), .Z(n1312) );
  XOR U2903 ( .A(n1399), .B(n1400), .Z(n1310) );
  ANDN U2904 ( .B(n1401), .A(n1402), .Z(n1399) );
  AND U2905 ( .A(b[11]), .B(a[101]), .Z(n1398) );
  XNOR U2906 ( .A(n1403), .B(n1315), .Z(n1317) );
  XOR U2907 ( .A(n1404), .B(n1405), .Z(n1315) );
  ANDN U2908 ( .B(n1406), .A(n1407), .Z(n1404) );
  AND U2909 ( .A(b[10]), .B(a[102]), .Z(n1403) );
  XNOR U2910 ( .A(n1408), .B(n1320), .Z(n1322) );
  XOR U2911 ( .A(n1409), .B(n1410), .Z(n1320) );
  ANDN U2912 ( .B(n1411), .A(n1412), .Z(n1409) );
  AND U2913 ( .A(b[9]), .B(a[103]), .Z(n1408) );
  XNOR U2914 ( .A(n1413), .B(n1325), .Z(n1327) );
  XOR U2915 ( .A(n1414), .B(n1415), .Z(n1325) );
  ANDN U2916 ( .B(n1416), .A(n1417), .Z(n1414) );
  AND U2917 ( .A(b[8]), .B(a[104]), .Z(n1413) );
  XNOR U2918 ( .A(n1418), .B(n1330), .Z(n1332) );
  XOR U2919 ( .A(n1419), .B(n1420), .Z(n1330) );
  ANDN U2920 ( .B(n1421), .A(n1422), .Z(n1419) );
  AND U2921 ( .A(b[7]), .B(a[105]), .Z(n1418) );
  XNOR U2922 ( .A(n1423), .B(n1335), .Z(n1337) );
  XOR U2923 ( .A(n1424), .B(n1425), .Z(n1335) );
  ANDN U2924 ( .B(n1426), .A(n1427), .Z(n1424) );
  AND U2925 ( .A(b[6]), .B(a[106]), .Z(n1423) );
  XNOR U2926 ( .A(n1428), .B(n1340), .Z(n1342) );
  XOR U2927 ( .A(n1429), .B(n1430), .Z(n1340) );
  ANDN U2928 ( .B(n1431), .A(n1432), .Z(n1429) );
  AND U2929 ( .A(b[5]), .B(a[107]), .Z(n1428) );
  XNOR U2930 ( .A(n1433), .B(n1345), .Z(n1347) );
  XOR U2931 ( .A(n1434), .B(n1435), .Z(n1345) );
  ANDN U2932 ( .B(n1436), .A(n1437), .Z(n1434) );
  AND U2933 ( .A(b[4]), .B(a[108]), .Z(n1433) );
  XNOR U2934 ( .A(n1438), .B(n1439), .Z(n1359) );
  NANDN U2935 ( .A(n1440), .B(n1441), .Z(n1439) );
  XNOR U2936 ( .A(n1442), .B(n1350), .Z(n1352) );
  XNOR U2937 ( .A(n1443), .B(n1444), .Z(n1350) );
  AND U2938 ( .A(n1445), .B(n1446), .Z(n1443) );
  AND U2939 ( .A(b[3]), .B(a[109]), .Z(n1442) );
  XNOR U2940 ( .A(n1447), .B(n1448), .Z(n1362) );
  NOR U2941 ( .A(n1449), .B(n1450), .Z(n1447) );
  XOR U2942 ( .A(n1450), .B(n1449), .Z(swire[111]) );
  XOR U2943 ( .A(sreg[239]), .B(n1448), .Z(n1449) );
  XOR U2944 ( .A(n1370), .B(n1451), .Z(n1450) );
  XNOR U2945 ( .A(n1369), .B(n1448), .Z(n1451) );
  XOR U2946 ( .A(n1452), .B(n1453), .Z(n1448) );
  NOR U2947 ( .A(n1454), .B(n1455), .Z(n1452) );
  NANDN U2948 ( .A(n179), .B(a[111]), .Z(n1369) );
  XNOR U2949 ( .A(n1440), .B(n1441), .Z(n1370) );
  XOR U2950 ( .A(n1438), .B(n1456), .Z(n1441) );
  NAND U2951 ( .A(b[1]), .B(a[110]), .Z(n1456) );
  XOR U2952 ( .A(n1446), .B(n1457), .Z(n1440) );
  XOR U2953 ( .A(n1438), .B(n1445), .Z(n1457) );
  XNOR U2954 ( .A(n1458), .B(n1444), .Z(n1445) );
  AND U2955 ( .A(b[2]), .B(a[109]), .Z(n1458) );
  NANDN U2956 ( .A(n1459), .B(n1460), .Z(n1438) );
  XOR U2957 ( .A(n1444), .B(n1436), .Z(n1461) );
  XNOR U2958 ( .A(n1435), .B(n1431), .Z(n1462) );
  XNOR U2959 ( .A(n1430), .B(n1426), .Z(n1463) );
  XNOR U2960 ( .A(n1425), .B(n1421), .Z(n1464) );
  XNOR U2961 ( .A(n1420), .B(n1416), .Z(n1465) );
  XNOR U2962 ( .A(n1415), .B(n1411), .Z(n1466) );
  XNOR U2963 ( .A(n1410), .B(n1406), .Z(n1467) );
  XNOR U2964 ( .A(n1405), .B(n1401), .Z(n1468) );
  XNOR U2965 ( .A(n1400), .B(n1396), .Z(n1469) );
  XOR U2966 ( .A(n1395), .B(n1392), .Z(n1470) );
  XOR U2967 ( .A(n1471), .B(n1472), .Z(n1392) );
  XOR U2968 ( .A(n1390), .B(n1473), .Z(n1472) );
  XOR U2969 ( .A(n1474), .B(n1475), .Z(n1473) );
  XOR U2970 ( .A(n1476), .B(n1477), .Z(n1475) );
  NAND U2971 ( .A(a[97]), .B(b[14]), .Z(n1477) );
  AND U2972 ( .A(a[96]), .B(b[15]), .Z(n1476) );
  XOR U2973 ( .A(n1478), .B(n1474), .Z(n1471) );
  XOR U2974 ( .A(n1479), .B(n1480), .Z(n1474) );
  NOR U2975 ( .A(n1481), .B(n1482), .Z(n1479) );
  AND U2976 ( .A(b[13]), .B(a[98]), .Z(n1478) );
  XNOR U2977 ( .A(n1483), .B(n1390), .Z(n1391) );
  XOR U2978 ( .A(n1484), .B(n1485), .Z(n1390) );
  ANDN U2979 ( .B(n1486), .A(n1487), .Z(n1484) );
  AND U2980 ( .A(b[12]), .B(a[99]), .Z(n1483) );
  XNOR U2981 ( .A(n1488), .B(n1395), .Z(n1397) );
  XOR U2982 ( .A(n1489), .B(n1490), .Z(n1395) );
  ANDN U2983 ( .B(n1491), .A(n1492), .Z(n1489) );
  AND U2984 ( .A(b[11]), .B(a[100]), .Z(n1488) );
  XNOR U2985 ( .A(n1493), .B(n1400), .Z(n1402) );
  XOR U2986 ( .A(n1494), .B(n1495), .Z(n1400) );
  ANDN U2987 ( .B(n1496), .A(n1497), .Z(n1494) );
  AND U2988 ( .A(b[10]), .B(a[101]), .Z(n1493) );
  XNOR U2989 ( .A(n1498), .B(n1405), .Z(n1407) );
  XOR U2990 ( .A(n1499), .B(n1500), .Z(n1405) );
  ANDN U2991 ( .B(n1501), .A(n1502), .Z(n1499) );
  AND U2992 ( .A(b[9]), .B(a[102]), .Z(n1498) );
  XNOR U2993 ( .A(n1503), .B(n1410), .Z(n1412) );
  XOR U2994 ( .A(n1504), .B(n1505), .Z(n1410) );
  ANDN U2995 ( .B(n1506), .A(n1507), .Z(n1504) );
  AND U2996 ( .A(b[8]), .B(a[103]), .Z(n1503) );
  XNOR U2997 ( .A(n1508), .B(n1415), .Z(n1417) );
  XOR U2998 ( .A(n1509), .B(n1510), .Z(n1415) );
  ANDN U2999 ( .B(n1511), .A(n1512), .Z(n1509) );
  AND U3000 ( .A(b[7]), .B(a[104]), .Z(n1508) );
  XNOR U3001 ( .A(n1513), .B(n1420), .Z(n1422) );
  XOR U3002 ( .A(n1514), .B(n1515), .Z(n1420) );
  ANDN U3003 ( .B(n1516), .A(n1517), .Z(n1514) );
  AND U3004 ( .A(b[6]), .B(a[105]), .Z(n1513) );
  XNOR U3005 ( .A(n1518), .B(n1425), .Z(n1427) );
  XOR U3006 ( .A(n1519), .B(n1520), .Z(n1425) );
  ANDN U3007 ( .B(n1521), .A(n1522), .Z(n1519) );
  AND U3008 ( .A(b[5]), .B(a[106]), .Z(n1518) );
  XNOR U3009 ( .A(n1523), .B(n1430), .Z(n1432) );
  XOR U3010 ( .A(n1524), .B(n1525), .Z(n1430) );
  ANDN U3011 ( .B(n1526), .A(n1527), .Z(n1524) );
  AND U3012 ( .A(b[4]), .B(a[107]), .Z(n1523) );
  XNOR U3013 ( .A(n1528), .B(n1529), .Z(n1444) );
  NANDN U3014 ( .A(n1530), .B(n1531), .Z(n1529) );
  XNOR U3015 ( .A(n1532), .B(n1435), .Z(n1437) );
  XNOR U3016 ( .A(n1533), .B(n1534), .Z(n1435) );
  AND U3017 ( .A(n1535), .B(n1536), .Z(n1533) );
  AND U3018 ( .A(b[3]), .B(a[108]), .Z(n1532) );
  XOR U3019 ( .A(n1455), .B(n1454), .Z(swire[110]) );
  XOR U3020 ( .A(sreg[238]), .B(n1453), .Z(n1454) );
  XOR U3021 ( .A(n1460), .B(n1537), .Z(n1455) );
  XNOR U3022 ( .A(n1459), .B(n1453), .Z(n1537) );
  XOR U3023 ( .A(n1538), .B(n1539), .Z(n1453) );
  NOR U3024 ( .A(n1540), .B(n1541), .Z(n1538) );
  NANDN U3025 ( .A(n179), .B(a[110]), .Z(n1459) );
  XNOR U3026 ( .A(n1530), .B(n1531), .Z(n1460) );
  XOR U3027 ( .A(n1528), .B(n1542), .Z(n1531) );
  NAND U3028 ( .A(b[1]), .B(a[109]), .Z(n1542) );
  XOR U3029 ( .A(n1536), .B(n1543), .Z(n1530) );
  XOR U3030 ( .A(n1528), .B(n1535), .Z(n1543) );
  XNOR U3031 ( .A(n1544), .B(n1534), .Z(n1535) );
  AND U3032 ( .A(b[2]), .B(a[108]), .Z(n1544) );
  NANDN U3033 ( .A(n1545), .B(n1546), .Z(n1528) );
  XOR U3034 ( .A(n1534), .B(n1526), .Z(n1547) );
  XNOR U3035 ( .A(n1525), .B(n1521), .Z(n1548) );
  XNOR U3036 ( .A(n1520), .B(n1516), .Z(n1549) );
  XNOR U3037 ( .A(n1515), .B(n1511), .Z(n1550) );
  XNOR U3038 ( .A(n1510), .B(n1506), .Z(n1551) );
  XNOR U3039 ( .A(n1505), .B(n1501), .Z(n1552) );
  XNOR U3040 ( .A(n1500), .B(n1496), .Z(n1553) );
  XNOR U3041 ( .A(n1495), .B(n1491), .Z(n1554) );
  XNOR U3042 ( .A(n1490), .B(n1486), .Z(n1555) );
  XOR U3043 ( .A(n1485), .B(n1482), .Z(n1556) );
  XOR U3044 ( .A(n1557), .B(n1558), .Z(n1482) );
  XOR U3045 ( .A(n1480), .B(n1559), .Z(n1558) );
  XOR U3046 ( .A(n1560), .B(n1561), .Z(n1559) );
  XOR U3047 ( .A(n1562), .B(n1563), .Z(n1561) );
  NAND U3048 ( .A(a[96]), .B(b[14]), .Z(n1563) );
  AND U3049 ( .A(a[95]), .B(b[15]), .Z(n1562) );
  XOR U3050 ( .A(n1564), .B(n1560), .Z(n1557) );
  XOR U3051 ( .A(n1565), .B(n1566), .Z(n1560) );
  NOR U3052 ( .A(n1567), .B(n1568), .Z(n1565) );
  AND U3053 ( .A(a[97]), .B(b[13]), .Z(n1564) );
  XNOR U3054 ( .A(n1569), .B(n1480), .Z(n1481) );
  XOR U3055 ( .A(n1570), .B(n1571), .Z(n1480) );
  ANDN U3056 ( .B(n1572), .A(n1573), .Z(n1570) );
  AND U3057 ( .A(b[12]), .B(a[98]), .Z(n1569) );
  XNOR U3058 ( .A(n1574), .B(n1485), .Z(n1487) );
  XOR U3059 ( .A(n1575), .B(n1576), .Z(n1485) );
  ANDN U3060 ( .B(n1577), .A(n1578), .Z(n1575) );
  AND U3061 ( .A(b[11]), .B(a[99]), .Z(n1574) );
  XNOR U3062 ( .A(n1579), .B(n1490), .Z(n1492) );
  XOR U3063 ( .A(n1580), .B(n1581), .Z(n1490) );
  ANDN U3064 ( .B(n1582), .A(n1583), .Z(n1580) );
  AND U3065 ( .A(b[10]), .B(a[100]), .Z(n1579) );
  XNOR U3066 ( .A(n1584), .B(n1495), .Z(n1497) );
  XOR U3067 ( .A(n1585), .B(n1586), .Z(n1495) );
  ANDN U3068 ( .B(n1587), .A(n1588), .Z(n1585) );
  AND U3069 ( .A(b[9]), .B(a[101]), .Z(n1584) );
  XNOR U3070 ( .A(n1589), .B(n1500), .Z(n1502) );
  XOR U3071 ( .A(n1590), .B(n1591), .Z(n1500) );
  ANDN U3072 ( .B(n1592), .A(n1593), .Z(n1590) );
  AND U3073 ( .A(b[8]), .B(a[102]), .Z(n1589) );
  XNOR U3074 ( .A(n1594), .B(n1505), .Z(n1507) );
  XOR U3075 ( .A(n1595), .B(n1596), .Z(n1505) );
  ANDN U3076 ( .B(n1597), .A(n1598), .Z(n1595) );
  AND U3077 ( .A(b[7]), .B(a[103]), .Z(n1594) );
  XNOR U3078 ( .A(n1599), .B(n1510), .Z(n1512) );
  XOR U3079 ( .A(n1600), .B(n1601), .Z(n1510) );
  ANDN U3080 ( .B(n1602), .A(n1603), .Z(n1600) );
  AND U3081 ( .A(b[6]), .B(a[104]), .Z(n1599) );
  XNOR U3082 ( .A(n1604), .B(n1515), .Z(n1517) );
  XOR U3083 ( .A(n1605), .B(n1606), .Z(n1515) );
  ANDN U3084 ( .B(n1607), .A(n1608), .Z(n1605) );
  AND U3085 ( .A(b[5]), .B(a[105]), .Z(n1604) );
  XNOR U3086 ( .A(n1609), .B(n1520), .Z(n1522) );
  XOR U3087 ( .A(n1610), .B(n1611), .Z(n1520) );
  ANDN U3088 ( .B(n1612), .A(n1613), .Z(n1610) );
  AND U3089 ( .A(b[4]), .B(a[106]), .Z(n1609) );
  XNOR U3090 ( .A(n1614), .B(n1615), .Z(n1534) );
  NANDN U3091 ( .A(n1616), .B(n1617), .Z(n1615) );
  XNOR U3092 ( .A(n1618), .B(n1525), .Z(n1527) );
  XNOR U3093 ( .A(n1619), .B(n1620), .Z(n1525) );
  AND U3094 ( .A(n1621), .B(n1622), .Z(n1619) );
  AND U3095 ( .A(b[3]), .B(a[107]), .Z(n1618) );
  XOR U3096 ( .A(n1541), .B(n1540), .Z(swire[109]) );
  XOR U3097 ( .A(sreg[237]), .B(n1539), .Z(n1540) );
  XOR U3098 ( .A(n1546), .B(n1623), .Z(n1541) );
  XNOR U3099 ( .A(n1545), .B(n1539), .Z(n1623) );
  XOR U3100 ( .A(n1624), .B(n1625), .Z(n1539) );
  NOR U3101 ( .A(n1626), .B(n1627), .Z(n1624) );
  NANDN U3102 ( .A(n179), .B(a[109]), .Z(n1545) );
  XNOR U3103 ( .A(n1616), .B(n1617), .Z(n1546) );
  XOR U3104 ( .A(n1614), .B(n1628), .Z(n1617) );
  NAND U3105 ( .A(b[1]), .B(a[108]), .Z(n1628) );
  XOR U3106 ( .A(n1622), .B(n1629), .Z(n1616) );
  XOR U3107 ( .A(n1614), .B(n1621), .Z(n1629) );
  XNOR U3108 ( .A(n1630), .B(n1620), .Z(n1621) );
  AND U3109 ( .A(b[2]), .B(a[107]), .Z(n1630) );
  NANDN U3110 ( .A(n1631), .B(n1632), .Z(n1614) );
  XOR U3111 ( .A(n1620), .B(n1612), .Z(n1633) );
  XNOR U3112 ( .A(n1611), .B(n1607), .Z(n1634) );
  XNOR U3113 ( .A(n1606), .B(n1602), .Z(n1635) );
  XNOR U3114 ( .A(n1601), .B(n1597), .Z(n1636) );
  XNOR U3115 ( .A(n1596), .B(n1592), .Z(n1637) );
  XNOR U3116 ( .A(n1591), .B(n1587), .Z(n1638) );
  XNOR U3117 ( .A(n1586), .B(n1582), .Z(n1639) );
  XNOR U3118 ( .A(n1581), .B(n1577), .Z(n1640) );
  XNOR U3119 ( .A(n1576), .B(n1572), .Z(n1641) );
  XOR U3120 ( .A(n1571), .B(n1568), .Z(n1642) );
  XOR U3121 ( .A(n1643), .B(n1644), .Z(n1568) );
  XOR U3122 ( .A(n1566), .B(n1645), .Z(n1644) );
  XOR U3123 ( .A(n1646), .B(n1647), .Z(n1645) );
  XOR U3124 ( .A(n1648), .B(n1649), .Z(n1647) );
  NAND U3125 ( .A(a[95]), .B(b[14]), .Z(n1649) );
  AND U3126 ( .A(a[94]), .B(b[15]), .Z(n1648) );
  XOR U3127 ( .A(n1650), .B(n1646), .Z(n1643) );
  XOR U3128 ( .A(n1651), .B(n1652), .Z(n1646) );
  NOR U3129 ( .A(n1653), .B(n1654), .Z(n1651) );
  AND U3130 ( .A(a[96]), .B(b[13]), .Z(n1650) );
  XNOR U3131 ( .A(n1655), .B(n1566), .Z(n1567) );
  XOR U3132 ( .A(n1656), .B(n1657), .Z(n1566) );
  ANDN U3133 ( .B(n1658), .A(n1659), .Z(n1656) );
  AND U3134 ( .A(a[97]), .B(b[12]), .Z(n1655) );
  XNOR U3135 ( .A(n1660), .B(n1571), .Z(n1573) );
  XOR U3136 ( .A(n1661), .B(n1662), .Z(n1571) );
  ANDN U3137 ( .B(n1663), .A(n1664), .Z(n1661) );
  AND U3138 ( .A(b[11]), .B(a[98]), .Z(n1660) );
  XNOR U3139 ( .A(n1665), .B(n1576), .Z(n1578) );
  XOR U3140 ( .A(n1666), .B(n1667), .Z(n1576) );
  ANDN U3141 ( .B(n1668), .A(n1669), .Z(n1666) );
  AND U3142 ( .A(b[10]), .B(a[99]), .Z(n1665) );
  XNOR U3143 ( .A(n1670), .B(n1581), .Z(n1583) );
  XOR U3144 ( .A(n1671), .B(n1672), .Z(n1581) );
  ANDN U3145 ( .B(n1673), .A(n1674), .Z(n1671) );
  AND U3146 ( .A(b[9]), .B(a[100]), .Z(n1670) );
  XNOR U3147 ( .A(n1675), .B(n1586), .Z(n1588) );
  XOR U3148 ( .A(n1676), .B(n1677), .Z(n1586) );
  ANDN U3149 ( .B(n1678), .A(n1679), .Z(n1676) );
  AND U3150 ( .A(b[8]), .B(a[101]), .Z(n1675) );
  XNOR U3151 ( .A(n1680), .B(n1591), .Z(n1593) );
  XOR U3152 ( .A(n1681), .B(n1682), .Z(n1591) );
  ANDN U3153 ( .B(n1683), .A(n1684), .Z(n1681) );
  AND U3154 ( .A(b[7]), .B(a[102]), .Z(n1680) );
  XNOR U3155 ( .A(n1685), .B(n1596), .Z(n1598) );
  XOR U3156 ( .A(n1686), .B(n1687), .Z(n1596) );
  ANDN U3157 ( .B(n1688), .A(n1689), .Z(n1686) );
  AND U3158 ( .A(b[6]), .B(a[103]), .Z(n1685) );
  XNOR U3159 ( .A(n1690), .B(n1601), .Z(n1603) );
  XOR U3160 ( .A(n1691), .B(n1692), .Z(n1601) );
  ANDN U3161 ( .B(n1693), .A(n1694), .Z(n1691) );
  AND U3162 ( .A(b[5]), .B(a[104]), .Z(n1690) );
  XNOR U3163 ( .A(n1695), .B(n1606), .Z(n1608) );
  XOR U3164 ( .A(n1696), .B(n1697), .Z(n1606) );
  ANDN U3165 ( .B(n1698), .A(n1699), .Z(n1696) );
  AND U3166 ( .A(b[4]), .B(a[105]), .Z(n1695) );
  XNOR U3167 ( .A(n1700), .B(n1701), .Z(n1620) );
  NANDN U3168 ( .A(n1702), .B(n1703), .Z(n1701) );
  XNOR U3169 ( .A(n1704), .B(n1611), .Z(n1613) );
  XNOR U3170 ( .A(n1705), .B(n1706), .Z(n1611) );
  AND U3171 ( .A(n1707), .B(n1708), .Z(n1705) );
  AND U3172 ( .A(b[3]), .B(a[106]), .Z(n1704) );
  XOR U3173 ( .A(n1627), .B(n1626), .Z(swire[108]) );
  XOR U3174 ( .A(sreg[236]), .B(n1625), .Z(n1626) );
  XOR U3175 ( .A(n1632), .B(n1709), .Z(n1627) );
  XNOR U3176 ( .A(n1631), .B(n1625), .Z(n1709) );
  XOR U3177 ( .A(n1710), .B(n1711), .Z(n1625) );
  NOR U3178 ( .A(n1712), .B(n1713), .Z(n1710) );
  NANDN U3179 ( .A(n179), .B(a[108]), .Z(n1631) );
  XNOR U3180 ( .A(n1702), .B(n1703), .Z(n1632) );
  XOR U3181 ( .A(n1700), .B(n1714), .Z(n1703) );
  NAND U3182 ( .A(b[1]), .B(a[107]), .Z(n1714) );
  XOR U3183 ( .A(n1708), .B(n1715), .Z(n1702) );
  XOR U3184 ( .A(n1700), .B(n1707), .Z(n1715) );
  XNOR U3185 ( .A(n1716), .B(n1706), .Z(n1707) );
  AND U3186 ( .A(b[2]), .B(a[106]), .Z(n1716) );
  NANDN U3187 ( .A(n1717), .B(n1718), .Z(n1700) );
  XOR U3188 ( .A(n1706), .B(n1698), .Z(n1719) );
  XNOR U3189 ( .A(n1697), .B(n1693), .Z(n1720) );
  XNOR U3190 ( .A(n1692), .B(n1688), .Z(n1721) );
  XNOR U3191 ( .A(n1687), .B(n1683), .Z(n1722) );
  XNOR U3192 ( .A(n1682), .B(n1678), .Z(n1723) );
  XNOR U3193 ( .A(n1677), .B(n1673), .Z(n1724) );
  XNOR U3194 ( .A(n1672), .B(n1668), .Z(n1725) );
  XNOR U3195 ( .A(n1667), .B(n1663), .Z(n1726) );
  XNOR U3196 ( .A(n1662), .B(n1658), .Z(n1727) );
  XOR U3197 ( .A(n1657), .B(n1654), .Z(n1728) );
  XOR U3198 ( .A(n1729), .B(n1730), .Z(n1654) );
  XOR U3199 ( .A(n1652), .B(n1731), .Z(n1730) );
  XOR U3200 ( .A(n1732), .B(n1733), .Z(n1731) );
  XOR U3201 ( .A(n1734), .B(n1735), .Z(n1733) );
  NAND U3202 ( .A(a[94]), .B(b[14]), .Z(n1735) );
  AND U3203 ( .A(a[93]), .B(b[15]), .Z(n1734) );
  XOR U3204 ( .A(n1736), .B(n1732), .Z(n1729) );
  XOR U3205 ( .A(n1737), .B(n1738), .Z(n1732) );
  NOR U3206 ( .A(n1739), .B(n1740), .Z(n1737) );
  AND U3207 ( .A(a[95]), .B(b[13]), .Z(n1736) );
  XNOR U3208 ( .A(n1741), .B(n1652), .Z(n1653) );
  XOR U3209 ( .A(n1742), .B(n1743), .Z(n1652) );
  ANDN U3210 ( .B(n1744), .A(n1745), .Z(n1742) );
  AND U3211 ( .A(a[96]), .B(b[12]), .Z(n1741) );
  XNOR U3212 ( .A(n1746), .B(n1657), .Z(n1659) );
  XOR U3213 ( .A(n1747), .B(n1748), .Z(n1657) );
  ANDN U3214 ( .B(n1749), .A(n1750), .Z(n1747) );
  AND U3215 ( .A(a[97]), .B(b[11]), .Z(n1746) );
  XNOR U3216 ( .A(n1751), .B(n1662), .Z(n1664) );
  XOR U3217 ( .A(n1752), .B(n1753), .Z(n1662) );
  ANDN U3218 ( .B(n1754), .A(n1755), .Z(n1752) );
  AND U3219 ( .A(b[10]), .B(a[98]), .Z(n1751) );
  XNOR U3220 ( .A(n1756), .B(n1667), .Z(n1669) );
  XOR U3221 ( .A(n1757), .B(n1758), .Z(n1667) );
  ANDN U3222 ( .B(n1759), .A(n1760), .Z(n1757) );
  AND U3223 ( .A(b[9]), .B(a[99]), .Z(n1756) );
  XNOR U3224 ( .A(n1761), .B(n1672), .Z(n1674) );
  XOR U3225 ( .A(n1762), .B(n1763), .Z(n1672) );
  ANDN U3226 ( .B(n1764), .A(n1765), .Z(n1762) );
  AND U3227 ( .A(b[8]), .B(a[100]), .Z(n1761) );
  XNOR U3228 ( .A(n1766), .B(n1677), .Z(n1679) );
  XOR U3229 ( .A(n1767), .B(n1768), .Z(n1677) );
  ANDN U3230 ( .B(n1769), .A(n1770), .Z(n1767) );
  AND U3231 ( .A(b[7]), .B(a[101]), .Z(n1766) );
  XNOR U3232 ( .A(n1771), .B(n1682), .Z(n1684) );
  XOR U3233 ( .A(n1772), .B(n1773), .Z(n1682) );
  ANDN U3234 ( .B(n1774), .A(n1775), .Z(n1772) );
  AND U3235 ( .A(b[6]), .B(a[102]), .Z(n1771) );
  XNOR U3236 ( .A(n1776), .B(n1687), .Z(n1689) );
  XOR U3237 ( .A(n1777), .B(n1778), .Z(n1687) );
  ANDN U3238 ( .B(n1779), .A(n1780), .Z(n1777) );
  AND U3239 ( .A(b[5]), .B(a[103]), .Z(n1776) );
  XNOR U3240 ( .A(n1781), .B(n1692), .Z(n1694) );
  XOR U3241 ( .A(n1782), .B(n1783), .Z(n1692) );
  ANDN U3242 ( .B(n1784), .A(n1785), .Z(n1782) );
  AND U3243 ( .A(b[4]), .B(a[104]), .Z(n1781) );
  XNOR U3244 ( .A(n1786), .B(n1787), .Z(n1706) );
  NANDN U3245 ( .A(n1788), .B(n1789), .Z(n1787) );
  XNOR U3246 ( .A(n1790), .B(n1697), .Z(n1699) );
  XNOR U3247 ( .A(n1791), .B(n1792), .Z(n1697) );
  AND U3248 ( .A(n1793), .B(n1794), .Z(n1791) );
  AND U3249 ( .A(b[3]), .B(a[105]), .Z(n1790) );
  XOR U3250 ( .A(n1713), .B(n1712), .Z(swire[107]) );
  XOR U3251 ( .A(sreg[235]), .B(n1711), .Z(n1712) );
  XOR U3252 ( .A(n1718), .B(n1795), .Z(n1713) );
  XNOR U3253 ( .A(n1717), .B(n1711), .Z(n1795) );
  XOR U3254 ( .A(n1796), .B(n1797), .Z(n1711) );
  NOR U3255 ( .A(n1798), .B(n1799), .Z(n1796) );
  NANDN U3256 ( .A(n179), .B(a[107]), .Z(n1717) );
  XNOR U3257 ( .A(n1788), .B(n1789), .Z(n1718) );
  XOR U3258 ( .A(n1786), .B(n1800), .Z(n1789) );
  NAND U3259 ( .A(b[1]), .B(a[106]), .Z(n1800) );
  XOR U3260 ( .A(n1794), .B(n1801), .Z(n1788) );
  XOR U3261 ( .A(n1786), .B(n1793), .Z(n1801) );
  XNOR U3262 ( .A(n1802), .B(n1792), .Z(n1793) );
  AND U3263 ( .A(b[2]), .B(a[105]), .Z(n1802) );
  NANDN U3264 ( .A(n1803), .B(n1804), .Z(n1786) );
  XOR U3265 ( .A(n1792), .B(n1784), .Z(n1805) );
  XNOR U3266 ( .A(n1783), .B(n1779), .Z(n1806) );
  XNOR U3267 ( .A(n1778), .B(n1774), .Z(n1807) );
  XNOR U3268 ( .A(n1773), .B(n1769), .Z(n1808) );
  XNOR U3269 ( .A(n1768), .B(n1764), .Z(n1809) );
  XNOR U3270 ( .A(n1763), .B(n1759), .Z(n1810) );
  XNOR U3271 ( .A(n1758), .B(n1754), .Z(n1811) );
  XNOR U3272 ( .A(n1753), .B(n1749), .Z(n1812) );
  XNOR U3273 ( .A(n1748), .B(n1744), .Z(n1813) );
  XOR U3274 ( .A(n1743), .B(n1740), .Z(n1814) );
  XOR U3275 ( .A(n1815), .B(n1816), .Z(n1740) );
  XOR U3276 ( .A(n1738), .B(n1817), .Z(n1816) );
  XOR U3277 ( .A(n1818), .B(n1819), .Z(n1817) );
  XOR U3278 ( .A(n1820), .B(n1821), .Z(n1819) );
  NAND U3279 ( .A(a[93]), .B(b[14]), .Z(n1821) );
  AND U3280 ( .A(a[92]), .B(b[15]), .Z(n1820) );
  XOR U3281 ( .A(n1822), .B(n1818), .Z(n1815) );
  XOR U3282 ( .A(n1823), .B(n1824), .Z(n1818) );
  NOR U3283 ( .A(n1825), .B(n1826), .Z(n1823) );
  AND U3284 ( .A(a[94]), .B(b[13]), .Z(n1822) );
  XNOR U3285 ( .A(n1827), .B(n1738), .Z(n1739) );
  XOR U3286 ( .A(n1828), .B(n1829), .Z(n1738) );
  ANDN U3287 ( .B(n1830), .A(n1831), .Z(n1828) );
  AND U3288 ( .A(a[95]), .B(b[12]), .Z(n1827) );
  XNOR U3289 ( .A(n1832), .B(n1743), .Z(n1745) );
  XOR U3290 ( .A(n1833), .B(n1834), .Z(n1743) );
  ANDN U3291 ( .B(n1835), .A(n1836), .Z(n1833) );
  AND U3292 ( .A(a[96]), .B(b[11]), .Z(n1832) );
  XNOR U3293 ( .A(n1837), .B(n1748), .Z(n1750) );
  XOR U3294 ( .A(n1838), .B(n1839), .Z(n1748) );
  ANDN U3295 ( .B(n1840), .A(n1841), .Z(n1838) );
  AND U3296 ( .A(a[97]), .B(b[10]), .Z(n1837) );
  XNOR U3297 ( .A(n1842), .B(n1753), .Z(n1755) );
  XOR U3298 ( .A(n1843), .B(n1844), .Z(n1753) );
  ANDN U3299 ( .B(n1845), .A(n1846), .Z(n1843) );
  AND U3300 ( .A(b[9]), .B(a[98]), .Z(n1842) );
  XNOR U3301 ( .A(n1847), .B(n1758), .Z(n1760) );
  XOR U3302 ( .A(n1848), .B(n1849), .Z(n1758) );
  ANDN U3303 ( .B(n1850), .A(n1851), .Z(n1848) );
  AND U3304 ( .A(b[8]), .B(a[99]), .Z(n1847) );
  XNOR U3305 ( .A(n1852), .B(n1763), .Z(n1765) );
  XOR U3306 ( .A(n1853), .B(n1854), .Z(n1763) );
  ANDN U3307 ( .B(n1855), .A(n1856), .Z(n1853) );
  AND U3308 ( .A(b[7]), .B(a[100]), .Z(n1852) );
  XNOR U3309 ( .A(n1857), .B(n1768), .Z(n1770) );
  XOR U3310 ( .A(n1858), .B(n1859), .Z(n1768) );
  ANDN U3311 ( .B(n1860), .A(n1861), .Z(n1858) );
  AND U3312 ( .A(b[6]), .B(a[101]), .Z(n1857) );
  XNOR U3313 ( .A(n1862), .B(n1773), .Z(n1775) );
  XOR U3314 ( .A(n1863), .B(n1864), .Z(n1773) );
  ANDN U3315 ( .B(n1865), .A(n1866), .Z(n1863) );
  AND U3316 ( .A(b[5]), .B(a[102]), .Z(n1862) );
  XNOR U3317 ( .A(n1867), .B(n1778), .Z(n1780) );
  XOR U3318 ( .A(n1868), .B(n1869), .Z(n1778) );
  ANDN U3319 ( .B(n1870), .A(n1871), .Z(n1868) );
  AND U3320 ( .A(b[4]), .B(a[103]), .Z(n1867) );
  XNOR U3321 ( .A(n1872), .B(n1873), .Z(n1792) );
  NANDN U3322 ( .A(n1874), .B(n1875), .Z(n1873) );
  XNOR U3323 ( .A(n1876), .B(n1783), .Z(n1785) );
  XNOR U3324 ( .A(n1877), .B(n1878), .Z(n1783) );
  AND U3325 ( .A(n1879), .B(n1880), .Z(n1877) );
  AND U3326 ( .A(b[3]), .B(a[104]), .Z(n1876) );
  XOR U3327 ( .A(n1799), .B(n1798), .Z(swire[106]) );
  XOR U3328 ( .A(sreg[234]), .B(n1797), .Z(n1798) );
  XOR U3329 ( .A(n1804), .B(n1881), .Z(n1799) );
  XNOR U3330 ( .A(n1803), .B(n1797), .Z(n1881) );
  XOR U3331 ( .A(n1882), .B(n1883), .Z(n1797) );
  NOR U3332 ( .A(n1884), .B(n1885), .Z(n1882) );
  NANDN U3333 ( .A(n179), .B(a[106]), .Z(n1803) );
  XNOR U3334 ( .A(n1874), .B(n1875), .Z(n1804) );
  XOR U3335 ( .A(n1872), .B(n1886), .Z(n1875) );
  NAND U3336 ( .A(b[1]), .B(a[105]), .Z(n1886) );
  XOR U3337 ( .A(n1880), .B(n1887), .Z(n1874) );
  XOR U3338 ( .A(n1872), .B(n1879), .Z(n1887) );
  XNOR U3339 ( .A(n1888), .B(n1878), .Z(n1879) );
  AND U3340 ( .A(b[2]), .B(a[104]), .Z(n1888) );
  NANDN U3341 ( .A(n1889), .B(n1890), .Z(n1872) );
  XOR U3342 ( .A(n1878), .B(n1870), .Z(n1891) );
  XNOR U3343 ( .A(n1869), .B(n1865), .Z(n1892) );
  XNOR U3344 ( .A(n1864), .B(n1860), .Z(n1893) );
  XNOR U3345 ( .A(n1859), .B(n1855), .Z(n1894) );
  XNOR U3346 ( .A(n1854), .B(n1850), .Z(n1895) );
  XNOR U3347 ( .A(n1849), .B(n1845), .Z(n1896) );
  XNOR U3348 ( .A(n1844), .B(n1840), .Z(n1897) );
  XNOR U3349 ( .A(n1839), .B(n1835), .Z(n1898) );
  XNOR U3350 ( .A(n1834), .B(n1830), .Z(n1899) );
  XOR U3351 ( .A(n1829), .B(n1826), .Z(n1900) );
  XOR U3352 ( .A(n1901), .B(n1902), .Z(n1826) );
  XOR U3353 ( .A(n1824), .B(n1903), .Z(n1902) );
  XOR U3354 ( .A(n1904), .B(n1905), .Z(n1903) );
  XOR U3355 ( .A(n1906), .B(n1907), .Z(n1905) );
  NAND U3356 ( .A(a[92]), .B(b[14]), .Z(n1907) );
  AND U3357 ( .A(a[91]), .B(b[15]), .Z(n1906) );
  XOR U3358 ( .A(n1908), .B(n1904), .Z(n1901) );
  XOR U3359 ( .A(n1909), .B(n1910), .Z(n1904) );
  NOR U3360 ( .A(n1911), .B(n1912), .Z(n1909) );
  AND U3361 ( .A(a[93]), .B(b[13]), .Z(n1908) );
  XNOR U3362 ( .A(n1913), .B(n1824), .Z(n1825) );
  XOR U3363 ( .A(n1914), .B(n1915), .Z(n1824) );
  ANDN U3364 ( .B(n1916), .A(n1917), .Z(n1914) );
  AND U3365 ( .A(a[94]), .B(b[12]), .Z(n1913) );
  XNOR U3366 ( .A(n1918), .B(n1829), .Z(n1831) );
  XOR U3367 ( .A(n1919), .B(n1920), .Z(n1829) );
  ANDN U3368 ( .B(n1921), .A(n1922), .Z(n1919) );
  AND U3369 ( .A(a[95]), .B(b[11]), .Z(n1918) );
  XNOR U3370 ( .A(n1923), .B(n1834), .Z(n1836) );
  XOR U3371 ( .A(n1924), .B(n1925), .Z(n1834) );
  ANDN U3372 ( .B(n1926), .A(n1927), .Z(n1924) );
  AND U3373 ( .A(a[96]), .B(b[10]), .Z(n1923) );
  XNOR U3374 ( .A(n1928), .B(n1839), .Z(n1841) );
  XOR U3375 ( .A(n1929), .B(n1930), .Z(n1839) );
  ANDN U3376 ( .B(n1931), .A(n1932), .Z(n1929) );
  AND U3377 ( .A(a[97]), .B(b[9]), .Z(n1928) );
  XNOR U3378 ( .A(n1933), .B(n1844), .Z(n1846) );
  XOR U3379 ( .A(n1934), .B(n1935), .Z(n1844) );
  ANDN U3380 ( .B(n1936), .A(n1937), .Z(n1934) );
  AND U3381 ( .A(b[8]), .B(a[98]), .Z(n1933) );
  XNOR U3382 ( .A(n1938), .B(n1849), .Z(n1851) );
  XOR U3383 ( .A(n1939), .B(n1940), .Z(n1849) );
  ANDN U3384 ( .B(n1941), .A(n1942), .Z(n1939) );
  AND U3385 ( .A(b[7]), .B(a[99]), .Z(n1938) );
  XNOR U3386 ( .A(n1943), .B(n1854), .Z(n1856) );
  XOR U3387 ( .A(n1944), .B(n1945), .Z(n1854) );
  ANDN U3388 ( .B(n1946), .A(n1947), .Z(n1944) );
  AND U3389 ( .A(b[6]), .B(a[100]), .Z(n1943) );
  XNOR U3390 ( .A(n1948), .B(n1859), .Z(n1861) );
  XOR U3391 ( .A(n1949), .B(n1950), .Z(n1859) );
  ANDN U3392 ( .B(n1951), .A(n1952), .Z(n1949) );
  AND U3393 ( .A(b[5]), .B(a[101]), .Z(n1948) );
  XNOR U3394 ( .A(n1953), .B(n1864), .Z(n1866) );
  XOR U3395 ( .A(n1954), .B(n1955), .Z(n1864) );
  ANDN U3396 ( .B(n1956), .A(n1957), .Z(n1954) );
  AND U3397 ( .A(b[4]), .B(a[102]), .Z(n1953) );
  XNOR U3398 ( .A(n1958), .B(n1959), .Z(n1878) );
  NANDN U3399 ( .A(n1960), .B(n1961), .Z(n1959) );
  XNOR U3400 ( .A(n1962), .B(n1869), .Z(n1871) );
  XNOR U3401 ( .A(n1963), .B(n1964), .Z(n1869) );
  AND U3402 ( .A(n1965), .B(n1966), .Z(n1963) );
  AND U3403 ( .A(b[3]), .B(a[103]), .Z(n1962) );
  XOR U3404 ( .A(n1885), .B(n1884), .Z(swire[105]) );
  XOR U3405 ( .A(sreg[233]), .B(n1883), .Z(n1884) );
  XOR U3406 ( .A(n1890), .B(n1967), .Z(n1885) );
  XNOR U3407 ( .A(n1889), .B(n1883), .Z(n1967) );
  XOR U3408 ( .A(n1968), .B(n1969), .Z(n1883) );
  NOR U3409 ( .A(n1970), .B(n1971), .Z(n1968) );
  NANDN U3410 ( .A(n179), .B(a[105]), .Z(n1889) );
  XNOR U3411 ( .A(n1960), .B(n1961), .Z(n1890) );
  XOR U3412 ( .A(n1958), .B(n1972), .Z(n1961) );
  NAND U3413 ( .A(b[1]), .B(a[104]), .Z(n1972) );
  XOR U3414 ( .A(n1966), .B(n1973), .Z(n1960) );
  XOR U3415 ( .A(n1958), .B(n1965), .Z(n1973) );
  XNOR U3416 ( .A(n1974), .B(n1964), .Z(n1965) );
  AND U3417 ( .A(b[2]), .B(a[103]), .Z(n1974) );
  NANDN U3418 ( .A(n1975), .B(n1976), .Z(n1958) );
  XOR U3419 ( .A(n1964), .B(n1956), .Z(n1977) );
  XNOR U3420 ( .A(n1955), .B(n1951), .Z(n1978) );
  XNOR U3421 ( .A(n1950), .B(n1946), .Z(n1979) );
  XNOR U3422 ( .A(n1945), .B(n1941), .Z(n1980) );
  XNOR U3423 ( .A(n1940), .B(n1936), .Z(n1981) );
  XNOR U3424 ( .A(n1935), .B(n1931), .Z(n1982) );
  XNOR U3425 ( .A(n1930), .B(n1926), .Z(n1983) );
  XNOR U3426 ( .A(n1925), .B(n1921), .Z(n1984) );
  XNOR U3427 ( .A(n1920), .B(n1916), .Z(n1985) );
  XOR U3428 ( .A(n1915), .B(n1912), .Z(n1986) );
  XOR U3429 ( .A(n1987), .B(n1988), .Z(n1912) );
  XOR U3430 ( .A(n1910), .B(n1989), .Z(n1988) );
  XOR U3431 ( .A(n1990), .B(n1991), .Z(n1989) );
  XOR U3432 ( .A(n1992), .B(n1993), .Z(n1991) );
  NAND U3433 ( .A(a[91]), .B(b[14]), .Z(n1993) );
  AND U3434 ( .A(a[90]), .B(b[15]), .Z(n1992) );
  XOR U3435 ( .A(n1994), .B(n1990), .Z(n1987) );
  XOR U3436 ( .A(n1995), .B(n1996), .Z(n1990) );
  NOR U3437 ( .A(n1997), .B(n1998), .Z(n1995) );
  AND U3438 ( .A(a[92]), .B(b[13]), .Z(n1994) );
  XNOR U3439 ( .A(n1999), .B(n1910), .Z(n1911) );
  XOR U3440 ( .A(n2000), .B(n2001), .Z(n1910) );
  ANDN U3441 ( .B(n2002), .A(n2003), .Z(n2000) );
  AND U3442 ( .A(a[93]), .B(b[12]), .Z(n1999) );
  XNOR U3443 ( .A(n2004), .B(n1915), .Z(n1917) );
  XOR U3444 ( .A(n2005), .B(n2006), .Z(n1915) );
  ANDN U3445 ( .B(n2007), .A(n2008), .Z(n2005) );
  AND U3446 ( .A(a[94]), .B(b[11]), .Z(n2004) );
  XNOR U3447 ( .A(n2009), .B(n1920), .Z(n1922) );
  XOR U3448 ( .A(n2010), .B(n2011), .Z(n1920) );
  ANDN U3449 ( .B(n2012), .A(n2013), .Z(n2010) );
  AND U3450 ( .A(a[95]), .B(b[10]), .Z(n2009) );
  XNOR U3451 ( .A(n2014), .B(n1925), .Z(n1927) );
  XOR U3452 ( .A(n2015), .B(n2016), .Z(n1925) );
  ANDN U3453 ( .B(n2017), .A(n2018), .Z(n2015) );
  AND U3454 ( .A(a[96]), .B(b[9]), .Z(n2014) );
  XNOR U3455 ( .A(n2019), .B(n1930), .Z(n1932) );
  XOR U3456 ( .A(n2020), .B(n2021), .Z(n1930) );
  ANDN U3457 ( .B(n2022), .A(n2023), .Z(n2020) );
  AND U3458 ( .A(a[97]), .B(b[8]), .Z(n2019) );
  XNOR U3459 ( .A(n2024), .B(n1935), .Z(n1937) );
  XOR U3460 ( .A(n2025), .B(n2026), .Z(n1935) );
  ANDN U3461 ( .B(n2027), .A(n2028), .Z(n2025) );
  AND U3462 ( .A(b[7]), .B(a[98]), .Z(n2024) );
  XNOR U3463 ( .A(n2029), .B(n1940), .Z(n1942) );
  XOR U3464 ( .A(n2030), .B(n2031), .Z(n1940) );
  ANDN U3465 ( .B(n2032), .A(n2033), .Z(n2030) );
  AND U3466 ( .A(b[6]), .B(a[99]), .Z(n2029) );
  XNOR U3467 ( .A(n2034), .B(n1945), .Z(n1947) );
  XOR U3468 ( .A(n2035), .B(n2036), .Z(n1945) );
  ANDN U3469 ( .B(n2037), .A(n2038), .Z(n2035) );
  AND U3470 ( .A(b[5]), .B(a[100]), .Z(n2034) );
  XNOR U3471 ( .A(n2039), .B(n1950), .Z(n1952) );
  XOR U3472 ( .A(n2040), .B(n2041), .Z(n1950) );
  ANDN U3473 ( .B(n2042), .A(n2043), .Z(n2040) );
  AND U3474 ( .A(b[4]), .B(a[101]), .Z(n2039) );
  XNOR U3475 ( .A(n2044), .B(n2045), .Z(n1964) );
  NANDN U3476 ( .A(n2046), .B(n2047), .Z(n2045) );
  XNOR U3477 ( .A(n2048), .B(n1955), .Z(n1957) );
  XNOR U3478 ( .A(n2049), .B(n2050), .Z(n1955) );
  AND U3479 ( .A(n2051), .B(n2052), .Z(n2049) );
  AND U3480 ( .A(b[3]), .B(a[102]), .Z(n2048) );
  XOR U3481 ( .A(n1971), .B(n1970), .Z(swire[104]) );
  XOR U3482 ( .A(sreg[232]), .B(n1969), .Z(n1970) );
  XOR U3483 ( .A(n1976), .B(n2053), .Z(n1971) );
  XNOR U3484 ( .A(n1975), .B(n1969), .Z(n2053) );
  XOR U3485 ( .A(n2054), .B(n2055), .Z(n1969) );
  NOR U3486 ( .A(n2056), .B(n2057), .Z(n2054) );
  NANDN U3487 ( .A(n179), .B(a[104]), .Z(n1975) );
  XNOR U3488 ( .A(n2046), .B(n2047), .Z(n1976) );
  XOR U3489 ( .A(n2044), .B(n2058), .Z(n2047) );
  NAND U3490 ( .A(b[1]), .B(a[103]), .Z(n2058) );
  XOR U3491 ( .A(n2052), .B(n2059), .Z(n2046) );
  XOR U3492 ( .A(n2044), .B(n2051), .Z(n2059) );
  XNOR U3493 ( .A(n2060), .B(n2050), .Z(n2051) );
  AND U3494 ( .A(b[2]), .B(a[102]), .Z(n2060) );
  NANDN U3495 ( .A(n2061), .B(n2062), .Z(n2044) );
  XOR U3496 ( .A(n2050), .B(n2042), .Z(n2063) );
  XNOR U3497 ( .A(n2041), .B(n2037), .Z(n2064) );
  XNOR U3498 ( .A(n2036), .B(n2032), .Z(n2065) );
  XNOR U3499 ( .A(n2031), .B(n2027), .Z(n2066) );
  XNOR U3500 ( .A(n2026), .B(n2022), .Z(n2067) );
  XNOR U3501 ( .A(n2021), .B(n2017), .Z(n2068) );
  XNOR U3502 ( .A(n2016), .B(n2012), .Z(n2069) );
  XNOR U3503 ( .A(n2011), .B(n2007), .Z(n2070) );
  XNOR U3504 ( .A(n2006), .B(n2002), .Z(n2071) );
  XOR U3505 ( .A(n2001), .B(n1998), .Z(n2072) );
  XOR U3506 ( .A(n2073), .B(n2074), .Z(n1998) );
  XOR U3507 ( .A(n1996), .B(n2075), .Z(n2074) );
  XOR U3508 ( .A(n2076), .B(n2077), .Z(n2075) );
  XOR U3509 ( .A(n2078), .B(n2079), .Z(n2077) );
  NAND U3510 ( .A(a[90]), .B(b[14]), .Z(n2079) );
  AND U3511 ( .A(a[89]), .B(b[15]), .Z(n2078) );
  XOR U3512 ( .A(n2080), .B(n2076), .Z(n2073) );
  XOR U3513 ( .A(n2081), .B(n2082), .Z(n2076) );
  NOR U3514 ( .A(n2083), .B(n2084), .Z(n2081) );
  AND U3515 ( .A(a[91]), .B(b[13]), .Z(n2080) );
  XNOR U3516 ( .A(n2085), .B(n1996), .Z(n1997) );
  XOR U3517 ( .A(n2086), .B(n2087), .Z(n1996) );
  ANDN U3518 ( .B(n2088), .A(n2089), .Z(n2086) );
  AND U3519 ( .A(a[92]), .B(b[12]), .Z(n2085) );
  XNOR U3520 ( .A(n2090), .B(n2001), .Z(n2003) );
  XOR U3521 ( .A(n2091), .B(n2092), .Z(n2001) );
  ANDN U3522 ( .B(n2093), .A(n2094), .Z(n2091) );
  AND U3523 ( .A(a[93]), .B(b[11]), .Z(n2090) );
  XNOR U3524 ( .A(n2095), .B(n2006), .Z(n2008) );
  XOR U3525 ( .A(n2096), .B(n2097), .Z(n2006) );
  ANDN U3526 ( .B(n2098), .A(n2099), .Z(n2096) );
  AND U3527 ( .A(a[94]), .B(b[10]), .Z(n2095) );
  XNOR U3528 ( .A(n2100), .B(n2011), .Z(n2013) );
  XOR U3529 ( .A(n2101), .B(n2102), .Z(n2011) );
  ANDN U3530 ( .B(n2103), .A(n2104), .Z(n2101) );
  AND U3531 ( .A(a[95]), .B(b[9]), .Z(n2100) );
  XNOR U3532 ( .A(n2105), .B(n2016), .Z(n2018) );
  XOR U3533 ( .A(n2106), .B(n2107), .Z(n2016) );
  ANDN U3534 ( .B(n2108), .A(n2109), .Z(n2106) );
  AND U3535 ( .A(a[96]), .B(b[8]), .Z(n2105) );
  XNOR U3536 ( .A(n2110), .B(n2021), .Z(n2023) );
  XOR U3537 ( .A(n2111), .B(n2112), .Z(n2021) );
  ANDN U3538 ( .B(n2113), .A(n2114), .Z(n2111) );
  AND U3539 ( .A(a[97]), .B(b[7]), .Z(n2110) );
  XNOR U3540 ( .A(n2115), .B(n2026), .Z(n2028) );
  XOR U3541 ( .A(n2116), .B(n2117), .Z(n2026) );
  ANDN U3542 ( .B(n2118), .A(n2119), .Z(n2116) );
  AND U3543 ( .A(b[6]), .B(a[98]), .Z(n2115) );
  XNOR U3544 ( .A(n2120), .B(n2031), .Z(n2033) );
  XOR U3545 ( .A(n2121), .B(n2122), .Z(n2031) );
  ANDN U3546 ( .B(n2123), .A(n2124), .Z(n2121) );
  AND U3547 ( .A(b[5]), .B(a[99]), .Z(n2120) );
  XNOR U3548 ( .A(n2125), .B(n2036), .Z(n2038) );
  XOR U3549 ( .A(n2126), .B(n2127), .Z(n2036) );
  ANDN U3550 ( .B(n2128), .A(n2129), .Z(n2126) );
  AND U3551 ( .A(b[4]), .B(a[100]), .Z(n2125) );
  XNOR U3552 ( .A(n2130), .B(n2131), .Z(n2050) );
  NANDN U3553 ( .A(n2132), .B(n2133), .Z(n2131) );
  XNOR U3554 ( .A(n2134), .B(n2041), .Z(n2043) );
  XNOR U3555 ( .A(n2135), .B(n2136), .Z(n2041) );
  AND U3556 ( .A(n2137), .B(n2138), .Z(n2135) );
  AND U3557 ( .A(b[3]), .B(a[101]), .Z(n2134) );
  XOR U3558 ( .A(n2057), .B(n2056), .Z(swire[103]) );
  XOR U3559 ( .A(sreg[231]), .B(n2055), .Z(n2056) );
  XOR U3560 ( .A(n2062), .B(n2139), .Z(n2057) );
  XNOR U3561 ( .A(n2061), .B(n2055), .Z(n2139) );
  XOR U3562 ( .A(n2140), .B(n2141), .Z(n2055) );
  NOR U3563 ( .A(n2142), .B(n2143), .Z(n2140) );
  NANDN U3564 ( .A(n179), .B(a[103]), .Z(n2061) );
  XNOR U3565 ( .A(n2132), .B(n2133), .Z(n2062) );
  XOR U3566 ( .A(n2130), .B(n2144), .Z(n2133) );
  NAND U3567 ( .A(b[1]), .B(a[102]), .Z(n2144) );
  XOR U3568 ( .A(n2138), .B(n2145), .Z(n2132) );
  XOR U3569 ( .A(n2130), .B(n2137), .Z(n2145) );
  XNOR U3570 ( .A(n2146), .B(n2136), .Z(n2137) );
  AND U3571 ( .A(b[2]), .B(a[101]), .Z(n2146) );
  NANDN U3572 ( .A(n2147), .B(n2148), .Z(n2130) );
  XOR U3573 ( .A(n2136), .B(n2128), .Z(n2149) );
  XNOR U3574 ( .A(n2127), .B(n2123), .Z(n2150) );
  XNOR U3575 ( .A(n2122), .B(n2118), .Z(n2151) );
  XNOR U3576 ( .A(n2117), .B(n2113), .Z(n2152) );
  XNOR U3577 ( .A(n2112), .B(n2108), .Z(n2153) );
  XNOR U3578 ( .A(n2107), .B(n2103), .Z(n2154) );
  XNOR U3579 ( .A(n2102), .B(n2098), .Z(n2155) );
  XNOR U3580 ( .A(n2097), .B(n2093), .Z(n2156) );
  XNOR U3581 ( .A(n2092), .B(n2088), .Z(n2157) );
  XOR U3582 ( .A(n2087), .B(n2084), .Z(n2158) );
  XOR U3583 ( .A(n2159), .B(n2160), .Z(n2084) );
  XOR U3584 ( .A(n2082), .B(n2161), .Z(n2160) );
  XOR U3585 ( .A(n2162), .B(n2163), .Z(n2161) );
  XOR U3586 ( .A(n2164), .B(n2165), .Z(n2163) );
  NAND U3587 ( .A(a[89]), .B(b[14]), .Z(n2165) );
  AND U3588 ( .A(a[88]), .B(b[15]), .Z(n2164) );
  XOR U3589 ( .A(n2166), .B(n2162), .Z(n2159) );
  XOR U3590 ( .A(n2167), .B(n2168), .Z(n2162) );
  NOR U3591 ( .A(n2169), .B(n2170), .Z(n2167) );
  AND U3592 ( .A(a[90]), .B(b[13]), .Z(n2166) );
  XNOR U3593 ( .A(n2171), .B(n2082), .Z(n2083) );
  XOR U3594 ( .A(n2172), .B(n2173), .Z(n2082) );
  ANDN U3595 ( .B(n2174), .A(n2175), .Z(n2172) );
  AND U3596 ( .A(a[91]), .B(b[12]), .Z(n2171) );
  XNOR U3597 ( .A(n2176), .B(n2087), .Z(n2089) );
  XOR U3598 ( .A(n2177), .B(n2178), .Z(n2087) );
  ANDN U3599 ( .B(n2179), .A(n2180), .Z(n2177) );
  AND U3600 ( .A(a[92]), .B(b[11]), .Z(n2176) );
  XNOR U3601 ( .A(n2181), .B(n2092), .Z(n2094) );
  XOR U3602 ( .A(n2182), .B(n2183), .Z(n2092) );
  ANDN U3603 ( .B(n2184), .A(n2185), .Z(n2182) );
  AND U3604 ( .A(a[93]), .B(b[10]), .Z(n2181) );
  XNOR U3605 ( .A(n2186), .B(n2097), .Z(n2099) );
  XOR U3606 ( .A(n2187), .B(n2188), .Z(n2097) );
  ANDN U3607 ( .B(n2189), .A(n2190), .Z(n2187) );
  AND U3608 ( .A(a[94]), .B(b[9]), .Z(n2186) );
  XNOR U3609 ( .A(n2191), .B(n2102), .Z(n2104) );
  XOR U3610 ( .A(n2192), .B(n2193), .Z(n2102) );
  ANDN U3611 ( .B(n2194), .A(n2195), .Z(n2192) );
  AND U3612 ( .A(a[95]), .B(b[8]), .Z(n2191) );
  XNOR U3613 ( .A(n2196), .B(n2107), .Z(n2109) );
  XOR U3614 ( .A(n2197), .B(n2198), .Z(n2107) );
  ANDN U3615 ( .B(n2199), .A(n2200), .Z(n2197) );
  AND U3616 ( .A(a[96]), .B(b[7]), .Z(n2196) );
  XNOR U3617 ( .A(n2201), .B(n2112), .Z(n2114) );
  XOR U3618 ( .A(n2202), .B(n2203), .Z(n2112) );
  ANDN U3619 ( .B(n2204), .A(n2205), .Z(n2202) );
  AND U3620 ( .A(a[97]), .B(b[6]), .Z(n2201) );
  XNOR U3621 ( .A(n2206), .B(n2117), .Z(n2119) );
  XOR U3622 ( .A(n2207), .B(n2208), .Z(n2117) );
  ANDN U3623 ( .B(n2209), .A(n2210), .Z(n2207) );
  AND U3624 ( .A(b[5]), .B(a[98]), .Z(n2206) );
  XNOR U3625 ( .A(n2211), .B(n2122), .Z(n2124) );
  XOR U3626 ( .A(n2212), .B(n2213), .Z(n2122) );
  ANDN U3627 ( .B(n2214), .A(n2215), .Z(n2212) );
  AND U3628 ( .A(b[4]), .B(a[99]), .Z(n2211) );
  XNOR U3629 ( .A(n2216), .B(n2217), .Z(n2136) );
  NANDN U3630 ( .A(n2218), .B(n2219), .Z(n2217) );
  XNOR U3631 ( .A(n2220), .B(n2127), .Z(n2129) );
  XNOR U3632 ( .A(n2221), .B(n2222), .Z(n2127) );
  AND U3633 ( .A(n2223), .B(n2224), .Z(n2221) );
  AND U3634 ( .A(b[3]), .B(a[100]), .Z(n2220) );
  XOR U3635 ( .A(n2143), .B(n2142), .Z(swire[102]) );
  XOR U3636 ( .A(sreg[230]), .B(n2141), .Z(n2142) );
  XOR U3637 ( .A(n2148), .B(n2225), .Z(n2143) );
  XNOR U3638 ( .A(n2147), .B(n2141), .Z(n2225) );
  XOR U3639 ( .A(n2226), .B(n2227), .Z(n2141) );
  NOR U3640 ( .A(n2228), .B(n2229), .Z(n2226) );
  NANDN U3641 ( .A(n179), .B(a[102]), .Z(n2147) );
  XNOR U3642 ( .A(n2218), .B(n2219), .Z(n2148) );
  XOR U3643 ( .A(n2216), .B(n2230), .Z(n2219) );
  NAND U3644 ( .A(b[1]), .B(a[101]), .Z(n2230) );
  XOR U3645 ( .A(n2224), .B(n2231), .Z(n2218) );
  XOR U3646 ( .A(n2216), .B(n2223), .Z(n2231) );
  XNOR U3647 ( .A(n2232), .B(n2222), .Z(n2223) );
  AND U3648 ( .A(b[2]), .B(a[100]), .Z(n2232) );
  NANDN U3649 ( .A(n2233), .B(n2234), .Z(n2216) );
  XOR U3650 ( .A(n2222), .B(n2214), .Z(n2235) );
  XNOR U3651 ( .A(n2213), .B(n2209), .Z(n2236) );
  XNOR U3652 ( .A(n2208), .B(n2204), .Z(n2237) );
  XNOR U3653 ( .A(n2203), .B(n2199), .Z(n2238) );
  XNOR U3654 ( .A(n2198), .B(n2194), .Z(n2239) );
  XNOR U3655 ( .A(n2193), .B(n2189), .Z(n2240) );
  XNOR U3656 ( .A(n2188), .B(n2184), .Z(n2241) );
  XNOR U3657 ( .A(n2183), .B(n2179), .Z(n2242) );
  XNOR U3658 ( .A(n2178), .B(n2174), .Z(n2243) );
  XOR U3659 ( .A(n2173), .B(n2170), .Z(n2244) );
  XOR U3660 ( .A(n2245), .B(n2246), .Z(n2170) );
  XOR U3661 ( .A(n2168), .B(n2247), .Z(n2246) );
  XOR U3662 ( .A(n2248), .B(n2249), .Z(n2247) );
  XOR U3663 ( .A(n2250), .B(n2251), .Z(n2249) );
  NAND U3664 ( .A(a[88]), .B(b[14]), .Z(n2251) );
  AND U3665 ( .A(a[87]), .B(b[15]), .Z(n2250) );
  XOR U3666 ( .A(n2252), .B(n2248), .Z(n2245) );
  XOR U3667 ( .A(n2253), .B(n2254), .Z(n2248) );
  NOR U3668 ( .A(n2255), .B(n2256), .Z(n2253) );
  AND U3669 ( .A(a[89]), .B(b[13]), .Z(n2252) );
  XNOR U3670 ( .A(n2257), .B(n2168), .Z(n2169) );
  XOR U3671 ( .A(n2258), .B(n2259), .Z(n2168) );
  ANDN U3672 ( .B(n2260), .A(n2261), .Z(n2258) );
  AND U3673 ( .A(a[90]), .B(b[12]), .Z(n2257) );
  XNOR U3674 ( .A(n2262), .B(n2173), .Z(n2175) );
  XOR U3675 ( .A(n2263), .B(n2264), .Z(n2173) );
  ANDN U3676 ( .B(n2265), .A(n2266), .Z(n2263) );
  AND U3677 ( .A(a[91]), .B(b[11]), .Z(n2262) );
  XNOR U3678 ( .A(n2267), .B(n2178), .Z(n2180) );
  XOR U3679 ( .A(n2268), .B(n2269), .Z(n2178) );
  ANDN U3680 ( .B(n2270), .A(n2271), .Z(n2268) );
  AND U3681 ( .A(a[92]), .B(b[10]), .Z(n2267) );
  XNOR U3682 ( .A(n2272), .B(n2183), .Z(n2185) );
  XOR U3683 ( .A(n2273), .B(n2274), .Z(n2183) );
  ANDN U3684 ( .B(n2275), .A(n2276), .Z(n2273) );
  AND U3685 ( .A(a[93]), .B(b[9]), .Z(n2272) );
  XNOR U3686 ( .A(n2277), .B(n2188), .Z(n2190) );
  XOR U3687 ( .A(n2278), .B(n2279), .Z(n2188) );
  ANDN U3688 ( .B(n2280), .A(n2281), .Z(n2278) );
  AND U3689 ( .A(a[94]), .B(b[8]), .Z(n2277) );
  XNOR U3690 ( .A(n2282), .B(n2193), .Z(n2195) );
  XOR U3691 ( .A(n2283), .B(n2284), .Z(n2193) );
  ANDN U3692 ( .B(n2285), .A(n2286), .Z(n2283) );
  AND U3693 ( .A(a[95]), .B(b[7]), .Z(n2282) );
  XNOR U3694 ( .A(n2287), .B(n2198), .Z(n2200) );
  XOR U3695 ( .A(n2288), .B(n2289), .Z(n2198) );
  ANDN U3696 ( .B(n2290), .A(n2291), .Z(n2288) );
  AND U3697 ( .A(a[96]), .B(b[6]), .Z(n2287) );
  XNOR U3698 ( .A(n2292), .B(n2203), .Z(n2205) );
  XOR U3699 ( .A(n2293), .B(n2294), .Z(n2203) );
  ANDN U3700 ( .B(n2295), .A(n2296), .Z(n2293) );
  AND U3701 ( .A(a[97]), .B(b[5]), .Z(n2292) );
  XNOR U3702 ( .A(n2297), .B(n2208), .Z(n2210) );
  XOR U3703 ( .A(n2298), .B(n2299), .Z(n2208) );
  ANDN U3704 ( .B(n2300), .A(n2301), .Z(n2298) );
  AND U3705 ( .A(b[4]), .B(a[98]), .Z(n2297) );
  XNOR U3706 ( .A(n2302), .B(n2303), .Z(n2222) );
  NANDN U3707 ( .A(n2304), .B(n2305), .Z(n2303) );
  XNOR U3708 ( .A(n2306), .B(n2213), .Z(n2215) );
  XNOR U3709 ( .A(n2307), .B(n2308), .Z(n2213) );
  AND U3710 ( .A(n2309), .B(n2310), .Z(n2307) );
  AND U3711 ( .A(b[3]), .B(a[99]), .Z(n2306) );
  XOR U3712 ( .A(n2229), .B(n2228), .Z(swire[101]) );
  XOR U3713 ( .A(sreg[229]), .B(n2227), .Z(n2228) );
  XOR U3714 ( .A(n2234), .B(n2311), .Z(n2229) );
  XNOR U3715 ( .A(n2233), .B(n2227), .Z(n2311) );
  XOR U3716 ( .A(n2312), .B(n2313), .Z(n2227) );
  NOR U3717 ( .A(n2314), .B(n2315), .Z(n2312) );
  NANDN U3718 ( .A(n179), .B(a[101]), .Z(n2233) );
  XNOR U3719 ( .A(n2304), .B(n2305), .Z(n2234) );
  XOR U3720 ( .A(n2302), .B(n2316), .Z(n2305) );
  NAND U3721 ( .A(b[1]), .B(a[100]), .Z(n2316) );
  XOR U3722 ( .A(n2310), .B(n2317), .Z(n2304) );
  XOR U3723 ( .A(n2302), .B(n2309), .Z(n2317) );
  XNOR U3724 ( .A(n2318), .B(n2308), .Z(n2309) );
  AND U3725 ( .A(b[2]), .B(a[99]), .Z(n2318) );
  NANDN U3726 ( .A(n2319), .B(n2320), .Z(n2302) );
  XOR U3727 ( .A(n2308), .B(n2300), .Z(n2321) );
  XNOR U3728 ( .A(n2299), .B(n2295), .Z(n2322) );
  XNOR U3729 ( .A(n2294), .B(n2290), .Z(n2323) );
  XNOR U3730 ( .A(n2289), .B(n2285), .Z(n2324) );
  XNOR U3731 ( .A(n2284), .B(n2280), .Z(n2325) );
  XNOR U3732 ( .A(n2279), .B(n2275), .Z(n2326) );
  XNOR U3733 ( .A(n2274), .B(n2270), .Z(n2327) );
  XNOR U3734 ( .A(n2269), .B(n2265), .Z(n2328) );
  XNOR U3735 ( .A(n2264), .B(n2260), .Z(n2329) );
  XOR U3736 ( .A(n2259), .B(n2256), .Z(n2330) );
  XOR U3737 ( .A(n2331), .B(n2332), .Z(n2256) );
  XOR U3738 ( .A(n2254), .B(n2333), .Z(n2332) );
  XOR U3739 ( .A(n2334), .B(n2335), .Z(n2333) );
  XOR U3740 ( .A(n2336), .B(n2337), .Z(n2335) );
  NAND U3741 ( .A(a[87]), .B(b[14]), .Z(n2337) );
  AND U3742 ( .A(a[86]), .B(b[15]), .Z(n2336) );
  XOR U3743 ( .A(n2338), .B(n2334), .Z(n2331) );
  XOR U3744 ( .A(n2339), .B(n2340), .Z(n2334) );
  NOR U3745 ( .A(n2341), .B(n2342), .Z(n2339) );
  AND U3746 ( .A(a[88]), .B(b[13]), .Z(n2338) );
  XNOR U3747 ( .A(n2343), .B(n2254), .Z(n2255) );
  XOR U3748 ( .A(n2344), .B(n2345), .Z(n2254) );
  ANDN U3749 ( .B(n2346), .A(n2347), .Z(n2344) );
  AND U3750 ( .A(a[89]), .B(b[12]), .Z(n2343) );
  XNOR U3751 ( .A(n2348), .B(n2259), .Z(n2261) );
  XOR U3752 ( .A(n2349), .B(n2350), .Z(n2259) );
  ANDN U3753 ( .B(n2351), .A(n2352), .Z(n2349) );
  AND U3754 ( .A(a[90]), .B(b[11]), .Z(n2348) );
  XNOR U3755 ( .A(n2353), .B(n2264), .Z(n2266) );
  XOR U3756 ( .A(n2354), .B(n2355), .Z(n2264) );
  ANDN U3757 ( .B(n2356), .A(n2357), .Z(n2354) );
  AND U3758 ( .A(a[91]), .B(b[10]), .Z(n2353) );
  XNOR U3759 ( .A(n2358), .B(n2269), .Z(n2271) );
  XOR U3760 ( .A(n2359), .B(n2360), .Z(n2269) );
  ANDN U3761 ( .B(n2361), .A(n2362), .Z(n2359) );
  AND U3762 ( .A(a[92]), .B(b[9]), .Z(n2358) );
  XNOR U3763 ( .A(n2363), .B(n2274), .Z(n2276) );
  XOR U3764 ( .A(n2364), .B(n2365), .Z(n2274) );
  ANDN U3765 ( .B(n2366), .A(n2367), .Z(n2364) );
  AND U3766 ( .A(a[93]), .B(b[8]), .Z(n2363) );
  XNOR U3767 ( .A(n2368), .B(n2279), .Z(n2281) );
  XOR U3768 ( .A(n2369), .B(n2370), .Z(n2279) );
  ANDN U3769 ( .B(n2371), .A(n2372), .Z(n2369) );
  AND U3770 ( .A(a[94]), .B(b[7]), .Z(n2368) );
  XNOR U3771 ( .A(n2373), .B(n2284), .Z(n2286) );
  XOR U3772 ( .A(n2374), .B(n2375), .Z(n2284) );
  ANDN U3773 ( .B(n2376), .A(n2377), .Z(n2374) );
  AND U3774 ( .A(a[95]), .B(b[6]), .Z(n2373) );
  XNOR U3775 ( .A(n2378), .B(n2289), .Z(n2291) );
  XOR U3776 ( .A(n2379), .B(n2380), .Z(n2289) );
  ANDN U3777 ( .B(n2381), .A(n2382), .Z(n2379) );
  AND U3778 ( .A(a[96]), .B(b[5]), .Z(n2378) );
  XNOR U3779 ( .A(n2383), .B(n2294), .Z(n2296) );
  XOR U3780 ( .A(n2384), .B(n2385), .Z(n2294) );
  ANDN U3781 ( .B(n2386), .A(n2387), .Z(n2384) );
  AND U3782 ( .A(a[97]), .B(b[4]), .Z(n2383) );
  XNOR U3783 ( .A(n2388), .B(n2389), .Z(n2308) );
  NANDN U3784 ( .A(n2390), .B(n2391), .Z(n2389) );
  XNOR U3785 ( .A(n2392), .B(n2299), .Z(n2301) );
  XNOR U3786 ( .A(n2393), .B(n2394), .Z(n2299) );
  AND U3787 ( .A(n2395), .B(n2396), .Z(n2393) );
  AND U3788 ( .A(b[3]), .B(a[98]), .Z(n2392) );
  XOR U3789 ( .A(n2315), .B(n2314), .Z(swire[100]) );
  XOR U3790 ( .A(sreg[228]), .B(n2313), .Z(n2314) );
  XOR U3791 ( .A(n2320), .B(n2397), .Z(n2315) );
  XNOR U3792 ( .A(n2319), .B(n2313), .Z(n2397) );
  XOR U3793 ( .A(n2398), .B(n2399), .Z(n2313) );
  ANDN U3794 ( .B(n2), .A(n1), .Z(n2398) );
  XOR U3795 ( .A(sreg[227]), .B(n2399), .Z(n1) );
  XOR U3796 ( .A(n2400), .B(n2401), .Z(n2) );
  XNOR U3797 ( .A(n2402), .B(n2399), .Z(n2401) );
  XOR U3798 ( .A(n2403), .B(n2404), .Z(n2399) );
  ANDN U3799 ( .B(n3), .A(n4), .Z(n2403) );
  XOR U3800 ( .A(sreg[226]), .B(n2404), .Z(n4) );
  XOR U3801 ( .A(n2405), .B(n2406), .Z(n3) );
  XNOR U3802 ( .A(n2407), .B(n2404), .Z(n2406) );
  XOR U3803 ( .A(n2408), .B(n2409), .Z(n2404) );
  ANDN U3804 ( .B(n5), .A(n6), .Z(n2408) );
  XOR U3805 ( .A(sreg[225]), .B(n2409), .Z(n6) );
  XOR U3806 ( .A(n2410), .B(n2411), .Z(n5) );
  XNOR U3807 ( .A(n2412), .B(n2409), .Z(n2411) );
  XOR U3808 ( .A(n2413), .B(n2414), .Z(n2409) );
  ANDN U3809 ( .B(n7), .A(n8), .Z(n2413) );
  XOR U3810 ( .A(sreg[224]), .B(n2414), .Z(n8) );
  XOR U3811 ( .A(n2415), .B(n2416), .Z(n7) );
  XNOR U3812 ( .A(n2417), .B(n2414), .Z(n2416) );
  XOR U3813 ( .A(n2418), .B(n2419), .Z(n2414) );
  ANDN U3814 ( .B(n9), .A(n10), .Z(n2418) );
  XOR U3815 ( .A(sreg[223]), .B(n2419), .Z(n10) );
  XOR U3816 ( .A(n2420), .B(n2421), .Z(n9) );
  XNOR U3817 ( .A(n2422), .B(n2419), .Z(n2421) );
  XOR U3818 ( .A(n2423), .B(n2424), .Z(n2419) );
  ANDN U3819 ( .B(n11), .A(n12), .Z(n2423) );
  XOR U3820 ( .A(sreg[222]), .B(n2424), .Z(n12) );
  XOR U3821 ( .A(n2425), .B(n2426), .Z(n11) );
  XNOR U3822 ( .A(n2427), .B(n2424), .Z(n2426) );
  XOR U3823 ( .A(n2428), .B(n2429), .Z(n2424) );
  ANDN U3824 ( .B(n13), .A(n14), .Z(n2428) );
  XOR U3825 ( .A(sreg[221]), .B(n2429), .Z(n14) );
  XOR U3826 ( .A(n2430), .B(n2431), .Z(n13) );
  XNOR U3827 ( .A(n2432), .B(n2429), .Z(n2431) );
  XOR U3828 ( .A(n2433), .B(n2434), .Z(n2429) );
  ANDN U3829 ( .B(n15), .A(n16), .Z(n2433) );
  XOR U3830 ( .A(sreg[220]), .B(n2434), .Z(n16) );
  XOR U3831 ( .A(n2435), .B(n2436), .Z(n15) );
  XNOR U3832 ( .A(n2437), .B(n2434), .Z(n2436) );
  XOR U3833 ( .A(n2438), .B(n2439), .Z(n2434) );
  ANDN U3834 ( .B(n17), .A(n18), .Z(n2438) );
  XOR U3835 ( .A(sreg[219]), .B(n2439), .Z(n18) );
  XOR U3836 ( .A(n2440), .B(n2441), .Z(n17) );
  XNOR U3837 ( .A(n2442), .B(n2439), .Z(n2441) );
  XOR U3838 ( .A(n2443), .B(n2444), .Z(n2439) );
  ANDN U3839 ( .B(n19), .A(n20), .Z(n2443) );
  XOR U3840 ( .A(sreg[218]), .B(n2444), .Z(n20) );
  XOR U3841 ( .A(n2445), .B(n2446), .Z(n19) );
  XNOR U3842 ( .A(n2447), .B(n2444), .Z(n2446) );
  XOR U3843 ( .A(n2448), .B(n2449), .Z(n2444) );
  ANDN U3844 ( .B(n21), .A(n22), .Z(n2448) );
  XOR U3845 ( .A(sreg[217]), .B(n2449), .Z(n22) );
  XOR U3846 ( .A(n2450), .B(n2451), .Z(n21) );
  XNOR U3847 ( .A(n2452), .B(n2449), .Z(n2451) );
  XOR U3848 ( .A(n2453), .B(n2454), .Z(n2449) );
  ANDN U3849 ( .B(n23), .A(n24), .Z(n2453) );
  XOR U3850 ( .A(sreg[216]), .B(n2454), .Z(n24) );
  XOR U3851 ( .A(n2455), .B(n2456), .Z(n23) );
  XNOR U3852 ( .A(n2457), .B(n2454), .Z(n2456) );
  XOR U3853 ( .A(n2458), .B(n2459), .Z(n2454) );
  ANDN U3854 ( .B(n25), .A(n26), .Z(n2458) );
  XOR U3855 ( .A(sreg[215]), .B(n2459), .Z(n26) );
  XOR U3856 ( .A(n2460), .B(n2461), .Z(n25) );
  XNOR U3857 ( .A(n2462), .B(n2459), .Z(n2461) );
  XOR U3858 ( .A(n2463), .B(n2464), .Z(n2459) );
  ANDN U3859 ( .B(n27), .A(n28), .Z(n2463) );
  XOR U3860 ( .A(sreg[214]), .B(n2464), .Z(n28) );
  XOR U3861 ( .A(n2465), .B(n2466), .Z(n27) );
  XNOR U3862 ( .A(n2467), .B(n2464), .Z(n2466) );
  XOR U3863 ( .A(n2468), .B(n2469), .Z(n2464) );
  ANDN U3864 ( .B(n29), .A(n30), .Z(n2468) );
  XOR U3865 ( .A(sreg[213]), .B(n2469), .Z(n30) );
  XOR U3866 ( .A(n2470), .B(n2471), .Z(n29) );
  XNOR U3867 ( .A(n2472), .B(n2469), .Z(n2471) );
  XOR U3868 ( .A(n2473), .B(n2474), .Z(n2469) );
  ANDN U3869 ( .B(n31), .A(n32), .Z(n2473) );
  XOR U3870 ( .A(sreg[212]), .B(n2474), .Z(n32) );
  XOR U3871 ( .A(n2475), .B(n2476), .Z(n31) );
  XNOR U3872 ( .A(n2477), .B(n2474), .Z(n2476) );
  XOR U3873 ( .A(n2478), .B(n2479), .Z(n2474) );
  ANDN U3874 ( .B(n33), .A(n34), .Z(n2478) );
  XOR U3875 ( .A(sreg[211]), .B(n2479), .Z(n34) );
  XOR U3876 ( .A(n2480), .B(n2481), .Z(n33) );
  XNOR U3877 ( .A(n2482), .B(n2479), .Z(n2481) );
  XOR U3878 ( .A(n2483), .B(n2484), .Z(n2479) );
  ANDN U3879 ( .B(n35), .A(n36), .Z(n2483) );
  XOR U3880 ( .A(sreg[210]), .B(n2484), .Z(n36) );
  XOR U3881 ( .A(n2485), .B(n2486), .Z(n35) );
  XNOR U3882 ( .A(n2487), .B(n2484), .Z(n2486) );
  XOR U3883 ( .A(n2488), .B(n2489), .Z(n2484) );
  ANDN U3884 ( .B(n37), .A(n38), .Z(n2488) );
  XOR U3885 ( .A(sreg[209]), .B(n2489), .Z(n38) );
  XOR U3886 ( .A(n2490), .B(n2491), .Z(n37) );
  XNOR U3887 ( .A(n2492), .B(n2489), .Z(n2491) );
  XOR U3888 ( .A(n2493), .B(n2494), .Z(n2489) );
  ANDN U3889 ( .B(n39), .A(n40), .Z(n2493) );
  XOR U3890 ( .A(sreg[208]), .B(n2494), .Z(n40) );
  XOR U3891 ( .A(n2495), .B(n2496), .Z(n39) );
  XNOR U3892 ( .A(n2497), .B(n2494), .Z(n2496) );
  XOR U3893 ( .A(n2498), .B(n2499), .Z(n2494) );
  ANDN U3894 ( .B(n41), .A(n42), .Z(n2498) );
  XOR U3895 ( .A(sreg[207]), .B(n2499), .Z(n42) );
  XOR U3896 ( .A(n2500), .B(n2501), .Z(n41) );
  XNOR U3897 ( .A(n2502), .B(n2499), .Z(n2501) );
  XOR U3898 ( .A(n2503), .B(n2504), .Z(n2499) );
  ANDN U3899 ( .B(n43), .A(n44), .Z(n2503) );
  XOR U3900 ( .A(sreg[206]), .B(n2504), .Z(n44) );
  XOR U3901 ( .A(n2505), .B(n2506), .Z(n43) );
  XNOR U3902 ( .A(n2507), .B(n2504), .Z(n2506) );
  XOR U3903 ( .A(n2508), .B(n2509), .Z(n2504) );
  ANDN U3904 ( .B(n45), .A(n46), .Z(n2508) );
  XOR U3905 ( .A(sreg[205]), .B(n2509), .Z(n46) );
  XOR U3906 ( .A(n2510), .B(n2511), .Z(n45) );
  XNOR U3907 ( .A(n2512), .B(n2509), .Z(n2511) );
  XOR U3908 ( .A(n2513), .B(n2514), .Z(n2509) );
  ANDN U3909 ( .B(n47), .A(n48), .Z(n2513) );
  XOR U3910 ( .A(sreg[204]), .B(n2514), .Z(n48) );
  XOR U3911 ( .A(n2515), .B(n2516), .Z(n47) );
  XNOR U3912 ( .A(n2517), .B(n2514), .Z(n2516) );
  XOR U3913 ( .A(n2518), .B(n2519), .Z(n2514) );
  ANDN U3914 ( .B(n49), .A(n50), .Z(n2518) );
  XOR U3915 ( .A(sreg[203]), .B(n2519), .Z(n50) );
  XOR U3916 ( .A(n2520), .B(n2521), .Z(n49) );
  XNOR U3917 ( .A(n2522), .B(n2519), .Z(n2521) );
  XOR U3918 ( .A(n2523), .B(n2524), .Z(n2519) );
  ANDN U3919 ( .B(n51), .A(n52), .Z(n2523) );
  XOR U3920 ( .A(sreg[202]), .B(n2524), .Z(n52) );
  XOR U3921 ( .A(n2525), .B(n2526), .Z(n51) );
  XNOR U3922 ( .A(n2527), .B(n2524), .Z(n2526) );
  XOR U3923 ( .A(n2528), .B(n2529), .Z(n2524) );
  ANDN U3924 ( .B(n53), .A(n54), .Z(n2528) );
  XOR U3925 ( .A(sreg[201]), .B(n2529), .Z(n54) );
  XOR U3926 ( .A(n2530), .B(n2531), .Z(n53) );
  XNOR U3927 ( .A(n2532), .B(n2529), .Z(n2531) );
  XOR U3928 ( .A(n2533), .B(n2534), .Z(n2529) );
  ANDN U3929 ( .B(n55), .A(n56), .Z(n2533) );
  XOR U3930 ( .A(sreg[200]), .B(n2534), .Z(n56) );
  XOR U3931 ( .A(n2535), .B(n2536), .Z(n55) );
  XNOR U3932 ( .A(n2537), .B(n2534), .Z(n2536) );
  XOR U3933 ( .A(n2538), .B(n2539), .Z(n2534) );
  ANDN U3934 ( .B(n57), .A(n58), .Z(n2538) );
  XOR U3935 ( .A(sreg[199]), .B(n2539), .Z(n58) );
  XOR U3936 ( .A(n2540), .B(n2541), .Z(n57) );
  XNOR U3937 ( .A(n2542), .B(n2539), .Z(n2541) );
  XOR U3938 ( .A(n2543), .B(n2544), .Z(n2539) );
  ANDN U3939 ( .B(n59), .A(n60), .Z(n2543) );
  XOR U3940 ( .A(sreg[198]), .B(n2544), .Z(n60) );
  XOR U3941 ( .A(n2545), .B(n2546), .Z(n59) );
  XNOR U3942 ( .A(n2547), .B(n2544), .Z(n2546) );
  XOR U3943 ( .A(n2548), .B(n2549), .Z(n2544) );
  ANDN U3944 ( .B(n61), .A(n62), .Z(n2548) );
  XOR U3945 ( .A(sreg[197]), .B(n2549), .Z(n62) );
  XOR U3946 ( .A(n2550), .B(n2551), .Z(n61) );
  XNOR U3947 ( .A(n2552), .B(n2549), .Z(n2551) );
  XOR U3948 ( .A(n2553), .B(n2554), .Z(n2549) );
  ANDN U3949 ( .B(n63), .A(n64), .Z(n2553) );
  XOR U3950 ( .A(sreg[196]), .B(n2554), .Z(n64) );
  XOR U3951 ( .A(n2555), .B(n2556), .Z(n63) );
  XNOR U3952 ( .A(n2557), .B(n2554), .Z(n2556) );
  XOR U3953 ( .A(n2558), .B(n2559), .Z(n2554) );
  ANDN U3954 ( .B(n65), .A(n66), .Z(n2558) );
  XOR U3955 ( .A(sreg[195]), .B(n2559), .Z(n66) );
  XOR U3956 ( .A(n2560), .B(n2561), .Z(n65) );
  XNOR U3957 ( .A(n2562), .B(n2559), .Z(n2561) );
  XOR U3958 ( .A(n2563), .B(n2564), .Z(n2559) );
  ANDN U3959 ( .B(n67), .A(n68), .Z(n2563) );
  XOR U3960 ( .A(sreg[194]), .B(n2564), .Z(n68) );
  XOR U3961 ( .A(n2565), .B(n2566), .Z(n67) );
  XNOR U3962 ( .A(n2567), .B(n2564), .Z(n2566) );
  XOR U3963 ( .A(n2568), .B(n2569), .Z(n2564) );
  ANDN U3964 ( .B(n69), .A(n70), .Z(n2568) );
  XOR U3965 ( .A(sreg[193]), .B(n2569), .Z(n70) );
  XOR U3966 ( .A(n2570), .B(n2571), .Z(n69) );
  XNOR U3967 ( .A(n2572), .B(n2569), .Z(n2571) );
  XOR U3968 ( .A(n2573), .B(n2574), .Z(n2569) );
  ANDN U3969 ( .B(n71), .A(n72), .Z(n2573) );
  XOR U3970 ( .A(sreg[192]), .B(n2574), .Z(n72) );
  XOR U3971 ( .A(n2575), .B(n2576), .Z(n71) );
  XNOR U3972 ( .A(n2577), .B(n2574), .Z(n2576) );
  XOR U3973 ( .A(n2578), .B(n2579), .Z(n2574) );
  ANDN U3974 ( .B(n73), .A(n74), .Z(n2578) );
  XOR U3975 ( .A(sreg[191]), .B(n2579), .Z(n74) );
  XOR U3976 ( .A(n2580), .B(n2581), .Z(n73) );
  XNOR U3977 ( .A(n2582), .B(n2579), .Z(n2581) );
  XOR U3978 ( .A(n2583), .B(n2584), .Z(n2579) );
  ANDN U3979 ( .B(n75), .A(n76), .Z(n2583) );
  XOR U3980 ( .A(sreg[190]), .B(n2584), .Z(n76) );
  XOR U3981 ( .A(n2585), .B(n2586), .Z(n75) );
  XNOR U3982 ( .A(n2587), .B(n2584), .Z(n2586) );
  XOR U3983 ( .A(n2588), .B(n2589), .Z(n2584) );
  ANDN U3984 ( .B(n77), .A(n78), .Z(n2588) );
  XOR U3985 ( .A(sreg[189]), .B(n2589), .Z(n78) );
  XOR U3986 ( .A(n2590), .B(n2591), .Z(n77) );
  XNOR U3987 ( .A(n2592), .B(n2589), .Z(n2591) );
  XOR U3988 ( .A(n2593), .B(n2594), .Z(n2589) );
  ANDN U3989 ( .B(n79), .A(n80), .Z(n2593) );
  XOR U3990 ( .A(sreg[188]), .B(n2594), .Z(n80) );
  XOR U3991 ( .A(n2595), .B(n2596), .Z(n79) );
  XNOR U3992 ( .A(n2597), .B(n2594), .Z(n2596) );
  XOR U3993 ( .A(n2598), .B(n2599), .Z(n2594) );
  ANDN U3994 ( .B(n81), .A(n82), .Z(n2598) );
  XOR U3995 ( .A(sreg[187]), .B(n2599), .Z(n82) );
  XOR U3996 ( .A(n2600), .B(n2601), .Z(n81) );
  XNOR U3997 ( .A(n2602), .B(n2599), .Z(n2601) );
  XOR U3998 ( .A(n2603), .B(n2604), .Z(n2599) );
  ANDN U3999 ( .B(n83), .A(n84), .Z(n2603) );
  XOR U4000 ( .A(sreg[186]), .B(n2604), .Z(n84) );
  XOR U4001 ( .A(n2605), .B(n2606), .Z(n83) );
  XNOR U4002 ( .A(n2607), .B(n2604), .Z(n2606) );
  XOR U4003 ( .A(n2608), .B(n2609), .Z(n2604) );
  ANDN U4004 ( .B(n85), .A(n86), .Z(n2608) );
  XOR U4005 ( .A(sreg[185]), .B(n2609), .Z(n86) );
  XOR U4006 ( .A(n2610), .B(n2611), .Z(n85) );
  XNOR U4007 ( .A(n2612), .B(n2609), .Z(n2611) );
  XOR U4008 ( .A(n2613), .B(n2614), .Z(n2609) );
  ANDN U4009 ( .B(n87), .A(n88), .Z(n2613) );
  XOR U4010 ( .A(sreg[184]), .B(n2614), .Z(n88) );
  XOR U4011 ( .A(n2615), .B(n2616), .Z(n87) );
  XNOR U4012 ( .A(n2617), .B(n2614), .Z(n2616) );
  XOR U4013 ( .A(n2618), .B(n2619), .Z(n2614) );
  ANDN U4014 ( .B(n89), .A(n90), .Z(n2618) );
  XOR U4015 ( .A(sreg[183]), .B(n2619), .Z(n90) );
  XOR U4016 ( .A(n2620), .B(n2621), .Z(n89) );
  XNOR U4017 ( .A(n2622), .B(n2619), .Z(n2621) );
  XOR U4018 ( .A(n2623), .B(n2624), .Z(n2619) );
  ANDN U4019 ( .B(n91), .A(n92), .Z(n2623) );
  XOR U4020 ( .A(sreg[182]), .B(n2624), .Z(n92) );
  XOR U4021 ( .A(n2625), .B(n2626), .Z(n91) );
  XNOR U4022 ( .A(n2627), .B(n2624), .Z(n2626) );
  XOR U4023 ( .A(n2628), .B(n2629), .Z(n2624) );
  ANDN U4024 ( .B(n93), .A(n94), .Z(n2628) );
  XOR U4025 ( .A(sreg[181]), .B(n2629), .Z(n94) );
  XOR U4026 ( .A(n2630), .B(n2631), .Z(n93) );
  XNOR U4027 ( .A(n2632), .B(n2629), .Z(n2631) );
  XOR U4028 ( .A(n2633), .B(n2634), .Z(n2629) );
  ANDN U4029 ( .B(n95), .A(n96), .Z(n2633) );
  XOR U4030 ( .A(sreg[180]), .B(n2634), .Z(n96) );
  XOR U4031 ( .A(n2635), .B(n2636), .Z(n95) );
  XNOR U4032 ( .A(n2637), .B(n2634), .Z(n2636) );
  XOR U4033 ( .A(n2638), .B(n2639), .Z(n2634) );
  ANDN U4034 ( .B(n97), .A(n98), .Z(n2638) );
  XOR U4035 ( .A(sreg[179]), .B(n2639), .Z(n98) );
  XOR U4036 ( .A(n2640), .B(n2641), .Z(n97) );
  XNOR U4037 ( .A(n2642), .B(n2639), .Z(n2641) );
  XOR U4038 ( .A(n2643), .B(n2644), .Z(n2639) );
  ANDN U4039 ( .B(n99), .A(n100), .Z(n2643) );
  XOR U4040 ( .A(sreg[178]), .B(n2644), .Z(n100) );
  XOR U4041 ( .A(n2645), .B(n2646), .Z(n99) );
  XNOR U4042 ( .A(n2647), .B(n2644), .Z(n2646) );
  XOR U4043 ( .A(n2648), .B(n2649), .Z(n2644) );
  ANDN U4044 ( .B(n101), .A(n102), .Z(n2648) );
  XOR U4045 ( .A(sreg[177]), .B(n2649), .Z(n102) );
  XOR U4046 ( .A(n2650), .B(n2651), .Z(n101) );
  XNOR U4047 ( .A(n2652), .B(n2649), .Z(n2651) );
  XOR U4048 ( .A(n2653), .B(n2654), .Z(n2649) );
  ANDN U4049 ( .B(n103), .A(n104), .Z(n2653) );
  XOR U4050 ( .A(sreg[176]), .B(n2654), .Z(n104) );
  XOR U4051 ( .A(n2655), .B(n2656), .Z(n103) );
  XNOR U4052 ( .A(n2657), .B(n2654), .Z(n2656) );
  XOR U4053 ( .A(n2658), .B(n2659), .Z(n2654) );
  ANDN U4054 ( .B(n105), .A(n106), .Z(n2658) );
  XOR U4055 ( .A(sreg[175]), .B(n2659), .Z(n106) );
  XOR U4056 ( .A(n2660), .B(n2661), .Z(n105) );
  XNOR U4057 ( .A(n2662), .B(n2659), .Z(n2661) );
  XOR U4058 ( .A(n2663), .B(n2664), .Z(n2659) );
  ANDN U4059 ( .B(n107), .A(n108), .Z(n2663) );
  XOR U4060 ( .A(sreg[174]), .B(n2664), .Z(n108) );
  XOR U4061 ( .A(n2665), .B(n2666), .Z(n107) );
  XNOR U4062 ( .A(n2667), .B(n2664), .Z(n2666) );
  XOR U4063 ( .A(n2668), .B(n2669), .Z(n2664) );
  ANDN U4064 ( .B(n109), .A(n110), .Z(n2668) );
  XOR U4065 ( .A(sreg[173]), .B(n2669), .Z(n110) );
  XOR U4066 ( .A(n2670), .B(n2671), .Z(n109) );
  XNOR U4067 ( .A(n2672), .B(n2669), .Z(n2671) );
  XOR U4068 ( .A(n2673), .B(n2674), .Z(n2669) );
  ANDN U4069 ( .B(n111), .A(n112), .Z(n2673) );
  XOR U4070 ( .A(sreg[172]), .B(n2674), .Z(n112) );
  XOR U4071 ( .A(n2675), .B(n2676), .Z(n111) );
  XNOR U4072 ( .A(n2677), .B(n2674), .Z(n2676) );
  XOR U4073 ( .A(n2678), .B(n2679), .Z(n2674) );
  ANDN U4074 ( .B(n113), .A(n114), .Z(n2678) );
  XOR U4075 ( .A(sreg[171]), .B(n2679), .Z(n114) );
  XOR U4076 ( .A(n2680), .B(n2681), .Z(n113) );
  XNOR U4077 ( .A(n2682), .B(n2679), .Z(n2681) );
  XOR U4078 ( .A(n2683), .B(n2684), .Z(n2679) );
  ANDN U4079 ( .B(n115), .A(n116), .Z(n2683) );
  XOR U4080 ( .A(sreg[170]), .B(n2684), .Z(n116) );
  XOR U4081 ( .A(n2685), .B(n2686), .Z(n115) );
  XNOR U4082 ( .A(n2687), .B(n2684), .Z(n2686) );
  XOR U4083 ( .A(n2688), .B(n2689), .Z(n2684) );
  ANDN U4084 ( .B(n117), .A(n118), .Z(n2688) );
  XOR U4085 ( .A(sreg[169]), .B(n2689), .Z(n118) );
  XOR U4086 ( .A(n2690), .B(n2691), .Z(n117) );
  XNOR U4087 ( .A(n2692), .B(n2689), .Z(n2691) );
  XOR U4088 ( .A(n2693), .B(n2694), .Z(n2689) );
  ANDN U4089 ( .B(n119), .A(n120), .Z(n2693) );
  XOR U4090 ( .A(sreg[168]), .B(n2694), .Z(n120) );
  XOR U4091 ( .A(n2695), .B(n2696), .Z(n119) );
  XNOR U4092 ( .A(n2697), .B(n2694), .Z(n2696) );
  XOR U4093 ( .A(n2698), .B(n2699), .Z(n2694) );
  ANDN U4094 ( .B(n121), .A(n122), .Z(n2698) );
  XOR U4095 ( .A(sreg[167]), .B(n2699), .Z(n122) );
  XOR U4096 ( .A(n2700), .B(n2701), .Z(n121) );
  XNOR U4097 ( .A(n2702), .B(n2699), .Z(n2701) );
  XOR U4098 ( .A(n2703), .B(n2704), .Z(n2699) );
  ANDN U4099 ( .B(n123), .A(n124), .Z(n2703) );
  XOR U4100 ( .A(sreg[166]), .B(n2704), .Z(n124) );
  XOR U4101 ( .A(n2705), .B(n2706), .Z(n123) );
  XNOR U4102 ( .A(n2707), .B(n2704), .Z(n2706) );
  XOR U4103 ( .A(n2708), .B(n2709), .Z(n2704) );
  ANDN U4104 ( .B(n125), .A(n126), .Z(n2708) );
  XOR U4105 ( .A(sreg[165]), .B(n2709), .Z(n126) );
  XOR U4106 ( .A(n2710), .B(n2711), .Z(n125) );
  XNOR U4107 ( .A(n2712), .B(n2709), .Z(n2711) );
  XOR U4108 ( .A(n2713), .B(n2714), .Z(n2709) );
  ANDN U4109 ( .B(n127), .A(n128), .Z(n2713) );
  XOR U4110 ( .A(sreg[164]), .B(n2714), .Z(n128) );
  XOR U4111 ( .A(n2715), .B(n2716), .Z(n127) );
  XNOR U4112 ( .A(n2717), .B(n2714), .Z(n2716) );
  XOR U4113 ( .A(n2718), .B(n2719), .Z(n2714) );
  ANDN U4114 ( .B(n129), .A(n130), .Z(n2718) );
  XOR U4115 ( .A(sreg[163]), .B(n2719), .Z(n130) );
  XOR U4116 ( .A(n2720), .B(n2721), .Z(n129) );
  XNOR U4117 ( .A(n2722), .B(n2719), .Z(n2721) );
  XOR U4118 ( .A(n2723), .B(n2724), .Z(n2719) );
  ANDN U4119 ( .B(n131), .A(n132), .Z(n2723) );
  XOR U4120 ( .A(sreg[162]), .B(n2724), .Z(n132) );
  XOR U4121 ( .A(n2725), .B(n2726), .Z(n131) );
  XNOR U4122 ( .A(n2727), .B(n2724), .Z(n2726) );
  XOR U4123 ( .A(n2728), .B(n2729), .Z(n2724) );
  ANDN U4124 ( .B(n133), .A(n134), .Z(n2728) );
  XOR U4125 ( .A(sreg[161]), .B(n2729), .Z(n134) );
  XOR U4126 ( .A(n2730), .B(n2731), .Z(n133) );
  XNOR U4127 ( .A(n2732), .B(n2729), .Z(n2731) );
  XOR U4128 ( .A(n2733), .B(n2734), .Z(n2729) );
  ANDN U4129 ( .B(n135), .A(n136), .Z(n2733) );
  XOR U4130 ( .A(sreg[160]), .B(n2734), .Z(n136) );
  XOR U4131 ( .A(n2735), .B(n2736), .Z(n135) );
  XNOR U4132 ( .A(n2737), .B(n2734), .Z(n2736) );
  XOR U4133 ( .A(n2738), .B(n2739), .Z(n2734) );
  ANDN U4134 ( .B(n137), .A(n138), .Z(n2738) );
  XOR U4135 ( .A(sreg[159]), .B(n2739), .Z(n138) );
  XOR U4136 ( .A(n2740), .B(n2741), .Z(n137) );
  XNOR U4137 ( .A(n2742), .B(n2739), .Z(n2741) );
  XOR U4138 ( .A(n2743), .B(n2744), .Z(n2739) );
  ANDN U4139 ( .B(n139), .A(n140), .Z(n2743) );
  XOR U4140 ( .A(sreg[158]), .B(n2744), .Z(n140) );
  XOR U4141 ( .A(n2745), .B(n2746), .Z(n139) );
  XNOR U4142 ( .A(n2747), .B(n2744), .Z(n2746) );
  XOR U4143 ( .A(n2748), .B(n2749), .Z(n2744) );
  ANDN U4144 ( .B(n141), .A(n142), .Z(n2748) );
  XOR U4145 ( .A(sreg[157]), .B(n2749), .Z(n142) );
  XOR U4146 ( .A(n2750), .B(n2751), .Z(n141) );
  XNOR U4147 ( .A(n2752), .B(n2749), .Z(n2751) );
  XOR U4148 ( .A(n2753), .B(n2754), .Z(n2749) );
  ANDN U4149 ( .B(n143), .A(n144), .Z(n2753) );
  XOR U4150 ( .A(sreg[156]), .B(n2754), .Z(n144) );
  XOR U4151 ( .A(n2755), .B(n2756), .Z(n143) );
  XNOR U4152 ( .A(n2757), .B(n2754), .Z(n2756) );
  XOR U4153 ( .A(n2758), .B(n2759), .Z(n2754) );
  ANDN U4154 ( .B(n145), .A(n146), .Z(n2758) );
  XOR U4155 ( .A(sreg[155]), .B(n2759), .Z(n146) );
  XOR U4156 ( .A(n2760), .B(n2761), .Z(n145) );
  XNOR U4157 ( .A(n2762), .B(n2759), .Z(n2761) );
  XOR U4158 ( .A(n2763), .B(n2764), .Z(n2759) );
  ANDN U4159 ( .B(n147), .A(n148), .Z(n2763) );
  XOR U4160 ( .A(sreg[154]), .B(n2764), .Z(n148) );
  XOR U4161 ( .A(n2765), .B(n2766), .Z(n147) );
  XNOR U4162 ( .A(n2767), .B(n2764), .Z(n2766) );
  XOR U4163 ( .A(n2768), .B(n2769), .Z(n2764) );
  ANDN U4164 ( .B(n149), .A(n150), .Z(n2768) );
  XOR U4165 ( .A(sreg[153]), .B(n2769), .Z(n150) );
  XOR U4166 ( .A(n2770), .B(n2771), .Z(n149) );
  XNOR U4167 ( .A(n2772), .B(n2769), .Z(n2771) );
  XOR U4168 ( .A(n2773), .B(n2774), .Z(n2769) );
  ANDN U4169 ( .B(n151), .A(n152), .Z(n2773) );
  XOR U4170 ( .A(sreg[152]), .B(n2774), .Z(n152) );
  XOR U4171 ( .A(n2775), .B(n2776), .Z(n151) );
  XNOR U4172 ( .A(n2777), .B(n2774), .Z(n2776) );
  XOR U4173 ( .A(n2778), .B(n2779), .Z(n2774) );
  ANDN U4174 ( .B(n153), .A(n154), .Z(n2778) );
  XOR U4175 ( .A(sreg[151]), .B(n2779), .Z(n154) );
  XOR U4176 ( .A(n2780), .B(n2781), .Z(n153) );
  XNOR U4177 ( .A(n2782), .B(n2779), .Z(n2781) );
  XOR U4178 ( .A(n2783), .B(n2784), .Z(n2779) );
  ANDN U4179 ( .B(n155), .A(n156), .Z(n2783) );
  XOR U4180 ( .A(sreg[150]), .B(n2784), .Z(n156) );
  XOR U4181 ( .A(n2785), .B(n2786), .Z(n155) );
  XNOR U4182 ( .A(n2787), .B(n2784), .Z(n2786) );
  XOR U4183 ( .A(n2788), .B(n2789), .Z(n2784) );
  ANDN U4184 ( .B(n157), .A(n158), .Z(n2788) );
  XOR U4185 ( .A(sreg[149]), .B(n2789), .Z(n158) );
  XOR U4186 ( .A(n2790), .B(n2791), .Z(n157) );
  XNOR U4187 ( .A(n2792), .B(n2789), .Z(n2791) );
  XOR U4188 ( .A(n2793), .B(n2794), .Z(n2789) );
  ANDN U4189 ( .B(n159), .A(n160), .Z(n2793) );
  XOR U4190 ( .A(sreg[148]), .B(n2794), .Z(n160) );
  XOR U4191 ( .A(n2795), .B(n2796), .Z(n159) );
  XNOR U4192 ( .A(n2797), .B(n2794), .Z(n2796) );
  XOR U4193 ( .A(n2798), .B(n2799), .Z(n2794) );
  ANDN U4194 ( .B(n161), .A(n162), .Z(n2798) );
  XOR U4195 ( .A(sreg[147]), .B(n2799), .Z(n162) );
  XOR U4196 ( .A(n2800), .B(n2801), .Z(n161) );
  XNOR U4197 ( .A(n2802), .B(n2799), .Z(n2801) );
  XOR U4198 ( .A(n2803), .B(n2804), .Z(n2799) );
  ANDN U4199 ( .B(n163), .A(n164), .Z(n2803) );
  XOR U4200 ( .A(sreg[146]), .B(n2804), .Z(n164) );
  XOR U4201 ( .A(n2805), .B(n2806), .Z(n163) );
  XNOR U4202 ( .A(n2807), .B(n2804), .Z(n2806) );
  XOR U4203 ( .A(n2808), .B(n2809), .Z(n2804) );
  ANDN U4204 ( .B(n165), .A(n166), .Z(n2808) );
  XOR U4205 ( .A(sreg[145]), .B(n2809), .Z(n166) );
  XOR U4206 ( .A(n2810), .B(n2811), .Z(n165) );
  XNOR U4207 ( .A(n2812), .B(n2809), .Z(n2811) );
  XOR U4208 ( .A(n2813), .B(n2814), .Z(n2809) );
  ANDN U4209 ( .B(n167), .A(n168), .Z(n2813) );
  XOR U4210 ( .A(sreg[144]), .B(n2814), .Z(n168) );
  XOR U4211 ( .A(n2815), .B(n2816), .Z(n167) );
  XNOR U4212 ( .A(n2817), .B(n2814), .Z(n2816) );
  XOR U4213 ( .A(n2818), .B(n2819), .Z(n2814) );
  ANDN U4214 ( .B(n2820), .A(n2821), .Z(n2818) );
  NANDN U4215 ( .A(n179), .B(a[100]), .Z(n2319) );
  XNOR U4216 ( .A(n2390), .B(n2391), .Z(n2320) );
  XOR U4217 ( .A(n2388), .B(n2822), .Z(n2391) );
  NAND U4218 ( .A(b[1]), .B(a[99]), .Z(n2822) );
  XOR U4219 ( .A(n2396), .B(n2823), .Z(n2390) );
  XOR U4220 ( .A(n2388), .B(n2395), .Z(n2823) );
  XNOR U4221 ( .A(n2824), .B(n2394), .Z(n2395) );
  AND U4222 ( .A(b[2]), .B(a[98]), .Z(n2824) );
  OR U4223 ( .A(n2402), .B(n2400), .Z(n2388) );
  XOR U4224 ( .A(n2825), .B(n2826), .Z(n2400) );
  NANDN U4225 ( .A(n179), .B(a[99]), .Z(n2402) );
  XOR U4226 ( .A(n2394), .B(n2386), .Z(n2827) );
  XNOR U4227 ( .A(n2385), .B(n2381), .Z(n2828) );
  XNOR U4228 ( .A(n2380), .B(n2376), .Z(n2829) );
  XNOR U4229 ( .A(n2375), .B(n2371), .Z(n2830) );
  XNOR U4230 ( .A(n2370), .B(n2366), .Z(n2831) );
  XNOR U4231 ( .A(n2365), .B(n2361), .Z(n2832) );
  XNOR U4232 ( .A(n2360), .B(n2356), .Z(n2833) );
  XNOR U4233 ( .A(n2355), .B(n2351), .Z(n2834) );
  XNOR U4234 ( .A(n2350), .B(n2346), .Z(n2835) );
  XOR U4235 ( .A(n2345), .B(n2342), .Z(n2836) );
  XOR U4236 ( .A(n2837), .B(n2838), .Z(n2342) );
  XOR U4237 ( .A(n2340), .B(n2839), .Z(n2838) );
  XNOR U4238 ( .A(n2840), .B(n2841), .Z(n2839) );
  XOR U4239 ( .A(n2842), .B(n2843), .Z(n2841) );
  NAND U4240 ( .A(a[86]), .B(b[14]), .Z(n2843) );
  AND U4241 ( .A(a[85]), .B(b[15]), .Z(n2842) );
  XNOR U4242 ( .A(n2844), .B(n2840), .Z(n2837) );
  XOR U4243 ( .A(n2845), .B(n2846), .Z(n2840) );
  NOR U4244 ( .A(n2847), .B(n2848), .Z(n2845) );
  AND U4245 ( .A(a[87]), .B(b[13]), .Z(n2844) );
  XNOR U4246 ( .A(n2849), .B(n2340), .Z(n2341) );
  XNOR U4247 ( .A(n2850), .B(n2851), .Z(n2340) );
  ANDN U4248 ( .B(n2852), .A(n2853), .Z(n2850) );
  AND U4249 ( .A(a[88]), .B(b[12]), .Z(n2849) );
  XNOR U4250 ( .A(n2854), .B(n2345), .Z(n2347) );
  XNOR U4251 ( .A(n2855), .B(n2856), .Z(n2345) );
  ANDN U4252 ( .B(n2857), .A(n2858), .Z(n2855) );
  AND U4253 ( .A(a[89]), .B(b[11]), .Z(n2854) );
  XNOR U4254 ( .A(n2859), .B(n2350), .Z(n2352) );
  XNOR U4255 ( .A(n2860), .B(n2861), .Z(n2350) );
  ANDN U4256 ( .B(n2862), .A(n2863), .Z(n2860) );
  AND U4257 ( .A(a[90]), .B(b[10]), .Z(n2859) );
  XNOR U4258 ( .A(n2864), .B(n2355), .Z(n2357) );
  XNOR U4259 ( .A(n2865), .B(n2866), .Z(n2355) );
  ANDN U4260 ( .B(n2867), .A(n2868), .Z(n2865) );
  AND U4261 ( .A(a[91]), .B(b[9]), .Z(n2864) );
  XNOR U4262 ( .A(n2869), .B(n2360), .Z(n2362) );
  XNOR U4263 ( .A(n2870), .B(n2871), .Z(n2360) );
  ANDN U4264 ( .B(n2872), .A(n2873), .Z(n2870) );
  AND U4265 ( .A(a[92]), .B(b[8]), .Z(n2869) );
  XNOR U4266 ( .A(n2874), .B(n2365), .Z(n2367) );
  XNOR U4267 ( .A(n2875), .B(n2876), .Z(n2365) );
  ANDN U4268 ( .B(n2877), .A(n2878), .Z(n2875) );
  AND U4269 ( .A(a[93]), .B(b[7]), .Z(n2874) );
  XNOR U4270 ( .A(n2879), .B(n2370), .Z(n2372) );
  XNOR U4271 ( .A(n2880), .B(n2881), .Z(n2370) );
  ANDN U4272 ( .B(n2882), .A(n2883), .Z(n2880) );
  AND U4273 ( .A(a[94]), .B(b[6]), .Z(n2879) );
  XNOR U4274 ( .A(n2884), .B(n2375), .Z(n2377) );
  XNOR U4275 ( .A(n2885), .B(n2886), .Z(n2375) );
  ANDN U4276 ( .B(n2887), .A(n2888), .Z(n2885) );
  AND U4277 ( .A(a[95]), .B(b[5]), .Z(n2884) );
  XNOR U4278 ( .A(n2889), .B(n2380), .Z(n2382) );
  XNOR U4279 ( .A(n2890), .B(n2891), .Z(n2380) );
  ANDN U4280 ( .B(n2892), .A(n2893), .Z(n2890) );
  AND U4281 ( .A(a[96]), .B(b[4]), .Z(n2889) );
  XNOR U4282 ( .A(n2894), .B(n2895), .Z(n2394) );
  NANDN U4283 ( .A(n2826), .B(n2825), .Z(n2895) );
  XOR U4284 ( .A(n2894), .B(n2896), .Z(n2825) );
  NAND U4285 ( .A(b[1]), .B(a[98]), .Z(n2896) );
  XOR U4286 ( .A(n2894), .B(n2898), .Z(n2897) );
  OR U4287 ( .A(n2407), .B(n2405), .Z(n2894) );
  XOR U4288 ( .A(n2900), .B(n2901), .Z(n2405) );
  NANDN U4289 ( .A(n179), .B(a[98]), .Z(n2407) );
  XNOR U4290 ( .A(n2902), .B(n2385), .Z(n2387) );
  XNOR U4291 ( .A(n2903), .B(n2904), .Z(n2385) );
  ANDN U4292 ( .B(n2898), .A(n2899), .Z(n2903) );
  XOR U4293 ( .A(n2905), .B(n2904), .Z(n2899) );
  IV U4294 ( .A(n2906), .Z(n2904) );
  AND U4295 ( .A(a[97]), .B(b[2]), .Z(n2905) );
  XNOR U4296 ( .A(n2892), .B(n2906), .Z(n2907) );
  XOR U4297 ( .A(n2908), .B(n2909), .Z(n2906) );
  NANDN U4298 ( .A(n2901), .B(n2900), .Z(n2909) );
  XOR U4299 ( .A(n2908), .B(n2910), .Z(n2900) );
  NAND U4300 ( .A(a[97]), .B(b[1]), .Z(n2910) );
  XOR U4301 ( .A(n2908), .B(n2912), .Z(n2911) );
  OR U4302 ( .A(n2412), .B(n2410), .Z(n2908) );
  XOR U4303 ( .A(n2914), .B(n2915), .Z(n2410) );
  NANDN U4304 ( .A(n179), .B(a[97]), .Z(n2412) );
  XNOR U4305 ( .A(n2887), .B(n2917), .Z(n2916) );
  XNOR U4306 ( .A(n2882), .B(n2919), .Z(n2918) );
  XNOR U4307 ( .A(n2877), .B(n2921), .Z(n2920) );
  XNOR U4308 ( .A(n2872), .B(n2923), .Z(n2922) );
  XNOR U4309 ( .A(n2867), .B(n2925), .Z(n2924) );
  XNOR U4310 ( .A(n2862), .B(n2927), .Z(n2926) );
  XNOR U4311 ( .A(n2857), .B(n2929), .Z(n2928) );
  XNOR U4312 ( .A(n2852), .B(n2931), .Z(n2930) );
  XOR U4313 ( .A(n2848), .B(n2933), .Z(n2932) );
  XOR U4314 ( .A(n2934), .B(n2935), .Z(n2848) );
  XNOR U4315 ( .A(n2936), .B(n2937), .Z(n2935) );
  XNOR U4316 ( .A(n2938), .B(n2939), .Z(n2936) );
  XOR U4317 ( .A(n2940), .B(n2941), .Z(n2939) );
  AND U4318 ( .A(b[15]), .B(a[84]), .Z(n2941) );
  AND U4319 ( .A(a[85]), .B(b[14]), .Z(n2940) );
  XNOR U4320 ( .A(n2942), .B(n2938), .Z(n2934) );
  XOR U4321 ( .A(n2943), .B(n2944), .Z(n2938) );
  NOR U4322 ( .A(n2945), .B(n2946), .Z(n2943) );
  AND U4323 ( .A(a[86]), .B(b[13]), .Z(n2942) );
  XOR U4324 ( .A(n2947), .B(n2846), .Z(n2847) );
  IV U4325 ( .A(n2937), .Z(n2846) );
  XOR U4326 ( .A(n2948), .B(n2949), .Z(n2937) );
  ANDN U4327 ( .B(n2950), .A(n2951), .Z(n2948) );
  AND U4328 ( .A(a[87]), .B(b[12]), .Z(n2947) );
  XOR U4329 ( .A(n2952), .B(n2851), .Z(n2853) );
  IV U4330 ( .A(n2933), .Z(n2851) );
  XOR U4331 ( .A(n2953), .B(n2954), .Z(n2933) );
  ANDN U4332 ( .B(n2955), .A(n2956), .Z(n2953) );
  AND U4333 ( .A(a[88]), .B(b[11]), .Z(n2952) );
  XOR U4334 ( .A(n2957), .B(n2856), .Z(n2858) );
  IV U4335 ( .A(n2931), .Z(n2856) );
  XOR U4336 ( .A(n2958), .B(n2959), .Z(n2931) );
  ANDN U4337 ( .B(n2960), .A(n2961), .Z(n2958) );
  AND U4338 ( .A(a[89]), .B(b[10]), .Z(n2957) );
  XOR U4339 ( .A(n2962), .B(n2861), .Z(n2863) );
  IV U4340 ( .A(n2929), .Z(n2861) );
  XOR U4341 ( .A(n2963), .B(n2964), .Z(n2929) );
  ANDN U4342 ( .B(n2965), .A(n2966), .Z(n2963) );
  AND U4343 ( .A(a[90]), .B(b[9]), .Z(n2962) );
  XOR U4344 ( .A(n2967), .B(n2866), .Z(n2868) );
  IV U4345 ( .A(n2927), .Z(n2866) );
  XOR U4346 ( .A(n2968), .B(n2969), .Z(n2927) );
  ANDN U4347 ( .B(n2970), .A(n2971), .Z(n2968) );
  AND U4348 ( .A(a[91]), .B(b[8]), .Z(n2967) );
  XOR U4349 ( .A(n2972), .B(n2871), .Z(n2873) );
  IV U4350 ( .A(n2925), .Z(n2871) );
  XOR U4351 ( .A(n2973), .B(n2974), .Z(n2925) );
  ANDN U4352 ( .B(n2975), .A(n2976), .Z(n2973) );
  AND U4353 ( .A(a[92]), .B(b[7]), .Z(n2972) );
  XOR U4354 ( .A(n2977), .B(n2876), .Z(n2878) );
  IV U4355 ( .A(n2923), .Z(n2876) );
  XOR U4356 ( .A(n2978), .B(n2979), .Z(n2923) );
  ANDN U4357 ( .B(n2980), .A(n2981), .Z(n2978) );
  AND U4358 ( .A(a[93]), .B(b[6]), .Z(n2977) );
  XOR U4359 ( .A(n2982), .B(n2881), .Z(n2883) );
  IV U4360 ( .A(n2921), .Z(n2881) );
  XOR U4361 ( .A(n2983), .B(n2984), .Z(n2921) );
  ANDN U4362 ( .B(n2985), .A(n2986), .Z(n2983) );
  AND U4363 ( .A(a[94]), .B(b[5]), .Z(n2982) );
  XOR U4364 ( .A(n2987), .B(n2886), .Z(n2888) );
  IV U4365 ( .A(n2919), .Z(n2886) );
  XOR U4366 ( .A(n2988), .B(n2989), .Z(n2919) );
  ANDN U4367 ( .B(n2990), .A(n2991), .Z(n2988) );
  AND U4368 ( .A(a[95]), .B(b[4]), .Z(n2987) );
  XOR U4369 ( .A(n2992), .B(n2891), .Z(n2893) );
  IV U4370 ( .A(n2917), .Z(n2891) );
  XOR U4371 ( .A(n2993), .B(n2994), .Z(n2917) );
  ANDN U4372 ( .B(n2912), .A(n2913), .Z(n2993) );
  AND U4373 ( .A(a[96]), .B(b[2]), .Z(n2995) );
  XNOR U4374 ( .A(n2990), .B(n2994), .Z(n2996) );
  XOR U4375 ( .A(n2997), .B(n2998), .Z(n2994) );
  NANDN U4376 ( .A(n2915), .B(n2914), .Z(n2998) );
  XOR U4377 ( .A(n2997), .B(n2999), .Z(n2914) );
  NAND U4378 ( .A(a[96]), .B(b[1]), .Z(n2999) );
  XOR U4379 ( .A(n2997), .B(n3001), .Z(n3000) );
  OR U4380 ( .A(n2417), .B(n2415), .Z(n2997) );
  XOR U4381 ( .A(n3003), .B(n3004), .Z(n2415) );
  NANDN U4382 ( .A(n179), .B(a[96]), .Z(n2417) );
  XNOR U4383 ( .A(n2985), .B(n2989), .Z(n3005) );
  XNOR U4384 ( .A(n2980), .B(n2984), .Z(n3006) );
  XNOR U4385 ( .A(n2975), .B(n2979), .Z(n3007) );
  XNOR U4386 ( .A(n2970), .B(n2974), .Z(n3008) );
  XNOR U4387 ( .A(n2965), .B(n2969), .Z(n3009) );
  XNOR U4388 ( .A(n2960), .B(n2964), .Z(n3010) );
  XNOR U4389 ( .A(n2955), .B(n2959), .Z(n3011) );
  XNOR U4390 ( .A(n2950), .B(n2954), .Z(n3012) );
  XOR U4391 ( .A(n2946), .B(n2949), .Z(n3013) );
  XOR U4392 ( .A(n3014), .B(n3015), .Z(n2946) );
  XNOR U4393 ( .A(n3016), .B(n3017), .Z(n3015) );
  XNOR U4394 ( .A(n3018), .B(n3019), .Z(n3016) );
  XOR U4395 ( .A(n3020), .B(n3021), .Z(n3019) );
  AND U4396 ( .A(b[14]), .B(a[84]), .Z(n3021) );
  AND U4397 ( .A(a[83]), .B(b[15]), .Z(n3020) );
  XNOR U4398 ( .A(n3022), .B(n3018), .Z(n3014) );
  XOR U4399 ( .A(n3023), .B(n3024), .Z(n3018) );
  NOR U4400 ( .A(n3025), .B(n3026), .Z(n3023) );
  AND U4401 ( .A(a[85]), .B(b[13]), .Z(n3022) );
  XOR U4402 ( .A(n3027), .B(n2944), .Z(n2945) );
  IV U4403 ( .A(n3017), .Z(n2944) );
  XOR U4404 ( .A(n3028), .B(n3029), .Z(n3017) );
  ANDN U4405 ( .B(n3030), .A(n3031), .Z(n3028) );
  AND U4406 ( .A(a[86]), .B(b[12]), .Z(n3027) );
  XOR U4407 ( .A(n3033), .B(n3034), .Z(n2949) );
  ANDN U4408 ( .B(n3035), .A(n3036), .Z(n3033) );
  AND U4409 ( .A(a[87]), .B(b[11]), .Z(n3032) );
  XOR U4410 ( .A(n3038), .B(n3039), .Z(n2954) );
  ANDN U4411 ( .B(n3040), .A(n3041), .Z(n3038) );
  AND U4412 ( .A(a[88]), .B(b[10]), .Z(n3037) );
  XOR U4413 ( .A(n3043), .B(n3044), .Z(n2959) );
  ANDN U4414 ( .B(n3045), .A(n3046), .Z(n3043) );
  AND U4415 ( .A(a[89]), .B(b[9]), .Z(n3042) );
  XOR U4416 ( .A(n3048), .B(n3049), .Z(n2964) );
  ANDN U4417 ( .B(n3050), .A(n3051), .Z(n3048) );
  AND U4418 ( .A(a[90]), .B(b[8]), .Z(n3047) );
  XOR U4419 ( .A(n3053), .B(n3054), .Z(n2969) );
  ANDN U4420 ( .B(n3055), .A(n3056), .Z(n3053) );
  AND U4421 ( .A(a[91]), .B(b[7]), .Z(n3052) );
  XOR U4422 ( .A(n3058), .B(n3059), .Z(n2974) );
  ANDN U4423 ( .B(n3060), .A(n3061), .Z(n3058) );
  AND U4424 ( .A(a[92]), .B(b[6]), .Z(n3057) );
  XOR U4425 ( .A(n3063), .B(n3064), .Z(n2979) );
  ANDN U4426 ( .B(n3065), .A(n3066), .Z(n3063) );
  AND U4427 ( .A(a[93]), .B(b[5]), .Z(n3062) );
  XOR U4428 ( .A(n3068), .B(n3069), .Z(n2984) );
  ANDN U4429 ( .B(n3070), .A(n3071), .Z(n3068) );
  AND U4430 ( .A(a[94]), .B(b[4]), .Z(n3067) );
  XOR U4431 ( .A(n3073), .B(n3074), .Z(n2989) );
  ANDN U4432 ( .B(n3001), .A(n3002), .Z(n3073) );
  AND U4433 ( .A(a[95]), .B(b[2]), .Z(n3075) );
  XNOR U4434 ( .A(n3070), .B(n3074), .Z(n3076) );
  XOR U4435 ( .A(n3077), .B(n3078), .Z(n3074) );
  NANDN U4436 ( .A(n3004), .B(n3003), .Z(n3078) );
  XOR U4437 ( .A(n3077), .B(n3079), .Z(n3003) );
  NAND U4438 ( .A(a[95]), .B(b[1]), .Z(n3079) );
  XOR U4439 ( .A(n3077), .B(n3081), .Z(n3080) );
  OR U4440 ( .A(n2422), .B(n2420), .Z(n3077) );
  XOR U4441 ( .A(n3083), .B(n3084), .Z(n2420) );
  NANDN U4442 ( .A(n179), .B(a[95]), .Z(n2422) );
  XNOR U4443 ( .A(n3065), .B(n3069), .Z(n3085) );
  XNOR U4444 ( .A(n3060), .B(n3064), .Z(n3086) );
  XNOR U4445 ( .A(n3055), .B(n3059), .Z(n3087) );
  XNOR U4446 ( .A(n3050), .B(n3054), .Z(n3088) );
  XNOR U4447 ( .A(n3045), .B(n3049), .Z(n3089) );
  XNOR U4448 ( .A(n3040), .B(n3044), .Z(n3090) );
  XNOR U4449 ( .A(n3035), .B(n3039), .Z(n3091) );
  XNOR U4450 ( .A(n3030), .B(n3034), .Z(n3092) );
  XOR U4451 ( .A(n3026), .B(n3029), .Z(n3093) );
  XOR U4452 ( .A(n3094), .B(n3095), .Z(n3026) );
  XNOR U4453 ( .A(n3096), .B(n3097), .Z(n3095) );
  XOR U4454 ( .A(n3098), .B(n3099), .Z(n3096) );
  AND U4455 ( .A(b[13]), .B(a[84]), .Z(n3098) );
  XOR U4456 ( .A(n3099), .B(n3100), .Z(n3094) );
  XOR U4457 ( .A(n3101), .B(n3102), .Z(n3100) );
  AND U4458 ( .A(a[83]), .B(b[14]), .Z(n3102) );
  AND U4459 ( .A(a[82]), .B(b[15]), .Z(n3101) );
  XOR U4460 ( .A(n3103), .B(n3104), .Z(n3099) );
  ANDN U4461 ( .B(n3105), .A(n3106), .Z(n3103) );
  XOR U4462 ( .A(n3107), .B(n3024), .Z(n3025) );
  IV U4463 ( .A(n3097), .Z(n3024) );
  XOR U4464 ( .A(n3108), .B(n3109), .Z(n3097) );
  NOR U4465 ( .A(n3110), .B(n3111), .Z(n3108) );
  AND U4466 ( .A(a[85]), .B(b[12]), .Z(n3107) );
  XOR U4467 ( .A(n3113), .B(n3114), .Z(n3029) );
  ANDN U4468 ( .B(n3115), .A(n3116), .Z(n3113) );
  AND U4469 ( .A(a[86]), .B(b[11]), .Z(n3112) );
  XOR U4470 ( .A(n3118), .B(n3119), .Z(n3034) );
  ANDN U4471 ( .B(n3120), .A(n3121), .Z(n3118) );
  AND U4472 ( .A(a[87]), .B(b[10]), .Z(n3117) );
  XOR U4473 ( .A(n3123), .B(n3124), .Z(n3039) );
  ANDN U4474 ( .B(n3125), .A(n3126), .Z(n3123) );
  AND U4475 ( .A(a[88]), .B(b[9]), .Z(n3122) );
  XOR U4476 ( .A(n3128), .B(n3129), .Z(n3044) );
  ANDN U4477 ( .B(n3130), .A(n3131), .Z(n3128) );
  AND U4478 ( .A(a[89]), .B(b[8]), .Z(n3127) );
  XOR U4479 ( .A(n3133), .B(n3134), .Z(n3049) );
  ANDN U4480 ( .B(n3135), .A(n3136), .Z(n3133) );
  AND U4481 ( .A(a[90]), .B(b[7]), .Z(n3132) );
  XOR U4482 ( .A(n3138), .B(n3139), .Z(n3054) );
  ANDN U4483 ( .B(n3140), .A(n3141), .Z(n3138) );
  AND U4484 ( .A(a[91]), .B(b[6]), .Z(n3137) );
  XOR U4485 ( .A(n3143), .B(n3144), .Z(n3059) );
  ANDN U4486 ( .B(n3145), .A(n3146), .Z(n3143) );
  AND U4487 ( .A(a[92]), .B(b[5]), .Z(n3142) );
  XOR U4488 ( .A(n3148), .B(n3149), .Z(n3064) );
  ANDN U4489 ( .B(n3150), .A(n3151), .Z(n3148) );
  AND U4490 ( .A(a[93]), .B(b[4]), .Z(n3147) );
  XOR U4491 ( .A(n3153), .B(n3154), .Z(n3069) );
  ANDN U4492 ( .B(n3081), .A(n3082), .Z(n3153) );
  AND U4493 ( .A(a[94]), .B(b[2]), .Z(n3155) );
  XNOR U4494 ( .A(n3150), .B(n3154), .Z(n3156) );
  XOR U4495 ( .A(n3157), .B(n3158), .Z(n3154) );
  NANDN U4496 ( .A(n3084), .B(n3083), .Z(n3158) );
  XOR U4497 ( .A(n3157), .B(n3159), .Z(n3083) );
  NAND U4498 ( .A(a[94]), .B(b[1]), .Z(n3159) );
  XOR U4499 ( .A(n3157), .B(n3161), .Z(n3160) );
  OR U4500 ( .A(n2427), .B(n2425), .Z(n3157) );
  XOR U4501 ( .A(n3163), .B(n3164), .Z(n2425) );
  NANDN U4502 ( .A(n179), .B(a[94]), .Z(n2427) );
  XNOR U4503 ( .A(n3145), .B(n3149), .Z(n3165) );
  XNOR U4504 ( .A(n3140), .B(n3144), .Z(n3166) );
  XNOR U4505 ( .A(n3135), .B(n3139), .Z(n3167) );
  XNOR U4506 ( .A(n3130), .B(n3134), .Z(n3168) );
  XNOR U4507 ( .A(n3125), .B(n3129), .Z(n3169) );
  XNOR U4508 ( .A(n3120), .B(n3124), .Z(n3170) );
  XNOR U4509 ( .A(n3115), .B(n3119), .Z(n3171) );
  XOR U4510 ( .A(n3111), .B(n3114), .Z(n3172) );
  XNOR U4511 ( .A(n3106), .B(n3173), .Z(n3111) );
  XNOR U4512 ( .A(n3105), .B(n3109), .Z(n3173) );
  XOR U4513 ( .A(n3174), .B(n3104), .Z(n3105) );
  AND U4514 ( .A(b[12]), .B(a[84]), .Z(n3174) );
  XOR U4515 ( .A(n3175), .B(n3176), .Z(n3106) );
  XOR U4516 ( .A(n3104), .B(n3177), .Z(n3176) );
  XOR U4517 ( .A(n3178), .B(n3179), .Z(n3177) );
  XOR U4518 ( .A(n3180), .B(n3181), .Z(n3179) );
  NAND U4519 ( .A(a[82]), .B(b[14]), .Z(n3181) );
  AND U4520 ( .A(a[81]), .B(b[15]), .Z(n3180) );
  XOR U4521 ( .A(n3182), .B(n3183), .Z(n3104) );
  ANDN U4522 ( .B(n3184), .A(n3185), .Z(n3182) );
  XOR U4523 ( .A(n3186), .B(n3178), .Z(n3175) );
  XOR U4524 ( .A(n3187), .B(n3188), .Z(n3178) );
  NOR U4525 ( .A(n3189), .B(n3190), .Z(n3187) );
  AND U4526 ( .A(a[83]), .B(b[13]), .Z(n3186) );
  XOR U4527 ( .A(n3192), .B(n3193), .Z(n3109) );
  ANDN U4528 ( .B(n3194), .A(n3195), .Z(n3192) );
  AND U4529 ( .A(a[85]), .B(b[11]), .Z(n3191) );
  XOR U4530 ( .A(n3197), .B(n3198), .Z(n3114) );
  ANDN U4531 ( .B(n3199), .A(n3200), .Z(n3197) );
  AND U4532 ( .A(a[86]), .B(b[10]), .Z(n3196) );
  XOR U4533 ( .A(n3202), .B(n3203), .Z(n3119) );
  ANDN U4534 ( .B(n3204), .A(n3205), .Z(n3202) );
  AND U4535 ( .A(a[87]), .B(b[9]), .Z(n3201) );
  XOR U4536 ( .A(n3207), .B(n3208), .Z(n3124) );
  ANDN U4537 ( .B(n3209), .A(n3210), .Z(n3207) );
  AND U4538 ( .A(a[88]), .B(b[8]), .Z(n3206) );
  XOR U4539 ( .A(n3212), .B(n3213), .Z(n3129) );
  ANDN U4540 ( .B(n3214), .A(n3215), .Z(n3212) );
  AND U4541 ( .A(a[89]), .B(b[7]), .Z(n3211) );
  XOR U4542 ( .A(n3217), .B(n3218), .Z(n3134) );
  ANDN U4543 ( .B(n3219), .A(n3220), .Z(n3217) );
  AND U4544 ( .A(a[90]), .B(b[6]), .Z(n3216) );
  XOR U4545 ( .A(n3222), .B(n3223), .Z(n3139) );
  ANDN U4546 ( .B(n3224), .A(n3225), .Z(n3222) );
  AND U4547 ( .A(a[91]), .B(b[5]), .Z(n3221) );
  XOR U4548 ( .A(n3227), .B(n3228), .Z(n3144) );
  ANDN U4549 ( .B(n3229), .A(n3230), .Z(n3227) );
  AND U4550 ( .A(a[92]), .B(b[4]), .Z(n3226) );
  XOR U4551 ( .A(n3232), .B(n3233), .Z(n3149) );
  ANDN U4552 ( .B(n3161), .A(n3162), .Z(n3232) );
  AND U4553 ( .A(a[93]), .B(b[2]), .Z(n3234) );
  XNOR U4554 ( .A(n3229), .B(n3233), .Z(n3235) );
  XOR U4555 ( .A(n3236), .B(n3237), .Z(n3233) );
  NANDN U4556 ( .A(n3164), .B(n3163), .Z(n3237) );
  XOR U4557 ( .A(n3236), .B(n3238), .Z(n3163) );
  NAND U4558 ( .A(a[93]), .B(b[1]), .Z(n3238) );
  XOR U4559 ( .A(n3236), .B(n3240), .Z(n3239) );
  OR U4560 ( .A(n2432), .B(n2430), .Z(n3236) );
  XOR U4561 ( .A(n3242), .B(n3243), .Z(n2430) );
  NANDN U4562 ( .A(n179), .B(a[93]), .Z(n2432) );
  XNOR U4563 ( .A(n3224), .B(n3228), .Z(n3244) );
  XNOR U4564 ( .A(n3219), .B(n3223), .Z(n3245) );
  XNOR U4565 ( .A(n3214), .B(n3218), .Z(n3246) );
  XNOR U4566 ( .A(n3209), .B(n3213), .Z(n3247) );
  XNOR U4567 ( .A(n3204), .B(n3208), .Z(n3248) );
  XNOR U4568 ( .A(n3199), .B(n3203), .Z(n3249) );
  XNOR U4569 ( .A(n3194), .B(n3198), .Z(n3250) );
  XNOR U4570 ( .A(n3184), .B(n3193), .Z(n3251) );
  XOR U4571 ( .A(n3252), .B(n3183), .Z(n3184) );
  AND U4572 ( .A(b[11]), .B(a[84]), .Z(n3252) );
  XOR U4573 ( .A(n3183), .B(n3190), .Z(n3253) );
  XOR U4574 ( .A(n3254), .B(n3255), .Z(n3190) );
  XOR U4575 ( .A(n3188), .B(n3256), .Z(n3255) );
  XOR U4576 ( .A(n3257), .B(n3258), .Z(n3256) );
  XOR U4577 ( .A(n3259), .B(n3260), .Z(n3258) );
  NAND U4578 ( .A(a[81]), .B(b[14]), .Z(n3260) );
  AND U4579 ( .A(a[80]), .B(b[15]), .Z(n3259) );
  XOR U4580 ( .A(n3261), .B(n3257), .Z(n3254) );
  XOR U4581 ( .A(n3262), .B(n3263), .Z(n3257) );
  NOR U4582 ( .A(n3264), .B(n3265), .Z(n3262) );
  AND U4583 ( .A(a[82]), .B(b[13]), .Z(n3261) );
  XOR U4584 ( .A(n3266), .B(n3267), .Z(n3183) );
  ANDN U4585 ( .B(n3268), .A(n3269), .Z(n3266) );
  XNOR U4586 ( .A(n3270), .B(n3188), .Z(n3189) );
  XOR U4587 ( .A(n3271), .B(n3272), .Z(n3188) );
  ANDN U4588 ( .B(n3273), .A(n3274), .Z(n3271) );
  AND U4589 ( .A(a[83]), .B(b[12]), .Z(n3270) );
  XOR U4590 ( .A(n3276), .B(n3277), .Z(n3193) );
  ANDN U4591 ( .B(n3278), .A(n3279), .Z(n3276) );
  AND U4592 ( .A(a[85]), .B(b[10]), .Z(n3275) );
  XOR U4593 ( .A(n3281), .B(n3282), .Z(n3198) );
  ANDN U4594 ( .B(n3283), .A(n3284), .Z(n3281) );
  AND U4595 ( .A(a[86]), .B(b[9]), .Z(n3280) );
  XOR U4596 ( .A(n3286), .B(n3287), .Z(n3203) );
  ANDN U4597 ( .B(n3288), .A(n3289), .Z(n3286) );
  AND U4598 ( .A(a[87]), .B(b[8]), .Z(n3285) );
  XOR U4599 ( .A(n3291), .B(n3292), .Z(n3208) );
  ANDN U4600 ( .B(n3293), .A(n3294), .Z(n3291) );
  AND U4601 ( .A(a[88]), .B(b[7]), .Z(n3290) );
  XOR U4602 ( .A(n3296), .B(n3297), .Z(n3213) );
  ANDN U4603 ( .B(n3298), .A(n3299), .Z(n3296) );
  AND U4604 ( .A(a[89]), .B(b[6]), .Z(n3295) );
  XOR U4605 ( .A(n3301), .B(n3302), .Z(n3218) );
  ANDN U4606 ( .B(n3303), .A(n3304), .Z(n3301) );
  AND U4607 ( .A(a[90]), .B(b[5]), .Z(n3300) );
  XOR U4608 ( .A(n3306), .B(n3307), .Z(n3223) );
  ANDN U4609 ( .B(n3308), .A(n3309), .Z(n3306) );
  AND U4610 ( .A(a[91]), .B(b[4]), .Z(n3305) );
  XOR U4611 ( .A(n3311), .B(n3312), .Z(n3228) );
  ANDN U4612 ( .B(n3240), .A(n3241), .Z(n3311) );
  AND U4613 ( .A(a[92]), .B(b[2]), .Z(n3313) );
  XNOR U4614 ( .A(n3308), .B(n3312), .Z(n3314) );
  XOR U4615 ( .A(n3315), .B(n3316), .Z(n3312) );
  NANDN U4616 ( .A(n3243), .B(n3242), .Z(n3316) );
  XOR U4617 ( .A(n3315), .B(n3317), .Z(n3242) );
  NAND U4618 ( .A(a[92]), .B(b[1]), .Z(n3317) );
  XOR U4619 ( .A(n3315), .B(n3319), .Z(n3318) );
  OR U4620 ( .A(n2437), .B(n2435), .Z(n3315) );
  XOR U4621 ( .A(n3321), .B(n3322), .Z(n2435) );
  NANDN U4622 ( .A(n179), .B(a[92]), .Z(n2437) );
  XNOR U4623 ( .A(n3303), .B(n3307), .Z(n3323) );
  XNOR U4624 ( .A(n3298), .B(n3302), .Z(n3324) );
  XNOR U4625 ( .A(n3293), .B(n3297), .Z(n3325) );
  XNOR U4626 ( .A(n3288), .B(n3292), .Z(n3326) );
  XNOR U4627 ( .A(n3283), .B(n3287), .Z(n3327) );
  XNOR U4628 ( .A(n3278), .B(n3282), .Z(n3328) );
  XNOR U4629 ( .A(n3268), .B(n3277), .Z(n3329) );
  XOR U4630 ( .A(n3330), .B(n3267), .Z(n3268) );
  AND U4631 ( .A(b[10]), .B(a[84]), .Z(n3330) );
  XNOR U4632 ( .A(n3267), .B(n3273), .Z(n3331) );
  XOR U4633 ( .A(n3272), .B(n3265), .Z(n3332) );
  XOR U4634 ( .A(n3333), .B(n3334), .Z(n3265) );
  XOR U4635 ( .A(n3263), .B(n3335), .Z(n3334) );
  XOR U4636 ( .A(n3336), .B(n3337), .Z(n3335) );
  XOR U4637 ( .A(n3338), .B(n3339), .Z(n3337) );
  NAND U4638 ( .A(a[80]), .B(b[14]), .Z(n3339) );
  AND U4639 ( .A(a[79]), .B(b[15]), .Z(n3338) );
  XOR U4640 ( .A(n3340), .B(n3336), .Z(n3333) );
  XOR U4641 ( .A(n3341), .B(n3342), .Z(n3336) );
  NOR U4642 ( .A(n3343), .B(n3344), .Z(n3341) );
  AND U4643 ( .A(a[81]), .B(b[13]), .Z(n3340) );
  XNOR U4644 ( .A(n3345), .B(n3263), .Z(n3264) );
  XOR U4645 ( .A(n3346), .B(n3347), .Z(n3263) );
  ANDN U4646 ( .B(n3348), .A(n3349), .Z(n3346) );
  AND U4647 ( .A(a[82]), .B(b[12]), .Z(n3345) );
  XOR U4648 ( .A(n3350), .B(n3351), .Z(n3267) );
  ANDN U4649 ( .B(n3352), .A(n3353), .Z(n3350) );
  XNOR U4650 ( .A(n3354), .B(n3272), .Z(n3274) );
  XOR U4651 ( .A(n3355), .B(n3356), .Z(n3272) );
  ANDN U4652 ( .B(n3357), .A(n3358), .Z(n3355) );
  AND U4653 ( .A(a[83]), .B(b[11]), .Z(n3354) );
  XOR U4654 ( .A(n3360), .B(n3361), .Z(n3277) );
  ANDN U4655 ( .B(n3362), .A(n3363), .Z(n3360) );
  AND U4656 ( .A(a[85]), .B(b[9]), .Z(n3359) );
  XOR U4657 ( .A(n3365), .B(n3366), .Z(n3282) );
  ANDN U4658 ( .B(n3367), .A(n3368), .Z(n3365) );
  AND U4659 ( .A(a[86]), .B(b[8]), .Z(n3364) );
  XOR U4660 ( .A(n3370), .B(n3371), .Z(n3287) );
  ANDN U4661 ( .B(n3372), .A(n3373), .Z(n3370) );
  AND U4662 ( .A(a[87]), .B(b[7]), .Z(n3369) );
  XOR U4663 ( .A(n3375), .B(n3376), .Z(n3292) );
  ANDN U4664 ( .B(n3377), .A(n3378), .Z(n3375) );
  AND U4665 ( .A(a[88]), .B(b[6]), .Z(n3374) );
  XOR U4666 ( .A(n3380), .B(n3381), .Z(n3297) );
  ANDN U4667 ( .B(n3382), .A(n3383), .Z(n3380) );
  AND U4668 ( .A(a[89]), .B(b[5]), .Z(n3379) );
  XOR U4669 ( .A(n3385), .B(n3386), .Z(n3302) );
  ANDN U4670 ( .B(n3387), .A(n3388), .Z(n3385) );
  AND U4671 ( .A(a[90]), .B(b[4]), .Z(n3384) );
  XOR U4672 ( .A(n3390), .B(n3391), .Z(n3307) );
  ANDN U4673 ( .B(n3319), .A(n3320), .Z(n3390) );
  AND U4674 ( .A(a[91]), .B(b[2]), .Z(n3392) );
  XNOR U4675 ( .A(n3387), .B(n3391), .Z(n3393) );
  XOR U4676 ( .A(n3394), .B(n3395), .Z(n3391) );
  NANDN U4677 ( .A(n3322), .B(n3321), .Z(n3395) );
  XOR U4678 ( .A(n3394), .B(n3396), .Z(n3321) );
  NAND U4679 ( .A(a[91]), .B(b[1]), .Z(n3396) );
  XOR U4680 ( .A(n3394), .B(n3398), .Z(n3397) );
  OR U4681 ( .A(n2442), .B(n2440), .Z(n3394) );
  XOR U4682 ( .A(n3400), .B(n3401), .Z(n2440) );
  NANDN U4683 ( .A(n179), .B(a[91]), .Z(n2442) );
  XNOR U4684 ( .A(n3382), .B(n3386), .Z(n3402) );
  XNOR U4685 ( .A(n3377), .B(n3381), .Z(n3403) );
  XNOR U4686 ( .A(n3372), .B(n3376), .Z(n3404) );
  XNOR U4687 ( .A(n3367), .B(n3371), .Z(n3405) );
  XNOR U4688 ( .A(n3362), .B(n3366), .Z(n3406) );
  XNOR U4689 ( .A(n3352), .B(n3361), .Z(n3407) );
  XOR U4690 ( .A(n3408), .B(n3351), .Z(n3352) );
  AND U4691 ( .A(b[9]), .B(a[84]), .Z(n3408) );
  XNOR U4692 ( .A(n3351), .B(n3357), .Z(n3409) );
  XNOR U4693 ( .A(n3356), .B(n3348), .Z(n3410) );
  XOR U4694 ( .A(n3347), .B(n3344), .Z(n3411) );
  XOR U4695 ( .A(n3412), .B(n3413), .Z(n3344) );
  XOR U4696 ( .A(n3342), .B(n3414), .Z(n3413) );
  XOR U4697 ( .A(n3415), .B(n3416), .Z(n3414) );
  XOR U4698 ( .A(n3417), .B(n3418), .Z(n3416) );
  NAND U4699 ( .A(a[79]), .B(b[14]), .Z(n3418) );
  AND U4700 ( .A(a[78]), .B(b[15]), .Z(n3417) );
  XOR U4701 ( .A(n3419), .B(n3415), .Z(n3412) );
  XOR U4702 ( .A(n3420), .B(n3421), .Z(n3415) );
  NOR U4703 ( .A(n3422), .B(n3423), .Z(n3420) );
  AND U4704 ( .A(a[80]), .B(b[13]), .Z(n3419) );
  XNOR U4705 ( .A(n3424), .B(n3342), .Z(n3343) );
  XOR U4706 ( .A(n3425), .B(n3426), .Z(n3342) );
  ANDN U4707 ( .B(n3427), .A(n3428), .Z(n3425) );
  AND U4708 ( .A(a[81]), .B(b[12]), .Z(n3424) );
  XNOR U4709 ( .A(n3429), .B(n3347), .Z(n3349) );
  XOR U4710 ( .A(n3430), .B(n3431), .Z(n3347) );
  ANDN U4711 ( .B(n3432), .A(n3433), .Z(n3430) );
  AND U4712 ( .A(a[82]), .B(b[11]), .Z(n3429) );
  XOR U4713 ( .A(n3434), .B(n3435), .Z(n3351) );
  ANDN U4714 ( .B(n3436), .A(n3437), .Z(n3434) );
  XNOR U4715 ( .A(n3438), .B(n3356), .Z(n3358) );
  XOR U4716 ( .A(n3439), .B(n3440), .Z(n3356) );
  ANDN U4717 ( .B(n3441), .A(n3442), .Z(n3439) );
  AND U4718 ( .A(a[83]), .B(b[10]), .Z(n3438) );
  XOR U4719 ( .A(n3444), .B(n3445), .Z(n3361) );
  ANDN U4720 ( .B(n3446), .A(n3447), .Z(n3444) );
  AND U4721 ( .A(a[85]), .B(b[8]), .Z(n3443) );
  XOR U4722 ( .A(n3449), .B(n3450), .Z(n3366) );
  ANDN U4723 ( .B(n3451), .A(n3452), .Z(n3449) );
  AND U4724 ( .A(a[86]), .B(b[7]), .Z(n3448) );
  XOR U4725 ( .A(n3454), .B(n3455), .Z(n3371) );
  ANDN U4726 ( .B(n3456), .A(n3457), .Z(n3454) );
  AND U4727 ( .A(a[87]), .B(b[6]), .Z(n3453) );
  XOR U4728 ( .A(n3459), .B(n3460), .Z(n3376) );
  ANDN U4729 ( .B(n3461), .A(n3462), .Z(n3459) );
  AND U4730 ( .A(a[88]), .B(b[5]), .Z(n3458) );
  XOR U4731 ( .A(n3464), .B(n3465), .Z(n3381) );
  ANDN U4732 ( .B(n3466), .A(n3467), .Z(n3464) );
  AND U4733 ( .A(a[89]), .B(b[4]), .Z(n3463) );
  XOR U4734 ( .A(n3469), .B(n3470), .Z(n3386) );
  ANDN U4735 ( .B(n3398), .A(n3399), .Z(n3469) );
  AND U4736 ( .A(a[90]), .B(b[2]), .Z(n3471) );
  XNOR U4737 ( .A(n3466), .B(n3470), .Z(n3472) );
  XOR U4738 ( .A(n3473), .B(n3474), .Z(n3470) );
  NANDN U4739 ( .A(n3401), .B(n3400), .Z(n3474) );
  XOR U4740 ( .A(n3473), .B(n3475), .Z(n3400) );
  NAND U4741 ( .A(a[90]), .B(b[1]), .Z(n3475) );
  XOR U4742 ( .A(n3473), .B(n3477), .Z(n3476) );
  OR U4743 ( .A(n2447), .B(n2445), .Z(n3473) );
  XOR U4744 ( .A(n3479), .B(n3480), .Z(n2445) );
  NANDN U4745 ( .A(n179), .B(a[90]), .Z(n2447) );
  XNOR U4746 ( .A(n3461), .B(n3465), .Z(n3481) );
  XNOR U4747 ( .A(n3456), .B(n3460), .Z(n3482) );
  XNOR U4748 ( .A(n3451), .B(n3455), .Z(n3483) );
  XNOR U4749 ( .A(n3446), .B(n3450), .Z(n3484) );
  XNOR U4750 ( .A(n3436), .B(n3445), .Z(n3485) );
  XOR U4751 ( .A(n3486), .B(n3435), .Z(n3436) );
  AND U4752 ( .A(b[8]), .B(a[84]), .Z(n3486) );
  XNOR U4753 ( .A(n3435), .B(n3441), .Z(n3487) );
  XNOR U4754 ( .A(n3440), .B(n3432), .Z(n3488) );
  XNOR U4755 ( .A(n3431), .B(n3427), .Z(n3489) );
  XOR U4756 ( .A(n3426), .B(n3423), .Z(n3490) );
  XOR U4757 ( .A(n3491), .B(n3492), .Z(n3423) );
  XOR U4758 ( .A(n3421), .B(n3493), .Z(n3492) );
  XOR U4759 ( .A(n3494), .B(n3495), .Z(n3493) );
  XOR U4760 ( .A(n3496), .B(n3497), .Z(n3495) );
  NAND U4761 ( .A(a[78]), .B(b[14]), .Z(n3497) );
  AND U4762 ( .A(a[77]), .B(b[15]), .Z(n3496) );
  XOR U4763 ( .A(n3498), .B(n3494), .Z(n3491) );
  XOR U4764 ( .A(n3499), .B(n3500), .Z(n3494) );
  NOR U4765 ( .A(n3501), .B(n3502), .Z(n3499) );
  AND U4766 ( .A(a[79]), .B(b[13]), .Z(n3498) );
  XNOR U4767 ( .A(n3503), .B(n3421), .Z(n3422) );
  XOR U4768 ( .A(n3504), .B(n3505), .Z(n3421) );
  ANDN U4769 ( .B(n3506), .A(n3507), .Z(n3504) );
  AND U4770 ( .A(a[80]), .B(b[12]), .Z(n3503) );
  XNOR U4771 ( .A(n3508), .B(n3426), .Z(n3428) );
  XOR U4772 ( .A(n3509), .B(n3510), .Z(n3426) );
  ANDN U4773 ( .B(n3511), .A(n3512), .Z(n3509) );
  AND U4774 ( .A(a[81]), .B(b[11]), .Z(n3508) );
  XNOR U4775 ( .A(n3513), .B(n3431), .Z(n3433) );
  XOR U4776 ( .A(n3514), .B(n3515), .Z(n3431) );
  ANDN U4777 ( .B(n3516), .A(n3517), .Z(n3514) );
  AND U4778 ( .A(a[82]), .B(b[10]), .Z(n3513) );
  XOR U4779 ( .A(n3518), .B(n3519), .Z(n3435) );
  ANDN U4780 ( .B(n3520), .A(n3521), .Z(n3518) );
  XNOR U4781 ( .A(n3522), .B(n3440), .Z(n3442) );
  XOR U4782 ( .A(n3523), .B(n3524), .Z(n3440) );
  ANDN U4783 ( .B(n3525), .A(n3526), .Z(n3523) );
  AND U4784 ( .A(a[83]), .B(b[9]), .Z(n3522) );
  XOR U4785 ( .A(n3528), .B(n3529), .Z(n3445) );
  ANDN U4786 ( .B(n3530), .A(n3531), .Z(n3528) );
  AND U4787 ( .A(a[85]), .B(b[7]), .Z(n3527) );
  XOR U4788 ( .A(n3533), .B(n3534), .Z(n3450) );
  ANDN U4789 ( .B(n3535), .A(n3536), .Z(n3533) );
  AND U4790 ( .A(a[86]), .B(b[6]), .Z(n3532) );
  XOR U4791 ( .A(n3538), .B(n3539), .Z(n3455) );
  ANDN U4792 ( .B(n3540), .A(n3541), .Z(n3538) );
  AND U4793 ( .A(a[87]), .B(b[5]), .Z(n3537) );
  XOR U4794 ( .A(n3543), .B(n3544), .Z(n3460) );
  ANDN U4795 ( .B(n3545), .A(n3546), .Z(n3543) );
  AND U4796 ( .A(a[88]), .B(b[4]), .Z(n3542) );
  XOR U4797 ( .A(n3548), .B(n3549), .Z(n3465) );
  ANDN U4798 ( .B(n3477), .A(n3478), .Z(n3548) );
  AND U4799 ( .A(a[89]), .B(b[2]), .Z(n3550) );
  XNOR U4800 ( .A(n3545), .B(n3549), .Z(n3551) );
  XOR U4801 ( .A(n3552), .B(n3553), .Z(n3549) );
  NANDN U4802 ( .A(n3480), .B(n3479), .Z(n3553) );
  XOR U4803 ( .A(n3552), .B(n3554), .Z(n3479) );
  NAND U4804 ( .A(a[89]), .B(b[1]), .Z(n3554) );
  XOR U4805 ( .A(n3552), .B(n3556), .Z(n3555) );
  OR U4806 ( .A(n2452), .B(n2450), .Z(n3552) );
  XOR U4807 ( .A(n3558), .B(n3559), .Z(n2450) );
  NANDN U4808 ( .A(n179), .B(a[89]), .Z(n2452) );
  XNOR U4809 ( .A(n3540), .B(n3544), .Z(n3560) );
  XNOR U4810 ( .A(n3535), .B(n3539), .Z(n3561) );
  XNOR U4811 ( .A(n3530), .B(n3534), .Z(n3562) );
  XNOR U4812 ( .A(n3520), .B(n3529), .Z(n3563) );
  XOR U4813 ( .A(n3564), .B(n3519), .Z(n3520) );
  AND U4814 ( .A(b[7]), .B(a[84]), .Z(n3564) );
  XNOR U4815 ( .A(n3519), .B(n3525), .Z(n3565) );
  XNOR U4816 ( .A(n3524), .B(n3516), .Z(n3566) );
  XNOR U4817 ( .A(n3515), .B(n3511), .Z(n3567) );
  XNOR U4818 ( .A(n3510), .B(n3506), .Z(n3568) );
  XOR U4819 ( .A(n3505), .B(n3502), .Z(n3569) );
  XOR U4820 ( .A(n3570), .B(n3571), .Z(n3502) );
  XOR U4821 ( .A(n3500), .B(n3572), .Z(n3571) );
  XOR U4822 ( .A(n3573), .B(n3574), .Z(n3572) );
  XOR U4823 ( .A(n3575), .B(n3576), .Z(n3574) );
  NAND U4824 ( .A(a[77]), .B(b[14]), .Z(n3576) );
  AND U4825 ( .A(a[76]), .B(b[15]), .Z(n3575) );
  XOR U4826 ( .A(n3577), .B(n3573), .Z(n3570) );
  XOR U4827 ( .A(n3578), .B(n3579), .Z(n3573) );
  NOR U4828 ( .A(n3580), .B(n3581), .Z(n3578) );
  AND U4829 ( .A(a[78]), .B(b[13]), .Z(n3577) );
  XNOR U4830 ( .A(n3582), .B(n3500), .Z(n3501) );
  XOR U4831 ( .A(n3583), .B(n3584), .Z(n3500) );
  ANDN U4832 ( .B(n3585), .A(n3586), .Z(n3583) );
  AND U4833 ( .A(a[79]), .B(b[12]), .Z(n3582) );
  XNOR U4834 ( .A(n3587), .B(n3505), .Z(n3507) );
  XOR U4835 ( .A(n3588), .B(n3589), .Z(n3505) );
  ANDN U4836 ( .B(n3590), .A(n3591), .Z(n3588) );
  AND U4837 ( .A(a[80]), .B(b[11]), .Z(n3587) );
  XNOR U4838 ( .A(n3592), .B(n3510), .Z(n3512) );
  XOR U4839 ( .A(n3593), .B(n3594), .Z(n3510) );
  ANDN U4840 ( .B(n3595), .A(n3596), .Z(n3593) );
  AND U4841 ( .A(a[81]), .B(b[10]), .Z(n3592) );
  XNOR U4842 ( .A(n3597), .B(n3515), .Z(n3517) );
  XOR U4843 ( .A(n3598), .B(n3599), .Z(n3515) );
  ANDN U4844 ( .B(n3600), .A(n3601), .Z(n3598) );
  AND U4845 ( .A(a[82]), .B(b[9]), .Z(n3597) );
  XOR U4846 ( .A(n3602), .B(n3603), .Z(n3519) );
  ANDN U4847 ( .B(n3604), .A(n3605), .Z(n3602) );
  XNOR U4848 ( .A(n3606), .B(n3524), .Z(n3526) );
  XOR U4849 ( .A(n3607), .B(n3608), .Z(n3524) );
  ANDN U4850 ( .B(n3609), .A(n3610), .Z(n3607) );
  AND U4851 ( .A(a[83]), .B(b[8]), .Z(n3606) );
  XOR U4852 ( .A(n3612), .B(n3613), .Z(n3529) );
  ANDN U4853 ( .B(n3614), .A(n3615), .Z(n3612) );
  AND U4854 ( .A(a[85]), .B(b[6]), .Z(n3611) );
  XOR U4855 ( .A(n3617), .B(n3618), .Z(n3534) );
  ANDN U4856 ( .B(n3619), .A(n3620), .Z(n3617) );
  AND U4857 ( .A(a[86]), .B(b[5]), .Z(n3616) );
  XOR U4858 ( .A(n3622), .B(n3623), .Z(n3539) );
  ANDN U4859 ( .B(n3624), .A(n3625), .Z(n3622) );
  AND U4860 ( .A(a[87]), .B(b[4]), .Z(n3621) );
  XOR U4861 ( .A(n3627), .B(n3628), .Z(n3544) );
  ANDN U4862 ( .B(n3556), .A(n3557), .Z(n3627) );
  AND U4863 ( .A(a[88]), .B(b[2]), .Z(n3629) );
  XNOR U4864 ( .A(n3624), .B(n3628), .Z(n3630) );
  XOR U4865 ( .A(n3631), .B(n3632), .Z(n3628) );
  NANDN U4866 ( .A(n3559), .B(n3558), .Z(n3632) );
  XOR U4867 ( .A(n3631), .B(n3633), .Z(n3558) );
  NAND U4868 ( .A(a[88]), .B(b[1]), .Z(n3633) );
  XOR U4869 ( .A(n3631), .B(n3635), .Z(n3634) );
  OR U4870 ( .A(n2457), .B(n2455), .Z(n3631) );
  XOR U4871 ( .A(n3637), .B(n3638), .Z(n2455) );
  NANDN U4872 ( .A(n179), .B(a[88]), .Z(n2457) );
  XNOR U4873 ( .A(n3619), .B(n3623), .Z(n3639) );
  XNOR U4874 ( .A(n3614), .B(n3618), .Z(n3640) );
  XNOR U4875 ( .A(n3604), .B(n3613), .Z(n3641) );
  XOR U4876 ( .A(n3642), .B(n3603), .Z(n3604) );
  AND U4877 ( .A(b[6]), .B(a[84]), .Z(n3642) );
  XNOR U4878 ( .A(n3603), .B(n3609), .Z(n3643) );
  XNOR U4879 ( .A(n3608), .B(n3600), .Z(n3644) );
  XNOR U4880 ( .A(n3599), .B(n3595), .Z(n3645) );
  XNOR U4881 ( .A(n3594), .B(n3590), .Z(n3646) );
  XNOR U4882 ( .A(n3589), .B(n3585), .Z(n3647) );
  XOR U4883 ( .A(n3584), .B(n3581), .Z(n3648) );
  XOR U4884 ( .A(n3649), .B(n3650), .Z(n3581) );
  XOR U4885 ( .A(n3579), .B(n3651), .Z(n3650) );
  XOR U4886 ( .A(n3652), .B(n3653), .Z(n3651) );
  XOR U4887 ( .A(n3654), .B(n3655), .Z(n3653) );
  NAND U4888 ( .A(a[76]), .B(b[14]), .Z(n3655) );
  AND U4889 ( .A(a[75]), .B(b[15]), .Z(n3654) );
  XOR U4890 ( .A(n3656), .B(n3652), .Z(n3649) );
  XOR U4891 ( .A(n3657), .B(n3658), .Z(n3652) );
  NOR U4892 ( .A(n3659), .B(n3660), .Z(n3657) );
  AND U4893 ( .A(a[77]), .B(b[13]), .Z(n3656) );
  XNOR U4894 ( .A(n3661), .B(n3579), .Z(n3580) );
  XOR U4895 ( .A(n3662), .B(n3663), .Z(n3579) );
  ANDN U4896 ( .B(n3664), .A(n3665), .Z(n3662) );
  AND U4897 ( .A(a[78]), .B(b[12]), .Z(n3661) );
  XNOR U4898 ( .A(n3666), .B(n3584), .Z(n3586) );
  XOR U4899 ( .A(n3667), .B(n3668), .Z(n3584) );
  ANDN U4900 ( .B(n3669), .A(n3670), .Z(n3667) );
  AND U4901 ( .A(a[79]), .B(b[11]), .Z(n3666) );
  XNOR U4902 ( .A(n3671), .B(n3589), .Z(n3591) );
  XOR U4903 ( .A(n3672), .B(n3673), .Z(n3589) );
  ANDN U4904 ( .B(n3674), .A(n3675), .Z(n3672) );
  AND U4905 ( .A(a[80]), .B(b[10]), .Z(n3671) );
  XNOR U4906 ( .A(n3676), .B(n3594), .Z(n3596) );
  XOR U4907 ( .A(n3677), .B(n3678), .Z(n3594) );
  ANDN U4908 ( .B(n3679), .A(n3680), .Z(n3677) );
  AND U4909 ( .A(a[81]), .B(b[9]), .Z(n3676) );
  XNOR U4910 ( .A(n3681), .B(n3599), .Z(n3601) );
  XOR U4911 ( .A(n3682), .B(n3683), .Z(n3599) );
  ANDN U4912 ( .B(n3684), .A(n3685), .Z(n3682) );
  AND U4913 ( .A(a[82]), .B(b[8]), .Z(n3681) );
  XOR U4914 ( .A(n3686), .B(n3687), .Z(n3603) );
  ANDN U4915 ( .B(n3688), .A(n3689), .Z(n3686) );
  XNOR U4916 ( .A(n3690), .B(n3608), .Z(n3610) );
  XOR U4917 ( .A(n3691), .B(n3692), .Z(n3608) );
  ANDN U4918 ( .B(n3693), .A(n3694), .Z(n3691) );
  AND U4919 ( .A(a[83]), .B(b[7]), .Z(n3690) );
  XOR U4920 ( .A(n3696), .B(n3697), .Z(n3613) );
  ANDN U4921 ( .B(n3698), .A(n3699), .Z(n3696) );
  AND U4922 ( .A(a[85]), .B(b[5]), .Z(n3695) );
  XOR U4923 ( .A(n3701), .B(n3702), .Z(n3618) );
  ANDN U4924 ( .B(n3703), .A(n3704), .Z(n3701) );
  AND U4925 ( .A(a[86]), .B(b[4]), .Z(n3700) );
  XOR U4926 ( .A(n3706), .B(n3707), .Z(n3623) );
  ANDN U4927 ( .B(n3635), .A(n3636), .Z(n3706) );
  AND U4928 ( .A(a[87]), .B(b[2]), .Z(n3708) );
  XNOR U4929 ( .A(n3703), .B(n3707), .Z(n3709) );
  XOR U4930 ( .A(n3710), .B(n3711), .Z(n3707) );
  NANDN U4931 ( .A(n3638), .B(n3637), .Z(n3711) );
  XOR U4932 ( .A(n3710), .B(n3712), .Z(n3637) );
  NAND U4933 ( .A(a[87]), .B(b[1]), .Z(n3712) );
  XOR U4934 ( .A(n3710), .B(n3714), .Z(n3713) );
  OR U4935 ( .A(n2462), .B(n2460), .Z(n3710) );
  XOR U4936 ( .A(n3716), .B(n3717), .Z(n2460) );
  NANDN U4937 ( .A(n179), .B(a[87]), .Z(n2462) );
  XNOR U4938 ( .A(n3698), .B(n3702), .Z(n3718) );
  XNOR U4939 ( .A(n3688), .B(n3697), .Z(n3719) );
  XOR U4940 ( .A(n3720), .B(n3687), .Z(n3688) );
  AND U4941 ( .A(b[5]), .B(a[84]), .Z(n3720) );
  XNOR U4942 ( .A(n3687), .B(n3693), .Z(n3721) );
  XNOR U4943 ( .A(n3692), .B(n3684), .Z(n3722) );
  XNOR U4944 ( .A(n3683), .B(n3679), .Z(n3723) );
  XNOR U4945 ( .A(n3678), .B(n3674), .Z(n3724) );
  XNOR U4946 ( .A(n3673), .B(n3669), .Z(n3725) );
  XNOR U4947 ( .A(n3668), .B(n3664), .Z(n3726) );
  XOR U4948 ( .A(n3663), .B(n3660), .Z(n3727) );
  XOR U4949 ( .A(n3728), .B(n3729), .Z(n3660) );
  XOR U4950 ( .A(n3658), .B(n3730), .Z(n3729) );
  XOR U4951 ( .A(n3731), .B(n3732), .Z(n3730) );
  XOR U4952 ( .A(n3733), .B(n3734), .Z(n3732) );
  NAND U4953 ( .A(a[75]), .B(b[14]), .Z(n3734) );
  AND U4954 ( .A(a[74]), .B(b[15]), .Z(n3733) );
  XOR U4955 ( .A(n3735), .B(n3731), .Z(n3728) );
  XOR U4956 ( .A(n3736), .B(n3737), .Z(n3731) );
  NOR U4957 ( .A(n3738), .B(n3739), .Z(n3736) );
  AND U4958 ( .A(a[76]), .B(b[13]), .Z(n3735) );
  XNOR U4959 ( .A(n3740), .B(n3658), .Z(n3659) );
  XOR U4960 ( .A(n3741), .B(n3742), .Z(n3658) );
  ANDN U4961 ( .B(n3743), .A(n3744), .Z(n3741) );
  AND U4962 ( .A(a[77]), .B(b[12]), .Z(n3740) );
  XNOR U4963 ( .A(n3745), .B(n3663), .Z(n3665) );
  XOR U4964 ( .A(n3746), .B(n3747), .Z(n3663) );
  ANDN U4965 ( .B(n3748), .A(n3749), .Z(n3746) );
  AND U4966 ( .A(a[78]), .B(b[11]), .Z(n3745) );
  XNOR U4967 ( .A(n3750), .B(n3668), .Z(n3670) );
  XOR U4968 ( .A(n3751), .B(n3752), .Z(n3668) );
  ANDN U4969 ( .B(n3753), .A(n3754), .Z(n3751) );
  AND U4970 ( .A(a[79]), .B(b[10]), .Z(n3750) );
  XNOR U4971 ( .A(n3755), .B(n3673), .Z(n3675) );
  XOR U4972 ( .A(n3756), .B(n3757), .Z(n3673) );
  ANDN U4973 ( .B(n3758), .A(n3759), .Z(n3756) );
  AND U4974 ( .A(a[80]), .B(b[9]), .Z(n3755) );
  XNOR U4975 ( .A(n3760), .B(n3678), .Z(n3680) );
  XOR U4976 ( .A(n3761), .B(n3762), .Z(n3678) );
  ANDN U4977 ( .B(n3763), .A(n3764), .Z(n3761) );
  AND U4978 ( .A(a[81]), .B(b[8]), .Z(n3760) );
  XNOR U4979 ( .A(n3765), .B(n3683), .Z(n3685) );
  XOR U4980 ( .A(n3766), .B(n3767), .Z(n3683) );
  ANDN U4981 ( .B(n3768), .A(n3769), .Z(n3766) );
  AND U4982 ( .A(a[82]), .B(b[7]), .Z(n3765) );
  XOR U4983 ( .A(n3770), .B(n3771), .Z(n3687) );
  ANDN U4984 ( .B(n3772), .A(n3773), .Z(n3770) );
  XNOR U4985 ( .A(n3774), .B(n3692), .Z(n3694) );
  XOR U4986 ( .A(n3775), .B(n3776), .Z(n3692) );
  ANDN U4987 ( .B(n3777), .A(n3778), .Z(n3775) );
  AND U4988 ( .A(a[83]), .B(b[6]), .Z(n3774) );
  XOR U4989 ( .A(n3780), .B(n3781), .Z(n3697) );
  ANDN U4990 ( .B(n3782), .A(n3783), .Z(n3780) );
  AND U4991 ( .A(a[85]), .B(b[4]), .Z(n3779) );
  XOR U4992 ( .A(n3785), .B(n3786), .Z(n3702) );
  ANDN U4993 ( .B(n3714), .A(n3715), .Z(n3785) );
  AND U4994 ( .A(a[86]), .B(b[2]), .Z(n3787) );
  XNOR U4995 ( .A(n3782), .B(n3786), .Z(n3788) );
  XOR U4996 ( .A(n3789), .B(n3790), .Z(n3786) );
  NANDN U4997 ( .A(n3717), .B(n3716), .Z(n3790) );
  XOR U4998 ( .A(n3789), .B(n3791), .Z(n3716) );
  NAND U4999 ( .A(a[86]), .B(b[1]), .Z(n3791) );
  XOR U5000 ( .A(n3789), .B(n3793), .Z(n3792) );
  OR U5001 ( .A(n2467), .B(n2465), .Z(n3789) );
  XOR U5002 ( .A(n3795), .B(n3796), .Z(n2465) );
  NANDN U5003 ( .A(n179), .B(a[86]), .Z(n2467) );
  XNOR U5004 ( .A(n3772), .B(n3781), .Z(n3797) );
  XOR U5005 ( .A(n3798), .B(n3771), .Z(n3772) );
  AND U5006 ( .A(b[4]), .B(a[84]), .Z(n3798) );
  XNOR U5007 ( .A(n3771), .B(n3777), .Z(n3799) );
  XNOR U5008 ( .A(n3776), .B(n3768), .Z(n3800) );
  XNOR U5009 ( .A(n3767), .B(n3763), .Z(n3801) );
  XNOR U5010 ( .A(n3762), .B(n3758), .Z(n3802) );
  XNOR U5011 ( .A(n3757), .B(n3753), .Z(n3803) );
  XNOR U5012 ( .A(n3752), .B(n3748), .Z(n3804) );
  XNOR U5013 ( .A(n3747), .B(n3743), .Z(n3805) );
  XOR U5014 ( .A(n3742), .B(n3739), .Z(n3806) );
  XOR U5015 ( .A(n3807), .B(n3808), .Z(n3739) );
  XOR U5016 ( .A(n3737), .B(n3809), .Z(n3808) );
  XOR U5017 ( .A(n3810), .B(n3811), .Z(n3809) );
  XOR U5018 ( .A(n3812), .B(n3813), .Z(n3811) );
  NAND U5019 ( .A(a[74]), .B(b[14]), .Z(n3813) );
  AND U5020 ( .A(a[73]), .B(b[15]), .Z(n3812) );
  XOR U5021 ( .A(n3814), .B(n3810), .Z(n3807) );
  XOR U5022 ( .A(n3815), .B(n3816), .Z(n3810) );
  NOR U5023 ( .A(n3817), .B(n3818), .Z(n3815) );
  AND U5024 ( .A(a[75]), .B(b[13]), .Z(n3814) );
  XNOR U5025 ( .A(n3819), .B(n3737), .Z(n3738) );
  XOR U5026 ( .A(n3820), .B(n3821), .Z(n3737) );
  ANDN U5027 ( .B(n3822), .A(n3823), .Z(n3820) );
  AND U5028 ( .A(a[76]), .B(b[12]), .Z(n3819) );
  XNOR U5029 ( .A(n3824), .B(n3742), .Z(n3744) );
  XOR U5030 ( .A(n3825), .B(n3826), .Z(n3742) );
  ANDN U5031 ( .B(n3827), .A(n3828), .Z(n3825) );
  AND U5032 ( .A(a[77]), .B(b[11]), .Z(n3824) );
  XNOR U5033 ( .A(n3829), .B(n3747), .Z(n3749) );
  XOR U5034 ( .A(n3830), .B(n3831), .Z(n3747) );
  ANDN U5035 ( .B(n3832), .A(n3833), .Z(n3830) );
  AND U5036 ( .A(a[78]), .B(b[10]), .Z(n3829) );
  XNOR U5037 ( .A(n3834), .B(n3752), .Z(n3754) );
  XOR U5038 ( .A(n3835), .B(n3836), .Z(n3752) );
  ANDN U5039 ( .B(n3837), .A(n3838), .Z(n3835) );
  AND U5040 ( .A(a[79]), .B(b[9]), .Z(n3834) );
  XNOR U5041 ( .A(n3839), .B(n3757), .Z(n3759) );
  XOR U5042 ( .A(n3840), .B(n3841), .Z(n3757) );
  ANDN U5043 ( .B(n3842), .A(n3843), .Z(n3840) );
  AND U5044 ( .A(a[80]), .B(b[8]), .Z(n3839) );
  XNOR U5045 ( .A(n3844), .B(n3762), .Z(n3764) );
  XOR U5046 ( .A(n3845), .B(n3846), .Z(n3762) );
  ANDN U5047 ( .B(n3847), .A(n3848), .Z(n3845) );
  AND U5048 ( .A(a[81]), .B(b[7]), .Z(n3844) );
  XNOR U5049 ( .A(n3849), .B(n3767), .Z(n3769) );
  XOR U5050 ( .A(n3850), .B(n3851), .Z(n3767) );
  ANDN U5051 ( .B(n3852), .A(n3853), .Z(n3850) );
  AND U5052 ( .A(a[82]), .B(b[6]), .Z(n3849) );
  XOR U5053 ( .A(n3854), .B(n3855), .Z(n3771) );
  ANDN U5054 ( .B(n3856), .A(n3857), .Z(n3854) );
  XNOR U5055 ( .A(n3858), .B(n3776), .Z(n3778) );
  XOR U5056 ( .A(n3859), .B(n3860), .Z(n3776) );
  ANDN U5057 ( .B(n3861), .A(n3862), .Z(n3859) );
  AND U5058 ( .A(a[83]), .B(b[5]), .Z(n3858) );
  XOR U5059 ( .A(n3864), .B(n3865), .Z(n3781) );
  ANDN U5060 ( .B(n3793), .A(n3794), .Z(n3864) );
  AND U5061 ( .A(a[85]), .B(b[2]), .Z(n3866) );
  XNOR U5062 ( .A(n3856), .B(n3865), .Z(n3867) );
  XOR U5063 ( .A(n3868), .B(n3869), .Z(n3865) );
  NANDN U5064 ( .A(n3796), .B(n3795), .Z(n3869) );
  XOR U5065 ( .A(n3868), .B(n3870), .Z(n3795) );
  NAND U5066 ( .A(a[85]), .B(b[1]), .Z(n3870) );
  XNOR U5067 ( .A(n3868), .B(n3872), .Z(n3871) );
  OR U5068 ( .A(n2472), .B(n2470), .Z(n3868) );
  NANDN U5069 ( .A(n179), .B(a[85]), .Z(n2472) );
  XOR U5070 ( .A(n3876), .B(n3855), .Z(n3856) );
  AND U5071 ( .A(b[3]), .B(a[84]), .Z(n3876) );
  XNOR U5072 ( .A(n3855), .B(n3861), .Z(n3877) );
  XNOR U5073 ( .A(n3860), .B(n3852), .Z(n3878) );
  XNOR U5074 ( .A(n3851), .B(n3847), .Z(n3879) );
  XNOR U5075 ( .A(n3846), .B(n3842), .Z(n3880) );
  XNOR U5076 ( .A(n3841), .B(n3837), .Z(n3881) );
  XNOR U5077 ( .A(n3836), .B(n3832), .Z(n3882) );
  XNOR U5078 ( .A(n3831), .B(n3827), .Z(n3883) );
  XNOR U5079 ( .A(n3826), .B(n3822), .Z(n3884) );
  XOR U5080 ( .A(n3821), .B(n3818), .Z(n3885) );
  XOR U5081 ( .A(n3886), .B(n3887), .Z(n3818) );
  XOR U5082 ( .A(n3816), .B(n3888), .Z(n3887) );
  XOR U5083 ( .A(n3889), .B(n3890), .Z(n3888) );
  XOR U5084 ( .A(n3891), .B(n3892), .Z(n3890) );
  NAND U5085 ( .A(a[73]), .B(b[14]), .Z(n3892) );
  AND U5086 ( .A(a[72]), .B(b[15]), .Z(n3891) );
  XOR U5087 ( .A(n3893), .B(n3889), .Z(n3886) );
  XOR U5088 ( .A(n3894), .B(n3895), .Z(n3889) );
  NOR U5089 ( .A(n3896), .B(n3897), .Z(n3894) );
  AND U5090 ( .A(a[74]), .B(b[13]), .Z(n3893) );
  XNOR U5091 ( .A(n3898), .B(n3816), .Z(n3817) );
  XOR U5092 ( .A(n3899), .B(n3900), .Z(n3816) );
  ANDN U5093 ( .B(n3901), .A(n3902), .Z(n3899) );
  AND U5094 ( .A(a[75]), .B(b[12]), .Z(n3898) );
  XNOR U5095 ( .A(n3903), .B(n3821), .Z(n3823) );
  XOR U5096 ( .A(n3904), .B(n3905), .Z(n3821) );
  ANDN U5097 ( .B(n3906), .A(n3907), .Z(n3904) );
  AND U5098 ( .A(a[76]), .B(b[11]), .Z(n3903) );
  XNOR U5099 ( .A(n3908), .B(n3826), .Z(n3828) );
  XOR U5100 ( .A(n3909), .B(n3910), .Z(n3826) );
  ANDN U5101 ( .B(n3911), .A(n3912), .Z(n3909) );
  AND U5102 ( .A(a[77]), .B(b[10]), .Z(n3908) );
  XNOR U5103 ( .A(n3913), .B(n3831), .Z(n3833) );
  XOR U5104 ( .A(n3914), .B(n3915), .Z(n3831) );
  ANDN U5105 ( .B(n3916), .A(n3917), .Z(n3914) );
  AND U5106 ( .A(a[78]), .B(b[9]), .Z(n3913) );
  XNOR U5107 ( .A(n3918), .B(n3836), .Z(n3838) );
  XOR U5108 ( .A(n3919), .B(n3920), .Z(n3836) );
  ANDN U5109 ( .B(n3921), .A(n3922), .Z(n3919) );
  AND U5110 ( .A(a[79]), .B(b[8]), .Z(n3918) );
  XNOR U5111 ( .A(n3923), .B(n3841), .Z(n3843) );
  XOR U5112 ( .A(n3924), .B(n3925), .Z(n3841) );
  ANDN U5113 ( .B(n3926), .A(n3927), .Z(n3924) );
  AND U5114 ( .A(a[80]), .B(b[7]), .Z(n3923) );
  XNOR U5115 ( .A(n3928), .B(n3846), .Z(n3848) );
  XOR U5116 ( .A(n3929), .B(n3930), .Z(n3846) );
  ANDN U5117 ( .B(n3931), .A(n3932), .Z(n3929) );
  AND U5118 ( .A(a[81]), .B(b[6]), .Z(n3928) );
  XNOR U5119 ( .A(n3933), .B(n3851), .Z(n3853) );
  XOR U5120 ( .A(n3934), .B(n3935), .Z(n3851) );
  ANDN U5121 ( .B(n3936), .A(n3937), .Z(n3934) );
  AND U5122 ( .A(a[82]), .B(b[5]), .Z(n3933) );
  XNOR U5123 ( .A(n3938), .B(n3939), .Z(n3855) );
  NOR U5124 ( .A(n3873), .B(n3872), .Z(n3938) );
  XOR U5125 ( .A(n3940), .B(n3939), .Z(n3872) );
  AND U5126 ( .A(b[2]), .B(a[84]), .Z(n3940) );
  XOR U5127 ( .A(n3939), .B(n3942), .Z(n3941) );
  XNOR U5128 ( .A(n3943), .B(n3944), .Z(n3939) );
  OR U5129 ( .A(n3874), .B(n3875), .Z(n3944) );
  XNOR U5130 ( .A(n3943), .B(n3946), .Z(n3945) );
  XNOR U5131 ( .A(n3943), .B(n3948), .Z(n3874) );
  NAND U5132 ( .A(b[1]), .B(a[84]), .Z(n3948) );
  OR U5133 ( .A(n2477), .B(n2475), .Z(n3943) );
  XOR U5134 ( .A(n3949), .B(n3950), .Z(n2475) );
  NANDN U5135 ( .A(n179), .B(a[84]), .Z(n2477) );
  XNOR U5136 ( .A(n3952), .B(n3860), .Z(n3862) );
  XOR U5137 ( .A(n3953), .B(n3954), .Z(n3860) );
  ANDN U5138 ( .B(n3942), .A(n3951), .Z(n3953) );
  XNOR U5139 ( .A(n3955), .B(n3954), .Z(n3951) );
  AND U5140 ( .A(a[83]), .B(b[3]), .Z(n3955) );
  XNOR U5141 ( .A(n3954), .B(n3936), .Z(n3956) );
  XNOR U5142 ( .A(n3935), .B(n3931), .Z(n3957) );
  XNOR U5143 ( .A(n3930), .B(n3926), .Z(n3958) );
  XNOR U5144 ( .A(n3925), .B(n3921), .Z(n3959) );
  XNOR U5145 ( .A(n3920), .B(n3916), .Z(n3960) );
  XNOR U5146 ( .A(n3915), .B(n3911), .Z(n3961) );
  XNOR U5147 ( .A(n3910), .B(n3906), .Z(n3962) );
  XNOR U5148 ( .A(n3905), .B(n3901), .Z(n3963) );
  XOR U5149 ( .A(n3900), .B(n3897), .Z(n3964) );
  XOR U5150 ( .A(n3965), .B(n3966), .Z(n3897) );
  XOR U5151 ( .A(n3895), .B(n3967), .Z(n3966) );
  XOR U5152 ( .A(n3968), .B(n3969), .Z(n3967) );
  XOR U5153 ( .A(n3970), .B(n3971), .Z(n3969) );
  NAND U5154 ( .A(a[72]), .B(b[14]), .Z(n3971) );
  AND U5155 ( .A(a[71]), .B(b[15]), .Z(n3970) );
  XOR U5156 ( .A(n3972), .B(n3968), .Z(n3965) );
  XOR U5157 ( .A(n3973), .B(n3974), .Z(n3968) );
  NOR U5158 ( .A(n3975), .B(n3976), .Z(n3973) );
  AND U5159 ( .A(a[73]), .B(b[13]), .Z(n3972) );
  XNOR U5160 ( .A(n3977), .B(n3895), .Z(n3896) );
  XOR U5161 ( .A(n3978), .B(n3979), .Z(n3895) );
  ANDN U5162 ( .B(n3980), .A(n3981), .Z(n3978) );
  AND U5163 ( .A(a[74]), .B(b[12]), .Z(n3977) );
  XNOR U5164 ( .A(n3982), .B(n3900), .Z(n3902) );
  XOR U5165 ( .A(n3983), .B(n3984), .Z(n3900) );
  ANDN U5166 ( .B(n3985), .A(n3986), .Z(n3983) );
  AND U5167 ( .A(a[75]), .B(b[11]), .Z(n3982) );
  XNOR U5168 ( .A(n3987), .B(n3905), .Z(n3907) );
  XOR U5169 ( .A(n3988), .B(n3989), .Z(n3905) );
  ANDN U5170 ( .B(n3990), .A(n3991), .Z(n3988) );
  AND U5171 ( .A(a[76]), .B(b[10]), .Z(n3987) );
  XNOR U5172 ( .A(n3992), .B(n3910), .Z(n3912) );
  XOR U5173 ( .A(n3993), .B(n3994), .Z(n3910) );
  ANDN U5174 ( .B(n3995), .A(n3996), .Z(n3993) );
  AND U5175 ( .A(a[77]), .B(b[9]), .Z(n3992) );
  XNOR U5176 ( .A(n3997), .B(n3915), .Z(n3917) );
  XOR U5177 ( .A(n3998), .B(n3999), .Z(n3915) );
  ANDN U5178 ( .B(n4000), .A(n4001), .Z(n3998) );
  AND U5179 ( .A(a[78]), .B(b[8]), .Z(n3997) );
  XNOR U5180 ( .A(n4002), .B(n3920), .Z(n3922) );
  XOR U5181 ( .A(n4003), .B(n4004), .Z(n3920) );
  ANDN U5182 ( .B(n4005), .A(n4006), .Z(n4003) );
  AND U5183 ( .A(a[79]), .B(b[7]), .Z(n4002) );
  XNOR U5184 ( .A(n4007), .B(n3925), .Z(n3927) );
  XOR U5185 ( .A(n4008), .B(n4009), .Z(n3925) );
  ANDN U5186 ( .B(n4010), .A(n4011), .Z(n4008) );
  AND U5187 ( .A(a[80]), .B(b[6]), .Z(n4007) );
  XNOR U5188 ( .A(n4012), .B(n3930), .Z(n3932) );
  XOR U5189 ( .A(n4013), .B(n4014), .Z(n3930) );
  ANDN U5190 ( .B(n4015), .A(n4016), .Z(n4013) );
  AND U5191 ( .A(a[81]), .B(b[5]), .Z(n4012) );
  XNOR U5192 ( .A(n4017), .B(n4018), .Z(n3954) );
  NOR U5193 ( .A(n3947), .B(n3946), .Z(n4017) );
  XOR U5194 ( .A(n4019), .B(n4018), .Z(n3946) );
  AND U5195 ( .A(a[83]), .B(b[2]), .Z(n4019) );
  XOR U5196 ( .A(n4018), .B(n4021), .Z(n4020) );
  XNOR U5197 ( .A(n4022), .B(n4023), .Z(n4018) );
  NANDN U5198 ( .A(n3950), .B(n3949), .Z(n4023) );
  XOR U5199 ( .A(n4022), .B(n4024), .Z(n3949) );
  NAND U5200 ( .A(a[83]), .B(b[1]), .Z(n4024) );
  XOR U5201 ( .A(n4022), .B(n4026), .Z(n4025) );
  OR U5202 ( .A(n2482), .B(n2480), .Z(n4022) );
  XOR U5203 ( .A(n4028), .B(n4029), .Z(n2480) );
  NANDN U5204 ( .A(n179), .B(a[83]), .Z(n2482) );
  XNOR U5205 ( .A(n4031), .B(n3935), .Z(n3937) );
  XOR U5206 ( .A(n4032), .B(n4033), .Z(n3935) );
  ANDN U5207 ( .B(n4021), .A(n4030), .Z(n4032) );
  XNOR U5208 ( .A(n4034), .B(n4033), .Z(n4030) );
  AND U5209 ( .A(a[82]), .B(b[3]), .Z(n4034) );
  XNOR U5210 ( .A(n4033), .B(n4015), .Z(n4035) );
  XNOR U5211 ( .A(n4014), .B(n4010), .Z(n4036) );
  XNOR U5212 ( .A(n4009), .B(n4005), .Z(n4037) );
  XNOR U5213 ( .A(n4004), .B(n4000), .Z(n4038) );
  XNOR U5214 ( .A(n3999), .B(n3995), .Z(n4039) );
  XNOR U5215 ( .A(n3994), .B(n3990), .Z(n4040) );
  XNOR U5216 ( .A(n3989), .B(n3985), .Z(n4041) );
  XNOR U5217 ( .A(n3984), .B(n3980), .Z(n4042) );
  XOR U5218 ( .A(n3979), .B(n3976), .Z(n4043) );
  XOR U5219 ( .A(n4044), .B(n4045), .Z(n3976) );
  XOR U5220 ( .A(n3974), .B(n4046), .Z(n4045) );
  XNOR U5221 ( .A(n4047), .B(n4048), .Z(n4046) );
  XOR U5222 ( .A(n4049), .B(n4050), .Z(n4048) );
  NAND U5223 ( .A(a[71]), .B(b[14]), .Z(n4050) );
  AND U5224 ( .A(a[70]), .B(b[15]), .Z(n4049) );
  XNOR U5225 ( .A(n4051), .B(n4047), .Z(n4044) );
  XOR U5226 ( .A(n4052), .B(n4053), .Z(n4047) );
  NOR U5227 ( .A(n4054), .B(n4055), .Z(n4052) );
  AND U5228 ( .A(a[72]), .B(b[13]), .Z(n4051) );
  XNOR U5229 ( .A(n4056), .B(n3974), .Z(n3975) );
  XNOR U5230 ( .A(n4057), .B(n4058), .Z(n3974) );
  ANDN U5231 ( .B(n4059), .A(n4060), .Z(n4057) );
  AND U5232 ( .A(a[73]), .B(b[12]), .Z(n4056) );
  XNOR U5233 ( .A(n4061), .B(n3979), .Z(n3981) );
  XNOR U5234 ( .A(n4062), .B(n4063), .Z(n3979) );
  ANDN U5235 ( .B(n4064), .A(n4065), .Z(n4062) );
  AND U5236 ( .A(a[74]), .B(b[11]), .Z(n4061) );
  XNOR U5237 ( .A(n4066), .B(n3984), .Z(n3986) );
  XNOR U5238 ( .A(n4067), .B(n4068), .Z(n3984) );
  ANDN U5239 ( .B(n4069), .A(n4070), .Z(n4067) );
  AND U5240 ( .A(a[75]), .B(b[10]), .Z(n4066) );
  XNOR U5241 ( .A(n4071), .B(n3989), .Z(n3991) );
  XNOR U5242 ( .A(n4072), .B(n4073), .Z(n3989) );
  ANDN U5243 ( .B(n4074), .A(n4075), .Z(n4072) );
  AND U5244 ( .A(a[76]), .B(b[9]), .Z(n4071) );
  XNOR U5245 ( .A(n4076), .B(n3994), .Z(n3996) );
  XNOR U5246 ( .A(n4077), .B(n4078), .Z(n3994) );
  ANDN U5247 ( .B(n4079), .A(n4080), .Z(n4077) );
  AND U5248 ( .A(a[77]), .B(b[8]), .Z(n4076) );
  XNOR U5249 ( .A(n4081), .B(n3999), .Z(n4001) );
  XNOR U5250 ( .A(n4082), .B(n4083), .Z(n3999) );
  ANDN U5251 ( .B(n4084), .A(n4085), .Z(n4082) );
  AND U5252 ( .A(a[78]), .B(b[7]), .Z(n4081) );
  XNOR U5253 ( .A(n4086), .B(n4004), .Z(n4006) );
  XNOR U5254 ( .A(n4087), .B(n4088), .Z(n4004) );
  ANDN U5255 ( .B(n4089), .A(n4090), .Z(n4087) );
  AND U5256 ( .A(a[79]), .B(b[6]), .Z(n4086) );
  XNOR U5257 ( .A(n4091), .B(n4009), .Z(n4011) );
  XNOR U5258 ( .A(n4092), .B(n4093), .Z(n4009) );
  ANDN U5259 ( .B(n4094), .A(n4095), .Z(n4092) );
  AND U5260 ( .A(a[80]), .B(b[5]), .Z(n4091) );
  XNOR U5261 ( .A(n4096), .B(n4097), .Z(n4033) );
  ANDN U5262 ( .B(n4026), .A(n4027), .Z(n4096) );
  XOR U5263 ( .A(n4098), .B(n4097), .Z(n4027) );
  IV U5264 ( .A(n4099), .Z(n4097) );
  AND U5265 ( .A(b[2]), .B(a[82]), .Z(n4098) );
  XNOR U5266 ( .A(n4101), .B(n4099), .Z(n4100) );
  XOR U5267 ( .A(n4102), .B(n4103), .Z(n4099) );
  NANDN U5268 ( .A(n4029), .B(n4028), .Z(n4103) );
  XOR U5269 ( .A(n4102), .B(n4104), .Z(n4028) );
  NAND U5270 ( .A(a[82]), .B(b[1]), .Z(n4104) );
  XOR U5271 ( .A(n4102), .B(n4106), .Z(n4105) );
  OR U5272 ( .A(n2487), .B(n2485), .Z(n4102) );
  XOR U5273 ( .A(n4108), .B(n4109), .Z(n2485) );
  NANDN U5274 ( .A(n179), .B(a[82]), .Z(n2487) );
  XNOR U5275 ( .A(n4111), .B(n4014), .Z(n4016) );
  XNOR U5276 ( .A(n4112), .B(n4113), .Z(n4014) );
  ANDN U5277 ( .B(n4101), .A(n4110), .Z(n4112) );
  XOR U5278 ( .A(n4114), .B(n4113), .Z(n4110) );
  IV U5279 ( .A(n4115), .Z(n4113) );
  AND U5280 ( .A(a[81]), .B(b[3]), .Z(n4114) );
  XNOR U5281 ( .A(n4094), .B(n4115), .Z(n4116) );
  XOR U5282 ( .A(n4117), .B(n4118), .Z(n4115) );
  ANDN U5283 ( .B(n4106), .A(n4107), .Z(n4117) );
  AND U5284 ( .A(b[2]), .B(a[81]), .Z(n4119) );
  XNOR U5285 ( .A(n4121), .B(n4118), .Z(n4120) );
  XOR U5286 ( .A(n4122), .B(n4123), .Z(n4118) );
  NANDN U5287 ( .A(n4109), .B(n4108), .Z(n4123) );
  XOR U5288 ( .A(n4122), .B(n4124), .Z(n4108) );
  NAND U5289 ( .A(a[81]), .B(b[1]), .Z(n4124) );
  XOR U5290 ( .A(n4122), .B(n4126), .Z(n4125) );
  OR U5291 ( .A(n2492), .B(n2490), .Z(n4122) );
  XOR U5292 ( .A(n4128), .B(n4129), .Z(n2490) );
  NANDN U5293 ( .A(n179), .B(a[81]), .Z(n2492) );
  XNOR U5294 ( .A(n4089), .B(n4132), .Z(n4131) );
  XNOR U5295 ( .A(n4084), .B(n4134), .Z(n4133) );
  XNOR U5296 ( .A(n4079), .B(n4136), .Z(n4135) );
  XNOR U5297 ( .A(n4074), .B(n4138), .Z(n4137) );
  XNOR U5298 ( .A(n4069), .B(n4140), .Z(n4139) );
  XNOR U5299 ( .A(n4064), .B(n4142), .Z(n4141) );
  XNOR U5300 ( .A(n4059), .B(n4144), .Z(n4143) );
  XOR U5301 ( .A(n4055), .B(n4146), .Z(n4145) );
  XOR U5302 ( .A(n4147), .B(n4148), .Z(n4055) );
  XNOR U5303 ( .A(n4149), .B(n4150), .Z(n4148) );
  XNOR U5304 ( .A(n4151), .B(n4152), .Z(n4149) );
  XOR U5305 ( .A(n4153), .B(n4154), .Z(n4152) );
  AND U5306 ( .A(b[15]), .B(a[69]), .Z(n4154) );
  AND U5307 ( .A(a[70]), .B(b[14]), .Z(n4153) );
  XNOR U5308 ( .A(n4155), .B(n4151), .Z(n4147) );
  XOR U5309 ( .A(n4156), .B(n4157), .Z(n4151) );
  NOR U5310 ( .A(n4158), .B(n4159), .Z(n4156) );
  AND U5311 ( .A(a[71]), .B(b[13]), .Z(n4155) );
  XOR U5312 ( .A(n4160), .B(n4053), .Z(n4054) );
  IV U5313 ( .A(n4150), .Z(n4053) );
  XOR U5314 ( .A(n4161), .B(n4162), .Z(n4150) );
  ANDN U5315 ( .B(n4163), .A(n4164), .Z(n4161) );
  AND U5316 ( .A(a[72]), .B(b[12]), .Z(n4160) );
  XOR U5317 ( .A(n4165), .B(n4058), .Z(n4060) );
  IV U5318 ( .A(n4146), .Z(n4058) );
  XOR U5319 ( .A(n4166), .B(n4167), .Z(n4146) );
  ANDN U5320 ( .B(n4168), .A(n4169), .Z(n4166) );
  AND U5321 ( .A(a[73]), .B(b[11]), .Z(n4165) );
  XOR U5322 ( .A(n4170), .B(n4063), .Z(n4065) );
  IV U5323 ( .A(n4144), .Z(n4063) );
  XOR U5324 ( .A(n4171), .B(n4172), .Z(n4144) );
  ANDN U5325 ( .B(n4173), .A(n4174), .Z(n4171) );
  AND U5326 ( .A(a[74]), .B(b[10]), .Z(n4170) );
  XOR U5327 ( .A(n4175), .B(n4068), .Z(n4070) );
  IV U5328 ( .A(n4142), .Z(n4068) );
  XOR U5329 ( .A(n4176), .B(n4177), .Z(n4142) );
  ANDN U5330 ( .B(n4178), .A(n4179), .Z(n4176) );
  AND U5331 ( .A(a[75]), .B(b[9]), .Z(n4175) );
  XOR U5332 ( .A(n4180), .B(n4073), .Z(n4075) );
  IV U5333 ( .A(n4140), .Z(n4073) );
  XOR U5334 ( .A(n4181), .B(n4182), .Z(n4140) );
  ANDN U5335 ( .B(n4183), .A(n4184), .Z(n4181) );
  AND U5336 ( .A(a[76]), .B(b[8]), .Z(n4180) );
  XOR U5337 ( .A(n4185), .B(n4078), .Z(n4080) );
  IV U5338 ( .A(n4138), .Z(n4078) );
  XOR U5339 ( .A(n4186), .B(n4187), .Z(n4138) );
  ANDN U5340 ( .B(n4188), .A(n4189), .Z(n4186) );
  AND U5341 ( .A(a[77]), .B(b[7]), .Z(n4185) );
  XOR U5342 ( .A(n4190), .B(n4083), .Z(n4085) );
  IV U5343 ( .A(n4136), .Z(n4083) );
  XOR U5344 ( .A(n4191), .B(n4192), .Z(n4136) );
  ANDN U5345 ( .B(n4193), .A(n4194), .Z(n4191) );
  AND U5346 ( .A(a[78]), .B(b[6]), .Z(n4190) );
  XOR U5347 ( .A(n4195), .B(n4088), .Z(n4090) );
  IV U5348 ( .A(n4134), .Z(n4088) );
  XOR U5349 ( .A(n4196), .B(n4197), .Z(n4134) );
  ANDN U5350 ( .B(n4198), .A(n4199), .Z(n4196) );
  AND U5351 ( .A(a[79]), .B(b[5]), .Z(n4195) );
  XOR U5352 ( .A(n4200), .B(n4093), .Z(n4095) );
  IV U5353 ( .A(n4132), .Z(n4093) );
  XOR U5354 ( .A(n4201), .B(n4202), .Z(n4132) );
  ANDN U5355 ( .B(n4121), .A(n4130), .Z(n4201) );
  AND U5356 ( .A(a[80]), .B(b[3]), .Z(n4203) );
  XNOR U5357 ( .A(n4198), .B(n4202), .Z(n4204) );
  XOR U5358 ( .A(n4205), .B(n4206), .Z(n4202) );
  ANDN U5359 ( .B(n4126), .A(n4127), .Z(n4205) );
  AND U5360 ( .A(b[2]), .B(a[80]), .Z(n4207) );
  XNOR U5361 ( .A(n4209), .B(n4206), .Z(n4208) );
  XOR U5362 ( .A(n4210), .B(n4211), .Z(n4206) );
  NANDN U5363 ( .A(n4129), .B(n4128), .Z(n4211) );
  XOR U5364 ( .A(n4210), .B(n4212), .Z(n4128) );
  NAND U5365 ( .A(a[80]), .B(b[1]), .Z(n4212) );
  XOR U5366 ( .A(n4210), .B(n4214), .Z(n4213) );
  OR U5367 ( .A(n2497), .B(n2495), .Z(n4210) );
  XOR U5368 ( .A(n4216), .B(n4217), .Z(n2495) );
  NANDN U5369 ( .A(n179), .B(a[80]), .Z(n2497) );
  XNOR U5370 ( .A(n4193), .B(n4197), .Z(n4219) );
  XNOR U5371 ( .A(n4188), .B(n4192), .Z(n4220) );
  XNOR U5372 ( .A(n4183), .B(n4187), .Z(n4221) );
  XNOR U5373 ( .A(n4178), .B(n4182), .Z(n4222) );
  XNOR U5374 ( .A(n4173), .B(n4177), .Z(n4223) );
  XNOR U5375 ( .A(n4168), .B(n4172), .Z(n4224) );
  XNOR U5376 ( .A(n4163), .B(n4167), .Z(n4225) );
  XOR U5377 ( .A(n4159), .B(n4162), .Z(n4226) );
  XOR U5378 ( .A(n4227), .B(n4228), .Z(n4159) );
  XNOR U5379 ( .A(n4229), .B(n4230), .Z(n4228) );
  XNOR U5380 ( .A(n4231), .B(n4232), .Z(n4229) );
  XOR U5381 ( .A(n4233), .B(n4234), .Z(n4232) );
  AND U5382 ( .A(b[14]), .B(a[69]), .Z(n4234) );
  AND U5383 ( .A(a[68]), .B(b[15]), .Z(n4233) );
  XNOR U5384 ( .A(n4235), .B(n4231), .Z(n4227) );
  XOR U5385 ( .A(n4236), .B(n4237), .Z(n4231) );
  NOR U5386 ( .A(n4238), .B(n4239), .Z(n4236) );
  AND U5387 ( .A(a[70]), .B(b[13]), .Z(n4235) );
  XOR U5388 ( .A(n4240), .B(n4157), .Z(n4158) );
  IV U5389 ( .A(n4230), .Z(n4157) );
  XOR U5390 ( .A(n4241), .B(n4242), .Z(n4230) );
  ANDN U5391 ( .B(n4243), .A(n4244), .Z(n4241) );
  AND U5392 ( .A(a[71]), .B(b[12]), .Z(n4240) );
  XOR U5393 ( .A(n4246), .B(n4247), .Z(n4162) );
  ANDN U5394 ( .B(n4248), .A(n4249), .Z(n4246) );
  AND U5395 ( .A(a[72]), .B(b[11]), .Z(n4245) );
  XOR U5396 ( .A(n4251), .B(n4252), .Z(n4167) );
  ANDN U5397 ( .B(n4253), .A(n4254), .Z(n4251) );
  AND U5398 ( .A(a[73]), .B(b[10]), .Z(n4250) );
  XOR U5399 ( .A(n4256), .B(n4257), .Z(n4172) );
  ANDN U5400 ( .B(n4258), .A(n4259), .Z(n4256) );
  AND U5401 ( .A(a[74]), .B(b[9]), .Z(n4255) );
  XOR U5402 ( .A(n4261), .B(n4262), .Z(n4177) );
  ANDN U5403 ( .B(n4263), .A(n4264), .Z(n4261) );
  AND U5404 ( .A(a[75]), .B(b[8]), .Z(n4260) );
  XOR U5405 ( .A(n4266), .B(n4267), .Z(n4182) );
  ANDN U5406 ( .B(n4268), .A(n4269), .Z(n4266) );
  AND U5407 ( .A(a[76]), .B(b[7]), .Z(n4265) );
  XOR U5408 ( .A(n4271), .B(n4272), .Z(n4187) );
  ANDN U5409 ( .B(n4273), .A(n4274), .Z(n4271) );
  AND U5410 ( .A(a[77]), .B(b[6]), .Z(n4270) );
  XOR U5411 ( .A(n4276), .B(n4277), .Z(n4192) );
  ANDN U5412 ( .B(n4278), .A(n4279), .Z(n4276) );
  AND U5413 ( .A(a[78]), .B(b[5]), .Z(n4275) );
  XOR U5414 ( .A(n4281), .B(n4282), .Z(n4197) );
  ANDN U5415 ( .B(n4209), .A(n4218), .Z(n4281) );
  AND U5416 ( .A(a[79]), .B(b[3]), .Z(n4283) );
  XNOR U5417 ( .A(n4278), .B(n4282), .Z(n4284) );
  XOR U5418 ( .A(n4285), .B(n4286), .Z(n4282) );
  ANDN U5419 ( .B(n4214), .A(n4215), .Z(n4285) );
  AND U5420 ( .A(b[2]), .B(a[79]), .Z(n4287) );
  XNOR U5421 ( .A(n4289), .B(n4286), .Z(n4288) );
  XOR U5422 ( .A(n4290), .B(n4291), .Z(n4286) );
  NANDN U5423 ( .A(n4217), .B(n4216), .Z(n4291) );
  XOR U5424 ( .A(n4290), .B(n4292), .Z(n4216) );
  NAND U5425 ( .A(a[79]), .B(b[1]), .Z(n4292) );
  XOR U5426 ( .A(n4290), .B(n4294), .Z(n4293) );
  OR U5427 ( .A(n2502), .B(n2500), .Z(n4290) );
  XOR U5428 ( .A(n4296), .B(n4297), .Z(n2500) );
  NANDN U5429 ( .A(n179), .B(a[79]), .Z(n2502) );
  XNOR U5430 ( .A(n4273), .B(n4277), .Z(n4299) );
  XNOR U5431 ( .A(n4268), .B(n4272), .Z(n4300) );
  XNOR U5432 ( .A(n4263), .B(n4267), .Z(n4301) );
  XNOR U5433 ( .A(n4258), .B(n4262), .Z(n4302) );
  XNOR U5434 ( .A(n4253), .B(n4257), .Z(n4303) );
  XNOR U5435 ( .A(n4248), .B(n4252), .Z(n4304) );
  XNOR U5436 ( .A(n4243), .B(n4247), .Z(n4305) );
  XOR U5437 ( .A(n4239), .B(n4242), .Z(n4306) );
  XOR U5438 ( .A(n4307), .B(n4308), .Z(n4239) );
  XNOR U5439 ( .A(n4309), .B(n4310), .Z(n4308) );
  XOR U5440 ( .A(n4311), .B(n4312), .Z(n4309) );
  AND U5441 ( .A(b[13]), .B(a[69]), .Z(n4311) );
  XOR U5442 ( .A(n4312), .B(n4313), .Z(n4307) );
  XOR U5443 ( .A(n4314), .B(n4315), .Z(n4313) );
  AND U5444 ( .A(a[68]), .B(b[14]), .Z(n4315) );
  AND U5445 ( .A(a[67]), .B(b[15]), .Z(n4314) );
  XOR U5446 ( .A(n4316), .B(n4317), .Z(n4312) );
  ANDN U5447 ( .B(n4318), .A(n4319), .Z(n4316) );
  XOR U5448 ( .A(n4320), .B(n4237), .Z(n4238) );
  IV U5449 ( .A(n4310), .Z(n4237) );
  XOR U5450 ( .A(n4321), .B(n4322), .Z(n4310) );
  NOR U5451 ( .A(n4323), .B(n4324), .Z(n4321) );
  AND U5452 ( .A(a[70]), .B(b[12]), .Z(n4320) );
  XOR U5453 ( .A(n4326), .B(n4327), .Z(n4242) );
  ANDN U5454 ( .B(n4328), .A(n4329), .Z(n4326) );
  AND U5455 ( .A(a[71]), .B(b[11]), .Z(n4325) );
  XOR U5456 ( .A(n4331), .B(n4332), .Z(n4247) );
  ANDN U5457 ( .B(n4333), .A(n4334), .Z(n4331) );
  AND U5458 ( .A(a[72]), .B(b[10]), .Z(n4330) );
  XOR U5459 ( .A(n4336), .B(n4337), .Z(n4252) );
  ANDN U5460 ( .B(n4338), .A(n4339), .Z(n4336) );
  AND U5461 ( .A(a[73]), .B(b[9]), .Z(n4335) );
  XOR U5462 ( .A(n4341), .B(n4342), .Z(n4257) );
  ANDN U5463 ( .B(n4343), .A(n4344), .Z(n4341) );
  AND U5464 ( .A(a[74]), .B(b[8]), .Z(n4340) );
  XOR U5465 ( .A(n4346), .B(n4347), .Z(n4262) );
  ANDN U5466 ( .B(n4348), .A(n4349), .Z(n4346) );
  AND U5467 ( .A(a[75]), .B(b[7]), .Z(n4345) );
  XOR U5468 ( .A(n4351), .B(n4352), .Z(n4267) );
  ANDN U5469 ( .B(n4353), .A(n4354), .Z(n4351) );
  AND U5470 ( .A(a[76]), .B(b[6]), .Z(n4350) );
  XOR U5471 ( .A(n4356), .B(n4357), .Z(n4272) );
  ANDN U5472 ( .B(n4358), .A(n4359), .Z(n4356) );
  AND U5473 ( .A(a[77]), .B(b[5]), .Z(n4355) );
  XOR U5474 ( .A(n4361), .B(n4362), .Z(n4277) );
  ANDN U5475 ( .B(n4289), .A(n4298), .Z(n4361) );
  AND U5476 ( .A(a[78]), .B(b[3]), .Z(n4363) );
  XNOR U5477 ( .A(n4358), .B(n4362), .Z(n4364) );
  XOR U5478 ( .A(n4365), .B(n4366), .Z(n4362) );
  ANDN U5479 ( .B(n4294), .A(n4295), .Z(n4365) );
  AND U5480 ( .A(b[2]), .B(a[78]), .Z(n4367) );
  XNOR U5481 ( .A(n4369), .B(n4366), .Z(n4368) );
  XOR U5482 ( .A(n4370), .B(n4371), .Z(n4366) );
  NANDN U5483 ( .A(n4297), .B(n4296), .Z(n4371) );
  XOR U5484 ( .A(n4370), .B(n4372), .Z(n4296) );
  NAND U5485 ( .A(a[78]), .B(b[1]), .Z(n4372) );
  XOR U5486 ( .A(n4370), .B(n4374), .Z(n4373) );
  OR U5487 ( .A(n2507), .B(n2505), .Z(n4370) );
  XOR U5488 ( .A(n4376), .B(n4377), .Z(n2505) );
  NANDN U5489 ( .A(n179), .B(a[78]), .Z(n2507) );
  XNOR U5490 ( .A(n4353), .B(n4357), .Z(n4379) );
  XNOR U5491 ( .A(n4348), .B(n4352), .Z(n4380) );
  XNOR U5492 ( .A(n4343), .B(n4347), .Z(n4381) );
  XNOR U5493 ( .A(n4338), .B(n4342), .Z(n4382) );
  XNOR U5494 ( .A(n4333), .B(n4337), .Z(n4383) );
  XNOR U5495 ( .A(n4328), .B(n4332), .Z(n4384) );
  XOR U5496 ( .A(n4324), .B(n4327), .Z(n4385) );
  XNOR U5497 ( .A(n4319), .B(n4386), .Z(n4324) );
  XNOR U5498 ( .A(n4318), .B(n4322), .Z(n4386) );
  XOR U5499 ( .A(n4387), .B(n4317), .Z(n4318) );
  AND U5500 ( .A(b[12]), .B(a[69]), .Z(n4387) );
  XOR U5501 ( .A(n4388), .B(n4389), .Z(n4319) );
  XOR U5502 ( .A(n4317), .B(n4390), .Z(n4389) );
  XOR U5503 ( .A(n4391), .B(n4392), .Z(n4390) );
  XOR U5504 ( .A(n4393), .B(n4394), .Z(n4392) );
  NAND U5505 ( .A(a[67]), .B(b[14]), .Z(n4394) );
  AND U5506 ( .A(a[66]), .B(b[15]), .Z(n4393) );
  XOR U5507 ( .A(n4395), .B(n4396), .Z(n4317) );
  ANDN U5508 ( .B(n4397), .A(n4398), .Z(n4395) );
  XOR U5509 ( .A(n4399), .B(n4391), .Z(n4388) );
  XOR U5510 ( .A(n4400), .B(n4401), .Z(n4391) );
  NOR U5511 ( .A(n4402), .B(n4403), .Z(n4400) );
  AND U5512 ( .A(a[68]), .B(b[13]), .Z(n4399) );
  XOR U5513 ( .A(n4405), .B(n4406), .Z(n4322) );
  ANDN U5514 ( .B(n4407), .A(n4408), .Z(n4405) );
  AND U5515 ( .A(a[70]), .B(b[11]), .Z(n4404) );
  XOR U5516 ( .A(n4410), .B(n4411), .Z(n4327) );
  ANDN U5517 ( .B(n4412), .A(n4413), .Z(n4410) );
  AND U5518 ( .A(a[71]), .B(b[10]), .Z(n4409) );
  XOR U5519 ( .A(n4415), .B(n4416), .Z(n4332) );
  ANDN U5520 ( .B(n4417), .A(n4418), .Z(n4415) );
  AND U5521 ( .A(a[72]), .B(b[9]), .Z(n4414) );
  XOR U5522 ( .A(n4420), .B(n4421), .Z(n4337) );
  ANDN U5523 ( .B(n4422), .A(n4423), .Z(n4420) );
  AND U5524 ( .A(a[73]), .B(b[8]), .Z(n4419) );
  XOR U5525 ( .A(n4425), .B(n4426), .Z(n4342) );
  ANDN U5526 ( .B(n4427), .A(n4428), .Z(n4425) );
  AND U5527 ( .A(a[74]), .B(b[7]), .Z(n4424) );
  XOR U5528 ( .A(n4430), .B(n4431), .Z(n4347) );
  ANDN U5529 ( .B(n4432), .A(n4433), .Z(n4430) );
  AND U5530 ( .A(a[75]), .B(b[6]), .Z(n4429) );
  XOR U5531 ( .A(n4435), .B(n4436), .Z(n4352) );
  ANDN U5532 ( .B(n4437), .A(n4438), .Z(n4435) );
  AND U5533 ( .A(a[76]), .B(b[5]), .Z(n4434) );
  XOR U5534 ( .A(n4440), .B(n4441), .Z(n4357) );
  ANDN U5535 ( .B(n4369), .A(n4378), .Z(n4440) );
  AND U5536 ( .A(a[77]), .B(b[3]), .Z(n4442) );
  XNOR U5537 ( .A(n4437), .B(n4441), .Z(n4443) );
  XOR U5538 ( .A(n4444), .B(n4445), .Z(n4441) );
  ANDN U5539 ( .B(n4374), .A(n4375), .Z(n4444) );
  AND U5540 ( .A(b[2]), .B(a[77]), .Z(n4446) );
  XNOR U5541 ( .A(n4448), .B(n4445), .Z(n4447) );
  XOR U5542 ( .A(n4449), .B(n4450), .Z(n4445) );
  NANDN U5543 ( .A(n4377), .B(n4376), .Z(n4450) );
  XOR U5544 ( .A(n4449), .B(n4451), .Z(n4376) );
  NAND U5545 ( .A(a[77]), .B(b[1]), .Z(n4451) );
  XOR U5546 ( .A(n4449), .B(n4453), .Z(n4452) );
  OR U5547 ( .A(n2512), .B(n2510), .Z(n4449) );
  XOR U5548 ( .A(n4455), .B(n4456), .Z(n2510) );
  NANDN U5549 ( .A(n179), .B(a[77]), .Z(n2512) );
  XNOR U5550 ( .A(n4432), .B(n4436), .Z(n4458) );
  XNOR U5551 ( .A(n4427), .B(n4431), .Z(n4459) );
  XNOR U5552 ( .A(n4422), .B(n4426), .Z(n4460) );
  XNOR U5553 ( .A(n4417), .B(n4421), .Z(n4461) );
  XNOR U5554 ( .A(n4412), .B(n4416), .Z(n4462) );
  XNOR U5555 ( .A(n4407), .B(n4411), .Z(n4463) );
  XNOR U5556 ( .A(n4397), .B(n4406), .Z(n4464) );
  XOR U5557 ( .A(n4465), .B(n4396), .Z(n4397) );
  AND U5558 ( .A(b[11]), .B(a[69]), .Z(n4465) );
  XOR U5559 ( .A(n4396), .B(n4403), .Z(n4466) );
  XOR U5560 ( .A(n4467), .B(n4468), .Z(n4403) );
  XOR U5561 ( .A(n4401), .B(n4469), .Z(n4468) );
  XOR U5562 ( .A(n4470), .B(n4471), .Z(n4469) );
  XOR U5563 ( .A(n4472), .B(n4473), .Z(n4471) );
  NAND U5564 ( .A(a[66]), .B(b[14]), .Z(n4473) );
  AND U5565 ( .A(a[65]), .B(b[15]), .Z(n4472) );
  XOR U5566 ( .A(n4474), .B(n4470), .Z(n4467) );
  XOR U5567 ( .A(n4475), .B(n4476), .Z(n4470) );
  NOR U5568 ( .A(n4477), .B(n4478), .Z(n4475) );
  AND U5569 ( .A(a[67]), .B(b[13]), .Z(n4474) );
  XOR U5570 ( .A(n4479), .B(n4480), .Z(n4396) );
  ANDN U5571 ( .B(n4481), .A(n4482), .Z(n4479) );
  XNOR U5572 ( .A(n4483), .B(n4401), .Z(n4402) );
  XOR U5573 ( .A(n4484), .B(n4485), .Z(n4401) );
  ANDN U5574 ( .B(n4486), .A(n4487), .Z(n4484) );
  AND U5575 ( .A(a[68]), .B(b[12]), .Z(n4483) );
  XOR U5576 ( .A(n4489), .B(n4490), .Z(n4406) );
  ANDN U5577 ( .B(n4491), .A(n4492), .Z(n4489) );
  AND U5578 ( .A(a[70]), .B(b[10]), .Z(n4488) );
  XOR U5579 ( .A(n4494), .B(n4495), .Z(n4411) );
  ANDN U5580 ( .B(n4496), .A(n4497), .Z(n4494) );
  AND U5581 ( .A(a[71]), .B(b[9]), .Z(n4493) );
  XOR U5582 ( .A(n4499), .B(n4500), .Z(n4416) );
  ANDN U5583 ( .B(n4501), .A(n4502), .Z(n4499) );
  AND U5584 ( .A(a[72]), .B(b[8]), .Z(n4498) );
  XOR U5585 ( .A(n4504), .B(n4505), .Z(n4421) );
  ANDN U5586 ( .B(n4506), .A(n4507), .Z(n4504) );
  AND U5587 ( .A(a[73]), .B(b[7]), .Z(n4503) );
  XOR U5588 ( .A(n4509), .B(n4510), .Z(n4426) );
  ANDN U5589 ( .B(n4511), .A(n4512), .Z(n4509) );
  AND U5590 ( .A(a[74]), .B(b[6]), .Z(n4508) );
  XOR U5591 ( .A(n4514), .B(n4515), .Z(n4431) );
  ANDN U5592 ( .B(n4516), .A(n4517), .Z(n4514) );
  AND U5593 ( .A(a[75]), .B(b[5]), .Z(n4513) );
  XOR U5594 ( .A(n4519), .B(n4520), .Z(n4436) );
  ANDN U5595 ( .B(n4448), .A(n4457), .Z(n4519) );
  AND U5596 ( .A(a[76]), .B(b[3]), .Z(n4521) );
  XNOR U5597 ( .A(n4516), .B(n4520), .Z(n4522) );
  XOR U5598 ( .A(n4523), .B(n4524), .Z(n4520) );
  ANDN U5599 ( .B(n4453), .A(n4454), .Z(n4523) );
  AND U5600 ( .A(b[2]), .B(a[76]), .Z(n4525) );
  XNOR U5601 ( .A(n4527), .B(n4524), .Z(n4526) );
  XOR U5602 ( .A(n4528), .B(n4529), .Z(n4524) );
  NANDN U5603 ( .A(n4456), .B(n4455), .Z(n4529) );
  XOR U5604 ( .A(n4528), .B(n4530), .Z(n4455) );
  NAND U5605 ( .A(a[76]), .B(b[1]), .Z(n4530) );
  XOR U5606 ( .A(n4528), .B(n4532), .Z(n4531) );
  OR U5607 ( .A(n2517), .B(n2515), .Z(n4528) );
  XOR U5608 ( .A(n4534), .B(n4535), .Z(n2515) );
  NANDN U5609 ( .A(n179), .B(a[76]), .Z(n2517) );
  XNOR U5610 ( .A(n4511), .B(n4515), .Z(n4537) );
  XNOR U5611 ( .A(n4506), .B(n4510), .Z(n4538) );
  XNOR U5612 ( .A(n4501), .B(n4505), .Z(n4539) );
  XNOR U5613 ( .A(n4496), .B(n4500), .Z(n4540) );
  XNOR U5614 ( .A(n4491), .B(n4495), .Z(n4541) );
  XNOR U5615 ( .A(n4481), .B(n4490), .Z(n4542) );
  XOR U5616 ( .A(n4543), .B(n4480), .Z(n4481) );
  AND U5617 ( .A(b[10]), .B(a[69]), .Z(n4543) );
  XNOR U5618 ( .A(n4480), .B(n4486), .Z(n4544) );
  XOR U5619 ( .A(n4485), .B(n4478), .Z(n4545) );
  XOR U5620 ( .A(n4546), .B(n4547), .Z(n4478) );
  XOR U5621 ( .A(n4476), .B(n4548), .Z(n4547) );
  XOR U5622 ( .A(n4549), .B(n4550), .Z(n4548) );
  XOR U5623 ( .A(n4551), .B(n4552), .Z(n4550) );
  NAND U5624 ( .A(a[65]), .B(b[14]), .Z(n4552) );
  AND U5625 ( .A(a[64]), .B(b[15]), .Z(n4551) );
  XOR U5626 ( .A(n4553), .B(n4549), .Z(n4546) );
  XOR U5627 ( .A(n4554), .B(n4555), .Z(n4549) );
  NOR U5628 ( .A(n4556), .B(n4557), .Z(n4554) );
  AND U5629 ( .A(a[66]), .B(b[13]), .Z(n4553) );
  XNOR U5630 ( .A(n4558), .B(n4476), .Z(n4477) );
  XOR U5631 ( .A(n4559), .B(n4560), .Z(n4476) );
  ANDN U5632 ( .B(n4561), .A(n4562), .Z(n4559) );
  AND U5633 ( .A(a[67]), .B(b[12]), .Z(n4558) );
  XOR U5634 ( .A(n4563), .B(n4564), .Z(n4480) );
  ANDN U5635 ( .B(n4565), .A(n4566), .Z(n4563) );
  XNOR U5636 ( .A(n4567), .B(n4485), .Z(n4487) );
  XOR U5637 ( .A(n4568), .B(n4569), .Z(n4485) );
  ANDN U5638 ( .B(n4570), .A(n4571), .Z(n4568) );
  AND U5639 ( .A(a[68]), .B(b[11]), .Z(n4567) );
  XOR U5640 ( .A(n4573), .B(n4574), .Z(n4490) );
  ANDN U5641 ( .B(n4575), .A(n4576), .Z(n4573) );
  AND U5642 ( .A(a[70]), .B(b[9]), .Z(n4572) );
  XOR U5643 ( .A(n4578), .B(n4579), .Z(n4495) );
  ANDN U5644 ( .B(n4580), .A(n4581), .Z(n4578) );
  AND U5645 ( .A(a[71]), .B(b[8]), .Z(n4577) );
  XOR U5646 ( .A(n4583), .B(n4584), .Z(n4500) );
  ANDN U5647 ( .B(n4585), .A(n4586), .Z(n4583) );
  AND U5648 ( .A(a[72]), .B(b[7]), .Z(n4582) );
  XOR U5649 ( .A(n4588), .B(n4589), .Z(n4505) );
  ANDN U5650 ( .B(n4590), .A(n4591), .Z(n4588) );
  AND U5651 ( .A(a[73]), .B(b[6]), .Z(n4587) );
  XOR U5652 ( .A(n4593), .B(n4594), .Z(n4510) );
  ANDN U5653 ( .B(n4595), .A(n4596), .Z(n4593) );
  AND U5654 ( .A(a[74]), .B(b[5]), .Z(n4592) );
  XOR U5655 ( .A(n4598), .B(n4599), .Z(n4515) );
  ANDN U5656 ( .B(n4527), .A(n4536), .Z(n4598) );
  AND U5657 ( .A(a[75]), .B(b[3]), .Z(n4600) );
  XNOR U5658 ( .A(n4595), .B(n4599), .Z(n4601) );
  XOR U5659 ( .A(n4602), .B(n4603), .Z(n4599) );
  ANDN U5660 ( .B(n4532), .A(n4533), .Z(n4602) );
  AND U5661 ( .A(b[2]), .B(a[75]), .Z(n4604) );
  XNOR U5662 ( .A(n4606), .B(n4603), .Z(n4605) );
  XOR U5663 ( .A(n4607), .B(n4608), .Z(n4603) );
  NANDN U5664 ( .A(n4535), .B(n4534), .Z(n4608) );
  XOR U5665 ( .A(n4607), .B(n4609), .Z(n4534) );
  NAND U5666 ( .A(a[75]), .B(b[1]), .Z(n4609) );
  XOR U5667 ( .A(n4607), .B(n4611), .Z(n4610) );
  OR U5668 ( .A(n2522), .B(n2520), .Z(n4607) );
  XOR U5669 ( .A(n4613), .B(n4614), .Z(n2520) );
  NANDN U5670 ( .A(n179), .B(a[75]), .Z(n2522) );
  XNOR U5671 ( .A(n4590), .B(n4594), .Z(n4616) );
  XNOR U5672 ( .A(n4585), .B(n4589), .Z(n4617) );
  XNOR U5673 ( .A(n4580), .B(n4584), .Z(n4618) );
  XNOR U5674 ( .A(n4575), .B(n4579), .Z(n4619) );
  XNOR U5675 ( .A(n4565), .B(n4574), .Z(n4620) );
  XOR U5676 ( .A(n4621), .B(n4564), .Z(n4565) );
  AND U5677 ( .A(b[9]), .B(a[69]), .Z(n4621) );
  XNOR U5678 ( .A(n4564), .B(n4570), .Z(n4622) );
  XNOR U5679 ( .A(n4569), .B(n4561), .Z(n4623) );
  XOR U5680 ( .A(n4560), .B(n4557), .Z(n4624) );
  XOR U5681 ( .A(n4625), .B(n4626), .Z(n4557) );
  XOR U5682 ( .A(n4555), .B(n4627), .Z(n4626) );
  XOR U5683 ( .A(n4628), .B(n4629), .Z(n4627) );
  XOR U5684 ( .A(n4630), .B(n4631), .Z(n4629) );
  NAND U5685 ( .A(a[64]), .B(b[14]), .Z(n4631) );
  AND U5686 ( .A(a[63]), .B(b[15]), .Z(n4630) );
  XOR U5687 ( .A(n4632), .B(n4628), .Z(n4625) );
  XOR U5688 ( .A(n4633), .B(n4634), .Z(n4628) );
  NOR U5689 ( .A(n4635), .B(n4636), .Z(n4633) );
  AND U5690 ( .A(a[65]), .B(b[13]), .Z(n4632) );
  XNOR U5691 ( .A(n4637), .B(n4555), .Z(n4556) );
  XOR U5692 ( .A(n4638), .B(n4639), .Z(n4555) );
  ANDN U5693 ( .B(n4640), .A(n4641), .Z(n4638) );
  AND U5694 ( .A(a[66]), .B(b[12]), .Z(n4637) );
  XNOR U5695 ( .A(n4642), .B(n4560), .Z(n4562) );
  XOR U5696 ( .A(n4643), .B(n4644), .Z(n4560) );
  ANDN U5697 ( .B(n4645), .A(n4646), .Z(n4643) );
  AND U5698 ( .A(a[67]), .B(b[11]), .Z(n4642) );
  XOR U5699 ( .A(n4647), .B(n4648), .Z(n4564) );
  ANDN U5700 ( .B(n4649), .A(n4650), .Z(n4647) );
  XNOR U5701 ( .A(n4651), .B(n4569), .Z(n4571) );
  XOR U5702 ( .A(n4652), .B(n4653), .Z(n4569) );
  ANDN U5703 ( .B(n4654), .A(n4655), .Z(n4652) );
  AND U5704 ( .A(a[68]), .B(b[10]), .Z(n4651) );
  XOR U5705 ( .A(n4657), .B(n4658), .Z(n4574) );
  ANDN U5706 ( .B(n4659), .A(n4660), .Z(n4657) );
  AND U5707 ( .A(a[70]), .B(b[8]), .Z(n4656) );
  XOR U5708 ( .A(n4662), .B(n4663), .Z(n4579) );
  ANDN U5709 ( .B(n4664), .A(n4665), .Z(n4662) );
  AND U5710 ( .A(a[71]), .B(b[7]), .Z(n4661) );
  XOR U5711 ( .A(n4667), .B(n4668), .Z(n4584) );
  ANDN U5712 ( .B(n4669), .A(n4670), .Z(n4667) );
  AND U5713 ( .A(a[72]), .B(b[6]), .Z(n4666) );
  XOR U5714 ( .A(n4672), .B(n4673), .Z(n4589) );
  ANDN U5715 ( .B(n4674), .A(n4675), .Z(n4672) );
  AND U5716 ( .A(a[73]), .B(b[5]), .Z(n4671) );
  XOR U5717 ( .A(n4677), .B(n4678), .Z(n4594) );
  ANDN U5718 ( .B(n4606), .A(n4615), .Z(n4677) );
  AND U5719 ( .A(a[74]), .B(b[3]), .Z(n4679) );
  XNOR U5720 ( .A(n4674), .B(n4678), .Z(n4680) );
  XOR U5721 ( .A(n4681), .B(n4682), .Z(n4678) );
  ANDN U5722 ( .B(n4611), .A(n4612), .Z(n4681) );
  AND U5723 ( .A(b[2]), .B(a[74]), .Z(n4683) );
  XNOR U5724 ( .A(n4685), .B(n4682), .Z(n4684) );
  XOR U5725 ( .A(n4686), .B(n4687), .Z(n4682) );
  NANDN U5726 ( .A(n4614), .B(n4613), .Z(n4687) );
  XOR U5727 ( .A(n4686), .B(n4688), .Z(n4613) );
  NAND U5728 ( .A(a[74]), .B(b[1]), .Z(n4688) );
  XOR U5729 ( .A(n4686), .B(n4690), .Z(n4689) );
  OR U5730 ( .A(n2527), .B(n2525), .Z(n4686) );
  XOR U5731 ( .A(n4692), .B(n4693), .Z(n2525) );
  NANDN U5732 ( .A(n179), .B(a[74]), .Z(n2527) );
  XNOR U5733 ( .A(n4669), .B(n4673), .Z(n4695) );
  XNOR U5734 ( .A(n4664), .B(n4668), .Z(n4696) );
  XNOR U5735 ( .A(n4659), .B(n4663), .Z(n4697) );
  XNOR U5736 ( .A(n4649), .B(n4658), .Z(n4698) );
  XOR U5737 ( .A(n4699), .B(n4648), .Z(n4649) );
  AND U5738 ( .A(b[8]), .B(a[69]), .Z(n4699) );
  XNOR U5739 ( .A(n4648), .B(n4654), .Z(n4700) );
  XNOR U5740 ( .A(n4653), .B(n4645), .Z(n4701) );
  XNOR U5741 ( .A(n4644), .B(n4640), .Z(n4702) );
  XOR U5742 ( .A(n4639), .B(n4636), .Z(n4703) );
  XOR U5743 ( .A(n4704), .B(n4705), .Z(n4636) );
  XOR U5744 ( .A(n4634), .B(n4706), .Z(n4705) );
  XOR U5745 ( .A(n4707), .B(n4708), .Z(n4706) );
  XOR U5746 ( .A(n4709), .B(n4710), .Z(n4708) );
  NAND U5747 ( .A(a[63]), .B(b[14]), .Z(n4710) );
  AND U5748 ( .A(a[62]), .B(b[15]), .Z(n4709) );
  XOR U5749 ( .A(n4711), .B(n4707), .Z(n4704) );
  XOR U5750 ( .A(n4712), .B(n4713), .Z(n4707) );
  NOR U5751 ( .A(n4714), .B(n4715), .Z(n4712) );
  AND U5752 ( .A(a[64]), .B(b[13]), .Z(n4711) );
  XNOR U5753 ( .A(n4716), .B(n4634), .Z(n4635) );
  XOR U5754 ( .A(n4717), .B(n4718), .Z(n4634) );
  ANDN U5755 ( .B(n4719), .A(n4720), .Z(n4717) );
  AND U5756 ( .A(a[65]), .B(b[12]), .Z(n4716) );
  XNOR U5757 ( .A(n4721), .B(n4639), .Z(n4641) );
  XOR U5758 ( .A(n4722), .B(n4723), .Z(n4639) );
  ANDN U5759 ( .B(n4724), .A(n4725), .Z(n4722) );
  AND U5760 ( .A(a[66]), .B(b[11]), .Z(n4721) );
  XNOR U5761 ( .A(n4726), .B(n4644), .Z(n4646) );
  XOR U5762 ( .A(n4727), .B(n4728), .Z(n4644) );
  ANDN U5763 ( .B(n4729), .A(n4730), .Z(n4727) );
  AND U5764 ( .A(a[67]), .B(b[10]), .Z(n4726) );
  XOR U5765 ( .A(n4731), .B(n4732), .Z(n4648) );
  ANDN U5766 ( .B(n4733), .A(n4734), .Z(n4731) );
  XNOR U5767 ( .A(n4735), .B(n4653), .Z(n4655) );
  XOR U5768 ( .A(n4736), .B(n4737), .Z(n4653) );
  ANDN U5769 ( .B(n4738), .A(n4739), .Z(n4736) );
  AND U5770 ( .A(a[68]), .B(b[9]), .Z(n4735) );
  XOR U5771 ( .A(n4741), .B(n4742), .Z(n4658) );
  ANDN U5772 ( .B(n4743), .A(n4744), .Z(n4741) );
  AND U5773 ( .A(a[70]), .B(b[7]), .Z(n4740) );
  XOR U5774 ( .A(n4746), .B(n4747), .Z(n4663) );
  ANDN U5775 ( .B(n4748), .A(n4749), .Z(n4746) );
  AND U5776 ( .A(a[71]), .B(b[6]), .Z(n4745) );
  XOR U5777 ( .A(n4751), .B(n4752), .Z(n4668) );
  ANDN U5778 ( .B(n4753), .A(n4754), .Z(n4751) );
  AND U5779 ( .A(a[72]), .B(b[5]), .Z(n4750) );
  XOR U5780 ( .A(n4756), .B(n4757), .Z(n4673) );
  ANDN U5781 ( .B(n4685), .A(n4694), .Z(n4756) );
  AND U5782 ( .A(a[73]), .B(b[3]), .Z(n4758) );
  XNOR U5783 ( .A(n4753), .B(n4757), .Z(n4759) );
  XOR U5784 ( .A(n4760), .B(n4761), .Z(n4757) );
  ANDN U5785 ( .B(n4690), .A(n4691), .Z(n4760) );
  AND U5786 ( .A(b[2]), .B(a[73]), .Z(n4762) );
  XNOR U5787 ( .A(n4764), .B(n4761), .Z(n4763) );
  XOR U5788 ( .A(n4765), .B(n4766), .Z(n4761) );
  NANDN U5789 ( .A(n4693), .B(n4692), .Z(n4766) );
  XOR U5790 ( .A(n4765), .B(n4767), .Z(n4692) );
  NAND U5791 ( .A(a[73]), .B(b[1]), .Z(n4767) );
  XOR U5792 ( .A(n4765), .B(n4769), .Z(n4768) );
  OR U5793 ( .A(n2532), .B(n2530), .Z(n4765) );
  XOR U5794 ( .A(n4771), .B(n4772), .Z(n2530) );
  NANDN U5795 ( .A(n179), .B(a[73]), .Z(n2532) );
  XNOR U5796 ( .A(n4748), .B(n4752), .Z(n4774) );
  XNOR U5797 ( .A(n4743), .B(n4747), .Z(n4775) );
  XNOR U5798 ( .A(n4733), .B(n4742), .Z(n4776) );
  XOR U5799 ( .A(n4777), .B(n4732), .Z(n4733) );
  AND U5800 ( .A(b[7]), .B(a[69]), .Z(n4777) );
  XNOR U5801 ( .A(n4732), .B(n4738), .Z(n4778) );
  XNOR U5802 ( .A(n4737), .B(n4729), .Z(n4779) );
  XNOR U5803 ( .A(n4728), .B(n4724), .Z(n4780) );
  XNOR U5804 ( .A(n4723), .B(n4719), .Z(n4781) );
  XOR U5805 ( .A(n4718), .B(n4715), .Z(n4782) );
  XOR U5806 ( .A(n4783), .B(n4784), .Z(n4715) );
  XOR U5807 ( .A(n4713), .B(n4785), .Z(n4784) );
  XOR U5808 ( .A(n4786), .B(n4787), .Z(n4785) );
  XOR U5809 ( .A(n4788), .B(n4789), .Z(n4787) );
  NAND U5810 ( .A(a[62]), .B(b[14]), .Z(n4789) );
  AND U5811 ( .A(a[61]), .B(b[15]), .Z(n4788) );
  XOR U5812 ( .A(n4790), .B(n4786), .Z(n4783) );
  XOR U5813 ( .A(n4791), .B(n4792), .Z(n4786) );
  NOR U5814 ( .A(n4793), .B(n4794), .Z(n4791) );
  AND U5815 ( .A(a[63]), .B(b[13]), .Z(n4790) );
  XNOR U5816 ( .A(n4795), .B(n4713), .Z(n4714) );
  XOR U5817 ( .A(n4796), .B(n4797), .Z(n4713) );
  ANDN U5818 ( .B(n4798), .A(n4799), .Z(n4796) );
  AND U5819 ( .A(a[64]), .B(b[12]), .Z(n4795) );
  XNOR U5820 ( .A(n4800), .B(n4718), .Z(n4720) );
  XOR U5821 ( .A(n4801), .B(n4802), .Z(n4718) );
  ANDN U5822 ( .B(n4803), .A(n4804), .Z(n4801) );
  AND U5823 ( .A(a[65]), .B(b[11]), .Z(n4800) );
  XNOR U5824 ( .A(n4805), .B(n4723), .Z(n4725) );
  XOR U5825 ( .A(n4806), .B(n4807), .Z(n4723) );
  ANDN U5826 ( .B(n4808), .A(n4809), .Z(n4806) );
  AND U5827 ( .A(a[66]), .B(b[10]), .Z(n4805) );
  XNOR U5828 ( .A(n4810), .B(n4728), .Z(n4730) );
  XOR U5829 ( .A(n4811), .B(n4812), .Z(n4728) );
  ANDN U5830 ( .B(n4813), .A(n4814), .Z(n4811) );
  AND U5831 ( .A(a[67]), .B(b[9]), .Z(n4810) );
  XOR U5832 ( .A(n4815), .B(n4816), .Z(n4732) );
  ANDN U5833 ( .B(n4817), .A(n4818), .Z(n4815) );
  XNOR U5834 ( .A(n4819), .B(n4737), .Z(n4739) );
  XOR U5835 ( .A(n4820), .B(n4821), .Z(n4737) );
  ANDN U5836 ( .B(n4822), .A(n4823), .Z(n4820) );
  AND U5837 ( .A(a[68]), .B(b[8]), .Z(n4819) );
  XOR U5838 ( .A(n4825), .B(n4826), .Z(n4742) );
  ANDN U5839 ( .B(n4827), .A(n4828), .Z(n4825) );
  AND U5840 ( .A(a[70]), .B(b[6]), .Z(n4824) );
  XOR U5841 ( .A(n4830), .B(n4831), .Z(n4747) );
  ANDN U5842 ( .B(n4832), .A(n4833), .Z(n4830) );
  AND U5843 ( .A(a[71]), .B(b[5]), .Z(n4829) );
  XOR U5844 ( .A(n4835), .B(n4836), .Z(n4752) );
  ANDN U5845 ( .B(n4764), .A(n4773), .Z(n4835) );
  AND U5846 ( .A(a[72]), .B(b[3]), .Z(n4837) );
  XNOR U5847 ( .A(n4832), .B(n4836), .Z(n4838) );
  XOR U5848 ( .A(n4839), .B(n4840), .Z(n4836) );
  ANDN U5849 ( .B(n4769), .A(n4770), .Z(n4839) );
  AND U5850 ( .A(b[2]), .B(a[72]), .Z(n4841) );
  XNOR U5851 ( .A(n4843), .B(n4840), .Z(n4842) );
  XOR U5852 ( .A(n4844), .B(n4845), .Z(n4840) );
  NANDN U5853 ( .A(n4772), .B(n4771), .Z(n4845) );
  XOR U5854 ( .A(n4844), .B(n4846), .Z(n4771) );
  NAND U5855 ( .A(a[72]), .B(b[1]), .Z(n4846) );
  XOR U5856 ( .A(n4844), .B(n4848), .Z(n4847) );
  OR U5857 ( .A(n2537), .B(n2535), .Z(n4844) );
  XOR U5858 ( .A(n4850), .B(n4851), .Z(n2535) );
  NANDN U5859 ( .A(n179), .B(a[72]), .Z(n2537) );
  XNOR U5860 ( .A(n4827), .B(n4831), .Z(n4853) );
  XNOR U5861 ( .A(n4817), .B(n4826), .Z(n4854) );
  XOR U5862 ( .A(n4855), .B(n4816), .Z(n4817) );
  AND U5863 ( .A(b[6]), .B(a[69]), .Z(n4855) );
  XNOR U5864 ( .A(n4816), .B(n4822), .Z(n4856) );
  XNOR U5865 ( .A(n4821), .B(n4813), .Z(n4857) );
  XNOR U5866 ( .A(n4812), .B(n4808), .Z(n4858) );
  XNOR U5867 ( .A(n4807), .B(n4803), .Z(n4859) );
  XNOR U5868 ( .A(n4802), .B(n4798), .Z(n4860) );
  XOR U5869 ( .A(n4797), .B(n4794), .Z(n4861) );
  XOR U5870 ( .A(n4862), .B(n4863), .Z(n4794) );
  XOR U5871 ( .A(n4792), .B(n4864), .Z(n4863) );
  XOR U5872 ( .A(n4865), .B(n4866), .Z(n4864) );
  XOR U5873 ( .A(n4867), .B(n4868), .Z(n4866) );
  NAND U5874 ( .A(a[61]), .B(b[14]), .Z(n4868) );
  AND U5875 ( .A(a[60]), .B(b[15]), .Z(n4867) );
  XOR U5876 ( .A(n4869), .B(n4865), .Z(n4862) );
  XOR U5877 ( .A(n4870), .B(n4871), .Z(n4865) );
  NOR U5878 ( .A(n4872), .B(n4873), .Z(n4870) );
  AND U5879 ( .A(a[62]), .B(b[13]), .Z(n4869) );
  XNOR U5880 ( .A(n4874), .B(n4792), .Z(n4793) );
  XOR U5881 ( .A(n4875), .B(n4876), .Z(n4792) );
  ANDN U5882 ( .B(n4877), .A(n4878), .Z(n4875) );
  AND U5883 ( .A(a[63]), .B(b[12]), .Z(n4874) );
  XNOR U5884 ( .A(n4879), .B(n4797), .Z(n4799) );
  XOR U5885 ( .A(n4880), .B(n4881), .Z(n4797) );
  ANDN U5886 ( .B(n4882), .A(n4883), .Z(n4880) );
  AND U5887 ( .A(a[64]), .B(b[11]), .Z(n4879) );
  XNOR U5888 ( .A(n4884), .B(n4802), .Z(n4804) );
  XOR U5889 ( .A(n4885), .B(n4886), .Z(n4802) );
  ANDN U5890 ( .B(n4887), .A(n4888), .Z(n4885) );
  AND U5891 ( .A(a[65]), .B(b[10]), .Z(n4884) );
  XNOR U5892 ( .A(n4889), .B(n4807), .Z(n4809) );
  XOR U5893 ( .A(n4890), .B(n4891), .Z(n4807) );
  ANDN U5894 ( .B(n4892), .A(n4893), .Z(n4890) );
  AND U5895 ( .A(a[66]), .B(b[9]), .Z(n4889) );
  XNOR U5896 ( .A(n4894), .B(n4812), .Z(n4814) );
  XOR U5897 ( .A(n4895), .B(n4896), .Z(n4812) );
  ANDN U5898 ( .B(n4897), .A(n4898), .Z(n4895) );
  AND U5899 ( .A(a[67]), .B(b[8]), .Z(n4894) );
  XOR U5900 ( .A(n4899), .B(n4900), .Z(n4816) );
  ANDN U5901 ( .B(n4901), .A(n4902), .Z(n4899) );
  XNOR U5902 ( .A(n4903), .B(n4821), .Z(n4823) );
  XOR U5903 ( .A(n4904), .B(n4905), .Z(n4821) );
  ANDN U5904 ( .B(n4906), .A(n4907), .Z(n4904) );
  AND U5905 ( .A(a[68]), .B(b[7]), .Z(n4903) );
  XOR U5906 ( .A(n4909), .B(n4910), .Z(n4826) );
  ANDN U5907 ( .B(n4911), .A(n4912), .Z(n4909) );
  AND U5908 ( .A(a[70]), .B(b[5]), .Z(n4908) );
  XOR U5909 ( .A(n4914), .B(n4915), .Z(n4831) );
  ANDN U5910 ( .B(n4843), .A(n4852), .Z(n4914) );
  AND U5911 ( .A(a[71]), .B(b[3]), .Z(n4916) );
  XNOR U5912 ( .A(n4911), .B(n4915), .Z(n4917) );
  XOR U5913 ( .A(n4918), .B(n4919), .Z(n4915) );
  ANDN U5914 ( .B(n4848), .A(n4849), .Z(n4918) );
  AND U5915 ( .A(b[2]), .B(a[71]), .Z(n4920) );
  XNOR U5916 ( .A(n4922), .B(n4919), .Z(n4921) );
  XOR U5917 ( .A(n4923), .B(n4924), .Z(n4919) );
  NANDN U5918 ( .A(n4851), .B(n4850), .Z(n4924) );
  XOR U5919 ( .A(n4923), .B(n4925), .Z(n4850) );
  NAND U5920 ( .A(a[71]), .B(b[1]), .Z(n4925) );
  XOR U5921 ( .A(n4923), .B(n4927), .Z(n4926) );
  OR U5922 ( .A(n2542), .B(n2540), .Z(n4923) );
  XOR U5923 ( .A(n4929), .B(n4930), .Z(n2540) );
  NANDN U5924 ( .A(n179), .B(a[71]), .Z(n2542) );
  XNOR U5925 ( .A(n4901), .B(n4910), .Z(n4932) );
  XOR U5926 ( .A(n4933), .B(n4900), .Z(n4901) );
  AND U5927 ( .A(b[5]), .B(a[69]), .Z(n4933) );
  XNOR U5928 ( .A(n4900), .B(n4906), .Z(n4934) );
  XNOR U5929 ( .A(n4905), .B(n4897), .Z(n4935) );
  XNOR U5930 ( .A(n4896), .B(n4892), .Z(n4936) );
  XNOR U5931 ( .A(n4891), .B(n4887), .Z(n4937) );
  XNOR U5932 ( .A(n4886), .B(n4882), .Z(n4938) );
  XNOR U5933 ( .A(n4881), .B(n4877), .Z(n4939) );
  XOR U5934 ( .A(n4876), .B(n4873), .Z(n4940) );
  XOR U5935 ( .A(n4941), .B(n4942), .Z(n4873) );
  XOR U5936 ( .A(n4871), .B(n4943), .Z(n4942) );
  XOR U5937 ( .A(n4944), .B(n4945), .Z(n4943) );
  XOR U5938 ( .A(n4946), .B(n4947), .Z(n4945) );
  NAND U5939 ( .A(a[60]), .B(b[14]), .Z(n4947) );
  AND U5940 ( .A(a[59]), .B(b[15]), .Z(n4946) );
  XOR U5941 ( .A(n4948), .B(n4944), .Z(n4941) );
  XOR U5942 ( .A(n4949), .B(n4950), .Z(n4944) );
  NOR U5943 ( .A(n4951), .B(n4952), .Z(n4949) );
  AND U5944 ( .A(a[61]), .B(b[13]), .Z(n4948) );
  XNOR U5945 ( .A(n4953), .B(n4871), .Z(n4872) );
  XOR U5946 ( .A(n4954), .B(n4955), .Z(n4871) );
  ANDN U5947 ( .B(n4956), .A(n4957), .Z(n4954) );
  AND U5948 ( .A(a[62]), .B(b[12]), .Z(n4953) );
  XNOR U5949 ( .A(n4958), .B(n4876), .Z(n4878) );
  XOR U5950 ( .A(n4959), .B(n4960), .Z(n4876) );
  ANDN U5951 ( .B(n4961), .A(n4962), .Z(n4959) );
  AND U5952 ( .A(a[63]), .B(b[11]), .Z(n4958) );
  XNOR U5953 ( .A(n4963), .B(n4881), .Z(n4883) );
  XOR U5954 ( .A(n4964), .B(n4965), .Z(n4881) );
  ANDN U5955 ( .B(n4966), .A(n4967), .Z(n4964) );
  AND U5956 ( .A(a[64]), .B(b[10]), .Z(n4963) );
  XNOR U5957 ( .A(n4968), .B(n4886), .Z(n4888) );
  XOR U5958 ( .A(n4969), .B(n4970), .Z(n4886) );
  ANDN U5959 ( .B(n4971), .A(n4972), .Z(n4969) );
  AND U5960 ( .A(a[65]), .B(b[9]), .Z(n4968) );
  XNOR U5961 ( .A(n4973), .B(n4891), .Z(n4893) );
  XOR U5962 ( .A(n4974), .B(n4975), .Z(n4891) );
  ANDN U5963 ( .B(n4976), .A(n4977), .Z(n4974) );
  AND U5964 ( .A(a[66]), .B(b[8]), .Z(n4973) );
  XNOR U5965 ( .A(n4978), .B(n4896), .Z(n4898) );
  XOR U5966 ( .A(n4979), .B(n4980), .Z(n4896) );
  ANDN U5967 ( .B(n4981), .A(n4982), .Z(n4979) );
  AND U5968 ( .A(a[67]), .B(b[7]), .Z(n4978) );
  XOR U5969 ( .A(n4983), .B(n4984), .Z(n4900) );
  ANDN U5970 ( .B(n4985), .A(n4986), .Z(n4983) );
  XNOR U5971 ( .A(n4987), .B(n4905), .Z(n4907) );
  XOR U5972 ( .A(n4988), .B(n4989), .Z(n4905) );
  ANDN U5973 ( .B(n4990), .A(n4991), .Z(n4988) );
  AND U5974 ( .A(a[68]), .B(b[6]), .Z(n4987) );
  XOR U5975 ( .A(n4993), .B(n4994), .Z(n4910) );
  ANDN U5976 ( .B(n4922), .A(n4931), .Z(n4993) );
  AND U5977 ( .A(a[70]), .B(b[3]), .Z(n4995) );
  XNOR U5978 ( .A(n4985), .B(n4994), .Z(n4996) );
  XOR U5979 ( .A(n4997), .B(n4998), .Z(n4994) );
  ANDN U5980 ( .B(n4927), .A(n4928), .Z(n4997) );
  AND U5981 ( .A(b[2]), .B(a[70]), .Z(n4999) );
  XNOR U5982 ( .A(n5001), .B(n4998), .Z(n5000) );
  XOR U5983 ( .A(n5002), .B(n5003), .Z(n4998) );
  NANDN U5984 ( .A(n4930), .B(n4929), .Z(n5003) );
  XOR U5985 ( .A(n5002), .B(n5004), .Z(n4929) );
  NAND U5986 ( .A(a[70]), .B(b[1]), .Z(n5004) );
  XNOR U5987 ( .A(n5002), .B(n5006), .Z(n5005) );
  OR U5988 ( .A(n2547), .B(n2545), .Z(n5002) );
  NANDN U5989 ( .A(n179), .B(a[70]), .Z(n2547) );
  XOR U5990 ( .A(n5011), .B(n4984), .Z(n4985) );
  AND U5991 ( .A(b[4]), .B(a[69]), .Z(n5011) );
  XNOR U5992 ( .A(n4984), .B(n4990), .Z(n5012) );
  XNOR U5993 ( .A(n4989), .B(n4981), .Z(n5013) );
  XNOR U5994 ( .A(n4980), .B(n4976), .Z(n5014) );
  XNOR U5995 ( .A(n4975), .B(n4971), .Z(n5015) );
  XNOR U5996 ( .A(n4970), .B(n4966), .Z(n5016) );
  XNOR U5997 ( .A(n4965), .B(n4961), .Z(n5017) );
  XNOR U5998 ( .A(n4960), .B(n4956), .Z(n5018) );
  XOR U5999 ( .A(n4955), .B(n4952), .Z(n5019) );
  XOR U6000 ( .A(n5020), .B(n5021), .Z(n4952) );
  XOR U6001 ( .A(n4950), .B(n5022), .Z(n5021) );
  XOR U6002 ( .A(n5023), .B(n5024), .Z(n5022) );
  XOR U6003 ( .A(n5025), .B(n5026), .Z(n5024) );
  NAND U6004 ( .A(a[59]), .B(b[14]), .Z(n5026) );
  AND U6005 ( .A(a[58]), .B(b[15]), .Z(n5025) );
  XOR U6006 ( .A(n5027), .B(n5023), .Z(n5020) );
  XOR U6007 ( .A(n5028), .B(n5029), .Z(n5023) );
  NOR U6008 ( .A(n5030), .B(n5031), .Z(n5028) );
  AND U6009 ( .A(a[60]), .B(b[13]), .Z(n5027) );
  XNOR U6010 ( .A(n5032), .B(n4950), .Z(n4951) );
  XOR U6011 ( .A(n5033), .B(n5034), .Z(n4950) );
  ANDN U6012 ( .B(n5035), .A(n5036), .Z(n5033) );
  AND U6013 ( .A(a[61]), .B(b[12]), .Z(n5032) );
  XNOR U6014 ( .A(n5037), .B(n4955), .Z(n4957) );
  XOR U6015 ( .A(n5038), .B(n5039), .Z(n4955) );
  ANDN U6016 ( .B(n5040), .A(n5041), .Z(n5038) );
  AND U6017 ( .A(a[62]), .B(b[11]), .Z(n5037) );
  XNOR U6018 ( .A(n5042), .B(n4960), .Z(n4962) );
  XOR U6019 ( .A(n5043), .B(n5044), .Z(n4960) );
  ANDN U6020 ( .B(n5045), .A(n5046), .Z(n5043) );
  AND U6021 ( .A(a[63]), .B(b[10]), .Z(n5042) );
  XNOR U6022 ( .A(n5047), .B(n4965), .Z(n4967) );
  XOR U6023 ( .A(n5048), .B(n5049), .Z(n4965) );
  ANDN U6024 ( .B(n5050), .A(n5051), .Z(n5048) );
  AND U6025 ( .A(a[64]), .B(b[9]), .Z(n5047) );
  XNOR U6026 ( .A(n5052), .B(n4970), .Z(n4972) );
  XOR U6027 ( .A(n5053), .B(n5054), .Z(n4970) );
  ANDN U6028 ( .B(n5055), .A(n5056), .Z(n5053) );
  AND U6029 ( .A(a[65]), .B(b[8]), .Z(n5052) );
  XNOR U6030 ( .A(n5057), .B(n4975), .Z(n4977) );
  XOR U6031 ( .A(n5058), .B(n5059), .Z(n4975) );
  ANDN U6032 ( .B(n5060), .A(n5061), .Z(n5058) );
  AND U6033 ( .A(a[66]), .B(b[7]), .Z(n5057) );
  XNOR U6034 ( .A(n5062), .B(n4980), .Z(n4982) );
  XOR U6035 ( .A(n5063), .B(n5064), .Z(n4980) );
  ANDN U6036 ( .B(n5065), .A(n5066), .Z(n5063) );
  AND U6037 ( .A(a[67]), .B(b[6]), .Z(n5062) );
  XOR U6038 ( .A(n5067), .B(n5068), .Z(n4984) );
  ANDN U6039 ( .B(n5001), .A(n5010), .Z(n5067) );
  XNOR U6040 ( .A(n5068), .B(n5070), .Z(n5069) );
  XOR U6041 ( .A(n5072), .B(n5068), .Z(n5001) );
  XNOR U6042 ( .A(n5073), .B(n5074), .Z(n5068) );
  NOR U6043 ( .A(n5007), .B(n5006), .Z(n5073) );
  XOR U6044 ( .A(n5075), .B(n5074), .Z(n5006) );
  AND U6045 ( .A(b[2]), .B(a[69]), .Z(n5075) );
  XOR U6046 ( .A(n5074), .B(n5077), .Z(n5076) );
  XNOR U6047 ( .A(n5078), .B(n5079), .Z(n5074) );
  OR U6048 ( .A(n5008), .B(n5009), .Z(n5079) );
  XNOR U6049 ( .A(n5078), .B(n5081), .Z(n5080) );
  XNOR U6050 ( .A(n5078), .B(n5083), .Z(n5008) );
  NAND U6051 ( .A(b[1]), .B(a[69]), .Z(n5083) );
  OR U6052 ( .A(n2552), .B(n2550), .Z(n5078) );
  XOR U6053 ( .A(n5084), .B(n5085), .Z(n2550) );
  NANDN U6054 ( .A(n179), .B(a[69]), .Z(n2552) );
  AND U6055 ( .A(b[3]), .B(a[69]), .Z(n5072) );
  XNOR U6056 ( .A(n5087), .B(n4989), .Z(n4991) );
  XOR U6057 ( .A(n5088), .B(n5089), .Z(n4989) );
  ANDN U6058 ( .B(n5070), .A(n5071), .Z(n5088) );
  XNOR U6059 ( .A(n5090), .B(n5089), .Z(n5071) );
  AND U6060 ( .A(a[68]), .B(b[4]), .Z(n5090) );
  XNOR U6061 ( .A(n5089), .B(n5065), .Z(n5091) );
  XNOR U6062 ( .A(n5064), .B(n5060), .Z(n5092) );
  XNOR U6063 ( .A(n5059), .B(n5055), .Z(n5093) );
  XNOR U6064 ( .A(n5054), .B(n5050), .Z(n5094) );
  XNOR U6065 ( .A(n5049), .B(n5045), .Z(n5095) );
  XNOR U6066 ( .A(n5044), .B(n5040), .Z(n5096) );
  XNOR U6067 ( .A(n5039), .B(n5035), .Z(n5097) );
  XOR U6068 ( .A(n5034), .B(n5031), .Z(n5098) );
  XOR U6069 ( .A(n5099), .B(n5100), .Z(n5031) );
  XOR U6070 ( .A(n5029), .B(n5101), .Z(n5100) );
  XOR U6071 ( .A(n5102), .B(n5103), .Z(n5101) );
  XOR U6072 ( .A(n5104), .B(n5105), .Z(n5103) );
  NAND U6073 ( .A(a[58]), .B(b[14]), .Z(n5105) );
  AND U6074 ( .A(a[57]), .B(b[15]), .Z(n5104) );
  XOR U6075 ( .A(n5106), .B(n5102), .Z(n5099) );
  XOR U6076 ( .A(n5107), .B(n5108), .Z(n5102) );
  NOR U6077 ( .A(n5109), .B(n5110), .Z(n5107) );
  AND U6078 ( .A(a[59]), .B(b[13]), .Z(n5106) );
  XNOR U6079 ( .A(n5111), .B(n5029), .Z(n5030) );
  XOR U6080 ( .A(n5112), .B(n5113), .Z(n5029) );
  ANDN U6081 ( .B(n5114), .A(n5115), .Z(n5112) );
  AND U6082 ( .A(a[60]), .B(b[12]), .Z(n5111) );
  XNOR U6083 ( .A(n5116), .B(n5034), .Z(n5036) );
  XOR U6084 ( .A(n5117), .B(n5118), .Z(n5034) );
  ANDN U6085 ( .B(n5119), .A(n5120), .Z(n5117) );
  AND U6086 ( .A(a[61]), .B(b[11]), .Z(n5116) );
  XNOR U6087 ( .A(n5121), .B(n5039), .Z(n5041) );
  XOR U6088 ( .A(n5122), .B(n5123), .Z(n5039) );
  ANDN U6089 ( .B(n5124), .A(n5125), .Z(n5122) );
  AND U6090 ( .A(a[62]), .B(b[10]), .Z(n5121) );
  XNOR U6091 ( .A(n5126), .B(n5044), .Z(n5046) );
  XOR U6092 ( .A(n5127), .B(n5128), .Z(n5044) );
  ANDN U6093 ( .B(n5129), .A(n5130), .Z(n5127) );
  AND U6094 ( .A(a[63]), .B(b[9]), .Z(n5126) );
  XNOR U6095 ( .A(n5131), .B(n5049), .Z(n5051) );
  XOR U6096 ( .A(n5132), .B(n5133), .Z(n5049) );
  ANDN U6097 ( .B(n5134), .A(n5135), .Z(n5132) );
  AND U6098 ( .A(a[64]), .B(b[8]), .Z(n5131) );
  XNOR U6099 ( .A(n5136), .B(n5054), .Z(n5056) );
  XOR U6100 ( .A(n5137), .B(n5138), .Z(n5054) );
  ANDN U6101 ( .B(n5139), .A(n5140), .Z(n5137) );
  AND U6102 ( .A(a[65]), .B(b[7]), .Z(n5136) );
  XNOR U6103 ( .A(n5141), .B(n5059), .Z(n5061) );
  XOR U6104 ( .A(n5142), .B(n5143), .Z(n5059) );
  ANDN U6105 ( .B(n5144), .A(n5145), .Z(n5142) );
  AND U6106 ( .A(a[66]), .B(b[6]), .Z(n5141) );
  XOR U6107 ( .A(n5146), .B(n5147), .Z(n5089) );
  ANDN U6108 ( .B(n5077), .A(n5086), .Z(n5146) );
  XNOR U6109 ( .A(n5148), .B(n5147), .Z(n5086) );
  AND U6110 ( .A(a[68]), .B(b[3]), .Z(n5148) );
  XNOR U6111 ( .A(n5147), .B(n5150), .Z(n5149) );
  XNOR U6112 ( .A(n5151), .B(n5152), .Z(n5147) );
  NOR U6113 ( .A(n5082), .B(n5081), .Z(n5151) );
  XOR U6114 ( .A(n5153), .B(n5152), .Z(n5081) );
  AND U6115 ( .A(b[2]), .B(a[68]), .Z(n5153) );
  XOR U6116 ( .A(n5152), .B(n5155), .Z(n5154) );
  XNOR U6117 ( .A(n5156), .B(n5157), .Z(n5152) );
  NANDN U6118 ( .A(n5085), .B(n5084), .Z(n5157) );
  XOR U6119 ( .A(n5156), .B(n5158), .Z(n5084) );
  NAND U6120 ( .A(a[68]), .B(b[1]), .Z(n5158) );
  XOR U6121 ( .A(n5156), .B(n5160), .Z(n5159) );
  OR U6122 ( .A(n2557), .B(n2555), .Z(n5156) );
  XOR U6123 ( .A(n5162), .B(n5163), .Z(n2555) );
  NANDN U6124 ( .A(n179), .B(a[68]), .Z(n2557) );
  XNOR U6125 ( .A(n5166), .B(n5064), .Z(n5066) );
  XOR U6126 ( .A(n5167), .B(n5168), .Z(n5064) );
  ANDN U6127 ( .B(n5150), .A(n5165), .Z(n5167) );
  XNOR U6128 ( .A(n5169), .B(n5168), .Z(n5165) );
  AND U6129 ( .A(a[67]), .B(b[4]), .Z(n5169) );
  XNOR U6130 ( .A(n5168), .B(n5144), .Z(n5170) );
  XNOR U6131 ( .A(n5143), .B(n5139), .Z(n5171) );
  XNOR U6132 ( .A(n5138), .B(n5134), .Z(n5172) );
  XNOR U6133 ( .A(n5133), .B(n5129), .Z(n5173) );
  XNOR U6134 ( .A(n5128), .B(n5124), .Z(n5174) );
  XNOR U6135 ( .A(n5123), .B(n5119), .Z(n5175) );
  XNOR U6136 ( .A(n5118), .B(n5114), .Z(n5176) );
  XOR U6137 ( .A(n5113), .B(n5110), .Z(n5177) );
  XOR U6138 ( .A(n5178), .B(n5179), .Z(n5110) );
  XOR U6139 ( .A(n5108), .B(n5180), .Z(n5179) );
  XOR U6140 ( .A(n5181), .B(n5182), .Z(n5180) );
  XOR U6141 ( .A(n5183), .B(n5184), .Z(n5182) );
  NAND U6142 ( .A(a[57]), .B(b[14]), .Z(n5184) );
  AND U6143 ( .A(a[56]), .B(b[15]), .Z(n5183) );
  XOR U6144 ( .A(n5185), .B(n5181), .Z(n5178) );
  XOR U6145 ( .A(n5186), .B(n5187), .Z(n5181) );
  NOR U6146 ( .A(n5188), .B(n5189), .Z(n5186) );
  AND U6147 ( .A(a[58]), .B(b[13]), .Z(n5185) );
  XNOR U6148 ( .A(n5190), .B(n5108), .Z(n5109) );
  XOR U6149 ( .A(n5191), .B(n5192), .Z(n5108) );
  ANDN U6150 ( .B(n5193), .A(n5194), .Z(n5191) );
  AND U6151 ( .A(a[59]), .B(b[12]), .Z(n5190) );
  XNOR U6152 ( .A(n5195), .B(n5113), .Z(n5115) );
  XOR U6153 ( .A(n5196), .B(n5197), .Z(n5113) );
  ANDN U6154 ( .B(n5198), .A(n5199), .Z(n5196) );
  AND U6155 ( .A(a[60]), .B(b[11]), .Z(n5195) );
  XNOR U6156 ( .A(n5200), .B(n5118), .Z(n5120) );
  XOR U6157 ( .A(n5201), .B(n5202), .Z(n5118) );
  ANDN U6158 ( .B(n5203), .A(n5204), .Z(n5201) );
  AND U6159 ( .A(a[61]), .B(b[10]), .Z(n5200) );
  XNOR U6160 ( .A(n5205), .B(n5123), .Z(n5125) );
  XOR U6161 ( .A(n5206), .B(n5207), .Z(n5123) );
  ANDN U6162 ( .B(n5208), .A(n5209), .Z(n5206) );
  AND U6163 ( .A(a[62]), .B(b[9]), .Z(n5205) );
  XNOR U6164 ( .A(n5210), .B(n5128), .Z(n5130) );
  XOR U6165 ( .A(n5211), .B(n5212), .Z(n5128) );
  ANDN U6166 ( .B(n5213), .A(n5214), .Z(n5211) );
  AND U6167 ( .A(a[63]), .B(b[8]), .Z(n5210) );
  XNOR U6168 ( .A(n5215), .B(n5133), .Z(n5135) );
  XOR U6169 ( .A(n5216), .B(n5217), .Z(n5133) );
  ANDN U6170 ( .B(n5218), .A(n5219), .Z(n5216) );
  AND U6171 ( .A(a[64]), .B(b[7]), .Z(n5215) );
  XNOR U6172 ( .A(n5220), .B(n5138), .Z(n5140) );
  XOR U6173 ( .A(n5221), .B(n5222), .Z(n5138) );
  ANDN U6174 ( .B(n5223), .A(n5224), .Z(n5221) );
  AND U6175 ( .A(a[65]), .B(b[6]), .Z(n5220) );
  XOR U6176 ( .A(n5225), .B(n5226), .Z(n5168) );
  ANDN U6177 ( .B(n5155), .A(n5164), .Z(n5225) );
  XNOR U6178 ( .A(n5227), .B(n5226), .Z(n5164) );
  AND U6179 ( .A(a[67]), .B(b[3]), .Z(n5227) );
  XNOR U6180 ( .A(n5226), .B(n5229), .Z(n5228) );
  XNOR U6181 ( .A(n5230), .B(n5231), .Z(n5226) );
  ANDN U6182 ( .B(n5160), .A(n5161), .Z(n5230) );
  XOR U6183 ( .A(n5232), .B(n5231), .Z(n5161) );
  IV U6184 ( .A(n5233), .Z(n5231) );
  AND U6185 ( .A(b[2]), .B(a[67]), .Z(n5232) );
  XNOR U6186 ( .A(n5235), .B(n5233), .Z(n5234) );
  XOR U6187 ( .A(n5236), .B(n5237), .Z(n5233) );
  NANDN U6188 ( .A(n5163), .B(n5162), .Z(n5237) );
  XOR U6189 ( .A(n5236), .B(n5238), .Z(n5162) );
  NAND U6190 ( .A(a[67]), .B(b[1]), .Z(n5238) );
  XOR U6191 ( .A(n5236), .B(n5240), .Z(n5239) );
  OR U6192 ( .A(n2562), .B(n2560), .Z(n5236) );
  XOR U6193 ( .A(n5242), .B(n5243), .Z(n2560) );
  NANDN U6194 ( .A(n179), .B(a[67]), .Z(n2562) );
  XNOR U6195 ( .A(n5246), .B(n5143), .Z(n5145) );
  XOR U6196 ( .A(n5247), .B(n5248), .Z(n5143) );
  ANDN U6197 ( .B(n5229), .A(n5245), .Z(n5247) );
  XNOR U6198 ( .A(n5249), .B(n5248), .Z(n5245) );
  AND U6199 ( .A(a[66]), .B(b[4]), .Z(n5249) );
  XNOR U6200 ( .A(n5248), .B(n5223), .Z(n5250) );
  XNOR U6201 ( .A(n5222), .B(n5218), .Z(n5251) );
  XNOR U6202 ( .A(n5217), .B(n5213), .Z(n5252) );
  XNOR U6203 ( .A(n5212), .B(n5208), .Z(n5253) );
  XNOR U6204 ( .A(n5207), .B(n5203), .Z(n5254) );
  XNOR U6205 ( .A(n5202), .B(n5198), .Z(n5255) );
  XNOR U6206 ( .A(n5197), .B(n5193), .Z(n5256) );
  XOR U6207 ( .A(n5192), .B(n5189), .Z(n5257) );
  XOR U6208 ( .A(n5258), .B(n5259), .Z(n5189) );
  XOR U6209 ( .A(n5187), .B(n5260), .Z(n5259) );
  XNOR U6210 ( .A(n5261), .B(n5262), .Z(n5260) );
  XOR U6211 ( .A(n5263), .B(n5264), .Z(n5262) );
  NAND U6212 ( .A(a[56]), .B(b[14]), .Z(n5264) );
  AND U6213 ( .A(a[55]), .B(b[15]), .Z(n5263) );
  XNOR U6214 ( .A(n5265), .B(n5261), .Z(n5258) );
  XOR U6215 ( .A(n5266), .B(n5267), .Z(n5261) );
  NOR U6216 ( .A(n5268), .B(n5269), .Z(n5266) );
  AND U6217 ( .A(a[57]), .B(b[13]), .Z(n5265) );
  XNOR U6218 ( .A(n5270), .B(n5187), .Z(n5188) );
  XNOR U6219 ( .A(n5271), .B(n5272), .Z(n5187) );
  ANDN U6220 ( .B(n5273), .A(n5274), .Z(n5271) );
  AND U6221 ( .A(a[58]), .B(b[12]), .Z(n5270) );
  XNOR U6222 ( .A(n5275), .B(n5192), .Z(n5194) );
  XNOR U6223 ( .A(n5276), .B(n5277), .Z(n5192) );
  ANDN U6224 ( .B(n5278), .A(n5279), .Z(n5276) );
  AND U6225 ( .A(a[59]), .B(b[11]), .Z(n5275) );
  XNOR U6226 ( .A(n5280), .B(n5197), .Z(n5199) );
  XNOR U6227 ( .A(n5281), .B(n5282), .Z(n5197) );
  ANDN U6228 ( .B(n5283), .A(n5284), .Z(n5281) );
  AND U6229 ( .A(a[60]), .B(b[10]), .Z(n5280) );
  XNOR U6230 ( .A(n5285), .B(n5202), .Z(n5204) );
  XNOR U6231 ( .A(n5286), .B(n5287), .Z(n5202) );
  ANDN U6232 ( .B(n5288), .A(n5289), .Z(n5286) );
  AND U6233 ( .A(a[61]), .B(b[9]), .Z(n5285) );
  XNOR U6234 ( .A(n5290), .B(n5207), .Z(n5209) );
  XNOR U6235 ( .A(n5291), .B(n5292), .Z(n5207) );
  ANDN U6236 ( .B(n5293), .A(n5294), .Z(n5291) );
  AND U6237 ( .A(a[62]), .B(b[8]), .Z(n5290) );
  XNOR U6238 ( .A(n5295), .B(n5212), .Z(n5214) );
  XNOR U6239 ( .A(n5296), .B(n5297), .Z(n5212) );
  ANDN U6240 ( .B(n5298), .A(n5299), .Z(n5296) );
  AND U6241 ( .A(a[63]), .B(b[7]), .Z(n5295) );
  XNOR U6242 ( .A(n5300), .B(n5217), .Z(n5219) );
  XNOR U6243 ( .A(n5301), .B(n5302), .Z(n5217) );
  ANDN U6244 ( .B(n5303), .A(n5304), .Z(n5301) );
  AND U6245 ( .A(a[64]), .B(b[6]), .Z(n5300) );
  XNOR U6246 ( .A(n5305), .B(n5306), .Z(n5248) );
  ANDN U6247 ( .B(n5235), .A(n5244), .Z(n5305) );
  XOR U6248 ( .A(n5307), .B(n5306), .Z(n5244) );
  IV U6249 ( .A(n5308), .Z(n5306) );
  AND U6250 ( .A(a[66]), .B(b[3]), .Z(n5307) );
  XNOR U6251 ( .A(n5310), .B(n5308), .Z(n5309) );
  XOR U6252 ( .A(n5311), .B(n5312), .Z(n5308) );
  ANDN U6253 ( .B(n5240), .A(n5241), .Z(n5311) );
  AND U6254 ( .A(b[2]), .B(a[66]), .Z(n5313) );
  XNOR U6255 ( .A(n5315), .B(n5312), .Z(n5314) );
  XOR U6256 ( .A(n5316), .B(n5317), .Z(n5312) );
  NANDN U6257 ( .A(n5243), .B(n5242), .Z(n5317) );
  XOR U6258 ( .A(n5316), .B(n5318), .Z(n5242) );
  NAND U6259 ( .A(a[66]), .B(b[1]), .Z(n5318) );
  XOR U6260 ( .A(n5316), .B(n5320), .Z(n5319) );
  OR U6261 ( .A(n2567), .B(n2565), .Z(n5316) );
  XOR U6262 ( .A(n5322), .B(n5323), .Z(n2565) );
  NANDN U6263 ( .A(n179), .B(a[66]), .Z(n2567) );
  XNOR U6264 ( .A(n5326), .B(n5222), .Z(n5224) );
  XNOR U6265 ( .A(n5327), .B(n5328), .Z(n5222) );
  ANDN U6266 ( .B(n5310), .A(n5325), .Z(n5327) );
  XOR U6267 ( .A(n5329), .B(n5328), .Z(n5325) );
  IV U6268 ( .A(n5330), .Z(n5328) );
  AND U6269 ( .A(a[65]), .B(b[4]), .Z(n5329) );
  XNOR U6270 ( .A(n5303), .B(n5330), .Z(n5331) );
  XOR U6271 ( .A(n5332), .B(n5333), .Z(n5330) );
  ANDN U6272 ( .B(n5315), .A(n5324), .Z(n5332) );
  AND U6273 ( .A(a[65]), .B(b[3]), .Z(n5334) );
  XNOR U6274 ( .A(n5336), .B(n5333), .Z(n5335) );
  XOR U6275 ( .A(n5337), .B(n5338), .Z(n5333) );
  ANDN U6276 ( .B(n5320), .A(n5321), .Z(n5337) );
  AND U6277 ( .A(b[2]), .B(a[65]), .Z(n5339) );
  XNOR U6278 ( .A(n5341), .B(n5338), .Z(n5340) );
  XOR U6279 ( .A(n5342), .B(n5343), .Z(n5338) );
  NANDN U6280 ( .A(n5323), .B(n5322), .Z(n5343) );
  XOR U6281 ( .A(n5342), .B(n5344), .Z(n5322) );
  NAND U6282 ( .A(a[65]), .B(b[1]), .Z(n5344) );
  XOR U6283 ( .A(n5342), .B(n5346), .Z(n5345) );
  OR U6284 ( .A(n2572), .B(n2570), .Z(n5342) );
  XOR U6285 ( .A(n5348), .B(n5349), .Z(n2570) );
  NANDN U6286 ( .A(n179), .B(a[65]), .Z(n2572) );
  XNOR U6287 ( .A(n5298), .B(n5353), .Z(n5352) );
  XNOR U6288 ( .A(n5293), .B(n5355), .Z(n5354) );
  XNOR U6289 ( .A(n5288), .B(n5357), .Z(n5356) );
  XNOR U6290 ( .A(n5283), .B(n5359), .Z(n5358) );
  XNOR U6291 ( .A(n5278), .B(n5361), .Z(n5360) );
  XNOR U6292 ( .A(n5273), .B(n5363), .Z(n5362) );
  XOR U6293 ( .A(n5269), .B(n5365), .Z(n5364) );
  XOR U6294 ( .A(n5366), .B(n5367), .Z(n5269) );
  XNOR U6295 ( .A(n5368), .B(n5369), .Z(n5367) );
  XNOR U6296 ( .A(n5370), .B(n5371), .Z(n5368) );
  XOR U6297 ( .A(n5372), .B(n5373), .Z(n5371) );
  AND U6298 ( .A(b[15]), .B(a[54]), .Z(n5373) );
  AND U6299 ( .A(a[55]), .B(b[14]), .Z(n5372) );
  XNOR U6300 ( .A(n5374), .B(n5370), .Z(n5366) );
  XOR U6301 ( .A(n5375), .B(n5376), .Z(n5370) );
  NOR U6302 ( .A(n5377), .B(n5378), .Z(n5375) );
  AND U6303 ( .A(a[56]), .B(b[13]), .Z(n5374) );
  XOR U6304 ( .A(n5379), .B(n5267), .Z(n5268) );
  IV U6305 ( .A(n5369), .Z(n5267) );
  XOR U6306 ( .A(n5380), .B(n5381), .Z(n5369) );
  ANDN U6307 ( .B(n5382), .A(n5383), .Z(n5380) );
  AND U6308 ( .A(a[57]), .B(b[12]), .Z(n5379) );
  XOR U6309 ( .A(n5384), .B(n5272), .Z(n5274) );
  IV U6310 ( .A(n5365), .Z(n5272) );
  XOR U6311 ( .A(n5385), .B(n5386), .Z(n5365) );
  ANDN U6312 ( .B(n5387), .A(n5388), .Z(n5385) );
  AND U6313 ( .A(a[58]), .B(b[11]), .Z(n5384) );
  XOR U6314 ( .A(n5389), .B(n5277), .Z(n5279) );
  IV U6315 ( .A(n5363), .Z(n5277) );
  XOR U6316 ( .A(n5390), .B(n5391), .Z(n5363) );
  ANDN U6317 ( .B(n5392), .A(n5393), .Z(n5390) );
  AND U6318 ( .A(a[59]), .B(b[10]), .Z(n5389) );
  XOR U6319 ( .A(n5394), .B(n5282), .Z(n5284) );
  IV U6320 ( .A(n5361), .Z(n5282) );
  XOR U6321 ( .A(n5395), .B(n5396), .Z(n5361) );
  ANDN U6322 ( .B(n5397), .A(n5398), .Z(n5395) );
  AND U6323 ( .A(a[60]), .B(b[9]), .Z(n5394) );
  XOR U6324 ( .A(n5399), .B(n5287), .Z(n5289) );
  IV U6325 ( .A(n5359), .Z(n5287) );
  XOR U6326 ( .A(n5400), .B(n5401), .Z(n5359) );
  ANDN U6327 ( .B(n5402), .A(n5403), .Z(n5400) );
  AND U6328 ( .A(a[61]), .B(b[8]), .Z(n5399) );
  XOR U6329 ( .A(n5404), .B(n5292), .Z(n5294) );
  IV U6330 ( .A(n5357), .Z(n5292) );
  XOR U6331 ( .A(n5405), .B(n5406), .Z(n5357) );
  ANDN U6332 ( .B(n5407), .A(n5408), .Z(n5405) );
  AND U6333 ( .A(a[62]), .B(b[7]), .Z(n5404) );
  XOR U6334 ( .A(n5409), .B(n5297), .Z(n5299) );
  IV U6335 ( .A(n5355), .Z(n5297) );
  XOR U6336 ( .A(n5410), .B(n5411), .Z(n5355) );
  ANDN U6337 ( .B(n5412), .A(n5413), .Z(n5410) );
  AND U6338 ( .A(a[63]), .B(b[6]), .Z(n5409) );
  XOR U6339 ( .A(n5414), .B(n5302), .Z(n5304) );
  IV U6340 ( .A(n5353), .Z(n5302) );
  XOR U6341 ( .A(n5415), .B(n5416), .Z(n5353) );
  ANDN U6342 ( .B(n5336), .A(n5351), .Z(n5415) );
  AND U6343 ( .A(a[64]), .B(b[4]), .Z(n5417) );
  XNOR U6344 ( .A(n5412), .B(n5416), .Z(n5418) );
  XOR U6345 ( .A(n5419), .B(n5420), .Z(n5416) );
  ANDN U6346 ( .B(n5341), .A(n5350), .Z(n5419) );
  AND U6347 ( .A(a[64]), .B(b[3]), .Z(n5421) );
  XNOR U6348 ( .A(n5423), .B(n5420), .Z(n5422) );
  XOR U6349 ( .A(n5424), .B(n5425), .Z(n5420) );
  ANDN U6350 ( .B(n5346), .A(n5347), .Z(n5424) );
  AND U6351 ( .A(b[2]), .B(a[64]), .Z(n5426) );
  XNOR U6352 ( .A(n5428), .B(n5425), .Z(n5427) );
  XOR U6353 ( .A(n5429), .B(n5430), .Z(n5425) );
  NANDN U6354 ( .A(n5349), .B(n5348), .Z(n5430) );
  XOR U6355 ( .A(n5429), .B(n5431), .Z(n5348) );
  NAND U6356 ( .A(a[64]), .B(b[1]), .Z(n5431) );
  XOR U6357 ( .A(n5429), .B(n5433), .Z(n5432) );
  OR U6358 ( .A(n2577), .B(n2575), .Z(n5429) );
  XOR U6359 ( .A(n5435), .B(n5436), .Z(n2575) );
  NANDN U6360 ( .A(n179), .B(a[64]), .Z(n2577) );
  XNOR U6361 ( .A(n5407), .B(n5411), .Z(n5439) );
  XNOR U6362 ( .A(n5402), .B(n5406), .Z(n5440) );
  XNOR U6363 ( .A(n5397), .B(n5401), .Z(n5441) );
  XNOR U6364 ( .A(n5392), .B(n5396), .Z(n5442) );
  XNOR U6365 ( .A(n5387), .B(n5391), .Z(n5443) );
  XNOR U6366 ( .A(n5382), .B(n5386), .Z(n5444) );
  XOR U6367 ( .A(n5378), .B(n5381), .Z(n5445) );
  XOR U6368 ( .A(n5446), .B(n5447), .Z(n5378) );
  XNOR U6369 ( .A(n5448), .B(n5449), .Z(n5447) );
  XNOR U6370 ( .A(n5450), .B(n5451), .Z(n5448) );
  XOR U6371 ( .A(n5452), .B(n5453), .Z(n5451) );
  AND U6372 ( .A(b[14]), .B(a[54]), .Z(n5453) );
  AND U6373 ( .A(a[53]), .B(b[15]), .Z(n5452) );
  XNOR U6374 ( .A(n5454), .B(n5450), .Z(n5446) );
  XOR U6375 ( .A(n5455), .B(n5456), .Z(n5450) );
  NOR U6376 ( .A(n5457), .B(n5458), .Z(n5455) );
  AND U6377 ( .A(a[55]), .B(b[13]), .Z(n5454) );
  XOR U6378 ( .A(n5459), .B(n5376), .Z(n5377) );
  IV U6379 ( .A(n5449), .Z(n5376) );
  XOR U6380 ( .A(n5460), .B(n5461), .Z(n5449) );
  ANDN U6381 ( .B(n5462), .A(n5463), .Z(n5460) );
  AND U6382 ( .A(a[56]), .B(b[12]), .Z(n5459) );
  XOR U6383 ( .A(n5465), .B(n5466), .Z(n5381) );
  ANDN U6384 ( .B(n5467), .A(n5468), .Z(n5465) );
  AND U6385 ( .A(a[57]), .B(b[11]), .Z(n5464) );
  XOR U6386 ( .A(n5470), .B(n5471), .Z(n5386) );
  ANDN U6387 ( .B(n5472), .A(n5473), .Z(n5470) );
  AND U6388 ( .A(a[58]), .B(b[10]), .Z(n5469) );
  XOR U6389 ( .A(n5475), .B(n5476), .Z(n5391) );
  ANDN U6390 ( .B(n5477), .A(n5478), .Z(n5475) );
  AND U6391 ( .A(a[59]), .B(b[9]), .Z(n5474) );
  XOR U6392 ( .A(n5480), .B(n5481), .Z(n5396) );
  ANDN U6393 ( .B(n5482), .A(n5483), .Z(n5480) );
  AND U6394 ( .A(a[60]), .B(b[8]), .Z(n5479) );
  XOR U6395 ( .A(n5485), .B(n5486), .Z(n5401) );
  ANDN U6396 ( .B(n5487), .A(n5488), .Z(n5485) );
  AND U6397 ( .A(a[61]), .B(b[7]), .Z(n5484) );
  XOR U6398 ( .A(n5490), .B(n5491), .Z(n5406) );
  ANDN U6399 ( .B(n5492), .A(n5493), .Z(n5490) );
  AND U6400 ( .A(a[62]), .B(b[6]), .Z(n5489) );
  XOR U6401 ( .A(n5495), .B(n5496), .Z(n5411) );
  ANDN U6402 ( .B(n5423), .A(n5438), .Z(n5495) );
  AND U6403 ( .A(a[63]), .B(b[4]), .Z(n5497) );
  XNOR U6404 ( .A(n5492), .B(n5496), .Z(n5498) );
  XOR U6405 ( .A(n5499), .B(n5500), .Z(n5496) );
  ANDN U6406 ( .B(n5428), .A(n5437), .Z(n5499) );
  AND U6407 ( .A(a[63]), .B(b[3]), .Z(n5501) );
  XNOR U6408 ( .A(n5503), .B(n5500), .Z(n5502) );
  XOR U6409 ( .A(n5504), .B(n5505), .Z(n5500) );
  ANDN U6410 ( .B(n5433), .A(n5434), .Z(n5504) );
  AND U6411 ( .A(b[2]), .B(a[63]), .Z(n5506) );
  XNOR U6412 ( .A(n5508), .B(n5505), .Z(n5507) );
  XOR U6413 ( .A(n5509), .B(n5510), .Z(n5505) );
  NANDN U6414 ( .A(n5436), .B(n5435), .Z(n5510) );
  XOR U6415 ( .A(n5509), .B(n5511), .Z(n5435) );
  NAND U6416 ( .A(a[63]), .B(b[1]), .Z(n5511) );
  XOR U6417 ( .A(n5509), .B(n5513), .Z(n5512) );
  OR U6418 ( .A(n2582), .B(n2580), .Z(n5509) );
  XOR U6419 ( .A(n5515), .B(n5516), .Z(n2580) );
  NANDN U6420 ( .A(n179), .B(a[63]), .Z(n2582) );
  XNOR U6421 ( .A(n5487), .B(n5491), .Z(n5519) );
  XNOR U6422 ( .A(n5482), .B(n5486), .Z(n5520) );
  XNOR U6423 ( .A(n5477), .B(n5481), .Z(n5521) );
  XNOR U6424 ( .A(n5472), .B(n5476), .Z(n5522) );
  XNOR U6425 ( .A(n5467), .B(n5471), .Z(n5523) );
  XNOR U6426 ( .A(n5462), .B(n5466), .Z(n5524) );
  XOR U6427 ( .A(n5458), .B(n5461), .Z(n5525) );
  XOR U6428 ( .A(n5526), .B(n5527), .Z(n5458) );
  XNOR U6429 ( .A(n5528), .B(n5529), .Z(n5527) );
  XOR U6430 ( .A(n5530), .B(n5531), .Z(n5528) );
  AND U6431 ( .A(b[13]), .B(a[54]), .Z(n5530) );
  XOR U6432 ( .A(n5531), .B(n5532), .Z(n5526) );
  XOR U6433 ( .A(n5533), .B(n5534), .Z(n5532) );
  AND U6434 ( .A(a[53]), .B(b[14]), .Z(n5534) );
  AND U6435 ( .A(a[52]), .B(b[15]), .Z(n5533) );
  XOR U6436 ( .A(n5535), .B(n5536), .Z(n5531) );
  ANDN U6437 ( .B(n5537), .A(n5538), .Z(n5535) );
  XOR U6438 ( .A(n5539), .B(n5456), .Z(n5457) );
  IV U6439 ( .A(n5529), .Z(n5456) );
  XOR U6440 ( .A(n5540), .B(n5541), .Z(n5529) );
  NOR U6441 ( .A(n5542), .B(n5543), .Z(n5540) );
  AND U6442 ( .A(a[55]), .B(b[12]), .Z(n5539) );
  XOR U6443 ( .A(n5545), .B(n5546), .Z(n5461) );
  ANDN U6444 ( .B(n5547), .A(n5548), .Z(n5545) );
  AND U6445 ( .A(a[56]), .B(b[11]), .Z(n5544) );
  XOR U6446 ( .A(n5550), .B(n5551), .Z(n5466) );
  ANDN U6447 ( .B(n5552), .A(n5553), .Z(n5550) );
  AND U6448 ( .A(a[57]), .B(b[10]), .Z(n5549) );
  XOR U6449 ( .A(n5555), .B(n5556), .Z(n5471) );
  ANDN U6450 ( .B(n5557), .A(n5558), .Z(n5555) );
  AND U6451 ( .A(a[58]), .B(b[9]), .Z(n5554) );
  XOR U6452 ( .A(n5560), .B(n5561), .Z(n5476) );
  ANDN U6453 ( .B(n5562), .A(n5563), .Z(n5560) );
  AND U6454 ( .A(a[59]), .B(b[8]), .Z(n5559) );
  XOR U6455 ( .A(n5565), .B(n5566), .Z(n5481) );
  ANDN U6456 ( .B(n5567), .A(n5568), .Z(n5565) );
  AND U6457 ( .A(a[60]), .B(b[7]), .Z(n5564) );
  XOR U6458 ( .A(n5570), .B(n5571), .Z(n5486) );
  ANDN U6459 ( .B(n5572), .A(n5573), .Z(n5570) );
  AND U6460 ( .A(a[61]), .B(b[6]), .Z(n5569) );
  XOR U6461 ( .A(n5575), .B(n5576), .Z(n5491) );
  ANDN U6462 ( .B(n5503), .A(n5518), .Z(n5575) );
  AND U6463 ( .A(a[62]), .B(b[4]), .Z(n5577) );
  XNOR U6464 ( .A(n5572), .B(n5576), .Z(n5578) );
  XOR U6465 ( .A(n5579), .B(n5580), .Z(n5576) );
  ANDN U6466 ( .B(n5508), .A(n5517), .Z(n5579) );
  AND U6467 ( .A(a[62]), .B(b[3]), .Z(n5581) );
  XNOR U6468 ( .A(n5583), .B(n5580), .Z(n5582) );
  XOR U6469 ( .A(n5584), .B(n5585), .Z(n5580) );
  ANDN U6470 ( .B(n5513), .A(n5514), .Z(n5584) );
  AND U6471 ( .A(b[2]), .B(a[62]), .Z(n5586) );
  XNOR U6472 ( .A(n5588), .B(n5585), .Z(n5587) );
  XOR U6473 ( .A(n5589), .B(n5590), .Z(n5585) );
  NANDN U6474 ( .A(n5516), .B(n5515), .Z(n5590) );
  XOR U6475 ( .A(n5589), .B(n5591), .Z(n5515) );
  NAND U6476 ( .A(a[62]), .B(b[1]), .Z(n5591) );
  XOR U6477 ( .A(n5589), .B(n5593), .Z(n5592) );
  OR U6478 ( .A(n2587), .B(n2585), .Z(n5589) );
  XOR U6479 ( .A(n5595), .B(n5596), .Z(n2585) );
  NANDN U6480 ( .A(n179), .B(a[62]), .Z(n2587) );
  XNOR U6481 ( .A(n5567), .B(n5571), .Z(n5599) );
  XNOR U6482 ( .A(n5562), .B(n5566), .Z(n5600) );
  XNOR U6483 ( .A(n5557), .B(n5561), .Z(n5601) );
  XNOR U6484 ( .A(n5552), .B(n5556), .Z(n5602) );
  XNOR U6485 ( .A(n5547), .B(n5551), .Z(n5603) );
  XOR U6486 ( .A(n5543), .B(n5546), .Z(n5604) );
  XNOR U6487 ( .A(n5538), .B(n5605), .Z(n5543) );
  XNOR U6488 ( .A(n5537), .B(n5541), .Z(n5605) );
  XOR U6489 ( .A(n5606), .B(n5536), .Z(n5537) );
  AND U6490 ( .A(b[12]), .B(a[54]), .Z(n5606) );
  XOR U6491 ( .A(n5607), .B(n5608), .Z(n5538) );
  XOR U6492 ( .A(n5536), .B(n5609), .Z(n5608) );
  XOR U6493 ( .A(n5610), .B(n5611), .Z(n5609) );
  XOR U6494 ( .A(n5612), .B(n5613), .Z(n5611) );
  NAND U6495 ( .A(a[52]), .B(b[14]), .Z(n5613) );
  AND U6496 ( .A(a[51]), .B(b[15]), .Z(n5612) );
  XOR U6497 ( .A(n5614), .B(n5615), .Z(n5536) );
  ANDN U6498 ( .B(n5616), .A(n5617), .Z(n5614) );
  XOR U6499 ( .A(n5618), .B(n5610), .Z(n5607) );
  XOR U6500 ( .A(n5619), .B(n5620), .Z(n5610) );
  NOR U6501 ( .A(n5621), .B(n5622), .Z(n5619) );
  AND U6502 ( .A(a[53]), .B(b[13]), .Z(n5618) );
  XOR U6503 ( .A(n5624), .B(n5625), .Z(n5541) );
  ANDN U6504 ( .B(n5626), .A(n5627), .Z(n5624) );
  AND U6505 ( .A(a[55]), .B(b[11]), .Z(n5623) );
  XOR U6506 ( .A(n5629), .B(n5630), .Z(n5546) );
  ANDN U6507 ( .B(n5631), .A(n5632), .Z(n5629) );
  AND U6508 ( .A(a[56]), .B(b[10]), .Z(n5628) );
  XOR U6509 ( .A(n5634), .B(n5635), .Z(n5551) );
  ANDN U6510 ( .B(n5636), .A(n5637), .Z(n5634) );
  AND U6511 ( .A(a[57]), .B(b[9]), .Z(n5633) );
  XOR U6512 ( .A(n5639), .B(n5640), .Z(n5556) );
  ANDN U6513 ( .B(n5641), .A(n5642), .Z(n5639) );
  AND U6514 ( .A(a[58]), .B(b[8]), .Z(n5638) );
  XOR U6515 ( .A(n5644), .B(n5645), .Z(n5561) );
  ANDN U6516 ( .B(n5646), .A(n5647), .Z(n5644) );
  AND U6517 ( .A(a[59]), .B(b[7]), .Z(n5643) );
  XOR U6518 ( .A(n5649), .B(n5650), .Z(n5566) );
  ANDN U6519 ( .B(n5651), .A(n5652), .Z(n5649) );
  AND U6520 ( .A(a[60]), .B(b[6]), .Z(n5648) );
  XOR U6521 ( .A(n5654), .B(n5655), .Z(n5571) );
  ANDN U6522 ( .B(n5583), .A(n5598), .Z(n5654) );
  AND U6523 ( .A(a[61]), .B(b[4]), .Z(n5656) );
  XNOR U6524 ( .A(n5651), .B(n5655), .Z(n5657) );
  XOR U6525 ( .A(n5658), .B(n5659), .Z(n5655) );
  ANDN U6526 ( .B(n5588), .A(n5597), .Z(n5658) );
  AND U6527 ( .A(a[61]), .B(b[3]), .Z(n5660) );
  XNOR U6528 ( .A(n5662), .B(n5659), .Z(n5661) );
  XOR U6529 ( .A(n5663), .B(n5664), .Z(n5659) );
  ANDN U6530 ( .B(n5593), .A(n5594), .Z(n5663) );
  AND U6531 ( .A(b[2]), .B(a[61]), .Z(n5665) );
  XNOR U6532 ( .A(n5667), .B(n5664), .Z(n5666) );
  XOR U6533 ( .A(n5668), .B(n5669), .Z(n5664) );
  NANDN U6534 ( .A(n5596), .B(n5595), .Z(n5669) );
  XOR U6535 ( .A(n5668), .B(n5670), .Z(n5595) );
  NAND U6536 ( .A(a[61]), .B(b[1]), .Z(n5670) );
  XOR U6537 ( .A(n5668), .B(n5672), .Z(n5671) );
  OR U6538 ( .A(n2592), .B(n2590), .Z(n5668) );
  XOR U6539 ( .A(n5674), .B(n5675), .Z(n2590) );
  NANDN U6540 ( .A(n179), .B(a[61]), .Z(n2592) );
  XNOR U6541 ( .A(n5646), .B(n5650), .Z(n5678) );
  XNOR U6542 ( .A(n5641), .B(n5645), .Z(n5679) );
  XNOR U6543 ( .A(n5636), .B(n5640), .Z(n5680) );
  XNOR U6544 ( .A(n5631), .B(n5635), .Z(n5681) );
  XNOR U6545 ( .A(n5626), .B(n5630), .Z(n5682) );
  XNOR U6546 ( .A(n5616), .B(n5625), .Z(n5683) );
  XOR U6547 ( .A(n5684), .B(n5615), .Z(n5616) );
  AND U6548 ( .A(b[11]), .B(a[54]), .Z(n5684) );
  XOR U6549 ( .A(n5615), .B(n5622), .Z(n5685) );
  XOR U6550 ( .A(n5686), .B(n5687), .Z(n5622) );
  XOR U6551 ( .A(n5620), .B(n5688), .Z(n5687) );
  XOR U6552 ( .A(n5689), .B(n5690), .Z(n5688) );
  XOR U6553 ( .A(n5691), .B(n5692), .Z(n5690) );
  NAND U6554 ( .A(a[51]), .B(b[14]), .Z(n5692) );
  AND U6555 ( .A(a[50]), .B(b[15]), .Z(n5691) );
  XOR U6556 ( .A(n5693), .B(n5689), .Z(n5686) );
  XOR U6557 ( .A(n5694), .B(n5695), .Z(n5689) );
  NOR U6558 ( .A(n5696), .B(n5697), .Z(n5694) );
  AND U6559 ( .A(a[52]), .B(b[13]), .Z(n5693) );
  XOR U6560 ( .A(n5698), .B(n5699), .Z(n5615) );
  ANDN U6561 ( .B(n5700), .A(n5701), .Z(n5698) );
  XNOR U6562 ( .A(n5702), .B(n5620), .Z(n5621) );
  XOR U6563 ( .A(n5703), .B(n5704), .Z(n5620) );
  ANDN U6564 ( .B(n5705), .A(n5706), .Z(n5703) );
  AND U6565 ( .A(a[53]), .B(b[12]), .Z(n5702) );
  XOR U6566 ( .A(n5708), .B(n5709), .Z(n5625) );
  ANDN U6567 ( .B(n5710), .A(n5711), .Z(n5708) );
  AND U6568 ( .A(a[55]), .B(b[10]), .Z(n5707) );
  XOR U6569 ( .A(n5713), .B(n5714), .Z(n5630) );
  ANDN U6570 ( .B(n5715), .A(n5716), .Z(n5713) );
  AND U6571 ( .A(a[56]), .B(b[9]), .Z(n5712) );
  XOR U6572 ( .A(n5718), .B(n5719), .Z(n5635) );
  ANDN U6573 ( .B(n5720), .A(n5721), .Z(n5718) );
  AND U6574 ( .A(a[57]), .B(b[8]), .Z(n5717) );
  XOR U6575 ( .A(n5723), .B(n5724), .Z(n5640) );
  ANDN U6576 ( .B(n5725), .A(n5726), .Z(n5723) );
  AND U6577 ( .A(a[58]), .B(b[7]), .Z(n5722) );
  XOR U6578 ( .A(n5728), .B(n5729), .Z(n5645) );
  ANDN U6579 ( .B(n5730), .A(n5731), .Z(n5728) );
  AND U6580 ( .A(a[59]), .B(b[6]), .Z(n5727) );
  XOR U6581 ( .A(n5733), .B(n5734), .Z(n5650) );
  ANDN U6582 ( .B(n5662), .A(n5677), .Z(n5733) );
  AND U6583 ( .A(a[60]), .B(b[4]), .Z(n5735) );
  XNOR U6584 ( .A(n5730), .B(n5734), .Z(n5736) );
  XOR U6585 ( .A(n5737), .B(n5738), .Z(n5734) );
  ANDN U6586 ( .B(n5667), .A(n5676), .Z(n5737) );
  AND U6587 ( .A(a[60]), .B(b[3]), .Z(n5739) );
  XNOR U6588 ( .A(n5741), .B(n5738), .Z(n5740) );
  XOR U6589 ( .A(n5742), .B(n5743), .Z(n5738) );
  ANDN U6590 ( .B(n5672), .A(n5673), .Z(n5742) );
  AND U6591 ( .A(b[2]), .B(a[60]), .Z(n5744) );
  XNOR U6592 ( .A(n5746), .B(n5743), .Z(n5745) );
  XOR U6593 ( .A(n5747), .B(n5748), .Z(n5743) );
  NANDN U6594 ( .A(n5675), .B(n5674), .Z(n5748) );
  XOR U6595 ( .A(n5747), .B(n5749), .Z(n5674) );
  NAND U6596 ( .A(a[60]), .B(b[1]), .Z(n5749) );
  XOR U6597 ( .A(n5747), .B(n5751), .Z(n5750) );
  OR U6598 ( .A(n2597), .B(n2595), .Z(n5747) );
  XOR U6599 ( .A(n5753), .B(n5754), .Z(n2595) );
  NANDN U6600 ( .A(n179), .B(a[60]), .Z(n2597) );
  XNOR U6601 ( .A(n5725), .B(n5729), .Z(n5757) );
  XNOR U6602 ( .A(n5720), .B(n5724), .Z(n5758) );
  XNOR U6603 ( .A(n5715), .B(n5719), .Z(n5759) );
  XNOR U6604 ( .A(n5710), .B(n5714), .Z(n5760) );
  XNOR U6605 ( .A(n5700), .B(n5709), .Z(n5761) );
  XOR U6606 ( .A(n5762), .B(n5699), .Z(n5700) );
  AND U6607 ( .A(b[10]), .B(a[54]), .Z(n5762) );
  XNOR U6608 ( .A(n5699), .B(n5705), .Z(n5763) );
  XOR U6609 ( .A(n5704), .B(n5697), .Z(n5764) );
  XOR U6610 ( .A(n5765), .B(n5766), .Z(n5697) );
  XOR U6611 ( .A(n5695), .B(n5767), .Z(n5766) );
  XOR U6612 ( .A(n5768), .B(n5769), .Z(n5767) );
  XOR U6613 ( .A(n5770), .B(n5771), .Z(n5769) );
  NAND U6614 ( .A(a[50]), .B(b[14]), .Z(n5771) );
  AND U6615 ( .A(a[49]), .B(b[15]), .Z(n5770) );
  XOR U6616 ( .A(n5772), .B(n5768), .Z(n5765) );
  XOR U6617 ( .A(n5773), .B(n5774), .Z(n5768) );
  NOR U6618 ( .A(n5775), .B(n5776), .Z(n5773) );
  AND U6619 ( .A(a[51]), .B(b[13]), .Z(n5772) );
  XNOR U6620 ( .A(n5777), .B(n5695), .Z(n5696) );
  XOR U6621 ( .A(n5778), .B(n5779), .Z(n5695) );
  ANDN U6622 ( .B(n5780), .A(n5781), .Z(n5778) );
  AND U6623 ( .A(a[52]), .B(b[12]), .Z(n5777) );
  XOR U6624 ( .A(n5782), .B(n5783), .Z(n5699) );
  ANDN U6625 ( .B(n5784), .A(n5785), .Z(n5782) );
  XNOR U6626 ( .A(n5786), .B(n5704), .Z(n5706) );
  XOR U6627 ( .A(n5787), .B(n5788), .Z(n5704) );
  ANDN U6628 ( .B(n5789), .A(n5790), .Z(n5787) );
  AND U6629 ( .A(a[53]), .B(b[11]), .Z(n5786) );
  XOR U6630 ( .A(n5792), .B(n5793), .Z(n5709) );
  ANDN U6631 ( .B(n5794), .A(n5795), .Z(n5792) );
  AND U6632 ( .A(a[55]), .B(b[9]), .Z(n5791) );
  XOR U6633 ( .A(n5797), .B(n5798), .Z(n5714) );
  ANDN U6634 ( .B(n5799), .A(n5800), .Z(n5797) );
  AND U6635 ( .A(a[56]), .B(b[8]), .Z(n5796) );
  XOR U6636 ( .A(n5802), .B(n5803), .Z(n5719) );
  ANDN U6637 ( .B(n5804), .A(n5805), .Z(n5802) );
  AND U6638 ( .A(a[57]), .B(b[7]), .Z(n5801) );
  XOR U6639 ( .A(n5807), .B(n5808), .Z(n5724) );
  ANDN U6640 ( .B(n5809), .A(n5810), .Z(n5807) );
  AND U6641 ( .A(a[58]), .B(b[6]), .Z(n5806) );
  XOR U6642 ( .A(n5812), .B(n5813), .Z(n5729) );
  ANDN U6643 ( .B(n5741), .A(n5756), .Z(n5812) );
  AND U6644 ( .A(a[59]), .B(b[4]), .Z(n5814) );
  XNOR U6645 ( .A(n5809), .B(n5813), .Z(n5815) );
  XOR U6646 ( .A(n5816), .B(n5817), .Z(n5813) );
  ANDN U6647 ( .B(n5746), .A(n5755), .Z(n5816) );
  AND U6648 ( .A(a[59]), .B(b[3]), .Z(n5818) );
  XNOR U6649 ( .A(n5820), .B(n5817), .Z(n5819) );
  XOR U6650 ( .A(n5821), .B(n5822), .Z(n5817) );
  ANDN U6651 ( .B(n5751), .A(n5752), .Z(n5821) );
  AND U6652 ( .A(b[2]), .B(a[59]), .Z(n5823) );
  XNOR U6653 ( .A(n5825), .B(n5822), .Z(n5824) );
  XOR U6654 ( .A(n5826), .B(n5827), .Z(n5822) );
  NANDN U6655 ( .A(n5754), .B(n5753), .Z(n5827) );
  XOR U6656 ( .A(n5826), .B(n5828), .Z(n5753) );
  NAND U6657 ( .A(a[59]), .B(b[1]), .Z(n5828) );
  XOR U6658 ( .A(n5826), .B(n5830), .Z(n5829) );
  OR U6659 ( .A(n2602), .B(n2600), .Z(n5826) );
  XOR U6660 ( .A(n5832), .B(n5833), .Z(n2600) );
  NANDN U6661 ( .A(n179), .B(a[59]), .Z(n2602) );
  XNOR U6662 ( .A(n5804), .B(n5808), .Z(n5836) );
  XNOR U6663 ( .A(n5799), .B(n5803), .Z(n5837) );
  XNOR U6664 ( .A(n5794), .B(n5798), .Z(n5838) );
  XNOR U6665 ( .A(n5784), .B(n5793), .Z(n5839) );
  XOR U6666 ( .A(n5840), .B(n5783), .Z(n5784) );
  AND U6667 ( .A(b[9]), .B(a[54]), .Z(n5840) );
  XNOR U6668 ( .A(n5783), .B(n5789), .Z(n5841) );
  XNOR U6669 ( .A(n5788), .B(n5780), .Z(n5842) );
  XOR U6670 ( .A(n5779), .B(n5776), .Z(n5843) );
  XOR U6671 ( .A(n5844), .B(n5845), .Z(n5776) );
  XOR U6672 ( .A(n5774), .B(n5846), .Z(n5845) );
  XOR U6673 ( .A(n5847), .B(n5848), .Z(n5846) );
  XOR U6674 ( .A(n5849), .B(n5850), .Z(n5848) );
  NAND U6675 ( .A(a[49]), .B(b[14]), .Z(n5850) );
  AND U6676 ( .A(a[48]), .B(b[15]), .Z(n5849) );
  XOR U6677 ( .A(n5851), .B(n5847), .Z(n5844) );
  XOR U6678 ( .A(n5852), .B(n5853), .Z(n5847) );
  NOR U6679 ( .A(n5854), .B(n5855), .Z(n5852) );
  AND U6680 ( .A(a[50]), .B(b[13]), .Z(n5851) );
  XNOR U6681 ( .A(n5856), .B(n5774), .Z(n5775) );
  XOR U6682 ( .A(n5857), .B(n5858), .Z(n5774) );
  ANDN U6683 ( .B(n5859), .A(n5860), .Z(n5857) );
  AND U6684 ( .A(a[51]), .B(b[12]), .Z(n5856) );
  XNOR U6685 ( .A(n5861), .B(n5779), .Z(n5781) );
  XOR U6686 ( .A(n5862), .B(n5863), .Z(n5779) );
  ANDN U6687 ( .B(n5864), .A(n5865), .Z(n5862) );
  AND U6688 ( .A(a[52]), .B(b[11]), .Z(n5861) );
  XOR U6689 ( .A(n5866), .B(n5867), .Z(n5783) );
  ANDN U6690 ( .B(n5868), .A(n5869), .Z(n5866) );
  XNOR U6691 ( .A(n5870), .B(n5788), .Z(n5790) );
  XOR U6692 ( .A(n5871), .B(n5872), .Z(n5788) );
  ANDN U6693 ( .B(n5873), .A(n5874), .Z(n5871) );
  AND U6694 ( .A(a[53]), .B(b[10]), .Z(n5870) );
  XOR U6695 ( .A(n5876), .B(n5877), .Z(n5793) );
  ANDN U6696 ( .B(n5878), .A(n5879), .Z(n5876) );
  AND U6697 ( .A(a[55]), .B(b[8]), .Z(n5875) );
  XOR U6698 ( .A(n5881), .B(n5882), .Z(n5798) );
  ANDN U6699 ( .B(n5883), .A(n5884), .Z(n5881) );
  AND U6700 ( .A(a[56]), .B(b[7]), .Z(n5880) );
  XOR U6701 ( .A(n5886), .B(n5887), .Z(n5803) );
  ANDN U6702 ( .B(n5888), .A(n5889), .Z(n5886) );
  AND U6703 ( .A(a[57]), .B(b[6]), .Z(n5885) );
  XOR U6704 ( .A(n5891), .B(n5892), .Z(n5808) );
  ANDN U6705 ( .B(n5820), .A(n5835), .Z(n5891) );
  AND U6706 ( .A(a[58]), .B(b[4]), .Z(n5893) );
  XNOR U6707 ( .A(n5888), .B(n5892), .Z(n5894) );
  XOR U6708 ( .A(n5895), .B(n5896), .Z(n5892) );
  ANDN U6709 ( .B(n5825), .A(n5834), .Z(n5895) );
  AND U6710 ( .A(a[58]), .B(b[3]), .Z(n5897) );
  XNOR U6711 ( .A(n5899), .B(n5896), .Z(n5898) );
  XOR U6712 ( .A(n5900), .B(n5901), .Z(n5896) );
  ANDN U6713 ( .B(n5830), .A(n5831), .Z(n5900) );
  AND U6714 ( .A(b[2]), .B(a[58]), .Z(n5902) );
  XNOR U6715 ( .A(n5904), .B(n5901), .Z(n5903) );
  XOR U6716 ( .A(n5905), .B(n5906), .Z(n5901) );
  NANDN U6717 ( .A(n5833), .B(n5832), .Z(n5906) );
  XOR U6718 ( .A(n5905), .B(n5907), .Z(n5832) );
  NAND U6719 ( .A(a[58]), .B(b[1]), .Z(n5907) );
  XOR U6720 ( .A(n5905), .B(n5909), .Z(n5908) );
  OR U6721 ( .A(n2607), .B(n2605), .Z(n5905) );
  XOR U6722 ( .A(n5911), .B(n5912), .Z(n2605) );
  NANDN U6723 ( .A(n179), .B(a[58]), .Z(n2607) );
  XNOR U6724 ( .A(n5883), .B(n5887), .Z(n5915) );
  XNOR U6725 ( .A(n5878), .B(n5882), .Z(n5916) );
  XNOR U6726 ( .A(n5868), .B(n5877), .Z(n5917) );
  XOR U6727 ( .A(n5918), .B(n5867), .Z(n5868) );
  AND U6728 ( .A(b[8]), .B(a[54]), .Z(n5918) );
  XNOR U6729 ( .A(n5867), .B(n5873), .Z(n5919) );
  XNOR U6730 ( .A(n5872), .B(n5864), .Z(n5920) );
  XNOR U6731 ( .A(n5863), .B(n5859), .Z(n5921) );
  XOR U6732 ( .A(n5858), .B(n5855), .Z(n5922) );
  XOR U6733 ( .A(n5923), .B(n5924), .Z(n5855) );
  XOR U6734 ( .A(n5853), .B(n5925), .Z(n5924) );
  XOR U6735 ( .A(n5926), .B(n5927), .Z(n5925) );
  XOR U6736 ( .A(n5928), .B(n5929), .Z(n5927) );
  NAND U6737 ( .A(a[48]), .B(b[14]), .Z(n5929) );
  AND U6738 ( .A(a[47]), .B(b[15]), .Z(n5928) );
  XOR U6739 ( .A(n5930), .B(n5926), .Z(n5923) );
  XOR U6740 ( .A(n5931), .B(n5932), .Z(n5926) );
  NOR U6741 ( .A(n5933), .B(n5934), .Z(n5931) );
  AND U6742 ( .A(a[49]), .B(b[13]), .Z(n5930) );
  XNOR U6743 ( .A(n5935), .B(n5853), .Z(n5854) );
  XOR U6744 ( .A(n5936), .B(n5937), .Z(n5853) );
  ANDN U6745 ( .B(n5938), .A(n5939), .Z(n5936) );
  AND U6746 ( .A(a[50]), .B(b[12]), .Z(n5935) );
  XNOR U6747 ( .A(n5940), .B(n5858), .Z(n5860) );
  XOR U6748 ( .A(n5941), .B(n5942), .Z(n5858) );
  ANDN U6749 ( .B(n5943), .A(n5944), .Z(n5941) );
  AND U6750 ( .A(a[51]), .B(b[11]), .Z(n5940) );
  XNOR U6751 ( .A(n5945), .B(n5863), .Z(n5865) );
  XOR U6752 ( .A(n5946), .B(n5947), .Z(n5863) );
  ANDN U6753 ( .B(n5948), .A(n5949), .Z(n5946) );
  AND U6754 ( .A(a[52]), .B(b[10]), .Z(n5945) );
  XOR U6755 ( .A(n5950), .B(n5951), .Z(n5867) );
  ANDN U6756 ( .B(n5952), .A(n5953), .Z(n5950) );
  XNOR U6757 ( .A(n5954), .B(n5872), .Z(n5874) );
  XOR U6758 ( .A(n5955), .B(n5956), .Z(n5872) );
  ANDN U6759 ( .B(n5957), .A(n5958), .Z(n5955) );
  AND U6760 ( .A(a[53]), .B(b[9]), .Z(n5954) );
  XOR U6761 ( .A(n5960), .B(n5961), .Z(n5877) );
  ANDN U6762 ( .B(n5962), .A(n5963), .Z(n5960) );
  AND U6763 ( .A(a[55]), .B(b[7]), .Z(n5959) );
  XOR U6764 ( .A(n5965), .B(n5966), .Z(n5882) );
  ANDN U6765 ( .B(n5967), .A(n5968), .Z(n5965) );
  AND U6766 ( .A(a[56]), .B(b[6]), .Z(n5964) );
  XOR U6767 ( .A(n5970), .B(n5971), .Z(n5887) );
  ANDN U6768 ( .B(n5899), .A(n5914), .Z(n5970) );
  AND U6769 ( .A(a[57]), .B(b[4]), .Z(n5972) );
  XNOR U6770 ( .A(n5967), .B(n5971), .Z(n5973) );
  XOR U6771 ( .A(n5974), .B(n5975), .Z(n5971) );
  ANDN U6772 ( .B(n5904), .A(n5913), .Z(n5974) );
  AND U6773 ( .A(a[57]), .B(b[3]), .Z(n5976) );
  XNOR U6774 ( .A(n5978), .B(n5975), .Z(n5977) );
  XOR U6775 ( .A(n5979), .B(n5980), .Z(n5975) );
  ANDN U6776 ( .B(n5909), .A(n5910), .Z(n5979) );
  AND U6777 ( .A(b[2]), .B(a[57]), .Z(n5981) );
  XNOR U6778 ( .A(n5983), .B(n5980), .Z(n5982) );
  XOR U6779 ( .A(n5984), .B(n5985), .Z(n5980) );
  NANDN U6780 ( .A(n5912), .B(n5911), .Z(n5985) );
  XOR U6781 ( .A(n5984), .B(n5986), .Z(n5911) );
  NAND U6782 ( .A(a[57]), .B(b[1]), .Z(n5986) );
  XOR U6783 ( .A(n5984), .B(n5988), .Z(n5987) );
  OR U6784 ( .A(n2612), .B(n2610), .Z(n5984) );
  XOR U6785 ( .A(n5990), .B(n5991), .Z(n2610) );
  NANDN U6786 ( .A(n179), .B(a[57]), .Z(n2612) );
  XNOR U6787 ( .A(n5962), .B(n5966), .Z(n5994) );
  XNOR U6788 ( .A(n5952), .B(n5961), .Z(n5995) );
  XOR U6789 ( .A(n5996), .B(n5951), .Z(n5952) );
  AND U6790 ( .A(b[7]), .B(a[54]), .Z(n5996) );
  XNOR U6791 ( .A(n5951), .B(n5957), .Z(n5997) );
  XNOR U6792 ( .A(n5956), .B(n5948), .Z(n5998) );
  XNOR U6793 ( .A(n5947), .B(n5943), .Z(n5999) );
  XNOR U6794 ( .A(n5942), .B(n5938), .Z(n6000) );
  XOR U6795 ( .A(n5937), .B(n5934), .Z(n6001) );
  XOR U6796 ( .A(n6002), .B(n6003), .Z(n5934) );
  XOR U6797 ( .A(n5932), .B(n6004), .Z(n6003) );
  XOR U6798 ( .A(n6005), .B(n6006), .Z(n6004) );
  XOR U6799 ( .A(n6007), .B(n6008), .Z(n6006) );
  NAND U6800 ( .A(a[47]), .B(b[14]), .Z(n6008) );
  AND U6801 ( .A(a[46]), .B(b[15]), .Z(n6007) );
  XOR U6802 ( .A(n6009), .B(n6005), .Z(n6002) );
  XOR U6803 ( .A(n6010), .B(n6011), .Z(n6005) );
  NOR U6804 ( .A(n6012), .B(n6013), .Z(n6010) );
  AND U6805 ( .A(a[48]), .B(b[13]), .Z(n6009) );
  XNOR U6806 ( .A(n6014), .B(n5932), .Z(n5933) );
  XOR U6807 ( .A(n6015), .B(n6016), .Z(n5932) );
  ANDN U6808 ( .B(n6017), .A(n6018), .Z(n6015) );
  AND U6809 ( .A(a[49]), .B(b[12]), .Z(n6014) );
  XNOR U6810 ( .A(n6019), .B(n5937), .Z(n5939) );
  XOR U6811 ( .A(n6020), .B(n6021), .Z(n5937) );
  ANDN U6812 ( .B(n6022), .A(n6023), .Z(n6020) );
  AND U6813 ( .A(a[50]), .B(b[11]), .Z(n6019) );
  XNOR U6814 ( .A(n6024), .B(n5942), .Z(n5944) );
  XOR U6815 ( .A(n6025), .B(n6026), .Z(n5942) );
  ANDN U6816 ( .B(n6027), .A(n6028), .Z(n6025) );
  AND U6817 ( .A(a[51]), .B(b[10]), .Z(n6024) );
  XNOR U6818 ( .A(n6029), .B(n5947), .Z(n5949) );
  XOR U6819 ( .A(n6030), .B(n6031), .Z(n5947) );
  ANDN U6820 ( .B(n6032), .A(n6033), .Z(n6030) );
  AND U6821 ( .A(a[52]), .B(b[9]), .Z(n6029) );
  XOR U6822 ( .A(n6034), .B(n6035), .Z(n5951) );
  ANDN U6823 ( .B(n6036), .A(n6037), .Z(n6034) );
  XNOR U6824 ( .A(n6038), .B(n5956), .Z(n5958) );
  XOR U6825 ( .A(n6039), .B(n6040), .Z(n5956) );
  ANDN U6826 ( .B(n6041), .A(n6042), .Z(n6039) );
  AND U6827 ( .A(a[53]), .B(b[8]), .Z(n6038) );
  XOR U6828 ( .A(n6044), .B(n6045), .Z(n5961) );
  ANDN U6829 ( .B(n6046), .A(n6047), .Z(n6044) );
  AND U6830 ( .A(a[55]), .B(b[6]), .Z(n6043) );
  XOR U6831 ( .A(n6049), .B(n6050), .Z(n5966) );
  ANDN U6832 ( .B(n5978), .A(n5993), .Z(n6049) );
  AND U6833 ( .A(a[56]), .B(b[4]), .Z(n6051) );
  XNOR U6834 ( .A(n6046), .B(n6050), .Z(n6052) );
  XOR U6835 ( .A(n6053), .B(n6054), .Z(n6050) );
  ANDN U6836 ( .B(n5983), .A(n5992), .Z(n6053) );
  AND U6837 ( .A(a[56]), .B(b[3]), .Z(n6055) );
  XNOR U6838 ( .A(n6057), .B(n6054), .Z(n6056) );
  XOR U6839 ( .A(n6058), .B(n6059), .Z(n6054) );
  ANDN U6840 ( .B(n5988), .A(n5989), .Z(n6058) );
  AND U6841 ( .A(b[2]), .B(a[56]), .Z(n6060) );
  XNOR U6842 ( .A(n6062), .B(n6059), .Z(n6061) );
  XOR U6843 ( .A(n6063), .B(n6064), .Z(n6059) );
  NANDN U6844 ( .A(n5991), .B(n5990), .Z(n6064) );
  XOR U6845 ( .A(n6063), .B(n6065), .Z(n5990) );
  NAND U6846 ( .A(a[56]), .B(b[1]), .Z(n6065) );
  XOR U6847 ( .A(n6063), .B(n6067), .Z(n6066) );
  OR U6848 ( .A(n2617), .B(n2615), .Z(n6063) );
  XOR U6849 ( .A(n6069), .B(n6070), .Z(n2615) );
  NANDN U6850 ( .A(n179), .B(a[56]), .Z(n2617) );
  XNOR U6851 ( .A(n6036), .B(n6045), .Z(n6073) );
  XOR U6852 ( .A(n6074), .B(n6035), .Z(n6036) );
  AND U6853 ( .A(b[6]), .B(a[54]), .Z(n6074) );
  XNOR U6854 ( .A(n6035), .B(n6041), .Z(n6075) );
  XNOR U6855 ( .A(n6040), .B(n6032), .Z(n6076) );
  XNOR U6856 ( .A(n6031), .B(n6027), .Z(n6077) );
  XNOR U6857 ( .A(n6026), .B(n6022), .Z(n6078) );
  XNOR U6858 ( .A(n6021), .B(n6017), .Z(n6079) );
  XOR U6859 ( .A(n6016), .B(n6013), .Z(n6080) );
  XOR U6860 ( .A(n6081), .B(n6082), .Z(n6013) );
  XOR U6861 ( .A(n6011), .B(n6083), .Z(n6082) );
  XOR U6862 ( .A(n6084), .B(n6085), .Z(n6083) );
  XOR U6863 ( .A(n6086), .B(n6087), .Z(n6085) );
  NAND U6864 ( .A(a[46]), .B(b[14]), .Z(n6087) );
  AND U6865 ( .A(a[45]), .B(b[15]), .Z(n6086) );
  XOR U6866 ( .A(n6088), .B(n6084), .Z(n6081) );
  XOR U6867 ( .A(n6089), .B(n6090), .Z(n6084) );
  NOR U6868 ( .A(n6091), .B(n6092), .Z(n6089) );
  AND U6869 ( .A(a[47]), .B(b[13]), .Z(n6088) );
  XNOR U6870 ( .A(n6093), .B(n6011), .Z(n6012) );
  XOR U6871 ( .A(n6094), .B(n6095), .Z(n6011) );
  ANDN U6872 ( .B(n6096), .A(n6097), .Z(n6094) );
  AND U6873 ( .A(a[48]), .B(b[12]), .Z(n6093) );
  XNOR U6874 ( .A(n6098), .B(n6016), .Z(n6018) );
  XOR U6875 ( .A(n6099), .B(n6100), .Z(n6016) );
  ANDN U6876 ( .B(n6101), .A(n6102), .Z(n6099) );
  AND U6877 ( .A(a[49]), .B(b[11]), .Z(n6098) );
  XNOR U6878 ( .A(n6103), .B(n6021), .Z(n6023) );
  XOR U6879 ( .A(n6104), .B(n6105), .Z(n6021) );
  ANDN U6880 ( .B(n6106), .A(n6107), .Z(n6104) );
  AND U6881 ( .A(a[50]), .B(b[10]), .Z(n6103) );
  XNOR U6882 ( .A(n6108), .B(n6026), .Z(n6028) );
  XOR U6883 ( .A(n6109), .B(n6110), .Z(n6026) );
  ANDN U6884 ( .B(n6111), .A(n6112), .Z(n6109) );
  AND U6885 ( .A(a[51]), .B(b[9]), .Z(n6108) );
  XNOR U6886 ( .A(n6113), .B(n6031), .Z(n6033) );
  XOR U6887 ( .A(n6114), .B(n6115), .Z(n6031) );
  ANDN U6888 ( .B(n6116), .A(n6117), .Z(n6114) );
  AND U6889 ( .A(a[52]), .B(b[8]), .Z(n6113) );
  XOR U6890 ( .A(n6118), .B(n6119), .Z(n6035) );
  ANDN U6891 ( .B(n6120), .A(n6121), .Z(n6118) );
  XNOR U6892 ( .A(n6122), .B(n6040), .Z(n6042) );
  XOR U6893 ( .A(n6123), .B(n6124), .Z(n6040) );
  ANDN U6894 ( .B(n6125), .A(n6126), .Z(n6123) );
  AND U6895 ( .A(a[53]), .B(b[7]), .Z(n6122) );
  XOR U6896 ( .A(n6128), .B(n6129), .Z(n6045) );
  ANDN U6897 ( .B(n6057), .A(n6072), .Z(n6128) );
  AND U6898 ( .A(a[55]), .B(b[4]), .Z(n6130) );
  XNOR U6899 ( .A(n6120), .B(n6129), .Z(n6131) );
  XOR U6900 ( .A(n6132), .B(n6133), .Z(n6129) );
  ANDN U6901 ( .B(n6062), .A(n6071), .Z(n6132) );
  AND U6902 ( .A(a[55]), .B(b[3]), .Z(n6134) );
  XNOR U6903 ( .A(n6136), .B(n6133), .Z(n6135) );
  XOR U6904 ( .A(n6137), .B(n6138), .Z(n6133) );
  ANDN U6905 ( .B(n6067), .A(n6068), .Z(n6137) );
  AND U6906 ( .A(b[2]), .B(a[55]), .Z(n6139) );
  XNOR U6907 ( .A(n6141), .B(n6138), .Z(n6140) );
  XOR U6908 ( .A(n6142), .B(n6143), .Z(n6138) );
  NANDN U6909 ( .A(n6070), .B(n6069), .Z(n6143) );
  XOR U6910 ( .A(n6142), .B(n6144), .Z(n6069) );
  NAND U6911 ( .A(a[55]), .B(b[1]), .Z(n6144) );
  XNOR U6912 ( .A(n6142), .B(n6146), .Z(n6145) );
  OR U6913 ( .A(n2622), .B(n2620), .Z(n6142) );
  NANDN U6914 ( .A(n179), .B(a[55]), .Z(n2622) );
  XOR U6915 ( .A(n6152), .B(n6119), .Z(n6120) );
  AND U6916 ( .A(b[5]), .B(a[54]), .Z(n6152) );
  XNOR U6917 ( .A(n6119), .B(n6125), .Z(n6153) );
  XNOR U6918 ( .A(n6124), .B(n6116), .Z(n6154) );
  XNOR U6919 ( .A(n6115), .B(n6111), .Z(n6155) );
  XNOR U6920 ( .A(n6110), .B(n6106), .Z(n6156) );
  XNOR U6921 ( .A(n6105), .B(n6101), .Z(n6157) );
  XNOR U6922 ( .A(n6100), .B(n6096), .Z(n6158) );
  XOR U6923 ( .A(n6095), .B(n6092), .Z(n6159) );
  XOR U6924 ( .A(n6160), .B(n6161), .Z(n6092) );
  XOR U6925 ( .A(n6090), .B(n6162), .Z(n6161) );
  XOR U6926 ( .A(n6163), .B(n6164), .Z(n6162) );
  XOR U6927 ( .A(n6165), .B(n6166), .Z(n6164) );
  NAND U6928 ( .A(a[45]), .B(b[14]), .Z(n6166) );
  AND U6929 ( .A(a[44]), .B(b[15]), .Z(n6165) );
  XOR U6930 ( .A(n6167), .B(n6163), .Z(n6160) );
  XOR U6931 ( .A(n6168), .B(n6169), .Z(n6163) );
  NOR U6932 ( .A(n6170), .B(n6171), .Z(n6168) );
  AND U6933 ( .A(a[46]), .B(b[13]), .Z(n6167) );
  XNOR U6934 ( .A(n6172), .B(n6090), .Z(n6091) );
  XOR U6935 ( .A(n6173), .B(n6174), .Z(n6090) );
  ANDN U6936 ( .B(n6175), .A(n6176), .Z(n6173) );
  AND U6937 ( .A(a[47]), .B(b[12]), .Z(n6172) );
  XNOR U6938 ( .A(n6177), .B(n6095), .Z(n6097) );
  XOR U6939 ( .A(n6178), .B(n6179), .Z(n6095) );
  ANDN U6940 ( .B(n6180), .A(n6181), .Z(n6178) );
  AND U6941 ( .A(a[48]), .B(b[11]), .Z(n6177) );
  XNOR U6942 ( .A(n6182), .B(n6100), .Z(n6102) );
  XOR U6943 ( .A(n6183), .B(n6184), .Z(n6100) );
  ANDN U6944 ( .B(n6185), .A(n6186), .Z(n6183) );
  AND U6945 ( .A(a[49]), .B(b[10]), .Z(n6182) );
  XNOR U6946 ( .A(n6187), .B(n6105), .Z(n6107) );
  XOR U6947 ( .A(n6188), .B(n6189), .Z(n6105) );
  ANDN U6948 ( .B(n6190), .A(n6191), .Z(n6188) );
  AND U6949 ( .A(a[50]), .B(b[9]), .Z(n6187) );
  XNOR U6950 ( .A(n6192), .B(n6110), .Z(n6112) );
  XOR U6951 ( .A(n6193), .B(n6194), .Z(n6110) );
  ANDN U6952 ( .B(n6195), .A(n6196), .Z(n6193) );
  AND U6953 ( .A(a[51]), .B(b[8]), .Z(n6192) );
  XNOR U6954 ( .A(n6197), .B(n6115), .Z(n6117) );
  XOR U6955 ( .A(n6198), .B(n6199), .Z(n6115) );
  ANDN U6956 ( .B(n6200), .A(n6201), .Z(n6198) );
  AND U6957 ( .A(a[52]), .B(b[7]), .Z(n6197) );
  XOR U6958 ( .A(n6202), .B(n6203), .Z(n6119) );
  ANDN U6959 ( .B(n6136), .A(n6151), .Z(n6202) );
  XNOR U6960 ( .A(n6203), .B(n6205), .Z(n6204) );
  XOR U6961 ( .A(n6207), .B(n6203), .Z(n6136) );
  XOR U6962 ( .A(n6208), .B(n6209), .Z(n6203) );
  ANDN U6963 ( .B(n6141), .A(n6150), .Z(n6208) );
  XNOR U6964 ( .A(n6209), .B(n6211), .Z(n6210) );
  XOR U6965 ( .A(n6213), .B(n6209), .Z(n6141) );
  XNOR U6966 ( .A(n6214), .B(n6215), .Z(n6209) );
  NOR U6967 ( .A(n6147), .B(n6146), .Z(n6214) );
  XOR U6968 ( .A(n6216), .B(n6215), .Z(n6146) );
  AND U6969 ( .A(b[2]), .B(a[54]), .Z(n6216) );
  XOR U6970 ( .A(n6215), .B(n6218), .Z(n6217) );
  XNOR U6971 ( .A(n6219), .B(n6220), .Z(n6215) );
  OR U6972 ( .A(n6148), .B(n6149), .Z(n6220) );
  XNOR U6973 ( .A(n6219), .B(n6222), .Z(n6221) );
  XNOR U6974 ( .A(n6219), .B(n6224), .Z(n6148) );
  NAND U6975 ( .A(b[1]), .B(a[54]), .Z(n6224) );
  OR U6976 ( .A(n2627), .B(n2625), .Z(n6219) );
  XOR U6977 ( .A(n6225), .B(n6226), .Z(n2625) );
  NANDN U6978 ( .A(n179), .B(a[54]), .Z(n2627) );
  AND U6979 ( .A(b[3]), .B(a[54]), .Z(n6213) );
  AND U6980 ( .A(b[4]), .B(a[54]), .Z(n6207) );
  XNOR U6981 ( .A(n6228), .B(n6124), .Z(n6126) );
  XOR U6982 ( .A(n6229), .B(n6230), .Z(n6124) );
  ANDN U6983 ( .B(n6205), .A(n6206), .Z(n6229) );
  XNOR U6984 ( .A(n6231), .B(n6230), .Z(n6206) );
  AND U6985 ( .A(a[53]), .B(b[5]), .Z(n6231) );
  XNOR U6986 ( .A(n6230), .B(n6200), .Z(n6232) );
  XNOR U6987 ( .A(n6199), .B(n6195), .Z(n6233) );
  XNOR U6988 ( .A(n6194), .B(n6190), .Z(n6234) );
  XNOR U6989 ( .A(n6189), .B(n6185), .Z(n6235) );
  XNOR U6990 ( .A(n6184), .B(n6180), .Z(n6236) );
  XNOR U6991 ( .A(n6179), .B(n6175), .Z(n6237) );
  XOR U6992 ( .A(n6174), .B(n6171), .Z(n6238) );
  XOR U6993 ( .A(n6239), .B(n6240), .Z(n6171) );
  XOR U6994 ( .A(n6169), .B(n6241), .Z(n6240) );
  XOR U6995 ( .A(n6242), .B(n6243), .Z(n6241) );
  XOR U6996 ( .A(n6244), .B(n6245), .Z(n6243) );
  NAND U6997 ( .A(a[44]), .B(b[14]), .Z(n6245) );
  AND U6998 ( .A(a[43]), .B(b[15]), .Z(n6244) );
  XOR U6999 ( .A(n6246), .B(n6242), .Z(n6239) );
  XOR U7000 ( .A(n6247), .B(n6248), .Z(n6242) );
  NOR U7001 ( .A(n6249), .B(n6250), .Z(n6247) );
  AND U7002 ( .A(a[45]), .B(b[13]), .Z(n6246) );
  XNOR U7003 ( .A(n6251), .B(n6169), .Z(n6170) );
  XOR U7004 ( .A(n6252), .B(n6253), .Z(n6169) );
  ANDN U7005 ( .B(n6254), .A(n6255), .Z(n6252) );
  AND U7006 ( .A(a[46]), .B(b[12]), .Z(n6251) );
  XNOR U7007 ( .A(n6256), .B(n6174), .Z(n6176) );
  XOR U7008 ( .A(n6257), .B(n6258), .Z(n6174) );
  ANDN U7009 ( .B(n6259), .A(n6260), .Z(n6257) );
  AND U7010 ( .A(a[47]), .B(b[11]), .Z(n6256) );
  XNOR U7011 ( .A(n6261), .B(n6179), .Z(n6181) );
  XOR U7012 ( .A(n6262), .B(n6263), .Z(n6179) );
  ANDN U7013 ( .B(n6264), .A(n6265), .Z(n6262) );
  AND U7014 ( .A(a[48]), .B(b[10]), .Z(n6261) );
  XNOR U7015 ( .A(n6266), .B(n6184), .Z(n6186) );
  XOR U7016 ( .A(n6267), .B(n6268), .Z(n6184) );
  ANDN U7017 ( .B(n6269), .A(n6270), .Z(n6267) );
  AND U7018 ( .A(a[49]), .B(b[9]), .Z(n6266) );
  XNOR U7019 ( .A(n6271), .B(n6189), .Z(n6191) );
  XOR U7020 ( .A(n6272), .B(n6273), .Z(n6189) );
  ANDN U7021 ( .B(n6274), .A(n6275), .Z(n6272) );
  AND U7022 ( .A(a[50]), .B(b[8]), .Z(n6271) );
  XNOR U7023 ( .A(n6276), .B(n6194), .Z(n6196) );
  XOR U7024 ( .A(n6277), .B(n6278), .Z(n6194) );
  ANDN U7025 ( .B(n6279), .A(n6280), .Z(n6277) );
  AND U7026 ( .A(a[51]), .B(b[7]), .Z(n6276) );
  XOR U7027 ( .A(n6281), .B(n6282), .Z(n6230) );
  ANDN U7028 ( .B(n6211), .A(n6212), .Z(n6281) );
  XNOR U7029 ( .A(n6283), .B(n6282), .Z(n6212) );
  AND U7030 ( .A(a[53]), .B(b[4]), .Z(n6283) );
  XNOR U7031 ( .A(n6282), .B(n6285), .Z(n6284) );
  XOR U7032 ( .A(n6286), .B(n6287), .Z(n6282) );
  ANDN U7033 ( .B(n6218), .A(n6227), .Z(n6286) );
  XNOR U7034 ( .A(n6288), .B(n6287), .Z(n6227) );
  AND U7035 ( .A(a[53]), .B(b[3]), .Z(n6288) );
  XNOR U7036 ( .A(n6287), .B(n6290), .Z(n6289) );
  XNOR U7037 ( .A(n6291), .B(n6292), .Z(n6287) );
  NOR U7038 ( .A(n6223), .B(n6222), .Z(n6291) );
  XOR U7039 ( .A(n6293), .B(n6292), .Z(n6222) );
  AND U7040 ( .A(b[2]), .B(a[53]), .Z(n6293) );
  XOR U7041 ( .A(n6292), .B(n6295), .Z(n6294) );
  XNOR U7042 ( .A(n6296), .B(n6297), .Z(n6292) );
  NANDN U7043 ( .A(n6226), .B(n6225), .Z(n6297) );
  XOR U7044 ( .A(n6296), .B(n6298), .Z(n6225) );
  NAND U7045 ( .A(a[53]), .B(b[1]), .Z(n6298) );
  XOR U7046 ( .A(n6296), .B(n6300), .Z(n6299) );
  OR U7047 ( .A(n2632), .B(n2630), .Z(n6296) );
  XOR U7048 ( .A(n6302), .B(n6303), .Z(n2630) );
  NANDN U7049 ( .A(n179), .B(a[53]), .Z(n2632) );
  XNOR U7050 ( .A(n6307), .B(n6199), .Z(n6201) );
  XOR U7051 ( .A(n6308), .B(n6309), .Z(n6199) );
  ANDN U7052 ( .B(n6285), .A(n6306), .Z(n6308) );
  XNOR U7053 ( .A(n6310), .B(n6309), .Z(n6306) );
  AND U7054 ( .A(a[52]), .B(b[5]), .Z(n6310) );
  XNOR U7055 ( .A(n6309), .B(n6279), .Z(n6311) );
  XNOR U7056 ( .A(n6278), .B(n6274), .Z(n6312) );
  XNOR U7057 ( .A(n6273), .B(n6269), .Z(n6313) );
  XNOR U7058 ( .A(n6268), .B(n6264), .Z(n6314) );
  XNOR U7059 ( .A(n6263), .B(n6259), .Z(n6315) );
  XNOR U7060 ( .A(n6258), .B(n6254), .Z(n6316) );
  XOR U7061 ( .A(n6253), .B(n6250), .Z(n6317) );
  XOR U7062 ( .A(n6318), .B(n6319), .Z(n6250) );
  XOR U7063 ( .A(n6248), .B(n6320), .Z(n6319) );
  XOR U7064 ( .A(n6321), .B(n6322), .Z(n6320) );
  XOR U7065 ( .A(n6323), .B(n6324), .Z(n6322) );
  NAND U7066 ( .A(a[43]), .B(b[14]), .Z(n6324) );
  AND U7067 ( .A(a[42]), .B(b[15]), .Z(n6323) );
  XOR U7068 ( .A(n6325), .B(n6321), .Z(n6318) );
  XOR U7069 ( .A(n6326), .B(n6327), .Z(n6321) );
  NOR U7070 ( .A(n6328), .B(n6329), .Z(n6326) );
  AND U7071 ( .A(a[44]), .B(b[13]), .Z(n6325) );
  XNOR U7072 ( .A(n6330), .B(n6248), .Z(n6249) );
  XOR U7073 ( .A(n6331), .B(n6332), .Z(n6248) );
  ANDN U7074 ( .B(n6333), .A(n6334), .Z(n6331) );
  AND U7075 ( .A(a[45]), .B(b[12]), .Z(n6330) );
  XNOR U7076 ( .A(n6335), .B(n6253), .Z(n6255) );
  XOR U7077 ( .A(n6336), .B(n6337), .Z(n6253) );
  ANDN U7078 ( .B(n6338), .A(n6339), .Z(n6336) );
  AND U7079 ( .A(a[46]), .B(b[11]), .Z(n6335) );
  XNOR U7080 ( .A(n6340), .B(n6258), .Z(n6260) );
  XOR U7081 ( .A(n6341), .B(n6342), .Z(n6258) );
  ANDN U7082 ( .B(n6343), .A(n6344), .Z(n6341) );
  AND U7083 ( .A(a[47]), .B(b[10]), .Z(n6340) );
  XNOR U7084 ( .A(n6345), .B(n6263), .Z(n6265) );
  XOR U7085 ( .A(n6346), .B(n6347), .Z(n6263) );
  ANDN U7086 ( .B(n6348), .A(n6349), .Z(n6346) );
  AND U7087 ( .A(a[48]), .B(b[9]), .Z(n6345) );
  XNOR U7088 ( .A(n6350), .B(n6268), .Z(n6270) );
  XOR U7089 ( .A(n6351), .B(n6352), .Z(n6268) );
  ANDN U7090 ( .B(n6353), .A(n6354), .Z(n6351) );
  AND U7091 ( .A(a[49]), .B(b[8]), .Z(n6350) );
  XNOR U7092 ( .A(n6355), .B(n6273), .Z(n6275) );
  XOR U7093 ( .A(n6356), .B(n6357), .Z(n6273) );
  ANDN U7094 ( .B(n6358), .A(n6359), .Z(n6356) );
  AND U7095 ( .A(a[50]), .B(b[7]), .Z(n6355) );
  XOR U7096 ( .A(n6360), .B(n6361), .Z(n6309) );
  ANDN U7097 ( .B(n6290), .A(n6305), .Z(n6360) );
  XNOR U7098 ( .A(n6362), .B(n6361), .Z(n6305) );
  AND U7099 ( .A(a[52]), .B(b[4]), .Z(n6362) );
  XNOR U7100 ( .A(n6361), .B(n6364), .Z(n6363) );
  XOR U7101 ( .A(n6365), .B(n6366), .Z(n6361) );
  ANDN U7102 ( .B(n6295), .A(n6304), .Z(n6365) );
  XNOR U7103 ( .A(n6367), .B(n6366), .Z(n6304) );
  AND U7104 ( .A(a[52]), .B(b[3]), .Z(n6367) );
  XNOR U7105 ( .A(n6366), .B(n6369), .Z(n6368) );
  XNOR U7106 ( .A(n6370), .B(n6371), .Z(n6366) );
  ANDN U7107 ( .B(n6300), .A(n6301), .Z(n6370) );
  XOR U7108 ( .A(n6372), .B(n6371), .Z(n6301) );
  IV U7109 ( .A(n6373), .Z(n6371) );
  AND U7110 ( .A(b[2]), .B(a[52]), .Z(n6372) );
  XNOR U7111 ( .A(n6375), .B(n6373), .Z(n6374) );
  XOR U7112 ( .A(n6376), .B(n6377), .Z(n6373) );
  NANDN U7113 ( .A(n6303), .B(n6302), .Z(n6377) );
  XOR U7114 ( .A(n6376), .B(n6378), .Z(n6302) );
  NAND U7115 ( .A(a[52]), .B(b[1]), .Z(n6378) );
  XOR U7116 ( .A(n6376), .B(n6380), .Z(n6379) );
  OR U7117 ( .A(n2637), .B(n2635), .Z(n6376) );
  XOR U7118 ( .A(n6382), .B(n6383), .Z(n2635) );
  NANDN U7119 ( .A(n179), .B(a[52]), .Z(n2637) );
  XNOR U7120 ( .A(n6387), .B(n6278), .Z(n6280) );
  XOR U7121 ( .A(n6388), .B(n6389), .Z(n6278) );
  ANDN U7122 ( .B(n6364), .A(n6386), .Z(n6388) );
  XNOR U7123 ( .A(n6390), .B(n6389), .Z(n6386) );
  AND U7124 ( .A(a[51]), .B(b[5]), .Z(n6390) );
  XNOR U7125 ( .A(n6389), .B(n6358), .Z(n6391) );
  XNOR U7126 ( .A(n6357), .B(n6353), .Z(n6392) );
  XNOR U7127 ( .A(n6352), .B(n6348), .Z(n6393) );
  XNOR U7128 ( .A(n6347), .B(n6343), .Z(n6394) );
  XNOR U7129 ( .A(n6342), .B(n6338), .Z(n6395) );
  XNOR U7130 ( .A(n6337), .B(n6333), .Z(n6396) );
  XOR U7131 ( .A(n6332), .B(n6329), .Z(n6397) );
  XOR U7132 ( .A(n6398), .B(n6399), .Z(n6329) );
  XOR U7133 ( .A(n6327), .B(n6400), .Z(n6399) );
  XOR U7134 ( .A(n6401), .B(n6402), .Z(n6400) );
  XOR U7135 ( .A(n6403), .B(n6404), .Z(n6402) );
  NAND U7136 ( .A(a[42]), .B(b[14]), .Z(n6404) );
  AND U7137 ( .A(a[41]), .B(b[15]), .Z(n6403) );
  XOR U7138 ( .A(n6405), .B(n6401), .Z(n6398) );
  XOR U7139 ( .A(n6406), .B(n6407), .Z(n6401) );
  NOR U7140 ( .A(n6408), .B(n6409), .Z(n6406) );
  AND U7141 ( .A(a[43]), .B(b[13]), .Z(n6405) );
  XNOR U7142 ( .A(n6410), .B(n6327), .Z(n6328) );
  XOR U7143 ( .A(n6411), .B(n6412), .Z(n6327) );
  ANDN U7144 ( .B(n6413), .A(n6414), .Z(n6411) );
  AND U7145 ( .A(a[44]), .B(b[12]), .Z(n6410) );
  XNOR U7146 ( .A(n6415), .B(n6332), .Z(n6334) );
  XOR U7147 ( .A(n6416), .B(n6417), .Z(n6332) );
  ANDN U7148 ( .B(n6418), .A(n6419), .Z(n6416) );
  AND U7149 ( .A(a[45]), .B(b[11]), .Z(n6415) );
  XNOR U7150 ( .A(n6420), .B(n6337), .Z(n6339) );
  XOR U7151 ( .A(n6421), .B(n6422), .Z(n6337) );
  ANDN U7152 ( .B(n6423), .A(n6424), .Z(n6421) );
  AND U7153 ( .A(a[46]), .B(b[10]), .Z(n6420) );
  XNOR U7154 ( .A(n6425), .B(n6342), .Z(n6344) );
  XOR U7155 ( .A(n6426), .B(n6427), .Z(n6342) );
  ANDN U7156 ( .B(n6428), .A(n6429), .Z(n6426) );
  AND U7157 ( .A(a[47]), .B(b[9]), .Z(n6425) );
  XNOR U7158 ( .A(n6430), .B(n6347), .Z(n6349) );
  XOR U7159 ( .A(n6431), .B(n6432), .Z(n6347) );
  ANDN U7160 ( .B(n6433), .A(n6434), .Z(n6431) );
  AND U7161 ( .A(a[48]), .B(b[8]), .Z(n6430) );
  XNOR U7162 ( .A(n6435), .B(n6352), .Z(n6354) );
  XOR U7163 ( .A(n6436), .B(n6437), .Z(n6352) );
  ANDN U7164 ( .B(n6438), .A(n6439), .Z(n6436) );
  AND U7165 ( .A(a[49]), .B(b[7]), .Z(n6435) );
  XOR U7166 ( .A(n6440), .B(n6441), .Z(n6389) );
  ANDN U7167 ( .B(n6369), .A(n6385), .Z(n6440) );
  XNOR U7168 ( .A(n6442), .B(n6441), .Z(n6385) );
  AND U7169 ( .A(a[51]), .B(b[4]), .Z(n6442) );
  XNOR U7170 ( .A(n6441), .B(n6444), .Z(n6443) );
  XNOR U7171 ( .A(n6445), .B(n6446), .Z(n6441) );
  ANDN U7172 ( .B(n6375), .A(n6384), .Z(n6445) );
  XOR U7173 ( .A(n6447), .B(n6446), .Z(n6384) );
  IV U7174 ( .A(n6448), .Z(n6446) );
  AND U7175 ( .A(a[51]), .B(b[3]), .Z(n6447) );
  XNOR U7176 ( .A(n6450), .B(n6448), .Z(n6449) );
  XOR U7177 ( .A(n6451), .B(n6452), .Z(n6448) );
  ANDN U7178 ( .B(n6380), .A(n6381), .Z(n6451) );
  AND U7179 ( .A(b[2]), .B(a[51]), .Z(n6453) );
  XNOR U7180 ( .A(n6455), .B(n6452), .Z(n6454) );
  XOR U7181 ( .A(n6456), .B(n6457), .Z(n6452) );
  NANDN U7182 ( .A(n6383), .B(n6382), .Z(n6457) );
  XOR U7183 ( .A(n6456), .B(n6458), .Z(n6382) );
  NAND U7184 ( .A(a[51]), .B(b[1]), .Z(n6458) );
  XOR U7185 ( .A(n6456), .B(n6460), .Z(n6459) );
  OR U7186 ( .A(n2642), .B(n2640), .Z(n6456) );
  XOR U7187 ( .A(n6462), .B(n6463), .Z(n2640) );
  NANDN U7188 ( .A(n179), .B(a[51]), .Z(n2642) );
  XNOR U7189 ( .A(n6467), .B(n6357), .Z(n6359) );
  XOR U7190 ( .A(n6468), .B(n6469), .Z(n6357) );
  ANDN U7191 ( .B(n6444), .A(n6466), .Z(n6468) );
  XNOR U7192 ( .A(n6470), .B(n6469), .Z(n6466) );
  AND U7193 ( .A(a[50]), .B(b[5]), .Z(n6470) );
  XNOR U7194 ( .A(n6469), .B(n6438), .Z(n6471) );
  XNOR U7195 ( .A(n6437), .B(n6433), .Z(n6472) );
  XNOR U7196 ( .A(n6432), .B(n6428), .Z(n6473) );
  XNOR U7197 ( .A(n6427), .B(n6423), .Z(n6474) );
  XNOR U7198 ( .A(n6422), .B(n6418), .Z(n6475) );
  XNOR U7199 ( .A(n6417), .B(n6413), .Z(n6476) );
  XOR U7200 ( .A(n6412), .B(n6409), .Z(n6477) );
  XOR U7201 ( .A(n6478), .B(n6479), .Z(n6409) );
  XOR U7202 ( .A(n6407), .B(n6480), .Z(n6479) );
  XNOR U7203 ( .A(n6481), .B(n6482), .Z(n6480) );
  XOR U7204 ( .A(n6483), .B(n6484), .Z(n6482) );
  NAND U7205 ( .A(a[41]), .B(b[14]), .Z(n6484) );
  AND U7206 ( .A(a[40]), .B(b[15]), .Z(n6483) );
  XNOR U7207 ( .A(n6485), .B(n6481), .Z(n6478) );
  XOR U7208 ( .A(n6486), .B(n6487), .Z(n6481) );
  NOR U7209 ( .A(n6488), .B(n6489), .Z(n6486) );
  AND U7210 ( .A(a[42]), .B(b[13]), .Z(n6485) );
  XNOR U7211 ( .A(n6490), .B(n6407), .Z(n6408) );
  XNOR U7212 ( .A(n6491), .B(n6492), .Z(n6407) );
  ANDN U7213 ( .B(n6493), .A(n6494), .Z(n6491) );
  AND U7214 ( .A(a[43]), .B(b[12]), .Z(n6490) );
  XNOR U7215 ( .A(n6495), .B(n6412), .Z(n6414) );
  XNOR U7216 ( .A(n6496), .B(n6497), .Z(n6412) );
  ANDN U7217 ( .B(n6498), .A(n6499), .Z(n6496) );
  AND U7218 ( .A(a[44]), .B(b[11]), .Z(n6495) );
  XNOR U7219 ( .A(n6500), .B(n6417), .Z(n6419) );
  XNOR U7220 ( .A(n6501), .B(n6502), .Z(n6417) );
  ANDN U7221 ( .B(n6503), .A(n6504), .Z(n6501) );
  AND U7222 ( .A(a[45]), .B(b[10]), .Z(n6500) );
  XNOR U7223 ( .A(n6505), .B(n6422), .Z(n6424) );
  XNOR U7224 ( .A(n6506), .B(n6507), .Z(n6422) );
  ANDN U7225 ( .B(n6508), .A(n6509), .Z(n6506) );
  AND U7226 ( .A(a[46]), .B(b[9]), .Z(n6505) );
  XNOR U7227 ( .A(n6510), .B(n6427), .Z(n6429) );
  XNOR U7228 ( .A(n6511), .B(n6512), .Z(n6427) );
  ANDN U7229 ( .B(n6513), .A(n6514), .Z(n6511) );
  AND U7230 ( .A(a[47]), .B(b[8]), .Z(n6510) );
  XNOR U7231 ( .A(n6515), .B(n6432), .Z(n6434) );
  XNOR U7232 ( .A(n6516), .B(n6517), .Z(n6432) );
  ANDN U7233 ( .B(n6518), .A(n6519), .Z(n6516) );
  AND U7234 ( .A(a[48]), .B(b[7]), .Z(n6515) );
  XNOR U7235 ( .A(n6520), .B(n6521), .Z(n6469) );
  ANDN U7236 ( .B(n6450), .A(n6465), .Z(n6520) );
  XOR U7237 ( .A(n6522), .B(n6521), .Z(n6465) );
  IV U7238 ( .A(n6523), .Z(n6521) );
  AND U7239 ( .A(a[50]), .B(b[4]), .Z(n6522) );
  XNOR U7240 ( .A(n6525), .B(n6523), .Z(n6524) );
  XOR U7241 ( .A(n6526), .B(n6527), .Z(n6523) );
  ANDN U7242 ( .B(n6455), .A(n6464), .Z(n6526) );
  AND U7243 ( .A(a[50]), .B(b[3]), .Z(n6528) );
  XNOR U7244 ( .A(n6530), .B(n6527), .Z(n6529) );
  XOR U7245 ( .A(n6531), .B(n6532), .Z(n6527) );
  ANDN U7246 ( .B(n6460), .A(n6461), .Z(n6531) );
  AND U7247 ( .A(b[2]), .B(a[50]), .Z(n6533) );
  XNOR U7248 ( .A(n6535), .B(n6532), .Z(n6534) );
  XOR U7249 ( .A(n6536), .B(n6537), .Z(n6532) );
  NANDN U7250 ( .A(n6463), .B(n6462), .Z(n6537) );
  XOR U7251 ( .A(n6536), .B(n6538), .Z(n6462) );
  NAND U7252 ( .A(a[50]), .B(b[1]), .Z(n6538) );
  XOR U7253 ( .A(n6536), .B(n6540), .Z(n6539) );
  OR U7254 ( .A(n2647), .B(n2645), .Z(n6536) );
  XOR U7255 ( .A(n6542), .B(n6543), .Z(n2645) );
  NANDN U7256 ( .A(n179), .B(a[50]), .Z(n2647) );
  XNOR U7257 ( .A(n6547), .B(n6437), .Z(n6439) );
  XNOR U7258 ( .A(n6548), .B(n6549), .Z(n6437) );
  ANDN U7259 ( .B(n6525), .A(n6546), .Z(n6548) );
  XOR U7260 ( .A(n6550), .B(n6549), .Z(n6546) );
  IV U7261 ( .A(n6551), .Z(n6549) );
  AND U7262 ( .A(a[49]), .B(b[5]), .Z(n6550) );
  XNOR U7263 ( .A(n6518), .B(n6551), .Z(n6552) );
  XOR U7264 ( .A(n6553), .B(n6554), .Z(n6551) );
  ANDN U7265 ( .B(n6530), .A(n6545), .Z(n6553) );
  AND U7266 ( .A(a[49]), .B(b[4]), .Z(n6555) );
  XNOR U7267 ( .A(n6557), .B(n6554), .Z(n6556) );
  XOR U7268 ( .A(n6558), .B(n6559), .Z(n6554) );
  ANDN U7269 ( .B(n6535), .A(n6544), .Z(n6558) );
  AND U7270 ( .A(a[49]), .B(b[3]), .Z(n6560) );
  XNOR U7271 ( .A(n6562), .B(n6559), .Z(n6561) );
  XOR U7272 ( .A(n6563), .B(n6564), .Z(n6559) );
  ANDN U7273 ( .B(n6540), .A(n6541), .Z(n6563) );
  AND U7274 ( .A(b[2]), .B(a[49]), .Z(n6565) );
  XNOR U7275 ( .A(n6567), .B(n6564), .Z(n6566) );
  XOR U7276 ( .A(n6568), .B(n6569), .Z(n6564) );
  NANDN U7277 ( .A(n6543), .B(n6542), .Z(n6569) );
  XOR U7278 ( .A(n6568), .B(n6570), .Z(n6542) );
  NAND U7279 ( .A(a[49]), .B(b[1]), .Z(n6570) );
  XOR U7280 ( .A(n6568), .B(n6572), .Z(n6571) );
  OR U7281 ( .A(n2652), .B(n2650), .Z(n6568) );
  XOR U7282 ( .A(n6574), .B(n6575), .Z(n2650) );
  NANDN U7283 ( .A(n179), .B(a[49]), .Z(n2652) );
  XNOR U7284 ( .A(n6513), .B(n6580), .Z(n6579) );
  XNOR U7285 ( .A(n6508), .B(n6582), .Z(n6581) );
  XNOR U7286 ( .A(n6503), .B(n6584), .Z(n6583) );
  XNOR U7287 ( .A(n6498), .B(n6586), .Z(n6585) );
  XNOR U7288 ( .A(n6493), .B(n6588), .Z(n6587) );
  XOR U7289 ( .A(n6489), .B(n6590), .Z(n6589) );
  XOR U7290 ( .A(n6591), .B(n6592), .Z(n6489) );
  XNOR U7291 ( .A(n6593), .B(n6594), .Z(n6592) );
  XNOR U7292 ( .A(n6595), .B(n6596), .Z(n6593) );
  XOR U7293 ( .A(n6597), .B(n6598), .Z(n6596) );
  AND U7294 ( .A(b[15]), .B(a[39]), .Z(n6598) );
  AND U7295 ( .A(a[40]), .B(b[14]), .Z(n6597) );
  XNOR U7296 ( .A(n6599), .B(n6595), .Z(n6591) );
  XOR U7297 ( .A(n6600), .B(n6601), .Z(n6595) );
  NOR U7298 ( .A(n6602), .B(n6603), .Z(n6600) );
  AND U7299 ( .A(a[41]), .B(b[13]), .Z(n6599) );
  XOR U7300 ( .A(n6604), .B(n6487), .Z(n6488) );
  IV U7301 ( .A(n6594), .Z(n6487) );
  XOR U7302 ( .A(n6605), .B(n6606), .Z(n6594) );
  ANDN U7303 ( .B(n6607), .A(n6608), .Z(n6605) );
  AND U7304 ( .A(a[42]), .B(b[12]), .Z(n6604) );
  XOR U7305 ( .A(n6609), .B(n6492), .Z(n6494) );
  IV U7306 ( .A(n6590), .Z(n6492) );
  XOR U7307 ( .A(n6610), .B(n6611), .Z(n6590) );
  ANDN U7308 ( .B(n6612), .A(n6613), .Z(n6610) );
  AND U7309 ( .A(a[43]), .B(b[11]), .Z(n6609) );
  XOR U7310 ( .A(n6614), .B(n6497), .Z(n6499) );
  IV U7311 ( .A(n6588), .Z(n6497) );
  XOR U7312 ( .A(n6615), .B(n6616), .Z(n6588) );
  ANDN U7313 ( .B(n6617), .A(n6618), .Z(n6615) );
  AND U7314 ( .A(a[44]), .B(b[10]), .Z(n6614) );
  XOR U7315 ( .A(n6619), .B(n6502), .Z(n6504) );
  IV U7316 ( .A(n6586), .Z(n6502) );
  XOR U7317 ( .A(n6620), .B(n6621), .Z(n6586) );
  ANDN U7318 ( .B(n6622), .A(n6623), .Z(n6620) );
  AND U7319 ( .A(a[45]), .B(b[9]), .Z(n6619) );
  XOR U7320 ( .A(n6624), .B(n6507), .Z(n6509) );
  IV U7321 ( .A(n6584), .Z(n6507) );
  XOR U7322 ( .A(n6625), .B(n6626), .Z(n6584) );
  ANDN U7323 ( .B(n6627), .A(n6628), .Z(n6625) );
  AND U7324 ( .A(a[46]), .B(b[8]), .Z(n6624) );
  XOR U7325 ( .A(n6629), .B(n6512), .Z(n6514) );
  IV U7326 ( .A(n6582), .Z(n6512) );
  XOR U7327 ( .A(n6630), .B(n6631), .Z(n6582) );
  ANDN U7328 ( .B(n6632), .A(n6633), .Z(n6630) );
  AND U7329 ( .A(a[47]), .B(b[7]), .Z(n6629) );
  XOR U7330 ( .A(n6634), .B(n6517), .Z(n6519) );
  IV U7331 ( .A(n6580), .Z(n6517) );
  XOR U7332 ( .A(n6635), .B(n6636), .Z(n6580) );
  ANDN U7333 ( .B(n6557), .A(n6578), .Z(n6635) );
  AND U7334 ( .A(a[48]), .B(b[5]), .Z(n6637) );
  XNOR U7335 ( .A(n6632), .B(n6636), .Z(n6638) );
  XOR U7336 ( .A(n6639), .B(n6640), .Z(n6636) );
  ANDN U7337 ( .B(n6562), .A(n6577), .Z(n6639) );
  AND U7338 ( .A(a[48]), .B(b[4]), .Z(n6641) );
  XNOR U7339 ( .A(n6643), .B(n6640), .Z(n6642) );
  XOR U7340 ( .A(n6644), .B(n6645), .Z(n6640) );
  ANDN U7341 ( .B(n6567), .A(n6576), .Z(n6644) );
  AND U7342 ( .A(a[48]), .B(b[3]), .Z(n6646) );
  XNOR U7343 ( .A(n6648), .B(n6645), .Z(n6647) );
  XOR U7344 ( .A(n6649), .B(n6650), .Z(n6645) );
  ANDN U7345 ( .B(n6572), .A(n6573), .Z(n6649) );
  AND U7346 ( .A(b[2]), .B(a[48]), .Z(n6651) );
  XNOR U7347 ( .A(n6653), .B(n6650), .Z(n6652) );
  XOR U7348 ( .A(n6654), .B(n6655), .Z(n6650) );
  NANDN U7349 ( .A(n6575), .B(n6574), .Z(n6655) );
  XOR U7350 ( .A(n6654), .B(n6656), .Z(n6574) );
  NAND U7351 ( .A(a[48]), .B(b[1]), .Z(n6656) );
  XOR U7352 ( .A(n6654), .B(n6658), .Z(n6657) );
  OR U7353 ( .A(n2657), .B(n2655), .Z(n6654) );
  XOR U7354 ( .A(n6660), .B(n6661), .Z(n2655) );
  NANDN U7355 ( .A(n179), .B(a[48]), .Z(n2657) );
  XNOR U7356 ( .A(n6627), .B(n6631), .Z(n6665) );
  XNOR U7357 ( .A(n6622), .B(n6626), .Z(n6666) );
  XNOR U7358 ( .A(n6617), .B(n6621), .Z(n6667) );
  XNOR U7359 ( .A(n6612), .B(n6616), .Z(n6668) );
  XNOR U7360 ( .A(n6607), .B(n6611), .Z(n6669) );
  XOR U7361 ( .A(n6603), .B(n6606), .Z(n6670) );
  XOR U7362 ( .A(n6671), .B(n6672), .Z(n6603) );
  XNOR U7363 ( .A(n6673), .B(n6674), .Z(n6672) );
  XNOR U7364 ( .A(n6675), .B(n6676), .Z(n6673) );
  XOR U7365 ( .A(n6677), .B(n6678), .Z(n6676) );
  AND U7366 ( .A(b[14]), .B(a[39]), .Z(n6678) );
  AND U7367 ( .A(a[38]), .B(b[15]), .Z(n6677) );
  XNOR U7368 ( .A(n6679), .B(n6675), .Z(n6671) );
  XOR U7369 ( .A(n6680), .B(n6681), .Z(n6675) );
  NOR U7370 ( .A(n6682), .B(n6683), .Z(n6680) );
  AND U7371 ( .A(a[40]), .B(b[13]), .Z(n6679) );
  XOR U7372 ( .A(n6684), .B(n6601), .Z(n6602) );
  IV U7373 ( .A(n6674), .Z(n6601) );
  XOR U7374 ( .A(n6685), .B(n6686), .Z(n6674) );
  ANDN U7375 ( .B(n6687), .A(n6688), .Z(n6685) );
  AND U7376 ( .A(a[41]), .B(b[12]), .Z(n6684) );
  XOR U7377 ( .A(n6690), .B(n6691), .Z(n6606) );
  ANDN U7378 ( .B(n6692), .A(n6693), .Z(n6690) );
  AND U7379 ( .A(a[42]), .B(b[11]), .Z(n6689) );
  XOR U7380 ( .A(n6695), .B(n6696), .Z(n6611) );
  ANDN U7381 ( .B(n6697), .A(n6698), .Z(n6695) );
  AND U7382 ( .A(a[43]), .B(b[10]), .Z(n6694) );
  XOR U7383 ( .A(n6700), .B(n6701), .Z(n6616) );
  ANDN U7384 ( .B(n6702), .A(n6703), .Z(n6700) );
  AND U7385 ( .A(a[44]), .B(b[9]), .Z(n6699) );
  XOR U7386 ( .A(n6705), .B(n6706), .Z(n6621) );
  ANDN U7387 ( .B(n6707), .A(n6708), .Z(n6705) );
  AND U7388 ( .A(a[45]), .B(b[8]), .Z(n6704) );
  XOR U7389 ( .A(n6710), .B(n6711), .Z(n6626) );
  ANDN U7390 ( .B(n6712), .A(n6713), .Z(n6710) );
  AND U7391 ( .A(a[46]), .B(b[7]), .Z(n6709) );
  XOR U7392 ( .A(n6715), .B(n6716), .Z(n6631) );
  ANDN U7393 ( .B(n6643), .A(n6664), .Z(n6715) );
  AND U7394 ( .A(a[47]), .B(b[5]), .Z(n6717) );
  XNOR U7395 ( .A(n6712), .B(n6716), .Z(n6718) );
  XOR U7396 ( .A(n6719), .B(n6720), .Z(n6716) );
  ANDN U7397 ( .B(n6648), .A(n6663), .Z(n6719) );
  AND U7398 ( .A(a[47]), .B(b[4]), .Z(n6721) );
  XNOR U7399 ( .A(n6723), .B(n6720), .Z(n6722) );
  XOR U7400 ( .A(n6724), .B(n6725), .Z(n6720) );
  ANDN U7401 ( .B(n6653), .A(n6662), .Z(n6724) );
  AND U7402 ( .A(a[47]), .B(b[3]), .Z(n6726) );
  XNOR U7403 ( .A(n6728), .B(n6725), .Z(n6727) );
  XOR U7404 ( .A(n6729), .B(n6730), .Z(n6725) );
  ANDN U7405 ( .B(n6658), .A(n6659), .Z(n6729) );
  AND U7406 ( .A(b[2]), .B(a[47]), .Z(n6731) );
  XNOR U7407 ( .A(n6733), .B(n6730), .Z(n6732) );
  XOR U7408 ( .A(n6734), .B(n6735), .Z(n6730) );
  NANDN U7409 ( .A(n6661), .B(n6660), .Z(n6735) );
  XOR U7410 ( .A(n6734), .B(n6736), .Z(n6660) );
  NAND U7411 ( .A(a[47]), .B(b[1]), .Z(n6736) );
  XOR U7412 ( .A(n6734), .B(n6738), .Z(n6737) );
  OR U7413 ( .A(n2662), .B(n2660), .Z(n6734) );
  XOR U7414 ( .A(n6740), .B(n6741), .Z(n2660) );
  NANDN U7415 ( .A(n179), .B(a[47]), .Z(n2662) );
  XNOR U7416 ( .A(n6707), .B(n6711), .Z(n6745) );
  XNOR U7417 ( .A(n6702), .B(n6706), .Z(n6746) );
  XNOR U7418 ( .A(n6697), .B(n6701), .Z(n6747) );
  XNOR U7419 ( .A(n6692), .B(n6696), .Z(n6748) );
  XNOR U7420 ( .A(n6687), .B(n6691), .Z(n6749) );
  XOR U7421 ( .A(n6683), .B(n6686), .Z(n6750) );
  XOR U7422 ( .A(n6751), .B(n6752), .Z(n6683) );
  XNOR U7423 ( .A(n6753), .B(n6754), .Z(n6752) );
  XOR U7424 ( .A(n6755), .B(n6756), .Z(n6753) );
  AND U7425 ( .A(b[13]), .B(a[39]), .Z(n6755) );
  XOR U7426 ( .A(n6756), .B(n6757), .Z(n6751) );
  XOR U7427 ( .A(n6758), .B(n6759), .Z(n6757) );
  AND U7428 ( .A(a[38]), .B(b[14]), .Z(n6759) );
  AND U7429 ( .A(a[37]), .B(b[15]), .Z(n6758) );
  XOR U7430 ( .A(n6760), .B(n6761), .Z(n6756) );
  ANDN U7431 ( .B(n6762), .A(n6763), .Z(n6760) );
  XOR U7432 ( .A(n6764), .B(n6681), .Z(n6682) );
  IV U7433 ( .A(n6754), .Z(n6681) );
  XOR U7434 ( .A(n6765), .B(n6766), .Z(n6754) );
  NOR U7435 ( .A(n6767), .B(n6768), .Z(n6765) );
  AND U7436 ( .A(a[40]), .B(b[12]), .Z(n6764) );
  XOR U7437 ( .A(n6770), .B(n6771), .Z(n6686) );
  ANDN U7438 ( .B(n6772), .A(n6773), .Z(n6770) );
  AND U7439 ( .A(a[41]), .B(b[11]), .Z(n6769) );
  XOR U7440 ( .A(n6775), .B(n6776), .Z(n6691) );
  ANDN U7441 ( .B(n6777), .A(n6778), .Z(n6775) );
  AND U7442 ( .A(a[42]), .B(b[10]), .Z(n6774) );
  XOR U7443 ( .A(n6780), .B(n6781), .Z(n6696) );
  ANDN U7444 ( .B(n6782), .A(n6783), .Z(n6780) );
  AND U7445 ( .A(a[43]), .B(b[9]), .Z(n6779) );
  XOR U7446 ( .A(n6785), .B(n6786), .Z(n6701) );
  ANDN U7447 ( .B(n6787), .A(n6788), .Z(n6785) );
  AND U7448 ( .A(a[44]), .B(b[8]), .Z(n6784) );
  XOR U7449 ( .A(n6790), .B(n6791), .Z(n6706) );
  ANDN U7450 ( .B(n6792), .A(n6793), .Z(n6790) );
  AND U7451 ( .A(a[45]), .B(b[7]), .Z(n6789) );
  XOR U7452 ( .A(n6795), .B(n6796), .Z(n6711) );
  ANDN U7453 ( .B(n6723), .A(n6744), .Z(n6795) );
  AND U7454 ( .A(a[46]), .B(b[5]), .Z(n6797) );
  XNOR U7455 ( .A(n6792), .B(n6796), .Z(n6798) );
  XOR U7456 ( .A(n6799), .B(n6800), .Z(n6796) );
  ANDN U7457 ( .B(n6728), .A(n6743), .Z(n6799) );
  AND U7458 ( .A(a[46]), .B(b[4]), .Z(n6801) );
  XNOR U7459 ( .A(n6803), .B(n6800), .Z(n6802) );
  XOR U7460 ( .A(n6804), .B(n6805), .Z(n6800) );
  ANDN U7461 ( .B(n6733), .A(n6742), .Z(n6804) );
  AND U7462 ( .A(a[46]), .B(b[3]), .Z(n6806) );
  XNOR U7463 ( .A(n6808), .B(n6805), .Z(n6807) );
  XOR U7464 ( .A(n6809), .B(n6810), .Z(n6805) );
  ANDN U7465 ( .B(n6738), .A(n6739), .Z(n6809) );
  AND U7466 ( .A(b[2]), .B(a[46]), .Z(n6811) );
  XNOR U7467 ( .A(n6813), .B(n6810), .Z(n6812) );
  XOR U7468 ( .A(n6814), .B(n6815), .Z(n6810) );
  NANDN U7469 ( .A(n6741), .B(n6740), .Z(n6815) );
  XOR U7470 ( .A(n6814), .B(n6816), .Z(n6740) );
  NAND U7471 ( .A(a[46]), .B(b[1]), .Z(n6816) );
  XOR U7472 ( .A(n6814), .B(n6818), .Z(n6817) );
  OR U7473 ( .A(n2667), .B(n2665), .Z(n6814) );
  XOR U7474 ( .A(n6820), .B(n6821), .Z(n2665) );
  NANDN U7475 ( .A(n179), .B(a[46]), .Z(n2667) );
  XNOR U7476 ( .A(n6787), .B(n6791), .Z(n6825) );
  XNOR U7477 ( .A(n6782), .B(n6786), .Z(n6826) );
  XNOR U7478 ( .A(n6777), .B(n6781), .Z(n6827) );
  XNOR U7479 ( .A(n6772), .B(n6776), .Z(n6828) );
  XOR U7480 ( .A(n6768), .B(n6771), .Z(n6829) );
  XNOR U7481 ( .A(n6763), .B(n6830), .Z(n6768) );
  XNOR U7482 ( .A(n6762), .B(n6766), .Z(n6830) );
  XOR U7483 ( .A(n6831), .B(n6761), .Z(n6762) );
  AND U7484 ( .A(b[12]), .B(a[39]), .Z(n6831) );
  XOR U7485 ( .A(n6832), .B(n6833), .Z(n6763) );
  XOR U7486 ( .A(n6761), .B(n6834), .Z(n6833) );
  XOR U7487 ( .A(n6835), .B(n6836), .Z(n6834) );
  XOR U7488 ( .A(n6837), .B(n6838), .Z(n6836) );
  NAND U7489 ( .A(a[37]), .B(b[14]), .Z(n6838) );
  AND U7490 ( .A(a[36]), .B(b[15]), .Z(n6837) );
  XOR U7491 ( .A(n6839), .B(n6840), .Z(n6761) );
  ANDN U7492 ( .B(n6841), .A(n6842), .Z(n6839) );
  XOR U7493 ( .A(n6843), .B(n6835), .Z(n6832) );
  XOR U7494 ( .A(n6844), .B(n6845), .Z(n6835) );
  NOR U7495 ( .A(n6846), .B(n6847), .Z(n6844) );
  AND U7496 ( .A(a[38]), .B(b[13]), .Z(n6843) );
  XOR U7497 ( .A(n6849), .B(n6850), .Z(n6766) );
  ANDN U7498 ( .B(n6851), .A(n6852), .Z(n6849) );
  AND U7499 ( .A(a[40]), .B(b[11]), .Z(n6848) );
  XOR U7500 ( .A(n6854), .B(n6855), .Z(n6771) );
  ANDN U7501 ( .B(n6856), .A(n6857), .Z(n6854) );
  AND U7502 ( .A(a[41]), .B(b[10]), .Z(n6853) );
  XOR U7503 ( .A(n6859), .B(n6860), .Z(n6776) );
  ANDN U7504 ( .B(n6861), .A(n6862), .Z(n6859) );
  AND U7505 ( .A(a[42]), .B(b[9]), .Z(n6858) );
  XOR U7506 ( .A(n6864), .B(n6865), .Z(n6781) );
  ANDN U7507 ( .B(n6866), .A(n6867), .Z(n6864) );
  AND U7508 ( .A(a[43]), .B(b[8]), .Z(n6863) );
  XOR U7509 ( .A(n6869), .B(n6870), .Z(n6786) );
  ANDN U7510 ( .B(n6871), .A(n6872), .Z(n6869) );
  AND U7511 ( .A(a[44]), .B(b[7]), .Z(n6868) );
  XOR U7512 ( .A(n6874), .B(n6875), .Z(n6791) );
  ANDN U7513 ( .B(n6803), .A(n6824), .Z(n6874) );
  AND U7514 ( .A(a[45]), .B(b[5]), .Z(n6876) );
  XNOR U7515 ( .A(n6871), .B(n6875), .Z(n6877) );
  XOR U7516 ( .A(n6878), .B(n6879), .Z(n6875) );
  ANDN U7517 ( .B(n6808), .A(n6823), .Z(n6878) );
  AND U7518 ( .A(a[45]), .B(b[4]), .Z(n6880) );
  XNOR U7519 ( .A(n6882), .B(n6879), .Z(n6881) );
  XOR U7520 ( .A(n6883), .B(n6884), .Z(n6879) );
  ANDN U7521 ( .B(n6813), .A(n6822), .Z(n6883) );
  AND U7522 ( .A(a[45]), .B(b[3]), .Z(n6885) );
  XNOR U7523 ( .A(n6887), .B(n6884), .Z(n6886) );
  XOR U7524 ( .A(n6888), .B(n6889), .Z(n6884) );
  ANDN U7525 ( .B(n6818), .A(n6819), .Z(n6888) );
  AND U7526 ( .A(b[2]), .B(a[45]), .Z(n6890) );
  XNOR U7527 ( .A(n6892), .B(n6889), .Z(n6891) );
  XOR U7528 ( .A(n6893), .B(n6894), .Z(n6889) );
  NANDN U7529 ( .A(n6821), .B(n6820), .Z(n6894) );
  XOR U7530 ( .A(n6893), .B(n6895), .Z(n6820) );
  NAND U7531 ( .A(a[45]), .B(b[1]), .Z(n6895) );
  XOR U7532 ( .A(n6893), .B(n6897), .Z(n6896) );
  OR U7533 ( .A(n2672), .B(n2670), .Z(n6893) );
  XOR U7534 ( .A(n6899), .B(n6900), .Z(n2670) );
  NANDN U7535 ( .A(n179), .B(a[45]), .Z(n2672) );
  XNOR U7536 ( .A(n6866), .B(n6870), .Z(n6904) );
  XNOR U7537 ( .A(n6861), .B(n6865), .Z(n6905) );
  XNOR U7538 ( .A(n6856), .B(n6860), .Z(n6906) );
  XNOR U7539 ( .A(n6851), .B(n6855), .Z(n6907) );
  XNOR U7540 ( .A(n6841), .B(n6850), .Z(n6908) );
  XOR U7541 ( .A(n6909), .B(n6840), .Z(n6841) );
  AND U7542 ( .A(b[11]), .B(a[39]), .Z(n6909) );
  XOR U7543 ( .A(n6840), .B(n6847), .Z(n6910) );
  XOR U7544 ( .A(n6911), .B(n6912), .Z(n6847) );
  XOR U7545 ( .A(n6845), .B(n6913), .Z(n6912) );
  XOR U7546 ( .A(n6914), .B(n6915), .Z(n6913) );
  XOR U7547 ( .A(n6916), .B(n6917), .Z(n6915) );
  NAND U7548 ( .A(a[36]), .B(b[14]), .Z(n6917) );
  AND U7549 ( .A(a[35]), .B(b[15]), .Z(n6916) );
  XOR U7550 ( .A(n6918), .B(n6914), .Z(n6911) );
  XOR U7551 ( .A(n6919), .B(n6920), .Z(n6914) );
  NOR U7552 ( .A(n6921), .B(n6922), .Z(n6919) );
  AND U7553 ( .A(a[37]), .B(b[13]), .Z(n6918) );
  XOR U7554 ( .A(n6923), .B(n6924), .Z(n6840) );
  ANDN U7555 ( .B(n6925), .A(n6926), .Z(n6923) );
  XNOR U7556 ( .A(n6927), .B(n6845), .Z(n6846) );
  XOR U7557 ( .A(n6928), .B(n6929), .Z(n6845) );
  ANDN U7558 ( .B(n6930), .A(n6931), .Z(n6928) );
  AND U7559 ( .A(a[38]), .B(b[12]), .Z(n6927) );
  XOR U7560 ( .A(n6933), .B(n6934), .Z(n6850) );
  ANDN U7561 ( .B(n6935), .A(n6936), .Z(n6933) );
  AND U7562 ( .A(a[40]), .B(b[10]), .Z(n6932) );
  XOR U7563 ( .A(n6938), .B(n6939), .Z(n6855) );
  ANDN U7564 ( .B(n6940), .A(n6941), .Z(n6938) );
  AND U7565 ( .A(a[41]), .B(b[9]), .Z(n6937) );
  XOR U7566 ( .A(n6943), .B(n6944), .Z(n6860) );
  ANDN U7567 ( .B(n6945), .A(n6946), .Z(n6943) );
  AND U7568 ( .A(a[42]), .B(b[8]), .Z(n6942) );
  XOR U7569 ( .A(n6948), .B(n6949), .Z(n6865) );
  ANDN U7570 ( .B(n6950), .A(n6951), .Z(n6948) );
  AND U7571 ( .A(a[43]), .B(b[7]), .Z(n6947) );
  XOR U7572 ( .A(n6953), .B(n6954), .Z(n6870) );
  ANDN U7573 ( .B(n6882), .A(n6903), .Z(n6953) );
  AND U7574 ( .A(a[44]), .B(b[5]), .Z(n6955) );
  XNOR U7575 ( .A(n6950), .B(n6954), .Z(n6956) );
  XOR U7576 ( .A(n6957), .B(n6958), .Z(n6954) );
  ANDN U7577 ( .B(n6887), .A(n6902), .Z(n6957) );
  AND U7578 ( .A(a[44]), .B(b[4]), .Z(n6959) );
  XNOR U7579 ( .A(n6961), .B(n6958), .Z(n6960) );
  XOR U7580 ( .A(n6962), .B(n6963), .Z(n6958) );
  ANDN U7581 ( .B(n6892), .A(n6901), .Z(n6962) );
  AND U7582 ( .A(a[44]), .B(b[3]), .Z(n6964) );
  XNOR U7583 ( .A(n6966), .B(n6963), .Z(n6965) );
  XOR U7584 ( .A(n6967), .B(n6968), .Z(n6963) );
  ANDN U7585 ( .B(n6897), .A(n6898), .Z(n6967) );
  AND U7586 ( .A(b[2]), .B(a[44]), .Z(n6969) );
  XNOR U7587 ( .A(n6971), .B(n6968), .Z(n6970) );
  XOR U7588 ( .A(n6972), .B(n6973), .Z(n6968) );
  NANDN U7589 ( .A(n6900), .B(n6899), .Z(n6973) );
  XOR U7590 ( .A(n6972), .B(n6974), .Z(n6899) );
  NAND U7591 ( .A(a[44]), .B(b[1]), .Z(n6974) );
  XOR U7592 ( .A(n6972), .B(n6976), .Z(n6975) );
  OR U7593 ( .A(n2677), .B(n2675), .Z(n6972) );
  XOR U7594 ( .A(n6978), .B(n6979), .Z(n2675) );
  NANDN U7595 ( .A(n179), .B(a[44]), .Z(n2677) );
  XNOR U7596 ( .A(n6945), .B(n6949), .Z(n6983) );
  XNOR U7597 ( .A(n6940), .B(n6944), .Z(n6984) );
  XNOR U7598 ( .A(n6935), .B(n6939), .Z(n6985) );
  XNOR U7599 ( .A(n6925), .B(n6934), .Z(n6986) );
  XOR U7600 ( .A(n6987), .B(n6924), .Z(n6925) );
  AND U7601 ( .A(b[10]), .B(a[39]), .Z(n6987) );
  XNOR U7602 ( .A(n6924), .B(n6930), .Z(n6988) );
  XOR U7603 ( .A(n6929), .B(n6922), .Z(n6989) );
  XOR U7604 ( .A(n6990), .B(n6991), .Z(n6922) );
  XOR U7605 ( .A(n6920), .B(n6992), .Z(n6991) );
  XOR U7606 ( .A(n6993), .B(n6994), .Z(n6992) );
  XOR U7607 ( .A(n6995), .B(n6996), .Z(n6994) );
  NAND U7608 ( .A(a[35]), .B(b[14]), .Z(n6996) );
  AND U7609 ( .A(a[34]), .B(b[15]), .Z(n6995) );
  XOR U7610 ( .A(n6997), .B(n6993), .Z(n6990) );
  XOR U7611 ( .A(n6998), .B(n6999), .Z(n6993) );
  NOR U7612 ( .A(n7000), .B(n7001), .Z(n6998) );
  AND U7613 ( .A(a[36]), .B(b[13]), .Z(n6997) );
  XNOR U7614 ( .A(n7002), .B(n6920), .Z(n6921) );
  XOR U7615 ( .A(n7003), .B(n7004), .Z(n6920) );
  ANDN U7616 ( .B(n7005), .A(n7006), .Z(n7003) );
  AND U7617 ( .A(a[37]), .B(b[12]), .Z(n7002) );
  XOR U7618 ( .A(n7007), .B(n7008), .Z(n6924) );
  ANDN U7619 ( .B(n7009), .A(n7010), .Z(n7007) );
  XNOR U7620 ( .A(n7011), .B(n6929), .Z(n6931) );
  XOR U7621 ( .A(n7012), .B(n7013), .Z(n6929) );
  ANDN U7622 ( .B(n7014), .A(n7015), .Z(n7012) );
  AND U7623 ( .A(a[38]), .B(b[11]), .Z(n7011) );
  XOR U7624 ( .A(n7017), .B(n7018), .Z(n6934) );
  ANDN U7625 ( .B(n7019), .A(n7020), .Z(n7017) );
  AND U7626 ( .A(a[40]), .B(b[9]), .Z(n7016) );
  XOR U7627 ( .A(n7022), .B(n7023), .Z(n6939) );
  ANDN U7628 ( .B(n7024), .A(n7025), .Z(n7022) );
  AND U7629 ( .A(a[41]), .B(b[8]), .Z(n7021) );
  XOR U7630 ( .A(n7027), .B(n7028), .Z(n6944) );
  ANDN U7631 ( .B(n7029), .A(n7030), .Z(n7027) );
  AND U7632 ( .A(a[42]), .B(b[7]), .Z(n7026) );
  XOR U7633 ( .A(n7032), .B(n7033), .Z(n6949) );
  ANDN U7634 ( .B(n6961), .A(n6982), .Z(n7032) );
  AND U7635 ( .A(a[43]), .B(b[5]), .Z(n7034) );
  XNOR U7636 ( .A(n7029), .B(n7033), .Z(n7035) );
  XOR U7637 ( .A(n7036), .B(n7037), .Z(n7033) );
  ANDN U7638 ( .B(n6966), .A(n6981), .Z(n7036) );
  AND U7639 ( .A(a[43]), .B(b[4]), .Z(n7038) );
  XNOR U7640 ( .A(n7040), .B(n7037), .Z(n7039) );
  XOR U7641 ( .A(n7041), .B(n7042), .Z(n7037) );
  ANDN U7642 ( .B(n6971), .A(n6980), .Z(n7041) );
  AND U7643 ( .A(a[43]), .B(b[3]), .Z(n7043) );
  XNOR U7644 ( .A(n7045), .B(n7042), .Z(n7044) );
  XOR U7645 ( .A(n7046), .B(n7047), .Z(n7042) );
  ANDN U7646 ( .B(n6976), .A(n6977), .Z(n7046) );
  AND U7647 ( .A(b[2]), .B(a[43]), .Z(n7048) );
  XNOR U7648 ( .A(n7050), .B(n7047), .Z(n7049) );
  XOR U7649 ( .A(n7051), .B(n7052), .Z(n7047) );
  NANDN U7650 ( .A(n6979), .B(n6978), .Z(n7052) );
  XOR U7651 ( .A(n7051), .B(n7053), .Z(n6978) );
  NAND U7652 ( .A(a[43]), .B(b[1]), .Z(n7053) );
  XOR U7653 ( .A(n7051), .B(n7055), .Z(n7054) );
  OR U7654 ( .A(n2682), .B(n2680), .Z(n7051) );
  XOR U7655 ( .A(n7057), .B(n7058), .Z(n2680) );
  NANDN U7656 ( .A(n179), .B(a[43]), .Z(n2682) );
  XNOR U7657 ( .A(n7024), .B(n7028), .Z(n7062) );
  XNOR U7658 ( .A(n7019), .B(n7023), .Z(n7063) );
  XNOR U7659 ( .A(n7009), .B(n7018), .Z(n7064) );
  XOR U7660 ( .A(n7065), .B(n7008), .Z(n7009) );
  AND U7661 ( .A(b[9]), .B(a[39]), .Z(n7065) );
  XNOR U7662 ( .A(n7008), .B(n7014), .Z(n7066) );
  XNOR U7663 ( .A(n7013), .B(n7005), .Z(n7067) );
  XOR U7664 ( .A(n7004), .B(n7001), .Z(n7068) );
  XOR U7665 ( .A(n7069), .B(n7070), .Z(n7001) );
  XOR U7666 ( .A(n6999), .B(n7071), .Z(n7070) );
  XOR U7667 ( .A(n7072), .B(n7073), .Z(n7071) );
  XOR U7668 ( .A(n7074), .B(n7075), .Z(n7073) );
  NAND U7669 ( .A(a[34]), .B(b[14]), .Z(n7075) );
  AND U7670 ( .A(a[33]), .B(b[15]), .Z(n7074) );
  XOR U7671 ( .A(n7076), .B(n7072), .Z(n7069) );
  XOR U7672 ( .A(n7077), .B(n7078), .Z(n7072) );
  NOR U7673 ( .A(n7079), .B(n7080), .Z(n7077) );
  AND U7674 ( .A(a[35]), .B(b[13]), .Z(n7076) );
  XNOR U7675 ( .A(n7081), .B(n6999), .Z(n7000) );
  XOR U7676 ( .A(n7082), .B(n7083), .Z(n6999) );
  ANDN U7677 ( .B(n7084), .A(n7085), .Z(n7082) );
  AND U7678 ( .A(a[36]), .B(b[12]), .Z(n7081) );
  XNOR U7679 ( .A(n7086), .B(n7004), .Z(n7006) );
  XOR U7680 ( .A(n7087), .B(n7088), .Z(n7004) );
  ANDN U7681 ( .B(n7089), .A(n7090), .Z(n7087) );
  AND U7682 ( .A(a[37]), .B(b[11]), .Z(n7086) );
  XOR U7683 ( .A(n7091), .B(n7092), .Z(n7008) );
  ANDN U7684 ( .B(n7093), .A(n7094), .Z(n7091) );
  XNOR U7685 ( .A(n7095), .B(n7013), .Z(n7015) );
  XOR U7686 ( .A(n7096), .B(n7097), .Z(n7013) );
  ANDN U7687 ( .B(n7098), .A(n7099), .Z(n7096) );
  AND U7688 ( .A(a[38]), .B(b[10]), .Z(n7095) );
  XOR U7689 ( .A(n7101), .B(n7102), .Z(n7018) );
  ANDN U7690 ( .B(n7103), .A(n7104), .Z(n7101) );
  AND U7691 ( .A(a[40]), .B(b[8]), .Z(n7100) );
  XOR U7692 ( .A(n7106), .B(n7107), .Z(n7023) );
  ANDN U7693 ( .B(n7108), .A(n7109), .Z(n7106) );
  AND U7694 ( .A(a[41]), .B(b[7]), .Z(n7105) );
  XOR U7695 ( .A(n7111), .B(n7112), .Z(n7028) );
  ANDN U7696 ( .B(n7040), .A(n7061), .Z(n7111) );
  AND U7697 ( .A(a[42]), .B(b[5]), .Z(n7113) );
  XNOR U7698 ( .A(n7108), .B(n7112), .Z(n7114) );
  XOR U7699 ( .A(n7115), .B(n7116), .Z(n7112) );
  ANDN U7700 ( .B(n7045), .A(n7060), .Z(n7115) );
  AND U7701 ( .A(a[42]), .B(b[4]), .Z(n7117) );
  XNOR U7702 ( .A(n7119), .B(n7116), .Z(n7118) );
  XOR U7703 ( .A(n7120), .B(n7121), .Z(n7116) );
  ANDN U7704 ( .B(n7050), .A(n7059), .Z(n7120) );
  AND U7705 ( .A(a[42]), .B(b[3]), .Z(n7122) );
  XNOR U7706 ( .A(n7124), .B(n7121), .Z(n7123) );
  XOR U7707 ( .A(n7125), .B(n7126), .Z(n7121) );
  ANDN U7708 ( .B(n7055), .A(n7056), .Z(n7125) );
  AND U7709 ( .A(b[2]), .B(a[42]), .Z(n7127) );
  XNOR U7710 ( .A(n7129), .B(n7126), .Z(n7128) );
  XOR U7711 ( .A(n7130), .B(n7131), .Z(n7126) );
  NANDN U7712 ( .A(n7058), .B(n7057), .Z(n7131) );
  XOR U7713 ( .A(n7130), .B(n7132), .Z(n7057) );
  NAND U7714 ( .A(a[42]), .B(b[1]), .Z(n7132) );
  XOR U7715 ( .A(n7130), .B(n7134), .Z(n7133) );
  OR U7716 ( .A(n2687), .B(n2685), .Z(n7130) );
  XOR U7717 ( .A(n7136), .B(n7137), .Z(n2685) );
  NANDN U7718 ( .A(n179), .B(a[42]), .Z(n2687) );
  XNOR U7719 ( .A(n7103), .B(n7107), .Z(n7141) );
  XNOR U7720 ( .A(n7093), .B(n7102), .Z(n7142) );
  XOR U7721 ( .A(n7143), .B(n7092), .Z(n7093) );
  AND U7722 ( .A(b[8]), .B(a[39]), .Z(n7143) );
  XNOR U7723 ( .A(n7092), .B(n7098), .Z(n7144) );
  XNOR U7724 ( .A(n7097), .B(n7089), .Z(n7145) );
  XNOR U7725 ( .A(n7088), .B(n7084), .Z(n7146) );
  XOR U7726 ( .A(n7083), .B(n7080), .Z(n7147) );
  XOR U7727 ( .A(n7148), .B(n7149), .Z(n7080) );
  XOR U7728 ( .A(n7078), .B(n7150), .Z(n7149) );
  XOR U7729 ( .A(n7151), .B(n7152), .Z(n7150) );
  XOR U7730 ( .A(n7153), .B(n7154), .Z(n7152) );
  NAND U7731 ( .A(a[33]), .B(b[14]), .Z(n7154) );
  AND U7732 ( .A(a[32]), .B(b[15]), .Z(n7153) );
  XOR U7733 ( .A(n7155), .B(n7151), .Z(n7148) );
  XOR U7734 ( .A(n7156), .B(n7157), .Z(n7151) );
  NOR U7735 ( .A(n7158), .B(n7159), .Z(n7156) );
  AND U7736 ( .A(a[34]), .B(b[13]), .Z(n7155) );
  XNOR U7737 ( .A(n7160), .B(n7078), .Z(n7079) );
  XOR U7738 ( .A(n7161), .B(n7162), .Z(n7078) );
  ANDN U7739 ( .B(n7163), .A(n7164), .Z(n7161) );
  AND U7740 ( .A(a[35]), .B(b[12]), .Z(n7160) );
  XNOR U7741 ( .A(n7165), .B(n7083), .Z(n7085) );
  XOR U7742 ( .A(n7166), .B(n7167), .Z(n7083) );
  ANDN U7743 ( .B(n7168), .A(n7169), .Z(n7166) );
  AND U7744 ( .A(a[36]), .B(b[11]), .Z(n7165) );
  XNOR U7745 ( .A(n7170), .B(n7088), .Z(n7090) );
  XOR U7746 ( .A(n7171), .B(n7172), .Z(n7088) );
  ANDN U7747 ( .B(n7173), .A(n7174), .Z(n7171) );
  AND U7748 ( .A(a[37]), .B(b[10]), .Z(n7170) );
  XOR U7749 ( .A(n7175), .B(n7176), .Z(n7092) );
  ANDN U7750 ( .B(n7177), .A(n7178), .Z(n7175) );
  XNOR U7751 ( .A(n7179), .B(n7097), .Z(n7099) );
  XOR U7752 ( .A(n7180), .B(n7181), .Z(n7097) );
  ANDN U7753 ( .B(n7182), .A(n7183), .Z(n7180) );
  AND U7754 ( .A(a[38]), .B(b[9]), .Z(n7179) );
  XOR U7755 ( .A(n7185), .B(n7186), .Z(n7102) );
  ANDN U7756 ( .B(n7187), .A(n7188), .Z(n7185) );
  AND U7757 ( .A(a[40]), .B(b[7]), .Z(n7184) );
  XOR U7758 ( .A(n7190), .B(n7191), .Z(n7107) );
  ANDN U7759 ( .B(n7119), .A(n7140), .Z(n7190) );
  AND U7760 ( .A(a[41]), .B(b[5]), .Z(n7192) );
  XNOR U7761 ( .A(n7187), .B(n7191), .Z(n7193) );
  XOR U7762 ( .A(n7194), .B(n7195), .Z(n7191) );
  ANDN U7763 ( .B(n7124), .A(n7139), .Z(n7194) );
  AND U7764 ( .A(a[41]), .B(b[4]), .Z(n7196) );
  XNOR U7765 ( .A(n7198), .B(n7195), .Z(n7197) );
  XOR U7766 ( .A(n7199), .B(n7200), .Z(n7195) );
  ANDN U7767 ( .B(n7129), .A(n7138), .Z(n7199) );
  AND U7768 ( .A(a[41]), .B(b[3]), .Z(n7201) );
  XNOR U7769 ( .A(n7203), .B(n7200), .Z(n7202) );
  XOR U7770 ( .A(n7204), .B(n7205), .Z(n7200) );
  ANDN U7771 ( .B(n7134), .A(n7135), .Z(n7204) );
  AND U7772 ( .A(b[2]), .B(a[41]), .Z(n7206) );
  XNOR U7773 ( .A(n7208), .B(n7205), .Z(n7207) );
  XOR U7774 ( .A(n7209), .B(n7210), .Z(n7205) );
  NANDN U7775 ( .A(n7137), .B(n7136), .Z(n7210) );
  XOR U7776 ( .A(n7209), .B(n7211), .Z(n7136) );
  NAND U7777 ( .A(a[41]), .B(b[1]), .Z(n7211) );
  XOR U7778 ( .A(n7209), .B(n7213), .Z(n7212) );
  OR U7779 ( .A(n2692), .B(n2690), .Z(n7209) );
  XOR U7780 ( .A(n7215), .B(n7216), .Z(n2690) );
  NANDN U7781 ( .A(n179), .B(a[41]), .Z(n2692) );
  XNOR U7782 ( .A(n7177), .B(n7186), .Z(n7220) );
  XOR U7783 ( .A(n7221), .B(n7176), .Z(n7177) );
  AND U7784 ( .A(b[7]), .B(a[39]), .Z(n7221) );
  XNOR U7785 ( .A(n7176), .B(n7182), .Z(n7222) );
  XNOR U7786 ( .A(n7181), .B(n7173), .Z(n7223) );
  XNOR U7787 ( .A(n7172), .B(n7168), .Z(n7224) );
  XNOR U7788 ( .A(n7167), .B(n7163), .Z(n7225) );
  XOR U7789 ( .A(n7162), .B(n7159), .Z(n7226) );
  XOR U7790 ( .A(n7227), .B(n7228), .Z(n7159) );
  XOR U7791 ( .A(n7157), .B(n7229), .Z(n7228) );
  XOR U7792 ( .A(n7230), .B(n7231), .Z(n7229) );
  XOR U7793 ( .A(n7232), .B(n7233), .Z(n7231) );
  NAND U7794 ( .A(a[32]), .B(b[14]), .Z(n7233) );
  AND U7795 ( .A(a[31]), .B(b[15]), .Z(n7232) );
  XOR U7796 ( .A(n7234), .B(n7230), .Z(n7227) );
  XOR U7797 ( .A(n7235), .B(n7236), .Z(n7230) );
  NOR U7798 ( .A(n7237), .B(n7238), .Z(n7235) );
  AND U7799 ( .A(a[33]), .B(b[13]), .Z(n7234) );
  XNOR U7800 ( .A(n7239), .B(n7157), .Z(n7158) );
  XOR U7801 ( .A(n7240), .B(n7241), .Z(n7157) );
  ANDN U7802 ( .B(n7242), .A(n7243), .Z(n7240) );
  AND U7803 ( .A(a[34]), .B(b[12]), .Z(n7239) );
  XNOR U7804 ( .A(n7244), .B(n7162), .Z(n7164) );
  XOR U7805 ( .A(n7245), .B(n7246), .Z(n7162) );
  ANDN U7806 ( .B(n7247), .A(n7248), .Z(n7245) );
  AND U7807 ( .A(a[35]), .B(b[11]), .Z(n7244) );
  XNOR U7808 ( .A(n7249), .B(n7167), .Z(n7169) );
  XOR U7809 ( .A(n7250), .B(n7251), .Z(n7167) );
  ANDN U7810 ( .B(n7252), .A(n7253), .Z(n7250) );
  AND U7811 ( .A(a[36]), .B(b[10]), .Z(n7249) );
  XNOR U7812 ( .A(n7254), .B(n7172), .Z(n7174) );
  XOR U7813 ( .A(n7255), .B(n7256), .Z(n7172) );
  ANDN U7814 ( .B(n7257), .A(n7258), .Z(n7255) );
  AND U7815 ( .A(a[37]), .B(b[9]), .Z(n7254) );
  XOR U7816 ( .A(n7259), .B(n7260), .Z(n7176) );
  ANDN U7817 ( .B(n7261), .A(n7262), .Z(n7259) );
  XNOR U7818 ( .A(n7263), .B(n7181), .Z(n7183) );
  XOR U7819 ( .A(n7264), .B(n7265), .Z(n7181) );
  ANDN U7820 ( .B(n7266), .A(n7267), .Z(n7264) );
  AND U7821 ( .A(a[38]), .B(b[8]), .Z(n7263) );
  XOR U7822 ( .A(n7269), .B(n7270), .Z(n7186) );
  ANDN U7823 ( .B(n7198), .A(n7219), .Z(n7269) );
  AND U7824 ( .A(a[40]), .B(b[5]), .Z(n7271) );
  XNOR U7825 ( .A(n7261), .B(n7270), .Z(n7272) );
  XOR U7826 ( .A(n7273), .B(n7274), .Z(n7270) );
  ANDN U7827 ( .B(n7203), .A(n7218), .Z(n7273) );
  AND U7828 ( .A(a[40]), .B(b[4]), .Z(n7275) );
  XNOR U7829 ( .A(n7277), .B(n7274), .Z(n7276) );
  XOR U7830 ( .A(n7278), .B(n7279), .Z(n7274) );
  ANDN U7831 ( .B(n7208), .A(n7217), .Z(n7278) );
  AND U7832 ( .A(a[40]), .B(b[3]), .Z(n7280) );
  XNOR U7833 ( .A(n7282), .B(n7279), .Z(n7281) );
  XOR U7834 ( .A(n7283), .B(n7284), .Z(n7279) );
  ANDN U7835 ( .B(n7213), .A(n7214), .Z(n7283) );
  AND U7836 ( .A(b[2]), .B(a[40]), .Z(n7285) );
  XNOR U7837 ( .A(n7287), .B(n7284), .Z(n7286) );
  XOR U7838 ( .A(n7288), .B(n7289), .Z(n7284) );
  NANDN U7839 ( .A(n7216), .B(n7215), .Z(n7289) );
  XOR U7840 ( .A(n7288), .B(n7290), .Z(n7215) );
  NAND U7841 ( .A(a[40]), .B(b[1]), .Z(n7290) );
  XNOR U7842 ( .A(n7288), .B(n7292), .Z(n7291) );
  OR U7843 ( .A(n2697), .B(n2695), .Z(n7288) );
  NANDN U7844 ( .A(n179), .B(a[40]), .Z(n2697) );
  XOR U7845 ( .A(n7299), .B(n7260), .Z(n7261) );
  AND U7846 ( .A(b[6]), .B(a[39]), .Z(n7299) );
  XNOR U7847 ( .A(n7260), .B(n7266), .Z(n7300) );
  XNOR U7848 ( .A(n7265), .B(n7257), .Z(n7301) );
  XNOR U7849 ( .A(n7256), .B(n7252), .Z(n7302) );
  XNOR U7850 ( .A(n7251), .B(n7247), .Z(n7303) );
  XNOR U7851 ( .A(n7246), .B(n7242), .Z(n7304) );
  XOR U7852 ( .A(n7241), .B(n7238), .Z(n7305) );
  XOR U7853 ( .A(n7306), .B(n7307), .Z(n7238) );
  XOR U7854 ( .A(n7236), .B(n7308), .Z(n7307) );
  XOR U7855 ( .A(n7309), .B(n7310), .Z(n7308) );
  XOR U7856 ( .A(n7311), .B(n7312), .Z(n7310) );
  NAND U7857 ( .A(a[31]), .B(b[14]), .Z(n7312) );
  AND U7858 ( .A(a[30]), .B(b[15]), .Z(n7311) );
  XOR U7859 ( .A(n7313), .B(n7309), .Z(n7306) );
  XOR U7860 ( .A(n7314), .B(n7315), .Z(n7309) );
  NOR U7861 ( .A(n7316), .B(n7317), .Z(n7314) );
  AND U7862 ( .A(a[32]), .B(b[13]), .Z(n7313) );
  XNOR U7863 ( .A(n7318), .B(n7236), .Z(n7237) );
  XOR U7864 ( .A(n7319), .B(n7320), .Z(n7236) );
  ANDN U7865 ( .B(n7321), .A(n7322), .Z(n7319) );
  AND U7866 ( .A(a[33]), .B(b[12]), .Z(n7318) );
  XNOR U7867 ( .A(n7323), .B(n7241), .Z(n7243) );
  XOR U7868 ( .A(n7324), .B(n7325), .Z(n7241) );
  ANDN U7869 ( .B(n7326), .A(n7327), .Z(n7324) );
  AND U7870 ( .A(a[34]), .B(b[11]), .Z(n7323) );
  XNOR U7871 ( .A(n7328), .B(n7246), .Z(n7248) );
  XOR U7872 ( .A(n7329), .B(n7330), .Z(n7246) );
  ANDN U7873 ( .B(n7331), .A(n7332), .Z(n7329) );
  AND U7874 ( .A(a[35]), .B(b[10]), .Z(n7328) );
  XNOR U7875 ( .A(n7333), .B(n7251), .Z(n7253) );
  XOR U7876 ( .A(n7334), .B(n7335), .Z(n7251) );
  ANDN U7877 ( .B(n7336), .A(n7337), .Z(n7334) );
  AND U7878 ( .A(a[36]), .B(b[9]), .Z(n7333) );
  XNOR U7879 ( .A(n7338), .B(n7256), .Z(n7258) );
  XOR U7880 ( .A(n7339), .B(n7340), .Z(n7256) );
  ANDN U7881 ( .B(n7341), .A(n7342), .Z(n7339) );
  AND U7882 ( .A(a[37]), .B(b[8]), .Z(n7338) );
  XOR U7883 ( .A(n7343), .B(n7344), .Z(n7260) );
  ANDN U7884 ( .B(n7277), .A(n7298), .Z(n7343) );
  XNOR U7885 ( .A(n7344), .B(n7346), .Z(n7345) );
  XOR U7886 ( .A(n7348), .B(n7344), .Z(n7277) );
  XOR U7887 ( .A(n7349), .B(n7350), .Z(n7344) );
  ANDN U7888 ( .B(n7282), .A(n7297), .Z(n7349) );
  XNOR U7889 ( .A(n7350), .B(n7352), .Z(n7351) );
  XOR U7890 ( .A(n7354), .B(n7350), .Z(n7282) );
  XOR U7891 ( .A(n7355), .B(n7356), .Z(n7350) );
  ANDN U7892 ( .B(n7287), .A(n7296), .Z(n7355) );
  XNOR U7893 ( .A(n7356), .B(n7358), .Z(n7357) );
  XOR U7894 ( .A(n7360), .B(n7356), .Z(n7287) );
  XNOR U7895 ( .A(n7361), .B(n7362), .Z(n7356) );
  NOR U7896 ( .A(n7293), .B(n7292), .Z(n7361) );
  XOR U7897 ( .A(n7363), .B(n7362), .Z(n7292) );
  AND U7898 ( .A(b[2]), .B(a[39]), .Z(n7363) );
  XOR U7899 ( .A(n7362), .B(n7365), .Z(n7364) );
  XNOR U7900 ( .A(n7366), .B(n7367), .Z(n7362) );
  OR U7901 ( .A(n7294), .B(n7295), .Z(n7367) );
  XNOR U7902 ( .A(n7366), .B(n7369), .Z(n7368) );
  XNOR U7903 ( .A(n7366), .B(n7371), .Z(n7294) );
  NAND U7904 ( .A(b[1]), .B(a[39]), .Z(n7371) );
  OR U7905 ( .A(n2702), .B(n2700), .Z(n7366) );
  XOR U7906 ( .A(n7372), .B(n7373), .Z(n2700) );
  NANDN U7907 ( .A(n179), .B(a[39]), .Z(n2702) );
  AND U7908 ( .A(b[3]), .B(a[39]), .Z(n7360) );
  AND U7909 ( .A(b[4]), .B(a[39]), .Z(n7354) );
  AND U7910 ( .A(b[5]), .B(a[39]), .Z(n7348) );
  XNOR U7911 ( .A(n7375), .B(n7265), .Z(n7267) );
  XOR U7912 ( .A(n7376), .B(n7377), .Z(n7265) );
  ANDN U7913 ( .B(n7346), .A(n7347), .Z(n7376) );
  XNOR U7914 ( .A(n7378), .B(n7377), .Z(n7347) );
  AND U7915 ( .A(a[38]), .B(b[6]), .Z(n7378) );
  XNOR U7916 ( .A(n7377), .B(n7341), .Z(n7379) );
  XNOR U7917 ( .A(n7340), .B(n7336), .Z(n7380) );
  XNOR U7918 ( .A(n7335), .B(n7331), .Z(n7381) );
  XNOR U7919 ( .A(n7330), .B(n7326), .Z(n7382) );
  XNOR U7920 ( .A(n7325), .B(n7321), .Z(n7383) );
  XOR U7921 ( .A(n7320), .B(n7317), .Z(n7384) );
  XOR U7922 ( .A(n7385), .B(n7386), .Z(n7317) );
  XOR U7923 ( .A(n7315), .B(n7387), .Z(n7386) );
  XOR U7924 ( .A(n7388), .B(n7389), .Z(n7387) );
  XOR U7925 ( .A(n7390), .B(n7391), .Z(n7389) );
  NAND U7926 ( .A(a[30]), .B(b[14]), .Z(n7391) );
  AND U7927 ( .A(a[29]), .B(b[15]), .Z(n7390) );
  XOR U7928 ( .A(n7392), .B(n7388), .Z(n7385) );
  XOR U7929 ( .A(n7393), .B(n7394), .Z(n7388) );
  NOR U7930 ( .A(n7395), .B(n7396), .Z(n7393) );
  AND U7931 ( .A(a[31]), .B(b[13]), .Z(n7392) );
  XNOR U7932 ( .A(n7397), .B(n7315), .Z(n7316) );
  XOR U7933 ( .A(n7398), .B(n7399), .Z(n7315) );
  ANDN U7934 ( .B(n7400), .A(n7401), .Z(n7398) );
  AND U7935 ( .A(a[32]), .B(b[12]), .Z(n7397) );
  XNOR U7936 ( .A(n7402), .B(n7320), .Z(n7322) );
  XOR U7937 ( .A(n7403), .B(n7404), .Z(n7320) );
  ANDN U7938 ( .B(n7405), .A(n7406), .Z(n7403) );
  AND U7939 ( .A(a[33]), .B(b[11]), .Z(n7402) );
  XNOR U7940 ( .A(n7407), .B(n7325), .Z(n7327) );
  XOR U7941 ( .A(n7408), .B(n7409), .Z(n7325) );
  ANDN U7942 ( .B(n7410), .A(n7411), .Z(n7408) );
  AND U7943 ( .A(a[34]), .B(b[10]), .Z(n7407) );
  XNOR U7944 ( .A(n7412), .B(n7330), .Z(n7332) );
  XOR U7945 ( .A(n7413), .B(n7414), .Z(n7330) );
  ANDN U7946 ( .B(n7415), .A(n7416), .Z(n7413) );
  AND U7947 ( .A(a[35]), .B(b[9]), .Z(n7412) );
  XNOR U7948 ( .A(n7417), .B(n7335), .Z(n7337) );
  XOR U7949 ( .A(n7418), .B(n7419), .Z(n7335) );
  ANDN U7950 ( .B(n7420), .A(n7421), .Z(n7418) );
  AND U7951 ( .A(a[36]), .B(b[8]), .Z(n7417) );
  XOR U7952 ( .A(n7422), .B(n7423), .Z(n7377) );
  ANDN U7953 ( .B(n7352), .A(n7353), .Z(n7422) );
  XNOR U7954 ( .A(n7424), .B(n7423), .Z(n7353) );
  AND U7955 ( .A(a[38]), .B(b[5]), .Z(n7424) );
  XNOR U7956 ( .A(n7423), .B(n7426), .Z(n7425) );
  XOR U7957 ( .A(n7427), .B(n7428), .Z(n7423) );
  ANDN U7958 ( .B(n7358), .A(n7359), .Z(n7427) );
  XNOR U7959 ( .A(n7429), .B(n7428), .Z(n7359) );
  AND U7960 ( .A(a[38]), .B(b[4]), .Z(n7429) );
  XNOR U7961 ( .A(n7428), .B(n7431), .Z(n7430) );
  XOR U7962 ( .A(n7432), .B(n7433), .Z(n7428) );
  ANDN U7963 ( .B(n7365), .A(n7374), .Z(n7432) );
  XNOR U7964 ( .A(n7434), .B(n7433), .Z(n7374) );
  AND U7965 ( .A(a[38]), .B(b[3]), .Z(n7434) );
  XNOR U7966 ( .A(n7433), .B(n7436), .Z(n7435) );
  XNOR U7967 ( .A(n7437), .B(n7438), .Z(n7433) );
  NOR U7968 ( .A(n7370), .B(n7369), .Z(n7437) );
  XOR U7969 ( .A(n7439), .B(n7438), .Z(n7369) );
  AND U7970 ( .A(b[2]), .B(a[38]), .Z(n7439) );
  XOR U7971 ( .A(n7438), .B(n7441), .Z(n7440) );
  XNOR U7972 ( .A(n7442), .B(n7443), .Z(n7438) );
  NANDN U7973 ( .A(n7373), .B(n7372), .Z(n7443) );
  XOR U7974 ( .A(n7442), .B(n7444), .Z(n7372) );
  NAND U7975 ( .A(a[38]), .B(b[1]), .Z(n7444) );
  XOR U7976 ( .A(n7442), .B(n7446), .Z(n7445) );
  OR U7977 ( .A(n2707), .B(n2705), .Z(n7442) );
  XOR U7978 ( .A(n7448), .B(n7449), .Z(n2705) );
  NANDN U7979 ( .A(n179), .B(a[38]), .Z(n2707) );
  XNOR U7980 ( .A(n7454), .B(n7340), .Z(n7342) );
  XOR U7981 ( .A(n7455), .B(n7456), .Z(n7340) );
  ANDN U7982 ( .B(n7426), .A(n7453), .Z(n7455) );
  XNOR U7983 ( .A(n7457), .B(n7456), .Z(n7453) );
  AND U7984 ( .A(a[37]), .B(b[6]), .Z(n7457) );
  XNOR U7985 ( .A(n7456), .B(n7420), .Z(n7458) );
  XNOR U7986 ( .A(n7419), .B(n7415), .Z(n7459) );
  XNOR U7987 ( .A(n7414), .B(n7410), .Z(n7460) );
  XNOR U7988 ( .A(n7409), .B(n7405), .Z(n7461) );
  XNOR U7989 ( .A(n7404), .B(n7400), .Z(n7462) );
  XOR U7990 ( .A(n7399), .B(n7396), .Z(n7463) );
  XOR U7991 ( .A(n7464), .B(n7465), .Z(n7396) );
  XOR U7992 ( .A(n7394), .B(n7466), .Z(n7465) );
  XOR U7993 ( .A(n7467), .B(n7468), .Z(n7466) );
  XOR U7994 ( .A(n7469), .B(n7470), .Z(n7468) );
  NAND U7995 ( .A(a[29]), .B(b[14]), .Z(n7470) );
  AND U7996 ( .A(a[28]), .B(b[15]), .Z(n7469) );
  XOR U7997 ( .A(n7471), .B(n7467), .Z(n7464) );
  XOR U7998 ( .A(n7472), .B(n7473), .Z(n7467) );
  NOR U7999 ( .A(n7474), .B(n7475), .Z(n7472) );
  AND U8000 ( .A(a[30]), .B(b[13]), .Z(n7471) );
  XNOR U8001 ( .A(n7476), .B(n7394), .Z(n7395) );
  XOR U8002 ( .A(n7477), .B(n7478), .Z(n7394) );
  ANDN U8003 ( .B(n7479), .A(n7480), .Z(n7477) );
  AND U8004 ( .A(a[31]), .B(b[12]), .Z(n7476) );
  XNOR U8005 ( .A(n7481), .B(n7399), .Z(n7401) );
  XOR U8006 ( .A(n7482), .B(n7483), .Z(n7399) );
  ANDN U8007 ( .B(n7484), .A(n7485), .Z(n7482) );
  AND U8008 ( .A(a[32]), .B(b[11]), .Z(n7481) );
  XNOR U8009 ( .A(n7486), .B(n7404), .Z(n7406) );
  XOR U8010 ( .A(n7487), .B(n7488), .Z(n7404) );
  ANDN U8011 ( .B(n7489), .A(n7490), .Z(n7487) );
  AND U8012 ( .A(a[33]), .B(b[10]), .Z(n7486) );
  XNOR U8013 ( .A(n7491), .B(n7409), .Z(n7411) );
  XOR U8014 ( .A(n7492), .B(n7493), .Z(n7409) );
  ANDN U8015 ( .B(n7494), .A(n7495), .Z(n7492) );
  AND U8016 ( .A(a[34]), .B(b[9]), .Z(n7491) );
  XNOR U8017 ( .A(n7496), .B(n7414), .Z(n7416) );
  XOR U8018 ( .A(n7497), .B(n7498), .Z(n7414) );
  ANDN U8019 ( .B(n7499), .A(n7500), .Z(n7497) );
  AND U8020 ( .A(a[35]), .B(b[8]), .Z(n7496) );
  XOR U8021 ( .A(n7501), .B(n7502), .Z(n7456) );
  ANDN U8022 ( .B(n7431), .A(n7452), .Z(n7501) );
  XNOR U8023 ( .A(n7503), .B(n7502), .Z(n7452) );
  AND U8024 ( .A(a[37]), .B(b[5]), .Z(n7503) );
  XNOR U8025 ( .A(n7502), .B(n7505), .Z(n7504) );
  XOR U8026 ( .A(n7506), .B(n7507), .Z(n7502) );
  ANDN U8027 ( .B(n7436), .A(n7451), .Z(n7506) );
  XNOR U8028 ( .A(n7508), .B(n7507), .Z(n7451) );
  AND U8029 ( .A(a[37]), .B(b[4]), .Z(n7508) );
  XNOR U8030 ( .A(n7507), .B(n7510), .Z(n7509) );
  XOR U8031 ( .A(n7511), .B(n7512), .Z(n7507) );
  ANDN U8032 ( .B(n7441), .A(n7450), .Z(n7511) );
  XNOR U8033 ( .A(n7513), .B(n7512), .Z(n7450) );
  AND U8034 ( .A(a[37]), .B(b[3]), .Z(n7513) );
  XNOR U8035 ( .A(n7512), .B(n7515), .Z(n7514) );
  XNOR U8036 ( .A(n7516), .B(n7517), .Z(n7512) );
  ANDN U8037 ( .B(n7446), .A(n7447), .Z(n7516) );
  XOR U8038 ( .A(n7518), .B(n7517), .Z(n7447) );
  IV U8039 ( .A(n7519), .Z(n7517) );
  AND U8040 ( .A(b[2]), .B(a[37]), .Z(n7518) );
  XNOR U8041 ( .A(n7521), .B(n7519), .Z(n7520) );
  XOR U8042 ( .A(n7522), .B(n7523), .Z(n7519) );
  NANDN U8043 ( .A(n7449), .B(n7448), .Z(n7523) );
  XOR U8044 ( .A(n7522), .B(n7524), .Z(n7448) );
  NAND U8045 ( .A(a[37]), .B(b[1]), .Z(n7524) );
  XOR U8046 ( .A(n7522), .B(n7526), .Z(n7525) );
  OR U8047 ( .A(n2712), .B(n2710), .Z(n7522) );
  XOR U8048 ( .A(n7528), .B(n7529), .Z(n2710) );
  NANDN U8049 ( .A(n179), .B(a[37]), .Z(n2712) );
  XNOR U8050 ( .A(n7534), .B(n7419), .Z(n7421) );
  XOR U8051 ( .A(n7535), .B(n7536), .Z(n7419) );
  ANDN U8052 ( .B(n7505), .A(n7533), .Z(n7535) );
  XNOR U8053 ( .A(n7537), .B(n7536), .Z(n7533) );
  AND U8054 ( .A(a[36]), .B(b[6]), .Z(n7537) );
  XNOR U8055 ( .A(n7536), .B(n7499), .Z(n7538) );
  XNOR U8056 ( .A(n7498), .B(n7494), .Z(n7539) );
  XNOR U8057 ( .A(n7493), .B(n7489), .Z(n7540) );
  XNOR U8058 ( .A(n7488), .B(n7484), .Z(n7541) );
  XNOR U8059 ( .A(n7483), .B(n7479), .Z(n7542) );
  XOR U8060 ( .A(n7478), .B(n7475), .Z(n7543) );
  XOR U8061 ( .A(n7544), .B(n7545), .Z(n7475) );
  XOR U8062 ( .A(n7473), .B(n7546), .Z(n7545) );
  XOR U8063 ( .A(n7547), .B(n7548), .Z(n7546) );
  XOR U8064 ( .A(n7549), .B(n7550), .Z(n7548) );
  NAND U8065 ( .A(a[28]), .B(b[14]), .Z(n7550) );
  AND U8066 ( .A(a[27]), .B(b[15]), .Z(n7549) );
  XOR U8067 ( .A(n7551), .B(n7547), .Z(n7544) );
  XOR U8068 ( .A(n7552), .B(n7553), .Z(n7547) );
  NOR U8069 ( .A(n7554), .B(n7555), .Z(n7552) );
  AND U8070 ( .A(a[29]), .B(b[13]), .Z(n7551) );
  XNOR U8071 ( .A(n7556), .B(n7473), .Z(n7474) );
  XOR U8072 ( .A(n7557), .B(n7558), .Z(n7473) );
  ANDN U8073 ( .B(n7559), .A(n7560), .Z(n7557) );
  AND U8074 ( .A(a[30]), .B(b[12]), .Z(n7556) );
  XNOR U8075 ( .A(n7561), .B(n7478), .Z(n7480) );
  XOR U8076 ( .A(n7562), .B(n7563), .Z(n7478) );
  ANDN U8077 ( .B(n7564), .A(n7565), .Z(n7562) );
  AND U8078 ( .A(a[31]), .B(b[11]), .Z(n7561) );
  XNOR U8079 ( .A(n7566), .B(n7483), .Z(n7485) );
  XOR U8080 ( .A(n7567), .B(n7568), .Z(n7483) );
  ANDN U8081 ( .B(n7569), .A(n7570), .Z(n7567) );
  AND U8082 ( .A(a[32]), .B(b[10]), .Z(n7566) );
  XNOR U8083 ( .A(n7571), .B(n7488), .Z(n7490) );
  XOR U8084 ( .A(n7572), .B(n7573), .Z(n7488) );
  ANDN U8085 ( .B(n7574), .A(n7575), .Z(n7572) );
  AND U8086 ( .A(a[33]), .B(b[9]), .Z(n7571) );
  XNOR U8087 ( .A(n7576), .B(n7493), .Z(n7495) );
  XOR U8088 ( .A(n7577), .B(n7578), .Z(n7493) );
  ANDN U8089 ( .B(n7579), .A(n7580), .Z(n7577) );
  AND U8090 ( .A(a[34]), .B(b[8]), .Z(n7576) );
  XOR U8091 ( .A(n7581), .B(n7582), .Z(n7536) );
  ANDN U8092 ( .B(n7510), .A(n7532), .Z(n7581) );
  XNOR U8093 ( .A(n7583), .B(n7582), .Z(n7532) );
  AND U8094 ( .A(a[36]), .B(b[5]), .Z(n7583) );
  XNOR U8095 ( .A(n7582), .B(n7585), .Z(n7584) );
  XOR U8096 ( .A(n7586), .B(n7587), .Z(n7582) );
  ANDN U8097 ( .B(n7515), .A(n7531), .Z(n7586) );
  XNOR U8098 ( .A(n7588), .B(n7587), .Z(n7531) );
  AND U8099 ( .A(a[36]), .B(b[4]), .Z(n7588) );
  XNOR U8100 ( .A(n7587), .B(n7590), .Z(n7589) );
  XNOR U8101 ( .A(n7591), .B(n7592), .Z(n7587) );
  ANDN U8102 ( .B(n7521), .A(n7530), .Z(n7591) );
  XOR U8103 ( .A(n7593), .B(n7592), .Z(n7530) );
  IV U8104 ( .A(n7594), .Z(n7592) );
  AND U8105 ( .A(a[36]), .B(b[3]), .Z(n7593) );
  XNOR U8106 ( .A(n7596), .B(n7594), .Z(n7595) );
  XOR U8107 ( .A(n7597), .B(n7598), .Z(n7594) );
  ANDN U8108 ( .B(n7526), .A(n7527), .Z(n7597) );
  AND U8109 ( .A(b[2]), .B(a[36]), .Z(n7599) );
  XNOR U8110 ( .A(n7601), .B(n7598), .Z(n7600) );
  XOR U8111 ( .A(n7602), .B(n7603), .Z(n7598) );
  NANDN U8112 ( .A(n7529), .B(n7528), .Z(n7603) );
  XOR U8113 ( .A(n7602), .B(n7604), .Z(n7528) );
  NAND U8114 ( .A(a[36]), .B(b[1]), .Z(n7604) );
  XOR U8115 ( .A(n7602), .B(n7606), .Z(n7605) );
  OR U8116 ( .A(n2717), .B(n2715), .Z(n7602) );
  XOR U8117 ( .A(n7608), .B(n7609), .Z(n2715) );
  NANDN U8118 ( .A(n179), .B(a[36]), .Z(n2717) );
  XNOR U8119 ( .A(n7614), .B(n7498), .Z(n7500) );
  XOR U8120 ( .A(n7615), .B(n7616), .Z(n7498) );
  ANDN U8121 ( .B(n7585), .A(n7613), .Z(n7615) );
  XNOR U8122 ( .A(n7617), .B(n7616), .Z(n7613) );
  AND U8123 ( .A(a[35]), .B(b[6]), .Z(n7617) );
  XNOR U8124 ( .A(n7616), .B(n7579), .Z(n7618) );
  XNOR U8125 ( .A(n7578), .B(n7574), .Z(n7619) );
  XNOR U8126 ( .A(n7573), .B(n7569), .Z(n7620) );
  XNOR U8127 ( .A(n7568), .B(n7564), .Z(n7621) );
  XNOR U8128 ( .A(n7563), .B(n7559), .Z(n7622) );
  XOR U8129 ( .A(n7558), .B(n7555), .Z(n7623) );
  XOR U8130 ( .A(n7624), .B(n7625), .Z(n7555) );
  XOR U8131 ( .A(n7553), .B(n7626), .Z(n7625) );
  XOR U8132 ( .A(n7627), .B(n7628), .Z(n7626) );
  XOR U8133 ( .A(n7629), .B(n7630), .Z(n7628) );
  NAND U8134 ( .A(a[27]), .B(b[14]), .Z(n7630) );
  AND U8135 ( .A(a[26]), .B(b[15]), .Z(n7629) );
  XOR U8136 ( .A(n7631), .B(n7627), .Z(n7624) );
  XOR U8137 ( .A(n7632), .B(n7633), .Z(n7627) );
  NOR U8138 ( .A(n7634), .B(n7635), .Z(n7632) );
  AND U8139 ( .A(a[28]), .B(b[13]), .Z(n7631) );
  XNOR U8140 ( .A(n7636), .B(n7553), .Z(n7554) );
  XOR U8141 ( .A(n7637), .B(n7638), .Z(n7553) );
  ANDN U8142 ( .B(n7639), .A(n7640), .Z(n7637) );
  AND U8143 ( .A(a[29]), .B(b[12]), .Z(n7636) );
  XNOR U8144 ( .A(n7641), .B(n7558), .Z(n7560) );
  XOR U8145 ( .A(n7642), .B(n7643), .Z(n7558) );
  ANDN U8146 ( .B(n7644), .A(n7645), .Z(n7642) );
  AND U8147 ( .A(a[30]), .B(b[11]), .Z(n7641) );
  XNOR U8148 ( .A(n7646), .B(n7563), .Z(n7565) );
  XOR U8149 ( .A(n7647), .B(n7648), .Z(n7563) );
  ANDN U8150 ( .B(n7649), .A(n7650), .Z(n7647) );
  AND U8151 ( .A(a[31]), .B(b[10]), .Z(n7646) );
  XNOR U8152 ( .A(n7651), .B(n7568), .Z(n7570) );
  XOR U8153 ( .A(n7652), .B(n7653), .Z(n7568) );
  ANDN U8154 ( .B(n7654), .A(n7655), .Z(n7652) );
  AND U8155 ( .A(a[32]), .B(b[9]), .Z(n7651) );
  XNOR U8156 ( .A(n7656), .B(n7573), .Z(n7575) );
  XOR U8157 ( .A(n7657), .B(n7658), .Z(n7573) );
  ANDN U8158 ( .B(n7659), .A(n7660), .Z(n7657) );
  AND U8159 ( .A(a[33]), .B(b[8]), .Z(n7656) );
  XOR U8160 ( .A(n7661), .B(n7662), .Z(n7616) );
  ANDN U8161 ( .B(n7590), .A(n7612), .Z(n7661) );
  XNOR U8162 ( .A(n7663), .B(n7662), .Z(n7612) );
  AND U8163 ( .A(a[35]), .B(b[5]), .Z(n7663) );
  XNOR U8164 ( .A(n7662), .B(n7665), .Z(n7664) );
  XNOR U8165 ( .A(n7666), .B(n7667), .Z(n7662) );
  ANDN U8166 ( .B(n7596), .A(n7611), .Z(n7666) );
  XOR U8167 ( .A(n7668), .B(n7667), .Z(n7611) );
  IV U8168 ( .A(n7669), .Z(n7667) );
  AND U8169 ( .A(a[35]), .B(b[4]), .Z(n7668) );
  XNOR U8170 ( .A(n7671), .B(n7669), .Z(n7670) );
  XOR U8171 ( .A(n7672), .B(n7673), .Z(n7669) );
  ANDN U8172 ( .B(n7601), .A(n7610), .Z(n7672) );
  AND U8173 ( .A(a[35]), .B(b[3]), .Z(n7674) );
  XNOR U8174 ( .A(n7676), .B(n7673), .Z(n7675) );
  XOR U8175 ( .A(n7677), .B(n7678), .Z(n7673) );
  ANDN U8176 ( .B(n7606), .A(n7607), .Z(n7677) );
  AND U8177 ( .A(b[2]), .B(a[35]), .Z(n7679) );
  XNOR U8178 ( .A(n7681), .B(n7678), .Z(n7680) );
  XOR U8179 ( .A(n7682), .B(n7683), .Z(n7678) );
  NANDN U8180 ( .A(n7609), .B(n7608), .Z(n7683) );
  XOR U8181 ( .A(n7682), .B(n7684), .Z(n7608) );
  NAND U8182 ( .A(a[35]), .B(b[1]), .Z(n7684) );
  XOR U8183 ( .A(n7682), .B(n7686), .Z(n7685) );
  OR U8184 ( .A(n2722), .B(n2720), .Z(n7682) );
  XOR U8185 ( .A(n7688), .B(n7689), .Z(n2720) );
  NANDN U8186 ( .A(n179), .B(a[35]), .Z(n2722) );
  XNOR U8187 ( .A(n7694), .B(n7578), .Z(n7580) );
  XOR U8188 ( .A(n7695), .B(n7696), .Z(n7578) );
  ANDN U8189 ( .B(n7665), .A(n7693), .Z(n7695) );
  XNOR U8190 ( .A(n7697), .B(n7696), .Z(n7693) );
  AND U8191 ( .A(a[34]), .B(b[6]), .Z(n7697) );
  XNOR U8192 ( .A(n7696), .B(n7659), .Z(n7698) );
  XNOR U8193 ( .A(n7658), .B(n7654), .Z(n7699) );
  XNOR U8194 ( .A(n7653), .B(n7649), .Z(n7700) );
  XNOR U8195 ( .A(n7648), .B(n7644), .Z(n7701) );
  XNOR U8196 ( .A(n7643), .B(n7639), .Z(n7702) );
  XOR U8197 ( .A(n7638), .B(n7635), .Z(n7703) );
  XOR U8198 ( .A(n7704), .B(n7705), .Z(n7635) );
  XOR U8199 ( .A(n7633), .B(n7706), .Z(n7705) );
  XNOR U8200 ( .A(n7707), .B(n7708), .Z(n7706) );
  XOR U8201 ( .A(n7709), .B(n7710), .Z(n7708) );
  NAND U8202 ( .A(a[26]), .B(b[14]), .Z(n7710) );
  AND U8203 ( .A(a[25]), .B(b[15]), .Z(n7709) );
  XNOR U8204 ( .A(n7711), .B(n7707), .Z(n7704) );
  XOR U8205 ( .A(n7712), .B(n7713), .Z(n7707) );
  NOR U8206 ( .A(n7714), .B(n7715), .Z(n7712) );
  AND U8207 ( .A(a[27]), .B(b[13]), .Z(n7711) );
  XNOR U8208 ( .A(n7716), .B(n7633), .Z(n7634) );
  XNOR U8209 ( .A(n7717), .B(n7718), .Z(n7633) );
  ANDN U8210 ( .B(n7719), .A(n7720), .Z(n7717) );
  AND U8211 ( .A(a[28]), .B(b[12]), .Z(n7716) );
  XNOR U8212 ( .A(n7721), .B(n7638), .Z(n7640) );
  XNOR U8213 ( .A(n7722), .B(n7723), .Z(n7638) );
  ANDN U8214 ( .B(n7724), .A(n7725), .Z(n7722) );
  AND U8215 ( .A(a[29]), .B(b[11]), .Z(n7721) );
  XNOR U8216 ( .A(n7726), .B(n7643), .Z(n7645) );
  XNOR U8217 ( .A(n7727), .B(n7728), .Z(n7643) );
  ANDN U8218 ( .B(n7729), .A(n7730), .Z(n7727) );
  AND U8219 ( .A(a[30]), .B(b[10]), .Z(n7726) );
  XNOR U8220 ( .A(n7731), .B(n7648), .Z(n7650) );
  XNOR U8221 ( .A(n7732), .B(n7733), .Z(n7648) );
  ANDN U8222 ( .B(n7734), .A(n7735), .Z(n7732) );
  AND U8223 ( .A(a[31]), .B(b[9]), .Z(n7731) );
  XNOR U8224 ( .A(n7736), .B(n7653), .Z(n7655) );
  XNOR U8225 ( .A(n7737), .B(n7738), .Z(n7653) );
  ANDN U8226 ( .B(n7739), .A(n7740), .Z(n7737) );
  AND U8227 ( .A(a[32]), .B(b[8]), .Z(n7736) );
  XNOR U8228 ( .A(n7741), .B(n7742), .Z(n7696) );
  ANDN U8229 ( .B(n7671), .A(n7692), .Z(n7741) );
  XOR U8230 ( .A(n7743), .B(n7742), .Z(n7692) );
  IV U8231 ( .A(n7744), .Z(n7742) );
  AND U8232 ( .A(a[34]), .B(b[5]), .Z(n7743) );
  XNOR U8233 ( .A(n7746), .B(n7744), .Z(n7745) );
  XOR U8234 ( .A(n7747), .B(n7748), .Z(n7744) );
  ANDN U8235 ( .B(n7676), .A(n7691), .Z(n7747) );
  AND U8236 ( .A(a[34]), .B(b[4]), .Z(n7749) );
  XNOR U8237 ( .A(n7751), .B(n7748), .Z(n7750) );
  XOR U8238 ( .A(n7752), .B(n7753), .Z(n7748) );
  ANDN U8239 ( .B(n7681), .A(n7690), .Z(n7752) );
  AND U8240 ( .A(a[34]), .B(b[3]), .Z(n7754) );
  XNOR U8241 ( .A(n7756), .B(n7753), .Z(n7755) );
  XOR U8242 ( .A(n7757), .B(n7758), .Z(n7753) );
  ANDN U8243 ( .B(n7686), .A(n7687), .Z(n7757) );
  AND U8244 ( .A(b[2]), .B(a[34]), .Z(n7759) );
  XNOR U8245 ( .A(n7761), .B(n7758), .Z(n7760) );
  XOR U8246 ( .A(n7762), .B(n7763), .Z(n7758) );
  NANDN U8247 ( .A(n7689), .B(n7688), .Z(n7763) );
  XOR U8248 ( .A(n7762), .B(n7764), .Z(n7688) );
  NAND U8249 ( .A(a[34]), .B(b[1]), .Z(n7764) );
  XOR U8250 ( .A(n7762), .B(n7766), .Z(n7765) );
  OR U8251 ( .A(n2727), .B(n2725), .Z(n7762) );
  XOR U8252 ( .A(n7768), .B(n7769), .Z(n2725) );
  NANDN U8253 ( .A(n179), .B(a[34]), .Z(n2727) );
  XNOR U8254 ( .A(n7774), .B(n7658), .Z(n7660) );
  XNOR U8255 ( .A(n7775), .B(n7776), .Z(n7658) );
  ANDN U8256 ( .B(n7746), .A(n7773), .Z(n7775) );
  XOR U8257 ( .A(n7777), .B(n7776), .Z(n7773) );
  IV U8258 ( .A(n7778), .Z(n7776) );
  AND U8259 ( .A(a[33]), .B(b[6]), .Z(n7777) );
  XNOR U8260 ( .A(n7739), .B(n7778), .Z(n7779) );
  XOR U8261 ( .A(n7780), .B(n7781), .Z(n7778) );
  ANDN U8262 ( .B(n7751), .A(n7772), .Z(n7780) );
  AND U8263 ( .A(a[33]), .B(b[5]), .Z(n7782) );
  XNOR U8264 ( .A(n7784), .B(n7781), .Z(n7783) );
  XOR U8265 ( .A(n7785), .B(n7786), .Z(n7781) );
  ANDN U8266 ( .B(n7756), .A(n7771), .Z(n7785) );
  AND U8267 ( .A(a[33]), .B(b[4]), .Z(n7787) );
  XNOR U8268 ( .A(n7789), .B(n7786), .Z(n7788) );
  XOR U8269 ( .A(n7790), .B(n7791), .Z(n7786) );
  ANDN U8270 ( .B(n7761), .A(n7770), .Z(n7790) );
  AND U8271 ( .A(a[33]), .B(b[3]), .Z(n7792) );
  XNOR U8272 ( .A(n7794), .B(n7791), .Z(n7793) );
  XOR U8273 ( .A(n7795), .B(n7796), .Z(n7791) );
  ANDN U8274 ( .B(n7766), .A(n7767), .Z(n7795) );
  AND U8275 ( .A(b[2]), .B(a[33]), .Z(n7797) );
  XNOR U8276 ( .A(n7799), .B(n7796), .Z(n7798) );
  XOR U8277 ( .A(n7800), .B(n7801), .Z(n7796) );
  NANDN U8278 ( .A(n7769), .B(n7768), .Z(n7801) );
  XOR U8279 ( .A(n7800), .B(n7802), .Z(n7768) );
  NAND U8280 ( .A(a[33]), .B(b[1]), .Z(n7802) );
  XOR U8281 ( .A(n7800), .B(n7804), .Z(n7803) );
  OR U8282 ( .A(n2732), .B(n2730), .Z(n7800) );
  XOR U8283 ( .A(n7806), .B(n7807), .Z(n2730) );
  NANDN U8284 ( .A(n179), .B(a[33]), .Z(n2732) );
  XNOR U8285 ( .A(n7734), .B(n7813), .Z(n7812) );
  XNOR U8286 ( .A(n7729), .B(n7815), .Z(n7814) );
  XNOR U8287 ( .A(n7724), .B(n7817), .Z(n7816) );
  XNOR U8288 ( .A(n7719), .B(n7819), .Z(n7818) );
  XOR U8289 ( .A(n7715), .B(n7821), .Z(n7820) );
  XOR U8290 ( .A(n7822), .B(n7823), .Z(n7715) );
  XNOR U8291 ( .A(n7824), .B(n7825), .Z(n7823) );
  XNOR U8292 ( .A(n7826), .B(n7827), .Z(n7824) );
  XOR U8293 ( .A(n7828), .B(n7829), .Z(n7827) );
  AND U8294 ( .A(b[15]), .B(a[24]), .Z(n7829) );
  AND U8295 ( .A(a[25]), .B(b[14]), .Z(n7828) );
  XNOR U8296 ( .A(n7830), .B(n7826), .Z(n7822) );
  XOR U8297 ( .A(n7831), .B(n7832), .Z(n7826) );
  NOR U8298 ( .A(n7833), .B(n7834), .Z(n7831) );
  AND U8299 ( .A(a[26]), .B(b[13]), .Z(n7830) );
  XOR U8300 ( .A(n7835), .B(n7713), .Z(n7714) );
  IV U8301 ( .A(n7825), .Z(n7713) );
  XOR U8302 ( .A(n7836), .B(n7837), .Z(n7825) );
  ANDN U8303 ( .B(n7838), .A(n7839), .Z(n7836) );
  AND U8304 ( .A(a[27]), .B(b[12]), .Z(n7835) );
  XOR U8305 ( .A(n7840), .B(n7718), .Z(n7720) );
  IV U8306 ( .A(n7821), .Z(n7718) );
  XOR U8307 ( .A(n7841), .B(n7842), .Z(n7821) );
  ANDN U8308 ( .B(n7843), .A(n7844), .Z(n7841) );
  AND U8309 ( .A(a[28]), .B(b[11]), .Z(n7840) );
  XOR U8310 ( .A(n7845), .B(n7723), .Z(n7725) );
  IV U8311 ( .A(n7819), .Z(n7723) );
  XOR U8312 ( .A(n7846), .B(n7847), .Z(n7819) );
  ANDN U8313 ( .B(n7848), .A(n7849), .Z(n7846) );
  AND U8314 ( .A(a[29]), .B(b[10]), .Z(n7845) );
  XOR U8315 ( .A(n7850), .B(n7728), .Z(n7730) );
  IV U8316 ( .A(n7817), .Z(n7728) );
  XOR U8317 ( .A(n7851), .B(n7852), .Z(n7817) );
  ANDN U8318 ( .B(n7853), .A(n7854), .Z(n7851) );
  AND U8319 ( .A(a[30]), .B(b[9]), .Z(n7850) );
  XOR U8320 ( .A(n7855), .B(n7733), .Z(n7735) );
  IV U8321 ( .A(n7815), .Z(n7733) );
  XOR U8322 ( .A(n7856), .B(n7857), .Z(n7815) );
  ANDN U8323 ( .B(n7858), .A(n7859), .Z(n7856) );
  AND U8324 ( .A(a[31]), .B(b[8]), .Z(n7855) );
  XOR U8325 ( .A(n7860), .B(n7738), .Z(n7740) );
  IV U8326 ( .A(n7813), .Z(n7738) );
  XOR U8327 ( .A(n7861), .B(n7862), .Z(n7813) );
  ANDN U8328 ( .B(n7784), .A(n7811), .Z(n7861) );
  AND U8329 ( .A(a[32]), .B(b[6]), .Z(n7863) );
  XNOR U8330 ( .A(n7858), .B(n7862), .Z(n7864) );
  XOR U8331 ( .A(n7865), .B(n7866), .Z(n7862) );
  ANDN U8332 ( .B(n7789), .A(n7810), .Z(n7865) );
  AND U8333 ( .A(a[32]), .B(b[5]), .Z(n7867) );
  XNOR U8334 ( .A(n7869), .B(n7866), .Z(n7868) );
  XOR U8335 ( .A(n7870), .B(n7871), .Z(n7866) );
  ANDN U8336 ( .B(n7794), .A(n7809), .Z(n7870) );
  AND U8337 ( .A(a[32]), .B(b[4]), .Z(n7872) );
  XNOR U8338 ( .A(n7874), .B(n7871), .Z(n7873) );
  XOR U8339 ( .A(n7875), .B(n7876), .Z(n7871) );
  ANDN U8340 ( .B(n7799), .A(n7808), .Z(n7875) );
  AND U8341 ( .A(a[32]), .B(b[3]), .Z(n7877) );
  XNOR U8342 ( .A(n7879), .B(n7876), .Z(n7878) );
  XOR U8343 ( .A(n7880), .B(n7881), .Z(n7876) );
  ANDN U8344 ( .B(n7804), .A(n7805), .Z(n7880) );
  AND U8345 ( .A(b[2]), .B(a[32]), .Z(n7882) );
  XNOR U8346 ( .A(n7884), .B(n7881), .Z(n7883) );
  XOR U8347 ( .A(n7885), .B(n7886), .Z(n7881) );
  NANDN U8348 ( .A(n7807), .B(n7806), .Z(n7886) );
  XOR U8349 ( .A(n7885), .B(n7887), .Z(n7806) );
  NAND U8350 ( .A(a[32]), .B(b[1]), .Z(n7887) );
  XOR U8351 ( .A(n7885), .B(n7889), .Z(n7888) );
  OR U8352 ( .A(n2737), .B(n2735), .Z(n7885) );
  XOR U8353 ( .A(n7891), .B(n7892), .Z(n2735) );
  NANDN U8354 ( .A(n179), .B(a[32]), .Z(n2737) );
  XNOR U8355 ( .A(n7853), .B(n7857), .Z(n7897) );
  XNOR U8356 ( .A(n7848), .B(n7852), .Z(n7898) );
  XNOR U8357 ( .A(n7843), .B(n7847), .Z(n7899) );
  XNOR U8358 ( .A(n7838), .B(n7842), .Z(n7900) );
  XOR U8359 ( .A(n7834), .B(n7837), .Z(n7901) );
  XOR U8360 ( .A(n7902), .B(n7903), .Z(n7834) );
  XNOR U8361 ( .A(n7904), .B(n7905), .Z(n7903) );
  XNOR U8362 ( .A(n7906), .B(n7907), .Z(n7904) );
  XOR U8363 ( .A(n7908), .B(n7909), .Z(n7907) );
  AND U8364 ( .A(b[14]), .B(a[24]), .Z(n7909) );
  AND U8365 ( .A(a[23]), .B(b[15]), .Z(n7908) );
  XNOR U8366 ( .A(n7910), .B(n7906), .Z(n7902) );
  XOR U8367 ( .A(n7911), .B(n7912), .Z(n7906) );
  NOR U8368 ( .A(n7913), .B(n7914), .Z(n7911) );
  AND U8369 ( .A(a[25]), .B(b[13]), .Z(n7910) );
  XOR U8370 ( .A(n7915), .B(n7832), .Z(n7833) );
  IV U8371 ( .A(n7905), .Z(n7832) );
  XOR U8372 ( .A(n7916), .B(n7917), .Z(n7905) );
  ANDN U8373 ( .B(n7918), .A(n7919), .Z(n7916) );
  AND U8374 ( .A(a[26]), .B(b[12]), .Z(n7915) );
  XOR U8375 ( .A(n7921), .B(n7922), .Z(n7837) );
  ANDN U8376 ( .B(n7923), .A(n7924), .Z(n7921) );
  AND U8377 ( .A(a[27]), .B(b[11]), .Z(n7920) );
  XOR U8378 ( .A(n7926), .B(n7927), .Z(n7842) );
  ANDN U8379 ( .B(n7928), .A(n7929), .Z(n7926) );
  AND U8380 ( .A(a[28]), .B(b[10]), .Z(n7925) );
  XOR U8381 ( .A(n7931), .B(n7932), .Z(n7847) );
  ANDN U8382 ( .B(n7933), .A(n7934), .Z(n7931) );
  AND U8383 ( .A(a[29]), .B(b[9]), .Z(n7930) );
  XOR U8384 ( .A(n7936), .B(n7937), .Z(n7852) );
  ANDN U8385 ( .B(n7938), .A(n7939), .Z(n7936) );
  AND U8386 ( .A(a[30]), .B(b[8]), .Z(n7935) );
  XOR U8387 ( .A(n7941), .B(n7942), .Z(n7857) );
  ANDN U8388 ( .B(n7869), .A(n7896), .Z(n7941) );
  AND U8389 ( .A(a[31]), .B(b[6]), .Z(n7943) );
  XNOR U8390 ( .A(n7938), .B(n7942), .Z(n7944) );
  XOR U8391 ( .A(n7945), .B(n7946), .Z(n7942) );
  ANDN U8392 ( .B(n7874), .A(n7895), .Z(n7945) );
  AND U8393 ( .A(a[31]), .B(b[5]), .Z(n7947) );
  XNOR U8394 ( .A(n7949), .B(n7946), .Z(n7948) );
  XOR U8395 ( .A(n7950), .B(n7951), .Z(n7946) );
  ANDN U8396 ( .B(n7879), .A(n7894), .Z(n7950) );
  AND U8397 ( .A(a[31]), .B(b[4]), .Z(n7952) );
  XNOR U8398 ( .A(n7954), .B(n7951), .Z(n7953) );
  XOR U8399 ( .A(n7955), .B(n7956), .Z(n7951) );
  ANDN U8400 ( .B(n7884), .A(n7893), .Z(n7955) );
  AND U8401 ( .A(a[31]), .B(b[3]), .Z(n7957) );
  XNOR U8402 ( .A(n7959), .B(n7956), .Z(n7958) );
  XOR U8403 ( .A(n7960), .B(n7961), .Z(n7956) );
  ANDN U8404 ( .B(n7889), .A(n7890), .Z(n7960) );
  AND U8405 ( .A(b[2]), .B(a[31]), .Z(n7962) );
  XNOR U8406 ( .A(n7964), .B(n7961), .Z(n7963) );
  XOR U8407 ( .A(n7965), .B(n7966), .Z(n7961) );
  NANDN U8408 ( .A(n7892), .B(n7891), .Z(n7966) );
  XOR U8409 ( .A(n7965), .B(n7967), .Z(n7891) );
  NAND U8410 ( .A(a[31]), .B(b[1]), .Z(n7967) );
  XOR U8411 ( .A(n7965), .B(n7969), .Z(n7968) );
  OR U8412 ( .A(n2742), .B(n2740), .Z(n7965) );
  XOR U8413 ( .A(n7971), .B(n7972), .Z(n2740) );
  NANDN U8414 ( .A(n179), .B(a[31]), .Z(n2742) );
  XNOR U8415 ( .A(n7933), .B(n7937), .Z(n7977) );
  XNOR U8416 ( .A(n7928), .B(n7932), .Z(n7978) );
  XNOR U8417 ( .A(n7923), .B(n7927), .Z(n7979) );
  XNOR U8418 ( .A(n7918), .B(n7922), .Z(n7980) );
  XOR U8419 ( .A(n7914), .B(n7917), .Z(n7981) );
  XOR U8420 ( .A(n7982), .B(n7983), .Z(n7914) );
  XNOR U8421 ( .A(n7984), .B(n7985), .Z(n7983) );
  XOR U8422 ( .A(n7986), .B(n7987), .Z(n7984) );
  AND U8423 ( .A(b[13]), .B(a[24]), .Z(n7986) );
  XOR U8424 ( .A(n7987), .B(n7988), .Z(n7982) );
  XOR U8425 ( .A(n7989), .B(n7990), .Z(n7988) );
  AND U8426 ( .A(a[23]), .B(b[14]), .Z(n7990) );
  AND U8427 ( .A(a[22]), .B(b[15]), .Z(n7989) );
  XOR U8428 ( .A(n7991), .B(n7992), .Z(n7987) );
  ANDN U8429 ( .B(n7993), .A(n7994), .Z(n7991) );
  XOR U8430 ( .A(n7995), .B(n7912), .Z(n7913) );
  IV U8431 ( .A(n7985), .Z(n7912) );
  XOR U8432 ( .A(n7996), .B(n7997), .Z(n7985) );
  NOR U8433 ( .A(n7998), .B(n7999), .Z(n7996) );
  AND U8434 ( .A(a[25]), .B(b[12]), .Z(n7995) );
  XOR U8435 ( .A(n8001), .B(n8002), .Z(n7917) );
  ANDN U8436 ( .B(n8003), .A(n8004), .Z(n8001) );
  AND U8437 ( .A(a[26]), .B(b[11]), .Z(n8000) );
  XOR U8438 ( .A(n8006), .B(n8007), .Z(n7922) );
  ANDN U8439 ( .B(n8008), .A(n8009), .Z(n8006) );
  AND U8440 ( .A(a[27]), .B(b[10]), .Z(n8005) );
  XOR U8441 ( .A(n8011), .B(n8012), .Z(n7927) );
  ANDN U8442 ( .B(n8013), .A(n8014), .Z(n8011) );
  AND U8443 ( .A(a[28]), .B(b[9]), .Z(n8010) );
  XOR U8444 ( .A(n8016), .B(n8017), .Z(n7932) );
  ANDN U8445 ( .B(n8018), .A(n8019), .Z(n8016) );
  AND U8446 ( .A(a[29]), .B(b[8]), .Z(n8015) );
  XOR U8447 ( .A(n8021), .B(n8022), .Z(n7937) );
  ANDN U8448 ( .B(n7949), .A(n7976), .Z(n8021) );
  AND U8449 ( .A(a[30]), .B(b[6]), .Z(n8023) );
  XNOR U8450 ( .A(n8018), .B(n8022), .Z(n8024) );
  XOR U8451 ( .A(n8025), .B(n8026), .Z(n8022) );
  ANDN U8452 ( .B(n7954), .A(n7975), .Z(n8025) );
  AND U8453 ( .A(a[30]), .B(b[5]), .Z(n8027) );
  XNOR U8454 ( .A(n8029), .B(n8026), .Z(n8028) );
  XOR U8455 ( .A(n8030), .B(n8031), .Z(n8026) );
  ANDN U8456 ( .B(n7959), .A(n7974), .Z(n8030) );
  AND U8457 ( .A(a[30]), .B(b[4]), .Z(n8032) );
  XNOR U8458 ( .A(n8034), .B(n8031), .Z(n8033) );
  XOR U8459 ( .A(n8035), .B(n8036), .Z(n8031) );
  ANDN U8460 ( .B(n7964), .A(n7973), .Z(n8035) );
  AND U8461 ( .A(a[30]), .B(b[3]), .Z(n8037) );
  XNOR U8462 ( .A(n8039), .B(n8036), .Z(n8038) );
  XOR U8463 ( .A(n8040), .B(n8041), .Z(n8036) );
  ANDN U8464 ( .B(n7969), .A(n7970), .Z(n8040) );
  AND U8465 ( .A(b[2]), .B(a[30]), .Z(n8042) );
  XNOR U8466 ( .A(n8044), .B(n8041), .Z(n8043) );
  XOR U8467 ( .A(n8045), .B(n8046), .Z(n8041) );
  NANDN U8468 ( .A(n7972), .B(n7971), .Z(n8046) );
  XOR U8469 ( .A(n8045), .B(n8047), .Z(n7971) );
  NAND U8470 ( .A(a[30]), .B(b[1]), .Z(n8047) );
  XOR U8471 ( .A(n8045), .B(n8049), .Z(n8048) );
  OR U8472 ( .A(n2747), .B(n2745), .Z(n8045) );
  XOR U8473 ( .A(n8051), .B(n8052), .Z(n2745) );
  NANDN U8474 ( .A(n179), .B(a[30]), .Z(n2747) );
  XNOR U8475 ( .A(n8013), .B(n8017), .Z(n8057) );
  XNOR U8476 ( .A(n8008), .B(n8012), .Z(n8058) );
  XNOR U8477 ( .A(n8003), .B(n8007), .Z(n8059) );
  XOR U8478 ( .A(n7999), .B(n8002), .Z(n8060) );
  XNOR U8479 ( .A(n7994), .B(n8061), .Z(n7999) );
  XNOR U8480 ( .A(n7993), .B(n7997), .Z(n8061) );
  XOR U8481 ( .A(n8062), .B(n7992), .Z(n7993) );
  AND U8482 ( .A(b[12]), .B(a[24]), .Z(n8062) );
  XOR U8483 ( .A(n8063), .B(n8064), .Z(n7994) );
  XOR U8484 ( .A(n7992), .B(n8065), .Z(n8064) );
  XOR U8485 ( .A(n8066), .B(n8067), .Z(n8065) );
  XOR U8486 ( .A(n8068), .B(n8069), .Z(n8067) );
  NAND U8487 ( .A(a[22]), .B(b[14]), .Z(n8069) );
  AND U8488 ( .A(a[21]), .B(b[15]), .Z(n8068) );
  XOR U8489 ( .A(n8070), .B(n8071), .Z(n7992) );
  ANDN U8490 ( .B(n8072), .A(n8073), .Z(n8070) );
  XOR U8491 ( .A(n8074), .B(n8066), .Z(n8063) );
  XOR U8492 ( .A(n8075), .B(n8076), .Z(n8066) );
  NOR U8493 ( .A(n8077), .B(n8078), .Z(n8075) );
  AND U8494 ( .A(a[23]), .B(b[13]), .Z(n8074) );
  XOR U8495 ( .A(n8080), .B(n8081), .Z(n7997) );
  ANDN U8496 ( .B(n8082), .A(n8083), .Z(n8080) );
  AND U8497 ( .A(a[25]), .B(b[11]), .Z(n8079) );
  XOR U8498 ( .A(n8085), .B(n8086), .Z(n8002) );
  ANDN U8499 ( .B(n8087), .A(n8088), .Z(n8085) );
  AND U8500 ( .A(a[26]), .B(b[10]), .Z(n8084) );
  XOR U8501 ( .A(n8090), .B(n8091), .Z(n8007) );
  ANDN U8502 ( .B(n8092), .A(n8093), .Z(n8090) );
  AND U8503 ( .A(a[27]), .B(b[9]), .Z(n8089) );
  XOR U8504 ( .A(n8095), .B(n8096), .Z(n8012) );
  ANDN U8505 ( .B(n8097), .A(n8098), .Z(n8095) );
  AND U8506 ( .A(a[28]), .B(b[8]), .Z(n8094) );
  XOR U8507 ( .A(n8100), .B(n8101), .Z(n8017) );
  ANDN U8508 ( .B(n8029), .A(n8056), .Z(n8100) );
  AND U8509 ( .A(a[29]), .B(b[6]), .Z(n8102) );
  XNOR U8510 ( .A(n8097), .B(n8101), .Z(n8103) );
  XOR U8511 ( .A(n8104), .B(n8105), .Z(n8101) );
  ANDN U8512 ( .B(n8034), .A(n8055), .Z(n8104) );
  AND U8513 ( .A(a[29]), .B(b[5]), .Z(n8106) );
  XNOR U8514 ( .A(n8108), .B(n8105), .Z(n8107) );
  XOR U8515 ( .A(n8109), .B(n8110), .Z(n8105) );
  ANDN U8516 ( .B(n8039), .A(n8054), .Z(n8109) );
  AND U8517 ( .A(a[29]), .B(b[4]), .Z(n8111) );
  XNOR U8518 ( .A(n8113), .B(n8110), .Z(n8112) );
  XOR U8519 ( .A(n8114), .B(n8115), .Z(n8110) );
  ANDN U8520 ( .B(n8044), .A(n8053), .Z(n8114) );
  AND U8521 ( .A(a[29]), .B(b[3]), .Z(n8116) );
  XNOR U8522 ( .A(n8118), .B(n8115), .Z(n8117) );
  XOR U8523 ( .A(n8119), .B(n8120), .Z(n8115) );
  ANDN U8524 ( .B(n8049), .A(n8050), .Z(n8119) );
  AND U8525 ( .A(b[2]), .B(a[29]), .Z(n8121) );
  XNOR U8526 ( .A(n8123), .B(n8120), .Z(n8122) );
  XOR U8527 ( .A(n8124), .B(n8125), .Z(n8120) );
  NANDN U8528 ( .A(n8052), .B(n8051), .Z(n8125) );
  XOR U8529 ( .A(n8124), .B(n8126), .Z(n8051) );
  NAND U8530 ( .A(a[29]), .B(b[1]), .Z(n8126) );
  XOR U8531 ( .A(n8124), .B(n8128), .Z(n8127) );
  OR U8532 ( .A(n2752), .B(n2750), .Z(n8124) );
  XOR U8533 ( .A(n8130), .B(n8131), .Z(n2750) );
  NANDN U8534 ( .A(n179), .B(a[29]), .Z(n2752) );
  XNOR U8535 ( .A(n8092), .B(n8096), .Z(n8136) );
  XNOR U8536 ( .A(n8087), .B(n8091), .Z(n8137) );
  XNOR U8537 ( .A(n8082), .B(n8086), .Z(n8138) );
  XNOR U8538 ( .A(n8072), .B(n8081), .Z(n8139) );
  XOR U8539 ( .A(n8140), .B(n8071), .Z(n8072) );
  AND U8540 ( .A(b[11]), .B(a[24]), .Z(n8140) );
  XOR U8541 ( .A(n8071), .B(n8078), .Z(n8141) );
  XOR U8542 ( .A(n8142), .B(n8143), .Z(n8078) );
  XOR U8543 ( .A(n8076), .B(n8144), .Z(n8143) );
  XOR U8544 ( .A(n8145), .B(n8146), .Z(n8144) );
  XOR U8545 ( .A(n8147), .B(n8148), .Z(n8146) );
  NAND U8546 ( .A(a[21]), .B(b[14]), .Z(n8148) );
  AND U8547 ( .A(a[20]), .B(b[15]), .Z(n8147) );
  XOR U8548 ( .A(n8149), .B(n8145), .Z(n8142) );
  XOR U8549 ( .A(n8150), .B(n8151), .Z(n8145) );
  NOR U8550 ( .A(n8152), .B(n8153), .Z(n8150) );
  AND U8551 ( .A(a[22]), .B(b[13]), .Z(n8149) );
  XOR U8552 ( .A(n8154), .B(n8155), .Z(n8071) );
  ANDN U8553 ( .B(n8156), .A(n8157), .Z(n8154) );
  XNOR U8554 ( .A(n8158), .B(n8076), .Z(n8077) );
  XOR U8555 ( .A(n8159), .B(n8160), .Z(n8076) );
  ANDN U8556 ( .B(n8161), .A(n8162), .Z(n8159) );
  AND U8557 ( .A(a[23]), .B(b[12]), .Z(n8158) );
  XOR U8558 ( .A(n8164), .B(n8165), .Z(n8081) );
  ANDN U8559 ( .B(n8166), .A(n8167), .Z(n8164) );
  AND U8560 ( .A(a[25]), .B(b[10]), .Z(n8163) );
  XOR U8561 ( .A(n8169), .B(n8170), .Z(n8086) );
  ANDN U8562 ( .B(n8171), .A(n8172), .Z(n8169) );
  AND U8563 ( .A(a[26]), .B(b[9]), .Z(n8168) );
  XOR U8564 ( .A(n8174), .B(n8175), .Z(n8091) );
  ANDN U8565 ( .B(n8176), .A(n8177), .Z(n8174) );
  AND U8566 ( .A(a[27]), .B(b[8]), .Z(n8173) );
  XOR U8567 ( .A(n8179), .B(n8180), .Z(n8096) );
  ANDN U8568 ( .B(n8108), .A(n8135), .Z(n8179) );
  AND U8569 ( .A(a[28]), .B(b[6]), .Z(n8181) );
  XNOR U8570 ( .A(n8176), .B(n8180), .Z(n8182) );
  XOR U8571 ( .A(n8183), .B(n8184), .Z(n8180) );
  ANDN U8572 ( .B(n8113), .A(n8134), .Z(n8183) );
  AND U8573 ( .A(a[28]), .B(b[5]), .Z(n8185) );
  XNOR U8574 ( .A(n8187), .B(n8184), .Z(n8186) );
  XOR U8575 ( .A(n8188), .B(n8189), .Z(n8184) );
  ANDN U8576 ( .B(n8118), .A(n8133), .Z(n8188) );
  AND U8577 ( .A(a[28]), .B(b[4]), .Z(n8190) );
  XNOR U8578 ( .A(n8192), .B(n8189), .Z(n8191) );
  XOR U8579 ( .A(n8193), .B(n8194), .Z(n8189) );
  ANDN U8580 ( .B(n8123), .A(n8132), .Z(n8193) );
  AND U8581 ( .A(a[28]), .B(b[3]), .Z(n8195) );
  XNOR U8582 ( .A(n8197), .B(n8194), .Z(n8196) );
  XOR U8583 ( .A(n8198), .B(n8199), .Z(n8194) );
  ANDN U8584 ( .B(n8128), .A(n8129), .Z(n8198) );
  AND U8585 ( .A(b[2]), .B(a[28]), .Z(n8200) );
  XNOR U8586 ( .A(n8202), .B(n8199), .Z(n8201) );
  XOR U8587 ( .A(n8203), .B(n8204), .Z(n8199) );
  NANDN U8588 ( .A(n8131), .B(n8130), .Z(n8204) );
  XOR U8589 ( .A(n8203), .B(n8205), .Z(n8130) );
  NAND U8590 ( .A(a[28]), .B(b[1]), .Z(n8205) );
  XOR U8591 ( .A(n8203), .B(n8207), .Z(n8206) );
  OR U8592 ( .A(n2757), .B(n2755), .Z(n8203) );
  XOR U8593 ( .A(n8209), .B(n8210), .Z(n2755) );
  NANDN U8594 ( .A(n179), .B(a[28]), .Z(n2757) );
  XNOR U8595 ( .A(n8171), .B(n8175), .Z(n8215) );
  XNOR U8596 ( .A(n8166), .B(n8170), .Z(n8216) );
  XNOR U8597 ( .A(n8156), .B(n8165), .Z(n8217) );
  XOR U8598 ( .A(n8218), .B(n8155), .Z(n8156) );
  AND U8599 ( .A(b[10]), .B(a[24]), .Z(n8218) );
  XNOR U8600 ( .A(n8155), .B(n8161), .Z(n8219) );
  XOR U8601 ( .A(n8160), .B(n8153), .Z(n8220) );
  XOR U8602 ( .A(n8221), .B(n8222), .Z(n8153) );
  XOR U8603 ( .A(n8151), .B(n8223), .Z(n8222) );
  XOR U8604 ( .A(n8224), .B(n8225), .Z(n8223) );
  XOR U8605 ( .A(n8226), .B(n8227), .Z(n8225) );
  NAND U8606 ( .A(a[20]), .B(b[14]), .Z(n8227) );
  AND U8607 ( .A(a[19]), .B(b[15]), .Z(n8226) );
  XOR U8608 ( .A(n8228), .B(n8224), .Z(n8221) );
  XOR U8609 ( .A(n8229), .B(n8230), .Z(n8224) );
  NOR U8610 ( .A(n8231), .B(n8232), .Z(n8229) );
  AND U8611 ( .A(a[21]), .B(b[13]), .Z(n8228) );
  XNOR U8612 ( .A(n8233), .B(n8151), .Z(n8152) );
  XOR U8613 ( .A(n8234), .B(n8235), .Z(n8151) );
  ANDN U8614 ( .B(n8236), .A(n8237), .Z(n8234) );
  AND U8615 ( .A(a[22]), .B(b[12]), .Z(n8233) );
  XOR U8616 ( .A(n8238), .B(n8239), .Z(n8155) );
  ANDN U8617 ( .B(n8240), .A(n8241), .Z(n8238) );
  XNOR U8618 ( .A(n8242), .B(n8160), .Z(n8162) );
  XOR U8619 ( .A(n8243), .B(n8244), .Z(n8160) );
  ANDN U8620 ( .B(n8245), .A(n8246), .Z(n8243) );
  AND U8621 ( .A(a[23]), .B(b[11]), .Z(n8242) );
  XOR U8622 ( .A(n8248), .B(n8249), .Z(n8165) );
  ANDN U8623 ( .B(n8250), .A(n8251), .Z(n8248) );
  AND U8624 ( .A(a[25]), .B(b[9]), .Z(n8247) );
  XOR U8625 ( .A(n8253), .B(n8254), .Z(n8170) );
  ANDN U8626 ( .B(n8255), .A(n8256), .Z(n8253) );
  AND U8627 ( .A(a[26]), .B(b[8]), .Z(n8252) );
  XOR U8628 ( .A(n8258), .B(n8259), .Z(n8175) );
  ANDN U8629 ( .B(n8187), .A(n8214), .Z(n8258) );
  AND U8630 ( .A(a[27]), .B(b[6]), .Z(n8260) );
  XNOR U8631 ( .A(n8255), .B(n8259), .Z(n8261) );
  XOR U8632 ( .A(n8262), .B(n8263), .Z(n8259) );
  ANDN U8633 ( .B(n8192), .A(n8213), .Z(n8262) );
  AND U8634 ( .A(a[27]), .B(b[5]), .Z(n8264) );
  XNOR U8635 ( .A(n8266), .B(n8263), .Z(n8265) );
  XOR U8636 ( .A(n8267), .B(n8268), .Z(n8263) );
  ANDN U8637 ( .B(n8197), .A(n8212), .Z(n8267) );
  AND U8638 ( .A(a[27]), .B(b[4]), .Z(n8269) );
  XNOR U8639 ( .A(n8271), .B(n8268), .Z(n8270) );
  XOR U8640 ( .A(n8272), .B(n8273), .Z(n8268) );
  ANDN U8641 ( .B(n8202), .A(n8211), .Z(n8272) );
  AND U8642 ( .A(a[27]), .B(b[3]), .Z(n8274) );
  XNOR U8643 ( .A(n8276), .B(n8273), .Z(n8275) );
  XOR U8644 ( .A(n8277), .B(n8278), .Z(n8273) );
  ANDN U8645 ( .B(n8207), .A(n8208), .Z(n8277) );
  AND U8646 ( .A(b[2]), .B(a[27]), .Z(n8279) );
  XNOR U8647 ( .A(n8281), .B(n8278), .Z(n8280) );
  XOR U8648 ( .A(n8282), .B(n8283), .Z(n8278) );
  NANDN U8649 ( .A(n8210), .B(n8209), .Z(n8283) );
  XOR U8650 ( .A(n8282), .B(n8284), .Z(n8209) );
  NAND U8651 ( .A(a[27]), .B(b[1]), .Z(n8284) );
  XOR U8652 ( .A(n8282), .B(n8286), .Z(n8285) );
  OR U8653 ( .A(n2762), .B(n2760), .Z(n8282) );
  XOR U8654 ( .A(n8288), .B(n8289), .Z(n2760) );
  NANDN U8655 ( .A(n179), .B(a[27]), .Z(n2762) );
  XNOR U8656 ( .A(n8250), .B(n8254), .Z(n8294) );
  XNOR U8657 ( .A(n8240), .B(n8249), .Z(n8295) );
  XOR U8658 ( .A(n8296), .B(n8239), .Z(n8240) );
  AND U8659 ( .A(b[9]), .B(a[24]), .Z(n8296) );
  XNOR U8660 ( .A(n8239), .B(n8245), .Z(n8297) );
  XNOR U8661 ( .A(n8244), .B(n8236), .Z(n8298) );
  XOR U8662 ( .A(n8235), .B(n8232), .Z(n8299) );
  XOR U8663 ( .A(n8300), .B(n8301), .Z(n8232) );
  XOR U8664 ( .A(n8230), .B(n8302), .Z(n8301) );
  XOR U8665 ( .A(n8303), .B(n8304), .Z(n8302) );
  XOR U8666 ( .A(n8305), .B(n8306), .Z(n8304) );
  NAND U8667 ( .A(a[19]), .B(b[14]), .Z(n8306) );
  AND U8668 ( .A(a[18]), .B(b[15]), .Z(n8305) );
  XOR U8669 ( .A(n8307), .B(n8303), .Z(n8300) );
  XOR U8670 ( .A(n8308), .B(n8309), .Z(n8303) );
  NOR U8671 ( .A(n8310), .B(n8311), .Z(n8308) );
  AND U8672 ( .A(a[20]), .B(b[13]), .Z(n8307) );
  XNOR U8673 ( .A(n8312), .B(n8230), .Z(n8231) );
  XOR U8674 ( .A(n8313), .B(n8314), .Z(n8230) );
  ANDN U8675 ( .B(n8315), .A(n8316), .Z(n8313) );
  AND U8676 ( .A(a[21]), .B(b[12]), .Z(n8312) );
  XNOR U8677 ( .A(n8317), .B(n8235), .Z(n8237) );
  XOR U8678 ( .A(n8318), .B(n8319), .Z(n8235) );
  ANDN U8679 ( .B(n8320), .A(n8321), .Z(n8318) );
  AND U8680 ( .A(a[22]), .B(b[11]), .Z(n8317) );
  XOR U8681 ( .A(n8322), .B(n8323), .Z(n8239) );
  ANDN U8682 ( .B(n8324), .A(n8325), .Z(n8322) );
  XNOR U8683 ( .A(n8326), .B(n8244), .Z(n8246) );
  XOR U8684 ( .A(n8327), .B(n8328), .Z(n8244) );
  ANDN U8685 ( .B(n8329), .A(n8330), .Z(n8327) );
  AND U8686 ( .A(a[23]), .B(b[10]), .Z(n8326) );
  XOR U8687 ( .A(n8332), .B(n8333), .Z(n8249) );
  ANDN U8688 ( .B(n8334), .A(n8335), .Z(n8332) );
  AND U8689 ( .A(a[25]), .B(b[8]), .Z(n8331) );
  XOR U8690 ( .A(n8337), .B(n8338), .Z(n8254) );
  ANDN U8691 ( .B(n8266), .A(n8293), .Z(n8337) );
  AND U8692 ( .A(a[26]), .B(b[6]), .Z(n8339) );
  XNOR U8693 ( .A(n8334), .B(n8338), .Z(n8340) );
  XOR U8694 ( .A(n8341), .B(n8342), .Z(n8338) );
  ANDN U8695 ( .B(n8271), .A(n8292), .Z(n8341) );
  AND U8696 ( .A(a[26]), .B(b[5]), .Z(n8343) );
  XNOR U8697 ( .A(n8345), .B(n8342), .Z(n8344) );
  XOR U8698 ( .A(n8346), .B(n8347), .Z(n8342) );
  ANDN U8699 ( .B(n8276), .A(n8291), .Z(n8346) );
  AND U8700 ( .A(a[26]), .B(b[4]), .Z(n8348) );
  XNOR U8701 ( .A(n8350), .B(n8347), .Z(n8349) );
  XOR U8702 ( .A(n8351), .B(n8352), .Z(n8347) );
  ANDN U8703 ( .B(n8281), .A(n8290), .Z(n8351) );
  AND U8704 ( .A(a[26]), .B(b[3]), .Z(n8353) );
  XNOR U8705 ( .A(n8355), .B(n8352), .Z(n8354) );
  XOR U8706 ( .A(n8356), .B(n8357), .Z(n8352) );
  ANDN U8707 ( .B(n8286), .A(n8287), .Z(n8356) );
  AND U8708 ( .A(b[2]), .B(a[26]), .Z(n8358) );
  XNOR U8709 ( .A(n8360), .B(n8357), .Z(n8359) );
  XOR U8710 ( .A(n8361), .B(n8362), .Z(n8357) );
  NANDN U8711 ( .A(n8289), .B(n8288), .Z(n8362) );
  XOR U8712 ( .A(n8361), .B(n8363), .Z(n8288) );
  NAND U8713 ( .A(a[26]), .B(b[1]), .Z(n8363) );
  XOR U8714 ( .A(n8361), .B(n8365), .Z(n8364) );
  OR U8715 ( .A(n2767), .B(n2765), .Z(n8361) );
  XOR U8716 ( .A(n8367), .B(n8368), .Z(n2765) );
  NANDN U8717 ( .A(n179), .B(a[26]), .Z(n2767) );
  XNOR U8718 ( .A(n8324), .B(n8333), .Z(n8373) );
  XOR U8719 ( .A(n8374), .B(n8323), .Z(n8324) );
  AND U8720 ( .A(b[8]), .B(a[24]), .Z(n8374) );
  XNOR U8721 ( .A(n8323), .B(n8329), .Z(n8375) );
  XNOR U8722 ( .A(n8328), .B(n8320), .Z(n8376) );
  XNOR U8723 ( .A(n8319), .B(n8315), .Z(n8377) );
  XOR U8724 ( .A(n8314), .B(n8311), .Z(n8378) );
  XOR U8725 ( .A(n8379), .B(n8380), .Z(n8311) );
  XOR U8726 ( .A(n8309), .B(n8381), .Z(n8380) );
  XOR U8727 ( .A(n8382), .B(n8383), .Z(n8381) );
  XOR U8728 ( .A(n8384), .B(n8385), .Z(n8383) );
  NAND U8729 ( .A(a[18]), .B(b[14]), .Z(n8385) );
  AND U8730 ( .A(a[17]), .B(b[15]), .Z(n8384) );
  XOR U8731 ( .A(n8386), .B(n8382), .Z(n8379) );
  XOR U8732 ( .A(n8387), .B(n8388), .Z(n8382) );
  NOR U8733 ( .A(n8389), .B(n8390), .Z(n8387) );
  AND U8734 ( .A(a[19]), .B(b[13]), .Z(n8386) );
  XNOR U8735 ( .A(n8391), .B(n8309), .Z(n8310) );
  XOR U8736 ( .A(n8392), .B(n8393), .Z(n8309) );
  ANDN U8737 ( .B(n8394), .A(n8395), .Z(n8392) );
  AND U8738 ( .A(a[20]), .B(b[12]), .Z(n8391) );
  XNOR U8739 ( .A(n8396), .B(n8314), .Z(n8316) );
  XOR U8740 ( .A(n8397), .B(n8398), .Z(n8314) );
  ANDN U8741 ( .B(n8399), .A(n8400), .Z(n8397) );
  AND U8742 ( .A(a[21]), .B(b[11]), .Z(n8396) );
  XNOR U8743 ( .A(n8401), .B(n8319), .Z(n8321) );
  XOR U8744 ( .A(n8402), .B(n8403), .Z(n8319) );
  ANDN U8745 ( .B(n8404), .A(n8405), .Z(n8402) );
  AND U8746 ( .A(a[22]), .B(b[10]), .Z(n8401) );
  XOR U8747 ( .A(n8406), .B(n8407), .Z(n8323) );
  ANDN U8748 ( .B(n8408), .A(n8409), .Z(n8406) );
  XNOR U8749 ( .A(n8410), .B(n8328), .Z(n8330) );
  XOR U8750 ( .A(n8411), .B(n8412), .Z(n8328) );
  ANDN U8751 ( .B(n8413), .A(n8414), .Z(n8411) );
  AND U8752 ( .A(a[23]), .B(b[9]), .Z(n8410) );
  XOR U8753 ( .A(n8416), .B(n8417), .Z(n8333) );
  ANDN U8754 ( .B(n8345), .A(n8372), .Z(n8416) );
  AND U8755 ( .A(a[25]), .B(b[6]), .Z(n8418) );
  XNOR U8756 ( .A(n8408), .B(n8417), .Z(n8419) );
  XOR U8757 ( .A(n8420), .B(n8421), .Z(n8417) );
  ANDN U8758 ( .B(n8350), .A(n8371), .Z(n8420) );
  AND U8759 ( .A(a[25]), .B(b[5]), .Z(n8422) );
  XNOR U8760 ( .A(n8424), .B(n8421), .Z(n8423) );
  XOR U8761 ( .A(n8425), .B(n8426), .Z(n8421) );
  ANDN U8762 ( .B(n8355), .A(n8370), .Z(n8425) );
  AND U8763 ( .A(a[25]), .B(b[4]), .Z(n8427) );
  XNOR U8764 ( .A(n8429), .B(n8426), .Z(n8428) );
  XOR U8765 ( .A(n8430), .B(n8431), .Z(n8426) );
  ANDN U8766 ( .B(n8360), .A(n8369), .Z(n8430) );
  AND U8767 ( .A(a[25]), .B(b[3]), .Z(n8432) );
  XNOR U8768 ( .A(n8434), .B(n8431), .Z(n8433) );
  XOR U8769 ( .A(n8435), .B(n8436), .Z(n8431) );
  ANDN U8770 ( .B(n8365), .A(n8366), .Z(n8435) );
  AND U8771 ( .A(b[2]), .B(a[25]), .Z(n8437) );
  XNOR U8772 ( .A(n8439), .B(n8436), .Z(n8438) );
  XOR U8773 ( .A(n8440), .B(n8441), .Z(n8436) );
  NANDN U8774 ( .A(n8368), .B(n8367), .Z(n8441) );
  XOR U8775 ( .A(n8440), .B(n8442), .Z(n8367) );
  NAND U8776 ( .A(a[25]), .B(b[1]), .Z(n8442) );
  XNOR U8777 ( .A(n8440), .B(n8444), .Z(n8443) );
  OR U8778 ( .A(n2772), .B(n2770), .Z(n8440) );
  NANDN U8779 ( .A(n179), .B(a[25]), .Z(n2772) );
  XOR U8780 ( .A(n8452), .B(n8407), .Z(n8408) );
  AND U8781 ( .A(b[7]), .B(a[24]), .Z(n8452) );
  XNOR U8782 ( .A(n8407), .B(n8413), .Z(n8453) );
  XNOR U8783 ( .A(n8412), .B(n8404), .Z(n8454) );
  XNOR U8784 ( .A(n8403), .B(n8399), .Z(n8455) );
  XNOR U8785 ( .A(n8398), .B(n8394), .Z(n8456) );
  XOR U8786 ( .A(n8393), .B(n8390), .Z(n8457) );
  XOR U8787 ( .A(n8458), .B(n8459), .Z(n8390) );
  XOR U8788 ( .A(n8388), .B(n8460), .Z(n8459) );
  XOR U8789 ( .A(n8461), .B(n8462), .Z(n8460) );
  XOR U8790 ( .A(n8463), .B(n8464), .Z(n8462) );
  NAND U8791 ( .A(a[17]), .B(b[14]), .Z(n8464) );
  AND U8792 ( .A(a[16]), .B(b[15]), .Z(n8463) );
  XOR U8793 ( .A(n8465), .B(n8461), .Z(n8458) );
  XOR U8794 ( .A(n8466), .B(n8467), .Z(n8461) );
  NOR U8795 ( .A(n8468), .B(n8469), .Z(n8466) );
  AND U8796 ( .A(a[18]), .B(b[13]), .Z(n8465) );
  XNOR U8797 ( .A(n8470), .B(n8388), .Z(n8389) );
  XOR U8798 ( .A(n8471), .B(n8472), .Z(n8388) );
  ANDN U8799 ( .B(n8473), .A(n8474), .Z(n8471) );
  AND U8800 ( .A(a[19]), .B(b[12]), .Z(n8470) );
  XNOR U8801 ( .A(n8475), .B(n8393), .Z(n8395) );
  XOR U8802 ( .A(n8476), .B(n8477), .Z(n8393) );
  ANDN U8803 ( .B(n8478), .A(n8479), .Z(n8476) );
  AND U8804 ( .A(a[20]), .B(b[11]), .Z(n8475) );
  XNOR U8805 ( .A(n8480), .B(n8398), .Z(n8400) );
  XOR U8806 ( .A(n8481), .B(n8482), .Z(n8398) );
  ANDN U8807 ( .B(n8483), .A(n8484), .Z(n8481) );
  AND U8808 ( .A(a[21]), .B(b[10]), .Z(n8480) );
  XNOR U8809 ( .A(n8485), .B(n8403), .Z(n8405) );
  XOR U8810 ( .A(n8486), .B(n8487), .Z(n8403) );
  ANDN U8811 ( .B(n8488), .A(n8489), .Z(n8486) );
  AND U8812 ( .A(a[22]), .B(b[9]), .Z(n8485) );
  XOR U8813 ( .A(n8490), .B(n8491), .Z(n8407) );
  ANDN U8814 ( .B(n8424), .A(n8451), .Z(n8490) );
  XNOR U8815 ( .A(n8491), .B(n8493), .Z(n8492) );
  XOR U8816 ( .A(n8495), .B(n8491), .Z(n8424) );
  XOR U8817 ( .A(n8496), .B(n8497), .Z(n8491) );
  ANDN U8818 ( .B(n8429), .A(n8450), .Z(n8496) );
  XNOR U8819 ( .A(n8497), .B(n8499), .Z(n8498) );
  XOR U8820 ( .A(n8501), .B(n8497), .Z(n8429) );
  XOR U8821 ( .A(n8502), .B(n8503), .Z(n8497) );
  ANDN U8822 ( .B(n8434), .A(n8449), .Z(n8502) );
  XNOR U8823 ( .A(n8503), .B(n8505), .Z(n8504) );
  XOR U8824 ( .A(n8507), .B(n8503), .Z(n8434) );
  XOR U8825 ( .A(n8508), .B(n8509), .Z(n8503) );
  ANDN U8826 ( .B(n8439), .A(n8448), .Z(n8508) );
  XNOR U8827 ( .A(n8509), .B(n8511), .Z(n8510) );
  XOR U8828 ( .A(n8513), .B(n8509), .Z(n8439) );
  XNOR U8829 ( .A(n8514), .B(n8515), .Z(n8509) );
  NOR U8830 ( .A(n8445), .B(n8444), .Z(n8514) );
  XOR U8831 ( .A(n8516), .B(n8515), .Z(n8444) );
  AND U8832 ( .A(b[2]), .B(a[24]), .Z(n8516) );
  XOR U8833 ( .A(n8515), .B(n8518), .Z(n8517) );
  XNOR U8834 ( .A(n8519), .B(n8520), .Z(n8515) );
  OR U8835 ( .A(n8446), .B(n8447), .Z(n8520) );
  XNOR U8836 ( .A(n8519), .B(n8522), .Z(n8521) );
  XNOR U8837 ( .A(n8519), .B(n8524), .Z(n8446) );
  NAND U8838 ( .A(b[1]), .B(a[24]), .Z(n8524) );
  OR U8839 ( .A(n2777), .B(n2775), .Z(n8519) );
  XOR U8840 ( .A(n8525), .B(n8526), .Z(n2775) );
  NANDN U8841 ( .A(n179), .B(a[24]), .Z(n2777) );
  AND U8842 ( .A(b[3]), .B(a[24]), .Z(n8513) );
  AND U8843 ( .A(b[4]), .B(a[24]), .Z(n8507) );
  AND U8844 ( .A(b[5]), .B(a[24]), .Z(n8501) );
  AND U8845 ( .A(b[6]), .B(a[24]), .Z(n8495) );
  XNOR U8846 ( .A(n8528), .B(n8412), .Z(n8414) );
  XOR U8847 ( .A(n8529), .B(n8530), .Z(n8412) );
  ANDN U8848 ( .B(n8493), .A(n8494), .Z(n8529) );
  XNOR U8849 ( .A(n8531), .B(n8530), .Z(n8494) );
  AND U8850 ( .A(a[23]), .B(b[7]), .Z(n8531) );
  XNOR U8851 ( .A(n8530), .B(n8488), .Z(n8532) );
  XNOR U8852 ( .A(n8487), .B(n8483), .Z(n8533) );
  XNOR U8853 ( .A(n8482), .B(n8478), .Z(n8534) );
  XNOR U8854 ( .A(n8477), .B(n8473), .Z(n8535) );
  XOR U8855 ( .A(n8472), .B(n8469), .Z(n8536) );
  XOR U8856 ( .A(n8537), .B(n8538), .Z(n8469) );
  XOR U8857 ( .A(n8467), .B(n8539), .Z(n8538) );
  XOR U8858 ( .A(n8540), .B(n8541), .Z(n8539) );
  XOR U8859 ( .A(n8542), .B(n8543), .Z(n8541) );
  NAND U8860 ( .A(a[16]), .B(b[14]), .Z(n8543) );
  AND U8861 ( .A(a[15]), .B(b[15]), .Z(n8542) );
  XOR U8862 ( .A(n8544), .B(n8540), .Z(n8537) );
  XOR U8863 ( .A(n8545), .B(n8546), .Z(n8540) );
  NOR U8864 ( .A(n8547), .B(n8548), .Z(n8545) );
  AND U8865 ( .A(a[17]), .B(b[13]), .Z(n8544) );
  XNOR U8866 ( .A(n8549), .B(n8467), .Z(n8468) );
  XOR U8867 ( .A(n8550), .B(n8551), .Z(n8467) );
  ANDN U8868 ( .B(n8552), .A(n8553), .Z(n8550) );
  AND U8869 ( .A(a[18]), .B(b[12]), .Z(n8549) );
  XNOR U8870 ( .A(n8554), .B(n8472), .Z(n8474) );
  XOR U8871 ( .A(n8555), .B(n8556), .Z(n8472) );
  ANDN U8872 ( .B(n8557), .A(n8558), .Z(n8555) );
  AND U8873 ( .A(a[19]), .B(b[11]), .Z(n8554) );
  XNOR U8874 ( .A(n8559), .B(n8477), .Z(n8479) );
  XOR U8875 ( .A(n8560), .B(n8561), .Z(n8477) );
  ANDN U8876 ( .B(n8562), .A(n8563), .Z(n8560) );
  AND U8877 ( .A(a[20]), .B(b[10]), .Z(n8559) );
  XNOR U8878 ( .A(n8564), .B(n8482), .Z(n8484) );
  XOR U8879 ( .A(n8565), .B(n8566), .Z(n8482) );
  ANDN U8880 ( .B(n8567), .A(n8568), .Z(n8565) );
  AND U8881 ( .A(a[21]), .B(b[9]), .Z(n8564) );
  XOR U8882 ( .A(n8569), .B(n8570), .Z(n8530) );
  ANDN U8883 ( .B(n8499), .A(n8500), .Z(n8569) );
  XNOR U8884 ( .A(n8571), .B(n8570), .Z(n8500) );
  AND U8885 ( .A(a[23]), .B(b[6]), .Z(n8571) );
  XNOR U8886 ( .A(n8570), .B(n8573), .Z(n8572) );
  XOR U8887 ( .A(n8574), .B(n8575), .Z(n8570) );
  ANDN U8888 ( .B(n8505), .A(n8506), .Z(n8574) );
  XNOR U8889 ( .A(n8576), .B(n8575), .Z(n8506) );
  AND U8890 ( .A(a[23]), .B(b[5]), .Z(n8576) );
  XNOR U8891 ( .A(n8575), .B(n8578), .Z(n8577) );
  XOR U8892 ( .A(n8579), .B(n8580), .Z(n8575) );
  ANDN U8893 ( .B(n8511), .A(n8512), .Z(n8579) );
  XNOR U8894 ( .A(n8581), .B(n8580), .Z(n8512) );
  AND U8895 ( .A(a[23]), .B(b[4]), .Z(n8581) );
  XNOR U8896 ( .A(n8580), .B(n8583), .Z(n8582) );
  XOR U8897 ( .A(n8584), .B(n8585), .Z(n8580) );
  ANDN U8898 ( .B(n8518), .A(n8527), .Z(n8584) );
  XNOR U8899 ( .A(n8586), .B(n8585), .Z(n8527) );
  AND U8900 ( .A(a[23]), .B(b[3]), .Z(n8586) );
  XNOR U8901 ( .A(n8585), .B(n8588), .Z(n8587) );
  XNOR U8902 ( .A(n8589), .B(n8590), .Z(n8585) );
  NOR U8903 ( .A(n8523), .B(n8522), .Z(n8589) );
  XOR U8904 ( .A(n8591), .B(n8590), .Z(n8522) );
  AND U8905 ( .A(b[2]), .B(a[23]), .Z(n8591) );
  XOR U8906 ( .A(n8590), .B(n8593), .Z(n8592) );
  XNOR U8907 ( .A(n8594), .B(n8595), .Z(n8590) );
  NANDN U8908 ( .A(n8526), .B(n8525), .Z(n8595) );
  XOR U8909 ( .A(n8594), .B(n8596), .Z(n8525) );
  NAND U8910 ( .A(a[23]), .B(b[1]), .Z(n8596) );
  XOR U8911 ( .A(n8594), .B(n8598), .Z(n8597) );
  OR U8912 ( .A(n2782), .B(n2780), .Z(n8594) );
  XOR U8913 ( .A(n8600), .B(n8601), .Z(n2780) );
  NANDN U8914 ( .A(n179), .B(a[23]), .Z(n2782) );
  XNOR U8915 ( .A(n8607), .B(n8487), .Z(n8489) );
  XOR U8916 ( .A(n8608), .B(n8609), .Z(n8487) );
  ANDN U8917 ( .B(n8573), .A(n8606), .Z(n8608) );
  XNOR U8918 ( .A(n8610), .B(n8609), .Z(n8606) );
  AND U8919 ( .A(a[22]), .B(b[7]), .Z(n8610) );
  XNOR U8920 ( .A(n8609), .B(n8567), .Z(n8611) );
  XNOR U8921 ( .A(n8566), .B(n8562), .Z(n8612) );
  XNOR U8922 ( .A(n8561), .B(n8557), .Z(n8613) );
  XNOR U8923 ( .A(n8556), .B(n8552), .Z(n8614) );
  XOR U8924 ( .A(n8551), .B(n8548), .Z(n8615) );
  XOR U8925 ( .A(n8616), .B(n8617), .Z(n8548) );
  XOR U8926 ( .A(n8546), .B(n8618), .Z(n8617) );
  XOR U8927 ( .A(n8619), .B(n8620), .Z(n8618) );
  XOR U8928 ( .A(n8621), .B(n8622), .Z(n8620) );
  NAND U8929 ( .A(a[15]), .B(b[14]), .Z(n8622) );
  AND U8930 ( .A(a[14]), .B(b[15]), .Z(n8621) );
  XOR U8931 ( .A(n8623), .B(n8619), .Z(n8616) );
  XOR U8932 ( .A(n8624), .B(n8625), .Z(n8619) );
  NOR U8933 ( .A(n8626), .B(n8627), .Z(n8624) );
  AND U8934 ( .A(a[16]), .B(b[13]), .Z(n8623) );
  XNOR U8935 ( .A(n8628), .B(n8546), .Z(n8547) );
  XOR U8936 ( .A(n8629), .B(n8630), .Z(n8546) );
  ANDN U8937 ( .B(n8631), .A(n8632), .Z(n8629) );
  AND U8938 ( .A(a[17]), .B(b[12]), .Z(n8628) );
  XNOR U8939 ( .A(n8633), .B(n8551), .Z(n8553) );
  XOR U8940 ( .A(n8634), .B(n8635), .Z(n8551) );
  ANDN U8941 ( .B(n8636), .A(n8637), .Z(n8634) );
  AND U8942 ( .A(a[18]), .B(b[11]), .Z(n8633) );
  XNOR U8943 ( .A(n8638), .B(n8556), .Z(n8558) );
  XOR U8944 ( .A(n8639), .B(n8640), .Z(n8556) );
  ANDN U8945 ( .B(n8641), .A(n8642), .Z(n8639) );
  AND U8946 ( .A(a[19]), .B(b[10]), .Z(n8638) );
  XNOR U8947 ( .A(n8643), .B(n8561), .Z(n8563) );
  XOR U8948 ( .A(n8644), .B(n8645), .Z(n8561) );
  ANDN U8949 ( .B(n8646), .A(n8647), .Z(n8644) );
  AND U8950 ( .A(a[20]), .B(b[9]), .Z(n8643) );
  XOR U8951 ( .A(n8648), .B(n8649), .Z(n8609) );
  ANDN U8952 ( .B(n8578), .A(n8605), .Z(n8648) );
  XNOR U8953 ( .A(n8650), .B(n8649), .Z(n8605) );
  AND U8954 ( .A(a[22]), .B(b[6]), .Z(n8650) );
  XNOR U8955 ( .A(n8649), .B(n8652), .Z(n8651) );
  XOR U8956 ( .A(n8653), .B(n8654), .Z(n8649) );
  ANDN U8957 ( .B(n8583), .A(n8604), .Z(n8653) );
  XNOR U8958 ( .A(n8655), .B(n8654), .Z(n8604) );
  AND U8959 ( .A(a[22]), .B(b[5]), .Z(n8655) );
  XNOR U8960 ( .A(n8654), .B(n8657), .Z(n8656) );
  XOR U8961 ( .A(n8658), .B(n8659), .Z(n8654) );
  ANDN U8962 ( .B(n8588), .A(n8603), .Z(n8658) );
  XNOR U8963 ( .A(n8660), .B(n8659), .Z(n8603) );
  AND U8964 ( .A(a[22]), .B(b[4]), .Z(n8660) );
  XNOR U8965 ( .A(n8659), .B(n8662), .Z(n8661) );
  XOR U8966 ( .A(n8663), .B(n8664), .Z(n8659) );
  ANDN U8967 ( .B(n8593), .A(n8602), .Z(n8663) );
  XNOR U8968 ( .A(n8665), .B(n8664), .Z(n8602) );
  AND U8969 ( .A(a[22]), .B(b[3]), .Z(n8665) );
  XNOR U8970 ( .A(n8664), .B(n8667), .Z(n8666) );
  XNOR U8971 ( .A(n8668), .B(n8669), .Z(n8664) );
  ANDN U8972 ( .B(n8598), .A(n8599), .Z(n8668) );
  XOR U8973 ( .A(n8670), .B(n8669), .Z(n8599) );
  IV U8974 ( .A(n8671), .Z(n8669) );
  AND U8975 ( .A(b[2]), .B(a[22]), .Z(n8670) );
  XNOR U8976 ( .A(n8673), .B(n8671), .Z(n8672) );
  XOR U8977 ( .A(n8674), .B(n8675), .Z(n8671) );
  NANDN U8978 ( .A(n8601), .B(n8600), .Z(n8675) );
  XOR U8979 ( .A(n8674), .B(n8676), .Z(n8600) );
  NAND U8980 ( .A(a[22]), .B(b[1]), .Z(n8676) );
  XOR U8981 ( .A(n8674), .B(n8678), .Z(n8677) );
  OR U8982 ( .A(n2787), .B(n2785), .Z(n8674) );
  XOR U8983 ( .A(n8680), .B(n8681), .Z(n2785) );
  NANDN U8984 ( .A(n179), .B(a[22]), .Z(n2787) );
  XNOR U8985 ( .A(n8687), .B(n8566), .Z(n8568) );
  XOR U8986 ( .A(n8688), .B(n8689), .Z(n8566) );
  ANDN U8987 ( .B(n8652), .A(n8686), .Z(n8688) );
  XNOR U8988 ( .A(n8690), .B(n8689), .Z(n8686) );
  AND U8989 ( .A(a[21]), .B(b[7]), .Z(n8690) );
  XNOR U8990 ( .A(n8689), .B(n8646), .Z(n8691) );
  XNOR U8991 ( .A(n8645), .B(n8641), .Z(n8692) );
  XNOR U8992 ( .A(n8640), .B(n8636), .Z(n8693) );
  XNOR U8993 ( .A(n8635), .B(n8631), .Z(n8694) );
  XOR U8994 ( .A(n8630), .B(n8627), .Z(n8695) );
  XOR U8995 ( .A(n8696), .B(n8697), .Z(n8627) );
  XOR U8996 ( .A(n8625), .B(n8698), .Z(n8697) );
  XOR U8997 ( .A(n8699), .B(n8700), .Z(n8698) );
  XOR U8998 ( .A(n8701), .B(n8702), .Z(n8700) );
  NAND U8999 ( .A(b[14]), .B(a[14]), .Z(n8702) );
  AND U9000 ( .A(a[13]), .B(b[15]), .Z(n8701) );
  XOR U9001 ( .A(n8703), .B(n8699), .Z(n8696) );
  XOR U9002 ( .A(n8704), .B(n8705), .Z(n8699) );
  NOR U9003 ( .A(n8706), .B(n8707), .Z(n8704) );
  AND U9004 ( .A(a[15]), .B(b[13]), .Z(n8703) );
  XNOR U9005 ( .A(n8708), .B(n8625), .Z(n8626) );
  XOR U9006 ( .A(n8709), .B(n8710), .Z(n8625) );
  ANDN U9007 ( .B(n8711), .A(n8712), .Z(n8709) );
  AND U9008 ( .A(a[16]), .B(b[12]), .Z(n8708) );
  XNOR U9009 ( .A(n8713), .B(n8630), .Z(n8632) );
  XOR U9010 ( .A(n8714), .B(n8715), .Z(n8630) );
  ANDN U9011 ( .B(n8716), .A(n8717), .Z(n8714) );
  AND U9012 ( .A(a[17]), .B(b[11]), .Z(n8713) );
  XNOR U9013 ( .A(n8718), .B(n8635), .Z(n8637) );
  XOR U9014 ( .A(n8719), .B(n8720), .Z(n8635) );
  ANDN U9015 ( .B(n8721), .A(n8722), .Z(n8719) );
  AND U9016 ( .A(a[18]), .B(b[10]), .Z(n8718) );
  XNOR U9017 ( .A(n8723), .B(n8640), .Z(n8642) );
  XOR U9018 ( .A(n8724), .B(n8725), .Z(n8640) );
  ANDN U9019 ( .B(n8726), .A(n8727), .Z(n8724) );
  AND U9020 ( .A(a[19]), .B(b[9]), .Z(n8723) );
  XOR U9021 ( .A(n8728), .B(n8729), .Z(n8689) );
  ANDN U9022 ( .B(n8657), .A(n8685), .Z(n8728) );
  XNOR U9023 ( .A(n8730), .B(n8729), .Z(n8685) );
  AND U9024 ( .A(a[21]), .B(b[6]), .Z(n8730) );
  XNOR U9025 ( .A(n8729), .B(n8732), .Z(n8731) );
  XOR U9026 ( .A(n8733), .B(n8734), .Z(n8729) );
  ANDN U9027 ( .B(n8662), .A(n8684), .Z(n8733) );
  XNOR U9028 ( .A(n8735), .B(n8734), .Z(n8684) );
  AND U9029 ( .A(a[21]), .B(b[5]), .Z(n8735) );
  XNOR U9030 ( .A(n8734), .B(n8737), .Z(n8736) );
  XOR U9031 ( .A(n8738), .B(n8739), .Z(n8734) );
  ANDN U9032 ( .B(n8667), .A(n8683), .Z(n8738) );
  XNOR U9033 ( .A(n8740), .B(n8739), .Z(n8683) );
  AND U9034 ( .A(a[21]), .B(b[4]), .Z(n8740) );
  XNOR U9035 ( .A(n8739), .B(n8742), .Z(n8741) );
  XNOR U9036 ( .A(n8743), .B(n8744), .Z(n8739) );
  ANDN U9037 ( .B(n8673), .A(n8682), .Z(n8743) );
  XOR U9038 ( .A(n8745), .B(n8744), .Z(n8682) );
  IV U9039 ( .A(n8746), .Z(n8744) );
  AND U9040 ( .A(a[21]), .B(b[3]), .Z(n8745) );
  XNOR U9041 ( .A(n8748), .B(n8746), .Z(n8747) );
  XOR U9042 ( .A(n8749), .B(n8750), .Z(n8746) );
  ANDN U9043 ( .B(n8678), .A(n8679), .Z(n8749) );
  AND U9044 ( .A(b[2]), .B(a[21]), .Z(n8751) );
  XNOR U9045 ( .A(n8753), .B(n8750), .Z(n8752) );
  XOR U9046 ( .A(n8754), .B(n8755), .Z(n8750) );
  NANDN U9047 ( .A(n8681), .B(n8680), .Z(n8755) );
  XOR U9048 ( .A(n8754), .B(n8756), .Z(n8680) );
  NAND U9049 ( .A(a[21]), .B(b[1]), .Z(n8756) );
  XOR U9050 ( .A(n8754), .B(n8758), .Z(n8757) );
  OR U9051 ( .A(n2792), .B(n2790), .Z(n8754) );
  XOR U9052 ( .A(n8760), .B(n8761), .Z(n2790) );
  NANDN U9053 ( .A(n179), .B(a[21]), .Z(n2792) );
  XNOR U9054 ( .A(n8767), .B(n8645), .Z(n8647) );
  XOR U9055 ( .A(n8768), .B(n8769), .Z(n8645) );
  ANDN U9056 ( .B(n8732), .A(n8766), .Z(n8768) );
  XNOR U9057 ( .A(n8770), .B(n8769), .Z(n8766) );
  AND U9058 ( .A(a[20]), .B(b[7]), .Z(n8770) );
  XNOR U9059 ( .A(n8769), .B(n8726), .Z(n8771) );
  XNOR U9060 ( .A(n8725), .B(n8721), .Z(n8772) );
  XNOR U9061 ( .A(n8720), .B(n8716), .Z(n8773) );
  XNOR U9062 ( .A(n8715), .B(n8711), .Z(n8774) );
  XOR U9063 ( .A(n8710), .B(n8707), .Z(n8775) );
  XOR U9064 ( .A(n8776), .B(n8777), .Z(n8707) );
  XOR U9065 ( .A(n8705), .B(n8778), .Z(n8777) );
  XOR U9066 ( .A(n8779), .B(n8780), .Z(n8778) );
  XOR U9067 ( .A(n8781), .B(n8782), .Z(n8780) );
  NAND U9068 ( .A(a[13]), .B(b[14]), .Z(n8782) );
  AND U9069 ( .A(a[12]), .B(b[15]), .Z(n8781) );
  XOR U9070 ( .A(n8783), .B(n8779), .Z(n8776) );
  XOR U9071 ( .A(n8784), .B(n8785), .Z(n8779) );
  NOR U9072 ( .A(n8786), .B(n8787), .Z(n8784) );
  AND U9073 ( .A(b[13]), .B(a[14]), .Z(n8783) );
  XNOR U9074 ( .A(n8788), .B(n8705), .Z(n8706) );
  XOR U9075 ( .A(n8789), .B(n8790), .Z(n8705) );
  ANDN U9076 ( .B(n8791), .A(n8792), .Z(n8789) );
  AND U9077 ( .A(a[15]), .B(b[12]), .Z(n8788) );
  XNOR U9078 ( .A(n8793), .B(n8710), .Z(n8712) );
  XOR U9079 ( .A(n8794), .B(n8795), .Z(n8710) );
  ANDN U9080 ( .B(n8796), .A(n8797), .Z(n8794) );
  AND U9081 ( .A(a[16]), .B(b[11]), .Z(n8793) );
  XNOR U9082 ( .A(n8798), .B(n8715), .Z(n8717) );
  XOR U9083 ( .A(n8799), .B(n8800), .Z(n8715) );
  ANDN U9084 ( .B(n8801), .A(n8802), .Z(n8799) );
  AND U9085 ( .A(a[17]), .B(b[10]), .Z(n8798) );
  XNOR U9086 ( .A(n8803), .B(n8720), .Z(n8722) );
  XOR U9087 ( .A(n8804), .B(n8805), .Z(n8720) );
  ANDN U9088 ( .B(n8806), .A(n8807), .Z(n8804) );
  AND U9089 ( .A(a[18]), .B(b[9]), .Z(n8803) );
  XOR U9090 ( .A(n8808), .B(n8809), .Z(n8769) );
  ANDN U9091 ( .B(n8737), .A(n8765), .Z(n8808) );
  XNOR U9092 ( .A(n8810), .B(n8809), .Z(n8765) );
  AND U9093 ( .A(a[20]), .B(b[6]), .Z(n8810) );
  XNOR U9094 ( .A(n8809), .B(n8812), .Z(n8811) );
  XOR U9095 ( .A(n8813), .B(n8814), .Z(n8809) );
  ANDN U9096 ( .B(n8742), .A(n8764), .Z(n8813) );
  XNOR U9097 ( .A(n8815), .B(n8814), .Z(n8764) );
  AND U9098 ( .A(a[20]), .B(b[5]), .Z(n8815) );
  XNOR U9099 ( .A(n8814), .B(n8817), .Z(n8816) );
  XNOR U9100 ( .A(n8818), .B(n8819), .Z(n8814) );
  ANDN U9101 ( .B(n8748), .A(n8763), .Z(n8818) );
  XOR U9102 ( .A(n8820), .B(n8819), .Z(n8763) );
  IV U9103 ( .A(n8821), .Z(n8819) );
  AND U9104 ( .A(a[20]), .B(b[4]), .Z(n8820) );
  XNOR U9105 ( .A(n8823), .B(n8821), .Z(n8822) );
  XOR U9106 ( .A(n8824), .B(n8825), .Z(n8821) );
  ANDN U9107 ( .B(n8753), .A(n8762), .Z(n8824) );
  AND U9108 ( .A(a[20]), .B(b[3]), .Z(n8826) );
  XNOR U9109 ( .A(n8828), .B(n8825), .Z(n8827) );
  XOR U9110 ( .A(n8829), .B(n8830), .Z(n8825) );
  ANDN U9111 ( .B(n8758), .A(n8759), .Z(n8829) );
  AND U9112 ( .A(b[2]), .B(a[20]), .Z(n8831) );
  XNOR U9113 ( .A(n8833), .B(n8830), .Z(n8832) );
  XOR U9114 ( .A(n8834), .B(n8835), .Z(n8830) );
  NANDN U9115 ( .A(n8761), .B(n8760), .Z(n8835) );
  XOR U9116 ( .A(n8834), .B(n8836), .Z(n8760) );
  NAND U9117 ( .A(a[20]), .B(b[1]), .Z(n8836) );
  XOR U9118 ( .A(n8834), .B(n8838), .Z(n8837) );
  OR U9119 ( .A(n2797), .B(n2795), .Z(n8834) );
  XOR U9120 ( .A(n8840), .B(n8841), .Z(n2795) );
  NANDN U9121 ( .A(n179), .B(a[20]), .Z(n2797) );
  XNOR U9122 ( .A(n8847), .B(n8725), .Z(n8727) );
  XOR U9123 ( .A(n8848), .B(n8849), .Z(n8725) );
  ANDN U9124 ( .B(n8812), .A(n8846), .Z(n8848) );
  XNOR U9125 ( .A(n8850), .B(n8849), .Z(n8846) );
  AND U9126 ( .A(a[19]), .B(b[7]), .Z(n8850) );
  XNOR U9127 ( .A(n8849), .B(n8806), .Z(n8851) );
  XNOR U9128 ( .A(n8805), .B(n8801), .Z(n8852) );
  XNOR U9129 ( .A(n8800), .B(n8796), .Z(n8853) );
  XNOR U9130 ( .A(n8795), .B(n8791), .Z(n8854) );
  XOR U9131 ( .A(n8790), .B(n8787), .Z(n8855) );
  XOR U9132 ( .A(n8856), .B(n8857), .Z(n8787) );
  XOR U9133 ( .A(n8785), .B(n8858), .Z(n8857) );
  XOR U9134 ( .A(n8859), .B(n8860), .Z(n8858) );
  XOR U9135 ( .A(n8861), .B(n8862), .Z(n8860) );
  NAND U9136 ( .A(a[12]), .B(b[14]), .Z(n8862) );
  AND U9137 ( .A(a[11]), .B(b[15]), .Z(n8861) );
  XOR U9138 ( .A(n8863), .B(n8859), .Z(n8856) );
  XOR U9139 ( .A(n8864), .B(n8865), .Z(n8859) );
  NOR U9140 ( .A(n8866), .B(n8867), .Z(n8864) );
  AND U9141 ( .A(a[13]), .B(b[13]), .Z(n8863) );
  XNOR U9142 ( .A(n8868), .B(n8785), .Z(n8786) );
  XOR U9143 ( .A(n8869), .B(n8870), .Z(n8785) );
  ANDN U9144 ( .B(n8871), .A(n8872), .Z(n8869) );
  AND U9145 ( .A(b[12]), .B(a[14]), .Z(n8868) );
  XNOR U9146 ( .A(n8873), .B(n8790), .Z(n8792) );
  XOR U9147 ( .A(n8874), .B(n8875), .Z(n8790) );
  ANDN U9148 ( .B(n8876), .A(n8877), .Z(n8874) );
  AND U9149 ( .A(a[15]), .B(b[11]), .Z(n8873) );
  XNOR U9150 ( .A(n8878), .B(n8795), .Z(n8797) );
  XOR U9151 ( .A(n8879), .B(n8880), .Z(n8795) );
  ANDN U9152 ( .B(n8881), .A(n8882), .Z(n8879) );
  AND U9153 ( .A(a[16]), .B(b[10]), .Z(n8878) );
  XNOR U9154 ( .A(n8883), .B(n8800), .Z(n8802) );
  XOR U9155 ( .A(n8884), .B(n8885), .Z(n8800) );
  ANDN U9156 ( .B(n8886), .A(n8887), .Z(n8884) );
  AND U9157 ( .A(a[17]), .B(b[9]), .Z(n8883) );
  XOR U9158 ( .A(n8888), .B(n8889), .Z(n8849) );
  ANDN U9159 ( .B(n8817), .A(n8845), .Z(n8888) );
  XNOR U9160 ( .A(n8890), .B(n8889), .Z(n8845) );
  AND U9161 ( .A(a[19]), .B(b[6]), .Z(n8890) );
  XNOR U9162 ( .A(n8889), .B(n8892), .Z(n8891) );
  XNOR U9163 ( .A(n8893), .B(n8894), .Z(n8889) );
  ANDN U9164 ( .B(n8823), .A(n8844), .Z(n8893) );
  XOR U9165 ( .A(n8895), .B(n8894), .Z(n8844) );
  IV U9166 ( .A(n8896), .Z(n8894) );
  AND U9167 ( .A(a[19]), .B(b[5]), .Z(n8895) );
  XNOR U9168 ( .A(n8898), .B(n8896), .Z(n8897) );
  XOR U9169 ( .A(n8899), .B(n8900), .Z(n8896) );
  ANDN U9170 ( .B(n8828), .A(n8843), .Z(n8899) );
  AND U9171 ( .A(a[19]), .B(b[4]), .Z(n8901) );
  XNOR U9172 ( .A(n8903), .B(n8900), .Z(n8902) );
  XOR U9173 ( .A(n8904), .B(n8905), .Z(n8900) );
  ANDN U9174 ( .B(n8833), .A(n8842), .Z(n8904) );
  AND U9175 ( .A(a[19]), .B(b[3]), .Z(n8906) );
  XNOR U9176 ( .A(n8908), .B(n8905), .Z(n8907) );
  XOR U9177 ( .A(n8909), .B(n8910), .Z(n8905) );
  ANDN U9178 ( .B(n8838), .A(n8839), .Z(n8909) );
  AND U9179 ( .A(b[2]), .B(a[19]), .Z(n8911) );
  XNOR U9180 ( .A(n8913), .B(n8910), .Z(n8912) );
  XOR U9181 ( .A(n8914), .B(n8915), .Z(n8910) );
  NANDN U9182 ( .A(n8841), .B(n8840), .Z(n8915) );
  XOR U9183 ( .A(n8914), .B(n8916), .Z(n8840) );
  NAND U9184 ( .A(a[19]), .B(b[1]), .Z(n8916) );
  XOR U9185 ( .A(n8914), .B(n8918), .Z(n8917) );
  OR U9186 ( .A(n2802), .B(n2800), .Z(n8914) );
  XOR U9187 ( .A(n8920), .B(n8921), .Z(n2800) );
  NANDN U9188 ( .A(n179), .B(a[19]), .Z(n2802) );
  XNOR U9189 ( .A(n8927), .B(n8805), .Z(n8807) );
  XOR U9190 ( .A(n8928), .B(n8929), .Z(n8805) );
  ANDN U9191 ( .B(n8892), .A(n8926), .Z(n8928) );
  XNOR U9192 ( .A(n8930), .B(n8929), .Z(n8926) );
  AND U9193 ( .A(a[18]), .B(b[7]), .Z(n8930) );
  XNOR U9194 ( .A(n8929), .B(n8886), .Z(n8931) );
  XNOR U9195 ( .A(n8885), .B(n8881), .Z(n8932) );
  XNOR U9196 ( .A(n8880), .B(n8876), .Z(n8933) );
  XNOR U9197 ( .A(n8875), .B(n8871), .Z(n8934) );
  XOR U9198 ( .A(n8870), .B(n8867), .Z(n8935) );
  XOR U9199 ( .A(n8936), .B(n8937), .Z(n8867) );
  XOR U9200 ( .A(n8865), .B(n8938), .Z(n8937) );
  XNOR U9201 ( .A(n8939), .B(n8940), .Z(n8938) );
  XOR U9202 ( .A(n8941), .B(n8942), .Z(n8940) );
  NAND U9203 ( .A(a[11]), .B(b[14]), .Z(n8942) );
  AND U9204 ( .A(a[10]), .B(b[15]), .Z(n8941) );
  XNOR U9205 ( .A(n8943), .B(n8939), .Z(n8936) );
  XOR U9206 ( .A(n8944), .B(n8945), .Z(n8939) );
  NOR U9207 ( .A(n8946), .B(n8947), .Z(n8944) );
  AND U9208 ( .A(a[12]), .B(b[13]), .Z(n8943) );
  XNOR U9209 ( .A(n8948), .B(n8865), .Z(n8866) );
  XNOR U9210 ( .A(n8949), .B(n8950), .Z(n8865) );
  ANDN U9211 ( .B(n8951), .A(n8952), .Z(n8949) );
  AND U9212 ( .A(a[13]), .B(b[12]), .Z(n8948) );
  XNOR U9213 ( .A(n8953), .B(n8870), .Z(n8872) );
  XNOR U9214 ( .A(n8954), .B(n8955), .Z(n8870) );
  ANDN U9215 ( .B(n8956), .A(n8957), .Z(n8954) );
  AND U9216 ( .A(b[11]), .B(a[14]), .Z(n8953) );
  XNOR U9217 ( .A(n8958), .B(n8875), .Z(n8877) );
  XNOR U9218 ( .A(n8959), .B(n8960), .Z(n8875) );
  ANDN U9219 ( .B(n8961), .A(n8962), .Z(n8959) );
  AND U9220 ( .A(a[15]), .B(b[10]), .Z(n8958) );
  XNOR U9221 ( .A(n8963), .B(n8880), .Z(n8882) );
  XNOR U9222 ( .A(n8964), .B(n8965), .Z(n8880) );
  ANDN U9223 ( .B(n8966), .A(n8967), .Z(n8964) );
  AND U9224 ( .A(a[16]), .B(b[9]), .Z(n8963) );
  XNOR U9225 ( .A(n8968), .B(n8969), .Z(n8929) );
  ANDN U9226 ( .B(n8898), .A(n8925), .Z(n8968) );
  XOR U9227 ( .A(n8970), .B(n8969), .Z(n8925) );
  IV U9228 ( .A(n8971), .Z(n8969) );
  AND U9229 ( .A(a[18]), .B(b[6]), .Z(n8970) );
  XNOR U9230 ( .A(n8973), .B(n8971), .Z(n8972) );
  XOR U9231 ( .A(n8974), .B(n8975), .Z(n8971) );
  ANDN U9232 ( .B(n8903), .A(n8924), .Z(n8974) );
  AND U9233 ( .A(a[18]), .B(b[5]), .Z(n8976) );
  XNOR U9234 ( .A(n8978), .B(n8975), .Z(n8977) );
  XOR U9235 ( .A(n8979), .B(n8980), .Z(n8975) );
  ANDN U9236 ( .B(n8908), .A(n8923), .Z(n8979) );
  AND U9237 ( .A(a[18]), .B(b[4]), .Z(n8981) );
  XNOR U9238 ( .A(n8983), .B(n8980), .Z(n8982) );
  XOR U9239 ( .A(n8984), .B(n8985), .Z(n8980) );
  ANDN U9240 ( .B(n8913), .A(n8922), .Z(n8984) );
  AND U9241 ( .A(a[18]), .B(b[3]), .Z(n8986) );
  XNOR U9242 ( .A(n8988), .B(n8985), .Z(n8987) );
  XOR U9243 ( .A(n8989), .B(n8990), .Z(n8985) );
  ANDN U9244 ( .B(n8918), .A(n8919), .Z(n8989) );
  AND U9245 ( .A(b[2]), .B(a[18]), .Z(n8991) );
  XNOR U9246 ( .A(n8993), .B(n8990), .Z(n8992) );
  XOR U9247 ( .A(n8994), .B(n8995), .Z(n8990) );
  NANDN U9248 ( .A(n8921), .B(n8920), .Z(n8995) );
  XOR U9249 ( .A(n8994), .B(n8996), .Z(n8920) );
  NAND U9250 ( .A(a[18]), .B(b[1]), .Z(n8996) );
  XOR U9251 ( .A(n8994), .B(n8998), .Z(n8997) );
  OR U9252 ( .A(n2807), .B(n2805), .Z(n8994) );
  XOR U9253 ( .A(n9000), .B(n9001), .Z(n2805) );
  NANDN U9254 ( .A(n179), .B(a[18]), .Z(n2807) );
  XNOR U9255 ( .A(n9007), .B(n8885), .Z(n8887) );
  XNOR U9256 ( .A(n9008), .B(n9009), .Z(n8885) );
  ANDN U9257 ( .B(n8973), .A(n9006), .Z(n9008) );
  XOR U9258 ( .A(n9010), .B(n9009), .Z(n9006) );
  IV U9259 ( .A(n9011), .Z(n9009) );
  AND U9260 ( .A(a[17]), .B(b[7]), .Z(n9010) );
  XNOR U9261 ( .A(n8966), .B(n9011), .Z(n9012) );
  XOR U9262 ( .A(n9013), .B(n9014), .Z(n9011) );
  ANDN U9263 ( .B(n8978), .A(n9005), .Z(n9013) );
  AND U9264 ( .A(a[17]), .B(b[6]), .Z(n9015) );
  XNOR U9265 ( .A(n9017), .B(n9014), .Z(n9016) );
  XOR U9266 ( .A(n9018), .B(n9019), .Z(n9014) );
  ANDN U9267 ( .B(n8983), .A(n9004), .Z(n9018) );
  AND U9268 ( .A(a[17]), .B(b[5]), .Z(n9020) );
  XNOR U9269 ( .A(n9022), .B(n9019), .Z(n9021) );
  XOR U9270 ( .A(n9023), .B(n9024), .Z(n9019) );
  ANDN U9271 ( .B(n8988), .A(n9003), .Z(n9023) );
  AND U9272 ( .A(a[17]), .B(b[4]), .Z(n9025) );
  XNOR U9273 ( .A(n9027), .B(n9024), .Z(n9026) );
  XOR U9274 ( .A(n9028), .B(n9029), .Z(n9024) );
  ANDN U9275 ( .B(n8993), .A(n9002), .Z(n9028) );
  AND U9276 ( .A(a[17]), .B(b[3]), .Z(n9030) );
  XNOR U9277 ( .A(n9032), .B(n9029), .Z(n9031) );
  XOR U9278 ( .A(n9033), .B(n9034), .Z(n9029) );
  ANDN U9279 ( .B(n8998), .A(n8999), .Z(n9033) );
  AND U9280 ( .A(b[2]), .B(a[17]), .Z(n9035) );
  XNOR U9281 ( .A(n9037), .B(n9034), .Z(n9036) );
  XOR U9282 ( .A(n9038), .B(n9039), .Z(n9034) );
  NANDN U9283 ( .A(n9001), .B(n9000), .Z(n9039) );
  XOR U9284 ( .A(n9038), .B(n9040), .Z(n9000) );
  NAND U9285 ( .A(a[17]), .B(b[1]), .Z(n9040) );
  XOR U9286 ( .A(n9038), .B(n9042), .Z(n9041) );
  OR U9287 ( .A(n2812), .B(n2810), .Z(n9038) );
  XOR U9288 ( .A(n9044), .B(n9045), .Z(n2810) );
  NANDN U9289 ( .A(n179), .B(a[17]), .Z(n2812) );
  XNOR U9290 ( .A(n8961), .B(n9052), .Z(n9051) );
  XNOR U9291 ( .A(n8956), .B(n9054), .Z(n9053) );
  XNOR U9292 ( .A(n8951), .B(n9056), .Z(n9055) );
  XOR U9293 ( .A(n8947), .B(n9058), .Z(n9057) );
  XOR U9294 ( .A(n9059), .B(n9060), .Z(n8947) );
  XNOR U9295 ( .A(n9061), .B(n9062), .Z(n9060) );
  XNOR U9296 ( .A(n9063), .B(n9064), .Z(n9061) );
  XOR U9297 ( .A(n9065), .B(n9066), .Z(n9064) );
  AND U9298 ( .A(a[9]), .B(b[15]), .Z(n9066) );
  AND U9299 ( .A(a[10]), .B(b[14]), .Z(n9065) );
  XNOR U9300 ( .A(n9067), .B(n9063), .Z(n9059) );
  XOR U9301 ( .A(n9068), .B(n9069), .Z(n9063) );
  NOR U9302 ( .A(n9070), .B(n9071), .Z(n9068) );
  AND U9303 ( .A(a[11]), .B(b[13]), .Z(n9067) );
  XOR U9304 ( .A(n9072), .B(n8945), .Z(n8946) );
  IV U9305 ( .A(n9062), .Z(n8945) );
  XOR U9306 ( .A(n9073), .B(n9074), .Z(n9062) );
  ANDN U9307 ( .B(n9075), .A(n9076), .Z(n9073) );
  AND U9308 ( .A(b[12]), .B(a[12]), .Z(n9072) );
  XOR U9309 ( .A(n9077), .B(n8950), .Z(n8952) );
  IV U9310 ( .A(n9058), .Z(n8950) );
  XOR U9311 ( .A(n9078), .B(n9079), .Z(n9058) );
  ANDN U9312 ( .B(n9080), .A(n9081), .Z(n9078) );
  AND U9313 ( .A(a[13]), .B(b[11]), .Z(n9077) );
  XOR U9314 ( .A(n9082), .B(n8955), .Z(n8957) );
  IV U9315 ( .A(n9056), .Z(n8955) );
  XOR U9316 ( .A(n9083), .B(n9084), .Z(n9056) );
  ANDN U9317 ( .B(n9085), .A(n9086), .Z(n9083) );
  AND U9318 ( .A(b[10]), .B(a[14]), .Z(n9082) );
  XOR U9319 ( .A(n9087), .B(n8960), .Z(n8962) );
  IV U9320 ( .A(n9054), .Z(n8960) );
  XOR U9321 ( .A(n9088), .B(n9089), .Z(n9054) );
  ANDN U9322 ( .B(n9090), .A(n9091), .Z(n9088) );
  AND U9323 ( .A(a[15]), .B(b[9]), .Z(n9087) );
  XOR U9324 ( .A(n9092), .B(n8965), .Z(n8967) );
  IV U9325 ( .A(n9052), .Z(n8965) );
  XOR U9326 ( .A(n9093), .B(n9094), .Z(n9052) );
  ANDN U9327 ( .B(n9017), .A(n9050), .Z(n9093) );
  AND U9328 ( .A(a[16]), .B(b[7]), .Z(n9095) );
  XNOR U9329 ( .A(n9090), .B(n9094), .Z(n9096) );
  XOR U9330 ( .A(n9097), .B(n9098), .Z(n9094) );
  ANDN U9331 ( .B(n9022), .A(n9049), .Z(n9097) );
  AND U9332 ( .A(a[16]), .B(b[6]), .Z(n9099) );
  XNOR U9333 ( .A(n9101), .B(n9098), .Z(n9100) );
  XOR U9334 ( .A(n9102), .B(n9103), .Z(n9098) );
  ANDN U9335 ( .B(n9027), .A(n9048), .Z(n9102) );
  AND U9336 ( .A(a[16]), .B(b[5]), .Z(n9104) );
  XNOR U9337 ( .A(n9106), .B(n9103), .Z(n9105) );
  XOR U9338 ( .A(n9107), .B(n9108), .Z(n9103) );
  ANDN U9339 ( .B(n9032), .A(n9047), .Z(n9107) );
  AND U9340 ( .A(a[16]), .B(b[4]), .Z(n9109) );
  XNOR U9341 ( .A(n9111), .B(n9108), .Z(n9110) );
  XOR U9342 ( .A(n9112), .B(n9113), .Z(n9108) );
  ANDN U9343 ( .B(n9037), .A(n9046), .Z(n9112) );
  AND U9344 ( .A(a[16]), .B(b[3]), .Z(n9114) );
  XNOR U9345 ( .A(n9116), .B(n9113), .Z(n9115) );
  XOR U9346 ( .A(n9117), .B(n9118), .Z(n9113) );
  ANDN U9347 ( .B(n9042), .A(n9043), .Z(n9117) );
  AND U9348 ( .A(b[2]), .B(a[16]), .Z(n9119) );
  XNOR U9349 ( .A(n9121), .B(n9118), .Z(n9120) );
  XOR U9350 ( .A(n9122), .B(n9123), .Z(n9118) );
  NANDN U9351 ( .A(n9045), .B(n9044), .Z(n9123) );
  XOR U9352 ( .A(n9122), .B(n9124), .Z(n9044) );
  NAND U9353 ( .A(a[16]), .B(b[1]), .Z(n9124) );
  XOR U9354 ( .A(n9122), .B(n9126), .Z(n9125) );
  OR U9355 ( .A(n2817), .B(n2815), .Z(n9122) );
  XOR U9356 ( .A(n9128), .B(n9129), .Z(n2815) );
  NANDN U9357 ( .A(n179), .B(a[16]), .Z(n2817) );
  XNOR U9358 ( .A(n9085), .B(n9089), .Z(n9135) );
  XNOR U9359 ( .A(n9080), .B(n9084), .Z(n9136) );
  XNOR U9360 ( .A(n9075), .B(n9079), .Z(n9137) );
  XOR U9361 ( .A(n9071), .B(n9074), .Z(n9138) );
  XOR U9362 ( .A(n9139), .B(n9140), .Z(n9071) );
  XNOR U9363 ( .A(n9141), .B(n9142), .Z(n9140) );
  XNOR U9364 ( .A(n9143), .B(n9144), .Z(n9141) );
  XOR U9365 ( .A(n9145), .B(n9146), .Z(n9144) );
  AND U9366 ( .A(a[9]), .B(b[14]), .Z(n9146) );
  AND U9367 ( .A(a[8]), .B(b[15]), .Z(n9145) );
  XNOR U9368 ( .A(n9147), .B(n9143), .Z(n9139) );
  XOR U9369 ( .A(n9148), .B(n9149), .Z(n9143) );
  NOR U9370 ( .A(n9150), .B(n9151), .Z(n9148) );
  AND U9371 ( .A(a[10]), .B(b[13]), .Z(n9147) );
  XOR U9372 ( .A(n9152), .B(n9069), .Z(n9070) );
  IV U9373 ( .A(n9142), .Z(n9069) );
  XOR U9374 ( .A(n9153), .B(n9154), .Z(n9142) );
  ANDN U9375 ( .B(n9155), .A(n9156), .Z(n9153) );
  AND U9376 ( .A(a[11]), .B(b[12]), .Z(n9152) );
  XOR U9377 ( .A(n9158), .B(n9159), .Z(n9074) );
  ANDN U9378 ( .B(n9160), .A(n9161), .Z(n9158) );
  AND U9379 ( .A(b[11]), .B(a[12]), .Z(n9157) );
  XOR U9380 ( .A(n9163), .B(n9164), .Z(n9079) );
  ANDN U9381 ( .B(n9165), .A(n9166), .Z(n9163) );
  AND U9382 ( .A(a[13]), .B(b[10]), .Z(n9162) );
  XOR U9383 ( .A(n9168), .B(n9169), .Z(n9084) );
  ANDN U9384 ( .B(n9170), .A(n9171), .Z(n9168) );
  AND U9385 ( .A(b[9]), .B(a[14]), .Z(n9167) );
  XOR U9386 ( .A(n9173), .B(n9174), .Z(n9089) );
  ANDN U9387 ( .B(n9101), .A(n9134), .Z(n9173) );
  AND U9388 ( .A(a[15]), .B(b[7]), .Z(n9175) );
  XNOR U9389 ( .A(n9170), .B(n9174), .Z(n9176) );
  XOR U9390 ( .A(n9177), .B(n9178), .Z(n9174) );
  ANDN U9391 ( .B(n9106), .A(n9133), .Z(n9177) );
  AND U9392 ( .A(a[15]), .B(b[6]), .Z(n9179) );
  XNOR U9393 ( .A(n9181), .B(n9178), .Z(n9180) );
  XOR U9394 ( .A(n9182), .B(n9183), .Z(n9178) );
  ANDN U9395 ( .B(n9111), .A(n9132), .Z(n9182) );
  AND U9396 ( .A(a[15]), .B(b[5]), .Z(n9184) );
  XNOR U9397 ( .A(n9186), .B(n9183), .Z(n9185) );
  XOR U9398 ( .A(n9187), .B(n9188), .Z(n9183) );
  ANDN U9399 ( .B(n9116), .A(n9131), .Z(n9187) );
  AND U9400 ( .A(a[15]), .B(b[4]), .Z(n9189) );
  XNOR U9401 ( .A(n9191), .B(n9188), .Z(n9190) );
  XOR U9402 ( .A(n9192), .B(n9193), .Z(n9188) );
  ANDN U9403 ( .B(n9121), .A(n9130), .Z(n9192) );
  AND U9404 ( .A(a[15]), .B(b[3]), .Z(n9194) );
  XNOR U9405 ( .A(n9196), .B(n9193), .Z(n9195) );
  XOR U9406 ( .A(n9197), .B(n9198), .Z(n9193) );
  ANDN U9407 ( .B(n9126), .A(n9127), .Z(n9197) );
  AND U9408 ( .A(b[2]), .B(a[15]), .Z(n9199) );
  XNOR U9409 ( .A(n9201), .B(n9198), .Z(n9200) );
  XOR U9410 ( .A(n9202), .B(n9203), .Z(n9198) );
  NANDN U9411 ( .A(n9129), .B(n9128), .Z(n9203) );
  XOR U9412 ( .A(n9202), .B(n9204), .Z(n9128) );
  NAND U9413 ( .A(a[15]), .B(b[1]), .Z(n9204) );
  XOR U9414 ( .A(n9202), .B(n9206), .Z(n9205) );
  OR U9415 ( .A(n9208), .B(n9209), .Z(n9202) );
  XNOR U9416 ( .A(n9165), .B(n9169), .Z(n9215) );
  XNOR U9417 ( .A(n9160), .B(n9164), .Z(n9216) );
  XNOR U9418 ( .A(n9155), .B(n9159), .Z(n9217) );
  XOR U9419 ( .A(n9151), .B(n9154), .Z(n9218) );
  XOR U9420 ( .A(n9219), .B(n9220), .Z(n9151) );
  XNOR U9421 ( .A(n9221), .B(n9222), .Z(n9220) );
  XOR U9422 ( .A(n9223), .B(n9224), .Z(n9221) );
  AND U9423 ( .A(a[9]), .B(b[13]), .Z(n9223) );
  XOR U9424 ( .A(n9224), .B(n9225), .Z(n9219) );
  XOR U9425 ( .A(n9226), .B(n9227), .Z(n9225) );
  AND U9426 ( .A(a[8]), .B(b[14]), .Z(n9227) );
  AND U9427 ( .A(a[7]), .B(b[15]), .Z(n9226) );
  XOR U9428 ( .A(n9228), .B(n9229), .Z(n9224) );
  ANDN U9429 ( .B(n9230), .A(n9231), .Z(n9228) );
  XOR U9430 ( .A(n9232), .B(n9149), .Z(n9150) );
  IV U9431 ( .A(n9222), .Z(n9149) );
  XOR U9432 ( .A(n9233), .B(n9234), .Z(n9222) );
  NOR U9433 ( .A(n9235), .B(n9236), .Z(n9233) );
  AND U9434 ( .A(a[10]), .B(b[12]), .Z(n9232) );
  XOR U9435 ( .A(n9238), .B(n9239), .Z(n9154) );
  ANDN U9436 ( .B(n9240), .A(n9241), .Z(n9238) );
  AND U9437 ( .A(a[11]), .B(b[11]), .Z(n9237) );
  XOR U9438 ( .A(n9243), .B(n9244), .Z(n9159) );
  ANDN U9439 ( .B(n9245), .A(n9246), .Z(n9243) );
  AND U9440 ( .A(b[10]), .B(a[12]), .Z(n9242) );
  XOR U9441 ( .A(n9248), .B(n9249), .Z(n9164) );
  ANDN U9442 ( .B(n9250), .A(n9251), .Z(n9248) );
  AND U9443 ( .A(a[13]), .B(b[9]), .Z(n9247) );
  XOR U9444 ( .A(n9253), .B(n9254), .Z(n9169) );
  ANDN U9445 ( .B(n9181), .A(n9214), .Z(n9253) );
  AND U9446 ( .A(b[7]), .B(a[14]), .Z(n9255) );
  XNOR U9447 ( .A(n9250), .B(n9254), .Z(n9256) );
  XOR U9448 ( .A(n9257), .B(n9258), .Z(n9254) );
  ANDN U9449 ( .B(n9186), .A(n9213), .Z(n9257) );
  AND U9450 ( .A(b[6]), .B(a[14]), .Z(n9259) );
  XNOR U9451 ( .A(n9261), .B(n9258), .Z(n9260) );
  XOR U9452 ( .A(n9262), .B(n9263), .Z(n9258) );
  ANDN U9453 ( .B(n9191), .A(n9212), .Z(n9262) );
  AND U9454 ( .A(b[5]), .B(a[14]), .Z(n9264) );
  XNOR U9455 ( .A(n9266), .B(n9263), .Z(n9265) );
  XOR U9456 ( .A(n9267), .B(n9268), .Z(n9263) );
  ANDN U9457 ( .B(n9196), .A(n9211), .Z(n9267) );
  AND U9458 ( .A(b[4]), .B(a[14]), .Z(n9269) );
  XNOR U9459 ( .A(n9271), .B(n9268), .Z(n9270) );
  XOR U9460 ( .A(n9272), .B(n9273), .Z(n9268) );
  ANDN U9461 ( .B(n9201), .A(n9210), .Z(n9272) );
  AND U9462 ( .A(b[3]), .B(a[14]), .Z(n9274) );
  XNOR U9463 ( .A(n9276), .B(n9273), .Z(n9275) );
  XOR U9464 ( .A(n9277), .B(n9278), .Z(n9273) );
  ANDN U9465 ( .B(n9206), .A(n9207), .Z(n9277) );
  AND U9466 ( .A(b[2]), .B(a[14]), .Z(n9279) );
  XNOR U9467 ( .A(n9281), .B(n9278), .Z(n9280) );
  XOR U9468 ( .A(n9282), .B(n9283), .Z(n9278) );
  OR U9469 ( .A(n9284), .B(n9285), .Z(n9283) );
  XNOR U9470 ( .A(n9245), .B(n9249), .Z(n9291) );
  XNOR U9471 ( .A(n9240), .B(n9244), .Z(n9292) );
  XOR U9472 ( .A(n9236), .B(n9239), .Z(n9293) );
  XNOR U9473 ( .A(n9231), .B(n9294), .Z(n9236) );
  XNOR U9474 ( .A(n9230), .B(n9234), .Z(n9294) );
  XOR U9475 ( .A(n9295), .B(n9229), .Z(n9230) );
  AND U9476 ( .A(a[9]), .B(b[12]), .Z(n9295) );
  XOR U9477 ( .A(n9296), .B(n9297), .Z(n9231) );
  XOR U9478 ( .A(n9229), .B(n9298), .Z(n9297) );
  XOR U9479 ( .A(n9299), .B(n9300), .Z(n9298) );
  XOR U9480 ( .A(n9301), .B(n9302), .Z(n9300) );
  NAND U9481 ( .A(a[7]), .B(b[14]), .Z(n9302) );
  AND U9482 ( .A(a[6]), .B(b[15]), .Z(n9301) );
  XOR U9483 ( .A(n9303), .B(n9304), .Z(n9229) );
  ANDN U9484 ( .B(n9305), .A(n9306), .Z(n9303) );
  XOR U9485 ( .A(n9307), .B(n9299), .Z(n9296) );
  XOR U9486 ( .A(n9308), .B(n9309), .Z(n9299) );
  NOR U9487 ( .A(n9310), .B(n9311), .Z(n9308) );
  AND U9488 ( .A(a[8]), .B(b[13]), .Z(n9307) );
  XOR U9489 ( .A(n9313), .B(n9314), .Z(n9234) );
  ANDN U9490 ( .B(n9315), .A(n9316), .Z(n9313) );
  AND U9491 ( .A(a[10]), .B(b[11]), .Z(n9312) );
  XOR U9492 ( .A(n9318), .B(n9319), .Z(n9239) );
  ANDN U9493 ( .B(n9320), .A(n9321), .Z(n9318) );
  AND U9494 ( .A(a[11]), .B(b[10]), .Z(n9317) );
  XOR U9495 ( .A(n9323), .B(n9324), .Z(n9244) );
  ANDN U9496 ( .B(n9325), .A(n9326), .Z(n9323) );
  AND U9497 ( .A(b[9]), .B(a[12]), .Z(n9322) );
  XOR U9498 ( .A(n9328), .B(n9329), .Z(n9249) );
  ANDN U9499 ( .B(n9261), .A(n9290), .Z(n9328) );
  AND U9500 ( .A(a[13]), .B(b[7]), .Z(n9330) );
  XNOR U9501 ( .A(n9325), .B(n9329), .Z(n9331) );
  XOR U9502 ( .A(n9332), .B(n9333), .Z(n9329) );
  ANDN U9503 ( .B(n9266), .A(n9289), .Z(n9332) );
  AND U9504 ( .A(a[13]), .B(b[6]), .Z(n9334) );
  XNOR U9505 ( .A(n9336), .B(n9333), .Z(n9335) );
  XOR U9506 ( .A(n9337), .B(n9338), .Z(n9333) );
  ANDN U9507 ( .B(n9271), .A(n9288), .Z(n9337) );
  AND U9508 ( .A(a[13]), .B(b[5]), .Z(n9339) );
  XNOR U9509 ( .A(n9341), .B(n9338), .Z(n9340) );
  XOR U9510 ( .A(n9342), .B(n9343), .Z(n9338) );
  ANDN U9511 ( .B(n9276), .A(n9287), .Z(n9342) );
  AND U9512 ( .A(a[13]), .B(b[4]), .Z(n9344) );
  XNOR U9513 ( .A(n9346), .B(n9343), .Z(n9345) );
  XOR U9514 ( .A(n9347), .B(n9348), .Z(n9343) );
  ANDN U9515 ( .B(n9281), .A(n9286), .Z(n9347) );
  XNOR U9516 ( .A(n9349), .B(n9348), .Z(n9286) );
  AND U9517 ( .A(a[13]), .B(b[3]), .Z(n9349) );
  XNOR U9518 ( .A(n9351), .B(n9348), .Z(n9350) );
  XNOR U9519 ( .A(n9352), .B(n9353), .Z(n9348) );
  NOR U9520 ( .A(n9354), .B(n9355), .Z(n9352) );
  XNOR U9521 ( .A(n9320), .B(n9324), .Z(n9360) );
  XNOR U9522 ( .A(n9315), .B(n9319), .Z(n9361) );
  XNOR U9523 ( .A(n9305), .B(n9314), .Z(n9362) );
  XOR U9524 ( .A(n9363), .B(n9304), .Z(n9305) );
  AND U9525 ( .A(a[9]), .B(b[11]), .Z(n9363) );
  XOR U9526 ( .A(n9304), .B(n9311), .Z(n9364) );
  XOR U9527 ( .A(n9365), .B(n9366), .Z(n9311) );
  XOR U9528 ( .A(n9309), .B(n9367), .Z(n9366) );
  XOR U9529 ( .A(n9368), .B(n9369), .Z(n9367) );
  XOR U9530 ( .A(n9370), .B(n9371), .Z(n9369) );
  NAND U9531 ( .A(a[6]), .B(b[14]), .Z(n9371) );
  AND U9532 ( .A(a[5]), .B(b[15]), .Z(n9370) );
  XOR U9533 ( .A(n9372), .B(n9368), .Z(n9365) );
  XOR U9534 ( .A(n9373), .B(n9374), .Z(n9368) );
  NOR U9535 ( .A(n9375), .B(n9376), .Z(n9373) );
  AND U9536 ( .A(a[7]), .B(b[13]), .Z(n9372) );
  XOR U9537 ( .A(n9377), .B(n9378), .Z(n9304) );
  ANDN U9538 ( .B(n9379), .A(n9380), .Z(n9377) );
  XNOR U9539 ( .A(n9381), .B(n9309), .Z(n9310) );
  XOR U9540 ( .A(n9382), .B(n9383), .Z(n9309) );
  ANDN U9541 ( .B(n9384), .A(n9385), .Z(n9382) );
  AND U9542 ( .A(a[8]), .B(b[12]), .Z(n9381) );
  XOR U9543 ( .A(n9387), .B(n9388), .Z(n9314) );
  ANDN U9544 ( .B(n9389), .A(n9390), .Z(n9387) );
  AND U9545 ( .A(b[10]), .B(a[10]), .Z(n9386) );
  XOR U9546 ( .A(n9392), .B(n9393), .Z(n9319) );
  ANDN U9547 ( .B(n9394), .A(n9395), .Z(n9392) );
  AND U9548 ( .A(a[11]), .B(b[9]), .Z(n9391) );
  XOR U9549 ( .A(n9397), .B(n9398), .Z(n9324) );
  ANDN U9550 ( .B(n9336), .A(n9359), .Z(n9397) );
  AND U9551 ( .A(b[7]), .B(a[12]), .Z(n9399) );
  XNOR U9552 ( .A(n9394), .B(n9398), .Z(n9400) );
  XOR U9553 ( .A(n9401), .B(n9402), .Z(n9398) );
  ANDN U9554 ( .B(n9341), .A(n9358), .Z(n9401) );
  AND U9555 ( .A(b[6]), .B(a[12]), .Z(n9403) );
  XNOR U9556 ( .A(n9405), .B(n9402), .Z(n9404) );
  XOR U9557 ( .A(n9406), .B(n9407), .Z(n9402) );
  ANDN U9558 ( .B(n9346), .A(n9357), .Z(n9406) );
  AND U9559 ( .A(b[5]), .B(a[12]), .Z(n9408) );
  XNOR U9560 ( .A(n9410), .B(n9407), .Z(n9409) );
  XOR U9561 ( .A(n9411), .B(n9412), .Z(n9407) );
  ANDN U9562 ( .B(n9351), .A(n9356), .Z(n9411) );
  XNOR U9563 ( .A(n9413), .B(n9412), .Z(n9356) );
  AND U9564 ( .A(b[4]), .B(a[12]), .Z(n9413) );
  XNOR U9565 ( .A(n9415), .B(n9412), .Z(n9414) );
  XOR U9566 ( .A(n9416), .B(n9417), .Z(n9412) );
  ANDN U9567 ( .B(n9418), .A(n9419), .Z(n9416) );
  XNOR U9568 ( .A(n9389), .B(n9393), .Z(n9423) );
  XNOR U9569 ( .A(n9379), .B(n9388), .Z(n9424) );
  XOR U9570 ( .A(n9425), .B(n9378), .Z(n9379) );
  AND U9571 ( .A(a[9]), .B(b[10]), .Z(n9425) );
  XNOR U9572 ( .A(n9378), .B(n9384), .Z(n9426) );
  XOR U9573 ( .A(n9383), .B(n9376), .Z(n9427) );
  XOR U9574 ( .A(n9428), .B(n9429), .Z(n9376) );
  XOR U9575 ( .A(n9374), .B(n9430), .Z(n9429) );
  XOR U9576 ( .A(n9431), .B(n9432), .Z(n9430) );
  XOR U9577 ( .A(n9433), .B(n9434), .Z(n9432) );
  NAND U9578 ( .A(a[5]), .B(b[14]), .Z(n9434) );
  AND U9579 ( .A(a[4]), .B(b[15]), .Z(n9433) );
  XOR U9580 ( .A(n9435), .B(n9431), .Z(n9428) );
  XOR U9581 ( .A(n9436), .B(n9437), .Z(n9431) );
  NOR U9582 ( .A(n9438), .B(n9439), .Z(n9436) );
  AND U9583 ( .A(a[6]), .B(b[13]), .Z(n9435) );
  XNOR U9584 ( .A(n9440), .B(n9374), .Z(n9375) );
  XOR U9585 ( .A(n9441), .B(n9442), .Z(n9374) );
  ANDN U9586 ( .B(n9443), .A(n9444), .Z(n9441) );
  AND U9587 ( .A(a[7]), .B(b[12]), .Z(n9440) );
  XOR U9588 ( .A(n9445), .B(n9446), .Z(n9378) );
  ANDN U9589 ( .B(n9447), .A(n9448), .Z(n9445) );
  XNOR U9590 ( .A(n9449), .B(n9383), .Z(n9385) );
  XOR U9591 ( .A(n9450), .B(n9451), .Z(n9383) );
  ANDN U9592 ( .B(n9452), .A(n9453), .Z(n9450) );
  AND U9593 ( .A(a[8]), .B(b[11]), .Z(n9449) );
  XOR U9594 ( .A(n9455), .B(n9456), .Z(n9388) );
  ANDN U9595 ( .B(n9457), .A(n9458), .Z(n9455) );
  AND U9596 ( .A(b[9]), .B(a[10]), .Z(n9454) );
  XOR U9597 ( .A(n9460), .B(n9461), .Z(n9393) );
  ANDN U9598 ( .B(n9405), .A(n9422), .Z(n9460) );
  AND U9599 ( .A(a[11]), .B(b[7]), .Z(n9462) );
  XNOR U9600 ( .A(n9457), .B(n9461), .Z(n9463) );
  XOR U9601 ( .A(n9464), .B(n9465), .Z(n9461) );
  ANDN U9602 ( .B(n9410), .A(n9421), .Z(n9464) );
  AND U9603 ( .A(a[11]), .B(b[6]), .Z(n9466) );
  XNOR U9604 ( .A(n9468), .B(n9465), .Z(n9467) );
  XOR U9605 ( .A(n9469), .B(n9470), .Z(n9465) );
  ANDN U9606 ( .B(n9415), .A(n9420), .Z(n9469) );
  XNOR U9607 ( .A(n9471), .B(n9470), .Z(n9420) );
  AND U9608 ( .A(a[11]), .B(b[5]), .Z(n9471) );
  XNOR U9609 ( .A(n9473), .B(n9470), .Z(n9472) );
  XOR U9610 ( .A(n9474), .B(n9475), .Z(n9470) );
  ANDN U9611 ( .B(n9476), .A(n9477), .Z(n9474) );
  XNOR U9612 ( .A(n9447), .B(n9456), .Z(n9480) );
  XOR U9613 ( .A(n9481), .B(n9446), .Z(n9447) );
  AND U9614 ( .A(a[9]), .B(b[9]), .Z(n9481) );
  XNOR U9615 ( .A(n9446), .B(n9452), .Z(n9482) );
  XNOR U9616 ( .A(n9451), .B(n9443), .Z(n9483) );
  XOR U9617 ( .A(n9442), .B(n9439), .Z(n9484) );
  XOR U9618 ( .A(n9485), .B(n9486), .Z(n9439) );
  XOR U9619 ( .A(n9437), .B(n9487), .Z(n9486) );
  XOR U9620 ( .A(n9488), .B(n9489), .Z(n9487) );
  XOR U9621 ( .A(n9490), .B(n9491), .Z(n9489) );
  NAND U9622 ( .A(a[4]), .B(b[14]), .Z(n9491) );
  AND U9623 ( .A(a[3]), .B(b[15]), .Z(n9490) );
  XOR U9624 ( .A(n9492), .B(n9488), .Z(n9485) );
  XOR U9625 ( .A(n9493), .B(n9494), .Z(n9488) );
  NOR U9626 ( .A(n9495), .B(n9496), .Z(n9493) );
  AND U9627 ( .A(a[5]), .B(b[13]), .Z(n9492) );
  XNOR U9628 ( .A(n9497), .B(n9437), .Z(n9438) );
  XOR U9629 ( .A(n9498), .B(n9499), .Z(n9437) );
  ANDN U9630 ( .B(n9500), .A(n9501), .Z(n9498) );
  AND U9631 ( .A(a[6]), .B(b[12]), .Z(n9497) );
  XNOR U9632 ( .A(n9502), .B(n9442), .Z(n9444) );
  XOR U9633 ( .A(n9503), .B(n9504), .Z(n9442) );
  ANDN U9634 ( .B(n9505), .A(n9506), .Z(n9503) );
  AND U9635 ( .A(a[7]), .B(b[11]), .Z(n9502) );
  XOR U9636 ( .A(n9507), .B(n9508), .Z(n9446) );
  ANDN U9637 ( .B(n9509), .A(n9510), .Z(n9507) );
  XNOR U9638 ( .A(n9511), .B(n9451), .Z(n9453) );
  XOR U9639 ( .A(n9512), .B(n9513), .Z(n9451) );
  ANDN U9640 ( .B(n9514), .A(n9515), .Z(n9512) );
  AND U9641 ( .A(a[8]), .B(b[10]), .Z(n9511) );
  XOR U9642 ( .A(n9517), .B(n9518), .Z(n9456) );
  ANDN U9643 ( .B(n9468), .A(n9479), .Z(n9517) );
  AND U9644 ( .A(b[7]), .B(a[10]), .Z(n9519) );
  XNOR U9645 ( .A(n9509), .B(n9518), .Z(n9520) );
  XOR U9646 ( .A(n9521), .B(n9522), .Z(n9518) );
  ANDN U9647 ( .B(n9473), .A(n9478), .Z(n9521) );
  XNOR U9648 ( .A(n9523), .B(n9522), .Z(n9478) );
  AND U9649 ( .A(b[6]), .B(a[10]), .Z(n9523) );
  XNOR U9650 ( .A(n9525), .B(n9522), .Z(n9524) );
  XOR U9651 ( .A(n9526), .B(n9527), .Z(n9522) );
  ANDN U9652 ( .B(n9528), .A(n9529), .Z(n9526) );
  XOR U9653 ( .A(n9531), .B(n9508), .Z(n9509) );
  AND U9654 ( .A(a[9]), .B(b[8]), .Z(n9531) );
  XNOR U9655 ( .A(n9508), .B(n9514), .Z(n9532) );
  XNOR U9656 ( .A(n9513), .B(n9505), .Z(n9533) );
  XNOR U9657 ( .A(n9504), .B(n9500), .Z(n9534) );
  XOR U9658 ( .A(n9499), .B(n9496), .Z(n9535) );
  XOR U9659 ( .A(n9536), .B(n9537), .Z(n9496) );
  XOR U9660 ( .A(n9494), .B(n9538), .Z(n9537) );
  XOR U9661 ( .A(n9539), .B(n9540), .Z(n9538) );
  XOR U9662 ( .A(n9541), .B(n9542), .Z(n9540) );
  NAND U9663 ( .A(a[3]), .B(b[14]), .Z(n9542) );
  AND U9664 ( .A(a[2]), .B(b[15]), .Z(n9541) );
  XOR U9665 ( .A(n9543), .B(n9539), .Z(n9536) );
  XOR U9666 ( .A(n9544), .B(n9545), .Z(n9539) );
  NOR U9667 ( .A(n9546), .B(n9547), .Z(n9544) );
  AND U9668 ( .A(a[4]), .B(b[13]), .Z(n9543) );
  XNOR U9669 ( .A(n9548), .B(n9494), .Z(n9495) );
  XOR U9670 ( .A(n9549), .B(n9550), .Z(n9494) );
  ANDN U9671 ( .B(n9551), .A(n9552), .Z(n9549) );
  AND U9672 ( .A(a[5]), .B(b[12]), .Z(n9548) );
  XNOR U9673 ( .A(n9553), .B(n9499), .Z(n9501) );
  XOR U9674 ( .A(n9554), .B(n9555), .Z(n9499) );
  ANDN U9675 ( .B(n9556), .A(n9557), .Z(n9554) );
  AND U9676 ( .A(a[6]), .B(b[11]), .Z(n9553) );
  XNOR U9677 ( .A(n9558), .B(n9504), .Z(n9506) );
  XOR U9678 ( .A(n9559), .B(n9560), .Z(n9504) );
  ANDN U9679 ( .B(n9561), .A(n9562), .Z(n9559) );
  AND U9680 ( .A(a[7]), .B(b[10]), .Z(n9558) );
  XOR U9681 ( .A(n9563), .B(n9564), .Z(n9508) );
  ANDN U9682 ( .B(n9525), .A(n9530), .Z(n9563) );
  XNOR U9683 ( .A(n9564), .B(n9566), .Z(n9565) );
  XOR U9684 ( .A(n9568), .B(n9564), .Z(n9525) );
  XOR U9685 ( .A(n9569), .B(n9570), .Z(n9564) );
  ANDN U9686 ( .B(n9571), .A(n9572), .Z(n9569) );
  AND U9687 ( .A(a[9]), .B(b[7]), .Z(n9568) );
  XNOR U9688 ( .A(n9573), .B(n9513), .Z(n9515) );
  XOR U9689 ( .A(n9574), .B(n9575), .Z(n9513) );
  ANDN U9690 ( .B(n9566), .A(n9567), .Z(n9574) );
  XNOR U9691 ( .A(n9576), .B(n9575), .Z(n9567) );
  AND U9692 ( .A(b[8]), .B(a[8]), .Z(n9576) );
  XNOR U9693 ( .A(n9575), .B(n9561), .Z(n9577) );
  XNOR U9694 ( .A(n9560), .B(n9556), .Z(n9578) );
  XNOR U9695 ( .A(n9555), .B(n9551), .Z(n9579) );
  XOR U9696 ( .A(n9550), .B(n9547), .Z(n9580) );
  XOR U9697 ( .A(n9581), .B(n9582), .Z(n9547) );
  XOR U9698 ( .A(n9545), .B(n9583), .Z(n9582) );
  XOR U9699 ( .A(n9584), .B(n9585), .Z(n9583) );
  XOR U9700 ( .A(n9586), .B(n9587), .Z(n9585) );
  NAND U9701 ( .A(a[2]), .B(b[14]), .Z(n9587) );
  AND U9702 ( .A(a[1]), .B(b[15]), .Z(n9586) );
  XOR U9703 ( .A(n9588), .B(n9584), .Z(n9581) );
  XOR U9704 ( .A(n9589), .B(n9590), .Z(n9584) );
  NOR U9705 ( .A(n9591), .B(n9592), .Z(n9589) );
  AND U9706 ( .A(a[3]), .B(b[13]), .Z(n9588) );
  XNOR U9707 ( .A(n9593), .B(n9545), .Z(n9546) );
  XOR U9708 ( .A(n9594), .B(n9595), .Z(n9545) );
  ANDN U9709 ( .B(n9596), .A(n9597), .Z(n9594) );
  AND U9710 ( .A(a[4]), .B(b[12]), .Z(n9593) );
  XNOR U9711 ( .A(n9598), .B(n9550), .Z(n9552) );
  XOR U9712 ( .A(n9599), .B(n9600), .Z(n9550) );
  ANDN U9713 ( .B(n9601), .A(n9602), .Z(n9599) );
  AND U9714 ( .A(a[5]), .B(b[11]), .Z(n9598) );
  XNOR U9715 ( .A(n9603), .B(n9555), .Z(n9557) );
  XOR U9716 ( .A(n9604), .B(n9605), .Z(n9555) );
  ANDN U9717 ( .B(n9606), .A(n9607), .Z(n9604) );
  AND U9718 ( .A(a[6]), .B(b[10]), .Z(n9603) );
  XOR U9719 ( .A(n9608), .B(n9609), .Z(n9575) );
  ANDN U9720 ( .B(n9610), .A(n9611), .Z(n9608) );
  XNOR U9721 ( .A(n9612), .B(n9560), .Z(n9562) );
  XOR U9722 ( .A(n9613), .B(n9614), .Z(n9560) );
  ANDN U9723 ( .B(n9615), .A(n9616), .Z(n9613) );
  AND U9724 ( .A(a[7]), .B(b[9]), .Z(n9612) );
  AND U9725 ( .A(a[8]), .B(b[9]), .Z(n9573) );
  AND U9726 ( .A(b[8]), .B(a[10]), .Z(n9516) );
  AND U9727 ( .A(a[11]), .B(b[8]), .Z(n9459) );
  AND U9728 ( .A(b[8]), .B(a[12]), .Z(n9396) );
  AND U9729 ( .A(a[13]), .B(b[8]), .Z(n9327) );
  AND U9730 ( .A(b[8]), .B(a[14]), .Z(n9252) );
  AND U9731 ( .A(a[15]), .B(b[8]), .Z(n9172) );
  AND U9732 ( .A(a[16]), .B(b[8]), .Z(n9092) );
  AND U9733 ( .A(a[17]), .B(b[8]), .Z(n9007) );
  AND U9734 ( .A(a[18]), .B(b[8]), .Z(n8927) );
  AND U9735 ( .A(a[19]), .B(b[8]), .Z(n8847) );
  AND U9736 ( .A(a[20]), .B(b[8]), .Z(n8767) );
  AND U9737 ( .A(a[21]), .B(b[8]), .Z(n8687) );
  AND U9738 ( .A(a[22]), .B(b[8]), .Z(n8607) );
  AND U9739 ( .A(a[23]), .B(b[8]), .Z(n8528) );
  AND U9740 ( .A(a[25]), .B(b[7]), .Z(n8415) );
  AND U9741 ( .A(a[26]), .B(b[7]), .Z(n8336) );
  AND U9742 ( .A(a[27]), .B(b[7]), .Z(n8257) );
  AND U9743 ( .A(a[28]), .B(b[7]), .Z(n8178) );
  AND U9744 ( .A(a[29]), .B(b[7]), .Z(n8099) );
  AND U9745 ( .A(a[30]), .B(b[7]), .Z(n8020) );
  AND U9746 ( .A(a[31]), .B(b[7]), .Z(n7940) );
  AND U9747 ( .A(a[32]), .B(b[7]), .Z(n7860) );
  AND U9748 ( .A(a[33]), .B(b[7]), .Z(n7774) );
  AND U9749 ( .A(a[34]), .B(b[7]), .Z(n7694) );
  AND U9750 ( .A(a[35]), .B(b[7]), .Z(n7614) );
  AND U9751 ( .A(a[36]), .B(b[7]), .Z(n7534) );
  AND U9752 ( .A(a[37]), .B(b[7]), .Z(n7454) );
  AND U9753 ( .A(a[38]), .B(b[7]), .Z(n7375) );
  AND U9754 ( .A(a[40]), .B(b[6]), .Z(n7268) );
  AND U9755 ( .A(a[41]), .B(b[6]), .Z(n7189) );
  AND U9756 ( .A(a[42]), .B(b[6]), .Z(n7110) );
  AND U9757 ( .A(a[43]), .B(b[6]), .Z(n7031) );
  AND U9758 ( .A(a[44]), .B(b[6]), .Z(n6952) );
  AND U9759 ( .A(a[45]), .B(b[6]), .Z(n6873) );
  AND U9760 ( .A(a[46]), .B(b[6]), .Z(n6794) );
  AND U9761 ( .A(a[47]), .B(b[6]), .Z(n6714) );
  AND U9762 ( .A(a[48]), .B(b[6]), .Z(n6634) );
  AND U9763 ( .A(a[49]), .B(b[6]), .Z(n6547) );
  AND U9764 ( .A(a[50]), .B(b[6]), .Z(n6467) );
  AND U9765 ( .A(a[51]), .B(b[6]), .Z(n6387) );
  AND U9766 ( .A(a[52]), .B(b[6]), .Z(n6307) );
  AND U9767 ( .A(a[53]), .B(b[6]), .Z(n6228) );
  AND U9768 ( .A(a[55]), .B(b[5]), .Z(n6127) );
  AND U9769 ( .A(a[56]), .B(b[5]), .Z(n6048) );
  AND U9770 ( .A(a[57]), .B(b[5]), .Z(n5969) );
  AND U9771 ( .A(a[58]), .B(b[5]), .Z(n5890) );
  AND U9772 ( .A(a[59]), .B(b[5]), .Z(n5811) );
  AND U9773 ( .A(a[60]), .B(b[5]), .Z(n5732) );
  AND U9774 ( .A(a[61]), .B(b[5]), .Z(n5653) );
  AND U9775 ( .A(a[62]), .B(b[5]), .Z(n5574) );
  AND U9776 ( .A(a[63]), .B(b[5]), .Z(n5494) );
  AND U9777 ( .A(a[64]), .B(b[5]), .Z(n5414) );
  AND U9778 ( .A(a[65]), .B(b[5]), .Z(n5326) );
  AND U9779 ( .A(a[66]), .B(b[5]), .Z(n5246) );
  AND U9780 ( .A(a[67]), .B(b[5]), .Z(n5166) );
  AND U9781 ( .A(a[68]), .B(b[5]), .Z(n5087) );
  AND U9782 ( .A(a[70]), .B(b[4]), .Z(n4992) );
  AND U9783 ( .A(a[71]), .B(b[4]), .Z(n4913) );
  AND U9784 ( .A(a[72]), .B(b[4]), .Z(n4834) );
  AND U9785 ( .A(a[73]), .B(b[4]), .Z(n4755) );
  AND U9786 ( .A(a[74]), .B(b[4]), .Z(n4676) );
  AND U9787 ( .A(a[75]), .B(b[4]), .Z(n4597) );
  AND U9788 ( .A(a[76]), .B(b[4]), .Z(n4518) );
  AND U9789 ( .A(a[77]), .B(b[4]), .Z(n4439) );
  AND U9790 ( .A(a[78]), .B(b[4]), .Z(n4360) );
  AND U9791 ( .A(a[79]), .B(b[4]), .Z(n4280) );
  AND U9792 ( .A(a[80]), .B(b[4]), .Z(n4200) );
  AND U9793 ( .A(a[81]), .B(b[4]), .Z(n4111) );
  AND U9794 ( .A(a[82]), .B(b[4]), .Z(n4031) );
  AND U9795 ( .A(a[83]), .B(b[4]), .Z(n3952) );
  AND U9796 ( .A(a[85]), .B(b[3]), .Z(n3863) );
  AND U9797 ( .A(a[86]), .B(b[3]), .Z(n3784) );
  AND U9798 ( .A(a[87]), .B(b[3]), .Z(n3705) );
  AND U9799 ( .A(a[88]), .B(b[3]), .Z(n3626) );
  AND U9800 ( .A(a[89]), .B(b[3]), .Z(n3547) );
  AND U9801 ( .A(a[90]), .B(b[3]), .Z(n3468) );
  AND U9802 ( .A(a[91]), .B(b[3]), .Z(n3389) );
  AND U9803 ( .A(a[92]), .B(b[3]), .Z(n3310) );
  AND U9804 ( .A(a[93]), .B(b[3]), .Z(n3231) );
  AND U9805 ( .A(a[94]), .B(b[3]), .Z(n3152) );
  AND U9806 ( .A(a[95]), .B(b[3]), .Z(n3072) );
  AND U9807 ( .A(a[96]), .B(b[3]), .Z(n2992) );
  AND U9808 ( .A(a[97]), .B(b[3]), .Z(n2902) );
  XNOR U9809 ( .A(n2820), .B(n2821), .Z(c[127]) );
  XOR U9810 ( .A(sreg[143]), .B(n2819), .Z(n2821) );
  XOR U9811 ( .A(n9209), .B(n9617), .Z(n2820) );
  XNOR U9812 ( .A(n9208), .B(n2819), .Z(n9617) );
  XOR U9813 ( .A(n9618), .B(n9619), .Z(n2819) );
  ANDN U9814 ( .B(n9620), .A(n9621), .Z(n9618) );
  NANDN U9815 ( .A(n179), .B(a[15]), .Z(n9208) );
  XNOR U9816 ( .A(n9282), .B(n9622), .Z(n9284) );
  NAND U9817 ( .A(b[1]), .B(a[14]), .Z(n9622) );
  XNOR U9818 ( .A(n9282), .B(n9355), .Z(n9623) );
  XOR U9819 ( .A(n9624), .B(n9353), .Z(n9355) );
  AND U9820 ( .A(b[2]), .B(a[13]), .Z(n9624) );
  OR U9821 ( .A(n9625), .B(n9626), .Z(n9282) );
  XOR U9822 ( .A(n9353), .B(n9418), .Z(n9627) );
  XNOR U9823 ( .A(n9417), .B(n9476), .Z(n9628) );
  XNOR U9824 ( .A(n9475), .B(n9528), .Z(n9629) );
  XNOR U9825 ( .A(n9527), .B(n9571), .Z(n9630) );
  XNOR U9826 ( .A(n9570), .B(n9610), .Z(n9631) );
  XNOR U9827 ( .A(n9609), .B(n9615), .Z(n9632) );
  XNOR U9828 ( .A(n9614), .B(n9606), .Z(n9633) );
  XNOR U9829 ( .A(n9605), .B(n9601), .Z(n9634) );
  XNOR U9830 ( .A(n9600), .B(n9596), .Z(n9635) );
  XOR U9831 ( .A(n9595), .B(n9592), .Z(n9636) );
  XOR U9832 ( .A(n9637), .B(n9638), .Z(n9592) );
  XOR U9833 ( .A(n9590), .B(n9639), .Z(n9638) );
  XOR U9834 ( .A(n9640), .B(n9641), .Z(n9639) );
  XOR U9835 ( .A(n9642), .B(n9643), .Z(n9641) );
  NAND U9836 ( .A(a[1]), .B(b[14]), .Z(n9643) );
  AND U9837 ( .A(a[0]), .B(b[15]), .Z(n9642) );
  XOR U9838 ( .A(n9644), .B(n9640), .Z(n9637) );
  XOR U9839 ( .A(n9645), .B(n9646), .Z(n9640) );
  NOR U9840 ( .A(n9647), .B(n9648), .Z(n9645) );
  AND U9841 ( .A(a[2]), .B(b[13]), .Z(n9644) );
  XNOR U9842 ( .A(n9649), .B(n9590), .Z(n9591) );
  XOR U9843 ( .A(n9650), .B(n9651), .Z(n9590) );
  ANDN U9844 ( .B(n9652), .A(n9653), .Z(n9650) );
  AND U9845 ( .A(a[3]), .B(b[12]), .Z(n9649) );
  XNOR U9846 ( .A(n9654), .B(n9595), .Z(n9597) );
  XOR U9847 ( .A(n9655), .B(n9656), .Z(n9595) );
  ANDN U9848 ( .B(n9657), .A(n9658), .Z(n9655) );
  AND U9849 ( .A(a[4]), .B(b[11]), .Z(n9654) );
  XNOR U9850 ( .A(n9659), .B(n9600), .Z(n9602) );
  XOR U9851 ( .A(n9660), .B(n9661), .Z(n9600) );
  ANDN U9852 ( .B(n9662), .A(n9663), .Z(n9660) );
  AND U9853 ( .A(a[5]), .B(b[10]), .Z(n9659) );
  XNOR U9854 ( .A(n9664), .B(n9605), .Z(n9607) );
  XOR U9855 ( .A(n9665), .B(n9666), .Z(n9605) );
  ANDN U9856 ( .B(n9667), .A(n9668), .Z(n9665) );
  AND U9857 ( .A(a[6]), .B(b[9]), .Z(n9664) );
  XNOR U9858 ( .A(n9669), .B(n9614), .Z(n9616) );
  XOR U9859 ( .A(n9670), .B(n9671), .Z(n9614) );
  ANDN U9860 ( .B(n9672), .A(n9673), .Z(n9670) );
  AND U9861 ( .A(a[7]), .B(b[8]), .Z(n9669) );
  XNOR U9862 ( .A(n9674), .B(n9609), .Z(n9611) );
  XOR U9863 ( .A(n9675), .B(n9676), .Z(n9609) );
  ANDN U9864 ( .B(n9677), .A(n9678), .Z(n9675) );
  AND U9865 ( .A(b[7]), .B(a[8]), .Z(n9674) );
  XNOR U9866 ( .A(n9679), .B(n9570), .Z(n9572) );
  XOR U9867 ( .A(n9680), .B(n9681), .Z(n9570) );
  ANDN U9868 ( .B(n9682), .A(n9683), .Z(n9680) );
  AND U9869 ( .A(a[9]), .B(b[6]), .Z(n9679) );
  XNOR U9870 ( .A(n9684), .B(n9527), .Z(n9529) );
  XOR U9871 ( .A(n9685), .B(n9686), .Z(n9527) );
  ANDN U9872 ( .B(n9687), .A(n9688), .Z(n9685) );
  AND U9873 ( .A(b[5]), .B(a[10]), .Z(n9684) );
  XNOR U9874 ( .A(n9689), .B(n9475), .Z(n9477) );
  XOR U9875 ( .A(n9690), .B(n9691), .Z(n9475) );
  ANDN U9876 ( .B(n9692), .A(n9693), .Z(n9690) );
  AND U9877 ( .A(a[11]), .B(b[4]), .Z(n9689) );
  XNOR U9878 ( .A(n9694), .B(n9695), .Z(n9353) );
  OR U9879 ( .A(n9696), .B(n9697), .Z(n9695) );
  XNOR U9880 ( .A(n9698), .B(n9417), .Z(n9419) );
  XNOR U9881 ( .A(n9699), .B(n9700), .Z(n9417) );
  NOR U9882 ( .A(n9701), .B(n9702), .Z(n9699) );
  AND U9883 ( .A(b[3]), .B(a[12]), .Z(n9698) );
  XNOR U9884 ( .A(n9620), .B(n9621), .Z(c[126]) );
  XOR U9885 ( .A(sreg[142]), .B(n9619), .Z(n9621) );
  XOR U9886 ( .A(n9626), .B(n9703), .Z(n9620) );
  XNOR U9887 ( .A(n9625), .B(n9619), .Z(n9703) );
  XOR U9888 ( .A(n9704), .B(n9705), .Z(n9619) );
  ANDN U9889 ( .B(n9706), .A(n9707), .Z(n9704) );
  NANDN U9890 ( .A(n179), .B(a[14]), .Z(n9625) );
  XNOR U9891 ( .A(n9694), .B(n9708), .Z(n9696) );
  NAND U9892 ( .A(a[13]), .B(b[1]), .Z(n9708) );
  XNOR U9893 ( .A(n9694), .B(n9702), .Z(n9709) );
  XOR U9894 ( .A(n9710), .B(n9700), .Z(n9702) );
  AND U9895 ( .A(b[2]), .B(a[12]), .Z(n9710) );
  OR U9896 ( .A(n9711), .B(n9712), .Z(n9694) );
  XOR U9897 ( .A(n9700), .B(n9692), .Z(n9713) );
  XNOR U9898 ( .A(n9691), .B(n9687), .Z(n9714) );
  XNOR U9899 ( .A(n9686), .B(n9682), .Z(n9715) );
  XNOR U9900 ( .A(n9681), .B(n9677), .Z(n9716) );
  XNOR U9901 ( .A(n9676), .B(n9672), .Z(n9717) );
  XNOR U9902 ( .A(n9671), .B(n9667), .Z(n9718) );
  XNOR U9903 ( .A(n9666), .B(n9662), .Z(n9719) );
  XNOR U9904 ( .A(n9661), .B(n9657), .Z(n9720) );
  XNOR U9905 ( .A(n9656), .B(n9652), .Z(n9721) );
  XOR U9906 ( .A(n9651), .B(n9648), .Z(n9722) );
  XOR U9907 ( .A(n9723), .B(n9724), .Z(n9648) );
  XOR U9908 ( .A(n9646), .B(n9725), .Z(n9724) );
  XOR U9909 ( .A(n9726), .B(n9727), .Z(n9725) );
  AND U9910 ( .A(a[0]), .B(b[14]), .Z(n9726) );
  XNOR U9911 ( .A(n9728), .B(n9727), .Z(n9723) );
  XNOR U9912 ( .A(n9729), .B(n9730), .Z(n9727) );
  ANDN U9913 ( .B(n9731), .A(n9732), .Z(n9729) );
  AND U9914 ( .A(a[1]), .B(b[13]), .Z(n9728) );
  XNOR U9915 ( .A(n9733), .B(n9646), .Z(n9647) );
  XOR U9916 ( .A(n9734), .B(n9735), .Z(n9646) );
  ANDN U9917 ( .B(n9736), .A(n9737), .Z(n9734) );
  AND U9918 ( .A(a[2]), .B(b[12]), .Z(n9733) );
  XNOR U9919 ( .A(n9738), .B(n9651), .Z(n9653) );
  XOR U9920 ( .A(n9739), .B(n9740), .Z(n9651) );
  ANDN U9921 ( .B(n9741), .A(n9742), .Z(n9739) );
  AND U9922 ( .A(a[3]), .B(b[11]), .Z(n9738) );
  XNOR U9923 ( .A(n9743), .B(n9656), .Z(n9658) );
  XOR U9924 ( .A(n9744), .B(n9745), .Z(n9656) );
  ANDN U9925 ( .B(n9746), .A(n9747), .Z(n9744) );
  AND U9926 ( .A(a[4]), .B(b[10]), .Z(n9743) );
  XNOR U9927 ( .A(n9748), .B(n9661), .Z(n9663) );
  XOR U9928 ( .A(n9749), .B(n9750), .Z(n9661) );
  ANDN U9929 ( .B(n9751), .A(n9752), .Z(n9749) );
  AND U9930 ( .A(a[5]), .B(b[9]), .Z(n9748) );
  XNOR U9931 ( .A(n9753), .B(n9666), .Z(n9668) );
  XOR U9932 ( .A(n9754), .B(n9755), .Z(n9666) );
  ANDN U9933 ( .B(n9756), .A(n9757), .Z(n9754) );
  AND U9934 ( .A(a[6]), .B(b[8]), .Z(n9753) );
  XNOR U9935 ( .A(n9758), .B(n9671), .Z(n9673) );
  XOR U9936 ( .A(n9759), .B(n9760), .Z(n9671) );
  ANDN U9937 ( .B(n9761), .A(n9762), .Z(n9759) );
  AND U9938 ( .A(a[7]), .B(b[7]), .Z(n9758) );
  XNOR U9939 ( .A(n9763), .B(n9676), .Z(n9678) );
  XOR U9940 ( .A(n9764), .B(n9765), .Z(n9676) );
  ANDN U9941 ( .B(n9766), .A(n9767), .Z(n9764) );
  AND U9942 ( .A(b[6]), .B(a[8]), .Z(n9763) );
  XNOR U9943 ( .A(n9768), .B(n9681), .Z(n9683) );
  XOR U9944 ( .A(n9769), .B(n9770), .Z(n9681) );
  ANDN U9945 ( .B(n9771), .A(n9772), .Z(n9769) );
  AND U9946 ( .A(a[9]), .B(b[5]), .Z(n9768) );
  XNOR U9947 ( .A(n9773), .B(n9686), .Z(n9688) );
  XOR U9948 ( .A(n9774), .B(n9775), .Z(n9686) );
  ANDN U9949 ( .B(n9776), .A(n9777), .Z(n9774) );
  AND U9950 ( .A(b[4]), .B(a[10]), .Z(n9773) );
  XNOR U9951 ( .A(n9778), .B(n9779), .Z(n9700) );
  OR U9952 ( .A(n9780), .B(n9781), .Z(n9779) );
  XNOR U9953 ( .A(n9782), .B(n9691), .Z(n9693) );
  XNOR U9954 ( .A(n9783), .B(n9784), .Z(n9691) );
  NOR U9955 ( .A(n9785), .B(n9786), .Z(n9783) );
  AND U9956 ( .A(a[11]), .B(b[3]), .Z(n9782) );
  XNOR U9957 ( .A(n9706), .B(n9707), .Z(c[125]) );
  XOR U9958 ( .A(sreg[141]), .B(n9705), .Z(n9707) );
  XOR U9959 ( .A(n9712), .B(n9787), .Z(n9706) );
  XNOR U9960 ( .A(n9711), .B(n9705), .Z(n9787) );
  XOR U9961 ( .A(n9788), .B(n9789), .Z(n9705) );
  ANDN U9962 ( .B(n9790), .A(n9791), .Z(n9788) );
  NANDN U9963 ( .A(n179), .B(a[13]), .Z(n9711) );
  XNOR U9964 ( .A(n9778), .B(n9792), .Z(n9780) );
  NAND U9965 ( .A(b[1]), .B(a[12]), .Z(n9792) );
  XNOR U9966 ( .A(n9778), .B(n9786), .Z(n9793) );
  XOR U9967 ( .A(n9794), .B(n9784), .Z(n9786) );
  AND U9968 ( .A(b[2]), .B(a[11]), .Z(n9794) );
  OR U9969 ( .A(n9795), .B(n9796), .Z(n9778) );
  XOR U9970 ( .A(n9784), .B(n9776), .Z(n9797) );
  XNOR U9971 ( .A(n9775), .B(n9771), .Z(n9798) );
  XNOR U9972 ( .A(n9770), .B(n9766), .Z(n9799) );
  XNOR U9973 ( .A(n9765), .B(n9761), .Z(n9800) );
  XNOR U9974 ( .A(n9760), .B(n9756), .Z(n9801) );
  XNOR U9975 ( .A(n9755), .B(n9751), .Z(n9802) );
  XNOR U9976 ( .A(n9750), .B(n9746), .Z(n9803) );
  XNOR U9977 ( .A(n9745), .B(n9741), .Z(n9804) );
  XNOR U9978 ( .A(n9740), .B(n9736), .Z(n9805) );
  XNOR U9979 ( .A(n9735), .B(n9731), .Z(n9806) );
  XOR U9980 ( .A(n9807), .B(n9730), .Z(n9731) );
  AND U9981 ( .A(a[0]), .B(b[13]), .Z(n9807) );
  XNOR U9982 ( .A(n9808), .B(n9730), .Z(n9732) );
  XNOR U9983 ( .A(n9809), .B(n9810), .Z(n9730) );
  ANDN U9984 ( .B(n9811), .A(n9812), .Z(n9809) );
  AND U9985 ( .A(a[1]), .B(b[12]), .Z(n9808) );
  XNOR U9986 ( .A(n9813), .B(n9735), .Z(n9737) );
  XOR U9987 ( .A(n9814), .B(n9815), .Z(n9735) );
  ANDN U9988 ( .B(n9816), .A(n9817), .Z(n9814) );
  AND U9989 ( .A(a[2]), .B(b[11]), .Z(n9813) );
  XNOR U9990 ( .A(n9818), .B(n9740), .Z(n9742) );
  XOR U9991 ( .A(n9819), .B(n9820), .Z(n9740) );
  ANDN U9992 ( .B(n9821), .A(n9822), .Z(n9819) );
  AND U9993 ( .A(a[3]), .B(b[10]), .Z(n9818) );
  XNOR U9994 ( .A(n9823), .B(n9745), .Z(n9747) );
  XOR U9995 ( .A(n9824), .B(n9825), .Z(n9745) );
  ANDN U9996 ( .B(n9826), .A(n9827), .Z(n9824) );
  AND U9997 ( .A(a[4]), .B(b[9]), .Z(n9823) );
  XNOR U9998 ( .A(n9828), .B(n9750), .Z(n9752) );
  XOR U9999 ( .A(n9829), .B(n9830), .Z(n9750) );
  ANDN U10000 ( .B(n9831), .A(n9832), .Z(n9829) );
  AND U10001 ( .A(a[5]), .B(b[8]), .Z(n9828) );
  XNOR U10002 ( .A(n9833), .B(n9755), .Z(n9757) );
  XOR U10003 ( .A(n9834), .B(n9835), .Z(n9755) );
  ANDN U10004 ( .B(n9836), .A(n9837), .Z(n9834) );
  AND U10005 ( .A(a[6]), .B(b[7]), .Z(n9833) );
  XNOR U10006 ( .A(n9838), .B(n9760), .Z(n9762) );
  XOR U10007 ( .A(n9839), .B(n9840), .Z(n9760) );
  ANDN U10008 ( .B(n9841), .A(n9842), .Z(n9839) );
  AND U10009 ( .A(a[7]), .B(b[6]), .Z(n9838) );
  XNOR U10010 ( .A(n9843), .B(n9765), .Z(n9767) );
  XOR U10011 ( .A(n9844), .B(n9845), .Z(n9765) );
  ANDN U10012 ( .B(n9846), .A(n9847), .Z(n9844) );
  AND U10013 ( .A(b[5]), .B(a[8]), .Z(n9843) );
  XNOR U10014 ( .A(n9848), .B(n9770), .Z(n9772) );
  XOR U10015 ( .A(n9849), .B(n9850), .Z(n9770) );
  ANDN U10016 ( .B(n9851), .A(n9852), .Z(n9849) );
  AND U10017 ( .A(a[9]), .B(b[4]), .Z(n9848) );
  XNOR U10018 ( .A(n9853), .B(n9854), .Z(n9784) );
  OR U10019 ( .A(n9855), .B(n9856), .Z(n9854) );
  XNOR U10020 ( .A(n9857), .B(n9775), .Z(n9777) );
  XNOR U10021 ( .A(n9858), .B(n9859), .Z(n9775) );
  NOR U10022 ( .A(n9860), .B(n9861), .Z(n9858) );
  AND U10023 ( .A(b[3]), .B(a[10]), .Z(n9857) );
  XNOR U10024 ( .A(n9790), .B(n9791), .Z(c[124]) );
  XOR U10025 ( .A(sreg[140]), .B(n9789), .Z(n9791) );
  XOR U10026 ( .A(n9796), .B(n9862), .Z(n9790) );
  XNOR U10027 ( .A(n9795), .B(n9789), .Z(n9862) );
  XOR U10028 ( .A(n9863), .B(n9864), .Z(n9789) );
  ANDN U10029 ( .B(n9865), .A(n9866), .Z(n9863) );
  NANDN U10030 ( .A(n179), .B(a[12]), .Z(n9795) );
  XNOR U10031 ( .A(n9853), .B(n9867), .Z(n9855) );
  NAND U10032 ( .A(a[11]), .B(b[1]), .Z(n9867) );
  XNOR U10033 ( .A(n9853), .B(n9861), .Z(n9868) );
  XOR U10034 ( .A(n9869), .B(n9859), .Z(n9861) );
  AND U10035 ( .A(b[2]), .B(a[10]), .Z(n9869) );
  OR U10036 ( .A(n9870), .B(n9871), .Z(n9853) );
  XOR U10037 ( .A(n9859), .B(n9851), .Z(n9872) );
  XNOR U10038 ( .A(n9850), .B(n9846), .Z(n9873) );
  XNOR U10039 ( .A(n9845), .B(n9841), .Z(n9874) );
  XNOR U10040 ( .A(n9840), .B(n9836), .Z(n9875) );
  XNOR U10041 ( .A(n9835), .B(n9831), .Z(n9876) );
  XNOR U10042 ( .A(n9830), .B(n9826), .Z(n9877) );
  XNOR U10043 ( .A(n9825), .B(n9821), .Z(n9878) );
  XNOR U10044 ( .A(n9820), .B(n9816), .Z(n9879) );
  XNOR U10045 ( .A(n9815), .B(n9811), .Z(n9880) );
  XNOR U10046 ( .A(n9881), .B(n9810), .Z(n9811) );
  AND U10047 ( .A(a[0]), .B(b[12]), .Z(n9881) );
  XOR U10048 ( .A(n9882), .B(n9810), .Z(n9812) );
  XNOR U10049 ( .A(n9883), .B(n9884), .Z(n9810) );
  ANDN U10050 ( .B(n9885), .A(n9886), .Z(n9883) );
  AND U10051 ( .A(a[1]), .B(b[11]), .Z(n9882) );
  XNOR U10052 ( .A(n9887), .B(n9815), .Z(n9817) );
  XOR U10053 ( .A(n9888), .B(n9889), .Z(n9815) );
  ANDN U10054 ( .B(n9890), .A(n9891), .Z(n9888) );
  AND U10055 ( .A(a[2]), .B(b[10]), .Z(n9887) );
  XNOR U10056 ( .A(n9892), .B(n9820), .Z(n9822) );
  XOR U10057 ( .A(n9893), .B(n9894), .Z(n9820) );
  ANDN U10058 ( .B(n9895), .A(n9896), .Z(n9893) );
  AND U10059 ( .A(a[3]), .B(b[9]), .Z(n9892) );
  XNOR U10060 ( .A(n9897), .B(n9825), .Z(n9827) );
  XOR U10061 ( .A(n9898), .B(n9899), .Z(n9825) );
  ANDN U10062 ( .B(n9900), .A(n9901), .Z(n9898) );
  AND U10063 ( .A(a[4]), .B(b[8]), .Z(n9897) );
  XNOR U10064 ( .A(n9902), .B(n9830), .Z(n9832) );
  XOR U10065 ( .A(n9903), .B(n9904), .Z(n9830) );
  ANDN U10066 ( .B(n9905), .A(n9906), .Z(n9903) );
  AND U10067 ( .A(a[5]), .B(b[7]), .Z(n9902) );
  XNOR U10068 ( .A(n9907), .B(n9835), .Z(n9837) );
  XOR U10069 ( .A(n9908), .B(n9909), .Z(n9835) );
  ANDN U10070 ( .B(n9910), .A(n9911), .Z(n9908) );
  AND U10071 ( .A(b[6]), .B(a[6]), .Z(n9907) );
  XNOR U10072 ( .A(n9912), .B(n9840), .Z(n9842) );
  XOR U10073 ( .A(n9913), .B(n9914), .Z(n9840) );
  ANDN U10074 ( .B(n9915), .A(n9916), .Z(n9913) );
  AND U10075 ( .A(a[7]), .B(b[5]), .Z(n9912) );
  XNOR U10076 ( .A(n9917), .B(n9845), .Z(n9847) );
  XOR U10077 ( .A(n9918), .B(n9919), .Z(n9845) );
  ANDN U10078 ( .B(n9920), .A(n9921), .Z(n9918) );
  AND U10079 ( .A(b[4]), .B(a[8]), .Z(n9917) );
  XNOR U10080 ( .A(n9922), .B(n9923), .Z(n9859) );
  OR U10081 ( .A(n9924), .B(n9925), .Z(n9923) );
  XNOR U10082 ( .A(n9926), .B(n9850), .Z(n9852) );
  XNOR U10083 ( .A(n9927), .B(n9928), .Z(n9850) );
  NOR U10084 ( .A(n9929), .B(n9930), .Z(n9927) );
  AND U10085 ( .A(a[9]), .B(b[3]), .Z(n9926) );
  XNOR U10086 ( .A(n9865), .B(n9866), .Z(c[123]) );
  XOR U10087 ( .A(sreg[139]), .B(n9864), .Z(n9866) );
  XOR U10088 ( .A(n9871), .B(n9931), .Z(n9865) );
  XNOR U10089 ( .A(n9870), .B(n9864), .Z(n9931) );
  XOR U10090 ( .A(n9932), .B(n9933), .Z(n9864) );
  ANDN U10091 ( .B(n9934), .A(n9935), .Z(n9932) );
  NANDN U10092 ( .A(n179), .B(a[11]), .Z(n9870) );
  XNOR U10093 ( .A(n9922), .B(n9936), .Z(n9924) );
  NAND U10094 ( .A(b[1]), .B(a[10]), .Z(n9936) );
  XNOR U10095 ( .A(n9922), .B(n9930), .Z(n9937) );
  XOR U10096 ( .A(n9938), .B(n9928), .Z(n9930) );
  AND U10097 ( .A(b[2]), .B(a[9]), .Z(n9938) );
  OR U10098 ( .A(n9939), .B(n9940), .Z(n9922) );
  XOR U10099 ( .A(n9928), .B(n9920), .Z(n9941) );
  XNOR U10100 ( .A(n9919), .B(n9915), .Z(n9942) );
  XNOR U10101 ( .A(n9914), .B(n9910), .Z(n9943) );
  XNOR U10102 ( .A(n9909), .B(n9905), .Z(n9944) );
  XNOR U10103 ( .A(n9904), .B(n9900), .Z(n9945) );
  XNOR U10104 ( .A(n9899), .B(n9895), .Z(n9946) );
  XNOR U10105 ( .A(n9894), .B(n9890), .Z(n9947) );
  XNOR U10106 ( .A(n9889), .B(n9885), .Z(n9948) );
  XOR U10107 ( .A(n9949), .B(n9884), .Z(n9885) );
  AND U10108 ( .A(a[0]), .B(b[11]), .Z(n9949) );
  XNOR U10109 ( .A(n9950), .B(n9884), .Z(n9886) );
  XNOR U10110 ( .A(n9951), .B(n9952), .Z(n9884) );
  ANDN U10111 ( .B(n9953), .A(n9954), .Z(n9951) );
  AND U10112 ( .A(a[1]), .B(b[10]), .Z(n9950) );
  XNOR U10113 ( .A(n9955), .B(n9889), .Z(n9891) );
  XOR U10114 ( .A(n9956), .B(n9957), .Z(n9889) );
  ANDN U10115 ( .B(n9958), .A(n9959), .Z(n9956) );
  AND U10116 ( .A(a[2]), .B(b[9]), .Z(n9955) );
  XNOR U10117 ( .A(n9960), .B(n9894), .Z(n9896) );
  XOR U10118 ( .A(n9961), .B(n9962), .Z(n9894) );
  ANDN U10119 ( .B(n9963), .A(n9964), .Z(n9961) );
  AND U10120 ( .A(a[3]), .B(b[8]), .Z(n9960) );
  XNOR U10121 ( .A(n9965), .B(n9899), .Z(n9901) );
  XOR U10122 ( .A(n9966), .B(n9967), .Z(n9899) );
  ANDN U10123 ( .B(n9968), .A(n9969), .Z(n9966) );
  AND U10124 ( .A(a[4]), .B(b[7]), .Z(n9965) );
  XNOR U10125 ( .A(n9970), .B(n9904), .Z(n9906) );
  XOR U10126 ( .A(n9971), .B(n9972), .Z(n9904) );
  ANDN U10127 ( .B(n9973), .A(n9974), .Z(n9971) );
  AND U10128 ( .A(a[5]), .B(b[6]), .Z(n9970) );
  XNOR U10129 ( .A(n9975), .B(n9909), .Z(n9911) );
  XOR U10130 ( .A(n9976), .B(n9977), .Z(n9909) );
  ANDN U10131 ( .B(n9978), .A(n9979), .Z(n9976) );
  AND U10132 ( .A(b[5]), .B(a[6]), .Z(n9975) );
  XNOR U10133 ( .A(n9980), .B(n9914), .Z(n9916) );
  XOR U10134 ( .A(n9981), .B(n9982), .Z(n9914) );
  ANDN U10135 ( .B(n9983), .A(n9984), .Z(n9981) );
  AND U10136 ( .A(a[7]), .B(b[4]), .Z(n9980) );
  XNOR U10137 ( .A(n9985), .B(n9986), .Z(n9928) );
  OR U10138 ( .A(n9987), .B(n9988), .Z(n9986) );
  XNOR U10139 ( .A(n9989), .B(n9919), .Z(n9921) );
  XNOR U10140 ( .A(n9990), .B(n9991), .Z(n9919) );
  NOR U10141 ( .A(n9992), .B(n9993), .Z(n9990) );
  AND U10142 ( .A(b[3]), .B(a[8]), .Z(n9989) );
  XNOR U10143 ( .A(n9934), .B(n9935), .Z(c[122]) );
  XOR U10144 ( .A(sreg[138]), .B(n9933), .Z(n9935) );
  XOR U10145 ( .A(n9940), .B(n9994), .Z(n9934) );
  XNOR U10146 ( .A(n9939), .B(n9933), .Z(n9994) );
  XOR U10147 ( .A(n9995), .B(n9996), .Z(n9933) );
  ANDN U10148 ( .B(n9997), .A(n9998), .Z(n9995) );
  NANDN U10149 ( .A(n179), .B(a[10]), .Z(n9939) );
  XNOR U10150 ( .A(n9985), .B(n9999), .Z(n9987) );
  NAND U10151 ( .A(a[9]), .B(b[1]), .Z(n9999) );
  XNOR U10152 ( .A(n9985), .B(n9993), .Z(n10000) );
  XOR U10153 ( .A(n10001), .B(n9991), .Z(n9993) );
  AND U10154 ( .A(b[2]), .B(a[8]), .Z(n10001) );
  OR U10155 ( .A(n10002), .B(n10003), .Z(n9985) );
  XOR U10156 ( .A(n9991), .B(n9983), .Z(n10004) );
  XNOR U10157 ( .A(n9982), .B(n9978), .Z(n10005) );
  XNOR U10158 ( .A(n9977), .B(n9973), .Z(n10006) );
  XNOR U10159 ( .A(n9972), .B(n9968), .Z(n10007) );
  XNOR U10160 ( .A(n9967), .B(n9963), .Z(n10008) );
  XNOR U10161 ( .A(n9962), .B(n9958), .Z(n10009) );
  XNOR U10162 ( .A(n9957), .B(n9953), .Z(n10010) );
  XNOR U10163 ( .A(n10011), .B(n9952), .Z(n9953) );
  AND U10164 ( .A(a[0]), .B(b[10]), .Z(n10011) );
  XOR U10165 ( .A(n10012), .B(n9952), .Z(n9954) );
  XNOR U10166 ( .A(n10013), .B(n10014), .Z(n9952) );
  ANDN U10167 ( .B(n10015), .A(n10016), .Z(n10013) );
  AND U10168 ( .A(a[1]), .B(b[9]), .Z(n10012) );
  XNOR U10169 ( .A(n10017), .B(n9957), .Z(n9959) );
  XOR U10170 ( .A(n10018), .B(n10019), .Z(n9957) );
  ANDN U10171 ( .B(n10020), .A(n10021), .Z(n10018) );
  AND U10172 ( .A(a[2]), .B(b[8]), .Z(n10017) );
  XNOR U10173 ( .A(n10022), .B(n9962), .Z(n9964) );
  XOR U10174 ( .A(n10023), .B(n10024), .Z(n9962) );
  ANDN U10175 ( .B(n10025), .A(n10026), .Z(n10023) );
  AND U10176 ( .A(a[3]), .B(b[7]), .Z(n10022) );
  XNOR U10177 ( .A(n10027), .B(n9967), .Z(n9969) );
  XOR U10178 ( .A(n10028), .B(n10029), .Z(n9967) );
  ANDN U10179 ( .B(n10030), .A(n10031), .Z(n10028) );
  AND U10180 ( .A(a[4]), .B(b[6]), .Z(n10027) );
  XNOR U10181 ( .A(n10032), .B(n9972), .Z(n9974) );
  XOR U10182 ( .A(n10033), .B(n10034), .Z(n9972) );
  ANDN U10183 ( .B(n10035), .A(n10036), .Z(n10033) );
  AND U10184 ( .A(a[5]), .B(b[5]), .Z(n10032) );
  XNOR U10185 ( .A(n10037), .B(n9977), .Z(n9979) );
  XOR U10186 ( .A(n10038), .B(n10039), .Z(n9977) );
  ANDN U10187 ( .B(n10040), .A(n10041), .Z(n10038) );
  AND U10188 ( .A(b[4]), .B(a[6]), .Z(n10037) );
  XNOR U10189 ( .A(n10042), .B(n10043), .Z(n9991) );
  OR U10190 ( .A(n10044), .B(n10045), .Z(n10043) );
  XNOR U10191 ( .A(n10046), .B(n9982), .Z(n9984) );
  XNOR U10192 ( .A(n10047), .B(n10048), .Z(n9982) );
  NOR U10193 ( .A(n10049), .B(n10050), .Z(n10047) );
  AND U10194 ( .A(a[7]), .B(b[3]), .Z(n10046) );
  XNOR U10195 ( .A(n9997), .B(n9998), .Z(c[121]) );
  XOR U10196 ( .A(sreg[137]), .B(n9996), .Z(n9998) );
  XOR U10197 ( .A(n10003), .B(n10051), .Z(n9997) );
  XNOR U10198 ( .A(n10002), .B(n9996), .Z(n10051) );
  XOR U10199 ( .A(n10052), .B(n10053), .Z(n9996) );
  ANDN U10200 ( .B(n10054), .A(n10055), .Z(n10052) );
  NANDN U10201 ( .A(n179), .B(a[9]), .Z(n10002) );
  XNOR U10202 ( .A(n10042), .B(n10056), .Z(n10044) );
  NAND U10203 ( .A(b[1]), .B(a[8]), .Z(n10056) );
  XNOR U10204 ( .A(n10042), .B(n10050), .Z(n10057) );
  XOR U10205 ( .A(n10058), .B(n10048), .Z(n10050) );
  AND U10206 ( .A(b[2]), .B(a[7]), .Z(n10058) );
  OR U10207 ( .A(n10059), .B(n10060), .Z(n10042) );
  XOR U10208 ( .A(n10048), .B(n10040), .Z(n10061) );
  XNOR U10209 ( .A(n10039), .B(n10035), .Z(n10062) );
  XNOR U10210 ( .A(n10034), .B(n10030), .Z(n10063) );
  XNOR U10211 ( .A(n10029), .B(n10025), .Z(n10064) );
  XNOR U10212 ( .A(n10024), .B(n10020), .Z(n10065) );
  XNOR U10213 ( .A(n10019), .B(n10015), .Z(n10066) );
  XOR U10214 ( .A(n10067), .B(n10014), .Z(n10015) );
  AND U10215 ( .A(a[0]), .B(b[9]), .Z(n10067) );
  XNOR U10216 ( .A(n10068), .B(n10014), .Z(n10016) );
  XNOR U10217 ( .A(n10069), .B(n10070), .Z(n10014) );
  ANDN U10218 ( .B(n10071), .A(n10072), .Z(n10069) );
  AND U10219 ( .A(a[1]), .B(b[8]), .Z(n10068) );
  XNOR U10220 ( .A(n10073), .B(n10019), .Z(n10021) );
  XOR U10221 ( .A(n10074), .B(n10075), .Z(n10019) );
  ANDN U10222 ( .B(n10076), .A(n10077), .Z(n10074) );
  AND U10223 ( .A(a[2]), .B(b[7]), .Z(n10073) );
  XNOR U10224 ( .A(n10078), .B(n10024), .Z(n10026) );
  XOR U10225 ( .A(n10079), .B(n10080), .Z(n10024) );
  ANDN U10226 ( .B(n10081), .A(n10082), .Z(n10079) );
  AND U10227 ( .A(a[3]), .B(b[6]), .Z(n10078) );
  XNOR U10228 ( .A(n10083), .B(n10029), .Z(n10031) );
  XOR U10229 ( .A(n10084), .B(n10085), .Z(n10029) );
  ANDN U10230 ( .B(n10086), .A(n10087), .Z(n10084) );
  AND U10231 ( .A(a[4]), .B(b[5]), .Z(n10083) );
  XNOR U10232 ( .A(n10088), .B(n10034), .Z(n10036) );
  XOR U10233 ( .A(n10089), .B(n10090), .Z(n10034) );
  ANDN U10234 ( .B(n10091), .A(n10092), .Z(n10089) );
  AND U10235 ( .A(a[5]), .B(b[4]), .Z(n10088) );
  XNOR U10236 ( .A(n10093), .B(n10094), .Z(n10048) );
  OR U10237 ( .A(n10095), .B(n10096), .Z(n10094) );
  XNOR U10238 ( .A(n10097), .B(n10039), .Z(n10041) );
  XNOR U10239 ( .A(n10098), .B(n10099), .Z(n10039) );
  NOR U10240 ( .A(n10100), .B(n10101), .Z(n10098) );
  AND U10241 ( .A(b[3]), .B(a[6]), .Z(n10097) );
  XNOR U10242 ( .A(n10054), .B(n10055), .Z(c[120]) );
  XOR U10243 ( .A(sreg[136]), .B(n10053), .Z(n10055) );
  XOR U10244 ( .A(n10060), .B(n10102), .Z(n10054) );
  XNOR U10245 ( .A(n10059), .B(n10053), .Z(n10102) );
  XOR U10246 ( .A(n10103), .B(n10104), .Z(n10053) );
  ANDN U10247 ( .B(n10105), .A(n10106), .Z(n10103) );
  NANDN U10248 ( .A(n179), .B(a[8]), .Z(n10059) );
  XNOR U10249 ( .A(n10093), .B(n10107), .Z(n10095) );
  NAND U10250 ( .A(a[7]), .B(b[1]), .Z(n10107) );
  XNOR U10251 ( .A(n10093), .B(n10101), .Z(n10108) );
  XOR U10252 ( .A(n10109), .B(n10099), .Z(n10101) );
  AND U10253 ( .A(b[2]), .B(a[6]), .Z(n10109) );
  OR U10254 ( .A(n10110), .B(n10111), .Z(n10093) );
  XOR U10255 ( .A(n10099), .B(n10091), .Z(n10112) );
  XNOR U10256 ( .A(n10090), .B(n10086), .Z(n10113) );
  XNOR U10257 ( .A(n10085), .B(n10081), .Z(n10114) );
  XNOR U10258 ( .A(n10080), .B(n10076), .Z(n10115) );
  XNOR U10259 ( .A(n10075), .B(n10071), .Z(n10116) );
  XNOR U10260 ( .A(n10117), .B(n10070), .Z(n10071) );
  AND U10261 ( .A(a[0]), .B(b[8]), .Z(n10117) );
  XOR U10262 ( .A(n10118), .B(n10070), .Z(n10072) );
  XNOR U10263 ( .A(n10119), .B(n10120), .Z(n10070) );
  ANDN U10264 ( .B(n10121), .A(n10122), .Z(n10119) );
  AND U10265 ( .A(a[1]), .B(b[7]), .Z(n10118) );
  XNOR U10266 ( .A(n10123), .B(n10075), .Z(n10077) );
  XOR U10267 ( .A(n10124), .B(n10125), .Z(n10075) );
  ANDN U10268 ( .B(n10126), .A(n10127), .Z(n10124) );
  AND U10269 ( .A(a[2]), .B(b[6]), .Z(n10123) );
  XNOR U10270 ( .A(n10128), .B(n10080), .Z(n10082) );
  XOR U10271 ( .A(n10129), .B(n10130), .Z(n10080) );
  ANDN U10272 ( .B(n10131), .A(n10132), .Z(n10129) );
  AND U10273 ( .A(a[3]), .B(b[5]), .Z(n10128) );
  XNOR U10274 ( .A(n10133), .B(n10085), .Z(n10087) );
  XOR U10275 ( .A(n10134), .B(n10135), .Z(n10085) );
  ANDN U10276 ( .B(n10136), .A(n10137), .Z(n10134) );
  AND U10277 ( .A(b[4]), .B(a[4]), .Z(n10133) );
  XNOR U10278 ( .A(n10138), .B(n10139), .Z(n10099) );
  OR U10279 ( .A(n10140), .B(n10141), .Z(n10139) );
  XNOR U10280 ( .A(n10142), .B(n10090), .Z(n10092) );
  XNOR U10281 ( .A(n10143), .B(n10144), .Z(n10090) );
  NOR U10282 ( .A(n10145), .B(n10146), .Z(n10143) );
  AND U10283 ( .A(a[5]), .B(b[3]), .Z(n10142) );
  XNOR U10284 ( .A(n10105), .B(n10106), .Z(c[119]) );
  XOR U10285 ( .A(sreg[135]), .B(n10104), .Z(n10106) );
  XOR U10286 ( .A(n10111), .B(n10147), .Z(n10105) );
  XNOR U10287 ( .A(n10110), .B(n10104), .Z(n10147) );
  XOR U10288 ( .A(n10148), .B(n10149), .Z(n10104) );
  ANDN U10289 ( .B(n10150), .A(n10151), .Z(n10148) );
  NANDN U10290 ( .A(n179), .B(a[7]), .Z(n10110) );
  XNOR U10291 ( .A(n10138), .B(n10152), .Z(n10140) );
  NAND U10292 ( .A(b[1]), .B(a[6]), .Z(n10152) );
  XNOR U10293 ( .A(n10138), .B(n10146), .Z(n10153) );
  XOR U10294 ( .A(n10154), .B(n10144), .Z(n10146) );
  AND U10295 ( .A(b[2]), .B(a[5]), .Z(n10154) );
  OR U10296 ( .A(n10155), .B(n10156), .Z(n10138) );
  XOR U10297 ( .A(n10144), .B(n10136), .Z(n10157) );
  XNOR U10298 ( .A(n10135), .B(n10131), .Z(n10158) );
  XNOR U10299 ( .A(n10130), .B(n10126), .Z(n10159) );
  XNOR U10300 ( .A(n10125), .B(n10121), .Z(n10160) );
  XOR U10301 ( .A(n10161), .B(n10120), .Z(n10121) );
  AND U10302 ( .A(a[0]), .B(b[7]), .Z(n10161) );
  XNOR U10303 ( .A(n10162), .B(n10120), .Z(n10122) );
  XNOR U10304 ( .A(n10163), .B(n10164), .Z(n10120) );
  ANDN U10305 ( .B(n10165), .A(n10166), .Z(n10163) );
  AND U10306 ( .A(a[1]), .B(b[6]), .Z(n10162) );
  XNOR U10307 ( .A(n10167), .B(n10125), .Z(n10127) );
  XOR U10308 ( .A(n10168), .B(n10169), .Z(n10125) );
  ANDN U10309 ( .B(n10170), .A(n10171), .Z(n10168) );
  AND U10310 ( .A(a[2]), .B(b[5]), .Z(n10167) );
  XNOR U10311 ( .A(n10172), .B(n10130), .Z(n10132) );
  XOR U10312 ( .A(n10173), .B(n10174), .Z(n10130) );
  ANDN U10313 ( .B(n10175), .A(n10176), .Z(n10173) );
  AND U10314 ( .A(a[3]), .B(b[4]), .Z(n10172) );
  XNOR U10315 ( .A(n10177), .B(n10178), .Z(n10144) );
  OR U10316 ( .A(n10179), .B(n10180), .Z(n10178) );
  XNOR U10317 ( .A(n10181), .B(n10135), .Z(n10137) );
  XNOR U10318 ( .A(n10182), .B(n10183), .Z(n10135) );
  NOR U10319 ( .A(n10184), .B(n10185), .Z(n10182) );
  AND U10320 ( .A(b[3]), .B(a[4]), .Z(n10181) );
  XNOR U10321 ( .A(n10150), .B(n10151), .Z(c[118]) );
  XOR U10322 ( .A(sreg[134]), .B(n10149), .Z(n10151) );
  XOR U10323 ( .A(n10156), .B(n10186), .Z(n10150) );
  XNOR U10324 ( .A(n10155), .B(n10149), .Z(n10186) );
  XOR U10325 ( .A(n10187), .B(n10188), .Z(n10149) );
  ANDN U10326 ( .B(n10189), .A(n10190), .Z(n10187) );
  NANDN U10327 ( .A(n179), .B(a[6]), .Z(n10155) );
  XNOR U10328 ( .A(n10177), .B(n10191), .Z(n10179) );
  NAND U10329 ( .A(a[5]), .B(b[1]), .Z(n10191) );
  XNOR U10330 ( .A(n10177), .B(n10185), .Z(n10192) );
  XOR U10331 ( .A(n10193), .B(n10183), .Z(n10185) );
  AND U10332 ( .A(b[2]), .B(a[4]), .Z(n10193) );
  OR U10333 ( .A(n10194), .B(n10195), .Z(n10177) );
  XOR U10334 ( .A(n10183), .B(n10175), .Z(n10196) );
  XNOR U10335 ( .A(n10174), .B(n10170), .Z(n10197) );
  XNOR U10336 ( .A(n10169), .B(n10165), .Z(n10198) );
  XNOR U10337 ( .A(n10199), .B(n10164), .Z(n10165) );
  AND U10338 ( .A(a[0]), .B(b[6]), .Z(n10199) );
  XOR U10339 ( .A(n10200), .B(n10164), .Z(n10166) );
  XNOR U10340 ( .A(n10201), .B(n10202), .Z(n10164) );
  ANDN U10341 ( .B(n10203), .A(n10204), .Z(n10201) );
  AND U10342 ( .A(a[1]), .B(b[5]), .Z(n10200) );
  XNOR U10343 ( .A(n10205), .B(n10169), .Z(n10171) );
  XOR U10344 ( .A(n10206), .B(n10207), .Z(n10169) );
  ANDN U10345 ( .B(n10208), .A(n10209), .Z(n10206) );
  AND U10346 ( .A(a[2]), .B(b[4]), .Z(n10205) );
  XNOR U10347 ( .A(n10210), .B(n10211), .Z(n10183) );
  OR U10348 ( .A(n10212), .B(n10213), .Z(n10211) );
  XNOR U10349 ( .A(n10214), .B(n10174), .Z(n10176) );
  XNOR U10350 ( .A(n10215), .B(n10216), .Z(n10174) );
  NOR U10351 ( .A(n10217), .B(n10218), .Z(n10215) );
  AND U10352 ( .A(a[3]), .B(b[3]), .Z(n10214) );
  XNOR U10353 ( .A(n10189), .B(n10190), .Z(c[117]) );
  XOR U10354 ( .A(sreg[133]), .B(n10188), .Z(n10190) );
  XOR U10355 ( .A(n10195), .B(n10219), .Z(n10189) );
  XNOR U10356 ( .A(n10194), .B(n10188), .Z(n10219) );
  XOR U10357 ( .A(n10220), .B(n10221), .Z(n10188) );
  ANDN U10358 ( .B(n10222), .A(n10223), .Z(n10220) );
  NANDN U10359 ( .A(n179), .B(a[5]), .Z(n10194) );
  XNOR U10360 ( .A(n10210), .B(n10224), .Z(n10212) );
  NAND U10361 ( .A(b[1]), .B(a[4]), .Z(n10224) );
  XNOR U10362 ( .A(n10210), .B(n10218), .Z(n10225) );
  XOR U10363 ( .A(n10226), .B(n10216), .Z(n10218) );
  AND U10364 ( .A(b[2]), .B(a[3]), .Z(n10226) );
  OR U10365 ( .A(n10227), .B(n10228), .Z(n10210) );
  XOR U10366 ( .A(n10216), .B(n10208), .Z(n10229) );
  XNOR U10367 ( .A(n10207), .B(n10203), .Z(n10230) );
  XOR U10368 ( .A(n10231), .B(n10202), .Z(n10203) );
  AND U10369 ( .A(a[0]), .B(b[5]), .Z(n10231) );
  XNOR U10370 ( .A(n10232), .B(n10202), .Z(n10204) );
  XNOR U10371 ( .A(n10233), .B(n10234), .Z(n10202) );
  ANDN U10372 ( .B(n10235), .A(n10236), .Z(n10233) );
  AND U10373 ( .A(a[1]), .B(b[4]), .Z(n10232) );
  XNOR U10374 ( .A(n10237), .B(n10238), .Z(n10216) );
  OR U10375 ( .A(n10239), .B(n10240), .Z(n10238) );
  XNOR U10376 ( .A(n10241), .B(n10207), .Z(n10209) );
  XNOR U10377 ( .A(n10242), .B(n10243), .Z(n10207) );
  NOR U10378 ( .A(n10244), .B(n10245), .Z(n10242) );
  AND U10379 ( .A(a[2]), .B(b[3]), .Z(n10241) );
  XNOR U10380 ( .A(n10222), .B(n10223), .Z(c[116]) );
  XOR U10381 ( .A(sreg[132]), .B(n10221), .Z(n10223) );
  XOR U10382 ( .A(n10228), .B(n10246), .Z(n10222) );
  XNOR U10383 ( .A(n10227), .B(n10221), .Z(n10246) );
  XOR U10384 ( .A(n10247), .B(n10248), .Z(n10221) );
  ANDN U10385 ( .B(n10249), .A(n10250), .Z(n10247) );
  NANDN U10386 ( .A(n179), .B(a[4]), .Z(n10227) );
  XNOR U10387 ( .A(n10237), .B(n10251), .Z(n10239) );
  NAND U10388 ( .A(a[3]), .B(b[1]), .Z(n10251) );
  XNOR U10389 ( .A(n10237), .B(n10245), .Z(n10252) );
  XOR U10390 ( .A(n10253), .B(n10243), .Z(n10245) );
  AND U10391 ( .A(b[2]), .B(a[2]), .Z(n10253) );
  OR U10392 ( .A(n10254), .B(n10255), .Z(n10237) );
  XOR U10393 ( .A(n10243), .B(n10235), .Z(n10256) );
  XNOR U10394 ( .A(n10257), .B(n10234), .Z(n10235) );
  AND U10395 ( .A(a[0]), .B(b[4]), .Z(n10257) );
  XOR U10396 ( .A(n10258), .B(n10259), .Z(n10243) );
  OR U10397 ( .A(n10260), .B(n10261), .Z(n10259) );
  XOR U10398 ( .A(n10262), .B(n10234), .Z(n10236) );
  XOR U10399 ( .A(n10263), .B(n10264), .Z(n10234) );
  NOR U10400 ( .A(n10265), .B(n10266), .Z(n10263) );
  AND U10401 ( .A(a[1]), .B(b[3]), .Z(n10262) );
  XNOR U10402 ( .A(n10249), .B(n10250), .Z(c[115]) );
  XOR U10403 ( .A(sreg[131]), .B(n10248), .Z(n10250) );
  XOR U10404 ( .A(n10255), .B(n10267), .Z(n10249) );
  XNOR U10405 ( .A(n10254), .B(n10248), .Z(n10267) );
  XNOR U10406 ( .A(n10268), .B(n10269), .Z(n10248) );
  ANDN U10407 ( .B(n10270), .A(n10271), .Z(n10268) );
  NANDN U10408 ( .A(n179), .B(a[3]), .Z(n10254) );
  XOR U10409 ( .A(n10258), .B(n10272), .Z(n10260) );
  NAND U10410 ( .A(b[1]), .B(a[2]), .Z(n10272) );
  XOR U10411 ( .A(n10258), .B(n10266), .Z(n10273) );
  XNOR U10412 ( .A(n10274), .B(n10275), .Z(n10266) );
  AND U10413 ( .A(b[2]), .B(a[1]), .Z(n10274) );
  NOR U10414 ( .A(n10276), .B(n10277), .Z(n10258) );
  XOR U10415 ( .A(n10278), .B(n10264), .Z(n10265) );
  IV U10416 ( .A(n10275), .Z(n10264) );
  XOR U10417 ( .A(n10279), .B(n10280), .Z(n10275) );
  OR U10418 ( .A(n10281), .B(n10282), .Z(n10280) );
  AND U10419 ( .A(a[0]), .B(b[3]), .Z(n10278) );
  XNOR U10420 ( .A(n10270), .B(n10271), .Z(c[114]) );
  XNOR U10421 ( .A(sreg[130]), .B(n10269), .Z(n10271) );
  XNOR U10422 ( .A(n10277), .B(n10284), .Z(n10283) );
  IV U10423 ( .A(n10269), .Z(n10284) );
  XNOR U10424 ( .A(n10285), .B(n10286), .Z(n10269) );
  NAND U10425 ( .A(n10287), .B(n10288), .Z(n10286) );
  NANDN U10426 ( .A(n179), .B(a[2]), .Z(n10277) );
  NAND U10427 ( .A(a[1]), .B(b[1]), .Z(n10289) );
  XOR U10428 ( .A(n10290), .B(n10279), .Z(n10281) );
  NANDN U10429 ( .A(n10291), .B(n10292), .Z(n10279) );
  AND U10430 ( .A(b[2]), .B(a[0]), .Z(n10290) );
  XOR U10431 ( .A(n10287), .B(n10288), .Z(c[113]) );
  XOR U10432 ( .A(sreg[129]), .B(n10285), .Z(n10288) );
  XNOR U10433 ( .A(n10285), .B(n10293), .Z(n10287) );
  XOR U10434 ( .A(n10291), .B(n10292), .Z(n10293) );
  AND U10435 ( .A(a[1]), .B(b[0]), .Z(n10292) );
  NAND U10436 ( .A(b[1]), .B(a[0]), .Z(n10291) );
  ANDN U10437 ( .B(sreg[128]), .A(n10294), .Z(n10285) );
  XNOR U10438 ( .A(sreg[128]), .B(n10294), .Z(c[112]) );
  NANDN U10439 ( .A(n179), .B(a[0]), .Z(n10294) );
  IV U10440 ( .A(b[0]), .Z(n179) );
endmodule

