
module sum_N256_CC4 ( clk, rst, a, b, c );
  input [63:0] a;
  input [63:0] b;
  output [63:0] c;
  input clk, rst;
  wire   carry_on, carry_on_d, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255;

  DFF carry_on_reg ( .D(carry_on_d), .CLK(clk), .RST(rst), .Q(carry_on) );
  XOR U3 ( .A(a[3]), .B(n245), .Z(n107) );
  XOR U4 ( .A(a[6]), .B(n236), .Z(n8) );
  XOR U5 ( .A(a[9]), .B(n227), .Z(n5) );
  XOR U6 ( .A(a[12]), .B(n215), .Z(n217) );
  XOR U7 ( .A(a[15]), .B(n203), .Z(n205) );
  XOR U8 ( .A(a[18]), .B(n191), .Z(n193) );
  XOR U9 ( .A(a[21]), .B(n178), .Z(n180) );
  XOR U10 ( .A(a[24]), .B(n166), .Z(n168) );
  XOR U11 ( .A(a[27]), .B(n154), .Z(n156) );
  XOR U12 ( .A(a[30]), .B(n141), .Z(n143) );
  XOR U13 ( .A(a[33]), .B(n129), .Z(n131) );
  XOR U14 ( .A(a[36]), .B(n117), .Z(n119) );
  XOR U15 ( .A(a[39]), .B(n104), .Z(n106) );
  XOR U16 ( .A(a[42]), .B(n92), .Z(n94) );
  XOR U17 ( .A(a[45]), .B(n80), .Z(n82) );
  XOR U18 ( .A(a[48]), .B(n68), .Z(n70) );
  XOR U19 ( .A(a[51]), .B(n55), .Z(n57) );
  XOR U20 ( .A(a[54]), .B(n43), .Z(n45) );
  XOR U21 ( .A(a[57]), .B(n31), .Z(n33) );
  XOR U22 ( .A(a[60]), .B(n18), .Z(n20) );
  XOR U23 ( .A(a[1]), .B(n251), .Z(n189) );
  XOR U24 ( .A(a[4]), .B(n242), .Z(n66) );
  XOR U25 ( .A(a[7]), .B(n233), .Z(n7) );
  XOR U26 ( .A(a[10]), .B(n223), .Z(n225) );
  XOR U27 ( .A(a[13]), .B(n211), .Z(n213) );
  XOR U28 ( .A(a[16]), .B(n199), .Z(n201) );
  XOR U29 ( .A(a[19]), .B(n186), .Z(n188) );
  XOR U30 ( .A(a[22]), .B(n174), .Z(n176) );
  XOR U31 ( .A(a[25]), .B(n162), .Z(n164) );
  XOR U32 ( .A(a[28]), .B(n150), .Z(n152) );
  XOR U33 ( .A(a[31]), .B(n137), .Z(n139) );
  XOR U34 ( .A(a[34]), .B(n125), .Z(n127) );
  XOR U35 ( .A(a[37]), .B(n113), .Z(n115) );
  XOR U36 ( .A(a[40]), .B(n100), .Z(n102) );
  XOR U37 ( .A(a[43]), .B(n88), .Z(n90) );
  XOR U38 ( .A(a[46]), .B(n76), .Z(n78) );
  XOR U39 ( .A(a[49]), .B(n63), .Z(n65) );
  XOR U40 ( .A(a[52]), .B(n51), .Z(n53) );
  XOR U41 ( .A(a[55]), .B(n39), .Z(n41) );
  XOR U42 ( .A(a[58]), .B(n27), .Z(n29) );
  XOR U43 ( .A(a[61]), .B(n14), .Z(n16) );
  XOR U44 ( .A(a[2]), .B(n248), .Z(n148) );
  XOR U45 ( .A(a[5]), .B(n239), .Z(n25) );
  XOR U46 ( .A(a[8]), .B(n230), .Z(n6) );
  XOR U47 ( .A(a[11]), .B(n219), .Z(n221) );
  XOR U48 ( .A(a[14]), .B(n207), .Z(n209) );
  XOR U49 ( .A(a[17]), .B(n195), .Z(n197) );
  XOR U50 ( .A(a[20]), .B(n182), .Z(n184) );
  XOR U51 ( .A(a[23]), .B(n170), .Z(n172) );
  XOR U52 ( .A(a[26]), .B(n158), .Z(n160) );
  XOR U53 ( .A(a[29]), .B(n145), .Z(n147) );
  XOR U54 ( .A(a[32]), .B(n133), .Z(n135) );
  XOR U55 ( .A(a[35]), .B(n121), .Z(n123) );
  XOR U56 ( .A(a[38]), .B(n109), .Z(n111) );
  XOR U57 ( .A(a[41]), .B(n96), .Z(n98) );
  XOR U58 ( .A(a[44]), .B(n84), .Z(n86) );
  XOR U59 ( .A(a[47]), .B(n72), .Z(n74) );
  XOR U60 ( .A(a[50]), .B(n59), .Z(n61) );
  XOR U61 ( .A(a[53]), .B(n47), .Z(n49) );
  XOR U62 ( .A(a[56]), .B(n35), .Z(n37) );
  XOR U63 ( .A(a[59]), .B(n22), .Z(n24) );
  XOR U64 ( .A(a[62]), .B(n10), .Z(n12) );
  XOR U65 ( .A(n1), .B(n2), .Z(carry_on_d) );
  ANDN U66 ( .B(n3), .A(n4), .Z(n1) );
  XOR U67 ( .A(b[63]), .B(n2), .Z(n3) );
  XNOR U68 ( .A(b[9]), .B(n5), .Z(c[9]) );
  XNOR U69 ( .A(b[8]), .B(n6), .Z(c[8]) );
  XNOR U70 ( .A(b[7]), .B(n7), .Z(c[7]) );
  XNOR U71 ( .A(b[6]), .B(n8), .Z(c[6]) );
  XNOR U72 ( .A(b[63]), .B(n4), .Z(c[63]) );
  XNOR U73 ( .A(a[63]), .B(n2), .Z(n4) );
  XNOR U74 ( .A(n9), .B(n10), .Z(n2) );
  ANDN U75 ( .B(n11), .A(n12), .Z(n9) );
  XNOR U76 ( .A(b[62]), .B(n10), .Z(n11) );
  XNOR U77 ( .A(b[62]), .B(n12), .Z(c[62]) );
  XOR U78 ( .A(n13), .B(n14), .Z(n10) );
  ANDN U79 ( .B(n15), .A(n16), .Z(n13) );
  XNOR U80 ( .A(b[61]), .B(n14), .Z(n15) );
  XNOR U81 ( .A(b[61]), .B(n16), .Z(c[61]) );
  XOR U82 ( .A(n17), .B(n18), .Z(n14) );
  ANDN U83 ( .B(n19), .A(n20), .Z(n17) );
  XNOR U84 ( .A(b[60]), .B(n18), .Z(n19) );
  XNOR U85 ( .A(b[60]), .B(n20), .Z(c[60]) );
  XOR U86 ( .A(n21), .B(n22), .Z(n18) );
  ANDN U87 ( .B(n23), .A(n24), .Z(n21) );
  XNOR U88 ( .A(b[59]), .B(n22), .Z(n23) );
  XNOR U89 ( .A(b[5]), .B(n25), .Z(c[5]) );
  XNOR U90 ( .A(b[59]), .B(n24), .Z(c[59]) );
  XOR U91 ( .A(n26), .B(n27), .Z(n22) );
  ANDN U92 ( .B(n28), .A(n29), .Z(n26) );
  XNOR U93 ( .A(b[58]), .B(n27), .Z(n28) );
  XNOR U94 ( .A(b[58]), .B(n29), .Z(c[58]) );
  XOR U95 ( .A(n30), .B(n31), .Z(n27) );
  ANDN U96 ( .B(n32), .A(n33), .Z(n30) );
  XNOR U97 ( .A(b[57]), .B(n31), .Z(n32) );
  XNOR U98 ( .A(b[57]), .B(n33), .Z(c[57]) );
  XOR U99 ( .A(n34), .B(n35), .Z(n31) );
  ANDN U100 ( .B(n36), .A(n37), .Z(n34) );
  XNOR U101 ( .A(b[56]), .B(n35), .Z(n36) );
  XNOR U102 ( .A(b[56]), .B(n37), .Z(c[56]) );
  XOR U103 ( .A(n38), .B(n39), .Z(n35) );
  ANDN U104 ( .B(n40), .A(n41), .Z(n38) );
  XNOR U105 ( .A(b[55]), .B(n39), .Z(n40) );
  XNOR U106 ( .A(b[55]), .B(n41), .Z(c[55]) );
  XOR U107 ( .A(n42), .B(n43), .Z(n39) );
  ANDN U108 ( .B(n44), .A(n45), .Z(n42) );
  XNOR U109 ( .A(b[54]), .B(n43), .Z(n44) );
  XNOR U110 ( .A(b[54]), .B(n45), .Z(c[54]) );
  XOR U111 ( .A(n46), .B(n47), .Z(n43) );
  ANDN U112 ( .B(n48), .A(n49), .Z(n46) );
  XNOR U113 ( .A(b[53]), .B(n47), .Z(n48) );
  XNOR U114 ( .A(b[53]), .B(n49), .Z(c[53]) );
  XOR U115 ( .A(n50), .B(n51), .Z(n47) );
  ANDN U116 ( .B(n52), .A(n53), .Z(n50) );
  XNOR U117 ( .A(b[52]), .B(n51), .Z(n52) );
  XNOR U118 ( .A(b[52]), .B(n53), .Z(c[52]) );
  XOR U119 ( .A(n54), .B(n55), .Z(n51) );
  ANDN U120 ( .B(n56), .A(n57), .Z(n54) );
  XNOR U121 ( .A(b[51]), .B(n55), .Z(n56) );
  XNOR U122 ( .A(b[51]), .B(n57), .Z(c[51]) );
  XOR U123 ( .A(n58), .B(n59), .Z(n55) );
  ANDN U124 ( .B(n60), .A(n61), .Z(n58) );
  XNOR U125 ( .A(b[50]), .B(n59), .Z(n60) );
  XNOR U126 ( .A(b[50]), .B(n61), .Z(c[50]) );
  XOR U127 ( .A(n62), .B(n63), .Z(n59) );
  ANDN U128 ( .B(n64), .A(n65), .Z(n62) );
  XNOR U129 ( .A(b[49]), .B(n63), .Z(n64) );
  XNOR U130 ( .A(b[4]), .B(n66), .Z(c[4]) );
  XNOR U131 ( .A(b[49]), .B(n65), .Z(c[49]) );
  XOR U132 ( .A(n67), .B(n68), .Z(n63) );
  ANDN U133 ( .B(n69), .A(n70), .Z(n67) );
  XNOR U134 ( .A(b[48]), .B(n68), .Z(n69) );
  XNOR U135 ( .A(b[48]), .B(n70), .Z(c[48]) );
  XOR U136 ( .A(n71), .B(n72), .Z(n68) );
  ANDN U137 ( .B(n73), .A(n74), .Z(n71) );
  XNOR U138 ( .A(b[47]), .B(n72), .Z(n73) );
  XNOR U139 ( .A(b[47]), .B(n74), .Z(c[47]) );
  XOR U140 ( .A(n75), .B(n76), .Z(n72) );
  ANDN U141 ( .B(n77), .A(n78), .Z(n75) );
  XNOR U142 ( .A(b[46]), .B(n76), .Z(n77) );
  XNOR U143 ( .A(b[46]), .B(n78), .Z(c[46]) );
  XOR U144 ( .A(n79), .B(n80), .Z(n76) );
  ANDN U145 ( .B(n81), .A(n82), .Z(n79) );
  XNOR U146 ( .A(b[45]), .B(n80), .Z(n81) );
  XNOR U147 ( .A(b[45]), .B(n82), .Z(c[45]) );
  XOR U148 ( .A(n83), .B(n84), .Z(n80) );
  ANDN U149 ( .B(n85), .A(n86), .Z(n83) );
  XNOR U150 ( .A(b[44]), .B(n84), .Z(n85) );
  XNOR U151 ( .A(b[44]), .B(n86), .Z(c[44]) );
  XOR U152 ( .A(n87), .B(n88), .Z(n84) );
  ANDN U153 ( .B(n89), .A(n90), .Z(n87) );
  XNOR U154 ( .A(b[43]), .B(n88), .Z(n89) );
  XNOR U155 ( .A(b[43]), .B(n90), .Z(c[43]) );
  XOR U156 ( .A(n91), .B(n92), .Z(n88) );
  ANDN U157 ( .B(n93), .A(n94), .Z(n91) );
  XNOR U158 ( .A(b[42]), .B(n92), .Z(n93) );
  XNOR U159 ( .A(b[42]), .B(n94), .Z(c[42]) );
  XOR U160 ( .A(n95), .B(n96), .Z(n92) );
  ANDN U161 ( .B(n97), .A(n98), .Z(n95) );
  XNOR U162 ( .A(b[41]), .B(n96), .Z(n97) );
  XNOR U163 ( .A(b[41]), .B(n98), .Z(c[41]) );
  XOR U164 ( .A(n99), .B(n100), .Z(n96) );
  ANDN U165 ( .B(n101), .A(n102), .Z(n99) );
  XNOR U166 ( .A(b[40]), .B(n100), .Z(n101) );
  XNOR U167 ( .A(b[40]), .B(n102), .Z(c[40]) );
  XOR U168 ( .A(n103), .B(n104), .Z(n100) );
  ANDN U169 ( .B(n105), .A(n106), .Z(n103) );
  XNOR U170 ( .A(b[39]), .B(n104), .Z(n105) );
  XNOR U171 ( .A(b[3]), .B(n107), .Z(c[3]) );
  XNOR U172 ( .A(b[39]), .B(n106), .Z(c[39]) );
  XOR U173 ( .A(n108), .B(n109), .Z(n104) );
  ANDN U174 ( .B(n110), .A(n111), .Z(n108) );
  XNOR U175 ( .A(b[38]), .B(n109), .Z(n110) );
  XNOR U176 ( .A(b[38]), .B(n111), .Z(c[38]) );
  XOR U177 ( .A(n112), .B(n113), .Z(n109) );
  ANDN U178 ( .B(n114), .A(n115), .Z(n112) );
  XNOR U179 ( .A(b[37]), .B(n113), .Z(n114) );
  XNOR U180 ( .A(b[37]), .B(n115), .Z(c[37]) );
  XOR U181 ( .A(n116), .B(n117), .Z(n113) );
  ANDN U182 ( .B(n118), .A(n119), .Z(n116) );
  XNOR U183 ( .A(b[36]), .B(n117), .Z(n118) );
  XNOR U184 ( .A(b[36]), .B(n119), .Z(c[36]) );
  XOR U185 ( .A(n120), .B(n121), .Z(n117) );
  ANDN U186 ( .B(n122), .A(n123), .Z(n120) );
  XNOR U187 ( .A(b[35]), .B(n121), .Z(n122) );
  XNOR U188 ( .A(b[35]), .B(n123), .Z(c[35]) );
  XOR U189 ( .A(n124), .B(n125), .Z(n121) );
  ANDN U190 ( .B(n126), .A(n127), .Z(n124) );
  XNOR U191 ( .A(b[34]), .B(n125), .Z(n126) );
  XNOR U192 ( .A(b[34]), .B(n127), .Z(c[34]) );
  XOR U193 ( .A(n128), .B(n129), .Z(n125) );
  ANDN U194 ( .B(n130), .A(n131), .Z(n128) );
  XNOR U195 ( .A(b[33]), .B(n129), .Z(n130) );
  XNOR U196 ( .A(b[33]), .B(n131), .Z(c[33]) );
  XOR U197 ( .A(n132), .B(n133), .Z(n129) );
  ANDN U198 ( .B(n134), .A(n135), .Z(n132) );
  XNOR U199 ( .A(b[32]), .B(n133), .Z(n134) );
  XNOR U200 ( .A(b[32]), .B(n135), .Z(c[32]) );
  XOR U201 ( .A(n136), .B(n137), .Z(n133) );
  ANDN U202 ( .B(n138), .A(n139), .Z(n136) );
  XNOR U203 ( .A(b[31]), .B(n137), .Z(n138) );
  XNOR U204 ( .A(b[31]), .B(n139), .Z(c[31]) );
  XOR U205 ( .A(n140), .B(n141), .Z(n137) );
  ANDN U206 ( .B(n142), .A(n143), .Z(n140) );
  XNOR U207 ( .A(b[30]), .B(n141), .Z(n142) );
  XNOR U208 ( .A(b[30]), .B(n143), .Z(c[30]) );
  XOR U209 ( .A(n144), .B(n145), .Z(n141) );
  ANDN U210 ( .B(n146), .A(n147), .Z(n144) );
  XNOR U211 ( .A(b[29]), .B(n145), .Z(n146) );
  XNOR U212 ( .A(b[2]), .B(n148), .Z(c[2]) );
  XNOR U213 ( .A(b[29]), .B(n147), .Z(c[29]) );
  XOR U214 ( .A(n149), .B(n150), .Z(n145) );
  ANDN U215 ( .B(n151), .A(n152), .Z(n149) );
  XNOR U216 ( .A(b[28]), .B(n150), .Z(n151) );
  XNOR U217 ( .A(b[28]), .B(n152), .Z(c[28]) );
  XOR U218 ( .A(n153), .B(n154), .Z(n150) );
  ANDN U219 ( .B(n155), .A(n156), .Z(n153) );
  XNOR U220 ( .A(b[27]), .B(n154), .Z(n155) );
  XNOR U221 ( .A(b[27]), .B(n156), .Z(c[27]) );
  XOR U222 ( .A(n157), .B(n158), .Z(n154) );
  ANDN U223 ( .B(n159), .A(n160), .Z(n157) );
  XNOR U224 ( .A(b[26]), .B(n158), .Z(n159) );
  XNOR U225 ( .A(b[26]), .B(n160), .Z(c[26]) );
  XOR U226 ( .A(n161), .B(n162), .Z(n158) );
  ANDN U227 ( .B(n163), .A(n164), .Z(n161) );
  XNOR U228 ( .A(b[25]), .B(n162), .Z(n163) );
  XNOR U229 ( .A(b[25]), .B(n164), .Z(c[25]) );
  XOR U230 ( .A(n165), .B(n166), .Z(n162) );
  ANDN U231 ( .B(n167), .A(n168), .Z(n165) );
  XNOR U232 ( .A(b[24]), .B(n166), .Z(n167) );
  XNOR U233 ( .A(b[24]), .B(n168), .Z(c[24]) );
  XOR U234 ( .A(n169), .B(n170), .Z(n166) );
  ANDN U235 ( .B(n171), .A(n172), .Z(n169) );
  XNOR U236 ( .A(b[23]), .B(n170), .Z(n171) );
  XNOR U237 ( .A(b[23]), .B(n172), .Z(c[23]) );
  XOR U238 ( .A(n173), .B(n174), .Z(n170) );
  ANDN U239 ( .B(n175), .A(n176), .Z(n173) );
  XNOR U240 ( .A(b[22]), .B(n174), .Z(n175) );
  XNOR U241 ( .A(b[22]), .B(n176), .Z(c[22]) );
  XOR U242 ( .A(n177), .B(n178), .Z(n174) );
  ANDN U243 ( .B(n179), .A(n180), .Z(n177) );
  XNOR U244 ( .A(b[21]), .B(n178), .Z(n179) );
  XNOR U245 ( .A(b[21]), .B(n180), .Z(c[21]) );
  XOR U246 ( .A(n181), .B(n182), .Z(n178) );
  ANDN U247 ( .B(n183), .A(n184), .Z(n181) );
  XNOR U248 ( .A(b[20]), .B(n182), .Z(n183) );
  XNOR U249 ( .A(b[20]), .B(n184), .Z(c[20]) );
  XOR U250 ( .A(n185), .B(n186), .Z(n182) );
  ANDN U251 ( .B(n187), .A(n188), .Z(n185) );
  XNOR U252 ( .A(b[19]), .B(n186), .Z(n187) );
  XNOR U253 ( .A(b[1]), .B(n189), .Z(c[1]) );
  XNOR U254 ( .A(b[19]), .B(n188), .Z(c[19]) );
  XOR U255 ( .A(n190), .B(n191), .Z(n186) );
  ANDN U256 ( .B(n192), .A(n193), .Z(n190) );
  XNOR U257 ( .A(b[18]), .B(n191), .Z(n192) );
  XNOR U258 ( .A(b[18]), .B(n193), .Z(c[18]) );
  XOR U259 ( .A(n194), .B(n195), .Z(n191) );
  ANDN U260 ( .B(n196), .A(n197), .Z(n194) );
  XNOR U261 ( .A(b[17]), .B(n195), .Z(n196) );
  XNOR U262 ( .A(b[17]), .B(n197), .Z(c[17]) );
  XOR U263 ( .A(n198), .B(n199), .Z(n195) );
  ANDN U264 ( .B(n200), .A(n201), .Z(n198) );
  XNOR U265 ( .A(b[16]), .B(n199), .Z(n200) );
  XNOR U266 ( .A(b[16]), .B(n201), .Z(c[16]) );
  XOR U267 ( .A(n202), .B(n203), .Z(n199) );
  ANDN U268 ( .B(n204), .A(n205), .Z(n202) );
  XNOR U269 ( .A(b[15]), .B(n203), .Z(n204) );
  XNOR U270 ( .A(b[15]), .B(n205), .Z(c[15]) );
  XOR U271 ( .A(n206), .B(n207), .Z(n203) );
  ANDN U272 ( .B(n208), .A(n209), .Z(n206) );
  XNOR U273 ( .A(b[14]), .B(n207), .Z(n208) );
  XNOR U274 ( .A(b[14]), .B(n209), .Z(c[14]) );
  XOR U275 ( .A(n210), .B(n211), .Z(n207) );
  ANDN U276 ( .B(n212), .A(n213), .Z(n210) );
  XNOR U277 ( .A(b[13]), .B(n211), .Z(n212) );
  XNOR U278 ( .A(b[13]), .B(n213), .Z(c[13]) );
  XOR U279 ( .A(n214), .B(n215), .Z(n211) );
  ANDN U280 ( .B(n216), .A(n217), .Z(n214) );
  XNOR U281 ( .A(b[12]), .B(n215), .Z(n216) );
  XNOR U282 ( .A(b[12]), .B(n217), .Z(c[12]) );
  XOR U283 ( .A(n218), .B(n219), .Z(n215) );
  ANDN U284 ( .B(n220), .A(n221), .Z(n218) );
  XNOR U285 ( .A(b[11]), .B(n219), .Z(n220) );
  XNOR U286 ( .A(b[11]), .B(n221), .Z(c[11]) );
  XOR U287 ( .A(n222), .B(n223), .Z(n219) );
  ANDN U288 ( .B(n224), .A(n225), .Z(n222) );
  XNOR U289 ( .A(b[10]), .B(n223), .Z(n224) );
  XNOR U290 ( .A(b[10]), .B(n225), .Z(c[10]) );
  XOR U291 ( .A(n226), .B(n227), .Z(n223) );
  ANDN U292 ( .B(n228), .A(n5), .Z(n226) );
  XNOR U293 ( .A(b[9]), .B(n227), .Z(n228) );
  XOR U294 ( .A(n229), .B(n230), .Z(n227) );
  ANDN U295 ( .B(n231), .A(n6), .Z(n229) );
  XNOR U296 ( .A(b[8]), .B(n230), .Z(n231) );
  XOR U297 ( .A(n232), .B(n233), .Z(n230) );
  ANDN U298 ( .B(n234), .A(n7), .Z(n232) );
  XNOR U299 ( .A(b[7]), .B(n233), .Z(n234) );
  XOR U300 ( .A(n235), .B(n236), .Z(n233) );
  ANDN U301 ( .B(n237), .A(n8), .Z(n235) );
  XNOR U302 ( .A(b[6]), .B(n236), .Z(n237) );
  XOR U303 ( .A(n238), .B(n239), .Z(n236) );
  ANDN U304 ( .B(n240), .A(n25), .Z(n238) );
  XNOR U305 ( .A(b[5]), .B(n239), .Z(n240) );
  XOR U306 ( .A(n241), .B(n242), .Z(n239) );
  ANDN U307 ( .B(n243), .A(n66), .Z(n241) );
  XNOR U308 ( .A(b[4]), .B(n242), .Z(n243) );
  XOR U309 ( .A(n244), .B(n245), .Z(n242) );
  ANDN U310 ( .B(n246), .A(n107), .Z(n244) );
  XNOR U311 ( .A(b[3]), .B(n245), .Z(n246) );
  XOR U312 ( .A(n247), .B(n248), .Z(n245) );
  ANDN U313 ( .B(n249), .A(n148), .Z(n247) );
  XNOR U314 ( .A(b[2]), .B(n248), .Z(n249) );
  XOR U315 ( .A(n250), .B(n251), .Z(n248) );
  ANDN U316 ( .B(n252), .A(n189), .Z(n250) );
  XNOR U317 ( .A(b[1]), .B(n251), .Z(n252) );
  XOR U318 ( .A(carry_on), .B(n253), .Z(n251) );
  NANDN U319 ( .A(n254), .B(n255), .Z(n253) );
  XOR U320 ( .A(carry_on), .B(b[0]), .Z(n255) );
  XNOR U321 ( .A(b[0]), .B(n254), .Z(c[0]) );
  XNOR U322 ( .A(a[0]), .B(carry_on), .Z(n254) );
endmodule

