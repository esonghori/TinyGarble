
module hamming_N160_CC1 ( clk, rst, x, y, o );
  input [159:0] x;
  input [159:0] y;
  output [7:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988;

  NAND U161 ( .A(n257), .B(n256), .Z(n1) );
  XOR U162 ( .A(n256), .B(n257), .Z(n2) );
  NANDN U163 ( .A(n255), .B(n2), .Z(n3) );
  NAND U164 ( .A(n1), .B(n3), .Z(n575) );
  NAND U165 ( .A(n597), .B(n596), .Z(n4) );
  XOR U166 ( .A(n596), .B(n597), .Z(n5) );
  NANDN U167 ( .A(n595), .B(n5), .Z(n6) );
  NAND U168 ( .A(n4), .B(n6), .Z(n799) );
  NAND U169 ( .A(n454), .B(n453), .Z(n7) );
  XOR U170 ( .A(n453), .B(n454), .Z(n8) );
  NANDN U171 ( .A(n452), .B(n8), .Z(n9) );
  NAND U172 ( .A(n7), .B(n9), .Z(n617) );
  XOR U173 ( .A(n501), .B(n499), .Z(n10) );
  NANDN U174 ( .A(n500), .B(n10), .Z(n11) );
  NAND U175 ( .A(n501), .B(n499), .Z(n12) );
  AND U176 ( .A(n11), .B(n12), .Z(n641) );
  XNOR U177 ( .A(n672), .B(n673), .Z(n576) );
  XNOR U178 ( .A(n752), .B(n754), .Z(n13) );
  XNOR U179 ( .A(n753), .B(n13), .Z(n771) );
  XOR U180 ( .A(n801), .B(n800), .Z(n14) );
  NANDN U181 ( .A(n799), .B(n14), .Z(n15) );
  NAND U182 ( .A(n801), .B(n800), .Z(n16) );
  AND U183 ( .A(n15), .B(n16), .Z(n890) );
  XNOR U184 ( .A(n550), .B(n551), .Z(n366) );
  XNOR U185 ( .A(n663), .B(n664), .Z(n616) );
  NAND U186 ( .A(n149), .B(n147), .Z(n17) );
  XOR U187 ( .A(n147), .B(n149), .Z(n18) );
  NANDN U188 ( .A(n148), .B(n18), .Z(n19) );
  NAND U189 ( .A(n17), .B(n19), .Z(n604) );
  OR U190 ( .A(n248), .B(n247), .Z(n20) );
  NANDN U191 ( .A(n250), .B(n249), .Z(n21) );
  NAND U192 ( .A(n20), .B(n21), .Z(n734) );
  XNOR U193 ( .A(n706), .B(n707), .Z(n643) );
  XNOR U194 ( .A(n824), .B(n825), .Z(n851) );
  XOR U195 ( .A(n586), .B(n585), .Z(n22) );
  NANDN U196 ( .A(n584), .B(n22), .Z(n23) );
  NAND U197 ( .A(n586), .B(n585), .Z(n24) );
  AND U198 ( .A(n23), .B(n24), .Z(n837) );
  XOR U199 ( .A(n409), .B(n408), .Z(n25) );
  NANDN U200 ( .A(n407), .B(n25), .Z(n26) );
  NAND U201 ( .A(n409), .B(n408), .Z(n27) );
  AND U202 ( .A(n26), .B(n27), .Z(n591) );
  XOR U203 ( .A(n800), .B(n799), .Z(n28) );
  XNOR U204 ( .A(n801), .B(n28), .Z(n886) );
  NAND U205 ( .A(n771), .B(n769), .Z(n29) );
  XOR U206 ( .A(n769), .B(n771), .Z(n30) );
  NANDN U207 ( .A(n770), .B(n30), .Z(n31) );
  NAND U208 ( .A(n29), .B(n31), .Z(n881) );
  XNOR U209 ( .A(n722), .B(n723), .Z(n624) );
  NAND U210 ( .A(n541), .B(n539), .Z(n32) );
  XOR U211 ( .A(n539), .B(n541), .Z(n33) );
  NANDN U212 ( .A(n540), .B(n33), .Z(n34) );
  NAND U213 ( .A(n32), .B(n34), .Z(n599) );
  XNOR U214 ( .A(n642), .B(n643), .Z(n35) );
  XNOR U215 ( .A(n641), .B(n35), .Z(n755) );
  NAND U216 ( .A(n614), .B(n613), .Z(n36) );
  XOR U217 ( .A(n613), .B(n614), .Z(n37) );
  NANDN U218 ( .A(n615), .B(n37), .Z(n38) );
  NAND U219 ( .A(n36), .B(n38), .Z(n843) );
  XOR U220 ( .A(n612), .B(n610), .Z(n39) );
  NANDN U221 ( .A(n611), .B(n39), .Z(n40) );
  NAND U222 ( .A(n612), .B(n610), .Z(n41) );
  AND U223 ( .A(n40), .B(n41), .Z(n802) );
  NAND U224 ( .A(n719), .B(n717), .Z(n42) );
  XOR U225 ( .A(n717), .B(n719), .Z(n43) );
  NANDN U226 ( .A(n718), .B(n43), .Z(n44) );
  NAND U227 ( .A(n42), .B(n44), .Z(n854) );
  NAND U228 ( .A(n669), .B(n667), .Z(n45) );
  XOR U229 ( .A(n667), .B(n669), .Z(n46) );
  NANDN U230 ( .A(n668), .B(n46), .Z(n47) );
  NAND U231 ( .A(n45), .B(n47), .Z(n822) );
  XOR U232 ( .A(n583), .B(n582), .Z(n48) );
  NANDN U233 ( .A(n581), .B(n48), .Z(n49) );
  NAND U234 ( .A(n583), .B(n582), .Z(n50) );
  AND U235 ( .A(n49), .B(n50), .Z(n836) );
  NAND U236 ( .A(n647), .B(n646), .Z(n51) );
  XOR U237 ( .A(n646), .B(n647), .Z(n52) );
  NANDN U238 ( .A(n645), .B(n52), .Z(n53) );
  NAND U239 ( .A(n51), .B(n53), .Z(n875) );
  NAND U240 ( .A(n576), .B(n575), .Z(n54) );
  XOR U241 ( .A(n575), .B(n576), .Z(n55) );
  NANDN U242 ( .A(n574), .B(n55), .Z(n56) );
  NAND U243 ( .A(n54), .B(n56), .Z(n809) );
  XOR U244 ( .A(n830), .B(n831), .Z(n832) );
  XNOR U245 ( .A(n535), .B(n536), .Z(n457) );
  XOR U246 ( .A(n593), .B(n591), .Z(n57) );
  NAND U247 ( .A(n57), .B(n592), .Z(n58) );
  NAND U248 ( .A(n593), .B(n591), .Z(n59) );
  AND U249 ( .A(n58), .B(n59), .Z(n784) );
  NAND U250 ( .A(n754), .B(n752), .Z(n60) );
  XOR U251 ( .A(n752), .B(n754), .Z(n61) );
  NANDN U252 ( .A(n753), .B(n61), .Z(n62) );
  NAND U253 ( .A(n60), .B(n62), .Z(n794) );
  XNOR U254 ( .A(n880), .B(n881), .Z(n883) );
  NAND U255 ( .A(n888), .B(n887), .Z(n63) );
  XOR U256 ( .A(n887), .B(n888), .Z(n64) );
  NANDN U257 ( .A(n886), .B(n64), .Z(n65) );
  NAND U258 ( .A(n63), .B(n65), .Z(n940) );
  XNOR U259 ( .A(n656), .B(n657), .Z(n605) );
  XNOR U260 ( .A(n698), .B(n699), .Z(n601) );
  OR U261 ( .A(n252), .B(n251), .Z(n66) );
  NANDN U262 ( .A(n254), .B(n253), .Z(n67) );
  NAND U263 ( .A(n66), .B(n67), .Z(n733) );
  NAND U264 ( .A(n405), .B(n404), .Z(n68) );
  XOR U265 ( .A(n404), .B(n405), .Z(n69) );
  NANDN U266 ( .A(n406), .B(n69), .Z(n70) );
  NAND U267 ( .A(n68), .B(n70), .Z(n568) );
  XNOR U268 ( .A(n678), .B(n679), .Z(n618) );
  XOR U269 ( .A(n624), .B(n625), .Z(n756) );
  NANDN U270 ( .A(n580), .B(n579), .Z(n71) );
  NANDN U271 ( .A(n578), .B(n577), .Z(n72) );
  NAND U272 ( .A(n71), .B(n72), .Z(n838) );
  NAND U273 ( .A(n643), .B(n642), .Z(n73) );
  XOR U274 ( .A(n642), .B(n643), .Z(n74) );
  NANDN U275 ( .A(n641), .B(n74), .Z(n75) );
  NAND U276 ( .A(n73), .B(n75), .Z(n817) );
  XNOR U277 ( .A(n305), .B(n306), .Z(n308) );
  XOR U278 ( .A(n319), .B(n317), .Z(n76) );
  NANDN U279 ( .A(n318), .B(n76), .Z(n77) );
  NAND U280 ( .A(n319), .B(n317), .Z(n78) );
  AND U281 ( .A(n77), .B(n78), .Z(n614) );
  XOR U282 ( .A(n210), .B(n208), .Z(n79) );
  NANDN U283 ( .A(n209), .B(n79), .Z(n80) );
  NAND U284 ( .A(n210), .B(n208), .Z(n81) );
  AND U285 ( .A(n80), .B(n81), .Z(n753) );
  NAND U286 ( .A(n590), .B(n589), .Z(n82) );
  XOR U287 ( .A(n589), .B(n590), .Z(n83) );
  NAND U288 ( .A(n83), .B(n588), .Z(n84) );
  NAND U289 ( .A(n82), .B(n84), .Z(n787) );
  NAND U290 ( .A(n852), .B(n851), .Z(n85) );
  XOR U291 ( .A(n851), .B(n852), .Z(n86) );
  NANDN U292 ( .A(n853), .B(n86), .Z(n87) );
  NAND U293 ( .A(n85), .B(n87), .Z(n903) );
  XNOR U294 ( .A(n921), .B(n920), .Z(n919) );
  XOR U295 ( .A(n780), .B(n781), .Z(n887) );
  XNOR U296 ( .A(n301), .B(n300), .Z(n104) );
  XNOR U297 ( .A(n764), .B(n763), .Z(n765) );
  XOR U298 ( .A(n954), .B(n953), .Z(n88) );
  NANDN U299 ( .A(n952), .B(n88), .Z(n89) );
  NAND U300 ( .A(n954), .B(n953), .Z(n90) );
  AND U301 ( .A(n89), .B(n90), .Z(n975) );
  XNOR U302 ( .A(n883), .B(n882), .Z(n775) );
  XNOR U303 ( .A(x[84]), .B(y[84]), .Z(n132) );
  XNOR U304 ( .A(x[158]), .B(y[158]), .Z(n130) );
  XNOR U305 ( .A(x[82]), .B(y[82]), .Z(n129) );
  XNOR U306 ( .A(n130), .B(n129), .Z(n131) );
  XOR U307 ( .A(n132), .B(n131), .Z(n502) );
  IV U308 ( .A(n502), .Z(n503) );
  XNOR U309 ( .A(x[74]), .B(y[74]), .Z(n138) );
  XNOR U310 ( .A(x[72]), .B(y[72]), .Z(n136) );
  XNOR U311 ( .A(x[70]), .B(y[70]), .Z(n135) );
  XNOR U312 ( .A(n136), .B(n135), .Z(n137) );
  XOR U313 ( .A(n138), .B(n137), .Z(n506) );
  XNOR U314 ( .A(x[80]), .B(y[80]), .Z(n144) );
  XNOR U315 ( .A(x[78]), .B(y[78]), .Z(n142) );
  XNOR U316 ( .A(x[76]), .B(y[76]), .Z(n141) );
  XNOR U317 ( .A(n142), .B(n141), .Z(n143) );
  XOR U318 ( .A(n144), .B(n143), .Z(n504) );
  XNOR U319 ( .A(n506), .B(n504), .Z(n91) );
  XNOR U320 ( .A(n503), .B(n91), .Z(n262) );
  XNOR U321 ( .A(x[88]), .B(y[88]), .Z(n177) );
  XNOR U322 ( .A(x[156]), .B(y[156]), .Z(n175) );
  XNOR U323 ( .A(x[86]), .B(y[86]), .Z(n174) );
  XNOR U324 ( .A(n175), .B(n174), .Z(n176) );
  XOR U325 ( .A(n177), .B(n176), .Z(n269) );
  XNOR U326 ( .A(x[96]), .B(y[96]), .Z(n171) );
  XNOR U327 ( .A(x[152]), .B(y[152]), .Z(n169) );
  XNOR U328 ( .A(x[94]), .B(y[94]), .Z(n168) );
  XNOR U329 ( .A(n169), .B(n168), .Z(n170) );
  XNOR U330 ( .A(n171), .B(n170), .Z(n266) );
  IV U331 ( .A(n266), .Z(n265) );
  XNOR U332 ( .A(x[92]), .B(y[92]), .Z(n183) );
  XNOR U333 ( .A(x[154]), .B(y[154]), .Z(n181) );
  XNOR U334 ( .A(x[90]), .B(y[90]), .Z(n180) );
  XNOR U335 ( .A(n181), .B(n180), .Z(n182) );
  XOR U336 ( .A(n183), .B(n182), .Z(n267) );
  XNOR U337 ( .A(n265), .B(n267), .Z(n92) );
  XOR U338 ( .A(n269), .B(n92), .Z(n259) );
  XNOR U339 ( .A(x[104]), .B(y[104]), .Z(n336) );
  XNOR U340 ( .A(x[102]), .B(y[102]), .Z(n333) );
  XNOR U341 ( .A(x[148]), .B(y[148]), .Z(n334) );
  XOR U342 ( .A(n333), .B(n334), .Z(n335) );
  XOR U343 ( .A(n336), .B(n335), .Z(n257) );
  XNOR U344 ( .A(x[108]), .B(y[108]), .Z(n324) );
  XNOR U345 ( .A(x[146]), .B(y[146]), .Z(n322) );
  XNOR U346 ( .A(x[106]), .B(y[106]), .Z(n321) );
  XOR U347 ( .A(n322), .B(n321), .Z(n323) );
  XNOR U348 ( .A(n324), .B(n323), .Z(n255) );
  XNOR U349 ( .A(x[100]), .B(y[100]), .Z(n330) );
  XNOR U350 ( .A(x[150]), .B(y[150]), .Z(n328) );
  XNOR U351 ( .A(x[98]), .B(y[98]), .Z(n327) );
  XOR U352 ( .A(n328), .B(n327), .Z(n329) );
  XOR U353 ( .A(n330), .B(n329), .Z(n256) );
  XOR U354 ( .A(n255), .B(n256), .Z(n93) );
  XNOR U355 ( .A(n257), .B(n93), .Z(n260) );
  XOR U356 ( .A(n259), .B(n260), .Z(n261) );
  XNOR U357 ( .A(n262), .B(n261), .Z(n301) );
  XNOR U358 ( .A(x[2]), .B(y[2]), .Z(n477) );
  XNOR U359 ( .A(x[1]), .B(y[1]), .Z(n475) );
  XNOR U360 ( .A(x[0]), .B(y[0]), .Z(n474) );
  XOR U361 ( .A(n475), .B(n474), .Z(n476) );
  XNOR U362 ( .A(n477), .B(n476), .Z(n454) );
  XNOR U363 ( .A(x[14]), .B(y[14]), .Z(n419) );
  XNOR U364 ( .A(x[12]), .B(y[12]), .Z(n417) );
  XNOR U365 ( .A(x[10]), .B(y[10]), .Z(n416) );
  XNOR U366 ( .A(n417), .B(n416), .Z(n418) );
  XNOR U367 ( .A(n419), .B(n418), .Z(n452) );
  XNOR U368 ( .A(x[8]), .B(y[8]), .Z(n425) );
  XNOR U369 ( .A(x[6]), .B(y[6]), .Z(n423) );
  XNOR U370 ( .A(x[4]), .B(y[4]), .Z(n422) );
  XNOR U371 ( .A(n423), .B(n422), .Z(n424) );
  XOR U372 ( .A(n425), .B(n424), .Z(n453) );
  XOR U373 ( .A(n452), .B(n453), .Z(n94) );
  XOR U374 ( .A(n454), .B(n94), .Z(n210) );
  XNOR U375 ( .A(x[3]), .B(y[3]), .Z(n471) );
  XNOR U376 ( .A(x[7]), .B(y[7]), .Z(n469) );
  XNOR U377 ( .A(x[5]), .B(y[5]), .Z(n468) );
  XOR U378 ( .A(n469), .B(n468), .Z(n470) );
  XOR U379 ( .A(n471), .B(n470), .Z(n368) );
  XNOR U380 ( .A(x[9]), .B(y[9]), .Z(n545) );
  XNOR U381 ( .A(x[13]), .B(y[13]), .Z(n543) );
  XNOR U382 ( .A(x[11]), .B(y[11]), .Z(n542) );
  XOR U383 ( .A(n543), .B(n542), .Z(n544) );
  XOR U384 ( .A(n545), .B(n544), .Z(n367) );
  XNOR U385 ( .A(x[19]), .B(y[19]), .Z(n548) );
  XNOR U386 ( .A(x[17]), .B(y[17]), .Z(n549) );
  XNOR U387 ( .A(n548), .B(n549), .Z(n550) );
  XNOR U388 ( .A(x[15]), .B(y[15]), .Z(n551) );
  XOR U389 ( .A(n367), .B(n366), .Z(n369) );
  XNOR U390 ( .A(n368), .B(n369), .Z(n209) );
  XNOR U391 ( .A(x[21]), .B(y[21]), .Z(n518) );
  XNOR U392 ( .A(x[25]), .B(y[25]), .Z(n516) );
  XNOR U393 ( .A(x[23]), .B(y[23]), .Z(n515) );
  XOR U394 ( .A(n516), .B(n515), .Z(n517) );
  XOR U395 ( .A(n518), .B(n517), .Z(n313) );
  XNOR U396 ( .A(x[33]), .B(y[33]), .Z(n226) );
  XNOR U397 ( .A(x[37]), .B(y[37]), .Z(n224) );
  XNOR U398 ( .A(x[35]), .B(y[35]), .Z(n223) );
  XNOR U399 ( .A(n224), .B(n223), .Z(n225) );
  XNOR U400 ( .A(n226), .B(n225), .Z(n312) );
  XNOR U401 ( .A(x[27]), .B(y[27]), .Z(n524) );
  XNOR U402 ( .A(x[31]), .B(y[31]), .Z(n522) );
  XNOR U403 ( .A(x[29]), .B(y[29]), .Z(n521) );
  XOR U404 ( .A(n522), .B(n521), .Z(n523) );
  XOR U405 ( .A(n524), .B(n523), .Z(n311) );
  XOR U406 ( .A(n312), .B(n311), .Z(n314) );
  XOR U407 ( .A(n313), .B(n314), .Z(n208) );
  XOR U408 ( .A(n209), .B(n208), .Z(n95) );
  XOR U409 ( .A(n210), .B(n95), .Z(n299) );
  XNOR U410 ( .A(x[99]), .B(y[99]), .Z(n232) );
  XNOR U411 ( .A(x[103]), .B(y[103]), .Z(n230) );
  XNOR U412 ( .A(x[101]), .B(y[101]), .Z(n229) );
  XNOR U413 ( .A(n230), .B(n229), .Z(n231) );
  XNOR U414 ( .A(n232), .B(n231), .Z(n319) );
  XNOR U415 ( .A(x[149]), .B(y[149]), .Z(n387) );
  XNOR U416 ( .A(x[159]), .B(y[159]), .Z(n385) );
  XNOR U417 ( .A(x[153]), .B(y[153]), .Z(n384) );
  XNOR U418 ( .A(n385), .B(n384), .Z(n386) );
  XNOR U419 ( .A(n387), .B(n386), .Z(n317) );
  XNOR U420 ( .A(x[93]), .B(y[93]), .Z(n483) );
  XNOR U421 ( .A(x[97]), .B(y[97]), .Z(n481) );
  XNOR U422 ( .A(x[95]), .B(y[95]), .Z(n480) );
  XNOR U423 ( .A(n481), .B(n480), .Z(n482) );
  XOR U424 ( .A(n483), .B(n482), .Z(n318) );
  XOR U425 ( .A(n317), .B(n318), .Z(n96) );
  XNOR U426 ( .A(n319), .B(n96), .Z(n563) );
  XNOR U427 ( .A(x[117]), .B(y[117]), .Z(n530) );
  XNOR U428 ( .A(x[121]), .B(y[121]), .Z(n528) );
  XNOR U429 ( .A(x[119]), .B(y[119]), .Z(n527) );
  XNOR U430 ( .A(n528), .B(n527), .Z(n529) );
  XNOR U431 ( .A(n530), .B(n529), .Z(n149) );
  XNOR U432 ( .A(x[141]), .B(y[141]), .Z(n437) );
  XNOR U433 ( .A(x[145]), .B(y[145]), .Z(n435) );
  XNOR U434 ( .A(x[143]), .B(y[143]), .Z(n434) );
  XNOR U435 ( .A(n435), .B(n434), .Z(n436) );
  XNOR U436 ( .A(n437), .B(n436), .Z(n147) );
  XNOR U437 ( .A(x[123]), .B(y[123]), .Z(n557) );
  XNOR U438 ( .A(x[127]), .B(y[127]), .Z(n555) );
  XNOR U439 ( .A(x[125]), .B(y[125]), .Z(n554) );
  XNOR U440 ( .A(n555), .B(n554), .Z(n556) );
  XOR U441 ( .A(n557), .B(n556), .Z(n148) );
  XOR U442 ( .A(n147), .B(n148), .Z(n97) );
  XOR U443 ( .A(n149), .B(n97), .Z(n561) );
  XNOR U444 ( .A(x[57]), .B(y[57]), .Z(n238) );
  XNOR U445 ( .A(x[59]), .B(y[59]), .Z(n236) );
  XNOR U446 ( .A(x[61]), .B(y[61]), .Z(n235) );
  XNOR U447 ( .A(n236), .B(n235), .Z(n237) );
  XOR U448 ( .A(n238), .B(n237), .Z(n400) );
  XNOR U449 ( .A(x[63]), .B(y[63]), .Z(n244) );
  XNOR U450 ( .A(x[65]), .B(y[65]), .Z(n242) );
  XNOR U451 ( .A(x[67]), .B(y[67]), .Z(n241) );
  XNOR U452 ( .A(n242), .B(n241), .Z(n243) );
  XOR U453 ( .A(n244), .B(n243), .Z(n398) );
  XNOR U454 ( .A(x[69]), .B(y[69]), .Z(n495) );
  XNOR U455 ( .A(x[73]), .B(y[73]), .Z(n493) );
  XNOR U456 ( .A(x[71]), .B(y[71]), .Z(n492) );
  XNOR U457 ( .A(n493), .B(n492), .Z(n494) );
  XOR U458 ( .A(n495), .B(n494), .Z(n399) );
  XNOR U459 ( .A(n398), .B(n399), .Z(n401) );
  XOR U460 ( .A(n400), .B(n401), .Z(n562) );
  XNOR U461 ( .A(n561), .B(n562), .Z(n98) );
  XNOR U462 ( .A(n563), .B(n98), .Z(n298) );
  XOR U463 ( .A(n299), .B(n298), .Z(n300) );
  XNOR U464 ( .A(x[129]), .B(y[129]), .Z(n465) );
  XNOR U465 ( .A(x[133]), .B(y[133]), .Z(n462) );
  XNOR U466 ( .A(x[131]), .B(y[131]), .Z(n463) );
  XOR U467 ( .A(n462), .B(n463), .Z(n464) );
  XOR U468 ( .A(n465), .B(n464), .Z(n272) );
  XNOR U469 ( .A(x[135]), .B(y[135]), .Z(n431) );
  XNOR U470 ( .A(x[137]), .B(y[137]), .Z(n428) );
  XNOR U471 ( .A(x[139]), .B(y[139]), .Z(n429) );
  XOR U472 ( .A(n428), .B(n429), .Z(n430) );
  XNOR U473 ( .A(n431), .B(n430), .Z(n273) );
  XNOR U474 ( .A(n272), .B(n273), .Z(n274) );
  XNOR U475 ( .A(x[157]), .B(y[157]), .Z(n199) );
  XNOR U476 ( .A(x[155]), .B(y[155]), .Z(n200) );
  XNOR U477 ( .A(n199), .B(n200), .Z(n381) );
  XNOR U478 ( .A(x[151]), .B(y[151]), .Z(n379) );
  XNOR U479 ( .A(x[147]), .B(y[147]), .Z(n378) );
  XOR U480 ( .A(n379), .B(n378), .Z(n380) );
  XOR U481 ( .A(n381), .B(n380), .Z(n372) );
  XNOR U482 ( .A(x[111]), .B(y[111]), .Z(n214) );
  XNOR U483 ( .A(x[115]), .B(y[115]), .Z(n211) );
  XNOR U484 ( .A(x[113]), .B(y[113]), .Z(n212) );
  XOR U485 ( .A(n211), .B(n212), .Z(n213) );
  XNOR U486 ( .A(n214), .B(n213), .Z(n373) );
  XNOR U487 ( .A(n372), .B(n373), .Z(n374) );
  XNOR U488 ( .A(x[105]), .B(y[105]), .Z(n293) );
  XNOR U489 ( .A(x[109]), .B(y[109]), .Z(n291) );
  XNOR U490 ( .A(x[107]), .B(y[107]), .Z(n290) );
  XNOR U491 ( .A(n291), .B(n290), .Z(n292) );
  XNOR U492 ( .A(n293), .B(n292), .Z(n375) );
  XNOR U493 ( .A(n374), .B(n375), .Z(n275) );
  XOR U494 ( .A(n274), .B(n275), .Z(n409) );
  XNOR U495 ( .A(x[75]), .B(y[75]), .Z(n254) );
  XNOR U496 ( .A(x[79]), .B(y[79]), .Z(n252) );
  XNOR U497 ( .A(x[77]), .B(y[77]), .Z(n251) );
  XOR U498 ( .A(n252), .B(n251), .Z(n253) );
  XNOR U499 ( .A(n254), .B(n253), .Z(n307) );
  XNOR U500 ( .A(x[87]), .B(y[87]), .Z(n489) );
  XNOR U501 ( .A(x[91]), .B(y[91]), .Z(n486) );
  XNOR U502 ( .A(x[89]), .B(y[89]), .Z(n487) );
  XOR U503 ( .A(n486), .B(n487), .Z(n488) );
  XNOR U504 ( .A(n489), .B(n488), .Z(n305) );
  XNOR U505 ( .A(x[81]), .B(y[81]), .Z(n250) );
  XNOR U506 ( .A(x[85]), .B(y[85]), .Z(n248) );
  XNOR U507 ( .A(x[83]), .B(y[83]), .Z(n247) );
  XOR U508 ( .A(n248), .B(n247), .Z(n249) );
  XNOR U509 ( .A(n250), .B(n249), .Z(n306) );
  XOR U510 ( .A(n307), .B(n308), .Z(n407) );
  XNOR U511 ( .A(x[51]), .B(y[51]), .Z(n281) );
  XNOR U512 ( .A(x[55]), .B(y[55]), .Z(n279) );
  XNOR U513 ( .A(x[53]), .B(y[53]), .Z(n278) );
  XNOR U514 ( .A(n279), .B(n278), .Z(n280) );
  XOR U515 ( .A(n281), .B(n280), .Z(n406) );
  XNOR U516 ( .A(x[39]), .B(y[39]), .Z(n220) );
  XNOR U517 ( .A(x[43]), .B(y[43]), .Z(n217) );
  XNOR U518 ( .A(x[41]), .B(y[41]), .Z(n218) );
  XOR U519 ( .A(n217), .B(n218), .Z(n219) );
  XOR U520 ( .A(n220), .B(n219), .Z(n404) );
  XNOR U521 ( .A(x[45]), .B(y[45]), .Z(n287) );
  XNOR U522 ( .A(x[49]), .B(y[49]), .Z(n285) );
  XNOR U523 ( .A(x[47]), .B(y[47]), .Z(n284) );
  XNOR U524 ( .A(n285), .B(n284), .Z(n286) );
  XNOR U525 ( .A(n287), .B(n286), .Z(n405) );
  XNOR U526 ( .A(n404), .B(n405), .Z(n99) );
  XNOR U527 ( .A(n406), .B(n99), .Z(n408) );
  XOR U528 ( .A(n407), .B(n408), .Z(n100) );
  XOR U529 ( .A(n409), .B(n100), .Z(n105) );
  XOR U530 ( .A(n104), .B(n105), .Z(n106) );
  XNOR U531 ( .A(x[116]), .B(y[116]), .Z(n361) );
  XNOR U532 ( .A(x[142]), .B(y[142]), .Z(n359) );
  XNOR U533 ( .A(x[114]), .B(y[114]), .Z(n358) );
  XNOR U534 ( .A(n359), .B(n358), .Z(n360) );
  XOR U535 ( .A(n361), .B(n360), .Z(n541) );
  XNOR U536 ( .A(x[112]), .B(y[112]), .Z(n355) );
  XNOR U537 ( .A(x[144]), .B(y[144]), .Z(n353) );
  XNOR U538 ( .A(x[110]), .B(y[110]), .Z(n352) );
  XNOR U539 ( .A(n353), .B(n352), .Z(n354) );
  XNOR U540 ( .A(n355), .B(n354), .Z(n540) );
  XNOR U541 ( .A(x[128]), .B(y[128]), .Z(n196) );
  XNOR U542 ( .A(x[130]), .B(y[130]), .Z(n194) );
  XNOR U543 ( .A(x[126]), .B(y[126]), .Z(n193) );
  XNOR U544 ( .A(n194), .B(n193), .Z(n195) );
  XOR U545 ( .A(n196), .B(n195), .Z(n539) );
  XOR U546 ( .A(n540), .B(n539), .Z(n101) );
  XOR U547 ( .A(n541), .B(n101), .Z(n410) );
  XNOR U548 ( .A(x[132]), .B(y[132]), .Z(n204) );
  XNOR U549 ( .A(x[136]), .B(y[136]), .Z(n202) );
  XNOR U550 ( .A(x[134]), .B(y[134]), .Z(n201) );
  XNOR U551 ( .A(n202), .B(n201), .Z(n203) );
  XOR U552 ( .A(n204), .B(n203), .Z(n339) );
  IV U553 ( .A(n339), .Z(n340) );
  XNOR U554 ( .A(x[120]), .B(y[120]), .Z(n349) );
  XNOR U555 ( .A(x[140]), .B(y[140]), .Z(n347) );
  XNOR U556 ( .A(x[118]), .B(y[118]), .Z(n346) );
  XNOR U557 ( .A(n347), .B(n346), .Z(n348) );
  XNOR U558 ( .A(n349), .B(n348), .Z(n342) );
  XNOR U559 ( .A(x[124]), .B(y[124]), .Z(n190) );
  XNOR U560 ( .A(x[138]), .B(y[138]), .Z(n188) );
  XNOR U561 ( .A(x[122]), .B(y[122]), .Z(n187) );
  XNOR U562 ( .A(n188), .B(n187), .Z(n189) );
  XOR U563 ( .A(n190), .B(n189), .Z(n341) );
  XOR U564 ( .A(n342), .B(n341), .Z(n102) );
  XNOR U565 ( .A(n340), .B(n102), .Z(n411) );
  XOR U566 ( .A(n410), .B(n411), .Z(n412) );
  XNOR U567 ( .A(x[20]), .B(y[20]), .Z(n443) );
  XNOR U568 ( .A(x[18]), .B(y[18]), .Z(n441) );
  XNOR U569 ( .A(x[16]), .B(y[16]), .Z(n440) );
  XNOR U570 ( .A(n441), .B(n440), .Z(n442) );
  XNOR U571 ( .A(n443), .B(n442), .Z(n501) );
  XNOR U572 ( .A(x[32]), .B(y[32]), .Z(n393) );
  XNOR U573 ( .A(x[30]), .B(y[30]), .Z(n391) );
  XNOR U574 ( .A(x[28]), .B(y[28]), .Z(n390) );
  XNOR U575 ( .A(n391), .B(n390), .Z(n392) );
  XNOR U576 ( .A(n393), .B(n392), .Z(n499) );
  XNOR U577 ( .A(x[26]), .B(y[26]), .Z(n449) );
  XNOR U578 ( .A(x[24]), .B(y[24]), .Z(n447) );
  XNOR U579 ( .A(x[22]), .B(y[22]), .Z(n446) );
  XNOR U580 ( .A(n447), .B(n446), .Z(n448) );
  XOR U581 ( .A(n449), .B(n448), .Z(n500) );
  XOR U582 ( .A(n499), .B(n500), .Z(n103) );
  XNOR U583 ( .A(n501), .B(n103), .Z(n458) );
  XNOR U584 ( .A(x[50]), .B(y[50]), .Z(n125) );
  XNOR U585 ( .A(x[48]), .B(y[48]), .Z(n123) );
  XNOR U586 ( .A(x[46]), .B(y[46]), .Z(n122) );
  XNOR U587 ( .A(n123), .B(n122), .Z(n124) );
  XOR U588 ( .A(n125), .B(n124), .Z(n536) );
  XNOR U589 ( .A(x[44]), .B(y[44]), .Z(n119) );
  XNOR U590 ( .A(x[42]), .B(y[42]), .Z(n117) );
  XNOR U591 ( .A(x[40]), .B(y[40]), .Z(n116) );
  XNOR U592 ( .A(n117), .B(n116), .Z(n118) );
  XOR U593 ( .A(n119), .B(n118), .Z(n533) );
  XNOR U594 ( .A(x[38]), .B(y[38]), .Z(n113) );
  XNOR U595 ( .A(x[36]), .B(y[36]), .Z(n111) );
  XNOR U596 ( .A(x[34]), .B(y[34]), .Z(n110) );
  XNOR U597 ( .A(n111), .B(n110), .Z(n112) );
  XOR U598 ( .A(n113), .B(n112), .Z(n534) );
  XNOR U599 ( .A(n533), .B(n534), .Z(n535) );
  XNOR U600 ( .A(x[68]), .B(y[68]), .Z(n159) );
  XNOR U601 ( .A(x[66]), .B(y[66]), .Z(n157) );
  XNOR U602 ( .A(x[64]), .B(y[64]), .Z(n156) );
  XNOR U603 ( .A(n157), .B(n156), .Z(n158) );
  XOR U604 ( .A(n159), .B(n158), .Z(n512) );
  XNOR U605 ( .A(x[56]), .B(y[56]), .Z(n165) );
  XNOR U606 ( .A(x[54]), .B(y[54]), .Z(n163) );
  XNOR U607 ( .A(x[52]), .B(y[52]), .Z(n162) );
  XNOR U608 ( .A(n163), .B(n162), .Z(n164) );
  XOR U609 ( .A(n165), .B(n164), .Z(n509) );
  XNOR U610 ( .A(x[62]), .B(y[62]), .Z(n153) );
  XNOR U611 ( .A(x[60]), .B(y[60]), .Z(n151) );
  XNOR U612 ( .A(x[58]), .B(y[58]), .Z(n150) );
  XNOR U613 ( .A(n151), .B(n150), .Z(n152) );
  XOR U614 ( .A(n153), .B(n152), .Z(n510) );
  XNOR U615 ( .A(n509), .B(n510), .Z(n511) );
  XOR U616 ( .A(n512), .B(n511), .Z(n456) );
  XOR U617 ( .A(n457), .B(n456), .Z(n459) );
  XOR U618 ( .A(n458), .B(n459), .Z(n413) );
  XNOR U619 ( .A(n412), .B(n413), .Z(n107) );
  XNOR U620 ( .A(n106), .B(n107), .Z(o[0]) );
  NAND U621 ( .A(n105), .B(n104), .Z(n109) );
  NAND U622 ( .A(n107), .B(n106), .Z(n108) );
  NAND U623 ( .A(n109), .B(n108), .Z(n741) );
  OR U624 ( .A(n111), .B(n110), .Z(n115) );
  OR U625 ( .A(n113), .B(n112), .Z(n114) );
  NAND U626 ( .A(n115), .B(n114), .Z(n583) );
  OR U627 ( .A(n117), .B(n116), .Z(n121) );
  OR U628 ( .A(n119), .B(n118), .Z(n120) );
  NAND U629 ( .A(n121), .B(n120), .Z(n582) );
  OR U630 ( .A(n123), .B(n122), .Z(n127) );
  OR U631 ( .A(n125), .B(n124), .Z(n126) );
  AND U632 ( .A(n127), .B(n126), .Z(n581) );
  XOR U633 ( .A(n582), .B(n581), .Z(n128) );
  XNOR U634 ( .A(n583), .B(n128), .Z(n607) );
  OR U635 ( .A(n130), .B(n129), .Z(n134) );
  OR U636 ( .A(n132), .B(n131), .Z(n133) );
  NAND U637 ( .A(n134), .B(n133), .Z(n655) );
  OR U638 ( .A(n136), .B(n135), .Z(n140) );
  OR U639 ( .A(n138), .B(n137), .Z(n139) );
  NAND U640 ( .A(n140), .B(n139), .Z(n654) );
  XNOR U641 ( .A(n655), .B(n654), .Z(n656) );
  OR U642 ( .A(n142), .B(n141), .Z(n146) );
  OR U643 ( .A(n144), .B(n143), .Z(n145) );
  NAND U644 ( .A(n146), .B(n145), .Z(n657) );
  XNOR U645 ( .A(n605), .B(n604), .Z(n606) );
  XNOR U646 ( .A(n607), .B(n606), .Z(n754) );
  OR U647 ( .A(n151), .B(n150), .Z(n155) );
  OR U648 ( .A(n153), .B(n152), .Z(n154) );
  NAND U649 ( .A(n155), .B(n154), .Z(n651) );
  OR U650 ( .A(n157), .B(n156), .Z(n161) );
  OR U651 ( .A(n159), .B(n158), .Z(n160) );
  NAND U652 ( .A(n161), .B(n160), .Z(n649) );
  OR U653 ( .A(n163), .B(n162), .Z(n167) );
  OR U654 ( .A(n165), .B(n164), .Z(n166) );
  NAND U655 ( .A(n167), .B(n166), .Z(n648) );
  XNOR U656 ( .A(n649), .B(n648), .Z(n650) );
  XNOR U657 ( .A(n651), .B(n650), .Z(n638) );
  OR U658 ( .A(n169), .B(n168), .Z(n173) );
  OR U659 ( .A(n171), .B(n170), .Z(n172) );
  AND U660 ( .A(n173), .B(n172), .Z(n645) );
  OR U661 ( .A(n175), .B(n174), .Z(n179) );
  OR U662 ( .A(n177), .B(n176), .Z(n178) );
  NAND U663 ( .A(n179), .B(n178), .Z(n647) );
  OR U664 ( .A(n181), .B(n180), .Z(n185) );
  OR U665 ( .A(n183), .B(n182), .Z(n184) );
  NAND U666 ( .A(n185), .B(n184), .Z(n646) );
  XNOR U667 ( .A(n647), .B(n646), .Z(n186) );
  XOR U668 ( .A(n645), .B(n186), .Z(n636) );
  OR U669 ( .A(n188), .B(n187), .Z(n192) );
  OR U670 ( .A(n190), .B(n189), .Z(n191) );
  AND U671 ( .A(n192), .B(n191), .Z(n714) );
  OR U672 ( .A(n194), .B(n193), .Z(n198) );
  OR U673 ( .A(n196), .B(n195), .Z(n197) );
  AND U674 ( .A(n198), .B(n197), .Z(n710) );
  IV U675 ( .A(n710), .Z(n712) );
  OR U676 ( .A(n200), .B(n199), .Z(n702) );
  OR U677 ( .A(n202), .B(n201), .Z(n206) );
  OR U678 ( .A(n204), .B(n203), .Z(n205) );
  AND U679 ( .A(n206), .B(n205), .Z(n703) );
  XOR U680 ( .A(n702), .B(n703), .Z(n711) );
  XOR U681 ( .A(n712), .B(n711), .Z(n207) );
  XNOR U682 ( .A(n714), .B(n207), .Z(n635) );
  XOR U683 ( .A(n636), .B(n635), .Z(n637) );
  XNOR U684 ( .A(n638), .B(n637), .Z(n752) );
  OR U685 ( .A(n212), .B(n211), .Z(n216) );
  NANDN U686 ( .A(n214), .B(n213), .Z(n215) );
  AND U687 ( .A(n216), .B(n215), .Z(n673) );
  OR U688 ( .A(n218), .B(n217), .Z(n222) );
  NANDN U689 ( .A(n220), .B(n219), .Z(n221) );
  AND U690 ( .A(n222), .B(n221), .Z(n670) );
  OR U691 ( .A(n224), .B(n223), .Z(n228) );
  OR U692 ( .A(n226), .B(n225), .Z(n227) );
  AND U693 ( .A(n228), .B(n227), .Z(n671) );
  XNOR U694 ( .A(n670), .B(n671), .Z(n672) );
  OR U695 ( .A(n230), .B(n229), .Z(n234) );
  OR U696 ( .A(n232), .B(n231), .Z(n233) );
  NAND U697 ( .A(n234), .B(n233), .Z(n685) );
  OR U698 ( .A(n236), .B(n235), .Z(n240) );
  OR U699 ( .A(n238), .B(n237), .Z(n239) );
  NAND U700 ( .A(n240), .B(n239), .Z(n683) );
  OR U701 ( .A(n242), .B(n241), .Z(n246) );
  OR U702 ( .A(n244), .B(n243), .Z(n245) );
  NAND U703 ( .A(n246), .B(n245), .Z(n682) );
  XNOR U704 ( .A(n683), .B(n682), .Z(n684) );
  XNOR U705 ( .A(n685), .B(n684), .Z(n736) );
  XNOR U706 ( .A(n734), .B(n733), .Z(n735) );
  XNOR U707 ( .A(n736), .B(n735), .Z(n574) );
  XOR U708 ( .A(n574), .B(n575), .Z(n258) );
  XNOR U709 ( .A(n576), .B(n258), .Z(n588) );
  NAND U710 ( .A(n260), .B(n259), .Z(n264) );
  NAND U711 ( .A(n262), .B(n261), .Z(n263) );
  NAND U712 ( .A(n264), .B(n263), .Z(n590) );
  OR U713 ( .A(n267), .B(n265), .Z(n271) );
  ANDN U714 ( .B(n267), .A(n266), .Z(n268) );
  OR U715 ( .A(n269), .B(n268), .Z(n270) );
  NAND U716 ( .A(n271), .B(n270), .Z(n629) );
  NANDN U717 ( .A(n273), .B(n272), .Z(n277) );
  NANDN U718 ( .A(n275), .B(n274), .Z(n276) );
  AND U719 ( .A(n277), .B(n276), .Z(n630) );
  XOR U720 ( .A(n629), .B(n630), .Z(n632) );
  OR U721 ( .A(n279), .B(n278), .Z(n283) );
  OR U722 ( .A(n281), .B(n280), .Z(n282) );
  NAND U723 ( .A(n283), .B(n282), .Z(n669) );
  OR U724 ( .A(n285), .B(n284), .Z(n289) );
  OR U725 ( .A(n287), .B(n286), .Z(n288) );
  NAND U726 ( .A(n289), .B(n288), .Z(n667) );
  OR U727 ( .A(n291), .B(n290), .Z(n295) );
  OR U728 ( .A(n293), .B(n292), .Z(n294) );
  AND U729 ( .A(n295), .B(n294), .Z(n668) );
  XOR U730 ( .A(n667), .B(n668), .Z(n296) );
  XOR U731 ( .A(n669), .B(n296), .Z(n631) );
  XNOR U732 ( .A(n632), .B(n631), .Z(n589) );
  XOR U733 ( .A(n590), .B(n589), .Z(n297) );
  XOR U734 ( .A(n588), .B(n297), .Z(n770) );
  OR U735 ( .A(n299), .B(n298), .Z(n303) );
  NANDN U736 ( .A(n301), .B(n300), .Z(n302) );
  AND U737 ( .A(n303), .B(n302), .Z(n769) );
  XOR U738 ( .A(n770), .B(n769), .Z(n304) );
  XOR U739 ( .A(n771), .B(n304), .Z(n740) );
  XNOR U740 ( .A(n741), .B(n740), .Z(n742) );
  OR U741 ( .A(n306), .B(n305), .Z(n310) );
  OR U742 ( .A(n308), .B(n307), .Z(n309) );
  NAND U743 ( .A(n310), .B(n309), .Z(n615) );
  NAND U744 ( .A(n312), .B(n311), .Z(n316) );
  NAND U745 ( .A(n314), .B(n313), .Z(n315) );
  AND U746 ( .A(n316), .B(n315), .Z(n613) );
  XNOR U747 ( .A(n613), .B(n614), .Z(n320) );
  XOR U748 ( .A(n615), .B(n320), .Z(n748) );
  OR U749 ( .A(n322), .B(n321), .Z(n326) );
  NANDN U750 ( .A(n324), .B(n323), .Z(n325) );
  NAND U751 ( .A(n326), .B(n325), .Z(n578) );
  OR U752 ( .A(n328), .B(n327), .Z(n332) );
  NANDN U753 ( .A(n330), .B(n329), .Z(n331) );
  AND U754 ( .A(n332), .B(n331), .Z(n577) );
  XNOR U755 ( .A(n578), .B(n577), .Z(n579) );
  OR U756 ( .A(n334), .B(n333), .Z(n338) );
  NANDN U757 ( .A(n336), .B(n335), .Z(n337) );
  NAND U758 ( .A(n338), .B(n337), .Z(n580) );
  XOR U759 ( .A(n579), .B(n580), .Z(n610) );
  OR U760 ( .A(n341), .B(n339), .Z(n345) );
  ANDN U761 ( .B(n341), .A(n340), .Z(n343) );
  NANDN U762 ( .A(n343), .B(n342), .Z(n344) );
  NAND U763 ( .A(n345), .B(n344), .Z(n611) );
  OR U764 ( .A(n347), .B(n346), .Z(n351) );
  OR U765 ( .A(n349), .B(n348), .Z(n350) );
  AND U766 ( .A(n351), .B(n350), .Z(n689) );
  IV U767 ( .A(n689), .Z(n688) );
  OR U768 ( .A(n353), .B(n352), .Z(n357) );
  OR U769 ( .A(n355), .B(n354), .Z(n356) );
  NAND U770 ( .A(n357), .B(n356), .Z(n692) );
  OR U771 ( .A(n359), .B(n358), .Z(n363) );
  OR U772 ( .A(n361), .B(n360), .Z(n362) );
  NAND U773 ( .A(n363), .B(n362), .Z(n690) );
  XNOR U774 ( .A(n692), .B(n690), .Z(n364) );
  XNOR U775 ( .A(n688), .B(n364), .Z(n612) );
  XNOR U776 ( .A(n611), .B(n612), .Z(n365) );
  XNOR U777 ( .A(n610), .B(n365), .Z(n746) );
  NAND U778 ( .A(n367), .B(n366), .Z(n371) );
  NAND U779 ( .A(n369), .B(n368), .Z(n370) );
  AND U780 ( .A(n371), .B(n370), .Z(n718) );
  NANDN U781 ( .A(n373), .B(n372), .Z(n377) );
  NAND U782 ( .A(n375), .B(n374), .Z(n376) );
  NAND U783 ( .A(n377), .B(n376), .Z(n719) );
  OR U784 ( .A(n379), .B(n378), .Z(n383) );
  NANDN U785 ( .A(n381), .B(n380), .Z(n382) );
  NAND U786 ( .A(n383), .B(n382), .Z(n586) );
  OR U787 ( .A(n385), .B(n384), .Z(n389) );
  OR U788 ( .A(n387), .B(n386), .Z(n388) );
  NAND U789 ( .A(n389), .B(n388), .Z(n585) );
  OR U790 ( .A(n391), .B(n390), .Z(n395) );
  OR U791 ( .A(n393), .B(n392), .Z(n394) );
  AND U792 ( .A(n395), .B(n394), .Z(n584) );
  XOR U793 ( .A(n585), .B(n584), .Z(n396) );
  XOR U794 ( .A(n586), .B(n396), .Z(n717) );
  XOR U795 ( .A(n719), .B(n717), .Z(n397) );
  XNOR U796 ( .A(n718), .B(n397), .Z(n570) );
  OR U797 ( .A(n399), .B(n398), .Z(n403) );
  OR U798 ( .A(n401), .B(n400), .Z(n402) );
  NAND U799 ( .A(n403), .B(n402), .Z(n569) );
  XOR U800 ( .A(n569), .B(n568), .Z(n571) );
  XNOR U801 ( .A(n570), .B(n571), .Z(n747) );
  XOR U802 ( .A(n746), .B(n747), .Z(n749) );
  XNOR U803 ( .A(n748), .B(n749), .Z(n766) );
  NAND U804 ( .A(n411), .B(n410), .Z(n415) );
  NANDN U805 ( .A(n413), .B(n412), .Z(n414) );
  NAND U806 ( .A(n415), .B(n414), .Z(n593) );
  OR U807 ( .A(n417), .B(n416), .Z(n421) );
  OR U808 ( .A(n419), .B(n418), .Z(n420) );
  NAND U809 ( .A(n421), .B(n420), .Z(n677) );
  OR U810 ( .A(n423), .B(n422), .Z(n427) );
  OR U811 ( .A(n425), .B(n424), .Z(n426) );
  NAND U812 ( .A(n427), .B(n426), .Z(n676) );
  XNOR U813 ( .A(n677), .B(n676), .Z(n678) );
  OR U814 ( .A(n429), .B(n428), .Z(n433) );
  NANDN U815 ( .A(n431), .B(n430), .Z(n432) );
  NAND U816 ( .A(n433), .B(n432), .Z(n679) );
  OR U817 ( .A(n435), .B(n434), .Z(n439) );
  OR U818 ( .A(n437), .B(n436), .Z(n438) );
  AND U819 ( .A(n439), .B(n438), .Z(n664) );
  OR U820 ( .A(n441), .B(n440), .Z(n445) );
  OR U821 ( .A(n443), .B(n442), .Z(n444) );
  AND U822 ( .A(n445), .B(n444), .Z(n661) );
  OR U823 ( .A(n447), .B(n446), .Z(n451) );
  OR U824 ( .A(n449), .B(n448), .Z(n450) );
  AND U825 ( .A(n451), .B(n450), .Z(n662) );
  XNOR U826 ( .A(n661), .B(n662), .Z(n663) );
  XOR U827 ( .A(n616), .B(n617), .Z(n619) );
  XOR U828 ( .A(n618), .B(n619), .Z(n592) );
  XOR U829 ( .A(n593), .B(n592), .Z(n455) );
  XOR U830 ( .A(n591), .B(n455), .Z(n763) );
  NANDN U831 ( .A(n457), .B(n456), .Z(n461) );
  NANDN U832 ( .A(n459), .B(n458), .Z(n460) );
  AND U833 ( .A(n461), .B(n460), .Z(n595) );
  OR U834 ( .A(n463), .B(n462), .Z(n467) );
  NANDN U835 ( .A(n465), .B(n464), .Z(n466) );
  AND U836 ( .A(n467), .B(n466), .Z(n707) );
  OR U837 ( .A(n469), .B(n468), .Z(n473) );
  NANDN U838 ( .A(n471), .B(n470), .Z(n472) );
  AND U839 ( .A(n473), .B(n472), .Z(n704) );
  OR U840 ( .A(n475), .B(n474), .Z(n479) );
  NANDN U841 ( .A(n477), .B(n476), .Z(n478) );
  AND U842 ( .A(n479), .B(n478), .Z(n705) );
  XNOR U843 ( .A(n704), .B(n705), .Z(n706) );
  OR U844 ( .A(n481), .B(n480), .Z(n485) );
  OR U845 ( .A(n483), .B(n482), .Z(n484) );
  AND U846 ( .A(n485), .B(n484), .Z(n727) );
  IV U847 ( .A(n727), .Z(n726) );
  OR U848 ( .A(n487), .B(n486), .Z(n491) );
  NANDN U849 ( .A(n489), .B(n488), .Z(n490) );
  NAND U850 ( .A(n491), .B(n490), .Z(n730) );
  OR U851 ( .A(n493), .B(n492), .Z(n497) );
  OR U852 ( .A(n495), .B(n494), .Z(n496) );
  NAND U853 ( .A(n497), .B(n496), .Z(n728) );
  XNOR U854 ( .A(n730), .B(n728), .Z(n498) );
  XOR U855 ( .A(n726), .B(n498), .Z(n642) );
  IV U856 ( .A(n755), .Z(n757) );
  OR U857 ( .A(n504), .B(n502), .Z(n508) );
  ANDN U858 ( .B(n504), .A(n503), .Z(n505) );
  OR U859 ( .A(n506), .B(n505), .Z(n507) );
  NAND U860 ( .A(n508), .B(n507), .Z(n622) );
  OR U861 ( .A(n510), .B(n509), .Z(n514) );
  OR U862 ( .A(n512), .B(n511), .Z(n513) );
  AND U863 ( .A(n514), .B(n513), .Z(n623) );
  XOR U864 ( .A(n622), .B(n623), .Z(n625) );
  OR U865 ( .A(n516), .B(n515), .Z(n520) );
  NANDN U866 ( .A(n518), .B(n517), .Z(n519) );
  NAND U867 ( .A(n520), .B(n519), .Z(n721) );
  OR U868 ( .A(n522), .B(n521), .Z(n526) );
  NANDN U869 ( .A(n524), .B(n523), .Z(n525) );
  NAND U870 ( .A(n526), .B(n525), .Z(n720) );
  XNOR U871 ( .A(n721), .B(n720), .Z(n722) );
  OR U872 ( .A(n528), .B(n527), .Z(n532) );
  OR U873 ( .A(n530), .B(n529), .Z(n531) );
  NAND U874 ( .A(n532), .B(n531), .Z(n723) );
  OR U875 ( .A(n534), .B(n533), .Z(n538) );
  OR U876 ( .A(n536), .B(n535), .Z(n537) );
  AND U877 ( .A(n538), .B(n537), .Z(n598) );
  XOR U878 ( .A(n598), .B(n599), .Z(n600) );
  OR U879 ( .A(n543), .B(n542), .Z(n547) );
  NANDN U880 ( .A(n545), .B(n544), .Z(n546) );
  NAND U881 ( .A(n547), .B(n546), .Z(n697) );
  OR U882 ( .A(n549), .B(n548), .Z(n553) );
  OR U883 ( .A(n551), .B(n550), .Z(n552) );
  NAND U884 ( .A(n553), .B(n552), .Z(n696) );
  XNOR U885 ( .A(n697), .B(n696), .Z(n698) );
  OR U886 ( .A(n555), .B(n554), .Z(n559) );
  OR U887 ( .A(n557), .B(n556), .Z(n558) );
  NAND U888 ( .A(n559), .B(n558), .Z(n699) );
  XOR U889 ( .A(n600), .B(n601), .Z(n758) );
  XOR U890 ( .A(n756), .B(n758), .Z(n560) );
  XNOR U891 ( .A(n757), .B(n560), .Z(n597) );
  NANDN U892 ( .A(n561), .B(n562), .Z(n566) );
  NANDN U893 ( .A(n562), .B(n561), .Z(n564) );
  NAND U894 ( .A(n564), .B(n563), .Z(n565) );
  NAND U895 ( .A(n566), .B(n565), .Z(n596) );
  XOR U896 ( .A(n597), .B(n596), .Z(n567) );
  XOR U897 ( .A(n595), .B(n567), .Z(n764) );
  XOR U898 ( .A(n766), .B(n765), .Z(n743) );
  XNOR U899 ( .A(n742), .B(n743), .Z(o[1]) );
  NAND U900 ( .A(n569), .B(n568), .Z(n573) );
  NAND U901 ( .A(n571), .B(n570), .Z(n572) );
  NAND U902 ( .A(n573), .B(n572), .Z(n811) );
  IV U903 ( .A(n809), .Z(n808) );
  XNOR U904 ( .A(n836), .B(n837), .Z(n839) );
  XOR U905 ( .A(n838), .B(n839), .Z(n810) );
  XOR U906 ( .A(n808), .B(n810), .Z(n587) );
  XOR U907 ( .A(n811), .B(n587), .Z(n785) );
  IV U908 ( .A(n784), .Z(n786) );
  XNOR U909 ( .A(n787), .B(n786), .Z(n594) );
  XNOR U910 ( .A(n785), .B(n594), .Z(n888) );
  OR U911 ( .A(n599), .B(n598), .Z(n603) );
  NANDN U912 ( .A(n601), .B(n600), .Z(n602) );
  AND U913 ( .A(n603), .B(n602), .Z(n805) );
  NANDN U914 ( .A(n605), .B(n604), .Z(n609) );
  NANDN U915 ( .A(n607), .B(n606), .Z(n608) );
  AND U916 ( .A(n609), .B(n608), .Z(n803) );
  XNOR U917 ( .A(n803), .B(n802), .Z(n804) );
  XOR U918 ( .A(n805), .B(n804), .Z(n800) );
  IV U919 ( .A(n843), .Z(n844) );
  NANDN U920 ( .A(n617), .B(n616), .Z(n621) );
  OR U921 ( .A(n619), .B(n618), .Z(n620) );
  AND U922 ( .A(n621), .B(n620), .Z(n847) );
  NANDN U923 ( .A(n623), .B(n622), .Z(n627) );
  OR U924 ( .A(n625), .B(n624), .Z(n626) );
  AND U925 ( .A(n627), .B(n626), .Z(n845) );
  XNOR U926 ( .A(n847), .B(n845), .Z(n628) );
  XOR U927 ( .A(n844), .B(n628), .Z(n801) );
  NANDN U928 ( .A(n630), .B(n629), .Z(n634) );
  NANDN U929 ( .A(n632), .B(n631), .Z(n633) );
  NAND U930 ( .A(n634), .B(n633), .Z(n816) );
  OR U931 ( .A(n636), .B(n635), .Z(n640) );
  NANDN U932 ( .A(n638), .B(n637), .Z(n639) );
  NAND U933 ( .A(n640), .B(n639), .Z(n818) );
  IV U934 ( .A(n817), .Z(n815) );
  XNOR U935 ( .A(n818), .B(n815), .Z(n644) );
  XNOR U936 ( .A(n816), .B(n644), .Z(n779) );
  IV U937 ( .A(n875), .Z(n872) );
  OR U938 ( .A(n649), .B(n648), .Z(n653) );
  OR U939 ( .A(n651), .B(n650), .Z(n652) );
  NAND U940 ( .A(n653), .B(n652), .Z(n876) );
  OR U941 ( .A(n655), .B(n654), .Z(n659) );
  OR U942 ( .A(n657), .B(n656), .Z(n658) );
  AND U943 ( .A(n659), .B(n658), .Z(n873) );
  IV U944 ( .A(n873), .Z(n874) );
  XNOR U945 ( .A(n876), .B(n874), .Z(n660) );
  XOR U946 ( .A(n872), .B(n660), .Z(n853) );
  OR U947 ( .A(n662), .B(n661), .Z(n666) );
  OR U948 ( .A(n664), .B(n663), .Z(n665) );
  AND U949 ( .A(n666), .B(n665), .Z(n824) );
  OR U950 ( .A(n671), .B(n670), .Z(n675) );
  OR U951 ( .A(n673), .B(n672), .Z(n674) );
  AND U952 ( .A(n675), .B(n674), .Z(n823) );
  XOR U953 ( .A(n822), .B(n823), .Z(n825) );
  OR U954 ( .A(n677), .B(n676), .Z(n681) );
  OR U955 ( .A(n679), .B(n678), .Z(n680) );
  AND U956 ( .A(n681), .B(n680), .Z(n869) );
  OR U957 ( .A(n683), .B(n682), .Z(n687) );
  OR U958 ( .A(n685), .B(n684), .Z(n686) );
  AND U959 ( .A(n687), .B(n686), .Z(n867) );
  OR U960 ( .A(n690), .B(n688), .Z(n694) );
  ANDN U961 ( .B(n690), .A(n689), .Z(n691) );
  OR U962 ( .A(n692), .B(n691), .Z(n693) );
  NAND U963 ( .A(n694), .B(n693), .Z(n866) );
  XNOR U964 ( .A(n867), .B(n866), .Z(n868) );
  XNOR U965 ( .A(n869), .B(n868), .Z(n852) );
  XOR U966 ( .A(n851), .B(n852), .Z(n695) );
  XNOR U967 ( .A(n853), .B(n695), .Z(n778) );
  XOR U968 ( .A(n779), .B(n778), .Z(n781) );
  OR U969 ( .A(n697), .B(n696), .Z(n701) );
  OR U970 ( .A(n699), .B(n698), .Z(n700) );
  NAND U971 ( .A(n701), .B(n700), .Z(n833) );
  OR U972 ( .A(n703), .B(n702), .Z(n829) );
  OR U973 ( .A(n705), .B(n704), .Z(n709) );
  OR U974 ( .A(n707), .B(n706), .Z(n708) );
  AND U975 ( .A(n709), .B(n708), .Z(n828) );
  XOR U976 ( .A(n829), .B(n828), .Z(n830) );
  NANDN U977 ( .A(n710), .B(n711), .Z(n716) );
  NOR U978 ( .A(n712), .B(n711), .Z(n713) );
  OR U979 ( .A(n714), .B(n713), .Z(n715) );
  NAND U980 ( .A(n716), .B(n715), .Z(n831) );
  XNOR U981 ( .A(n833), .B(n832), .Z(n855) );
  XOR U982 ( .A(n855), .B(n854), .Z(n857) );
  OR U983 ( .A(n721), .B(n720), .Z(n725) );
  OR U984 ( .A(n723), .B(n722), .Z(n724) );
  AND U985 ( .A(n725), .B(n724), .Z(n862) );
  OR U986 ( .A(n728), .B(n726), .Z(n732) );
  ANDN U987 ( .B(n728), .A(n727), .Z(n729) );
  OR U988 ( .A(n730), .B(n729), .Z(n731) );
  NAND U989 ( .A(n732), .B(n731), .Z(n860) );
  OR U990 ( .A(n734), .B(n733), .Z(n738) );
  OR U991 ( .A(n736), .B(n735), .Z(n737) );
  AND U992 ( .A(n738), .B(n737), .Z(n861) );
  XOR U993 ( .A(n860), .B(n861), .Z(n863) );
  XOR U994 ( .A(n862), .B(n863), .Z(n856) );
  XOR U995 ( .A(n857), .B(n856), .Z(n780) );
  XNOR U996 ( .A(n886), .B(n887), .Z(n739) );
  XOR U997 ( .A(n888), .B(n739), .Z(n772) );
  NAND U998 ( .A(n741), .B(n740), .Z(n745) );
  OR U999 ( .A(n743), .B(n742), .Z(n744) );
  AND U1000 ( .A(n745), .B(n744), .Z(n773) );
  XNOR U1001 ( .A(n772), .B(n773), .Z(n774) );
  NANDN U1002 ( .A(n747), .B(n746), .Z(n751) );
  OR U1003 ( .A(n749), .B(n748), .Z(n750) );
  AND U1004 ( .A(n751), .B(n750), .Z(n793) );
  NANDN U1005 ( .A(n755), .B(n756), .Z(n761) );
  NOR U1006 ( .A(n757), .B(n756), .Z(n759) );
  OR U1007 ( .A(n759), .B(n758), .Z(n760) );
  AND U1008 ( .A(n761), .B(n760), .Z(n791) );
  IV U1009 ( .A(n791), .Z(n792) );
  XNOR U1010 ( .A(n794), .B(n792), .Z(n762) );
  XOR U1011 ( .A(n793), .B(n762), .Z(n882) );
  NANDN U1012 ( .A(n764), .B(n763), .Z(n768) );
  NANDN U1013 ( .A(n766), .B(n765), .Z(n767) );
  AND U1014 ( .A(n768), .B(n767), .Z(n880) );
  XNOR U1015 ( .A(n774), .B(n775), .Z(o[2]) );
  NANDN U1016 ( .A(n773), .B(n772), .Z(n777) );
  NAND U1017 ( .A(n775), .B(n774), .Z(n776) );
  NAND U1018 ( .A(n777), .B(n776), .Z(n945) );
  NANDN U1019 ( .A(n779), .B(n778), .Z(n783) );
  OR U1020 ( .A(n781), .B(n780), .Z(n782) );
  AND U1021 ( .A(n783), .B(n782), .Z(n898) );
  NANDN U1022 ( .A(n784), .B(n785), .Z(n790) );
  NOR U1023 ( .A(n786), .B(n785), .Z(n788) );
  NANDN U1024 ( .A(n788), .B(n787), .Z(n789) );
  NAND U1025 ( .A(n790), .B(n789), .Z(n899) );
  OR U1026 ( .A(n793), .B(n791), .Z(n797) );
  ANDN U1027 ( .B(n793), .A(n792), .Z(n795) );
  NANDN U1028 ( .A(n795), .B(n794), .Z(n796) );
  AND U1029 ( .A(n797), .B(n796), .Z(n896) );
  IV U1030 ( .A(n896), .Z(n897) );
  XNOR U1031 ( .A(n899), .B(n897), .Z(n798) );
  XNOR U1032 ( .A(n898), .B(n798), .Z(n946) );
  XNOR U1033 ( .A(n945), .B(n946), .Z(n947) );
  NANDN U1034 ( .A(n803), .B(n802), .Z(n807) );
  NANDN U1035 ( .A(n805), .B(n804), .Z(n806) );
  AND U1036 ( .A(n807), .B(n806), .Z(n911) );
  OR U1037 ( .A(n810), .B(n808), .Z(n814) );
  ANDN U1038 ( .B(n810), .A(n809), .Z(n812) );
  NANDN U1039 ( .A(n812), .B(n811), .Z(n813) );
  NAND U1040 ( .A(n814), .B(n813), .Z(n926) );
  NANDN U1041 ( .A(n815), .B(n816), .Z(n821) );
  NOR U1042 ( .A(n817), .B(n816), .Z(n819) );
  NANDN U1043 ( .A(n819), .B(n818), .Z(n820) );
  NAND U1044 ( .A(n821), .B(n820), .Z(n928) );
  NANDN U1045 ( .A(n823), .B(n822), .Z(n827) );
  OR U1046 ( .A(n825), .B(n824), .Z(n826) );
  AND U1047 ( .A(n827), .B(n826), .Z(n916) );
  OR U1048 ( .A(n829), .B(n828), .Z(n917) );
  XNOR U1049 ( .A(n916), .B(n917), .Z(n921) );
  OR U1050 ( .A(n831), .B(n830), .Z(n835) );
  NAND U1051 ( .A(n833), .B(n832), .Z(n834) );
  NAND U1052 ( .A(n835), .B(n834), .Z(n920) );
  NAND U1053 ( .A(n837), .B(n836), .Z(n841) );
  NANDN U1054 ( .A(n839), .B(n838), .Z(n840) );
  NAND U1055 ( .A(n841), .B(n840), .Z(n918) );
  XNOR U1056 ( .A(n919), .B(n918), .Z(n927) );
  IV U1057 ( .A(n927), .Z(n925) );
  XOR U1058 ( .A(n928), .B(n925), .Z(n842) );
  XOR U1059 ( .A(n926), .B(n842), .Z(n913) );
  OR U1060 ( .A(n845), .B(n843), .Z(n849) );
  ANDN U1061 ( .B(n845), .A(n844), .Z(n846) );
  OR U1062 ( .A(n847), .B(n846), .Z(n848) );
  AND U1063 ( .A(n849), .B(n848), .Z(n909) );
  IV U1064 ( .A(n909), .Z(n910) );
  XOR U1065 ( .A(n913), .B(n910), .Z(n850) );
  XNOR U1066 ( .A(n911), .B(n850), .Z(n891) );
  XOR U1067 ( .A(n890), .B(n891), .Z(n893) );
  NANDN U1068 ( .A(n855), .B(n854), .Z(n859) );
  NANDN U1069 ( .A(n857), .B(n856), .Z(n858) );
  AND U1070 ( .A(n859), .B(n858), .Z(n904) );
  XOR U1071 ( .A(n903), .B(n904), .Z(n906) );
  NANDN U1072 ( .A(n861), .B(n860), .Z(n865) );
  OR U1073 ( .A(n863), .B(n862), .Z(n864) );
  AND U1074 ( .A(n865), .B(n864), .Z(n934) );
  NANDN U1075 ( .A(n867), .B(n866), .Z(n871) );
  NANDN U1076 ( .A(n869), .B(n868), .Z(n870) );
  AND U1077 ( .A(n871), .B(n870), .Z(n933) );
  NANDN U1078 ( .A(n873), .B(n872), .Z(n879) );
  ANDN U1079 ( .B(n875), .A(n874), .Z(n877) );
  NANDN U1080 ( .A(n877), .B(n876), .Z(n878) );
  NAND U1081 ( .A(n879), .B(n878), .Z(n932) );
  XOR U1082 ( .A(n933), .B(n932), .Z(n935) );
  XNOR U1083 ( .A(n934), .B(n935), .Z(n905) );
  XNOR U1084 ( .A(n906), .B(n905), .Z(n892) );
  XOR U1085 ( .A(n893), .B(n892), .Z(n939) );
  OR U1086 ( .A(n881), .B(n880), .Z(n885) );
  NANDN U1087 ( .A(n883), .B(n882), .Z(n884) );
  NAND U1088 ( .A(n885), .B(n884), .Z(n941) );
  IV U1089 ( .A(n940), .Z(n938) );
  XNOR U1090 ( .A(n941), .B(n938), .Z(n889) );
  XNOR U1091 ( .A(n939), .B(n889), .Z(n948) );
  XOR U1092 ( .A(n947), .B(n948), .Z(o[3]) );
  NANDN U1093 ( .A(n891), .B(n890), .Z(n895) );
  OR U1094 ( .A(n893), .B(n892), .Z(n894) );
  AND U1095 ( .A(n895), .B(n894), .Z(n958) );
  OR U1096 ( .A(n898), .B(n896), .Z(n902) );
  ANDN U1097 ( .B(n898), .A(n897), .Z(n900) );
  NANDN U1098 ( .A(n900), .B(n899), .Z(n901) );
  NAND U1099 ( .A(n902), .B(n901), .Z(n955) );
  NANDN U1100 ( .A(n904), .B(n903), .Z(n908) );
  OR U1101 ( .A(n906), .B(n905), .Z(n907) );
  AND U1102 ( .A(n908), .B(n907), .Z(n972) );
  OR U1103 ( .A(n911), .B(n909), .Z(n915) );
  ANDN U1104 ( .B(n911), .A(n910), .Z(n912) );
  OR U1105 ( .A(n913), .B(n912), .Z(n914) );
  AND U1106 ( .A(n915), .B(n914), .Z(n970) );
  OR U1107 ( .A(n917), .B(n916), .Z(n968) );
  OR U1108 ( .A(n919), .B(n918), .Z(n967) );
  XNOR U1109 ( .A(n968), .B(n967), .Z(n924) );
  NOR U1110 ( .A(n921), .B(n920), .Z(n922) );
  NAND U1111 ( .A(n922), .B(n968), .Z(n923) );
  AND U1112 ( .A(n924), .B(n923), .Z(n964) );
  NANDN U1113 ( .A(n925), .B(n926), .Z(n931) );
  NOR U1114 ( .A(n927), .B(n926), .Z(n929) );
  NANDN U1115 ( .A(n929), .B(n928), .Z(n930) );
  NAND U1116 ( .A(n931), .B(n930), .Z(n962) );
  NANDN U1117 ( .A(n933), .B(n932), .Z(n937) );
  OR U1118 ( .A(n935), .B(n934), .Z(n936) );
  NAND U1119 ( .A(n937), .B(n936), .Z(n961) );
  XNOR U1120 ( .A(n962), .B(n961), .Z(n963) );
  XNOR U1121 ( .A(n964), .B(n963), .Z(n969) );
  XNOR U1122 ( .A(n970), .B(n969), .Z(n971) );
  XNOR U1123 ( .A(n972), .B(n971), .Z(n956) );
  XOR U1124 ( .A(n955), .B(n956), .Z(n957) );
  XOR U1125 ( .A(n958), .B(n957), .Z(n954) );
  NANDN U1126 ( .A(n938), .B(n939), .Z(n944) );
  NOR U1127 ( .A(n940), .B(n939), .Z(n942) );
  NANDN U1128 ( .A(n942), .B(n941), .Z(n943) );
  NAND U1129 ( .A(n944), .B(n943), .Z(n952) );
  NANDN U1130 ( .A(n946), .B(n945), .Z(n950) );
  NANDN U1131 ( .A(n948), .B(n947), .Z(n949) );
  AND U1132 ( .A(n950), .B(n949), .Z(n953) );
  XOR U1133 ( .A(n952), .B(n953), .Z(n951) );
  XNOR U1134 ( .A(n954), .B(n951), .Z(o[4]) );
  NAND U1135 ( .A(n956), .B(n955), .Z(n960) );
  NANDN U1136 ( .A(n958), .B(n957), .Z(n959) );
  AND U1137 ( .A(n960), .B(n959), .Z(n976) );
  XNOR U1138 ( .A(n975), .B(n976), .Z(n977) );
  OR U1139 ( .A(n962), .B(n961), .Z(n966) );
  OR U1140 ( .A(n964), .B(n963), .Z(n965) );
  AND U1141 ( .A(n966), .B(n965), .Z(n984) );
  OR U1142 ( .A(n968), .B(n967), .Z(n982) );
  NANDN U1143 ( .A(n970), .B(n969), .Z(n974) );
  NANDN U1144 ( .A(n972), .B(n971), .Z(n973) );
  NAND U1145 ( .A(n974), .B(n973), .Z(n981) );
  XOR U1146 ( .A(n982), .B(n981), .Z(n983) );
  XNOR U1147 ( .A(n984), .B(n983), .Z(n978) );
  XOR U1148 ( .A(n977), .B(n978), .Z(o[5]) );
  NANDN U1149 ( .A(n976), .B(n975), .Z(n980) );
  NANDN U1150 ( .A(n978), .B(n977), .Z(n979) );
  NAND U1151 ( .A(n980), .B(n979), .Z(n988) );
  OR U1152 ( .A(n982), .B(n981), .Z(n986) );
  NANDN U1153 ( .A(n984), .B(n983), .Z(n985) );
  AND U1154 ( .A(n986), .B(n985), .Z(n987) );
  XOR U1155 ( .A(n988), .B(n987), .Z(o[6]) );
  NOR U1156 ( .A(n988), .B(n987), .Z(o[7]) );
endmodule

