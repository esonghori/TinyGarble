
module sum ( a, b, c );
  input [255:0] a;
  input [255:0] b;
  output [256:0] c;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270;

  IV U2 ( .A(n2157), .Z(n2) );
  IV U3 ( .A(b[4]), .Z(n3) );
  NOR U4 ( .A(n2), .B(n3), .Z(n4) );
  XOR U5 ( .A(n2157), .B(n3), .Z(n5) );
  IV U6 ( .A(a[4]), .Z(n6) );
  NOR U7 ( .A(n5), .B(n6), .Z(n7) );
  NOR U8 ( .A(n4), .B(n7), .Z(n8) );
  IV U9 ( .A(n8), .Z(n2179) );
  IV U10 ( .A(n2223), .Z(n9) );
  IV U11 ( .A(b[7]), .Z(n10) );
  NOR U12 ( .A(n9), .B(n10), .Z(n11) );
  XOR U13 ( .A(n2223), .B(n10), .Z(n12) );
  IV U14 ( .A(a[7]), .Z(n13) );
  NOR U15 ( .A(n12), .B(n13), .Z(n14) );
  NOR U16 ( .A(n11), .B(n14), .Z(n15) );
  IV U17 ( .A(n15), .Z(n2245) );
  IV U18 ( .A(n1744), .Z(n16) );
  IV U19 ( .A(b[10]), .Z(n17) );
  NOR U20 ( .A(n16), .B(n17), .Z(n18) );
  XOR U21 ( .A(n1744), .B(n17), .Z(n19) );
  IV U22 ( .A(a[10]), .Z(n20) );
  NOR U23 ( .A(n19), .B(n20), .Z(n21) );
  NOR U24 ( .A(n18), .B(n21), .Z(n22) );
  IV U25 ( .A(n22), .Z(n1766) );
  IV U26 ( .A(n1810), .Z(n23) );
  IV U27 ( .A(b[13]), .Z(n24) );
  NOR U28 ( .A(n23), .B(n24), .Z(n25) );
  XOR U29 ( .A(n1810), .B(n24), .Z(n26) );
  IV U30 ( .A(a[13]), .Z(n27) );
  NOR U31 ( .A(n26), .B(n27), .Z(n28) );
  NOR U32 ( .A(n25), .B(n28), .Z(n29) );
  IV U33 ( .A(n29), .Z(n1832) );
  IV U34 ( .A(n1876), .Z(n30) );
  IV U35 ( .A(b[16]), .Z(n31) );
  NOR U36 ( .A(n30), .B(n31), .Z(n32) );
  XOR U37 ( .A(n1876), .B(n31), .Z(n33) );
  IV U38 ( .A(a[16]), .Z(n34) );
  NOR U39 ( .A(n33), .B(n34), .Z(n35) );
  NOR U40 ( .A(n32), .B(n35), .Z(n36) );
  IV U41 ( .A(n36), .Z(n1898) );
  IV U42 ( .A(n1942), .Z(n37) );
  IV U43 ( .A(b[19]), .Z(n38) );
  NOR U44 ( .A(n37), .B(n38), .Z(n39) );
  XOR U45 ( .A(n1942), .B(n38), .Z(n40) );
  IV U46 ( .A(a[19]), .Z(n41) );
  NOR U47 ( .A(n40), .B(n41), .Z(n42) );
  NOR U48 ( .A(n39), .B(n42), .Z(n43) );
  IV U49 ( .A(n43), .Z(n1966) );
  IV U50 ( .A(n2010), .Z(n44) );
  IV U51 ( .A(b[22]), .Z(n45) );
  NOR U52 ( .A(n44), .B(n45), .Z(n46) );
  XOR U53 ( .A(n2010), .B(n45), .Z(n47) );
  IV U54 ( .A(a[22]), .Z(n48) );
  NOR U55 ( .A(n47), .B(n48), .Z(n49) );
  NOR U56 ( .A(n46), .B(n49), .Z(n50) );
  IV U57 ( .A(n50), .Z(n2032) );
  IV U58 ( .A(n2102), .Z(n51) );
  IV U59 ( .A(b[25]), .Z(n52) );
  NOR U60 ( .A(n51), .B(n52), .Z(n53) );
  XOR U61 ( .A(n2102), .B(n52), .Z(n54) );
  IV U62 ( .A(a[25]), .Z(n55) );
  NOR U63 ( .A(n54), .B(n55), .Z(n56) );
  NOR U64 ( .A(n53), .B(n56), .Z(n57) );
  IV U65 ( .A(n57), .Z(n2104) );
  IV U66 ( .A(n2108), .Z(n58) );
  IV U67 ( .A(b[28]), .Z(n59) );
  NOR U68 ( .A(n58), .B(n59), .Z(n60) );
  XOR U69 ( .A(n2108), .B(n59), .Z(n61) );
  IV U70 ( .A(a[28]), .Z(n62) );
  NOR U71 ( .A(n61), .B(n62), .Z(n63) );
  NOR U72 ( .A(n60), .B(n63), .Z(n64) );
  IV U73 ( .A(n64), .Z(n2110) );
  IV U74 ( .A(n2117), .Z(n65) );
  IV U75 ( .A(b[31]), .Z(n66) );
  NOR U76 ( .A(n65), .B(n66), .Z(n67) );
  XOR U77 ( .A(n2117), .B(n66), .Z(n68) );
  IV U78 ( .A(a[31]), .Z(n69) );
  NOR U79 ( .A(n68), .B(n69), .Z(n70) );
  NOR U80 ( .A(n67), .B(n70), .Z(n71) );
  IV U81 ( .A(n71), .Z(n2119) );
  IV U82 ( .A(n2123), .Z(n72) );
  IV U83 ( .A(b[34]), .Z(n73) );
  NOR U84 ( .A(n72), .B(n73), .Z(n74) );
  XOR U85 ( .A(n2123), .B(n73), .Z(n75) );
  IV U86 ( .A(a[34]), .Z(n76) );
  NOR U87 ( .A(n75), .B(n76), .Z(n77) );
  NOR U88 ( .A(n74), .B(n77), .Z(n78) );
  IV U89 ( .A(n78), .Z(n2125) );
  IV U90 ( .A(n2129), .Z(n79) );
  IV U91 ( .A(b[37]), .Z(n80) );
  NOR U92 ( .A(n79), .B(n80), .Z(n81) );
  XOR U93 ( .A(n2129), .B(n80), .Z(n82) );
  IV U94 ( .A(a[37]), .Z(n83) );
  NOR U95 ( .A(n82), .B(n83), .Z(n84) );
  NOR U96 ( .A(n81), .B(n84), .Z(n85) );
  IV U97 ( .A(n85), .Z(n2131) );
  IV U98 ( .A(n2137), .Z(n86) );
  IV U99 ( .A(b[40]), .Z(n87) );
  NOR U100 ( .A(n86), .B(n87), .Z(n88) );
  XOR U101 ( .A(n2137), .B(n87), .Z(n89) );
  IV U102 ( .A(a[40]), .Z(n90) );
  NOR U103 ( .A(n89), .B(n90), .Z(n91) );
  NOR U104 ( .A(n88), .B(n91), .Z(n92) );
  IV U105 ( .A(n92), .Z(n2139) );
  IV U106 ( .A(n2143), .Z(n93) );
  IV U107 ( .A(b[43]), .Z(n94) );
  NOR U108 ( .A(n93), .B(n94), .Z(n95) );
  XOR U109 ( .A(n2143), .B(n94), .Z(n96) );
  IV U110 ( .A(a[43]), .Z(n97) );
  NOR U111 ( .A(n96), .B(n97), .Z(n98) );
  NOR U112 ( .A(n95), .B(n98), .Z(n99) );
  IV U113 ( .A(n99), .Z(n2145) );
  IV U114 ( .A(n2149), .Z(n100) );
  IV U115 ( .A(b[46]), .Z(n101) );
  NOR U116 ( .A(n100), .B(n101), .Z(n102) );
  XOR U117 ( .A(n2149), .B(n101), .Z(n103) );
  IV U118 ( .A(a[46]), .Z(n104) );
  NOR U119 ( .A(n103), .B(n104), .Z(n105) );
  NOR U120 ( .A(n102), .B(n105), .Z(n106) );
  IV U121 ( .A(n106), .Z(n2151) );
  IV U122 ( .A(n2155), .Z(n107) );
  IV U123 ( .A(b[49]), .Z(n108) );
  NOR U124 ( .A(n107), .B(n108), .Z(n109) );
  XOR U125 ( .A(n2155), .B(n108), .Z(n110) );
  IV U126 ( .A(a[49]), .Z(n111) );
  NOR U127 ( .A(n110), .B(n111), .Z(n112) );
  NOR U128 ( .A(n109), .B(n112), .Z(n113) );
  IV U129 ( .A(n113), .Z(n2159) );
  IV U130 ( .A(n2163), .Z(n114) );
  IV U131 ( .A(b[52]), .Z(n115) );
  NOR U132 ( .A(n114), .B(n115), .Z(n116) );
  XOR U133 ( .A(n2163), .B(n115), .Z(n117) );
  IV U134 ( .A(a[52]), .Z(n118) );
  NOR U135 ( .A(n117), .B(n118), .Z(n119) );
  NOR U136 ( .A(n116), .B(n119), .Z(n120) );
  IV U137 ( .A(n120), .Z(n2165) );
  IV U138 ( .A(n2169), .Z(n121) );
  IV U139 ( .A(b[55]), .Z(n122) );
  NOR U140 ( .A(n121), .B(n122), .Z(n123) );
  XOR U141 ( .A(n2169), .B(n122), .Z(n124) );
  IV U142 ( .A(a[55]), .Z(n125) );
  NOR U143 ( .A(n124), .B(n125), .Z(n126) );
  NOR U144 ( .A(n123), .B(n126), .Z(n127) );
  IV U145 ( .A(n127), .Z(n2171) );
  IV U146 ( .A(n2175), .Z(n128) );
  IV U147 ( .A(b[58]), .Z(n129) );
  NOR U148 ( .A(n128), .B(n129), .Z(n130) );
  XOR U149 ( .A(n2175), .B(n129), .Z(n131) );
  IV U150 ( .A(a[58]), .Z(n132) );
  NOR U151 ( .A(n131), .B(n132), .Z(n133) );
  NOR U152 ( .A(n130), .B(n133), .Z(n134) );
  IV U153 ( .A(n134), .Z(n2177) );
  IV U154 ( .A(n2183), .Z(n135) );
  IV U155 ( .A(b[61]), .Z(n136) );
  NOR U156 ( .A(n135), .B(n136), .Z(n137) );
  XOR U157 ( .A(n2183), .B(n136), .Z(n138) );
  IV U158 ( .A(a[61]), .Z(n139) );
  NOR U159 ( .A(n138), .B(n139), .Z(n140) );
  NOR U160 ( .A(n137), .B(n140), .Z(n141) );
  IV U161 ( .A(n141), .Z(n2185) );
  IV U162 ( .A(n2189), .Z(n142) );
  IV U163 ( .A(b[64]), .Z(n143) );
  NOR U164 ( .A(n142), .B(n143), .Z(n144) );
  XOR U165 ( .A(n2189), .B(n143), .Z(n145) );
  IV U166 ( .A(a[64]), .Z(n146) );
  NOR U167 ( .A(n145), .B(n146), .Z(n147) );
  NOR U168 ( .A(n144), .B(n147), .Z(n148) );
  IV U169 ( .A(n148), .Z(n2191) );
  IV U170 ( .A(n2195), .Z(n149) );
  IV U171 ( .A(b[67]), .Z(n150) );
  NOR U172 ( .A(n149), .B(n150), .Z(n151) );
  XOR U173 ( .A(n2195), .B(n150), .Z(n152) );
  IV U174 ( .A(a[67]), .Z(n153) );
  NOR U175 ( .A(n152), .B(n153), .Z(n154) );
  NOR U176 ( .A(n151), .B(n154), .Z(n155) );
  IV U177 ( .A(n155), .Z(n2197) );
  IV U178 ( .A(n2203), .Z(n156) );
  IV U179 ( .A(b[70]), .Z(n157) );
  NOR U180 ( .A(n156), .B(n157), .Z(n158) );
  XOR U181 ( .A(n2203), .B(n157), .Z(n159) );
  IV U182 ( .A(a[70]), .Z(n160) );
  NOR U183 ( .A(n159), .B(n160), .Z(n161) );
  NOR U184 ( .A(n158), .B(n161), .Z(n162) );
  IV U185 ( .A(n162), .Z(n2205) );
  IV U186 ( .A(n2209), .Z(n163) );
  IV U187 ( .A(b[73]), .Z(n164) );
  NOR U188 ( .A(n163), .B(n164), .Z(n165) );
  XOR U189 ( .A(n2209), .B(n164), .Z(n166) );
  IV U190 ( .A(a[73]), .Z(n167) );
  NOR U191 ( .A(n166), .B(n167), .Z(n168) );
  NOR U192 ( .A(n165), .B(n168), .Z(n169) );
  IV U193 ( .A(n169), .Z(n2211) );
  IV U194 ( .A(n2215), .Z(n170) );
  IV U195 ( .A(b[76]), .Z(n171) );
  NOR U196 ( .A(n170), .B(n171), .Z(n172) );
  XOR U197 ( .A(n2215), .B(n171), .Z(n173) );
  IV U198 ( .A(a[76]), .Z(n174) );
  NOR U199 ( .A(n173), .B(n174), .Z(n175) );
  NOR U200 ( .A(n172), .B(n175), .Z(n176) );
  IV U201 ( .A(n176), .Z(n2217) );
  IV U202 ( .A(n2221), .Z(n177) );
  IV U203 ( .A(b[79]), .Z(n178) );
  NOR U204 ( .A(n177), .B(n178), .Z(n179) );
  XOR U205 ( .A(n2221), .B(n178), .Z(n180) );
  IV U206 ( .A(a[79]), .Z(n181) );
  NOR U207 ( .A(n180), .B(n181), .Z(n182) );
  NOR U208 ( .A(n179), .B(n182), .Z(n183) );
  IV U209 ( .A(n183), .Z(n2225) );
  IV U210 ( .A(n2229), .Z(n184) );
  IV U211 ( .A(b[82]), .Z(n185) );
  NOR U212 ( .A(n184), .B(n185), .Z(n186) );
  XOR U213 ( .A(n2229), .B(n185), .Z(n187) );
  IV U214 ( .A(a[82]), .Z(n188) );
  NOR U215 ( .A(n187), .B(n188), .Z(n189) );
  NOR U216 ( .A(n186), .B(n189), .Z(n190) );
  IV U217 ( .A(n190), .Z(n2231) );
  IV U218 ( .A(n2235), .Z(n191) );
  IV U219 ( .A(b[85]), .Z(n192) );
  NOR U220 ( .A(n191), .B(n192), .Z(n193) );
  XOR U221 ( .A(n2235), .B(n192), .Z(n194) );
  IV U222 ( .A(a[85]), .Z(n195) );
  NOR U223 ( .A(n194), .B(n195), .Z(n196) );
  NOR U224 ( .A(n193), .B(n196), .Z(n197) );
  IV U225 ( .A(n197), .Z(n2237) );
  IV U226 ( .A(n2241), .Z(n198) );
  IV U227 ( .A(b[88]), .Z(n199) );
  NOR U228 ( .A(n198), .B(n199), .Z(n200) );
  XOR U229 ( .A(n2241), .B(n199), .Z(n201) );
  IV U230 ( .A(a[88]), .Z(n202) );
  NOR U231 ( .A(n201), .B(n202), .Z(n203) );
  NOR U232 ( .A(n200), .B(n203), .Z(n204) );
  IV U233 ( .A(n204), .Z(n2243) );
  IV U234 ( .A(n2249), .Z(n205) );
  IV U235 ( .A(b[91]), .Z(n206) );
  NOR U236 ( .A(n205), .B(n206), .Z(n207) );
  XOR U237 ( .A(n2249), .B(n206), .Z(n208) );
  IV U238 ( .A(a[91]), .Z(n209) );
  NOR U239 ( .A(n208), .B(n209), .Z(n210) );
  NOR U240 ( .A(n207), .B(n210), .Z(n211) );
  IV U241 ( .A(n211), .Z(n2251) );
  IV U242 ( .A(n2255), .Z(n212) );
  IV U243 ( .A(b[94]), .Z(n213) );
  NOR U244 ( .A(n212), .B(n213), .Z(n214) );
  XOR U245 ( .A(n2255), .B(n213), .Z(n215) );
  IV U246 ( .A(a[94]), .Z(n216) );
  NOR U247 ( .A(n215), .B(n216), .Z(n217) );
  NOR U248 ( .A(n214), .B(n217), .Z(n218) );
  IV U249 ( .A(n218), .Z(n2257) );
  IV U250 ( .A(n2261), .Z(n219) );
  IV U251 ( .A(b[97]), .Z(n220) );
  NOR U252 ( .A(n219), .B(n220), .Z(n221) );
  XOR U253 ( .A(n2261), .B(n220), .Z(n222) );
  IV U254 ( .A(a[97]), .Z(n223) );
  NOR U255 ( .A(n222), .B(n223), .Z(n224) );
  NOR U256 ( .A(n221), .B(n224), .Z(n225) );
  IV U257 ( .A(n225), .Z(n2263) );
  IV U258 ( .A(n1726), .Z(n226) );
  IV U259 ( .A(b[100]), .Z(n227) );
  NOR U260 ( .A(n226), .B(n227), .Z(n228) );
  XOR U261 ( .A(n1726), .B(n227), .Z(n229) );
  IV U262 ( .A(a[100]), .Z(n230) );
  NOR U263 ( .A(n229), .B(n230), .Z(n231) );
  NOR U264 ( .A(n228), .B(n231), .Z(n232) );
  IV U265 ( .A(n232), .Z(n1728) );
  IV U266 ( .A(n1732), .Z(n233) );
  IV U267 ( .A(b[103]), .Z(n234) );
  NOR U268 ( .A(n233), .B(n234), .Z(n235) );
  XOR U269 ( .A(n1732), .B(n234), .Z(n236) );
  IV U270 ( .A(a[103]), .Z(n237) );
  NOR U271 ( .A(n236), .B(n237), .Z(n238) );
  NOR U272 ( .A(n235), .B(n238), .Z(n239) );
  IV U273 ( .A(n239), .Z(n1734) );
  IV U274 ( .A(n1738), .Z(n240) );
  IV U275 ( .A(b[106]), .Z(n241) );
  NOR U276 ( .A(n240), .B(n241), .Z(n242) );
  XOR U277 ( .A(n1738), .B(n241), .Z(n243) );
  IV U278 ( .A(a[106]), .Z(n244) );
  NOR U279 ( .A(n243), .B(n244), .Z(n245) );
  NOR U280 ( .A(n242), .B(n245), .Z(n246) );
  IV U281 ( .A(n246), .Z(n1740) );
  IV U282 ( .A(n1746), .Z(n247) );
  IV U283 ( .A(b[109]), .Z(n248) );
  NOR U284 ( .A(n247), .B(n248), .Z(n249) );
  XOR U285 ( .A(n1746), .B(n248), .Z(n250) );
  IV U286 ( .A(a[109]), .Z(n251) );
  NOR U287 ( .A(n250), .B(n251), .Z(n252) );
  NOR U288 ( .A(n249), .B(n252), .Z(n253) );
  IV U289 ( .A(n253), .Z(n1748) );
  IV U290 ( .A(n1752), .Z(n254) );
  IV U291 ( .A(b[112]), .Z(n255) );
  NOR U292 ( .A(n254), .B(n255), .Z(n256) );
  XOR U293 ( .A(n1752), .B(n255), .Z(n257) );
  IV U294 ( .A(a[112]), .Z(n258) );
  NOR U295 ( .A(n257), .B(n258), .Z(n259) );
  NOR U296 ( .A(n256), .B(n259), .Z(n260) );
  IV U297 ( .A(n260), .Z(n1754) );
  IV U298 ( .A(n1758), .Z(n261) );
  IV U299 ( .A(b[115]), .Z(n262) );
  NOR U300 ( .A(n261), .B(n262), .Z(n263) );
  XOR U301 ( .A(n1758), .B(n262), .Z(n264) );
  IV U302 ( .A(a[115]), .Z(n265) );
  NOR U303 ( .A(n264), .B(n265), .Z(n266) );
  NOR U304 ( .A(n263), .B(n266), .Z(n267) );
  IV U305 ( .A(n267), .Z(n1760) );
  IV U306 ( .A(n1764), .Z(n268) );
  IV U307 ( .A(b[118]), .Z(n269) );
  NOR U308 ( .A(n268), .B(n269), .Z(n270) );
  XOR U309 ( .A(n1764), .B(n269), .Z(n271) );
  IV U310 ( .A(a[118]), .Z(n272) );
  NOR U311 ( .A(n271), .B(n272), .Z(n273) );
  NOR U312 ( .A(n270), .B(n273), .Z(n274) );
  IV U313 ( .A(n274), .Z(n1768) );
  IV U314 ( .A(n1772), .Z(n275) );
  IV U315 ( .A(b[121]), .Z(n276) );
  NOR U316 ( .A(n275), .B(n276), .Z(n277) );
  XOR U317 ( .A(n1772), .B(n276), .Z(n278) );
  IV U318 ( .A(a[121]), .Z(n279) );
  NOR U319 ( .A(n278), .B(n279), .Z(n280) );
  NOR U320 ( .A(n277), .B(n280), .Z(n281) );
  IV U321 ( .A(n281), .Z(n1774) );
  IV U322 ( .A(n1778), .Z(n282) );
  IV U323 ( .A(b[124]), .Z(n283) );
  NOR U324 ( .A(n282), .B(n283), .Z(n284) );
  XOR U325 ( .A(n1778), .B(n283), .Z(n285) );
  IV U326 ( .A(a[124]), .Z(n286) );
  NOR U327 ( .A(n285), .B(n286), .Z(n287) );
  NOR U328 ( .A(n284), .B(n287), .Z(n288) );
  IV U329 ( .A(n288), .Z(n1780) );
  IV U330 ( .A(n1784), .Z(n289) );
  IV U331 ( .A(b[127]), .Z(n290) );
  NOR U332 ( .A(n289), .B(n290), .Z(n291) );
  XOR U333 ( .A(n1784), .B(n290), .Z(n292) );
  IV U334 ( .A(a[127]), .Z(n293) );
  NOR U335 ( .A(n292), .B(n293), .Z(n294) );
  NOR U336 ( .A(n291), .B(n294), .Z(n295) );
  IV U337 ( .A(n295), .Z(n1786) );
  IV U338 ( .A(n1792), .Z(n296) );
  IV U339 ( .A(b[130]), .Z(n297) );
  NOR U340 ( .A(n296), .B(n297), .Z(n298) );
  XOR U341 ( .A(n1792), .B(n297), .Z(n299) );
  IV U342 ( .A(a[130]), .Z(n300) );
  NOR U343 ( .A(n299), .B(n300), .Z(n301) );
  NOR U344 ( .A(n298), .B(n301), .Z(n302) );
  IV U345 ( .A(n302), .Z(n1794) );
  IV U346 ( .A(n1798), .Z(n303) );
  IV U347 ( .A(b[133]), .Z(n304) );
  NOR U348 ( .A(n303), .B(n304), .Z(n305) );
  XOR U349 ( .A(n1798), .B(n304), .Z(n306) );
  IV U350 ( .A(a[133]), .Z(n307) );
  NOR U351 ( .A(n306), .B(n307), .Z(n308) );
  NOR U352 ( .A(n305), .B(n308), .Z(n309) );
  IV U353 ( .A(n309), .Z(n1800) );
  IV U354 ( .A(n1804), .Z(n310) );
  IV U355 ( .A(b[136]), .Z(n311) );
  NOR U356 ( .A(n310), .B(n311), .Z(n312) );
  XOR U357 ( .A(n1804), .B(n311), .Z(n313) );
  IV U358 ( .A(a[136]), .Z(n314) );
  NOR U359 ( .A(n313), .B(n314), .Z(n315) );
  NOR U360 ( .A(n312), .B(n315), .Z(n316) );
  IV U361 ( .A(n316), .Z(n1806) );
  IV U362 ( .A(n1812), .Z(n317) );
  IV U363 ( .A(b[139]), .Z(n318) );
  NOR U364 ( .A(n317), .B(n318), .Z(n319) );
  XOR U365 ( .A(n1812), .B(n318), .Z(n320) );
  IV U366 ( .A(a[139]), .Z(n321) );
  NOR U367 ( .A(n320), .B(n321), .Z(n322) );
  NOR U368 ( .A(n319), .B(n322), .Z(n323) );
  IV U369 ( .A(n323), .Z(n1814) );
  IV U370 ( .A(n1818), .Z(n324) );
  IV U371 ( .A(b[142]), .Z(n325) );
  NOR U372 ( .A(n324), .B(n325), .Z(n326) );
  XOR U373 ( .A(n1818), .B(n325), .Z(n327) );
  IV U374 ( .A(a[142]), .Z(n328) );
  NOR U375 ( .A(n327), .B(n328), .Z(n329) );
  NOR U376 ( .A(n326), .B(n329), .Z(n330) );
  IV U377 ( .A(n330), .Z(n1820) );
  IV U378 ( .A(n1824), .Z(n331) );
  IV U379 ( .A(b[145]), .Z(n332) );
  NOR U380 ( .A(n331), .B(n332), .Z(n333) );
  XOR U381 ( .A(n1824), .B(n332), .Z(n334) );
  IV U382 ( .A(a[145]), .Z(n335) );
  NOR U383 ( .A(n334), .B(n335), .Z(n336) );
  NOR U384 ( .A(n333), .B(n336), .Z(n337) );
  IV U385 ( .A(n337), .Z(n1826) );
  IV U386 ( .A(n1830), .Z(n338) );
  IV U387 ( .A(b[148]), .Z(n339) );
  NOR U388 ( .A(n338), .B(n339), .Z(n340) );
  XOR U389 ( .A(n1830), .B(n339), .Z(n341) );
  IV U390 ( .A(a[148]), .Z(n342) );
  NOR U391 ( .A(n341), .B(n342), .Z(n343) );
  NOR U392 ( .A(n340), .B(n343), .Z(n344) );
  IV U393 ( .A(n344), .Z(n1834) );
  IV U394 ( .A(n1838), .Z(n345) );
  IV U395 ( .A(b[151]), .Z(n346) );
  NOR U396 ( .A(n345), .B(n346), .Z(n347) );
  XOR U397 ( .A(n1838), .B(n346), .Z(n348) );
  IV U398 ( .A(a[151]), .Z(n349) );
  NOR U399 ( .A(n348), .B(n349), .Z(n350) );
  NOR U400 ( .A(n347), .B(n350), .Z(n351) );
  IV U401 ( .A(n351), .Z(n1840) );
  IV U402 ( .A(n1844), .Z(n352) );
  IV U403 ( .A(b[154]), .Z(n353) );
  NOR U404 ( .A(n352), .B(n353), .Z(n354) );
  XOR U405 ( .A(n1844), .B(n353), .Z(n355) );
  IV U406 ( .A(a[154]), .Z(n356) );
  NOR U407 ( .A(n355), .B(n356), .Z(n357) );
  NOR U408 ( .A(n354), .B(n357), .Z(n358) );
  IV U409 ( .A(n358), .Z(n1846) );
  IV U410 ( .A(n1850), .Z(n359) );
  IV U411 ( .A(b[157]), .Z(n360) );
  NOR U412 ( .A(n359), .B(n360), .Z(n361) );
  XOR U413 ( .A(n1850), .B(n360), .Z(n362) );
  IV U414 ( .A(a[157]), .Z(n363) );
  NOR U415 ( .A(n362), .B(n363), .Z(n364) );
  NOR U416 ( .A(n361), .B(n364), .Z(n365) );
  IV U417 ( .A(n365), .Z(n1852) );
  IV U418 ( .A(n1858), .Z(n366) );
  IV U419 ( .A(b[160]), .Z(n367) );
  NOR U420 ( .A(n366), .B(n367), .Z(n368) );
  XOR U421 ( .A(n1858), .B(n367), .Z(n369) );
  IV U422 ( .A(a[160]), .Z(n370) );
  NOR U423 ( .A(n369), .B(n370), .Z(n371) );
  NOR U424 ( .A(n368), .B(n371), .Z(n372) );
  IV U425 ( .A(n372), .Z(n1860) );
  IV U426 ( .A(n1864), .Z(n373) );
  IV U427 ( .A(b[163]), .Z(n374) );
  NOR U428 ( .A(n373), .B(n374), .Z(n375) );
  XOR U429 ( .A(n1864), .B(n374), .Z(n376) );
  IV U430 ( .A(a[163]), .Z(n377) );
  NOR U431 ( .A(n376), .B(n377), .Z(n378) );
  NOR U432 ( .A(n375), .B(n378), .Z(n379) );
  IV U433 ( .A(n379), .Z(n1866) );
  IV U434 ( .A(n1870), .Z(n380) );
  IV U435 ( .A(b[166]), .Z(n381) );
  NOR U436 ( .A(n380), .B(n381), .Z(n382) );
  XOR U437 ( .A(n1870), .B(n381), .Z(n383) );
  IV U438 ( .A(a[166]), .Z(n384) );
  NOR U439 ( .A(n383), .B(n384), .Z(n385) );
  NOR U440 ( .A(n382), .B(n385), .Z(n386) );
  IV U441 ( .A(n386), .Z(n1872) );
  IV U442 ( .A(n1878), .Z(n387) );
  IV U443 ( .A(b[169]), .Z(n388) );
  NOR U444 ( .A(n387), .B(n388), .Z(n389) );
  XOR U445 ( .A(n1878), .B(n388), .Z(n390) );
  IV U446 ( .A(a[169]), .Z(n391) );
  NOR U447 ( .A(n390), .B(n391), .Z(n392) );
  NOR U448 ( .A(n389), .B(n392), .Z(n393) );
  IV U449 ( .A(n393), .Z(n1880) );
  IV U450 ( .A(n1884), .Z(n394) );
  IV U451 ( .A(b[172]), .Z(n395) );
  NOR U452 ( .A(n394), .B(n395), .Z(n396) );
  XOR U453 ( .A(n1884), .B(n395), .Z(n397) );
  IV U454 ( .A(a[172]), .Z(n398) );
  NOR U455 ( .A(n397), .B(n398), .Z(n399) );
  NOR U456 ( .A(n396), .B(n399), .Z(n400) );
  IV U457 ( .A(n400), .Z(n1886) );
  IV U458 ( .A(n1890), .Z(n401) );
  IV U459 ( .A(b[175]), .Z(n402) );
  NOR U460 ( .A(n401), .B(n402), .Z(n403) );
  XOR U461 ( .A(n1890), .B(n402), .Z(n404) );
  IV U462 ( .A(a[175]), .Z(n405) );
  NOR U463 ( .A(n404), .B(n405), .Z(n406) );
  NOR U464 ( .A(n403), .B(n406), .Z(n407) );
  IV U465 ( .A(n407), .Z(n1892) );
  IV U466 ( .A(n1896), .Z(n408) );
  IV U467 ( .A(b[178]), .Z(n409) );
  NOR U468 ( .A(n408), .B(n409), .Z(n410) );
  XOR U469 ( .A(n1896), .B(n409), .Z(n411) );
  IV U470 ( .A(a[178]), .Z(n412) );
  NOR U471 ( .A(n411), .B(n412), .Z(n413) );
  NOR U472 ( .A(n410), .B(n413), .Z(n414) );
  IV U473 ( .A(n414), .Z(n1900) );
  IV U474 ( .A(n1904), .Z(n415) );
  IV U475 ( .A(b[181]), .Z(n416) );
  NOR U476 ( .A(n415), .B(n416), .Z(n417) );
  XOR U477 ( .A(n1904), .B(n416), .Z(n418) );
  IV U478 ( .A(a[181]), .Z(n419) );
  NOR U479 ( .A(n418), .B(n419), .Z(n420) );
  NOR U480 ( .A(n417), .B(n420), .Z(n421) );
  IV U481 ( .A(n421), .Z(n1906) );
  IV U482 ( .A(n1910), .Z(n422) );
  IV U483 ( .A(b[184]), .Z(n423) );
  NOR U484 ( .A(n422), .B(n423), .Z(n424) );
  XOR U485 ( .A(n1910), .B(n423), .Z(n425) );
  IV U486 ( .A(a[184]), .Z(n426) );
  NOR U487 ( .A(n425), .B(n426), .Z(n427) );
  NOR U488 ( .A(n424), .B(n427), .Z(n428) );
  IV U489 ( .A(n428), .Z(n1912) );
  IV U490 ( .A(n1916), .Z(n429) );
  IV U491 ( .A(b[187]), .Z(n430) );
  NOR U492 ( .A(n429), .B(n430), .Z(n431) );
  XOR U493 ( .A(n1916), .B(n430), .Z(n432) );
  IV U494 ( .A(a[187]), .Z(n433) );
  NOR U495 ( .A(n432), .B(n433), .Z(n434) );
  NOR U496 ( .A(n431), .B(n434), .Z(n435) );
  IV U497 ( .A(n435), .Z(n1918) );
  IV U498 ( .A(n1924), .Z(n436) );
  IV U499 ( .A(b[190]), .Z(n437) );
  NOR U500 ( .A(n436), .B(n437), .Z(n438) );
  XOR U501 ( .A(n1924), .B(n437), .Z(n439) );
  IV U502 ( .A(a[190]), .Z(n440) );
  NOR U503 ( .A(n439), .B(n440), .Z(n441) );
  NOR U504 ( .A(n438), .B(n441), .Z(n442) );
  IV U505 ( .A(n442), .Z(n1926) );
  IV U506 ( .A(n1930), .Z(n443) );
  IV U507 ( .A(b[193]), .Z(n444) );
  NOR U508 ( .A(n443), .B(n444), .Z(n445) );
  XOR U509 ( .A(n1930), .B(n444), .Z(n446) );
  IV U510 ( .A(a[193]), .Z(n447) );
  NOR U511 ( .A(n446), .B(n447), .Z(n448) );
  NOR U512 ( .A(n445), .B(n448), .Z(n449) );
  IV U513 ( .A(n449), .Z(n1932) );
  IV U514 ( .A(n1936), .Z(n450) );
  IV U515 ( .A(b[196]), .Z(n451) );
  NOR U516 ( .A(n450), .B(n451), .Z(n452) );
  XOR U517 ( .A(n1936), .B(n451), .Z(n453) );
  IV U518 ( .A(a[196]), .Z(n454) );
  NOR U519 ( .A(n453), .B(n454), .Z(n455) );
  NOR U520 ( .A(n452), .B(n455), .Z(n456) );
  IV U521 ( .A(n456), .Z(n1938) );
  IV U522 ( .A(n1946), .Z(n457) );
  IV U523 ( .A(b[199]), .Z(n458) );
  NOR U524 ( .A(n457), .B(n458), .Z(n459) );
  XOR U525 ( .A(n1946), .B(n458), .Z(n460) );
  IV U526 ( .A(a[199]), .Z(n461) );
  NOR U527 ( .A(n460), .B(n461), .Z(n462) );
  NOR U528 ( .A(n459), .B(n462), .Z(n463) );
  IV U529 ( .A(n463), .Z(n1948) );
  IV U530 ( .A(n1952), .Z(n464) );
  IV U531 ( .A(b[202]), .Z(n465) );
  NOR U532 ( .A(n464), .B(n465), .Z(n466) );
  XOR U533 ( .A(n1952), .B(n465), .Z(n467) );
  IV U534 ( .A(a[202]), .Z(n468) );
  NOR U535 ( .A(n467), .B(n468), .Z(n469) );
  NOR U536 ( .A(n466), .B(n469), .Z(n470) );
  IV U537 ( .A(n470), .Z(n1954) );
  IV U538 ( .A(n1958), .Z(n471) );
  IV U539 ( .A(b[205]), .Z(n472) );
  NOR U540 ( .A(n471), .B(n472), .Z(n473) );
  XOR U541 ( .A(n1958), .B(n472), .Z(n474) );
  IV U542 ( .A(a[205]), .Z(n475) );
  NOR U543 ( .A(n474), .B(n475), .Z(n476) );
  NOR U544 ( .A(n473), .B(n476), .Z(n477) );
  IV U545 ( .A(n477), .Z(n1960) );
  IV U546 ( .A(n1964), .Z(n478) );
  IV U547 ( .A(b[208]), .Z(n479) );
  NOR U548 ( .A(n478), .B(n479), .Z(n480) );
  XOR U549 ( .A(n1964), .B(n479), .Z(n481) );
  IV U550 ( .A(a[208]), .Z(n482) );
  NOR U551 ( .A(n481), .B(n482), .Z(n483) );
  NOR U552 ( .A(n480), .B(n483), .Z(n484) );
  IV U553 ( .A(n484), .Z(n1968) );
  IV U554 ( .A(n1972), .Z(n485) );
  IV U555 ( .A(b[211]), .Z(n486) );
  NOR U556 ( .A(n485), .B(n486), .Z(n487) );
  XOR U557 ( .A(n1972), .B(n486), .Z(n488) );
  IV U558 ( .A(a[211]), .Z(n489) );
  NOR U559 ( .A(n488), .B(n489), .Z(n490) );
  NOR U560 ( .A(n487), .B(n490), .Z(n491) );
  IV U561 ( .A(n491), .Z(n1974) );
  IV U562 ( .A(n1978), .Z(n492) );
  IV U563 ( .A(b[214]), .Z(n493) );
  NOR U564 ( .A(n492), .B(n493), .Z(n494) );
  XOR U565 ( .A(n1978), .B(n493), .Z(n495) );
  IV U566 ( .A(a[214]), .Z(n496) );
  NOR U567 ( .A(n495), .B(n496), .Z(n497) );
  NOR U568 ( .A(n494), .B(n497), .Z(n498) );
  IV U569 ( .A(n498), .Z(n1980) );
  IV U570 ( .A(n1984), .Z(n499) );
  IV U571 ( .A(b[217]), .Z(n500) );
  NOR U572 ( .A(n499), .B(n500), .Z(n501) );
  XOR U573 ( .A(n1984), .B(n500), .Z(n502) );
  IV U574 ( .A(a[217]), .Z(n503) );
  NOR U575 ( .A(n502), .B(n503), .Z(n504) );
  NOR U576 ( .A(n501), .B(n504), .Z(n505) );
  IV U577 ( .A(n505), .Z(n1986) );
  IV U578 ( .A(n1992), .Z(n506) );
  IV U579 ( .A(b[220]), .Z(n507) );
  NOR U580 ( .A(n506), .B(n507), .Z(n508) );
  XOR U581 ( .A(n1992), .B(n507), .Z(n509) );
  IV U582 ( .A(a[220]), .Z(n510) );
  NOR U583 ( .A(n509), .B(n510), .Z(n511) );
  NOR U584 ( .A(n508), .B(n511), .Z(n512) );
  IV U585 ( .A(n512), .Z(n1994) );
  IV U586 ( .A(n1998), .Z(n513) );
  IV U587 ( .A(b[223]), .Z(n514) );
  NOR U588 ( .A(n513), .B(n514), .Z(n515) );
  XOR U589 ( .A(n1998), .B(n514), .Z(n516) );
  IV U590 ( .A(a[223]), .Z(n517) );
  NOR U591 ( .A(n516), .B(n517), .Z(n518) );
  NOR U592 ( .A(n515), .B(n518), .Z(n519) );
  IV U593 ( .A(n519), .Z(n2000) );
  IV U594 ( .A(n2004), .Z(n520) );
  IV U595 ( .A(b[226]), .Z(n521) );
  NOR U596 ( .A(n520), .B(n521), .Z(n522) );
  XOR U597 ( .A(n2004), .B(n521), .Z(n523) );
  IV U598 ( .A(a[226]), .Z(n524) );
  NOR U599 ( .A(n523), .B(n524), .Z(n525) );
  NOR U600 ( .A(n522), .B(n525), .Z(n526) );
  IV U601 ( .A(n526), .Z(n2006) );
  IV U602 ( .A(n2012), .Z(n527) );
  IV U603 ( .A(b[229]), .Z(n528) );
  NOR U604 ( .A(n527), .B(n528), .Z(n529) );
  XOR U605 ( .A(n2012), .B(n528), .Z(n530) );
  IV U606 ( .A(a[229]), .Z(n531) );
  NOR U607 ( .A(n530), .B(n531), .Z(n532) );
  NOR U608 ( .A(n529), .B(n532), .Z(n533) );
  IV U609 ( .A(n533), .Z(n2014) );
  IV U610 ( .A(n2018), .Z(n534) );
  IV U611 ( .A(b[232]), .Z(n535) );
  NOR U612 ( .A(n534), .B(n535), .Z(n536) );
  XOR U613 ( .A(n2018), .B(n535), .Z(n537) );
  IV U614 ( .A(a[232]), .Z(n538) );
  NOR U615 ( .A(n537), .B(n538), .Z(n539) );
  NOR U616 ( .A(n536), .B(n539), .Z(n540) );
  IV U617 ( .A(n540), .Z(n2020) );
  IV U618 ( .A(n2024), .Z(n541) );
  IV U619 ( .A(b[235]), .Z(n542) );
  NOR U620 ( .A(n541), .B(n542), .Z(n543) );
  XOR U621 ( .A(n2024), .B(n542), .Z(n544) );
  IV U622 ( .A(a[235]), .Z(n545) );
  NOR U623 ( .A(n544), .B(n545), .Z(n546) );
  NOR U624 ( .A(n543), .B(n546), .Z(n547) );
  IV U625 ( .A(n547), .Z(n2026) );
  IV U626 ( .A(n2030), .Z(n548) );
  IV U627 ( .A(b[238]), .Z(n549) );
  NOR U628 ( .A(n548), .B(n549), .Z(n550) );
  XOR U629 ( .A(n2030), .B(n549), .Z(n551) );
  IV U630 ( .A(a[238]), .Z(n552) );
  NOR U631 ( .A(n551), .B(n552), .Z(n553) );
  NOR U632 ( .A(n550), .B(n553), .Z(n554) );
  IV U633 ( .A(n554), .Z(n2034) );
  IV U634 ( .A(n2038), .Z(n555) );
  IV U635 ( .A(b[241]), .Z(n556) );
  NOR U636 ( .A(n555), .B(n556), .Z(n557) );
  XOR U637 ( .A(n2038), .B(n556), .Z(n558) );
  IV U638 ( .A(a[241]), .Z(n559) );
  NOR U639 ( .A(n558), .B(n559), .Z(n560) );
  NOR U640 ( .A(n557), .B(n560), .Z(n561) );
  IV U641 ( .A(n561), .Z(n2040) );
  IV U642 ( .A(n2044), .Z(n562) );
  IV U643 ( .A(b[244]), .Z(n563) );
  NOR U644 ( .A(n562), .B(n563), .Z(n564) );
  XOR U645 ( .A(n2044), .B(n563), .Z(n565) );
  IV U646 ( .A(a[244]), .Z(n566) );
  NOR U647 ( .A(n565), .B(n566), .Z(n567) );
  NOR U648 ( .A(n564), .B(n567), .Z(n568) );
  IV U649 ( .A(n568), .Z(n2046) );
  IV U650 ( .A(n2179), .Z(n569) );
  IV U651 ( .A(b[5]), .Z(n570) );
  NOR U652 ( .A(n569), .B(n570), .Z(n571) );
  XOR U653 ( .A(n2179), .B(n570), .Z(n572) );
  IV U654 ( .A(a[5]), .Z(n573) );
  NOR U655 ( .A(n572), .B(n573), .Z(n574) );
  NOR U656 ( .A(n571), .B(n574), .Z(n575) );
  IV U657 ( .A(n575), .Z(n2201) );
  IV U658 ( .A(n2245), .Z(n576) );
  IV U659 ( .A(b[8]), .Z(n577) );
  NOR U660 ( .A(n576), .B(n577), .Z(n578) );
  XOR U661 ( .A(n2245), .B(n577), .Z(n579) );
  IV U662 ( .A(a[8]), .Z(n580) );
  NOR U663 ( .A(n579), .B(n580), .Z(n581) );
  NOR U664 ( .A(n578), .B(n581), .Z(n582) );
  IV U665 ( .A(n582), .Z(n2267) );
  IV U666 ( .A(n1766), .Z(n583) );
  IV U667 ( .A(b[11]), .Z(n584) );
  NOR U668 ( .A(n583), .B(n584), .Z(n585) );
  XOR U669 ( .A(n1766), .B(n584), .Z(n586) );
  IV U670 ( .A(a[11]), .Z(n587) );
  NOR U671 ( .A(n586), .B(n587), .Z(n588) );
  NOR U672 ( .A(n585), .B(n588), .Z(n589) );
  IV U673 ( .A(n589), .Z(n1788) );
  IV U674 ( .A(n1832), .Z(n590) );
  IV U675 ( .A(b[14]), .Z(n591) );
  NOR U676 ( .A(n590), .B(n591), .Z(n592) );
  XOR U677 ( .A(n1832), .B(n591), .Z(n593) );
  IV U678 ( .A(a[14]), .Z(n594) );
  NOR U679 ( .A(n593), .B(n594), .Z(n595) );
  NOR U680 ( .A(n592), .B(n595), .Z(n596) );
  IV U681 ( .A(n596), .Z(n1854) );
  IV U682 ( .A(n1898), .Z(n597) );
  IV U683 ( .A(b[17]), .Z(n598) );
  NOR U684 ( .A(n597), .B(n598), .Z(n599) );
  XOR U685 ( .A(n1898), .B(n598), .Z(n600) );
  IV U686 ( .A(a[17]), .Z(n601) );
  NOR U687 ( .A(n600), .B(n601), .Z(n602) );
  NOR U688 ( .A(n599), .B(n602), .Z(n603) );
  IV U689 ( .A(n603), .Z(n1920) );
  IV U690 ( .A(n1966), .Z(n604) );
  IV U691 ( .A(b[20]), .Z(n605) );
  NOR U692 ( .A(n604), .B(n605), .Z(n606) );
  XOR U693 ( .A(n1966), .B(n605), .Z(n607) );
  IV U694 ( .A(a[20]), .Z(n608) );
  NOR U695 ( .A(n607), .B(n608), .Z(n609) );
  NOR U696 ( .A(n606), .B(n609), .Z(n610) );
  IV U697 ( .A(n610), .Z(n1988) );
  IV U698 ( .A(n2032), .Z(n611) );
  IV U699 ( .A(b[23]), .Z(n612) );
  NOR U700 ( .A(n611), .B(n612), .Z(n613) );
  XOR U701 ( .A(n2032), .B(n612), .Z(n614) );
  IV U702 ( .A(a[23]), .Z(n615) );
  NOR U703 ( .A(n614), .B(n615), .Z(n616) );
  NOR U704 ( .A(n613), .B(n616), .Z(n617) );
  IV U705 ( .A(n617), .Z(n2063) );
  IV U706 ( .A(n2104), .Z(n618) );
  IV U707 ( .A(b[26]), .Z(n619) );
  NOR U708 ( .A(n618), .B(n619), .Z(n620) );
  XOR U709 ( .A(n2104), .B(n619), .Z(n621) );
  IV U710 ( .A(a[26]), .Z(n622) );
  NOR U711 ( .A(n621), .B(n622), .Z(n623) );
  NOR U712 ( .A(n620), .B(n623), .Z(n624) );
  IV U713 ( .A(n624), .Z(n2106) );
  IV U714 ( .A(n2110), .Z(n625) );
  IV U715 ( .A(b[29]), .Z(n626) );
  NOR U716 ( .A(n625), .B(n626), .Z(n627) );
  XOR U717 ( .A(n2110), .B(n626), .Z(n628) );
  IV U718 ( .A(a[29]), .Z(n629) );
  NOR U719 ( .A(n628), .B(n629), .Z(n630) );
  NOR U720 ( .A(n627), .B(n630), .Z(n631) );
  IV U721 ( .A(n631), .Z(n2115) );
  IV U722 ( .A(n2119), .Z(n632) );
  IV U723 ( .A(b[32]), .Z(n633) );
  NOR U724 ( .A(n632), .B(n633), .Z(n634) );
  XOR U725 ( .A(n2119), .B(n633), .Z(n635) );
  IV U726 ( .A(a[32]), .Z(n636) );
  NOR U727 ( .A(n635), .B(n636), .Z(n637) );
  NOR U728 ( .A(n634), .B(n637), .Z(n638) );
  IV U729 ( .A(n638), .Z(n2121) );
  IV U730 ( .A(n2125), .Z(n639) );
  IV U731 ( .A(b[35]), .Z(n640) );
  NOR U732 ( .A(n639), .B(n640), .Z(n641) );
  XOR U733 ( .A(n2125), .B(n640), .Z(n642) );
  IV U734 ( .A(a[35]), .Z(n643) );
  NOR U735 ( .A(n642), .B(n643), .Z(n644) );
  NOR U736 ( .A(n641), .B(n644), .Z(n645) );
  IV U737 ( .A(n645), .Z(n2127) );
  IV U738 ( .A(n2131), .Z(n646) );
  IV U739 ( .A(b[38]), .Z(n647) );
  NOR U740 ( .A(n646), .B(n647), .Z(n648) );
  XOR U741 ( .A(n2131), .B(n647), .Z(n649) );
  IV U742 ( .A(a[38]), .Z(n650) );
  NOR U743 ( .A(n649), .B(n650), .Z(n651) );
  NOR U744 ( .A(n648), .B(n651), .Z(n652) );
  IV U745 ( .A(n652), .Z(n2133) );
  IV U746 ( .A(n2139), .Z(n653) );
  IV U747 ( .A(b[41]), .Z(n654) );
  NOR U748 ( .A(n653), .B(n654), .Z(n655) );
  XOR U749 ( .A(n2139), .B(n654), .Z(n656) );
  IV U750 ( .A(a[41]), .Z(n657) );
  NOR U751 ( .A(n656), .B(n657), .Z(n658) );
  NOR U752 ( .A(n655), .B(n658), .Z(n659) );
  IV U753 ( .A(n659), .Z(n2141) );
  IV U754 ( .A(n2145), .Z(n660) );
  IV U755 ( .A(b[44]), .Z(n661) );
  NOR U756 ( .A(n660), .B(n661), .Z(n662) );
  XOR U757 ( .A(n2145), .B(n661), .Z(n663) );
  IV U758 ( .A(a[44]), .Z(n664) );
  NOR U759 ( .A(n663), .B(n664), .Z(n665) );
  NOR U760 ( .A(n662), .B(n665), .Z(n666) );
  IV U761 ( .A(n666), .Z(n2147) );
  IV U762 ( .A(n2151), .Z(n667) );
  IV U763 ( .A(b[47]), .Z(n668) );
  NOR U764 ( .A(n667), .B(n668), .Z(n669) );
  XOR U765 ( .A(n2151), .B(n668), .Z(n670) );
  IV U766 ( .A(a[47]), .Z(n671) );
  NOR U767 ( .A(n670), .B(n671), .Z(n672) );
  NOR U768 ( .A(n669), .B(n672), .Z(n673) );
  IV U769 ( .A(n673), .Z(n2153) );
  IV U770 ( .A(n2159), .Z(n674) );
  IV U771 ( .A(b[50]), .Z(n675) );
  NOR U772 ( .A(n674), .B(n675), .Z(n676) );
  XOR U773 ( .A(n2159), .B(n675), .Z(n677) );
  IV U774 ( .A(a[50]), .Z(n678) );
  NOR U775 ( .A(n677), .B(n678), .Z(n679) );
  NOR U776 ( .A(n676), .B(n679), .Z(n680) );
  IV U777 ( .A(n680), .Z(n2161) );
  IV U778 ( .A(n2165), .Z(n681) );
  IV U779 ( .A(b[53]), .Z(n682) );
  NOR U780 ( .A(n681), .B(n682), .Z(n683) );
  XOR U781 ( .A(n2165), .B(n682), .Z(n684) );
  IV U782 ( .A(a[53]), .Z(n685) );
  NOR U783 ( .A(n684), .B(n685), .Z(n686) );
  NOR U784 ( .A(n683), .B(n686), .Z(n687) );
  IV U785 ( .A(n687), .Z(n2167) );
  IV U786 ( .A(n2171), .Z(n688) );
  IV U787 ( .A(b[56]), .Z(n689) );
  NOR U788 ( .A(n688), .B(n689), .Z(n690) );
  XOR U789 ( .A(n2171), .B(n689), .Z(n691) );
  IV U790 ( .A(a[56]), .Z(n692) );
  NOR U791 ( .A(n691), .B(n692), .Z(n693) );
  NOR U792 ( .A(n690), .B(n693), .Z(n694) );
  IV U793 ( .A(n694), .Z(n2173) );
  IV U794 ( .A(n2177), .Z(n695) );
  IV U795 ( .A(b[59]), .Z(n696) );
  NOR U796 ( .A(n695), .B(n696), .Z(n697) );
  XOR U797 ( .A(n2177), .B(n696), .Z(n698) );
  IV U798 ( .A(a[59]), .Z(n699) );
  NOR U799 ( .A(n698), .B(n699), .Z(n700) );
  NOR U800 ( .A(n697), .B(n700), .Z(n701) );
  IV U801 ( .A(n701), .Z(n2181) );
  IV U802 ( .A(n2185), .Z(n702) );
  IV U803 ( .A(b[62]), .Z(n703) );
  NOR U804 ( .A(n702), .B(n703), .Z(n704) );
  XOR U805 ( .A(n2185), .B(n703), .Z(n705) );
  IV U806 ( .A(a[62]), .Z(n706) );
  NOR U807 ( .A(n705), .B(n706), .Z(n707) );
  NOR U808 ( .A(n704), .B(n707), .Z(n708) );
  IV U809 ( .A(n708), .Z(n2187) );
  IV U810 ( .A(n2191), .Z(n709) );
  IV U811 ( .A(b[65]), .Z(n710) );
  NOR U812 ( .A(n709), .B(n710), .Z(n711) );
  XOR U813 ( .A(n2191), .B(n710), .Z(n712) );
  IV U814 ( .A(a[65]), .Z(n713) );
  NOR U815 ( .A(n712), .B(n713), .Z(n714) );
  NOR U816 ( .A(n711), .B(n714), .Z(n715) );
  IV U817 ( .A(n715), .Z(n2193) );
  IV U818 ( .A(n2197), .Z(n716) );
  IV U819 ( .A(b[68]), .Z(n717) );
  NOR U820 ( .A(n716), .B(n717), .Z(n718) );
  XOR U821 ( .A(n2197), .B(n717), .Z(n719) );
  IV U822 ( .A(a[68]), .Z(n720) );
  NOR U823 ( .A(n719), .B(n720), .Z(n721) );
  NOR U824 ( .A(n718), .B(n721), .Z(n722) );
  IV U825 ( .A(n722), .Z(n2199) );
  IV U826 ( .A(n2205), .Z(n723) );
  IV U827 ( .A(b[71]), .Z(n724) );
  NOR U828 ( .A(n723), .B(n724), .Z(n725) );
  XOR U829 ( .A(n2205), .B(n724), .Z(n726) );
  IV U830 ( .A(a[71]), .Z(n727) );
  NOR U831 ( .A(n726), .B(n727), .Z(n728) );
  NOR U832 ( .A(n725), .B(n728), .Z(n729) );
  IV U833 ( .A(n729), .Z(n2207) );
  IV U834 ( .A(n2211), .Z(n730) );
  IV U835 ( .A(b[74]), .Z(n731) );
  NOR U836 ( .A(n730), .B(n731), .Z(n732) );
  XOR U837 ( .A(n2211), .B(n731), .Z(n733) );
  IV U838 ( .A(a[74]), .Z(n734) );
  NOR U839 ( .A(n733), .B(n734), .Z(n735) );
  NOR U840 ( .A(n732), .B(n735), .Z(n736) );
  IV U841 ( .A(n736), .Z(n2213) );
  IV U842 ( .A(n2217), .Z(n737) );
  IV U843 ( .A(b[77]), .Z(n738) );
  NOR U844 ( .A(n737), .B(n738), .Z(n739) );
  XOR U845 ( .A(n2217), .B(n738), .Z(n740) );
  IV U846 ( .A(a[77]), .Z(n741) );
  NOR U847 ( .A(n740), .B(n741), .Z(n742) );
  NOR U848 ( .A(n739), .B(n742), .Z(n743) );
  IV U849 ( .A(n743), .Z(n2219) );
  IV U850 ( .A(n2225), .Z(n744) );
  IV U851 ( .A(b[80]), .Z(n745) );
  NOR U852 ( .A(n744), .B(n745), .Z(n746) );
  XOR U853 ( .A(n2225), .B(n745), .Z(n747) );
  IV U854 ( .A(a[80]), .Z(n748) );
  NOR U855 ( .A(n747), .B(n748), .Z(n749) );
  NOR U856 ( .A(n746), .B(n749), .Z(n750) );
  IV U857 ( .A(n750), .Z(n2227) );
  IV U858 ( .A(n2231), .Z(n751) );
  IV U859 ( .A(b[83]), .Z(n752) );
  NOR U860 ( .A(n751), .B(n752), .Z(n753) );
  XOR U861 ( .A(n2231), .B(n752), .Z(n754) );
  IV U862 ( .A(a[83]), .Z(n755) );
  NOR U863 ( .A(n754), .B(n755), .Z(n756) );
  NOR U864 ( .A(n753), .B(n756), .Z(n757) );
  IV U865 ( .A(n757), .Z(n2233) );
  IV U866 ( .A(n2237), .Z(n758) );
  IV U867 ( .A(b[86]), .Z(n759) );
  NOR U868 ( .A(n758), .B(n759), .Z(n760) );
  XOR U869 ( .A(n2237), .B(n759), .Z(n761) );
  IV U870 ( .A(a[86]), .Z(n762) );
  NOR U871 ( .A(n761), .B(n762), .Z(n763) );
  NOR U872 ( .A(n760), .B(n763), .Z(n764) );
  IV U873 ( .A(n764), .Z(n2239) );
  IV U874 ( .A(n2243), .Z(n765) );
  IV U875 ( .A(b[89]), .Z(n766) );
  NOR U876 ( .A(n765), .B(n766), .Z(n767) );
  XOR U877 ( .A(n2243), .B(n766), .Z(n768) );
  IV U878 ( .A(a[89]), .Z(n769) );
  NOR U879 ( .A(n768), .B(n769), .Z(n770) );
  NOR U880 ( .A(n767), .B(n770), .Z(n771) );
  IV U881 ( .A(n771), .Z(n2247) );
  IV U882 ( .A(n2251), .Z(n772) );
  IV U883 ( .A(b[92]), .Z(n773) );
  NOR U884 ( .A(n772), .B(n773), .Z(n774) );
  XOR U885 ( .A(n2251), .B(n773), .Z(n775) );
  IV U886 ( .A(a[92]), .Z(n776) );
  NOR U887 ( .A(n775), .B(n776), .Z(n777) );
  NOR U888 ( .A(n774), .B(n777), .Z(n778) );
  IV U889 ( .A(n778), .Z(n2253) );
  IV U890 ( .A(n2257), .Z(n779) );
  IV U891 ( .A(b[95]), .Z(n780) );
  NOR U892 ( .A(n779), .B(n780), .Z(n781) );
  XOR U893 ( .A(n2257), .B(n780), .Z(n782) );
  IV U894 ( .A(a[95]), .Z(n783) );
  NOR U895 ( .A(n782), .B(n783), .Z(n784) );
  NOR U896 ( .A(n781), .B(n784), .Z(n785) );
  IV U897 ( .A(n785), .Z(n2259) );
  IV U898 ( .A(n2263), .Z(n786) );
  IV U899 ( .A(b[98]), .Z(n787) );
  NOR U900 ( .A(n786), .B(n787), .Z(n788) );
  XOR U901 ( .A(n2263), .B(n787), .Z(n789) );
  IV U902 ( .A(a[98]), .Z(n790) );
  NOR U903 ( .A(n789), .B(n790), .Z(n791) );
  NOR U904 ( .A(n788), .B(n791), .Z(n792) );
  IV U905 ( .A(n792), .Z(n2265) );
  IV U906 ( .A(n1728), .Z(n793) );
  IV U907 ( .A(b[101]), .Z(n794) );
  NOR U908 ( .A(n793), .B(n794), .Z(n795) );
  XOR U909 ( .A(n1728), .B(n794), .Z(n796) );
  IV U910 ( .A(a[101]), .Z(n797) );
  NOR U911 ( .A(n796), .B(n797), .Z(n798) );
  NOR U912 ( .A(n795), .B(n798), .Z(n799) );
  IV U913 ( .A(n799), .Z(n1730) );
  IV U914 ( .A(n1734), .Z(n800) );
  IV U915 ( .A(b[104]), .Z(n801) );
  NOR U916 ( .A(n800), .B(n801), .Z(n802) );
  XOR U917 ( .A(n1734), .B(n801), .Z(n803) );
  IV U918 ( .A(a[104]), .Z(n804) );
  NOR U919 ( .A(n803), .B(n804), .Z(n805) );
  NOR U920 ( .A(n802), .B(n805), .Z(n806) );
  IV U921 ( .A(n806), .Z(n1736) );
  IV U922 ( .A(n1740), .Z(n807) );
  IV U923 ( .A(b[107]), .Z(n808) );
  NOR U924 ( .A(n807), .B(n808), .Z(n809) );
  XOR U925 ( .A(n1740), .B(n808), .Z(n810) );
  IV U926 ( .A(a[107]), .Z(n811) );
  NOR U927 ( .A(n810), .B(n811), .Z(n812) );
  NOR U928 ( .A(n809), .B(n812), .Z(n813) );
  IV U929 ( .A(n813), .Z(n1742) );
  IV U930 ( .A(n1748), .Z(n814) );
  IV U931 ( .A(b[110]), .Z(n815) );
  NOR U932 ( .A(n814), .B(n815), .Z(n816) );
  XOR U933 ( .A(n1748), .B(n815), .Z(n817) );
  IV U934 ( .A(a[110]), .Z(n818) );
  NOR U935 ( .A(n817), .B(n818), .Z(n819) );
  NOR U936 ( .A(n816), .B(n819), .Z(n820) );
  IV U937 ( .A(n820), .Z(n1750) );
  IV U938 ( .A(n1754), .Z(n821) );
  IV U939 ( .A(b[113]), .Z(n822) );
  NOR U940 ( .A(n821), .B(n822), .Z(n823) );
  XOR U941 ( .A(n1754), .B(n822), .Z(n824) );
  IV U942 ( .A(a[113]), .Z(n825) );
  NOR U943 ( .A(n824), .B(n825), .Z(n826) );
  NOR U944 ( .A(n823), .B(n826), .Z(n827) );
  IV U945 ( .A(n827), .Z(n1756) );
  IV U946 ( .A(n1760), .Z(n828) );
  IV U947 ( .A(b[116]), .Z(n829) );
  NOR U948 ( .A(n828), .B(n829), .Z(n830) );
  XOR U949 ( .A(n1760), .B(n829), .Z(n831) );
  IV U950 ( .A(a[116]), .Z(n832) );
  NOR U951 ( .A(n831), .B(n832), .Z(n833) );
  NOR U952 ( .A(n830), .B(n833), .Z(n834) );
  IV U953 ( .A(n834), .Z(n1762) );
  IV U954 ( .A(n1768), .Z(n835) );
  IV U955 ( .A(b[119]), .Z(n836) );
  NOR U956 ( .A(n835), .B(n836), .Z(n837) );
  XOR U957 ( .A(n1768), .B(n836), .Z(n838) );
  IV U958 ( .A(a[119]), .Z(n839) );
  NOR U959 ( .A(n838), .B(n839), .Z(n840) );
  NOR U960 ( .A(n837), .B(n840), .Z(n841) );
  IV U961 ( .A(n841), .Z(n1770) );
  IV U962 ( .A(n1774), .Z(n842) );
  IV U963 ( .A(b[122]), .Z(n843) );
  NOR U964 ( .A(n842), .B(n843), .Z(n844) );
  XOR U965 ( .A(n1774), .B(n843), .Z(n845) );
  IV U966 ( .A(a[122]), .Z(n846) );
  NOR U967 ( .A(n845), .B(n846), .Z(n847) );
  NOR U968 ( .A(n844), .B(n847), .Z(n848) );
  IV U969 ( .A(n848), .Z(n1776) );
  IV U970 ( .A(n1780), .Z(n849) );
  IV U971 ( .A(b[125]), .Z(n850) );
  NOR U972 ( .A(n849), .B(n850), .Z(n851) );
  XOR U973 ( .A(n1780), .B(n850), .Z(n852) );
  IV U974 ( .A(a[125]), .Z(n853) );
  NOR U975 ( .A(n852), .B(n853), .Z(n854) );
  NOR U976 ( .A(n851), .B(n854), .Z(n855) );
  IV U977 ( .A(n855), .Z(n1782) );
  IV U978 ( .A(n1786), .Z(n856) );
  IV U979 ( .A(b[128]), .Z(n857) );
  NOR U980 ( .A(n856), .B(n857), .Z(n858) );
  XOR U981 ( .A(n1786), .B(n857), .Z(n859) );
  IV U982 ( .A(a[128]), .Z(n860) );
  NOR U983 ( .A(n859), .B(n860), .Z(n861) );
  NOR U984 ( .A(n858), .B(n861), .Z(n862) );
  IV U985 ( .A(n862), .Z(n1790) );
  IV U986 ( .A(n1794), .Z(n863) );
  IV U987 ( .A(b[131]), .Z(n864) );
  NOR U988 ( .A(n863), .B(n864), .Z(n865) );
  XOR U989 ( .A(n1794), .B(n864), .Z(n866) );
  IV U990 ( .A(a[131]), .Z(n867) );
  NOR U991 ( .A(n866), .B(n867), .Z(n868) );
  NOR U992 ( .A(n865), .B(n868), .Z(n869) );
  IV U993 ( .A(n869), .Z(n1796) );
  IV U994 ( .A(n1800), .Z(n870) );
  IV U995 ( .A(b[134]), .Z(n871) );
  NOR U996 ( .A(n870), .B(n871), .Z(n872) );
  XOR U997 ( .A(n1800), .B(n871), .Z(n873) );
  IV U998 ( .A(a[134]), .Z(n874) );
  NOR U999 ( .A(n873), .B(n874), .Z(n875) );
  NOR U1000 ( .A(n872), .B(n875), .Z(n876) );
  IV U1001 ( .A(n876), .Z(n1802) );
  IV U1002 ( .A(n1806), .Z(n877) );
  IV U1003 ( .A(b[137]), .Z(n878) );
  NOR U1004 ( .A(n877), .B(n878), .Z(n879) );
  XOR U1005 ( .A(n1806), .B(n878), .Z(n880) );
  IV U1006 ( .A(a[137]), .Z(n881) );
  NOR U1007 ( .A(n880), .B(n881), .Z(n882) );
  NOR U1008 ( .A(n879), .B(n882), .Z(n883) );
  IV U1009 ( .A(n883), .Z(n1808) );
  IV U1010 ( .A(n1814), .Z(n884) );
  IV U1011 ( .A(b[140]), .Z(n885) );
  NOR U1012 ( .A(n884), .B(n885), .Z(n886) );
  XOR U1013 ( .A(n1814), .B(n885), .Z(n887) );
  IV U1014 ( .A(a[140]), .Z(n888) );
  NOR U1015 ( .A(n887), .B(n888), .Z(n889) );
  NOR U1016 ( .A(n886), .B(n889), .Z(n890) );
  IV U1017 ( .A(n890), .Z(n1816) );
  IV U1018 ( .A(n1820), .Z(n891) );
  IV U1019 ( .A(b[143]), .Z(n892) );
  NOR U1020 ( .A(n891), .B(n892), .Z(n893) );
  XOR U1021 ( .A(n1820), .B(n892), .Z(n894) );
  IV U1022 ( .A(a[143]), .Z(n895) );
  NOR U1023 ( .A(n894), .B(n895), .Z(n896) );
  NOR U1024 ( .A(n893), .B(n896), .Z(n897) );
  IV U1025 ( .A(n897), .Z(n1822) );
  IV U1026 ( .A(n1826), .Z(n898) );
  IV U1027 ( .A(b[146]), .Z(n899) );
  NOR U1028 ( .A(n898), .B(n899), .Z(n900) );
  XOR U1029 ( .A(n1826), .B(n899), .Z(n901) );
  IV U1030 ( .A(a[146]), .Z(n902) );
  NOR U1031 ( .A(n901), .B(n902), .Z(n903) );
  NOR U1032 ( .A(n900), .B(n903), .Z(n904) );
  IV U1033 ( .A(n904), .Z(n1828) );
  IV U1034 ( .A(n1834), .Z(n905) );
  IV U1035 ( .A(b[149]), .Z(n906) );
  NOR U1036 ( .A(n905), .B(n906), .Z(n907) );
  XOR U1037 ( .A(n1834), .B(n906), .Z(n908) );
  IV U1038 ( .A(a[149]), .Z(n909) );
  NOR U1039 ( .A(n908), .B(n909), .Z(n910) );
  NOR U1040 ( .A(n907), .B(n910), .Z(n911) );
  IV U1041 ( .A(n911), .Z(n1836) );
  IV U1042 ( .A(n1840), .Z(n912) );
  IV U1043 ( .A(b[152]), .Z(n913) );
  NOR U1044 ( .A(n912), .B(n913), .Z(n914) );
  XOR U1045 ( .A(n1840), .B(n913), .Z(n915) );
  IV U1046 ( .A(a[152]), .Z(n916) );
  NOR U1047 ( .A(n915), .B(n916), .Z(n917) );
  NOR U1048 ( .A(n914), .B(n917), .Z(n918) );
  IV U1049 ( .A(n918), .Z(n1842) );
  IV U1050 ( .A(n1846), .Z(n919) );
  IV U1051 ( .A(b[155]), .Z(n920) );
  NOR U1052 ( .A(n919), .B(n920), .Z(n921) );
  XOR U1053 ( .A(n1846), .B(n920), .Z(n922) );
  IV U1054 ( .A(a[155]), .Z(n923) );
  NOR U1055 ( .A(n922), .B(n923), .Z(n924) );
  NOR U1056 ( .A(n921), .B(n924), .Z(n925) );
  IV U1057 ( .A(n925), .Z(n1848) );
  IV U1058 ( .A(n1852), .Z(n926) );
  IV U1059 ( .A(b[158]), .Z(n927) );
  NOR U1060 ( .A(n926), .B(n927), .Z(n928) );
  XOR U1061 ( .A(n1852), .B(n927), .Z(n929) );
  IV U1062 ( .A(a[158]), .Z(n930) );
  NOR U1063 ( .A(n929), .B(n930), .Z(n931) );
  NOR U1064 ( .A(n928), .B(n931), .Z(n932) );
  IV U1065 ( .A(n932), .Z(n1856) );
  IV U1066 ( .A(n1860), .Z(n933) );
  IV U1067 ( .A(b[161]), .Z(n934) );
  NOR U1068 ( .A(n933), .B(n934), .Z(n935) );
  XOR U1069 ( .A(n1860), .B(n934), .Z(n936) );
  IV U1070 ( .A(a[161]), .Z(n937) );
  NOR U1071 ( .A(n936), .B(n937), .Z(n938) );
  NOR U1072 ( .A(n935), .B(n938), .Z(n939) );
  IV U1073 ( .A(n939), .Z(n1862) );
  IV U1074 ( .A(n1866), .Z(n940) );
  IV U1075 ( .A(b[164]), .Z(n941) );
  NOR U1076 ( .A(n940), .B(n941), .Z(n942) );
  XOR U1077 ( .A(n1866), .B(n941), .Z(n943) );
  IV U1078 ( .A(a[164]), .Z(n944) );
  NOR U1079 ( .A(n943), .B(n944), .Z(n945) );
  NOR U1080 ( .A(n942), .B(n945), .Z(n946) );
  IV U1081 ( .A(n946), .Z(n1868) );
  IV U1082 ( .A(n1872), .Z(n947) );
  IV U1083 ( .A(b[167]), .Z(n948) );
  NOR U1084 ( .A(n947), .B(n948), .Z(n949) );
  XOR U1085 ( .A(n1872), .B(n948), .Z(n950) );
  IV U1086 ( .A(a[167]), .Z(n951) );
  NOR U1087 ( .A(n950), .B(n951), .Z(n952) );
  NOR U1088 ( .A(n949), .B(n952), .Z(n953) );
  IV U1089 ( .A(n953), .Z(n1874) );
  IV U1090 ( .A(n1880), .Z(n954) );
  IV U1091 ( .A(b[170]), .Z(n955) );
  NOR U1092 ( .A(n954), .B(n955), .Z(n956) );
  XOR U1093 ( .A(n1880), .B(n955), .Z(n957) );
  IV U1094 ( .A(a[170]), .Z(n958) );
  NOR U1095 ( .A(n957), .B(n958), .Z(n959) );
  NOR U1096 ( .A(n956), .B(n959), .Z(n960) );
  IV U1097 ( .A(n960), .Z(n1882) );
  IV U1098 ( .A(n1886), .Z(n961) );
  IV U1099 ( .A(b[173]), .Z(n962) );
  NOR U1100 ( .A(n961), .B(n962), .Z(n963) );
  XOR U1101 ( .A(n1886), .B(n962), .Z(n964) );
  IV U1102 ( .A(a[173]), .Z(n965) );
  NOR U1103 ( .A(n964), .B(n965), .Z(n966) );
  NOR U1104 ( .A(n963), .B(n966), .Z(n967) );
  IV U1105 ( .A(n967), .Z(n1888) );
  IV U1106 ( .A(n1892), .Z(n968) );
  IV U1107 ( .A(b[176]), .Z(n969) );
  NOR U1108 ( .A(n968), .B(n969), .Z(n970) );
  XOR U1109 ( .A(n1892), .B(n969), .Z(n971) );
  IV U1110 ( .A(a[176]), .Z(n972) );
  NOR U1111 ( .A(n971), .B(n972), .Z(n973) );
  NOR U1112 ( .A(n970), .B(n973), .Z(n974) );
  IV U1113 ( .A(n974), .Z(n1894) );
  IV U1114 ( .A(n1900), .Z(n975) );
  IV U1115 ( .A(b[179]), .Z(n976) );
  NOR U1116 ( .A(n975), .B(n976), .Z(n977) );
  XOR U1117 ( .A(n1900), .B(n976), .Z(n978) );
  IV U1118 ( .A(a[179]), .Z(n979) );
  NOR U1119 ( .A(n978), .B(n979), .Z(n980) );
  NOR U1120 ( .A(n977), .B(n980), .Z(n981) );
  IV U1121 ( .A(n981), .Z(n1902) );
  IV U1122 ( .A(n1906), .Z(n982) );
  IV U1123 ( .A(b[182]), .Z(n983) );
  NOR U1124 ( .A(n982), .B(n983), .Z(n984) );
  XOR U1125 ( .A(n1906), .B(n983), .Z(n985) );
  IV U1126 ( .A(a[182]), .Z(n986) );
  NOR U1127 ( .A(n985), .B(n986), .Z(n987) );
  NOR U1128 ( .A(n984), .B(n987), .Z(n988) );
  IV U1129 ( .A(n988), .Z(n1908) );
  IV U1130 ( .A(n1912), .Z(n989) );
  IV U1131 ( .A(b[185]), .Z(n990) );
  NOR U1132 ( .A(n989), .B(n990), .Z(n991) );
  XOR U1133 ( .A(n1912), .B(n990), .Z(n992) );
  IV U1134 ( .A(a[185]), .Z(n993) );
  NOR U1135 ( .A(n992), .B(n993), .Z(n994) );
  NOR U1136 ( .A(n991), .B(n994), .Z(n995) );
  IV U1137 ( .A(n995), .Z(n1914) );
  IV U1138 ( .A(n1918), .Z(n996) );
  IV U1139 ( .A(b[188]), .Z(n997) );
  NOR U1140 ( .A(n996), .B(n997), .Z(n998) );
  XOR U1141 ( .A(n1918), .B(n997), .Z(n999) );
  IV U1142 ( .A(a[188]), .Z(n1000) );
  NOR U1143 ( .A(n999), .B(n1000), .Z(n1001) );
  NOR U1144 ( .A(n998), .B(n1001), .Z(n1002) );
  IV U1145 ( .A(n1002), .Z(n1922) );
  IV U1146 ( .A(n1926), .Z(n1003) );
  IV U1147 ( .A(b[191]), .Z(n1004) );
  NOR U1148 ( .A(n1003), .B(n1004), .Z(n1005) );
  XOR U1149 ( .A(n1926), .B(n1004), .Z(n1006) );
  IV U1150 ( .A(a[191]), .Z(n1007) );
  NOR U1151 ( .A(n1006), .B(n1007), .Z(n1008) );
  NOR U1152 ( .A(n1005), .B(n1008), .Z(n1009) );
  IV U1153 ( .A(n1009), .Z(n1928) );
  IV U1154 ( .A(n1932), .Z(n1010) );
  IV U1155 ( .A(b[194]), .Z(n1011) );
  NOR U1156 ( .A(n1010), .B(n1011), .Z(n1012) );
  XOR U1157 ( .A(n1932), .B(n1011), .Z(n1013) );
  IV U1158 ( .A(a[194]), .Z(n1014) );
  NOR U1159 ( .A(n1013), .B(n1014), .Z(n1015) );
  NOR U1160 ( .A(n1012), .B(n1015), .Z(n1016) );
  IV U1161 ( .A(n1016), .Z(n1934) );
  IV U1162 ( .A(n1938), .Z(n1017) );
  IV U1163 ( .A(b[197]), .Z(n1018) );
  NOR U1164 ( .A(n1017), .B(n1018), .Z(n1019) );
  XOR U1165 ( .A(n1938), .B(n1018), .Z(n1020) );
  IV U1166 ( .A(a[197]), .Z(n1021) );
  NOR U1167 ( .A(n1020), .B(n1021), .Z(n1022) );
  NOR U1168 ( .A(n1019), .B(n1022), .Z(n1023) );
  IV U1169 ( .A(n1023), .Z(n1940) );
  IV U1170 ( .A(n1948), .Z(n1024) );
  IV U1171 ( .A(b[200]), .Z(n1025) );
  NOR U1172 ( .A(n1024), .B(n1025), .Z(n1026) );
  XOR U1173 ( .A(n1948), .B(n1025), .Z(n1027) );
  IV U1174 ( .A(a[200]), .Z(n1028) );
  NOR U1175 ( .A(n1027), .B(n1028), .Z(n1029) );
  NOR U1176 ( .A(n1026), .B(n1029), .Z(n1030) );
  IV U1177 ( .A(n1030), .Z(n1950) );
  IV U1178 ( .A(n1954), .Z(n1031) );
  IV U1179 ( .A(b[203]), .Z(n1032) );
  NOR U1180 ( .A(n1031), .B(n1032), .Z(n1033) );
  XOR U1181 ( .A(n1954), .B(n1032), .Z(n1034) );
  IV U1182 ( .A(a[203]), .Z(n1035) );
  NOR U1183 ( .A(n1034), .B(n1035), .Z(n1036) );
  NOR U1184 ( .A(n1033), .B(n1036), .Z(n1037) );
  IV U1185 ( .A(n1037), .Z(n1956) );
  IV U1186 ( .A(n1960), .Z(n1038) );
  IV U1187 ( .A(b[206]), .Z(n1039) );
  NOR U1188 ( .A(n1038), .B(n1039), .Z(n1040) );
  XOR U1189 ( .A(n1960), .B(n1039), .Z(n1041) );
  IV U1190 ( .A(a[206]), .Z(n1042) );
  NOR U1191 ( .A(n1041), .B(n1042), .Z(n1043) );
  NOR U1192 ( .A(n1040), .B(n1043), .Z(n1044) );
  IV U1193 ( .A(n1044), .Z(n1962) );
  IV U1194 ( .A(n1968), .Z(n1045) );
  IV U1195 ( .A(b[209]), .Z(n1046) );
  NOR U1196 ( .A(n1045), .B(n1046), .Z(n1047) );
  XOR U1197 ( .A(n1968), .B(n1046), .Z(n1048) );
  IV U1198 ( .A(a[209]), .Z(n1049) );
  NOR U1199 ( .A(n1048), .B(n1049), .Z(n1050) );
  NOR U1200 ( .A(n1047), .B(n1050), .Z(n1051) );
  IV U1201 ( .A(n1051), .Z(n1970) );
  IV U1202 ( .A(n1974), .Z(n1052) );
  IV U1203 ( .A(b[212]), .Z(n1053) );
  NOR U1204 ( .A(n1052), .B(n1053), .Z(n1054) );
  XOR U1205 ( .A(n1974), .B(n1053), .Z(n1055) );
  IV U1206 ( .A(a[212]), .Z(n1056) );
  NOR U1207 ( .A(n1055), .B(n1056), .Z(n1057) );
  NOR U1208 ( .A(n1054), .B(n1057), .Z(n1058) );
  IV U1209 ( .A(n1058), .Z(n1976) );
  IV U1210 ( .A(n1980), .Z(n1059) );
  IV U1211 ( .A(b[215]), .Z(n1060) );
  NOR U1212 ( .A(n1059), .B(n1060), .Z(n1061) );
  XOR U1213 ( .A(n1980), .B(n1060), .Z(n1062) );
  IV U1214 ( .A(a[215]), .Z(n1063) );
  NOR U1215 ( .A(n1062), .B(n1063), .Z(n1064) );
  NOR U1216 ( .A(n1061), .B(n1064), .Z(n1065) );
  IV U1217 ( .A(n1065), .Z(n1982) );
  IV U1218 ( .A(n1986), .Z(n1066) );
  IV U1219 ( .A(b[218]), .Z(n1067) );
  NOR U1220 ( .A(n1066), .B(n1067), .Z(n1068) );
  XOR U1221 ( .A(n1986), .B(n1067), .Z(n1069) );
  IV U1222 ( .A(a[218]), .Z(n1070) );
  NOR U1223 ( .A(n1069), .B(n1070), .Z(n1071) );
  NOR U1224 ( .A(n1068), .B(n1071), .Z(n1072) );
  IV U1225 ( .A(n1072), .Z(n1990) );
  IV U1226 ( .A(n1994), .Z(n1073) );
  IV U1227 ( .A(b[221]), .Z(n1074) );
  NOR U1228 ( .A(n1073), .B(n1074), .Z(n1075) );
  XOR U1229 ( .A(n1994), .B(n1074), .Z(n1076) );
  IV U1230 ( .A(a[221]), .Z(n1077) );
  NOR U1231 ( .A(n1076), .B(n1077), .Z(n1078) );
  NOR U1232 ( .A(n1075), .B(n1078), .Z(n1079) );
  IV U1233 ( .A(n1079), .Z(n1996) );
  IV U1234 ( .A(n2000), .Z(n1080) );
  IV U1235 ( .A(b[224]), .Z(n1081) );
  NOR U1236 ( .A(n1080), .B(n1081), .Z(n1082) );
  XOR U1237 ( .A(n2000), .B(n1081), .Z(n1083) );
  IV U1238 ( .A(a[224]), .Z(n1084) );
  NOR U1239 ( .A(n1083), .B(n1084), .Z(n1085) );
  NOR U1240 ( .A(n1082), .B(n1085), .Z(n1086) );
  IV U1241 ( .A(n1086), .Z(n2002) );
  IV U1242 ( .A(n2006), .Z(n1087) );
  IV U1243 ( .A(b[227]), .Z(n1088) );
  NOR U1244 ( .A(n1087), .B(n1088), .Z(n1089) );
  XOR U1245 ( .A(n2006), .B(n1088), .Z(n1090) );
  IV U1246 ( .A(a[227]), .Z(n1091) );
  NOR U1247 ( .A(n1090), .B(n1091), .Z(n1092) );
  NOR U1248 ( .A(n1089), .B(n1092), .Z(n1093) );
  IV U1249 ( .A(n1093), .Z(n2008) );
  IV U1250 ( .A(n2014), .Z(n1094) );
  IV U1251 ( .A(b[230]), .Z(n1095) );
  NOR U1252 ( .A(n1094), .B(n1095), .Z(n1096) );
  XOR U1253 ( .A(n2014), .B(n1095), .Z(n1097) );
  IV U1254 ( .A(a[230]), .Z(n1098) );
  NOR U1255 ( .A(n1097), .B(n1098), .Z(n1099) );
  NOR U1256 ( .A(n1096), .B(n1099), .Z(n1100) );
  IV U1257 ( .A(n1100), .Z(n2016) );
  IV U1258 ( .A(n2020), .Z(n1101) );
  IV U1259 ( .A(b[233]), .Z(n1102) );
  NOR U1260 ( .A(n1101), .B(n1102), .Z(n1103) );
  XOR U1261 ( .A(n2020), .B(n1102), .Z(n1104) );
  IV U1262 ( .A(a[233]), .Z(n1105) );
  NOR U1263 ( .A(n1104), .B(n1105), .Z(n1106) );
  NOR U1264 ( .A(n1103), .B(n1106), .Z(n1107) );
  IV U1265 ( .A(n1107), .Z(n2022) );
  IV U1266 ( .A(n2026), .Z(n1108) );
  IV U1267 ( .A(b[236]), .Z(n1109) );
  NOR U1268 ( .A(n1108), .B(n1109), .Z(n1110) );
  XOR U1269 ( .A(n2026), .B(n1109), .Z(n1111) );
  IV U1270 ( .A(a[236]), .Z(n1112) );
  NOR U1271 ( .A(n1111), .B(n1112), .Z(n1113) );
  NOR U1272 ( .A(n1110), .B(n1113), .Z(n1114) );
  IV U1273 ( .A(n1114), .Z(n2028) );
  IV U1274 ( .A(n2034), .Z(n1115) );
  IV U1275 ( .A(b[239]), .Z(n1116) );
  NOR U1276 ( .A(n1115), .B(n1116), .Z(n1117) );
  XOR U1277 ( .A(n2034), .B(n1116), .Z(n1118) );
  IV U1278 ( .A(a[239]), .Z(n1119) );
  NOR U1279 ( .A(n1118), .B(n1119), .Z(n1120) );
  NOR U1280 ( .A(n1117), .B(n1120), .Z(n1121) );
  IV U1281 ( .A(n1121), .Z(n2036) );
  IV U1282 ( .A(n2040), .Z(n1122) );
  IV U1283 ( .A(b[242]), .Z(n1123) );
  NOR U1284 ( .A(n1122), .B(n1123), .Z(n1124) );
  XOR U1285 ( .A(n2040), .B(n1123), .Z(n1125) );
  IV U1286 ( .A(a[242]), .Z(n1126) );
  NOR U1287 ( .A(n1125), .B(n1126), .Z(n1127) );
  NOR U1288 ( .A(n1124), .B(n1127), .Z(n1128) );
  IV U1289 ( .A(n1128), .Z(n2042) );
  IV U1290 ( .A(n2046), .Z(n1129) );
  IV U1291 ( .A(b[245]), .Z(n1130) );
  NOR U1292 ( .A(n1129), .B(n1130), .Z(n1131) );
  XOR U1293 ( .A(n2046), .B(n1130), .Z(n1132) );
  IV U1294 ( .A(a[245]), .Z(n1133) );
  NOR U1295 ( .A(n1132), .B(n1133), .Z(n1134) );
  NOR U1296 ( .A(n1131), .B(n1134), .Z(n1135) );
  IV U1297 ( .A(n1135), .Z(n2048) );
  IV U1298 ( .A(n2135), .Z(n1136) );
  IV U1299 ( .A(b[3]), .Z(n1137) );
  NOR U1300 ( .A(n1136), .B(n1137), .Z(n1138) );
  XOR U1301 ( .A(n2135), .B(n1137), .Z(n1139) );
  IV U1302 ( .A(a[3]), .Z(n1140) );
  NOR U1303 ( .A(n1139), .B(n1140), .Z(n1141) );
  NOR U1304 ( .A(n1138), .B(n1141), .Z(n1142) );
  IV U1305 ( .A(n1142), .Z(n2157) );
  IV U1306 ( .A(n2201), .Z(n1143) );
  IV U1307 ( .A(b[6]), .Z(n1144) );
  NOR U1308 ( .A(n1143), .B(n1144), .Z(n1145) );
  XOR U1309 ( .A(n2201), .B(n1144), .Z(n1146) );
  IV U1310 ( .A(a[6]), .Z(n1147) );
  NOR U1311 ( .A(n1146), .B(n1147), .Z(n1148) );
  NOR U1312 ( .A(n1145), .B(n1148), .Z(n1149) );
  IV U1313 ( .A(n1149), .Z(n2223) );
  IV U1314 ( .A(n2267), .Z(n1150) );
  IV U1315 ( .A(a[9]), .Z(n1151) );
  NOR U1316 ( .A(n1150), .B(n1151), .Z(n1152) );
  XOR U1317 ( .A(n2267), .B(n1151), .Z(n1153) );
  IV U1318 ( .A(b[9]), .Z(n1154) );
  NOR U1319 ( .A(n1153), .B(n1154), .Z(n1155) );
  NOR U1320 ( .A(n1152), .B(n1155), .Z(n1156) );
  IV U1321 ( .A(n1156), .Z(n1744) );
  IV U1322 ( .A(n1788), .Z(n1157) );
  IV U1323 ( .A(b[12]), .Z(n1158) );
  NOR U1324 ( .A(n1157), .B(n1158), .Z(n1159) );
  XOR U1325 ( .A(n1788), .B(n1158), .Z(n1160) );
  IV U1326 ( .A(a[12]), .Z(n1161) );
  NOR U1327 ( .A(n1160), .B(n1161), .Z(n1162) );
  NOR U1328 ( .A(n1159), .B(n1162), .Z(n1163) );
  IV U1329 ( .A(n1163), .Z(n1810) );
  IV U1330 ( .A(n1854), .Z(n1164) );
  IV U1331 ( .A(b[15]), .Z(n1165) );
  NOR U1332 ( .A(n1164), .B(n1165), .Z(n1166) );
  XOR U1333 ( .A(n1854), .B(n1165), .Z(n1167) );
  IV U1334 ( .A(a[15]), .Z(n1168) );
  NOR U1335 ( .A(n1167), .B(n1168), .Z(n1169) );
  NOR U1336 ( .A(n1166), .B(n1169), .Z(n1170) );
  IV U1337 ( .A(n1170), .Z(n1876) );
  IV U1338 ( .A(n1920), .Z(n1171) );
  IV U1339 ( .A(b[18]), .Z(n1172) );
  NOR U1340 ( .A(n1171), .B(n1172), .Z(n1173) );
  XOR U1341 ( .A(n1920), .B(n1172), .Z(n1174) );
  IV U1342 ( .A(a[18]), .Z(n1175) );
  NOR U1343 ( .A(n1174), .B(n1175), .Z(n1176) );
  NOR U1344 ( .A(n1173), .B(n1176), .Z(n1177) );
  IV U1345 ( .A(n1177), .Z(n1942) );
  IV U1346 ( .A(n1988), .Z(n1178) );
  IV U1347 ( .A(b[21]), .Z(n1179) );
  NOR U1348 ( .A(n1178), .B(n1179), .Z(n1180) );
  XOR U1349 ( .A(n1988), .B(n1179), .Z(n1181) );
  IV U1350 ( .A(a[21]), .Z(n1182) );
  NOR U1351 ( .A(n1181), .B(n1182), .Z(n1183) );
  NOR U1352 ( .A(n1180), .B(n1183), .Z(n1184) );
  IV U1353 ( .A(n1184), .Z(n2010) );
  IV U1354 ( .A(n2063), .Z(n1185) );
  IV U1355 ( .A(b[24]), .Z(n1186) );
  NOR U1356 ( .A(n1185), .B(n1186), .Z(n1187) );
  XOR U1357 ( .A(n2063), .B(n1186), .Z(n1188) );
  IV U1358 ( .A(a[24]), .Z(n1189) );
  NOR U1359 ( .A(n1188), .B(n1189), .Z(n1190) );
  NOR U1360 ( .A(n1187), .B(n1190), .Z(n1191) );
  IV U1361 ( .A(n1191), .Z(n2102) );
  IV U1362 ( .A(n2106), .Z(n1192) );
  IV U1363 ( .A(b[27]), .Z(n1193) );
  NOR U1364 ( .A(n1192), .B(n1193), .Z(n1194) );
  XOR U1365 ( .A(n2106), .B(n1193), .Z(n1195) );
  IV U1366 ( .A(a[27]), .Z(n1196) );
  NOR U1367 ( .A(n1195), .B(n1196), .Z(n1197) );
  NOR U1368 ( .A(n1194), .B(n1197), .Z(n1198) );
  IV U1369 ( .A(n1198), .Z(n2108) );
  IV U1370 ( .A(n2115), .Z(n1199) );
  IV U1371 ( .A(b[30]), .Z(n1200) );
  NOR U1372 ( .A(n1199), .B(n1200), .Z(n1201) );
  XOR U1373 ( .A(n2115), .B(n1200), .Z(n1202) );
  IV U1374 ( .A(a[30]), .Z(n1203) );
  NOR U1375 ( .A(n1202), .B(n1203), .Z(n1204) );
  NOR U1376 ( .A(n1201), .B(n1204), .Z(n1205) );
  IV U1377 ( .A(n1205), .Z(n2117) );
  IV U1378 ( .A(n2121), .Z(n1206) );
  IV U1379 ( .A(b[33]), .Z(n1207) );
  NOR U1380 ( .A(n1206), .B(n1207), .Z(n1208) );
  XOR U1381 ( .A(n2121), .B(n1207), .Z(n1209) );
  IV U1382 ( .A(a[33]), .Z(n1210) );
  NOR U1383 ( .A(n1209), .B(n1210), .Z(n1211) );
  NOR U1384 ( .A(n1208), .B(n1211), .Z(n1212) );
  IV U1385 ( .A(n1212), .Z(n2123) );
  IV U1386 ( .A(n2127), .Z(n1213) );
  IV U1387 ( .A(b[36]), .Z(n1214) );
  NOR U1388 ( .A(n1213), .B(n1214), .Z(n1215) );
  XOR U1389 ( .A(n2127), .B(n1214), .Z(n1216) );
  IV U1390 ( .A(a[36]), .Z(n1217) );
  NOR U1391 ( .A(n1216), .B(n1217), .Z(n1218) );
  NOR U1392 ( .A(n1215), .B(n1218), .Z(n1219) );
  IV U1393 ( .A(n1219), .Z(n2129) );
  IV U1394 ( .A(n2133), .Z(n1220) );
  IV U1395 ( .A(b[39]), .Z(n1221) );
  NOR U1396 ( .A(n1220), .B(n1221), .Z(n1222) );
  XOR U1397 ( .A(n2133), .B(n1221), .Z(n1223) );
  IV U1398 ( .A(a[39]), .Z(n1224) );
  NOR U1399 ( .A(n1223), .B(n1224), .Z(n1225) );
  NOR U1400 ( .A(n1222), .B(n1225), .Z(n1226) );
  IV U1401 ( .A(n1226), .Z(n2137) );
  IV U1402 ( .A(n2141), .Z(n1227) );
  IV U1403 ( .A(b[42]), .Z(n1228) );
  NOR U1404 ( .A(n1227), .B(n1228), .Z(n1229) );
  XOR U1405 ( .A(n2141), .B(n1228), .Z(n1230) );
  IV U1406 ( .A(a[42]), .Z(n1231) );
  NOR U1407 ( .A(n1230), .B(n1231), .Z(n1232) );
  NOR U1408 ( .A(n1229), .B(n1232), .Z(n1233) );
  IV U1409 ( .A(n1233), .Z(n2143) );
  IV U1410 ( .A(n2147), .Z(n1234) );
  IV U1411 ( .A(b[45]), .Z(n1235) );
  NOR U1412 ( .A(n1234), .B(n1235), .Z(n1236) );
  XOR U1413 ( .A(n2147), .B(n1235), .Z(n1237) );
  IV U1414 ( .A(a[45]), .Z(n1238) );
  NOR U1415 ( .A(n1237), .B(n1238), .Z(n1239) );
  NOR U1416 ( .A(n1236), .B(n1239), .Z(n1240) );
  IV U1417 ( .A(n1240), .Z(n2149) );
  IV U1418 ( .A(n2153), .Z(n1241) );
  IV U1419 ( .A(b[48]), .Z(n1242) );
  NOR U1420 ( .A(n1241), .B(n1242), .Z(n1243) );
  XOR U1421 ( .A(n2153), .B(n1242), .Z(n1244) );
  IV U1422 ( .A(a[48]), .Z(n1245) );
  NOR U1423 ( .A(n1244), .B(n1245), .Z(n1246) );
  NOR U1424 ( .A(n1243), .B(n1246), .Z(n1247) );
  IV U1425 ( .A(n1247), .Z(n2155) );
  IV U1426 ( .A(n2161), .Z(n1248) );
  IV U1427 ( .A(b[51]), .Z(n1249) );
  NOR U1428 ( .A(n1248), .B(n1249), .Z(n1250) );
  XOR U1429 ( .A(n2161), .B(n1249), .Z(n1251) );
  IV U1430 ( .A(a[51]), .Z(n1252) );
  NOR U1431 ( .A(n1251), .B(n1252), .Z(n1253) );
  NOR U1432 ( .A(n1250), .B(n1253), .Z(n1254) );
  IV U1433 ( .A(n1254), .Z(n2163) );
  IV U1434 ( .A(n2167), .Z(n1255) );
  IV U1435 ( .A(b[54]), .Z(n1256) );
  NOR U1436 ( .A(n1255), .B(n1256), .Z(n1257) );
  XOR U1437 ( .A(n2167), .B(n1256), .Z(n1258) );
  IV U1438 ( .A(a[54]), .Z(n1259) );
  NOR U1439 ( .A(n1258), .B(n1259), .Z(n1260) );
  NOR U1440 ( .A(n1257), .B(n1260), .Z(n1261) );
  IV U1441 ( .A(n1261), .Z(n2169) );
  IV U1442 ( .A(n2173), .Z(n1262) );
  IV U1443 ( .A(b[57]), .Z(n1263) );
  NOR U1444 ( .A(n1262), .B(n1263), .Z(n1264) );
  XOR U1445 ( .A(n2173), .B(n1263), .Z(n1265) );
  IV U1446 ( .A(a[57]), .Z(n1266) );
  NOR U1447 ( .A(n1265), .B(n1266), .Z(n1267) );
  NOR U1448 ( .A(n1264), .B(n1267), .Z(n1268) );
  IV U1449 ( .A(n1268), .Z(n2175) );
  IV U1450 ( .A(n2181), .Z(n1269) );
  IV U1451 ( .A(b[60]), .Z(n1270) );
  NOR U1452 ( .A(n1269), .B(n1270), .Z(n1271) );
  XOR U1453 ( .A(n2181), .B(n1270), .Z(n1272) );
  IV U1454 ( .A(a[60]), .Z(n1273) );
  NOR U1455 ( .A(n1272), .B(n1273), .Z(n1274) );
  NOR U1456 ( .A(n1271), .B(n1274), .Z(n1275) );
  IV U1457 ( .A(n1275), .Z(n2183) );
  IV U1458 ( .A(n2187), .Z(n1276) );
  IV U1459 ( .A(b[63]), .Z(n1277) );
  NOR U1460 ( .A(n1276), .B(n1277), .Z(n1278) );
  XOR U1461 ( .A(n2187), .B(n1277), .Z(n1279) );
  IV U1462 ( .A(a[63]), .Z(n1280) );
  NOR U1463 ( .A(n1279), .B(n1280), .Z(n1281) );
  NOR U1464 ( .A(n1278), .B(n1281), .Z(n1282) );
  IV U1465 ( .A(n1282), .Z(n2189) );
  IV U1466 ( .A(n2193), .Z(n1283) );
  IV U1467 ( .A(b[66]), .Z(n1284) );
  NOR U1468 ( .A(n1283), .B(n1284), .Z(n1285) );
  XOR U1469 ( .A(n2193), .B(n1284), .Z(n1286) );
  IV U1470 ( .A(a[66]), .Z(n1287) );
  NOR U1471 ( .A(n1286), .B(n1287), .Z(n1288) );
  NOR U1472 ( .A(n1285), .B(n1288), .Z(n1289) );
  IV U1473 ( .A(n1289), .Z(n2195) );
  IV U1474 ( .A(n2199), .Z(n1290) );
  IV U1475 ( .A(b[69]), .Z(n1291) );
  NOR U1476 ( .A(n1290), .B(n1291), .Z(n1292) );
  XOR U1477 ( .A(n2199), .B(n1291), .Z(n1293) );
  IV U1478 ( .A(a[69]), .Z(n1294) );
  NOR U1479 ( .A(n1293), .B(n1294), .Z(n1295) );
  NOR U1480 ( .A(n1292), .B(n1295), .Z(n1296) );
  IV U1481 ( .A(n1296), .Z(n2203) );
  IV U1482 ( .A(n2207), .Z(n1297) );
  IV U1483 ( .A(b[72]), .Z(n1298) );
  NOR U1484 ( .A(n1297), .B(n1298), .Z(n1299) );
  XOR U1485 ( .A(n2207), .B(n1298), .Z(n1300) );
  IV U1486 ( .A(a[72]), .Z(n1301) );
  NOR U1487 ( .A(n1300), .B(n1301), .Z(n1302) );
  NOR U1488 ( .A(n1299), .B(n1302), .Z(n1303) );
  IV U1489 ( .A(n1303), .Z(n2209) );
  IV U1490 ( .A(n2213), .Z(n1304) );
  IV U1491 ( .A(b[75]), .Z(n1305) );
  NOR U1492 ( .A(n1304), .B(n1305), .Z(n1306) );
  XOR U1493 ( .A(n2213), .B(n1305), .Z(n1307) );
  IV U1494 ( .A(a[75]), .Z(n1308) );
  NOR U1495 ( .A(n1307), .B(n1308), .Z(n1309) );
  NOR U1496 ( .A(n1306), .B(n1309), .Z(n1310) );
  IV U1497 ( .A(n1310), .Z(n2215) );
  IV U1498 ( .A(n2219), .Z(n1311) );
  IV U1499 ( .A(b[78]), .Z(n1312) );
  NOR U1500 ( .A(n1311), .B(n1312), .Z(n1313) );
  XOR U1501 ( .A(n2219), .B(n1312), .Z(n1314) );
  IV U1502 ( .A(a[78]), .Z(n1315) );
  NOR U1503 ( .A(n1314), .B(n1315), .Z(n1316) );
  NOR U1504 ( .A(n1313), .B(n1316), .Z(n1317) );
  IV U1505 ( .A(n1317), .Z(n2221) );
  IV U1506 ( .A(n2227), .Z(n1318) );
  IV U1507 ( .A(b[81]), .Z(n1319) );
  NOR U1508 ( .A(n1318), .B(n1319), .Z(n1320) );
  XOR U1509 ( .A(n2227), .B(n1319), .Z(n1321) );
  IV U1510 ( .A(a[81]), .Z(n1322) );
  NOR U1511 ( .A(n1321), .B(n1322), .Z(n1323) );
  NOR U1512 ( .A(n1320), .B(n1323), .Z(n1324) );
  IV U1513 ( .A(n1324), .Z(n2229) );
  IV U1514 ( .A(n2233), .Z(n1325) );
  IV U1515 ( .A(b[84]), .Z(n1326) );
  NOR U1516 ( .A(n1325), .B(n1326), .Z(n1327) );
  XOR U1517 ( .A(n2233), .B(n1326), .Z(n1328) );
  IV U1518 ( .A(a[84]), .Z(n1329) );
  NOR U1519 ( .A(n1328), .B(n1329), .Z(n1330) );
  NOR U1520 ( .A(n1327), .B(n1330), .Z(n1331) );
  IV U1521 ( .A(n1331), .Z(n2235) );
  IV U1522 ( .A(n2239), .Z(n1332) );
  IV U1523 ( .A(b[87]), .Z(n1333) );
  NOR U1524 ( .A(n1332), .B(n1333), .Z(n1334) );
  XOR U1525 ( .A(n2239), .B(n1333), .Z(n1335) );
  IV U1526 ( .A(a[87]), .Z(n1336) );
  NOR U1527 ( .A(n1335), .B(n1336), .Z(n1337) );
  NOR U1528 ( .A(n1334), .B(n1337), .Z(n1338) );
  IV U1529 ( .A(n1338), .Z(n2241) );
  IV U1530 ( .A(n2247), .Z(n1339) );
  IV U1531 ( .A(b[90]), .Z(n1340) );
  NOR U1532 ( .A(n1339), .B(n1340), .Z(n1341) );
  XOR U1533 ( .A(n2247), .B(n1340), .Z(n1342) );
  IV U1534 ( .A(a[90]), .Z(n1343) );
  NOR U1535 ( .A(n1342), .B(n1343), .Z(n1344) );
  NOR U1536 ( .A(n1341), .B(n1344), .Z(n1345) );
  IV U1537 ( .A(n1345), .Z(n2249) );
  IV U1538 ( .A(n2253), .Z(n1346) );
  IV U1539 ( .A(b[93]), .Z(n1347) );
  NOR U1540 ( .A(n1346), .B(n1347), .Z(n1348) );
  XOR U1541 ( .A(n2253), .B(n1347), .Z(n1349) );
  IV U1542 ( .A(a[93]), .Z(n1350) );
  NOR U1543 ( .A(n1349), .B(n1350), .Z(n1351) );
  NOR U1544 ( .A(n1348), .B(n1351), .Z(n1352) );
  IV U1545 ( .A(n1352), .Z(n2255) );
  IV U1546 ( .A(n2259), .Z(n1353) );
  IV U1547 ( .A(b[96]), .Z(n1354) );
  NOR U1548 ( .A(n1353), .B(n1354), .Z(n1355) );
  XOR U1549 ( .A(n2259), .B(n1354), .Z(n1356) );
  IV U1550 ( .A(a[96]), .Z(n1357) );
  NOR U1551 ( .A(n1356), .B(n1357), .Z(n1358) );
  NOR U1552 ( .A(n1355), .B(n1358), .Z(n1359) );
  IV U1553 ( .A(n1359), .Z(n2261) );
  IV U1554 ( .A(n2265), .Z(n1360) );
  IV U1555 ( .A(a[99]), .Z(n1361) );
  NOR U1556 ( .A(n1360), .B(n1361), .Z(n1362) );
  XOR U1557 ( .A(n2265), .B(n1361), .Z(n1363) );
  IV U1558 ( .A(b[99]), .Z(n1364) );
  NOR U1559 ( .A(n1363), .B(n1364), .Z(n1365) );
  NOR U1560 ( .A(n1362), .B(n1365), .Z(n1366) );
  IV U1561 ( .A(n1366), .Z(n1726) );
  IV U1562 ( .A(n1730), .Z(n1367) );
  IV U1563 ( .A(b[102]), .Z(n1368) );
  NOR U1564 ( .A(n1367), .B(n1368), .Z(n1369) );
  XOR U1565 ( .A(n1730), .B(n1368), .Z(n1370) );
  IV U1566 ( .A(a[102]), .Z(n1371) );
  NOR U1567 ( .A(n1370), .B(n1371), .Z(n1372) );
  NOR U1568 ( .A(n1369), .B(n1372), .Z(n1373) );
  IV U1569 ( .A(n1373), .Z(n1732) );
  IV U1570 ( .A(n1736), .Z(n1374) );
  IV U1571 ( .A(b[105]), .Z(n1375) );
  NOR U1572 ( .A(n1374), .B(n1375), .Z(n1376) );
  XOR U1573 ( .A(n1736), .B(n1375), .Z(n1377) );
  IV U1574 ( .A(a[105]), .Z(n1378) );
  NOR U1575 ( .A(n1377), .B(n1378), .Z(n1379) );
  NOR U1576 ( .A(n1376), .B(n1379), .Z(n1380) );
  IV U1577 ( .A(n1380), .Z(n1738) );
  IV U1578 ( .A(n1742), .Z(n1381) );
  IV U1579 ( .A(b[108]), .Z(n1382) );
  NOR U1580 ( .A(n1381), .B(n1382), .Z(n1383) );
  XOR U1581 ( .A(n1742), .B(n1382), .Z(n1384) );
  IV U1582 ( .A(a[108]), .Z(n1385) );
  NOR U1583 ( .A(n1384), .B(n1385), .Z(n1386) );
  NOR U1584 ( .A(n1383), .B(n1386), .Z(n1387) );
  IV U1585 ( .A(n1387), .Z(n1746) );
  IV U1586 ( .A(n1750), .Z(n1388) );
  IV U1587 ( .A(b[111]), .Z(n1389) );
  NOR U1588 ( .A(n1388), .B(n1389), .Z(n1390) );
  XOR U1589 ( .A(n1750), .B(n1389), .Z(n1391) );
  IV U1590 ( .A(a[111]), .Z(n1392) );
  NOR U1591 ( .A(n1391), .B(n1392), .Z(n1393) );
  NOR U1592 ( .A(n1390), .B(n1393), .Z(n1394) );
  IV U1593 ( .A(n1394), .Z(n1752) );
  IV U1594 ( .A(n1756), .Z(n1395) );
  IV U1595 ( .A(b[114]), .Z(n1396) );
  NOR U1596 ( .A(n1395), .B(n1396), .Z(n1397) );
  XOR U1597 ( .A(n1756), .B(n1396), .Z(n1398) );
  IV U1598 ( .A(a[114]), .Z(n1399) );
  NOR U1599 ( .A(n1398), .B(n1399), .Z(n1400) );
  NOR U1600 ( .A(n1397), .B(n1400), .Z(n1401) );
  IV U1601 ( .A(n1401), .Z(n1758) );
  IV U1602 ( .A(n1762), .Z(n1402) );
  IV U1603 ( .A(b[117]), .Z(n1403) );
  NOR U1604 ( .A(n1402), .B(n1403), .Z(n1404) );
  XOR U1605 ( .A(n1762), .B(n1403), .Z(n1405) );
  IV U1606 ( .A(a[117]), .Z(n1406) );
  NOR U1607 ( .A(n1405), .B(n1406), .Z(n1407) );
  NOR U1608 ( .A(n1404), .B(n1407), .Z(n1408) );
  IV U1609 ( .A(n1408), .Z(n1764) );
  IV U1610 ( .A(n1770), .Z(n1409) );
  IV U1611 ( .A(b[120]), .Z(n1410) );
  NOR U1612 ( .A(n1409), .B(n1410), .Z(n1411) );
  XOR U1613 ( .A(n1770), .B(n1410), .Z(n1412) );
  IV U1614 ( .A(a[120]), .Z(n1413) );
  NOR U1615 ( .A(n1412), .B(n1413), .Z(n1414) );
  NOR U1616 ( .A(n1411), .B(n1414), .Z(n1415) );
  IV U1617 ( .A(n1415), .Z(n1772) );
  IV U1618 ( .A(n1776), .Z(n1416) );
  IV U1619 ( .A(b[123]), .Z(n1417) );
  NOR U1620 ( .A(n1416), .B(n1417), .Z(n1418) );
  XOR U1621 ( .A(n1776), .B(n1417), .Z(n1419) );
  IV U1622 ( .A(a[123]), .Z(n1420) );
  NOR U1623 ( .A(n1419), .B(n1420), .Z(n1421) );
  NOR U1624 ( .A(n1418), .B(n1421), .Z(n1422) );
  IV U1625 ( .A(n1422), .Z(n1778) );
  IV U1626 ( .A(n1782), .Z(n1423) );
  IV U1627 ( .A(b[126]), .Z(n1424) );
  NOR U1628 ( .A(n1423), .B(n1424), .Z(n1425) );
  XOR U1629 ( .A(n1782), .B(n1424), .Z(n1426) );
  IV U1630 ( .A(a[126]), .Z(n1427) );
  NOR U1631 ( .A(n1426), .B(n1427), .Z(n1428) );
  NOR U1632 ( .A(n1425), .B(n1428), .Z(n1429) );
  IV U1633 ( .A(n1429), .Z(n1784) );
  IV U1634 ( .A(n1790), .Z(n1430) );
  IV U1635 ( .A(b[129]), .Z(n1431) );
  NOR U1636 ( .A(n1430), .B(n1431), .Z(n1432) );
  XOR U1637 ( .A(n1790), .B(n1431), .Z(n1433) );
  IV U1638 ( .A(a[129]), .Z(n1434) );
  NOR U1639 ( .A(n1433), .B(n1434), .Z(n1435) );
  NOR U1640 ( .A(n1432), .B(n1435), .Z(n1436) );
  IV U1641 ( .A(n1436), .Z(n1792) );
  IV U1642 ( .A(n1796), .Z(n1437) );
  IV U1643 ( .A(b[132]), .Z(n1438) );
  NOR U1644 ( .A(n1437), .B(n1438), .Z(n1439) );
  XOR U1645 ( .A(n1796), .B(n1438), .Z(n1440) );
  IV U1646 ( .A(a[132]), .Z(n1441) );
  NOR U1647 ( .A(n1440), .B(n1441), .Z(n1442) );
  NOR U1648 ( .A(n1439), .B(n1442), .Z(n1443) );
  IV U1649 ( .A(n1443), .Z(n1798) );
  IV U1650 ( .A(n1802), .Z(n1444) );
  IV U1651 ( .A(b[135]), .Z(n1445) );
  NOR U1652 ( .A(n1444), .B(n1445), .Z(n1446) );
  XOR U1653 ( .A(n1802), .B(n1445), .Z(n1447) );
  IV U1654 ( .A(a[135]), .Z(n1448) );
  NOR U1655 ( .A(n1447), .B(n1448), .Z(n1449) );
  NOR U1656 ( .A(n1446), .B(n1449), .Z(n1450) );
  IV U1657 ( .A(n1450), .Z(n1804) );
  IV U1658 ( .A(n1808), .Z(n1451) );
  IV U1659 ( .A(b[138]), .Z(n1452) );
  NOR U1660 ( .A(n1451), .B(n1452), .Z(n1453) );
  XOR U1661 ( .A(n1808), .B(n1452), .Z(n1454) );
  IV U1662 ( .A(a[138]), .Z(n1455) );
  NOR U1663 ( .A(n1454), .B(n1455), .Z(n1456) );
  NOR U1664 ( .A(n1453), .B(n1456), .Z(n1457) );
  IV U1665 ( .A(n1457), .Z(n1812) );
  IV U1666 ( .A(n1816), .Z(n1458) );
  IV U1667 ( .A(b[141]), .Z(n1459) );
  NOR U1668 ( .A(n1458), .B(n1459), .Z(n1460) );
  XOR U1669 ( .A(n1816), .B(n1459), .Z(n1461) );
  IV U1670 ( .A(a[141]), .Z(n1462) );
  NOR U1671 ( .A(n1461), .B(n1462), .Z(n1463) );
  NOR U1672 ( .A(n1460), .B(n1463), .Z(n1464) );
  IV U1673 ( .A(n1464), .Z(n1818) );
  IV U1674 ( .A(n1822), .Z(n1465) );
  IV U1675 ( .A(b[144]), .Z(n1466) );
  NOR U1676 ( .A(n1465), .B(n1466), .Z(n1467) );
  XOR U1677 ( .A(n1822), .B(n1466), .Z(n1468) );
  IV U1678 ( .A(a[144]), .Z(n1469) );
  NOR U1679 ( .A(n1468), .B(n1469), .Z(n1470) );
  NOR U1680 ( .A(n1467), .B(n1470), .Z(n1471) );
  IV U1681 ( .A(n1471), .Z(n1824) );
  IV U1682 ( .A(n1828), .Z(n1472) );
  IV U1683 ( .A(b[147]), .Z(n1473) );
  NOR U1684 ( .A(n1472), .B(n1473), .Z(n1474) );
  XOR U1685 ( .A(n1828), .B(n1473), .Z(n1475) );
  IV U1686 ( .A(a[147]), .Z(n1476) );
  NOR U1687 ( .A(n1475), .B(n1476), .Z(n1477) );
  NOR U1688 ( .A(n1474), .B(n1477), .Z(n1478) );
  IV U1689 ( .A(n1478), .Z(n1830) );
  IV U1690 ( .A(n1836), .Z(n1479) );
  IV U1691 ( .A(b[150]), .Z(n1480) );
  NOR U1692 ( .A(n1479), .B(n1480), .Z(n1481) );
  XOR U1693 ( .A(n1836), .B(n1480), .Z(n1482) );
  IV U1694 ( .A(a[150]), .Z(n1483) );
  NOR U1695 ( .A(n1482), .B(n1483), .Z(n1484) );
  NOR U1696 ( .A(n1481), .B(n1484), .Z(n1485) );
  IV U1697 ( .A(n1485), .Z(n1838) );
  IV U1698 ( .A(n1842), .Z(n1486) );
  IV U1699 ( .A(b[153]), .Z(n1487) );
  NOR U1700 ( .A(n1486), .B(n1487), .Z(n1488) );
  XOR U1701 ( .A(n1842), .B(n1487), .Z(n1489) );
  IV U1702 ( .A(a[153]), .Z(n1490) );
  NOR U1703 ( .A(n1489), .B(n1490), .Z(n1491) );
  NOR U1704 ( .A(n1488), .B(n1491), .Z(n1492) );
  IV U1705 ( .A(n1492), .Z(n1844) );
  IV U1706 ( .A(n1848), .Z(n1493) );
  IV U1707 ( .A(b[156]), .Z(n1494) );
  NOR U1708 ( .A(n1493), .B(n1494), .Z(n1495) );
  XOR U1709 ( .A(n1848), .B(n1494), .Z(n1496) );
  IV U1710 ( .A(a[156]), .Z(n1497) );
  NOR U1711 ( .A(n1496), .B(n1497), .Z(n1498) );
  NOR U1712 ( .A(n1495), .B(n1498), .Z(n1499) );
  IV U1713 ( .A(n1499), .Z(n1850) );
  IV U1714 ( .A(n1856), .Z(n1500) );
  IV U1715 ( .A(b[159]), .Z(n1501) );
  NOR U1716 ( .A(n1500), .B(n1501), .Z(n1502) );
  XOR U1717 ( .A(n1856), .B(n1501), .Z(n1503) );
  IV U1718 ( .A(a[159]), .Z(n1504) );
  NOR U1719 ( .A(n1503), .B(n1504), .Z(n1505) );
  NOR U1720 ( .A(n1502), .B(n1505), .Z(n1506) );
  IV U1721 ( .A(n1506), .Z(n1858) );
  IV U1722 ( .A(n1862), .Z(n1507) );
  IV U1723 ( .A(b[162]), .Z(n1508) );
  NOR U1724 ( .A(n1507), .B(n1508), .Z(n1509) );
  XOR U1725 ( .A(n1862), .B(n1508), .Z(n1510) );
  IV U1726 ( .A(a[162]), .Z(n1511) );
  NOR U1727 ( .A(n1510), .B(n1511), .Z(n1512) );
  NOR U1728 ( .A(n1509), .B(n1512), .Z(n1513) );
  IV U1729 ( .A(n1513), .Z(n1864) );
  IV U1730 ( .A(n1868), .Z(n1514) );
  IV U1731 ( .A(b[165]), .Z(n1515) );
  NOR U1732 ( .A(n1514), .B(n1515), .Z(n1516) );
  XOR U1733 ( .A(n1868), .B(n1515), .Z(n1517) );
  IV U1734 ( .A(a[165]), .Z(n1518) );
  NOR U1735 ( .A(n1517), .B(n1518), .Z(n1519) );
  NOR U1736 ( .A(n1516), .B(n1519), .Z(n1520) );
  IV U1737 ( .A(n1520), .Z(n1870) );
  IV U1738 ( .A(n1874), .Z(n1521) );
  IV U1739 ( .A(b[168]), .Z(n1522) );
  NOR U1740 ( .A(n1521), .B(n1522), .Z(n1523) );
  XOR U1741 ( .A(n1874), .B(n1522), .Z(n1524) );
  IV U1742 ( .A(a[168]), .Z(n1525) );
  NOR U1743 ( .A(n1524), .B(n1525), .Z(n1526) );
  NOR U1744 ( .A(n1523), .B(n1526), .Z(n1527) );
  IV U1745 ( .A(n1527), .Z(n1878) );
  IV U1746 ( .A(n1882), .Z(n1528) );
  IV U1747 ( .A(b[171]), .Z(n1529) );
  NOR U1748 ( .A(n1528), .B(n1529), .Z(n1530) );
  XOR U1749 ( .A(n1882), .B(n1529), .Z(n1531) );
  IV U1750 ( .A(a[171]), .Z(n1532) );
  NOR U1751 ( .A(n1531), .B(n1532), .Z(n1533) );
  NOR U1752 ( .A(n1530), .B(n1533), .Z(n1534) );
  IV U1753 ( .A(n1534), .Z(n1884) );
  IV U1754 ( .A(n1888), .Z(n1535) );
  IV U1755 ( .A(b[174]), .Z(n1536) );
  NOR U1756 ( .A(n1535), .B(n1536), .Z(n1537) );
  XOR U1757 ( .A(n1888), .B(n1536), .Z(n1538) );
  IV U1758 ( .A(a[174]), .Z(n1539) );
  NOR U1759 ( .A(n1538), .B(n1539), .Z(n1540) );
  NOR U1760 ( .A(n1537), .B(n1540), .Z(n1541) );
  IV U1761 ( .A(n1541), .Z(n1890) );
  IV U1762 ( .A(n1894), .Z(n1542) );
  IV U1763 ( .A(b[177]), .Z(n1543) );
  NOR U1764 ( .A(n1542), .B(n1543), .Z(n1544) );
  XOR U1765 ( .A(n1894), .B(n1543), .Z(n1545) );
  IV U1766 ( .A(a[177]), .Z(n1546) );
  NOR U1767 ( .A(n1545), .B(n1546), .Z(n1547) );
  NOR U1768 ( .A(n1544), .B(n1547), .Z(n1548) );
  IV U1769 ( .A(n1548), .Z(n1896) );
  IV U1770 ( .A(n1902), .Z(n1549) );
  IV U1771 ( .A(b[180]), .Z(n1550) );
  NOR U1772 ( .A(n1549), .B(n1550), .Z(n1551) );
  XOR U1773 ( .A(n1902), .B(n1550), .Z(n1552) );
  IV U1774 ( .A(a[180]), .Z(n1553) );
  NOR U1775 ( .A(n1552), .B(n1553), .Z(n1554) );
  NOR U1776 ( .A(n1551), .B(n1554), .Z(n1555) );
  IV U1777 ( .A(n1555), .Z(n1904) );
  IV U1778 ( .A(n1908), .Z(n1556) );
  IV U1779 ( .A(b[183]), .Z(n1557) );
  NOR U1780 ( .A(n1556), .B(n1557), .Z(n1558) );
  XOR U1781 ( .A(n1908), .B(n1557), .Z(n1559) );
  IV U1782 ( .A(a[183]), .Z(n1560) );
  NOR U1783 ( .A(n1559), .B(n1560), .Z(n1561) );
  NOR U1784 ( .A(n1558), .B(n1561), .Z(n1562) );
  IV U1785 ( .A(n1562), .Z(n1910) );
  IV U1786 ( .A(n1914), .Z(n1563) );
  IV U1787 ( .A(b[186]), .Z(n1564) );
  NOR U1788 ( .A(n1563), .B(n1564), .Z(n1565) );
  XOR U1789 ( .A(n1914), .B(n1564), .Z(n1566) );
  IV U1790 ( .A(a[186]), .Z(n1567) );
  NOR U1791 ( .A(n1566), .B(n1567), .Z(n1568) );
  NOR U1792 ( .A(n1565), .B(n1568), .Z(n1569) );
  IV U1793 ( .A(n1569), .Z(n1916) );
  IV U1794 ( .A(n1922), .Z(n1570) );
  IV U1795 ( .A(b[189]), .Z(n1571) );
  NOR U1796 ( .A(n1570), .B(n1571), .Z(n1572) );
  XOR U1797 ( .A(n1922), .B(n1571), .Z(n1573) );
  IV U1798 ( .A(a[189]), .Z(n1574) );
  NOR U1799 ( .A(n1573), .B(n1574), .Z(n1575) );
  NOR U1800 ( .A(n1572), .B(n1575), .Z(n1576) );
  IV U1801 ( .A(n1576), .Z(n1924) );
  IV U1802 ( .A(n1928), .Z(n1577) );
  IV U1803 ( .A(b[192]), .Z(n1578) );
  NOR U1804 ( .A(n1577), .B(n1578), .Z(n1579) );
  XOR U1805 ( .A(n1928), .B(n1578), .Z(n1580) );
  IV U1806 ( .A(a[192]), .Z(n1581) );
  NOR U1807 ( .A(n1580), .B(n1581), .Z(n1582) );
  NOR U1808 ( .A(n1579), .B(n1582), .Z(n1583) );
  IV U1809 ( .A(n1583), .Z(n1930) );
  IV U1810 ( .A(n1934), .Z(n1584) );
  IV U1811 ( .A(b[195]), .Z(n1585) );
  NOR U1812 ( .A(n1584), .B(n1585), .Z(n1586) );
  XOR U1813 ( .A(n1934), .B(n1585), .Z(n1587) );
  IV U1814 ( .A(a[195]), .Z(n1588) );
  NOR U1815 ( .A(n1587), .B(n1588), .Z(n1589) );
  NOR U1816 ( .A(n1586), .B(n1589), .Z(n1590) );
  IV U1817 ( .A(n1590), .Z(n1936) );
  IV U1818 ( .A(n1940), .Z(n1591) );
  IV U1819 ( .A(b[198]), .Z(n1592) );
  NOR U1820 ( .A(n1591), .B(n1592), .Z(n1593) );
  XOR U1821 ( .A(n1940), .B(n1592), .Z(n1594) );
  IV U1822 ( .A(a[198]), .Z(n1595) );
  NOR U1823 ( .A(n1594), .B(n1595), .Z(n1596) );
  NOR U1824 ( .A(n1593), .B(n1596), .Z(n1597) );
  IV U1825 ( .A(n1597), .Z(n1946) );
  IV U1826 ( .A(n1950), .Z(n1598) );
  IV U1827 ( .A(b[201]), .Z(n1599) );
  NOR U1828 ( .A(n1598), .B(n1599), .Z(n1600) );
  XOR U1829 ( .A(n1950), .B(n1599), .Z(n1601) );
  IV U1830 ( .A(a[201]), .Z(n1602) );
  NOR U1831 ( .A(n1601), .B(n1602), .Z(n1603) );
  NOR U1832 ( .A(n1600), .B(n1603), .Z(n1604) );
  IV U1833 ( .A(n1604), .Z(n1952) );
  IV U1834 ( .A(n1956), .Z(n1605) );
  IV U1835 ( .A(b[204]), .Z(n1606) );
  NOR U1836 ( .A(n1605), .B(n1606), .Z(n1607) );
  XOR U1837 ( .A(n1956), .B(n1606), .Z(n1608) );
  IV U1838 ( .A(a[204]), .Z(n1609) );
  NOR U1839 ( .A(n1608), .B(n1609), .Z(n1610) );
  NOR U1840 ( .A(n1607), .B(n1610), .Z(n1611) );
  IV U1841 ( .A(n1611), .Z(n1958) );
  IV U1842 ( .A(n1962), .Z(n1612) );
  IV U1843 ( .A(b[207]), .Z(n1613) );
  NOR U1844 ( .A(n1612), .B(n1613), .Z(n1614) );
  XOR U1845 ( .A(n1962), .B(n1613), .Z(n1615) );
  IV U1846 ( .A(a[207]), .Z(n1616) );
  NOR U1847 ( .A(n1615), .B(n1616), .Z(n1617) );
  NOR U1848 ( .A(n1614), .B(n1617), .Z(n1618) );
  IV U1849 ( .A(n1618), .Z(n1964) );
  IV U1850 ( .A(n1970), .Z(n1619) );
  IV U1851 ( .A(b[210]), .Z(n1620) );
  NOR U1852 ( .A(n1619), .B(n1620), .Z(n1621) );
  XOR U1853 ( .A(n1970), .B(n1620), .Z(n1622) );
  IV U1854 ( .A(a[210]), .Z(n1623) );
  NOR U1855 ( .A(n1622), .B(n1623), .Z(n1624) );
  NOR U1856 ( .A(n1621), .B(n1624), .Z(n1625) );
  IV U1857 ( .A(n1625), .Z(n1972) );
  IV U1858 ( .A(n1976), .Z(n1626) );
  IV U1859 ( .A(b[213]), .Z(n1627) );
  NOR U1860 ( .A(n1626), .B(n1627), .Z(n1628) );
  XOR U1861 ( .A(n1976), .B(n1627), .Z(n1629) );
  IV U1862 ( .A(a[213]), .Z(n1630) );
  NOR U1863 ( .A(n1629), .B(n1630), .Z(n1631) );
  NOR U1864 ( .A(n1628), .B(n1631), .Z(n1632) );
  IV U1865 ( .A(n1632), .Z(n1978) );
  IV U1866 ( .A(n1982), .Z(n1633) );
  IV U1867 ( .A(b[216]), .Z(n1634) );
  NOR U1868 ( .A(n1633), .B(n1634), .Z(n1635) );
  XOR U1869 ( .A(n1982), .B(n1634), .Z(n1636) );
  IV U1870 ( .A(a[216]), .Z(n1637) );
  NOR U1871 ( .A(n1636), .B(n1637), .Z(n1638) );
  NOR U1872 ( .A(n1635), .B(n1638), .Z(n1639) );
  IV U1873 ( .A(n1639), .Z(n1984) );
  IV U1874 ( .A(n1990), .Z(n1640) );
  IV U1875 ( .A(b[219]), .Z(n1641) );
  NOR U1876 ( .A(n1640), .B(n1641), .Z(n1642) );
  XOR U1877 ( .A(n1990), .B(n1641), .Z(n1643) );
  IV U1878 ( .A(a[219]), .Z(n1644) );
  NOR U1879 ( .A(n1643), .B(n1644), .Z(n1645) );
  NOR U1880 ( .A(n1642), .B(n1645), .Z(n1646) );
  IV U1881 ( .A(n1646), .Z(n1992) );
  IV U1882 ( .A(n1996), .Z(n1647) );
  IV U1883 ( .A(b[222]), .Z(n1648) );
  NOR U1884 ( .A(n1647), .B(n1648), .Z(n1649) );
  XOR U1885 ( .A(n1996), .B(n1648), .Z(n1650) );
  IV U1886 ( .A(a[222]), .Z(n1651) );
  NOR U1887 ( .A(n1650), .B(n1651), .Z(n1652) );
  NOR U1888 ( .A(n1649), .B(n1652), .Z(n1653) );
  IV U1889 ( .A(n1653), .Z(n1998) );
  IV U1890 ( .A(n2002), .Z(n1654) );
  IV U1891 ( .A(b[225]), .Z(n1655) );
  NOR U1892 ( .A(n1654), .B(n1655), .Z(n1656) );
  XOR U1893 ( .A(n2002), .B(n1655), .Z(n1657) );
  IV U1894 ( .A(a[225]), .Z(n1658) );
  NOR U1895 ( .A(n1657), .B(n1658), .Z(n1659) );
  NOR U1896 ( .A(n1656), .B(n1659), .Z(n1660) );
  IV U1897 ( .A(n1660), .Z(n2004) );
  IV U1898 ( .A(n2008), .Z(n1661) );
  IV U1899 ( .A(b[228]), .Z(n1662) );
  NOR U1900 ( .A(n1661), .B(n1662), .Z(n1663) );
  XOR U1901 ( .A(n2008), .B(n1662), .Z(n1664) );
  IV U1902 ( .A(a[228]), .Z(n1665) );
  NOR U1903 ( .A(n1664), .B(n1665), .Z(n1666) );
  NOR U1904 ( .A(n1663), .B(n1666), .Z(n1667) );
  IV U1905 ( .A(n1667), .Z(n2012) );
  IV U1906 ( .A(n2016), .Z(n1668) );
  IV U1907 ( .A(b[231]), .Z(n1669) );
  NOR U1908 ( .A(n1668), .B(n1669), .Z(n1670) );
  XOR U1909 ( .A(n2016), .B(n1669), .Z(n1671) );
  IV U1910 ( .A(a[231]), .Z(n1672) );
  NOR U1911 ( .A(n1671), .B(n1672), .Z(n1673) );
  NOR U1912 ( .A(n1670), .B(n1673), .Z(n1674) );
  IV U1913 ( .A(n1674), .Z(n2018) );
  IV U1914 ( .A(n2022), .Z(n1675) );
  IV U1915 ( .A(b[234]), .Z(n1676) );
  NOR U1916 ( .A(n1675), .B(n1676), .Z(n1677) );
  XOR U1917 ( .A(n2022), .B(n1676), .Z(n1678) );
  IV U1918 ( .A(a[234]), .Z(n1679) );
  NOR U1919 ( .A(n1678), .B(n1679), .Z(n1680) );
  NOR U1920 ( .A(n1677), .B(n1680), .Z(n1681) );
  IV U1921 ( .A(n1681), .Z(n2024) );
  IV U1922 ( .A(n2028), .Z(n1682) );
  IV U1923 ( .A(b[237]), .Z(n1683) );
  NOR U1924 ( .A(n1682), .B(n1683), .Z(n1684) );
  XOR U1925 ( .A(n2028), .B(n1683), .Z(n1685) );
  IV U1926 ( .A(a[237]), .Z(n1686) );
  NOR U1927 ( .A(n1685), .B(n1686), .Z(n1687) );
  NOR U1928 ( .A(n1684), .B(n1687), .Z(n1688) );
  IV U1929 ( .A(n1688), .Z(n2030) );
  IV U1930 ( .A(n2036), .Z(n1689) );
  IV U1931 ( .A(b[240]), .Z(n1690) );
  NOR U1932 ( .A(n1689), .B(n1690), .Z(n1691) );
  XOR U1933 ( .A(n2036), .B(n1690), .Z(n1692) );
  IV U1934 ( .A(a[240]), .Z(n1693) );
  NOR U1935 ( .A(n1692), .B(n1693), .Z(n1694) );
  NOR U1936 ( .A(n1691), .B(n1694), .Z(n1695) );
  IV U1937 ( .A(n1695), .Z(n2038) );
  IV U1938 ( .A(n2042), .Z(n1696) );
  IV U1939 ( .A(b[243]), .Z(n1697) );
  NOR U1940 ( .A(n1696), .B(n1697), .Z(n1698) );
  XOR U1941 ( .A(n2042), .B(n1697), .Z(n1699) );
  IV U1942 ( .A(a[243]), .Z(n1700) );
  NOR U1943 ( .A(n1699), .B(n1700), .Z(n1701) );
  NOR U1944 ( .A(n1698), .B(n1701), .Z(n1702) );
  IV U1945 ( .A(n1702), .Z(n2044) );
  IV U1946 ( .A(b[246]), .Z(n1703) );
  IV U1947 ( .A(a[246]), .Z(n1704) );
  IV U1948 ( .A(n2048), .Z(n1705) );
  NOR U1949 ( .A(n1705), .B(n1703), .Z(n1706) );
  XOR U1950 ( .A(n2048), .B(n1703), .Z(n1707) );
  NOR U1951 ( .A(n1707), .B(n1704), .Z(n1708) );
  NOR U1952 ( .A(n1706), .B(n1708), .Z(n1709) );
  IV U1953 ( .A(n1709), .Z(n2050) );
  IV U1954 ( .A(a[255]), .Z(n1710) );
  NOR U1955 ( .A(a[255]), .B(n2270), .Z(n1711) );
  NOR U1956 ( .A(n2269), .B(n1710), .Z(n1712) );
  NOR U1957 ( .A(b[255]), .B(n1712), .Z(n1713) );
  NOR U1958 ( .A(n1711), .B(n1713), .Z(c[256]) );
  XOR U1959 ( .A(a[0]), .B(b[0]), .Z(c[0]) );
  IV U1960 ( .A(a[1]), .Z(n1714) );
  IV U1961 ( .A(b[1]), .Z(n1715) );
  NOR U1962 ( .A(n1714), .B(n1715), .Z(n1720) );
  XOR U1963 ( .A(a[1]), .B(n1715), .Z(n1945) );
  IV U1964 ( .A(a[0]), .Z(n1717) );
  IV U1965 ( .A(b[0]), .Z(n1716) );
  NOR U1966 ( .A(n1717), .B(n1716), .Z(n1718) );
  IV U1967 ( .A(n1718), .Z(n1944) );
  NOR U1968 ( .A(n1945), .B(n1944), .Z(n1719) );
  NOR U1969 ( .A(n1720), .B(n1719), .Z(n2112) );
  IV U1970 ( .A(n2112), .Z(n1721) );
  NOR U1971 ( .A(a[2]), .B(n1721), .Z(n1724) );
  IV U1972 ( .A(a[2]), .Z(n2114) );
  NOR U1973 ( .A(n2112), .B(n2114), .Z(n1722) );
  NOR U1974 ( .A(b[2]), .B(n1722), .Z(n1723) );
  NOR U1975 ( .A(n1724), .B(n1723), .Z(n2135) );
  XOR U1976 ( .A(b[100]), .B(n1726), .Z(n1725) );
  XOR U1977 ( .A(a[100]), .B(n1725), .Z(c[100]) );
  XOR U1978 ( .A(b[101]), .B(n1728), .Z(n1727) );
  XOR U1979 ( .A(a[101]), .B(n1727), .Z(c[101]) );
  XOR U1980 ( .A(b[102]), .B(n1730), .Z(n1729) );
  XOR U1981 ( .A(a[102]), .B(n1729), .Z(c[102]) );
  XOR U1982 ( .A(b[103]), .B(n1732), .Z(n1731) );
  XOR U1983 ( .A(a[103]), .B(n1731), .Z(c[103]) );
  XOR U1984 ( .A(b[104]), .B(n1734), .Z(n1733) );
  XOR U1985 ( .A(a[104]), .B(n1733), .Z(c[104]) );
  XOR U1986 ( .A(b[105]), .B(n1736), .Z(n1735) );
  XOR U1987 ( .A(a[105]), .B(n1735), .Z(c[105]) );
  XOR U1988 ( .A(b[106]), .B(n1738), .Z(n1737) );
  XOR U1989 ( .A(a[106]), .B(n1737), .Z(c[106]) );
  XOR U1990 ( .A(b[107]), .B(n1740), .Z(n1739) );
  XOR U1991 ( .A(a[107]), .B(n1739), .Z(c[107]) );
  XOR U1992 ( .A(b[108]), .B(n1742), .Z(n1741) );
  XOR U1993 ( .A(a[108]), .B(n1741), .Z(c[108]) );
  XOR U1994 ( .A(b[109]), .B(n1746), .Z(n1743) );
  XOR U1995 ( .A(a[109]), .B(n1743), .Z(c[109]) );
  XOR U1996 ( .A(b[10]), .B(n1744), .Z(n1745) );
  XOR U1997 ( .A(a[10]), .B(n1745), .Z(c[10]) );
  XOR U1998 ( .A(b[110]), .B(n1748), .Z(n1747) );
  XOR U1999 ( .A(a[110]), .B(n1747), .Z(c[110]) );
  XOR U2000 ( .A(b[111]), .B(n1750), .Z(n1749) );
  XOR U2001 ( .A(a[111]), .B(n1749), .Z(c[111]) );
  XOR U2002 ( .A(b[112]), .B(n1752), .Z(n1751) );
  XOR U2003 ( .A(a[112]), .B(n1751), .Z(c[112]) );
  XOR U2004 ( .A(b[113]), .B(n1754), .Z(n1753) );
  XOR U2005 ( .A(a[113]), .B(n1753), .Z(c[113]) );
  XOR U2006 ( .A(b[114]), .B(n1756), .Z(n1755) );
  XOR U2007 ( .A(a[114]), .B(n1755), .Z(c[114]) );
  XOR U2008 ( .A(b[115]), .B(n1758), .Z(n1757) );
  XOR U2009 ( .A(a[115]), .B(n1757), .Z(c[115]) );
  XOR U2010 ( .A(b[116]), .B(n1760), .Z(n1759) );
  XOR U2011 ( .A(a[116]), .B(n1759), .Z(c[116]) );
  XOR U2012 ( .A(b[117]), .B(n1762), .Z(n1761) );
  XOR U2013 ( .A(a[117]), .B(n1761), .Z(c[117]) );
  XOR U2014 ( .A(b[118]), .B(n1764), .Z(n1763) );
  XOR U2015 ( .A(a[118]), .B(n1763), .Z(c[118]) );
  XOR U2016 ( .A(b[119]), .B(n1768), .Z(n1765) );
  XOR U2017 ( .A(a[119]), .B(n1765), .Z(c[119]) );
  XOR U2018 ( .A(b[11]), .B(n1766), .Z(n1767) );
  XOR U2019 ( .A(a[11]), .B(n1767), .Z(c[11]) );
  XOR U2020 ( .A(b[120]), .B(n1770), .Z(n1769) );
  XOR U2021 ( .A(a[120]), .B(n1769), .Z(c[120]) );
  XOR U2022 ( .A(b[121]), .B(n1772), .Z(n1771) );
  XOR U2023 ( .A(a[121]), .B(n1771), .Z(c[121]) );
  XOR U2024 ( .A(b[122]), .B(n1774), .Z(n1773) );
  XOR U2025 ( .A(a[122]), .B(n1773), .Z(c[122]) );
  XOR U2026 ( .A(b[123]), .B(n1776), .Z(n1775) );
  XOR U2027 ( .A(a[123]), .B(n1775), .Z(c[123]) );
  XOR U2028 ( .A(b[124]), .B(n1778), .Z(n1777) );
  XOR U2029 ( .A(a[124]), .B(n1777), .Z(c[124]) );
  XOR U2030 ( .A(b[125]), .B(n1780), .Z(n1779) );
  XOR U2031 ( .A(a[125]), .B(n1779), .Z(c[125]) );
  XOR U2032 ( .A(b[126]), .B(n1782), .Z(n1781) );
  XOR U2033 ( .A(a[126]), .B(n1781), .Z(c[126]) );
  XOR U2034 ( .A(b[127]), .B(n1784), .Z(n1783) );
  XOR U2035 ( .A(a[127]), .B(n1783), .Z(c[127]) );
  XOR U2036 ( .A(b[128]), .B(n1786), .Z(n1785) );
  XOR U2037 ( .A(a[128]), .B(n1785), .Z(c[128]) );
  XOR U2038 ( .A(b[129]), .B(n1790), .Z(n1787) );
  XOR U2039 ( .A(a[129]), .B(n1787), .Z(c[129]) );
  XOR U2040 ( .A(b[12]), .B(n1788), .Z(n1789) );
  XOR U2041 ( .A(a[12]), .B(n1789), .Z(c[12]) );
  XOR U2042 ( .A(b[130]), .B(n1792), .Z(n1791) );
  XOR U2043 ( .A(a[130]), .B(n1791), .Z(c[130]) );
  XOR U2044 ( .A(b[131]), .B(n1794), .Z(n1793) );
  XOR U2045 ( .A(a[131]), .B(n1793), .Z(c[131]) );
  XOR U2046 ( .A(b[132]), .B(n1796), .Z(n1795) );
  XOR U2047 ( .A(a[132]), .B(n1795), .Z(c[132]) );
  XOR U2048 ( .A(b[133]), .B(n1798), .Z(n1797) );
  XOR U2049 ( .A(a[133]), .B(n1797), .Z(c[133]) );
  XOR U2050 ( .A(b[134]), .B(n1800), .Z(n1799) );
  XOR U2051 ( .A(a[134]), .B(n1799), .Z(c[134]) );
  XOR U2052 ( .A(b[135]), .B(n1802), .Z(n1801) );
  XOR U2053 ( .A(a[135]), .B(n1801), .Z(c[135]) );
  XOR U2054 ( .A(b[136]), .B(n1804), .Z(n1803) );
  XOR U2055 ( .A(a[136]), .B(n1803), .Z(c[136]) );
  XOR U2056 ( .A(b[137]), .B(n1806), .Z(n1805) );
  XOR U2057 ( .A(a[137]), .B(n1805), .Z(c[137]) );
  XOR U2058 ( .A(b[138]), .B(n1808), .Z(n1807) );
  XOR U2059 ( .A(a[138]), .B(n1807), .Z(c[138]) );
  XOR U2060 ( .A(b[139]), .B(n1812), .Z(n1809) );
  XOR U2061 ( .A(a[139]), .B(n1809), .Z(c[139]) );
  XOR U2062 ( .A(b[13]), .B(n1810), .Z(n1811) );
  XOR U2063 ( .A(a[13]), .B(n1811), .Z(c[13]) );
  XOR U2064 ( .A(b[140]), .B(n1814), .Z(n1813) );
  XOR U2065 ( .A(a[140]), .B(n1813), .Z(c[140]) );
  XOR U2066 ( .A(b[141]), .B(n1816), .Z(n1815) );
  XOR U2067 ( .A(a[141]), .B(n1815), .Z(c[141]) );
  XOR U2068 ( .A(b[142]), .B(n1818), .Z(n1817) );
  XOR U2069 ( .A(a[142]), .B(n1817), .Z(c[142]) );
  XOR U2070 ( .A(b[143]), .B(n1820), .Z(n1819) );
  XOR U2071 ( .A(a[143]), .B(n1819), .Z(c[143]) );
  XOR U2072 ( .A(b[144]), .B(n1822), .Z(n1821) );
  XOR U2073 ( .A(a[144]), .B(n1821), .Z(c[144]) );
  XOR U2074 ( .A(b[145]), .B(n1824), .Z(n1823) );
  XOR U2075 ( .A(a[145]), .B(n1823), .Z(c[145]) );
  XOR U2076 ( .A(b[146]), .B(n1826), .Z(n1825) );
  XOR U2077 ( .A(a[146]), .B(n1825), .Z(c[146]) );
  XOR U2078 ( .A(b[147]), .B(n1828), .Z(n1827) );
  XOR U2079 ( .A(a[147]), .B(n1827), .Z(c[147]) );
  XOR U2080 ( .A(b[148]), .B(n1830), .Z(n1829) );
  XOR U2081 ( .A(a[148]), .B(n1829), .Z(c[148]) );
  XOR U2082 ( .A(b[149]), .B(n1834), .Z(n1831) );
  XOR U2083 ( .A(a[149]), .B(n1831), .Z(c[149]) );
  XOR U2084 ( .A(b[14]), .B(n1832), .Z(n1833) );
  XOR U2085 ( .A(a[14]), .B(n1833), .Z(c[14]) );
  XOR U2086 ( .A(b[150]), .B(n1836), .Z(n1835) );
  XOR U2087 ( .A(a[150]), .B(n1835), .Z(c[150]) );
  XOR U2088 ( .A(b[151]), .B(n1838), .Z(n1837) );
  XOR U2089 ( .A(a[151]), .B(n1837), .Z(c[151]) );
  XOR U2090 ( .A(b[152]), .B(n1840), .Z(n1839) );
  XOR U2091 ( .A(a[152]), .B(n1839), .Z(c[152]) );
  XOR U2092 ( .A(b[153]), .B(n1842), .Z(n1841) );
  XOR U2093 ( .A(a[153]), .B(n1841), .Z(c[153]) );
  XOR U2094 ( .A(b[154]), .B(n1844), .Z(n1843) );
  XOR U2095 ( .A(a[154]), .B(n1843), .Z(c[154]) );
  XOR U2096 ( .A(b[155]), .B(n1846), .Z(n1845) );
  XOR U2097 ( .A(a[155]), .B(n1845), .Z(c[155]) );
  XOR U2098 ( .A(b[156]), .B(n1848), .Z(n1847) );
  XOR U2099 ( .A(a[156]), .B(n1847), .Z(c[156]) );
  XOR U2100 ( .A(b[157]), .B(n1850), .Z(n1849) );
  XOR U2101 ( .A(a[157]), .B(n1849), .Z(c[157]) );
  XOR U2102 ( .A(b[158]), .B(n1852), .Z(n1851) );
  XOR U2103 ( .A(a[158]), .B(n1851), .Z(c[158]) );
  XOR U2104 ( .A(b[159]), .B(n1856), .Z(n1853) );
  XOR U2105 ( .A(a[159]), .B(n1853), .Z(c[159]) );
  XOR U2106 ( .A(b[15]), .B(n1854), .Z(n1855) );
  XOR U2107 ( .A(a[15]), .B(n1855), .Z(c[15]) );
  XOR U2108 ( .A(b[160]), .B(n1858), .Z(n1857) );
  XOR U2109 ( .A(a[160]), .B(n1857), .Z(c[160]) );
  XOR U2110 ( .A(b[161]), .B(n1860), .Z(n1859) );
  XOR U2111 ( .A(a[161]), .B(n1859), .Z(c[161]) );
  XOR U2112 ( .A(b[162]), .B(n1862), .Z(n1861) );
  XOR U2113 ( .A(a[162]), .B(n1861), .Z(c[162]) );
  XOR U2114 ( .A(b[163]), .B(n1864), .Z(n1863) );
  XOR U2115 ( .A(a[163]), .B(n1863), .Z(c[163]) );
  XOR U2116 ( .A(b[164]), .B(n1866), .Z(n1865) );
  XOR U2117 ( .A(a[164]), .B(n1865), .Z(c[164]) );
  XOR U2118 ( .A(b[165]), .B(n1868), .Z(n1867) );
  XOR U2119 ( .A(a[165]), .B(n1867), .Z(c[165]) );
  XOR U2120 ( .A(b[166]), .B(n1870), .Z(n1869) );
  XOR U2121 ( .A(a[166]), .B(n1869), .Z(c[166]) );
  XOR U2122 ( .A(b[167]), .B(n1872), .Z(n1871) );
  XOR U2123 ( .A(a[167]), .B(n1871), .Z(c[167]) );
  XOR U2124 ( .A(b[168]), .B(n1874), .Z(n1873) );
  XOR U2125 ( .A(a[168]), .B(n1873), .Z(c[168]) );
  XOR U2126 ( .A(b[169]), .B(n1878), .Z(n1875) );
  XOR U2127 ( .A(a[169]), .B(n1875), .Z(c[169]) );
  XOR U2128 ( .A(b[16]), .B(n1876), .Z(n1877) );
  XOR U2129 ( .A(a[16]), .B(n1877), .Z(c[16]) );
  XOR U2130 ( .A(b[170]), .B(n1880), .Z(n1879) );
  XOR U2131 ( .A(a[170]), .B(n1879), .Z(c[170]) );
  XOR U2132 ( .A(b[171]), .B(n1882), .Z(n1881) );
  XOR U2133 ( .A(a[171]), .B(n1881), .Z(c[171]) );
  XOR U2134 ( .A(b[172]), .B(n1884), .Z(n1883) );
  XOR U2135 ( .A(a[172]), .B(n1883), .Z(c[172]) );
  XOR U2136 ( .A(b[173]), .B(n1886), .Z(n1885) );
  XOR U2137 ( .A(a[173]), .B(n1885), .Z(c[173]) );
  XOR U2138 ( .A(b[174]), .B(n1888), .Z(n1887) );
  XOR U2139 ( .A(a[174]), .B(n1887), .Z(c[174]) );
  XOR U2140 ( .A(b[175]), .B(n1890), .Z(n1889) );
  XOR U2141 ( .A(a[175]), .B(n1889), .Z(c[175]) );
  XOR U2142 ( .A(b[176]), .B(n1892), .Z(n1891) );
  XOR U2143 ( .A(a[176]), .B(n1891), .Z(c[176]) );
  XOR U2144 ( .A(b[177]), .B(n1894), .Z(n1893) );
  XOR U2145 ( .A(a[177]), .B(n1893), .Z(c[177]) );
  XOR U2146 ( .A(b[178]), .B(n1896), .Z(n1895) );
  XOR U2147 ( .A(a[178]), .B(n1895), .Z(c[178]) );
  XOR U2148 ( .A(b[179]), .B(n1900), .Z(n1897) );
  XOR U2149 ( .A(a[179]), .B(n1897), .Z(c[179]) );
  XOR U2150 ( .A(b[17]), .B(n1898), .Z(n1899) );
  XOR U2151 ( .A(a[17]), .B(n1899), .Z(c[17]) );
  XOR U2152 ( .A(b[180]), .B(n1902), .Z(n1901) );
  XOR U2153 ( .A(a[180]), .B(n1901), .Z(c[180]) );
  XOR U2154 ( .A(b[181]), .B(n1904), .Z(n1903) );
  XOR U2155 ( .A(a[181]), .B(n1903), .Z(c[181]) );
  XOR U2156 ( .A(b[182]), .B(n1906), .Z(n1905) );
  XOR U2157 ( .A(a[182]), .B(n1905), .Z(c[182]) );
  XOR U2158 ( .A(b[183]), .B(n1908), .Z(n1907) );
  XOR U2159 ( .A(a[183]), .B(n1907), .Z(c[183]) );
  XOR U2160 ( .A(b[184]), .B(n1910), .Z(n1909) );
  XOR U2161 ( .A(a[184]), .B(n1909), .Z(c[184]) );
  XOR U2162 ( .A(b[185]), .B(n1912), .Z(n1911) );
  XOR U2163 ( .A(a[185]), .B(n1911), .Z(c[185]) );
  XOR U2164 ( .A(b[186]), .B(n1914), .Z(n1913) );
  XOR U2165 ( .A(a[186]), .B(n1913), .Z(c[186]) );
  XOR U2166 ( .A(b[187]), .B(n1916), .Z(n1915) );
  XOR U2167 ( .A(a[187]), .B(n1915), .Z(c[187]) );
  XOR U2168 ( .A(b[188]), .B(n1918), .Z(n1917) );
  XOR U2169 ( .A(a[188]), .B(n1917), .Z(c[188]) );
  XOR U2170 ( .A(b[189]), .B(n1922), .Z(n1919) );
  XOR U2171 ( .A(a[189]), .B(n1919), .Z(c[189]) );
  XOR U2172 ( .A(b[18]), .B(n1920), .Z(n1921) );
  XOR U2173 ( .A(a[18]), .B(n1921), .Z(c[18]) );
  XOR U2174 ( .A(b[190]), .B(n1924), .Z(n1923) );
  XOR U2175 ( .A(a[190]), .B(n1923), .Z(c[190]) );
  XOR U2176 ( .A(b[191]), .B(n1926), .Z(n1925) );
  XOR U2177 ( .A(a[191]), .B(n1925), .Z(c[191]) );
  XOR U2178 ( .A(b[192]), .B(n1928), .Z(n1927) );
  XOR U2179 ( .A(a[192]), .B(n1927), .Z(c[192]) );
  XOR U2180 ( .A(b[193]), .B(n1930), .Z(n1929) );
  XOR U2181 ( .A(a[193]), .B(n1929), .Z(c[193]) );
  XOR U2182 ( .A(b[194]), .B(n1932), .Z(n1931) );
  XOR U2183 ( .A(a[194]), .B(n1931), .Z(c[194]) );
  XOR U2184 ( .A(b[195]), .B(n1934), .Z(n1933) );
  XOR U2185 ( .A(a[195]), .B(n1933), .Z(c[195]) );
  XOR U2186 ( .A(b[196]), .B(n1936), .Z(n1935) );
  XOR U2187 ( .A(a[196]), .B(n1935), .Z(c[196]) );
  XOR U2188 ( .A(b[197]), .B(n1938), .Z(n1937) );
  XOR U2189 ( .A(a[197]), .B(n1937), .Z(c[197]) );
  XOR U2190 ( .A(b[198]), .B(n1940), .Z(n1939) );
  XOR U2191 ( .A(a[198]), .B(n1939), .Z(c[198]) );
  XOR U2192 ( .A(b[199]), .B(n1946), .Z(n1941) );
  XOR U2193 ( .A(a[199]), .B(n1941), .Z(c[199]) );
  XOR U2194 ( .A(b[19]), .B(n1942), .Z(n1943) );
  XOR U2195 ( .A(a[19]), .B(n1943), .Z(c[19]) );
  XOR U2196 ( .A(n1945), .B(n1944), .Z(c[1]) );
  XOR U2197 ( .A(b[200]), .B(n1948), .Z(n1947) );
  XOR U2198 ( .A(a[200]), .B(n1947), .Z(c[200]) );
  XOR U2199 ( .A(b[201]), .B(n1950), .Z(n1949) );
  XOR U2200 ( .A(a[201]), .B(n1949), .Z(c[201]) );
  XOR U2201 ( .A(b[202]), .B(n1952), .Z(n1951) );
  XOR U2202 ( .A(a[202]), .B(n1951), .Z(c[202]) );
  XOR U2203 ( .A(b[203]), .B(n1954), .Z(n1953) );
  XOR U2204 ( .A(a[203]), .B(n1953), .Z(c[203]) );
  XOR U2205 ( .A(b[204]), .B(n1956), .Z(n1955) );
  XOR U2206 ( .A(a[204]), .B(n1955), .Z(c[204]) );
  XOR U2207 ( .A(b[205]), .B(n1958), .Z(n1957) );
  XOR U2208 ( .A(a[205]), .B(n1957), .Z(c[205]) );
  XOR U2209 ( .A(b[206]), .B(n1960), .Z(n1959) );
  XOR U2210 ( .A(a[206]), .B(n1959), .Z(c[206]) );
  XOR U2211 ( .A(b[207]), .B(n1962), .Z(n1961) );
  XOR U2212 ( .A(a[207]), .B(n1961), .Z(c[207]) );
  XOR U2213 ( .A(b[208]), .B(n1964), .Z(n1963) );
  XOR U2214 ( .A(a[208]), .B(n1963), .Z(c[208]) );
  XOR U2215 ( .A(b[209]), .B(n1968), .Z(n1965) );
  XOR U2216 ( .A(a[209]), .B(n1965), .Z(c[209]) );
  XOR U2217 ( .A(b[20]), .B(n1966), .Z(n1967) );
  XOR U2218 ( .A(a[20]), .B(n1967), .Z(c[20]) );
  XOR U2219 ( .A(b[210]), .B(n1970), .Z(n1969) );
  XOR U2220 ( .A(a[210]), .B(n1969), .Z(c[210]) );
  XOR U2221 ( .A(b[211]), .B(n1972), .Z(n1971) );
  XOR U2222 ( .A(a[211]), .B(n1971), .Z(c[211]) );
  XOR U2223 ( .A(b[212]), .B(n1974), .Z(n1973) );
  XOR U2224 ( .A(a[212]), .B(n1973), .Z(c[212]) );
  XOR U2225 ( .A(b[213]), .B(n1976), .Z(n1975) );
  XOR U2226 ( .A(a[213]), .B(n1975), .Z(c[213]) );
  XOR U2227 ( .A(b[214]), .B(n1978), .Z(n1977) );
  XOR U2228 ( .A(a[214]), .B(n1977), .Z(c[214]) );
  XOR U2229 ( .A(b[215]), .B(n1980), .Z(n1979) );
  XOR U2230 ( .A(a[215]), .B(n1979), .Z(c[215]) );
  XOR U2231 ( .A(b[216]), .B(n1982), .Z(n1981) );
  XOR U2232 ( .A(a[216]), .B(n1981), .Z(c[216]) );
  XOR U2233 ( .A(b[217]), .B(n1984), .Z(n1983) );
  XOR U2234 ( .A(a[217]), .B(n1983), .Z(c[217]) );
  XOR U2235 ( .A(b[218]), .B(n1986), .Z(n1985) );
  XOR U2236 ( .A(a[218]), .B(n1985), .Z(c[218]) );
  XOR U2237 ( .A(b[219]), .B(n1990), .Z(n1987) );
  XOR U2238 ( .A(a[219]), .B(n1987), .Z(c[219]) );
  XOR U2239 ( .A(b[21]), .B(n1988), .Z(n1989) );
  XOR U2240 ( .A(a[21]), .B(n1989), .Z(c[21]) );
  XOR U2241 ( .A(b[220]), .B(n1992), .Z(n1991) );
  XOR U2242 ( .A(a[220]), .B(n1991), .Z(c[220]) );
  XOR U2243 ( .A(b[221]), .B(n1994), .Z(n1993) );
  XOR U2244 ( .A(a[221]), .B(n1993), .Z(c[221]) );
  XOR U2245 ( .A(b[222]), .B(n1996), .Z(n1995) );
  XOR U2246 ( .A(a[222]), .B(n1995), .Z(c[222]) );
  XOR U2247 ( .A(b[223]), .B(n1998), .Z(n1997) );
  XOR U2248 ( .A(a[223]), .B(n1997), .Z(c[223]) );
  XOR U2249 ( .A(b[224]), .B(n2000), .Z(n1999) );
  XOR U2250 ( .A(a[224]), .B(n1999), .Z(c[224]) );
  XOR U2251 ( .A(b[225]), .B(n2002), .Z(n2001) );
  XOR U2252 ( .A(a[225]), .B(n2001), .Z(c[225]) );
  XOR U2253 ( .A(b[226]), .B(n2004), .Z(n2003) );
  XOR U2254 ( .A(a[226]), .B(n2003), .Z(c[226]) );
  XOR U2255 ( .A(b[227]), .B(n2006), .Z(n2005) );
  XOR U2256 ( .A(a[227]), .B(n2005), .Z(c[227]) );
  XOR U2257 ( .A(b[228]), .B(n2008), .Z(n2007) );
  XOR U2258 ( .A(a[228]), .B(n2007), .Z(c[228]) );
  XOR U2259 ( .A(b[229]), .B(n2012), .Z(n2009) );
  XOR U2260 ( .A(a[229]), .B(n2009), .Z(c[229]) );
  XOR U2261 ( .A(b[22]), .B(n2010), .Z(n2011) );
  XOR U2262 ( .A(a[22]), .B(n2011), .Z(c[22]) );
  XOR U2263 ( .A(b[230]), .B(n2014), .Z(n2013) );
  XOR U2264 ( .A(a[230]), .B(n2013), .Z(c[230]) );
  XOR U2265 ( .A(b[231]), .B(n2016), .Z(n2015) );
  XOR U2266 ( .A(a[231]), .B(n2015), .Z(c[231]) );
  XOR U2267 ( .A(b[232]), .B(n2018), .Z(n2017) );
  XOR U2268 ( .A(a[232]), .B(n2017), .Z(c[232]) );
  XOR U2269 ( .A(b[233]), .B(n2020), .Z(n2019) );
  XOR U2270 ( .A(a[233]), .B(n2019), .Z(c[233]) );
  XOR U2271 ( .A(b[234]), .B(n2022), .Z(n2021) );
  XOR U2272 ( .A(a[234]), .B(n2021), .Z(c[234]) );
  XOR U2273 ( .A(b[235]), .B(n2024), .Z(n2023) );
  XOR U2274 ( .A(a[235]), .B(n2023), .Z(c[235]) );
  XOR U2275 ( .A(b[236]), .B(n2026), .Z(n2025) );
  XOR U2276 ( .A(a[236]), .B(n2025), .Z(c[236]) );
  XOR U2277 ( .A(b[237]), .B(n2028), .Z(n2027) );
  XOR U2278 ( .A(a[237]), .B(n2027), .Z(c[237]) );
  XOR U2279 ( .A(b[238]), .B(n2030), .Z(n2029) );
  XOR U2280 ( .A(a[238]), .B(n2029), .Z(c[238]) );
  XOR U2281 ( .A(b[239]), .B(n2034), .Z(n2031) );
  XOR U2282 ( .A(a[239]), .B(n2031), .Z(c[239]) );
  XOR U2283 ( .A(b[23]), .B(n2032), .Z(n2033) );
  XOR U2284 ( .A(a[23]), .B(n2033), .Z(c[23]) );
  XOR U2285 ( .A(b[240]), .B(n2036), .Z(n2035) );
  XOR U2286 ( .A(a[240]), .B(n2035), .Z(c[240]) );
  XOR U2287 ( .A(b[241]), .B(n2038), .Z(n2037) );
  XOR U2288 ( .A(a[241]), .B(n2037), .Z(c[241]) );
  XOR U2289 ( .A(b[242]), .B(n2040), .Z(n2039) );
  XOR U2290 ( .A(a[242]), .B(n2039), .Z(c[242]) );
  XOR U2291 ( .A(b[243]), .B(n2042), .Z(n2041) );
  XOR U2292 ( .A(a[243]), .B(n2041), .Z(c[243]) );
  XOR U2293 ( .A(b[244]), .B(n2044), .Z(n2043) );
  XOR U2294 ( .A(a[244]), .B(n2043), .Z(c[244]) );
  XOR U2295 ( .A(b[245]), .B(n2046), .Z(n2045) );
  XOR U2296 ( .A(a[245]), .B(n2045), .Z(c[245]) );
  XOR U2297 ( .A(b[246]), .B(n2048), .Z(n2047) );
  XOR U2298 ( .A(a[246]), .B(n2047), .Z(c[246]) );
  XOR U2299 ( .A(b[247]), .B(n2050), .Z(n2049) );
  XOR U2300 ( .A(a[247]), .B(n2049), .Z(c[247]) );
  IV U2301 ( .A(a[248]), .Z(n2057) );
  IV U2302 ( .A(n2050), .Z(n2053) );
  XOR U2303 ( .A(b[247]), .B(n2053), .Z(n2052) );
  IV U2304 ( .A(a[247]), .Z(n2051) );
  NOR U2305 ( .A(n2052), .B(n2051), .Z(n2056) );
  IV U2306 ( .A(b[247]), .Z(n2054) );
  NOR U2307 ( .A(n2054), .B(n2053), .Z(n2055) );
  NOR U2308 ( .A(n2056), .B(n2055), .Z(n2059) );
  XOR U2309 ( .A(b[248]), .B(n2059), .Z(n2058) );
  XOR U2310 ( .A(n2057), .B(n2058), .Z(c[248]) );
  IV U2311 ( .A(a[249]), .Z(n2065) );
  NOR U2312 ( .A(n2058), .B(n2057), .Z(n2062) );
  IV U2313 ( .A(b[248]), .Z(n2060) );
  NOR U2314 ( .A(n2060), .B(n2059), .Z(n2061) );
  NOR U2315 ( .A(n2062), .B(n2061), .Z(n2067) );
  XOR U2316 ( .A(b[249]), .B(n2067), .Z(n2066) );
  XOR U2317 ( .A(n2065), .B(n2066), .Z(c[249]) );
  XOR U2318 ( .A(b[24]), .B(n2063), .Z(n2064) );
  XOR U2319 ( .A(a[24]), .B(n2064), .Z(c[24]) );
  IV U2320 ( .A(a[250]), .Z(n2071) );
  NOR U2321 ( .A(n2066), .B(n2065), .Z(n2070) );
  IV U2322 ( .A(b[249]), .Z(n2068) );
  NOR U2323 ( .A(n2068), .B(n2067), .Z(n2069) );
  NOR U2324 ( .A(n2070), .B(n2069), .Z(n2073) );
  XOR U2325 ( .A(b[250]), .B(n2073), .Z(n2072) );
  XOR U2326 ( .A(n2071), .B(n2072), .Z(c[250]) );
  IV U2327 ( .A(a[251]), .Z(n2077) );
  NOR U2328 ( .A(n2072), .B(n2071), .Z(n2076) );
  IV U2329 ( .A(b[250]), .Z(n2074) );
  NOR U2330 ( .A(n2074), .B(n2073), .Z(n2075) );
  NOR U2331 ( .A(n2076), .B(n2075), .Z(n2079) );
  XOR U2332 ( .A(b[251]), .B(n2079), .Z(n2078) );
  XOR U2333 ( .A(n2077), .B(n2078), .Z(c[251]) );
  IV U2334 ( .A(a[252]), .Z(n2083) );
  NOR U2335 ( .A(n2078), .B(n2077), .Z(n2082) );
  IV U2336 ( .A(b[251]), .Z(n2080) );
  NOR U2337 ( .A(n2080), .B(n2079), .Z(n2081) );
  NOR U2338 ( .A(n2082), .B(n2081), .Z(n2085) );
  XOR U2339 ( .A(b[252]), .B(n2085), .Z(n2084) );
  XOR U2340 ( .A(n2083), .B(n2084), .Z(c[252]) );
  IV U2341 ( .A(a[253]), .Z(n2089) );
  NOR U2342 ( .A(n2084), .B(n2083), .Z(n2088) );
  IV U2343 ( .A(b[252]), .Z(n2086) );
  NOR U2344 ( .A(n2086), .B(n2085), .Z(n2087) );
  NOR U2345 ( .A(n2088), .B(n2087), .Z(n2091) );
  XOR U2346 ( .A(b[253]), .B(n2091), .Z(n2090) );
  XOR U2347 ( .A(n2089), .B(n2090), .Z(c[253]) );
  IV U2348 ( .A(a[254]), .Z(n2095) );
  NOR U2349 ( .A(n2090), .B(n2089), .Z(n2094) );
  IV U2350 ( .A(b[253]), .Z(n2092) );
  NOR U2351 ( .A(n2092), .B(n2091), .Z(n2093) );
  NOR U2352 ( .A(n2094), .B(n2093), .Z(n2097) );
  XOR U2353 ( .A(b[254]), .B(n2097), .Z(n2096) );
  XOR U2354 ( .A(n2095), .B(n2096), .Z(c[254]) );
  NOR U2355 ( .A(n2096), .B(n2095), .Z(n2100) );
  IV U2356 ( .A(b[254]), .Z(n2098) );
  NOR U2357 ( .A(n2098), .B(n2097), .Z(n2099) );
  NOR U2358 ( .A(n2100), .B(n2099), .Z(n2269) );
  IV U2359 ( .A(n2269), .Z(n2270) );
  XOR U2360 ( .A(a[255]), .B(n2270), .Z(n2101) );
  XOR U2361 ( .A(b[255]), .B(n2101), .Z(c[255]) );
  XOR U2362 ( .A(b[25]), .B(n2102), .Z(n2103) );
  XOR U2363 ( .A(a[25]), .B(n2103), .Z(c[25]) );
  XOR U2364 ( .A(b[26]), .B(n2104), .Z(n2105) );
  XOR U2365 ( .A(a[26]), .B(n2105), .Z(c[26]) );
  XOR U2366 ( .A(b[27]), .B(n2106), .Z(n2107) );
  XOR U2367 ( .A(a[27]), .B(n2107), .Z(c[27]) );
  XOR U2368 ( .A(b[28]), .B(n2108), .Z(n2109) );
  XOR U2369 ( .A(a[28]), .B(n2109), .Z(c[28]) );
  XOR U2370 ( .A(b[29]), .B(n2110), .Z(n2111) );
  XOR U2371 ( .A(a[29]), .B(n2111), .Z(c[29]) );
  XOR U2372 ( .A(b[2]), .B(n2112), .Z(n2113) );
  XOR U2373 ( .A(n2114), .B(n2113), .Z(c[2]) );
  XOR U2374 ( .A(b[30]), .B(n2115), .Z(n2116) );
  XOR U2375 ( .A(a[30]), .B(n2116), .Z(c[30]) );
  XOR U2376 ( .A(b[31]), .B(n2117), .Z(n2118) );
  XOR U2377 ( .A(a[31]), .B(n2118), .Z(c[31]) );
  XOR U2378 ( .A(b[32]), .B(n2119), .Z(n2120) );
  XOR U2379 ( .A(a[32]), .B(n2120), .Z(c[32]) );
  XOR U2380 ( .A(b[33]), .B(n2121), .Z(n2122) );
  XOR U2381 ( .A(a[33]), .B(n2122), .Z(c[33]) );
  XOR U2382 ( .A(b[34]), .B(n2123), .Z(n2124) );
  XOR U2383 ( .A(a[34]), .B(n2124), .Z(c[34]) );
  XOR U2384 ( .A(b[35]), .B(n2125), .Z(n2126) );
  XOR U2385 ( .A(a[35]), .B(n2126), .Z(c[35]) );
  XOR U2386 ( .A(b[36]), .B(n2127), .Z(n2128) );
  XOR U2387 ( .A(a[36]), .B(n2128), .Z(c[36]) );
  XOR U2388 ( .A(b[37]), .B(n2129), .Z(n2130) );
  XOR U2389 ( .A(a[37]), .B(n2130), .Z(c[37]) );
  XOR U2390 ( .A(b[38]), .B(n2131), .Z(n2132) );
  XOR U2391 ( .A(a[38]), .B(n2132), .Z(c[38]) );
  XOR U2392 ( .A(b[39]), .B(n2133), .Z(n2134) );
  XOR U2393 ( .A(a[39]), .B(n2134), .Z(c[39]) );
  XOR U2394 ( .A(b[3]), .B(n2135), .Z(n2136) );
  XOR U2395 ( .A(a[3]), .B(n2136), .Z(c[3]) );
  XOR U2396 ( .A(b[40]), .B(n2137), .Z(n2138) );
  XOR U2397 ( .A(a[40]), .B(n2138), .Z(c[40]) );
  XOR U2398 ( .A(b[41]), .B(n2139), .Z(n2140) );
  XOR U2399 ( .A(a[41]), .B(n2140), .Z(c[41]) );
  XOR U2400 ( .A(b[42]), .B(n2141), .Z(n2142) );
  XOR U2401 ( .A(a[42]), .B(n2142), .Z(c[42]) );
  XOR U2402 ( .A(b[43]), .B(n2143), .Z(n2144) );
  XOR U2403 ( .A(a[43]), .B(n2144), .Z(c[43]) );
  XOR U2404 ( .A(b[44]), .B(n2145), .Z(n2146) );
  XOR U2405 ( .A(a[44]), .B(n2146), .Z(c[44]) );
  XOR U2406 ( .A(b[45]), .B(n2147), .Z(n2148) );
  XOR U2407 ( .A(a[45]), .B(n2148), .Z(c[45]) );
  XOR U2408 ( .A(b[46]), .B(n2149), .Z(n2150) );
  XOR U2409 ( .A(a[46]), .B(n2150), .Z(c[46]) );
  XOR U2410 ( .A(b[47]), .B(n2151), .Z(n2152) );
  XOR U2411 ( .A(a[47]), .B(n2152), .Z(c[47]) );
  XOR U2412 ( .A(b[48]), .B(n2153), .Z(n2154) );
  XOR U2413 ( .A(a[48]), .B(n2154), .Z(c[48]) );
  XOR U2414 ( .A(b[49]), .B(n2155), .Z(n2156) );
  XOR U2415 ( .A(a[49]), .B(n2156), .Z(c[49]) );
  XOR U2416 ( .A(b[4]), .B(n2157), .Z(n2158) );
  XOR U2417 ( .A(a[4]), .B(n2158), .Z(c[4]) );
  XOR U2418 ( .A(b[50]), .B(n2159), .Z(n2160) );
  XOR U2419 ( .A(a[50]), .B(n2160), .Z(c[50]) );
  XOR U2420 ( .A(b[51]), .B(n2161), .Z(n2162) );
  XOR U2421 ( .A(a[51]), .B(n2162), .Z(c[51]) );
  XOR U2422 ( .A(b[52]), .B(n2163), .Z(n2164) );
  XOR U2423 ( .A(a[52]), .B(n2164), .Z(c[52]) );
  XOR U2424 ( .A(b[53]), .B(n2165), .Z(n2166) );
  XOR U2425 ( .A(a[53]), .B(n2166), .Z(c[53]) );
  XOR U2426 ( .A(b[54]), .B(n2167), .Z(n2168) );
  XOR U2427 ( .A(a[54]), .B(n2168), .Z(c[54]) );
  XOR U2428 ( .A(b[55]), .B(n2169), .Z(n2170) );
  XOR U2429 ( .A(a[55]), .B(n2170), .Z(c[55]) );
  XOR U2430 ( .A(b[56]), .B(n2171), .Z(n2172) );
  XOR U2431 ( .A(a[56]), .B(n2172), .Z(c[56]) );
  XOR U2432 ( .A(b[57]), .B(n2173), .Z(n2174) );
  XOR U2433 ( .A(a[57]), .B(n2174), .Z(c[57]) );
  XOR U2434 ( .A(b[58]), .B(n2175), .Z(n2176) );
  XOR U2435 ( .A(a[58]), .B(n2176), .Z(c[58]) );
  XOR U2436 ( .A(b[59]), .B(n2177), .Z(n2178) );
  XOR U2437 ( .A(a[59]), .B(n2178), .Z(c[59]) );
  XOR U2438 ( .A(b[5]), .B(n2179), .Z(n2180) );
  XOR U2439 ( .A(a[5]), .B(n2180), .Z(c[5]) );
  XOR U2440 ( .A(b[60]), .B(n2181), .Z(n2182) );
  XOR U2441 ( .A(a[60]), .B(n2182), .Z(c[60]) );
  XOR U2442 ( .A(b[61]), .B(n2183), .Z(n2184) );
  XOR U2443 ( .A(a[61]), .B(n2184), .Z(c[61]) );
  XOR U2444 ( .A(b[62]), .B(n2185), .Z(n2186) );
  XOR U2445 ( .A(a[62]), .B(n2186), .Z(c[62]) );
  XOR U2446 ( .A(b[63]), .B(n2187), .Z(n2188) );
  XOR U2447 ( .A(a[63]), .B(n2188), .Z(c[63]) );
  XOR U2448 ( .A(b[64]), .B(n2189), .Z(n2190) );
  XOR U2449 ( .A(a[64]), .B(n2190), .Z(c[64]) );
  XOR U2450 ( .A(b[65]), .B(n2191), .Z(n2192) );
  XOR U2451 ( .A(a[65]), .B(n2192), .Z(c[65]) );
  XOR U2452 ( .A(b[66]), .B(n2193), .Z(n2194) );
  XOR U2453 ( .A(a[66]), .B(n2194), .Z(c[66]) );
  XOR U2454 ( .A(b[67]), .B(n2195), .Z(n2196) );
  XOR U2455 ( .A(a[67]), .B(n2196), .Z(c[67]) );
  XOR U2456 ( .A(b[68]), .B(n2197), .Z(n2198) );
  XOR U2457 ( .A(a[68]), .B(n2198), .Z(c[68]) );
  XOR U2458 ( .A(b[69]), .B(n2199), .Z(n2200) );
  XOR U2459 ( .A(a[69]), .B(n2200), .Z(c[69]) );
  XOR U2460 ( .A(b[6]), .B(n2201), .Z(n2202) );
  XOR U2461 ( .A(a[6]), .B(n2202), .Z(c[6]) );
  XOR U2462 ( .A(b[70]), .B(n2203), .Z(n2204) );
  XOR U2463 ( .A(a[70]), .B(n2204), .Z(c[70]) );
  XOR U2464 ( .A(b[71]), .B(n2205), .Z(n2206) );
  XOR U2465 ( .A(a[71]), .B(n2206), .Z(c[71]) );
  XOR U2466 ( .A(b[72]), .B(n2207), .Z(n2208) );
  XOR U2467 ( .A(a[72]), .B(n2208), .Z(c[72]) );
  XOR U2468 ( .A(b[73]), .B(n2209), .Z(n2210) );
  XOR U2469 ( .A(a[73]), .B(n2210), .Z(c[73]) );
  XOR U2470 ( .A(b[74]), .B(n2211), .Z(n2212) );
  XOR U2471 ( .A(a[74]), .B(n2212), .Z(c[74]) );
  XOR U2472 ( .A(b[75]), .B(n2213), .Z(n2214) );
  XOR U2473 ( .A(a[75]), .B(n2214), .Z(c[75]) );
  XOR U2474 ( .A(b[76]), .B(n2215), .Z(n2216) );
  XOR U2475 ( .A(a[76]), .B(n2216), .Z(c[76]) );
  XOR U2476 ( .A(b[77]), .B(n2217), .Z(n2218) );
  XOR U2477 ( .A(a[77]), .B(n2218), .Z(c[77]) );
  XOR U2478 ( .A(b[78]), .B(n2219), .Z(n2220) );
  XOR U2479 ( .A(a[78]), .B(n2220), .Z(c[78]) );
  XOR U2480 ( .A(b[79]), .B(n2221), .Z(n2222) );
  XOR U2481 ( .A(a[79]), .B(n2222), .Z(c[79]) );
  XOR U2482 ( .A(b[7]), .B(n2223), .Z(n2224) );
  XOR U2483 ( .A(a[7]), .B(n2224), .Z(c[7]) );
  XOR U2484 ( .A(b[80]), .B(n2225), .Z(n2226) );
  XOR U2485 ( .A(a[80]), .B(n2226), .Z(c[80]) );
  XOR U2486 ( .A(b[81]), .B(n2227), .Z(n2228) );
  XOR U2487 ( .A(a[81]), .B(n2228), .Z(c[81]) );
  XOR U2488 ( .A(b[82]), .B(n2229), .Z(n2230) );
  XOR U2489 ( .A(a[82]), .B(n2230), .Z(c[82]) );
  XOR U2490 ( .A(b[83]), .B(n2231), .Z(n2232) );
  XOR U2491 ( .A(a[83]), .B(n2232), .Z(c[83]) );
  XOR U2492 ( .A(b[84]), .B(n2233), .Z(n2234) );
  XOR U2493 ( .A(a[84]), .B(n2234), .Z(c[84]) );
  XOR U2494 ( .A(b[85]), .B(n2235), .Z(n2236) );
  XOR U2495 ( .A(a[85]), .B(n2236), .Z(c[85]) );
  XOR U2496 ( .A(b[86]), .B(n2237), .Z(n2238) );
  XOR U2497 ( .A(a[86]), .B(n2238), .Z(c[86]) );
  XOR U2498 ( .A(b[87]), .B(n2239), .Z(n2240) );
  XOR U2499 ( .A(a[87]), .B(n2240), .Z(c[87]) );
  XOR U2500 ( .A(b[88]), .B(n2241), .Z(n2242) );
  XOR U2501 ( .A(a[88]), .B(n2242), .Z(c[88]) );
  XOR U2502 ( .A(b[89]), .B(n2243), .Z(n2244) );
  XOR U2503 ( .A(a[89]), .B(n2244), .Z(c[89]) );
  XOR U2504 ( .A(b[8]), .B(n2245), .Z(n2246) );
  XOR U2505 ( .A(a[8]), .B(n2246), .Z(c[8]) );
  XOR U2506 ( .A(b[90]), .B(n2247), .Z(n2248) );
  XOR U2507 ( .A(a[90]), .B(n2248), .Z(c[90]) );
  XOR U2508 ( .A(b[91]), .B(n2249), .Z(n2250) );
  XOR U2509 ( .A(a[91]), .B(n2250), .Z(c[91]) );
  XOR U2510 ( .A(b[92]), .B(n2251), .Z(n2252) );
  XOR U2511 ( .A(a[92]), .B(n2252), .Z(c[92]) );
  XOR U2512 ( .A(b[93]), .B(n2253), .Z(n2254) );
  XOR U2513 ( .A(a[93]), .B(n2254), .Z(c[93]) );
  XOR U2514 ( .A(b[94]), .B(n2255), .Z(n2256) );
  XOR U2515 ( .A(a[94]), .B(n2256), .Z(c[94]) );
  XOR U2516 ( .A(b[95]), .B(n2257), .Z(n2258) );
  XOR U2517 ( .A(a[95]), .B(n2258), .Z(c[95]) );
  XOR U2518 ( .A(b[96]), .B(n2259), .Z(n2260) );
  XOR U2519 ( .A(a[96]), .B(n2260), .Z(c[96]) );
  XOR U2520 ( .A(b[97]), .B(n2261), .Z(n2262) );
  XOR U2521 ( .A(a[97]), .B(n2262), .Z(c[97]) );
  XOR U2522 ( .A(b[98]), .B(n2263), .Z(n2264) );
  XOR U2523 ( .A(a[98]), .B(n2264), .Z(c[98]) );
  XOR U2524 ( .A(a[99]), .B(n2265), .Z(n2266) );
  XOR U2525 ( .A(b[99]), .B(n2266), .Z(c[99]) );
  XOR U2526 ( .A(a[9]), .B(n2267), .Z(n2268) );
  XOR U2527 ( .A(b[9]), .B(n2268), .Z(c[9]) );
endmodule

