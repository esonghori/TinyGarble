
module compare_N16384_CC256 ( clk, rst, x, y, g );
  input [63:0] x;
  input [63:0] y;
  input clk, rst;
  output g;
  wire   ci, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320;

  DFF ci_reg ( .D(g), .CLK(clk), .RST(rst), .I(1'b1), .Q(ci) );
  XOR U68 ( .A(y[3]), .B(n307), .Z(n308) );
  XOR U69 ( .A(y[7]), .B(n291), .Z(n292) );
  XOR U70 ( .A(y[11]), .B(n275), .Z(n276) );
  XOR U71 ( .A(y[15]), .B(n259), .Z(n260) );
  XOR U72 ( .A(y[19]), .B(n243), .Z(n244) );
  XOR U73 ( .A(y[23]), .B(n227), .Z(n228) );
  XOR U74 ( .A(y[27]), .B(n211), .Z(n212) );
  XOR U75 ( .A(y[31]), .B(n195), .Z(n196) );
  XOR U76 ( .A(y[35]), .B(n179), .Z(n180) );
  XOR U77 ( .A(y[39]), .B(n163), .Z(n164) );
  XOR U78 ( .A(y[43]), .B(n147), .Z(n148) );
  XOR U79 ( .A(y[47]), .B(n131), .Z(n132) );
  XOR U80 ( .A(y[51]), .B(n115), .Z(n116) );
  XOR U81 ( .A(y[55]), .B(n99), .Z(n100) );
  XOR U82 ( .A(y[59]), .B(n83), .Z(n84) );
  XOR U83 ( .A(y[4]), .B(n303), .Z(n304) );
  XOR U84 ( .A(y[8]), .B(n287), .Z(n288) );
  XOR U85 ( .A(y[12]), .B(n271), .Z(n272) );
  XOR U86 ( .A(y[16]), .B(n255), .Z(n256) );
  XOR U87 ( .A(y[20]), .B(n239), .Z(n240) );
  XOR U88 ( .A(y[24]), .B(n223), .Z(n224) );
  XOR U89 ( .A(y[28]), .B(n207), .Z(n208) );
  XOR U90 ( .A(y[32]), .B(n191), .Z(n192) );
  XOR U91 ( .A(y[36]), .B(n175), .Z(n176) );
  XOR U92 ( .A(y[40]), .B(n159), .Z(n160) );
  XOR U93 ( .A(y[44]), .B(n143), .Z(n144) );
  XOR U94 ( .A(y[48]), .B(n127), .Z(n128) );
  XOR U95 ( .A(y[52]), .B(n111), .Z(n112) );
  XOR U96 ( .A(y[56]), .B(n95), .Z(n96) );
  XOR U97 ( .A(y[60]), .B(n79), .Z(n80) );
  XOR U98 ( .A(y[5]), .B(n299), .Z(n300) );
  XOR U99 ( .A(y[9]), .B(n283), .Z(n284) );
  XOR U100 ( .A(y[13]), .B(n267), .Z(n268) );
  XOR U101 ( .A(y[17]), .B(n251), .Z(n252) );
  XOR U102 ( .A(y[21]), .B(n235), .Z(n236) );
  XOR U103 ( .A(y[25]), .B(n219), .Z(n220) );
  XOR U104 ( .A(y[29]), .B(n203), .Z(n204) );
  XOR U105 ( .A(y[33]), .B(n187), .Z(n188) );
  XOR U106 ( .A(y[37]), .B(n171), .Z(n172) );
  XOR U107 ( .A(y[41]), .B(n155), .Z(n156) );
  XOR U108 ( .A(y[45]), .B(n139), .Z(n140) );
  XOR U109 ( .A(y[49]), .B(n123), .Z(n124) );
  XOR U110 ( .A(y[53]), .B(n107), .Z(n108) );
  XOR U111 ( .A(y[57]), .B(n91), .Z(n92) );
  XOR U112 ( .A(y[61]), .B(n75), .Z(n76) );
  XOR U113 ( .A(y[2]), .B(n311), .Z(n312) );
  XOR U114 ( .A(y[6]), .B(n295), .Z(n296) );
  XOR U115 ( .A(y[10]), .B(n279), .Z(n280) );
  XOR U116 ( .A(y[14]), .B(n263), .Z(n264) );
  XOR U117 ( .A(y[18]), .B(n247), .Z(n248) );
  XOR U118 ( .A(y[22]), .B(n231), .Z(n232) );
  XOR U119 ( .A(y[26]), .B(n215), .Z(n216) );
  XOR U120 ( .A(y[30]), .B(n199), .Z(n200) );
  XOR U121 ( .A(y[34]), .B(n183), .Z(n184) );
  XOR U122 ( .A(y[38]), .B(n167), .Z(n168) );
  XOR U123 ( .A(y[42]), .B(n151), .Z(n152) );
  XOR U124 ( .A(y[46]), .B(n135), .Z(n136) );
  XOR U125 ( .A(y[50]), .B(n119), .Z(n120) );
  XOR U126 ( .A(y[54]), .B(n103), .Z(n104) );
  XOR U127 ( .A(y[58]), .B(n87), .Z(n88) );
  XOR U128 ( .A(y[62]), .B(n71), .Z(n72) );
  XOR U129 ( .A(n66), .B(n67), .Z(g) );
  AND U130 ( .A(n68), .B(n69), .Z(n66) );
  XOR U131 ( .A(x[63]), .B(n67), .Z(n69) );
  XNOR U132 ( .A(y[63]), .B(n67), .Z(n68) );
  XNOR U133 ( .A(n70), .B(n71), .Z(n67) );
  AND U134 ( .A(n72), .B(n73), .Z(n70) );
  XNOR U135 ( .A(x[62]), .B(n71), .Z(n73) );
  XOR U136 ( .A(n74), .B(n75), .Z(n71) );
  AND U137 ( .A(n76), .B(n77), .Z(n74) );
  XNOR U138 ( .A(x[61]), .B(n75), .Z(n77) );
  XOR U139 ( .A(n78), .B(n79), .Z(n75) );
  AND U140 ( .A(n80), .B(n81), .Z(n78) );
  XNOR U141 ( .A(x[60]), .B(n79), .Z(n81) );
  XOR U142 ( .A(n82), .B(n83), .Z(n79) );
  AND U143 ( .A(n84), .B(n85), .Z(n82) );
  XNOR U144 ( .A(x[59]), .B(n83), .Z(n85) );
  XOR U145 ( .A(n86), .B(n87), .Z(n83) );
  AND U146 ( .A(n88), .B(n89), .Z(n86) );
  XNOR U147 ( .A(x[58]), .B(n87), .Z(n89) );
  XOR U148 ( .A(n90), .B(n91), .Z(n87) );
  AND U149 ( .A(n92), .B(n93), .Z(n90) );
  XNOR U150 ( .A(x[57]), .B(n91), .Z(n93) );
  XOR U151 ( .A(n94), .B(n95), .Z(n91) );
  AND U152 ( .A(n96), .B(n97), .Z(n94) );
  XNOR U153 ( .A(x[56]), .B(n95), .Z(n97) );
  XOR U154 ( .A(n98), .B(n99), .Z(n95) );
  AND U155 ( .A(n100), .B(n101), .Z(n98) );
  XNOR U156 ( .A(x[55]), .B(n99), .Z(n101) );
  XOR U157 ( .A(n102), .B(n103), .Z(n99) );
  AND U158 ( .A(n104), .B(n105), .Z(n102) );
  XNOR U159 ( .A(x[54]), .B(n103), .Z(n105) );
  XOR U160 ( .A(n106), .B(n107), .Z(n103) );
  AND U161 ( .A(n108), .B(n109), .Z(n106) );
  XNOR U162 ( .A(x[53]), .B(n107), .Z(n109) );
  XOR U163 ( .A(n110), .B(n111), .Z(n107) );
  AND U164 ( .A(n112), .B(n113), .Z(n110) );
  XNOR U165 ( .A(x[52]), .B(n111), .Z(n113) );
  XOR U166 ( .A(n114), .B(n115), .Z(n111) );
  AND U167 ( .A(n116), .B(n117), .Z(n114) );
  XNOR U168 ( .A(x[51]), .B(n115), .Z(n117) );
  XOR U169 ( .A(n118), .B(n119), .Z(n115) );
  AND U170 ( .A(n120), .B(n121), .Z(n118) );
  XNOR U171 ( .A(x[50]), .B(n119), .Z(n121) );
  XOR U172 ( .A(n122), .B(n123), .Z(n119) );
  AND U173 ( .A(n124), .B(n125), .Z(n122) );
  XNOR U174 ( .A(x[49]), .B(n123), .Z(n125) );
  XOR U175 ( .A(n126), .B(n127), .Z(n123) );
  AND U176 ( .A(n128), .B(n129), .Z(n126) );
  XNOR U177 ( .A(x[48]), .B(n127), .Z(n129) );
  XOR U178 ( .A(n130), .B(n131), .Z(n127) );
  AND U179 ( .A(n132), .B(n133), .Z(n130) );
  XNOR U180 ( .A(x[47]), .B(n131), .Z(n133) );
  XOR U181 ( .A(n134), .B(n135), .Z(n131) );
  AND U182 ( .A(n136), .B(n137), .Z(n134) );
  XNOR U183 ( .A(x[46]), .B(n135), .Z(n137) );
  XOR U184 ( .A(n138), .B(n139), .Z(n135) );
  AND U185 ( .A(n140), .B(n141), .Z(n138) );
  XNOR U186 ( .A(x[45]), .B(n139), .Z(n141) );
  XOR U187 ( .A(n142), .B(n143), .Z(n139) );
  AND U188 ( .A(n144), .B(n145), .Z(n142) );
  XNOR U189 ( .A(x[44]), .B(n143), .Z(n145) );
  XOR U190 ( .A(n146), .B(n147), .Z(n143) );
  AND U191 ( .A(n148), .B(n149), .Z(n146) );
  XNOR U192 ( .A(x[43]), .B(n147), .Z(n149) );
  XOR U193 ( .A(n150), .B(n151), .Z(n147) );
  AND U194 ( .A(n152), .B(n153), .Z(n150) );
  XNOR U195 ( .A(x[42]), .B(n151), .Z(n153) );
  XOR U196 ( .A(n154), .B(n155), .Z(n151) );
  AND U197 ( .A(n156), .B(n157), .Z(n154) );
  XNOR U198 ( .A(x[41]), .B(n155), .Z(n157) );
  XOR U199 ( .A(n158), .B(n159), .Z(n155) );
  AND U200 ( .A(n160), .B(n161), .Z(n158) );
  XNOR U201 ( .A(x[40]), .B(n159), .Z(n161) );
  XOR U202 ( .A(n162), .B(n163), .Z(n159) );
  AND U203 ( .A(n164), .B(n165), .Z(n162) );
  XNOR U204 ( .A(x[39]), .B(n163), .Z(n165) );
  XOR U205 ( .A(n166), .B(n167), .Z(n163) );
  AND U206 ( .A(n168), .B(n169), .Z(n166) );
  XNOR U207 ( .A(x[38]), .B(n167), .Z(n169) );
  XOR U208 ( .A(n170), .B(n171), .Z(n167) );
  AND U209 ( .A(n172), .B(n173), .Z(n170) );
  XNOR U210 ( .A(x[37]), .B(n171), .Z(n173) );
  XOR U211 ( .A(n174), .B(n175), .Z(n171) );
  AND U212 ( .A(n176), .B(n177), .Z(n174) );
  XNOR U213 ( .A(x[36]), .B(n175), .Z(n177) );
  XOR U214 ( .A(n178), .B(n179), .Z(n175) );
  AND U215 ( .A(n180), .B(n181), .Z(n178) );
  XNOR U216 ( .A(x[35]), .B(n179), .Z(n181) );
  XOR U217 ( .A(n182), .B(n183), .Z(n179) );
  AND U218 ( .A(n184), .B(n185), .Z(n182) );
  XNOR U219 ( .A(x[34]), .B(n183), .Z(n185) );
  XOR U220 ( .A(n186), .B(n187), .Z(n183) );
  AND U221 ( .A(n188), .B(n189), .Z(n186) );
  XNOR U222 ( .A(x[33]), .B(n187), .Z(n189) );
  XOR U223 ( .A(n190), .B(n191), .Z(n187) );
  AND U224 ( .A(n192), .B(n193), .Z(n190) );
  XNOR U225 ( .A(x[32]), .B(n191), .Z(n193) );
  XOR U226 ( .A(n194), .B(n195), .Z(n191) );
  AND U227 ( .A(n196), .B(n197), .Z(n194) );
  XNOR U228 ( .A(x[31]), .B(n195), .Z(n197) );
  XOR U229 ( .A(n198), .B(n199), .Z(n195) );
  AND U230 ( .A(n200), .B(n201), .Z(n198) );
  XNOR U231 ( .A(x[30]), .B(n199), .Z(n201) );
  XOR U232 ( .A(n202), .B(n203), .Z(n199) );
  AND U233 ( .A(n204), .B(n205), .Z(n202) );
  XNOR U234 ( .A(x[29]), .B(n203), .Z(n205) );
  XOR U235 ( .A(n206), .B(n207), .Z(n203) );
  AND U236 ( .A(n208), .B(n209), .Z(n206) );
  XNOR U237 ( .A(x[28]), .B(n207), .Z(n209) );
  XOR U238 ( .A(n210), .B(n211), .Z(n207) );
  AND U239 ( .A(n212), .B(n213), .Z(n210) );
  XNOR U240 ( .A(x[27]), .B(n211), .Z(n213) );
  XOR U241 ( .A(n214), .B(n215), .Z(n211) );
  AND U242 ( .A(n216), .B(n217), .Z(n214) );
  XNOR U243 ( .A(x[26]), .B(n215), .Z(n217) );
  XOR U244 ( .A(n218), .B(n219), .Z(n215) );
  AND U245 ( .A(n220), .B(n221), .Z(n218) );
  XNOR U246 ( .A(x[25]), .B(n219), .Z(n221) );
  XOR U247 ( .A(n222), .B(n223), .Z(n219) );
  AND U248 ( .A(n224), .B(n225), .Z(n222) );
  XNOR U249 ( .A(x[24]), .B(n223), .Z(n225) );
  XOR U250 ( .A(n226), .B(n227), .Z(n223) );
  AND U251 ( .A(n228), .B(n229), .Z(n226) );
  XNOR U252 ( .A(x[23]), .B(n227), .Z(n229) );
  XOR U253 ( .A(n230), .B(n231), .Z(n227) );
  AND U254 ( .A(n232), .B(n233), .Z(n230) );
  XNOR U255 ( .A(x[22]), .B(n231), .Z(n233) );
  XOR U256 ( .A(n234), .B(n235), .Z(n231) );
  AND U257 ( .A(n236), .B(n237), .Z(n234) );
  XNOR U258 ( .A(x[21]), .B(n235), .Z(n237) );
  XOR U259 ( .A(n238), .B(n239), .Z(n235) );
  AND U260 ( .A(n240), .B(n241), .Z(n238) );
  XNOR U261 ( .A(x[20]), .B(n239), .Z(n241) );
  XOR U262 ( .A(n242), .B(n243), .Z(n239) );
  AND U263 ( .A(n244), .B(n245), .Z(n242) );
  XNOR U264 ( .A(x[19]), .B(n243), .Z(n245) );
  XOR U265 ( .A(n246), .B(n247), .Z(n243) );
  AND U266 ( .A(n248), .B(n249), .Z(n246) );
  XNOR U267 ( .A(x[18]), .B(n247), .Z(n249) );
  XOR U268 ( .A(n250), .B(n251), .Z(n247) );
  AND U269 ( .A(n252), .B(n253), .Z(n250) );
  XNOR U270 ( .A(x[17]), .B(n251), .Z(n253) );
  XOR U271 ( .A(n254), .B(n255), .Z(n251) );
  AND U272 ( .A(n256), .B(n257), .Z(n254) );
  XNOR U273 ( .A(x[16]), .B(n255), .Z(n257) );
  XOR U274 ( .A(n258), .B(n259), .Z(n255) );
  AND U275 ( .A(n260), .B(n261), .Z(n258) );
  XNOR U276 ( .A(x[15]), .B(n259), .Z(n261) );
  XOR U277 ( .A(n262), .B(n263), .Z(n259) );
  AND U278 ( .A(n264), .B(n265), .Z(n262) );
  XNOR U279 ( .A(x[14]), .B(n263), .Z(n265) );
  XOR U280 ( .A(n266), .B(n267), .Z(n263) );
  AND U281 ( .A(n268), .B(n269), .Z(n266) );
  XNOR U282 ( .A(x[13]), .B(n267), .Z(n269) );
  XOR U283 ( .A(n270), .B(n271), .Z(n267) );
  AND U284 ( .A(n272), .B(n273), .Z(n270) );
  XNOR U285 ( .A(x[12]), .B(n271), .Z(n273) );
  XOR U286 ( .A(n274), .B(n275), .Z(n271) );
  AND U287 ( .A(n276), .B(n277), .Z(n274) );
  XNOR U288 ( .A(x[11]), .B(n275), .Z(n277) );
  XOR U289 ( .A(n278), .B(n279), .Z(n275) );
  AND U290 ( .A(n280), .B(n281), .Z(n278) );
  XNOR U291 ( .A(x[10]), .B(n279), .Z(n281) );
  XOR U292 ( .A(n282), .B(n283), .Z(n279) );
  AND U293 ( .A(n284), .B(n285), .Z(n282) );
  XNOR U294 ( .A(x[9]), .B(n283), .Z(n285) );
  XOR U295 ( .A(n286), .B(n287), .Z(n283) );
  AND U296 ( .A(n288), .B(n289), .Z(n286) );
  XNOR U297 ( .A(x[8]), .B(n287), .Z(n289) );
  XOR U298 ( .A(n290), .B(n291), .Z(n287) );
  AND U299 ( .A(n292), .B(n293), .Z(n290) );
  XNOR U300 ( .A(x[7]), .B(n291), .Z(n293) );
  XOR U301 ( .A(n294), .B(n295), .Z(n291) );
  AND U302 ( .A(n296), .B(n297), .Z(n294) );
  XNOR U303 ( .A(x[6]), .B(n295), .Z(n297) );
  XOR U304 ( .A(n298), .B(n299), .Z(n295) );
  AND U305 ( .A(n300), .B(n301), .Z(n298) );
  XNOR U306 ( .A(x[5]), .B(n299), .Z(n301) );
  XOR U307 ( .A(n302), .B(n303), .Z(n299) );
  AND U308 ( .A(n304), .B(n305), .Z(n302) );
  XNOR U309 ( .A(x[4]), .B(n303), .Z(n305) );
  XOR U310 ( .A(n306), .B(n307), .Z(n303) );
  AND U311 ( .A(n308), .B(n309), .Z(n306) );
  XNOR U312 ( .A(x[3]), .B(n307), .Z(n309) );
  XOR U313 ( .A(n310), .B(n311), .Z(n307) );
  AND U314 ( .A(n312), .B(n313), .Z(n310) );
  XNOR U315 ( .A(x[2]), .B(n311), .Z(n313) );
  XOR U316 ( .A(n314), .B(n315), .Z(n311) );
  AND U317 ( .A(n316), .B(n317), .Z(n314) );
  XNOR U318 ( .A(x[1]), .B(n315), .Z(n317) );
  XOR U319 ( .A(y[1]), .B(n315), .Z(n316) );
  XOR U320 ( .A(ci), .B(n318), .Z(n315) );
  NANDN U321 ( .A(n319), .B(n320), .Z(n318) );
  XOR U322 ( .A(x[0]), .B(ci), .Z(n320) );
  XOR U323 ( .A(y[0]), .B(ci), .Z(n319) );
endmodule

