
module sum_N256_CC8 ( clk, rst, a, b, c );
  input [31:0] a;
  input [31:0] b;
  output [31:0] c;
  input clk, rst;
  wire   N66, N67, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472;
  wire   [1:0] carry_on;

  DFF \carry_on_reg[1]  ( .D(N67), .CLK(clk), .RST(rst), .Q(carry_on[1]) );
  DFF \carry_on_reg[0]  ( .D(N66), .CLK(clk), .RST(rst), .Q(carry_on[0]) );
  DFF \rc_reg[31]  ( .D(n128), .CLK(clk), .RST(1'b0), .Q(c[31]) );
  DFF \rc_reg[30]  ( .D(n127), .CLK(clk), .RST(1'b0), .Q(c[30]) );
  DFF \rc_reg[29]  ( .D(n126), .CLK(clk), .RST(1'b0), .Q(c[29]) );
  DFF \rc_reg[28]  ( .D(n125), .CLK(clk), .RST(1'b0), .Q(c[28]) );
  DFF \rc_reg[27]  ( .D(n124), .CLK(clk), .RST(1'b0), .Q(c[27]) );
  DFF \rc_reg[26]  ( .D(n123), .CLK(clk), .RST(1'b0), .Q(c[26]) );
  DFF \rc_reg[25]  ( .D(n122), .CLK(clk), .RST(1'b0), .Q(c[25]) );
  DFF \rc_reg[24]  ( .D(n121), .CLK(clk), .RST(1'b0), .Q(c[24]) );
  DFF \rc_reg[23]  ( .D(n120), .CLK(clk), .RST(1'b0), .Q(c[23]) );
  DFF \rc_reg[22]  ( .D(n119), .CLK(clk), .RST(1'b0), .Q(c[22]) );
  DFF \rc_reg[21]  ( .D(n118), .CLK(clk), .RST(1'b0), .Q(c[21]) );
  DFF \rc_reg[20]  ( .D(n117), .CLK(clk), .RST(1'b0), .Q(c[20]) );
  DFF \rc_reg[19]  ( .D(n116), .CLK(clk), .RST(1'b0), .Q(c[19]) );
  DFF \rc_reg[18]  ( .D(n115), .CLK(clk), .RST(1'b0), .Q(c[18]) );
  DFF \rc_reg[17]  ( .D(n114), .CLK(clk), .RST(1'b0), .Q(c[17]) );
  DFF \rc_reg[16]  ( .D(n113), .CLK(clk), .RST(1'b0), .Q(c[16]) );
  DFF \rc_reg[15]  ( .D(n112), .CLK(clk), .RST(1'b0), .Q(c[15]) );
  DFF \rc_reg[14]  ( .D(n111), .CLK(clk), .RST(1'b0), .Q(c[14]) );
  DFF \rc_reg[13]  ( .D(n110), .CLK(clk), .RST(1'b0), .Q(c[13]) );
  DFF \rc_reg[12]  ( .D(n109), .CLK(clk), .RST(1'b0), .Q(c[12]) );
  DFF \rc_reg[11]  ( .D(n108), .CLK(clk), .RST(1'b0), .Q(c[11]) );
  DFF \rc_reg[10]  ( .D(n107), .CLK(clk), .RST(1'b0), .Q(c[10]) );
  DFF \rc_reg[9]  ( .D(n106), .CLK(clk), .RST(1'b0), .Q(c[9]) );
  DFF \rc_reg[8]  ( .D(n105), .CLK(clk), .RST(1'b0), .Q(c[8]) );
  DFF \rc_reg[7]  ( .D(n104), .CLK(clk), .RST(1'b0), .Q(c[7]) );
  DFF \rc_reg[6]  ( .D(n103), .CLK(clk), .RST(1'b0), .Q(c[6]) );
  DFF \rc_reg[5]  ( .D(n102), .CLK(clk), .RST(1'b0), .Q(c[5]) );
  DFF \rc_reg[4]  ( .D(n101), .CLK(clk), .RST(1'b0), .Q(c[4]) );
  DFF \rc_reg[3]  ( .D(n100), .CLK(clk), .RST(1'b0), .Q(c[3]) );
  DFF \rc_reg[2]  ( .D(n99), .CLK(clk), .RST(1'b0), .Q(c[2]) );
  DFF \rc_reg[1]  ( .D(n98), .CLK(clk), .RST(1'b0), .Q(c[1]) );
  DFF \rc_reg[0]  ( .D(n97), .CLK(clk), .RST(1'b0), .Q(c[0]) );
  NANDN U131 ( .A(n305), .B(n306), .Z(n129) );
  NANDN U132 ( .A(n459), .B(n458), .Z(n130) );
  AND U133 ( .A(n129), .B(n130), .Z(n131) );
  NAND U134 ( .A(n464), .B(n463), .Z(n132) );
  NANDN U135 ( .A(n131), .B(n307), .Z(n133) );
  AND U136 ( .A(n132), .B(n133), .Z(n308) );
  XOR U137 ( .A(n188), .B(n187), .Z(n358) );
  XOR U138 ( .A(n212), .B(n211), .Z(n378) );
  XOR U139 ( .A(n236), .B(n235), .Z(n398) );
  XOR U140 ( .A(n260), .B(n259), .Z(n418) );
  XOR U141 ( .A(n284), .B(n283), .Z(n438) );
  XOR U142 ( .A(n151), .B(n150), .Z(n328) );
  XOR U143 ( .A(n176), .B(n175), .Z(n348) );
  XOR U144 ( .A(n200), .B(n199), .Z(n368) );
  XOR U145 ( .A(n224), .B(n223), .Z(n388) );
  XOR U146 ( .A(n248), .B(n247), .Z(n408) );
  XOR U147 ( .A(n272), .B(n271), .Z(n428) );
  XOR U148 ( .A(n296), .B(n295), .Z(n448) );
  AND U149 ( .A(b[31]), .B(a[31]), .Z(n313) );
  NAND U150 ( .A(a[29]), .B(b[29]), .Z(n307) );
  AND U151 ( .A(a[28]), .B(b[28]), .Z(n305) );
  XNOR U152 ( .A(a[1]), .B(b[1]), .Z(n136) );
  XNOR U153 ( .A(carry_on[1]), .B(n136), .Z(n319) );
  NAND U154 ( .A(a[0]), .B(b[0]), .Z(n135) );
  XOR U155 ( .A(a[0]), .B(b[0]), .Z(n314) );
  NAND U156 ( .A(n314), .B(carry_on[0]), .Z(n134) );
  NAND U157 ( .A(n135), .B(n134), .Z(n318) );
  NAND U158 ( .A(n319), .B(n318), .Z(n138) );
  ANDN U159 ( .B(carry_on[1]), .A(n136), .Z(n139) );
  ANDN U160 ( .B(n138), .A(n139), .Z(n137) );
  NAND U161 ( .A(a[1]), .B(b[1]), .Z(n140) );
  NAND U162 ( .A(n137), .B(n140), .Z(n144) );
  XNOR U163 ( .A(n140), .B(n138), .Z(n142) );
  NAND U164 ( .A(n140), .B(n139), .Z(n141) );
  NAND U165 ( .A(n142), .B(n141), .Z(n324) );
  XNOR U166 ( .A(a[2]), .B(b[2]), .Z(n323) );
  NAND U167 ( .A(n324), .B(n323), .Z(n143) );
  NAND U168 ( .A(n144), .B(n143), .Z(n150) );
  NAND U169 ( .A(a[2]), .B(b[2]), .Z(n151) );
  AND U170 ( .A(n150), .B(n151), .Z(n146) );
  XOR U171 ( .A(a[3]), .B(b[3]), .Z(n329) );
  ANDN U172 ( .B(n328), .A(n329), .Z(n145) );
  OR U173 ( .A(n146), .B(n145), .Z(n147) );
  AND U174 ( .A(a[3]), .B(b[3]), .Z(n149) );
  ANDN U175 ( .B(n147), .A(n149), .Z(n156) );
  NOR U176 ( .A(n151), .B(n150), .Z(n148) );
  XNOR U177 ( .A(n149), .B(n148), .Z(n154) );
  XOR U178 ( .A(n151), .B(n150), .Z(n152) );
  NAND U179 ( .A(n152), .B(n329), .Z(n153) );
  NAND U180 ( .A(n154), .B(n153), .Z(n334) );
  XNOR U181 ( .A(a[4]), .B(b[4]), .Z(n333) );
  NAND U182 ( .A(n334), .B(n333), .Z(n155) );
  NANDN U183 ( .A(n156), .B(n155), .Z(n163) );
  AND U184 ( .A(a[4]), .B(b[4]), .Z(n157) );
  IV U185 ( .A(n157), .Z(n164) );
  AND U186 ( .A(n163), .B(n164), .Z(n159) );
  XOR U187 ( .A(a[5]), .B(b[5]), .Z(n339) );
  XNOR U188 ( .A(n157), .B(n163), .Z(n338) );
  NANDN U189 ( .A(n339), .B(n338), .Z(n158) );
  NANDN U190 ( .A(n159), .B(n158), .Z(n160) );
  AND U191 ( .A(a[5]), .B(b[5]), .Z(n162) );
  ANDN U192 ( .B(n160), .A(n162), .Z(n169) );
  NOR U193 ( .A(n164), .B(n163), .Z(n161) );
  XNOR U194 ( .A(n162), .B(n161), .Z(n167) );
  XOR U195 ( .A(n164), .B(n163), .Z(n165) );
  NAND U196 ( .A(n165), .B(n339), .Z(n166) );
  NAND U197 ( .A(n167), .B(n166), .Z(n344) );
  XNOR U198 ( .A(a[6]), .B(b[6]), .Z(n343) );
  NAND U199 ( .A(n344), .B(n343), .Z(n168) );
  NANDN U200 ( .A(n169), .B(n168), .Z(n175) );
  NAND U201 ( .A(a[6]), .B(b[6]), .Z(n176) );
  AND U202 ( .A(n175), .B(n176), .Z(n171) );
  XOR U203 ( .A(a[7]), .B(b[7]), .Z(n349) );
  ANDN U204 ( .B(n348), .A(n349), .Z(n170) );
  OR U205 ( .A(n171), .B(n170), .Z(n172) );
  AND U206 ( .A(a[7]), .B(b[7]), .Z(n174) );
  ANDN U207 ( .B(n172), .A(n174), .Z(n181) );
  NOR U208 ( .A(n176), .B(n175), .Z(n173) );
  XNOR U209 ( .A(n174), .B(n173), .Z(n179) );
  XOR U210 ( .A(n176), .B(n175), .Z(n177) );
  NAND U211 ( .A(n177), .B(n349), .Z(n178) );
  NAND U212 ( .A(n179), .B(n178), .Z(n354) );
  XNOR U213 ( .A(a[8]), .B(b[8]), .Z(n353) );
  NAND U214 ( .A(n354), .B(n353), .Z(n180) );
  NANDN U215 ( .A(n181), .B(n180), .Z(n187) );
  NAND U216 ( .A(a[8]), .B(b[8]), .Z(n188) );
  AND U217 ( .A(n187), .B(n188), .Z(n183) );
  XOR U218 ( .A(a[9]), .B(b[9]), .Z(n359) );
  ANDN U219 ( .B(n358), .A(n359), .Z(n182) );
  OR U220 ( .A(n183), .B(n182), .Z(n184) );
  AND U221 ( .A(a[9]), .B(b[9]), .Z(n186) );
  ANDN U222 ( .B(n184), .A(n186), .Z(n193) );
  NOR U223 ( .A(n188), .B(n187), .Z(n185) );
  XNOR U224 ( .A(n186), .B(n185), .Z(n191) );
  XOR U225 ( .A(n188), .B(n187), .Z(n189) );
  NAND U226 ( .A(n189), .B(n359), .Z(n190) );
  NAND U227 ( .A(n191), .B(n190), .Z(n364) );
  XNOR U228 ( .A(a[10]), .B(b[10]), .Z(n363) );
  NAND U229 ( .A(n364), .B(n363), .Z(n192) );
  NANDN U230 ( .A(n193), .B(n192), .Z(n199) );
  NAND U231 ( .A(a[10]), .B(b[10]), .Z(n200) );
  AND U232 ( .A(n199), .B(n200), .Z(n195) );
  XOR U233 ( .A(a[11]), .B(b[11]), .Z(n369) );
  ANDN U234 ( .B(n368), .A(n369), .Z(n194) );
  OR U235 ( .A(n195), .B(n194), .Z(n196) );
  AND U236 ( .A(a[11]), .B(b[11]), .Z(n198) );
  ANDN U237 ( .B(n196), .A(n198), .Z(n205) );
  NOR U238 ( .A(n200), .B(n199), .Z(n197) );
  XNOR U239 ( .A(n198), .B(n197), .Z(n203) );
  XOR U240 ( .A(n200), .B(n199), .Z(n201) );
  NAND U241 ( .A(n201), .B(n369), .Z(n202) );
  NAND U242 ( .A(n203), .B(n202), .Z(n374) );
  XNOR U243 ( .A(a[12]), .B(b[12]), .Z(n373) );
  NAND U244 ( .A(n374), .B(n373), .Z(n204) );
  NANDN U245 ( .A(n205), .B(n204), .Z(n211) );
  NAND U246 ( .A(a[12]), .B(b[12]), .Z(n212) );
  AND U247 ( .A(n211), .B(n212), .Z(n207) );
  XOR U248 ( .A(a[13]), .B(b[13]), .Z(n379) );
  ANDN U249 ( .B(n378), .A(n379), .Z(n206) );
  OR U250 ( .A(n207), .B(n206), .Z(n208) );
  AND U251 ( .A(a[13]), .B(b[13]), .Z(n210) );
  ANDN U252 ( .B(n208), .A(n210), .Z(n217) );
  NOR U253 ( .A(n212), .B(n211), .Z(n209) );
  XNOR U254 ( .A(n210), .B(n209), .Z(n215) );
  XOR U255 ( .A(n212), .B(n211), .Z(n213) );
  NAND U256 ( .A(n213), .B(n379), .Z(n214) );
  NAND U257 ( .A(n215), .B(n214), .Z(n384) );
  XNOR U258 ( .A(a[14]), .B(b[14]), .Z(n383) );
  NAND U259 ( .A(n384), .B(n383), .Z(n216) );
  NANDN U260 ( .A(n217), .B(n216), .Z(n223) );
  NAND U261 ( .A(a[14]), .B(b[14]), .Z(n224) );
  AND U262 ( .A(n223), .B(n224), .Z(n219) );
  XOR U263 ( .A(a[15]), .B(b[15]), .Z(n389) );
  ANDN U264 ( .B(n388), .A(n389), .Z(n218) );
  OR U265 ( .A(n219), .B(n218), .Z(n220) );
  AND U266 ( .A(a[15]), .B(b[15]), .Z(n222) );
  ANDN U267 ( .B(n220), .A(n222), .Z(n229) );
  NOR U268 ( .A(n224), .B(n223), .Z(n221) );
  XNOR U269 ( .A(n222), .B(n221), .Z(n227) );
  XOR U270 ( .A(n224), .B(n223), .Z(n225) );
  NAND U271 ( .A(n225), .B(n389), .Z(n226) );
  NAND U272 ( .A(n227), .B(n226), .Z(n394) );
  XNOR U273 ( .A(a[16]), .B(b[16]), .Z(n393) );
  NAND U274 ( .A(n394), .B(n393), .Z(n228) );
  NANDN U275 ( .A(n229), .B(n228), .Z(n235) );
  NAND U276 ( .A(a[16]), .B(b[16]), .Z(n236) );
  AND U277 ( .A(n235), .B(n236), .Z(n231) );
  XOR U278 ( .A(a[17]), .B(b[17]), .Z(n399) );
  ANDN U279 ( .B(n398), .A(n399), .Z(n230) );
  OR U280 ( .A(n231), .B(n230), .Z(n232) );
  AND U281 ( .A(a[17]), .B(b[17]), .Z(n234) );
  ANDN U282 ( .B(n232), .A(n234), .Z(n241) );
  NOR U283 ( .A(n236), .B(n235), .Z(n233) );
  XNOR U284 ( .A(n234), .B(n233), .Z(n239) );
  XOR U285 ( .A(n236), .B(n235), .Z(n237) );
  NAND U286 ( .A(n237), .B(n399), .Z(n238) );
  NAND U287 ( .A(n239), .B(n238), .Z(n404) );
  XNOR U288 ( .A(a[18]), .B(b[18]), .Z(n403) );
  NAND U289 ( .A(n404), .B(n403), .Z(n240) );
  NANDN U290 ( .A(n241), .B(n240), .Z(n247) );
  NAND U291 ( .A(a[18]), .B(b[18]), .Z(n248) );
  AND U292 ( .A(n247), .B(n248), .Z(n243) );
  XOR U293 ( .A(a[19]), .B(b[19]), .Z(n409) );
  ANDN U294 ( .B(n408), .A(n409), .Z(n242) );
  OR U295 ( .A(n243), .B(n242), .Z(n244) );
  AND U296 ( .A(a[19]), .B(b[19]), .Z(n246) );
  ANDN U297 ( .B(n244), .A(n246), .Z(n253) );
  NOR U298 ( .A(n248), .B(n247), .Z(n245) );
  XNOR U299 ( .A(n246), .B(n245), .Z(n251) );
  XOR U300 ( .A(n248), .B(n247), .Z(n249) );
  NAND U301 ( .A(n249), .B(n409), .Z(n250) );
  NAND U302 ( .A(n251), .B(n250), .Z(n414) );
  XNOR U303 ( .A(a[20]), .B(b[20]), .Z(n413) );
  NAND U304 ( .A(n414), .B(n413), .Z(n252) );
  NANDN U305 ( .A(n253), .B(n252), .Z(n259) );
  NAND U306 ( .A(a[20]), .B(b[20]), .Z(n260) );
  AND U307 ( .A(n259), .B(n260), .Z(n255) );
  XOR U308 ( .A(a[21]), .B(b[21]), .Z(n419) );
  ANDN U309 ( .B(n418), .A(n419), .Z(n254) );
  OR U310 ( .A(n255), .B(n254), .Z(n256) );
  AND U311 ( .A(a[21]), .B(b[21]), .Z(n258) );
  ANDN U312 ( .B(n256), .A(n258), .Z(n265) );
  NOR U313 ( .A(n260), .B(n259), .Z(n257) );
  XNOR U314 ( .A(n258), .B(n257), .Z(n263) );
  XOR U315 ( .A(n260), .B(n259), .Z(n261) );
  NAND U316 ( .A(n261), .B(n419), .Z(n262) );
  NAND U317 ( .A(n263), .B(n262), .Z(n424) );
  XNOR U318 ( .A(a[22]), .B(b[22]), .Z(n423) );
  NAND U319 ( .A(n424), .B(n423), .Z(n264) );
  NANDN U320 ( .A(n265), .B(n264), .Z(n271) );
  NAND U321 ( .A(a[22]), .B(b[22]), .Z(n272) );
  AND U322 ( .A(n271), .B(n272), .Z(n267) );
  XOR U323 ( .A(a[23]), .B(b[23]), .Z(n429) );
  ANDN U324 ( .B(n428), .A(n429), .Z(n266) );
  OR U325 ( .A(n267), .B(n266), .Z(n268) );
  AND U326 ( .A(a[23]), .B(b[23]), .Z(n270) );
  ANDN U327 ( .B(n268), .A(n270), .Z(n277) );
  NOR U328 ( .A(n272), .B(n271), .Z(n269) );
  XNOR U329 ( .A(n270), .B(n269), .Z(n275) );
  XOR U330 ( .A(n272), .B(n271), .Z(n273) );
  NAND U331 ( .A(n273), .B(n429), .Z(n274) );
  NAND U332 ( .A(n275), .B(n274), .Z(n434) );
  XNOR U333 ( .A(a[24]), .B(b[24]), .Z(n433) );
  NAND U334 ( .A(n434), .B(n433), .Z(n276) );
  NANDN U335 ( .A(n277), .B(n276), .Z(n283) );
  NAND U336 ( .A(a[24]), .B(b[24]), .Z(n284) );
  AND U337 ( .A(n283), .B(n284), .Z(n279) );
  XOR U338 ( .A(a[25]), .B(b[25]), .Z(n439) );
  ANDN U339 ( .B(n438), .A(n439), .Z(n278) );
  OR U340 ( .A(n279), .B(n278), .Z(n280) );
  AND U341 ( .A(a[25]), .B(b[25]), .Z(n282) );
  ANDN U342 ( .B(n280), .A(n282), .Z(n289) );
  NOR U343 ( .A(n284), .B(n283), .Z(n281) );
  XNOR U344 ( .A(n282), .B(n281), .Z(n287) );
  XOR U345 ( .A(n284), .B(n283), .Z(n285) );
  NAND U346 ( .A(n285), .B(n439), .Z(n286) );
  NAND U347 ( .A(n287), .B(n286), .Z(n444) );
  XNOR U348 ( .A(a[26]), .B(b[26]), .Z(n443) );
  NAND U349 ( .A(n444), .B(n443), .Z(n288) );
  NANDN U350 ( .A(n289), .B(n288), .Z(n295) );
  NAND U351 ( .A(a[26]), .B(b[26]), .Z(n296) );
  AND U352 ( .A(n295), .B(n296), .Z(n291) );
  XOR U353 ( .A(a[27]), .B(b[27]), .Z(n449) );
  ANDN U354 ( .B(n448), .A(n449), .Z(n290) );
  OR U355 ( .A(n291), .B(n290), .Z(n292) );
  AND U356 ( .A(a[27]), .B(b[27]), .Z(n294) );
  ANDN U357 ( .B(n292), .A(n294), .Z(n301) );
  NOR U358 ( .A(n296), .B(n295), .Z(n293) );
  XNOR U359 ( .A(n294), .B(n293), .Z(n299) );
  XOR U360 ( .A(n296), .B(n295), .Z(n297) );
  NAND U361 ( .A(n297), .B(n449), .Z(n298) );
  NAND U362 ( .A(n299), .B(n298), .Z(n454) );
  XNOR U363 ( .A(a[28]), .B(b[28]), .Z(n453) );
  NAND U364 ( .A(n454), .B(n453), .Z(n300) );
  NANDN U365 ( .A(n301), .B(n300), .Z(n306) );
  ANDN U366 ( .B(n305), .A(n306), .Z(n302) );
  XOR U367 ( .A(n307), .B(n302), .Z(n304) );
  XOR U368 ( .A(a[29]), .B(b[29]), .Z(n459) );
  XNOR U369 ( .A(n305), .B(n306), .Z(n458) );
  NAND U370 ( .A(n459), .B(n458), .Z(n303) );
  NAND U371 ( .A(n304), .B(n303), .Z(n464) );
  XNOR U372 ( .A(a[30]), .B(b[30]), .Z(n463) );
  NAND U373 ( .A(a[30]), .B(b[30]), .Z(n309) );
  ANDN U374 ( .B(n308), .A(n309), .Z(n312) );
  XNOR U375 ( .A(n313), .B(n312), .Z(n311) );
  XNOR U376 ( .A(n309), .B(n308), .Z(n468) );
  XOR U377 ( .A(b[31]), .B(a[31]), .Z(n469) );
  NAND U378 ( .A(n468), .B(n469), .Z(n310) );
  NAND U379 ( .A(n311), .B(n310), .Z(N66) );
  AND U380 ( .A(n313), .B(n312), .Z(N67) );
  NAND U382 ( .A(c[0]), .B(rst), .Z(n317) );
  XOR U383 ( .A(n314), .B(carry_on[0]), .Z(n315) );
  NANDN U384 ( .A(rst), .B(n315), .Z(n316) );
  NAND U385 ( .A(n317), .B(n316), .Z(n97) );
  NAND U386 ( .A(c[1]), .B(rst), .Z(n322) );
  XOR U387 ( .A(n319), .B(n318), .Z(n320) );
  NANDN U388 ( .A(rst), .B(n320), .Z(n321) );
  NAND U389 ( .A(n322), .B(n321), .Z(n98) );
  NAND U390 ( .A(c[2]), .B(rst), .Z(n327) );
  XNOR U391 ( .A(n324), .B(n323), .Z(n325) );
  NANDN U392 ( .A(rst), .B(n325), .Z(n326) );
  NAND U393 ( .A(n327), .B(n326), .Z(n99) );
  NAND U394 ( .A(c[3]), .B(rst), .Z(n332) );
  XOR U395 ( .A(n329), .B(n328), .Z(n330) );
  NANDN U396 ( .A(rst), .B(n330), .Z(n331) );
  NAND U397 ( .A(n332), .B(n331), .Z(n100) );
  NAND U398 ( .A(c[4]), .B(rst), .Z(n337) );
  XNOR U399 ( .A(n334), .B(n333), .Z(n335) );
  NANDN U400 ( .A(rst), .B(n335), .Z(n336) );
  NAND U401 ( .A(n337), .B(n336), .Z(n101) );
  NAND U402 ( .A(c[5]), .B(rst), .Z(n342) );
  XOR U403 ( .A(n339), .B(n338), .Z(n340) );
  NANDN U404 ( .A(rst), .B(n340), .Z(n341) );
  NAND U405 ( .A(n342), .B(n341), .Z(n102) );
  NAND U406 ( .A(c[6]), .B(rst), .Z(n347) );
  XNOR U407 ( .A(n344), .B(n343), .Z(n345) );
  NANDN U408 ( .A(rst), .B(n345), .Z(n346) );
  NAND U409 ( .A(n347), .B(n346), .Z(n103) );
  NAND U410 ( .A(c[7]), .B(rst), .Z(n352) );
  XOR U411 ( .A(n349), .B(n348), .Z(n350) );
  NANDN U412 ( .A(rst), .B(n350), .Z(n351) );
  NAND U413 ( .A(n352), .B(n351), .Z(n104) );
  NAND U414 ( .A(c[8]), .B(rst), .Z(n357) );
  XNOR U415 ( .A(n354), .B(n353), .Z(n355) );
  NANDN U416 ( .A(rst), .B(n355), .Z(n356) );
  NAND U417 ( .A(n357), .B(n356), .Z(n105) );
  NAND U418 ( .A(c[9]), .B(rst), .Z(n362) );
  XOR U419 ( .A(n359), .B(n358), .Z(n360) );
  NANDN U420 ( .A(rst), .B(n360), .Z(n361) );
  NAND U421 ( .A(n362), .B(n361), .Z(n106) );
  NAND U422 ( .A(c[10]), .B(rst), .Z(n367) );
  XNOR U423 ( .A(n364), .B(n363), .Z(n365) );
  NANDN U424 ( .A(rst), .B(n365), .Z(n366) );
  NAND U425 ( .A(n367), .B(n366), .Z(n107) );
  NAND U426 ( .A(c[11]), .B(rst), .Z(n372) );
  XOR U427 ( .A(n369), .B(n368), .Z(n370) );
  NANDN U428 ( .A(rst), .B(n370), .Z(n371) );
  NAND U429 ( .A(n372), .B(n371), .Z(n108) );
  NAND U430 ( .A(c[12]), .B(rst), .Z(n377) );
  XNOR U431 ( .A(n374), .B(n373), .Z(n375) );
  NANDN U432 ( .A(rst), .B(n375), .Z(n376) );
  NAND U433 ( .A(n377), .B(n376), .Z(n109) );
  NAND U434 ( .A(c[13]), .B(rst), .Z(n382) );
  XOR U435 ( .A(n379), .B(n378), .Z(n380) );
  NANDN U436 ( .A(rst), .B(n380), .Z(n381) );
  NAND U437 ( .A(n382), .B(n381), .Z(n110) );
  NAND U438 ( .A(c[14]), .B(rst), .Z(n387) );
  XNOR U439 ( .A(n384), .B(n383), .Z(n385) );
  NANDN U440 ( .A(rst), .B(n385), .Z(n386) );
  NAND U441 ( .A(n387), .B(n386), .Z(n111) );
  NAND U442 ( .A(c[15]), .B(rst), .Z(n392) );
  XOR U443 ( .A(n389), .B(n388), .Z(n390) );
  NANDN U444 ( .A(rst), .B(n390), .Z(n391) );
  NAND U445 ( .A(n392), .B(n391), .Z(n112) );
  NAND U446 ( .A(c[16]), .B(rst), .Z(n397) );
  XNOR U447 ( .A(n394), .B(n393), .Z(n395) );
  NANDN U448 ( .A(rst), .B(n395), .Z(n396) );
  NAND U449 ( .A(n397), .B(n396), .Z(n113) );
  NAND U450 ( .A(c[17]), .B(rst), .Z(n402) );
  XOR U451 ( .A(n399), .B(n398), .Z(n400) );
  NANDN U452 ( .A(rst), .B(n400), .Z(n401) );
  NAND U453 ( .A(n402), .B(n401), .Z(n114) );
  NAND U454 ( .A(c[18]), .B(rst), .Z(n407) );
  XNOR U455 ( .A(n404), .B(n403), .Z(n405) );
  NANDN U456 ( .A(rst), .B(n405), .Z(n406) );
  NAND U457 ( .A(n407), .B(n406), .Z(n115) );
  NAND U458 ( .A(c[19]), .B(rst), .Z(n412) );
  XOR U459 ( .A(n409), .B(n408), .Z(n410) );
  NANDN U460 ( .A(rst), .B(n410), .Z(n411) );
  NAND U461 ( .A(n412), .B(n411), .Z(n116) );
  NAND U462 ( .A(c[20]), .B(rst), .Z(n417) );
  XNOR U463 ( .A(n414), .B(n413), .Z(n415) );
  NANDN U464 ( .A(rst), .B(n415), .Z(n416) );
  NAND U465 ( .A(n417), .B(n416), .Z(n117) );
  NAND U466 ( .A(c[21]), .B(rst), .Z(n422) );
  XOR U467 ( .A(n419), .B(n418), .Z(n420) );
  NANDN U468 ( .A(rst), .B(n420), .Z(n421) );
  NAND U469 ( .A(n422), .B(n421), .Z(n118) );
  NAND U470 ( .A(c[22]), .B(rst), .Z(n427) );
  XNOR U471 ( .A(n424), .B(n423), .Z(n425) );
  NANDN U472 ( .A(rst), .B(n425), .Z(n426) );
  NAND U473 ( .A(n427), .B(n426), .Z(n119) );
  NAND U474 ( .A(c[23]), .B(rst), .Z(n432) );
  XOR U475 ( .A(n429), .B(n428), .Z(n430) );
  NANDN U476 ( .A(rst), .B(n430), .Z(n431) );
  NAND U477 ( .A(n432), .B(n431), .Z(n120) );
  NAND U478 ( .A(c[24]), .B(rst), .Z(n437) );
  XNOR U479 ( .A(n434), .B(n433), .Z(n435) );
  NANDN U480 ( .A(rst), .B(n435), .Z(n436) );
  NAND U481 ( .A(n437), .B(n436), .Z(n121) );
  NAND U482 ( .A(c[25]), .B(rst), .Z(n442) );
  XOR U483 ( .A(n439), .B(n438), .Z(n440) );
  NANDN U484 ( .A(rst), .B(n440), .Z(n441) );
  NAND U485 ( .A(n442), .B(n441), .Z(n122) );
  NAND U486 ( .A(c[26]), .B(rst), .Z(n447) );
  XNOR U487 ( .A(n444), .B(n443), .Z(n445) );
  NANDN U488 ( .A(rst), .B(n445), .Z(n446) );
  NAND U489 ( .A(n447), .B(n446), .Z(n123) );
  NAND U490 ( .A(c[27]), .B(rst), .Z(n452) );
  XOR U491 ( .A(n449), .B(n448), .Z(n450) );
  NANDN U492 ( .A(rst), .B(n450), .Z(n451) );
  NAND U493 ( .A(n452), .B(n451), .Z(n124) );
  NAND U494 ( .A(c[28]), .B(rst), .Z(n457) );
  XNOR U495 ( .A(n454), .B(n453), .Z(n455) );
  NANDN U496 ( .A(rst), .B(n455), .Z(n456) );
  NAND U497 ( .A(n457), .B(n456), .Z(n125) );
  NAND U498 ( .A(c[29]), .B(rst), .Z(n462) );
  XOR U499 ( .A(n459), .B(n458), .Z(n460) );
  NANDN U500 ( .A(rst), .B(n460), .Z(n461) );
  NAND U501 ( .A(n462), .B(n461), .Z(n126) );
  NAND U502 ( .A(c[30]), .B(rst), .Z(n467) );
  XNOR U503 ( .A(n464), .B(n463), .Z(n465) );
  NANDN U504 ( .A(rst), .B(n465), .Z(n466) );
  NAND U505 ( .A(n467), .B(n466), .Z(n127) );
  NAND U506 ( .A(c[31]), .B(rst), .Z(n472) );
  XOR U507 ( .A(n469), .B(n468), .Z(n470) );
  NANDN U508 ( .A(rst), .B(n470), .Z(n471) );
  NAND U509 ( .A(n472), .B(n471), .Z(n128) );
endmodule

