
module stackMachine_N32 ( clk, rst, x, opcode, o );
  input [31:0] x;
  input [2:0] opcode;
  output [31:0] o;
  input clk, rst;
  wire   \stack[7][31] , \stack[7][30] , \stack[7][29] , \stack[7][28] ,
         \stack[7][27] , \stack[7][26] , \stack[7][25] , \stack[7][24] ,
         \stack[7][23] , \stack[7][22] , \stack[7][21] , \stack[7][20] ,
         \stack[7][19] , \stack[7][18] , \stack[7][17] , \stack[7][16] ,
         \stack[7][15] , \stack[7][14] , \stack[7][13] , \stack[7][12] ,
         \stack[7][11] , \stack[7][10] , \stack[7][9] , \stack[7][8] ,
         \stack[7][7] , \stack[7][6] , \stack[7][5] , \stack[7][4] ,
         \stack[7][3] , \stack[7][2] , \stack[7][1] , \stack[7][0] ,
         \stack[6][31] , \stack[6][30] , \stack[6][29] , \stack[6][28] ,
         \stack[6][27] , \stack[6][26] , \stack[6][25] , \stack[6][24] ,
         \stack[6][23] , \stack[6][22] , \stack[6][21] , \stack[6][20] ,
         \stack[6][19] , \stack[6][18] , \stack[6][17] , \stack[6][16] ,
         \stack[6][15] , \stack[6][14] , \stack[6][13] , \stack[6][12] ,
         \stack[6][11] , \stack[6][10] , \stack[6][9] , \stack[6][8] ,
         \stack[6][7] , \stack[6][6] , \stack[6][5] , \stack[6][4] ,
         \stack[6][3] , \stack[6][2] , \stack[6][1] , \stack[6][0] ,
         \stack[5][31] , \stack[5][30] , \stack[5][29] , \stack[5][28] ,
         \stack[5][27] , \stack[5][26] , \stack[5][25] , \stack[5][24] ,
         \stack[5][23] , \stack[5][22] , \stack[5][21] , \stack[5][20] ,
         \stack[5][19] , \stack[5][18] , \stack[5][17] , \stack[5][16] ,
         \stack[5][15] , \stack[5][14] , \stack[5][13] , \stack[5][12] ,
         \stack[5][11] , \stack[5][10] , \stack[5][9] , \stack[5][8] ,
         \stack[5][7] , \stack[5][6] , \stack[5][5] , \stack[5][4] ,
         \stack[5][3] , \stack[5][2] , \stack[5][1] , \stack[5][0] ,
         \stack[4][31] , \stack[4][30] , \stack[4][29] , \stack[4][28] ,
         \stack[4][27] , \stack[4][26] , \stack[4][25] , \stack[4][24] ,
         \stack[4][23] , \stack[4][22] , \stack[4][21] , \stack[4][20] ,
         \stack[4][19] , \stack[4][18] , \stack[4][17] , \stack[4][16] ,
         \stack[4][15] , \stack[4][14] , \stack[4][13] , \stack[4][12] ,
         \stack[4][11] , \stack[4][10] , \stack[4][9] , \stack[4][8] ,
         \stack[4][7] , \stack[4][6] , \stack[4][5] , \stack[4][4] ,
         \stack[4][3] , \stack[4][2] , \stack[4][1] , \stack[4][0] ,
         \stack[3][31] , \stack[3][30] , \stack[3][29] , \stack[3][28] ,
         \stack[3][27] , \stack[3][26] , \stack[3][25] , \stack[3][24] ,
         \stack[3][23] , \stack[3][22] , \stack[3][21] , \stack[3][20] ,
         \stack[3][19] , \stack[3][18] , \stack[3][17] , \stack[3][16] ,
         \stack[3][15] , \stack[3][14] , \stack[3][13] , \stack[3][12] ,
         \stack[3][11] , \stack[3][10] , \stack[3][9] , \stack[3][8] ,
         \stack[3][7] , \stack[3][6] , \stack[3][5] , \stack[3][4] ,
         \stack[3][3] , \stack[3][2] , \stack[3][1] , \stack[3][0] ,
         \stack[2][31] , \stack[2][30] , \stack[2][29] , \stack[2][28] ,
         \stack[2][27] , \stack[2][26] , \stack[2][25] , \stack[2][24] ,
         \stack[2][23] , \stack[2][22] , \stack[2][21] , \stack[2][20] ,
         \stack[2][19] , \stack[2][18] , \stack[2][17] , \stack[2][16] ,
         \stack[2][15] , \stack[2][14] , \stack[2][13] , \stack[2][12] ,
         \stack[2][11] , \stack[2][10] , \stack[2][9] , \stack[2][8] ,
         \stack[2][7] , \stack[2][6] , \stack[2][5] , \stack[2][4] ,
         \stack[2][3] , \stack[2][2] , \stack[2][1] , \stack[2][0] ,
         \stack[1][31] , \stack[1][30] , \stack[1][29] , \stack[1][28] ,
         \stack[1][27] , \stack[1][26] , \stack[1][25] , \stack[1][24] ,
         \stack[1][23] , \stack[1][22] , \stack[1][21] , \stack[1][20] ,
         \stack[1][19] , \stack[1][18] , \stack[1][17] , \stack[1][16] ,
         \stack[1][15] , \stack[1][14] , \stack[1][13] , \stack[1][12] ,
         \stack[1][11] , \stack[1][10] , \stack[1][9] , \stack[1][8] ,
         \stack[1][7] , \stack[1][6] , \stack[1][5] , \stack[1][4] ,
         \stack[1][3] , \stack[1][2] , \stack[1][1] , \stack[1][0] ,
         \C3/DATA5_0 , \C3/DATA5_1 , \C3/DATA5_2 , \C3/DATA5_3 , \C3/DATA5_4 ,
         \C3/DATA5_5 , \C3/DATA5_6 , \C3/DATA5_7 , \C3/DATA5_8 , \C3/DATA5_9 ,
         \C3/DATA5_10 , \C3/DATA5_11 , \C3/DATA5_12 , \C3/DATA5_13 ,
         \C3/DATA5_14 , \C3/DATA5_15 , \C3/DATA5_16 , \C3/DATA5_17 ,
         \C3/DATA5_18 , \C3/DATA5_19 , \C3/DATA5_20 , \C3/DATA5_21 ,
         \C3/DATA5_22 , \C3/DATA5_23 , \C3/DATA5_24 , \C3/DATA5_25 ,
         \C3/DATA5_26 , \C3/DATA5_27 , \C3/DATA5_28 , \C3/DATA5_29 ,
         \C3/DATA5_30 , \C3/DATA5_31 , n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, \C1/Z_0 , \U1/RSOP_16/C3/Z_31 , \U1/RSOP_16/C3/Z_30 ,
         \U1/RSOP_16/C3/Z_29 , \U1/RSOP_16/C3/Z_28 , \U1/RSOP_16/C3/Z_27 ,
         \U1/RSOP_16/C3/Z_26 , \U1/RSOP_16/C3/Z_25 , \U1/RSOP_16/C3/Z_24 ,
         \U1/RSOP_16/C3/Z_23 , \U1/RSOP_16/C3/Z_22 , \U1/RSOP_16/C3/Z_21 ,
         \U1/RSOP_16/C3/Z_20 , \U1/RSOP_16/C3/Z_19 , \U1/RSOP_16/C3/Z_18 ,
         \U1/RSOP_16/C3/Z_17 , \U1/RSOP_16/C3/Z_16 , \U1/RSOP_16/C3/Z_15 ,
         \U1/RSOP_16/C3/Z_14 , \U1/RSOP_16/C3/Z_13 , \U1/RSOP_16/C3/Z_12 ,
         \U1/RSOP_16/C3/Z_11 , \U1/RSOP_16/C3/Z_10 , \U1/RSOP_16/C3/Z_9 ,
         \U1/RSOP_16/C3/Z_8 , \U1/RSOP_16/C3/Z_7 , \U1/RSOP_16/C3/Z_6 ,
         \U1/RSOP_16/C3/Z_5 , \U1/RSOP_16/C3/Z_4 , \U1/RSOP_16/C3/Z_3 ,
         \U1/RSOP_16/C3/Z_2 , \U1/RSOP_16/C3/Z_1 , \U1/RSOP_16/C3/Z_0 ,
         \U1/RSOP_16/C2/Z_31 , \U1/RSOP_16/C2/Z_30 , \U1/RSOP_16/C2/Z_29 ,
         \U1/RSOP_16/C2/Z_28 , \U1/RSOP_16/C2/Z_27 , \U1/RSOP_16/C2/Z_26 ,
         \U1/RSOP_16/C2/Z_25 , \U1/RSOP_16/C2/Z_24 , \U1/RSOP_16/C2/Z_23 ,
         \U1/RSOP_16/C2/Z_22 , \U1/RSOP_16/C2/Z_21 , \U1/RSOP_16/C2/Z_20 ,
         \U1/RSOP_16/C2/Z_19 , \U1/RSOP_16/C2/Z_18 , \U1/RSOP_16/C2/Z_17 ,
         \U1/RSOP_16/C2/Z_16 , \U1/RSOP_16/C2/Z_15 , \U1/RSOP_16/C2/Z_14 ,
         \U1/RSOP_16/C2/Z_13 , \U1/RSOP_16/C2/Z_12 , \U1/RSOP_16/C2/Z_11 ,
         \U1/RSOP_16/C2/Z_10 , \U1/RSOP_16/C2/Z_9 , \U1/RSOP_16/C2/Z_8 ,
         \U1/RSOP_16/C2/Z_7 , \U1/RSOP_16/C2/Z_6 , \U1/RSOP_16/C2/Z_5 ,
         \U1/RSOP_16/C2/Z_4 , \U1/RSOP_16/C2/Z_3 , \U1/RSOP_16/C2/Z_2 ,
         \U1/RSOP_16/C2/Z_1 , \U1/RSOP_16/C2/Z_0 , \DP_OP_25_64_5665/n336 ,
         \DP_OP_25_64_5665/n335 , \DP_OP_25_64_5665/n334 ,
         \DP_OP_25_64_5665/n333 , \DP_OP_25_64_5665/n332 ,
         \DP_OP_25_64_5665/n331 , \DP_OP_25_64_5665/n330 ,
         \DP_OP_25_64_5665/n329 , \DP_OP_25_64_5665/n328 ,
         \DP_OP_25_64_5665/n327 , \DP_OP_25_64_5665/n326 ,
         \DP_OP_25_64_5665/n325 , \DP_OP_25_64_5665/n324 ,
         \DP_OP_25_64_5665/n323 , \DP_OP_25_64_5665/n322 ,
         \DP_OP_25_64_5665/n321 , \DP_OP_25_64_5665/n320 ,
         \DP_OP_25_64_5665/n319 , \DP_OP_25_64_5665/n318 ,
         \DP_OP_25_64_5665/n317 , \DP_OP_25_64_5665/n316 ,
         \DP_OP_25_64_5665/n315 , \DP_OP_25_64_5665/n314 ,
         \DP_OP_25_64_5665/n313 , \DP_OP_25_64_5665/n312 ,
         \DP_OP_25_64_5665/n311 , \DP_OP_25_64_5665/n310 ,
         \DP_OP_25_64_5665/n309 , \DP_OP_25_64_5665/n308 ,
         \DP_OP_25_64_5665/n307 , \DP_OP_25_64_5665/n306 ,
         \DP_OP_25_64_5665/n305 , \DP_OP_25_64_5665/n300 ,
         \DP_OP_25_64_5665/n299 , \DP_OP_25_64_5665/n298 ,
         \DP_OP_25_64_5665/n297 , \DP_OP_25_64_5665/n296 ,
         \DP_OP_25_64_5665/n295 , \DP_OP_25_64_5665/n294 ,
         \DP_OP_25_64_5665/n293 , \DP_OP_25_64_5665/n292 ,
         \DP_OP_25_64_5665/n291 , \DP_OP_25_64_5665/n290 ,
         \DP_OP_25_64_5665/n289 , \DP_OP_25_64_5665/n288 ,
         \DP_OP_25_64_5665/n287 , \DP_OP_25_64_5665/n286 ,
         \DP_OP_25_64_5665/n285 , \DP_OP_25_64_5665/n284 ,
         \DP_OP_25_64_5665/n283 , \DP_OP_25_64_5665/n282 ,
         \DP_OP_25_64_5665/n281 , \DP_OP_25_64_5665/n280 ,
         \DP_OP_25_64_5665/n279 , \DP_OP_25_64_5665/n278 ,
         \DP_OP_25_64_5665/n277 , \DP_OP_25_64_5665/n276 ,
         \DP_OP_25_64_5665/n275 , \DP_OP_25_64_5665/n274 ,
         \DP_OP_25_64_5665/n273 , \DP_OP_25_64_5665/n272 ,
         \DP_OP_25_64_5665/n271 , \DP_OP_25_64_5665/n270 ,
         \DP_OP_25_64_5665/n269 , \DP_OP_25_64_5665/n268 ,
         \DP_OP_25_64_5665/n267 , \DP_OP_25_64_5665/n266 ,
         \DP_OP_25_64_5665/n265 , \DP_OP_25_64_5665/n264 ,
         \DP_OP_25_64_5665/n263 , \DP_OP_25_64_5665/n262 ,
         \DP_OP_25_64_5665/n261 , \DP_OP_25_64_5665/n260 ,
         \DP_OP_25_64_5665/n259 , \DP_OP_25_64_5665/n258 ,
         \DP_OP_25_64_5665/n257 , \DP_OP_25_64_5665/n256 ,
         \DP_OP_25_64_5665/n255 , \DP_OP_25_64_5665/n254 ,
         \DP_OP_25_64_5665/n253 , \DP_OP_25_64_5665/n252 ,
         \DP_OP_25_64_5665/n251 , \DP_OP_25_64_5665/n250 ,
         \DP_OP_25_64_5665/n249 , \DP_OP_25_64_5665/n248 ,
         \DP_OP_25_64_5665/n247 , \DP_OP_25_64_5665/n246 ,
         \DP_OP_25_64_5665/n245 , \DP_OP_25_64_5665/n244 ,
         \DP_OP_25_64_5665/n243 , \DP_OP_25_64_5665/n242 ,
         \DP_OP_25_64_5665/n241 , \DP_OP_25_64_5665/n240 ,
         \DP_OP_25_64_5665/n239 , \DP_OP_25_64_5665/n238 ,
         \DP_OP_25_64_5665/n236 , \DP_OP_25_64_5665/n235 ,
         \DP_OP_25_64_5665/n229 , \DP_OP_25_64_5665/n228 ,
         \DP_OP_25_64_5665/n222 , \DP_OP_25_64_5665/n221 ,
         \DP_OP_25_64_5665/n215 , \DP_OP_25_64_5665/n214 ,
         \DP_OP_25_64_5665/n208 , \DP_OP_25_64_5665/n207 ,
         \DP_OP_25_64_5665/n201 , \DP_OP_25_64_5665/n200 ,
         \DP_OP_25_64_5665/n194 , \DP_OP_25_64_5665/n193 ,
         \DP_OP_25_64_5665/n187 , \DP_OP_25_64_5665/n186 ,
         \DP_OP_25_64_5665/n180 , \DP_OP_25_64_5665/n179 ,
         \DP_OP_25_64_5665/n173 , \DP_OP_25_64_5665/n172 ,
         \DP_OP_25_64_5665/n166 , \DP_OP_25_64_5665/n165 ,
         \DP_OP_25_64_5665/n159 , \DP_OP_25_64_5665/n158 ,
         \DP_OP_25_64_5665/n152 , \DP_OP_25_64_5665/n151 ,
         \DP_OP_25_64_5665/n145 , \DP_OP_25_64_5665/n144 ,
         \DP_OP_25_64_5665/n138 , \DP_OP_25_64_5665/n137 ,
         \DP_OP_25_64_5665/n131 , \DP_OP_25_64_5665/n130 ,
         \DP_OP_25_64_5665/n124 , \DP_OP_25_64_5665/n123 ,
         \DP_OP_25_64_5665/n117 , \DP_OP_25_64_5665/n116 ,
         \DP_OP_25_64_5665/n110 , \DP_OP_25_64_5665/n109 ,
         \DP_OP_25_64_5665/n103 , \DP_OP_25_64_5665/n102 ,
         \DP_OP_25_64_5665/n96 , \DP_OP_25_64_5665/n95 ,
         \DP_OP_25_64_5665/n89 , \DP_OP_25_64_5665/n88 ,
         \DP_OP_25_64_5665/n82 , \DP_OP_25_64_5665/n81 ,
         \DP_OP_25_64_5665/n57 , \DP_OP_25_64_5665/n56 ,
         \DP_OP_25_64_5665/n50 , \DP_OP_25_64_5665/n49 ,
         \DP_OP_25_64_5665/n43 , \DP_OP_25_64_5665/n42 ,
         \DP_OP_25_64_5665/n36 , \DP_OP_25_64_5665/n35 ,
         \DP_OP_25_64_5665/n29 , \DP_OP_25_64_5665/n28 ,
         \DP_OP_25_64_5665/n22 , \DP_OP_25_64_5665/n21 ,
         \DP_OP_25_64_5665/n15 , \DP_OP_25_64_5665/n14 , \DP_OP_25_64_5665/n8 ,
         \DP_OP_25_64_5665/n5 , n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675;

  DFF \stack_reg[0][0]  ( .D(n1320), .CLK(clk), .RST(rst), .Q(o[0]) );
  DFF \stack_reg[1][0]  ( .D(n1319), .CLK(clk), .RST(rst), .Q(\stack[1][0] )
         );
  DFF \stack_reg[0][1]  ( .D(n1318), .CLK(clk), .RST(rst), .Q(o[1]) );
  DFF \stack_reg[1][1]  ( .D(n1317), .CLK(clk), .RST(rst), .Q(\stack[1][1] )
         );
  DFF \stack_reg[2][1]  ( .D(n1316), .CLK(clk), .RST(rst), .Q(\stack[2][1] )
         );
  DFF \stack_reg[3][1]  ( .D(n1315), .CLK(clk), .RST(rst), .Q(\stack[3][1] )
         );
  DFF \stack_reg[4][1]  ( .D(n1314), .CLK(clk), .RST(rst), .Q(\stack[4][1] )
         );
  DFF \stack_reg[5][1]  ( .D(n1313), .CLK(clk), .RST(rst), .Q(\stack[5][1] )
         );
  DFF \stack_reg[6][1]  ( .D(n1312), .CLK(clk), .RST(rst), .Q(\stack[6][1] )
         );
  DFF \stack_reg[7][1]  ( .D(n1311), .CLK(clk), .RST(rst), .Q(\stack[7][1] )
         );
  DFF \stack_reg[0][2]  ( .D(n1310), .CLK(clk), .RST(rst), .Q(o[2]) );
  DFF \stack_reg[1][2]  ( .D(n1309), .CLK(clk), .RST(rst), .Q(\stack[1][2] )
         );
  DFF \stack_reg[2][2]  ( .D(n1308), .CLK(clk), .RST(rst), .Q(\stack[2][2] )
         );
  DFF \stack_reg[3][2]  ( .D(n1307), .CLK(clk), .RST(rst), .Q(\stack[3][2] )
         );
  DFF \stack_reg[4][2]  ( .D(n1306), .CLK(clk), .RST(rst), .Q(\stack[4][2] )
         );
  DFF \stack_reg[5][2]  ( .D(n1305), .CLK(clk), .RST(rst), .Q(\stack[5][2] )
         );
  DFF \stack_reg[6][2]  ( .D(n1304), .CLK(clk), .RST(rst), .Q(\stack[6][2] )
         );
  DFF \stack_reg[7][2]  ( .D(n1303), .CLK(clk), .RST(rst), .Q(\stack[7][2] )
         );
  DFF \stack_reg[0][3]  ( .D(n1302), .CLK(clk), .RST(rst), .Q(o[3]) );
  DFF \stack_reg[1][3]  ( .D(n1301), .CLK(clk), .RST(rst), .Q(\stack[1][3] )
         );
  DFF \stack_reg[2][3]  ( .D(n1300), .CLK(clk), .RST(rst), .Q(\stack[2][3] )
         );
  DFF \stack_reg[3][3]  ( .D(n1299), .CLK(clk), .RST(rst), .Q(\stack[3][3] )
         );
  DFF \stack_reg[4][3]  ( .D(n1298), .CLK(clk), .RST(rst), .Q(\stack[4][3] )
         );
  DFF \stack_reg[5][3]  ( .D(n1297), .CLK(clk), .RST(rst), .Q(\stack[5][3] )
         );
  DFF \stack_reg[6][3]  ( .D(n1296), .CLK(clk), .RST(rst), .Q(\stack[6][3] )
         );
  DFF \stack_reg[7][3]  ( .D(n1295), .CLK(clk), .RST(rst), .Q(\stack[7][3] )
         );
  DFF \stack_reg[0][4]  ( .D(n1294), .CLK(clk), .RST(rst), .Q(o[4]) );
  DFF \stack_reg[1][4]  ( .D(n1293), .CLK(clk), .RST(rst), .Q(\stack[1][4] )
         );
  DFF \stack_reg[2][4]  ( .D(n1292), .CLK(clk), .RST(rst), .Q(\stack[2][4] )
         );
  DFF \stack_reg[3][4]  ( .D(n1291), .CLK(clk), .RST(rst), .Q(\stack[3][4] )
         );
  DFF \stack_reg[4][4]  ( .D(n1290), .CLK(clk), .RST(rst), .Q(\stack[4][4] )
         );
  DFF \stack_reg[5][4]  ( .D(n1289), .CLK(clk), .RST(rst), .Q(\stack[5][4] )
         );
  DFF \stack_reg[6][4]  ( .D(n1288), .CLK(clk), .RST(rst), .Q(\stack[6][4] )
         );
  DFF \stack_reg[7][4]  ( .D(n1287), .CLK(clk), .RST(rst), .Q(\stack[7][4] )
         );
  DFF \stack_reg[0][5]  ( .D(n1286), .CLK(clk), .RST(rst), .Q(o[5]) );
  DFF \stack_reg[1][5]  ( .D(n1285), .CLK(clk), .RST(rst), .Q(\stack[1][5] )
         );
  DFF \stack_reg[2][5]  ( .D(n1284), .CLK(clk), .RST(rst), .Q(\stack[2][5] )
         );
  DFF \stack_reg[3][5]  ( .D(n1283), .CLK(clk), .RST(rst), .Q(\stack[3][5] )
         );
  DFF \stack_reg[4][5]  ( .D(n1282), .CLK(clk), .RST(rst), .Q(\stack[4][5] )
         );
  DFF \stack_reg[5][5]  ( .D(n1281), .CLK(clk), .RST(rst), .Q(\stack[5][5] )
         );
  DFF \stack_reg[6][5]  ( .D(n1280), .CLK(clk), .RST(rst), .Q(\stack[6][5] )
         );
  DFF \stack_reg[7][5]  ( .D(n1279), .CLK(clk), .RST(rst), .Q(\stack[7][5] )
         );
  DFF \stack_reg[0][6]  ( .D(n1278), .CLK(clk), .RST(rst), .Q(o[6]) );
  DFF \stack_reg[1][6]  ( .D(n1277), .CLK(clk), .RST(rst), .Q(\stack[1][6] )
         );
  DFF \stack_reg[2][6]  ( .D(n1276), .CLK(clk), .RST(rst), .Q(\stack[2][6] )
         );
  DFF \stack_reg[3][6]  ( .D(n1275), .CLK(clk), .RST(rst), .Q(\stack[3][6] )
         );
  DFF \stack_reg[4][6]  ( .D(n1274), .CLK(clk), .RST(rst), .Q(\stack[4][6] )
         );
  DFF \stack_reg[5][6]  ( .D(n1273), .CLK(clk), .RST(rst), .Q(\stack[5][6] )
         );
  DFF \stack_reg[6][6]  ( .D(n1272), .CLK(clk), .RST(rst), .Q(\stack[6][6] )
         );
  DFF \stack_reg[7][6]  ( .D(n1271), .CLK(clk), .RST(rst), .Q(\stack[7][6] )
         );
  DFF \stack_reg[0][7]  ( .D(n1270), .CLK(clk), .RST(rst), .Q(o[7]) );
  DFF \stack_reg[1][7]  ( .D(n1269), .CLK(clk), .RST(rst), .Q(\stack[1][7] )
         );
  DFF \stack_reg[2][7]  ( .D(n1268), .CLK(clk), .RST(rst), .Q(\stack[2][7] )
         );
  DFF \stack_reg[3][7]  ( .D(n1267), .CLK(clk), .RST(rst), .Q(\stack[3][7] )
         );
  DFF \stack_reg[4][7]  ( .D(n1266), .CLK(clk), .RST(rst), .Q(\stack[4][7] )
         );
  DFF \stack_reg[5][7]  ( .D(n1265), .CLK(clk), .RST(rst), .Q(\stack[5][7] )
         );
  DFF \stack_reg[6][7]  ( .D(n1264), .CLK(clk), .RST(rst), .Q(\stack[6][7] )
         );
  DFF \stack_reg[7][7]  ( .D(n1263), .CLK(clk), .RST(rst), .Q(\stack[7][7] )
         );
  DFF \stack_reg[0][8]  ( .D(n1262), .CLK(clk), .RST(rst), .Q(o[8]) );
  DFF \stack_reg[1][8]  ( .D(n1261), .CLK(clk), .RST(rst), .Q(\stack[1][8] )
         );
  DFF \stack_reg[2][8]  ( .D(n1260), .CLK(clk), .RST(rst), .Q(\stack[2][8] )
         );
  DFF \stack_reg[3][8]  ( .D(n1259), .CLK(clk), .RST(rst), .Q(\stack[3][8] )
         );
  DFF \stack_reg[4][8]  ( .D(n1258), .CLK(clk), .RST(rst), .Q(\stack[4][8] )
         );
  DFF \stack_reg[5][8]  ( .D(n1257), .CLK(clk), .RST(rst), .Q(\stack[5][8] )
         );
  DFF \stack_reg[6][8]  ( .D(n1256), .CLK(clk), .RST(rst), .Q(\stack[6][8] )
         );
  DFF \stack_reg[7][8]  ( .D(n1255), .CLK(clk), .RST(rst), .Q(\stack[7][8] )
         );
  DFF \stack_reg[0][9]  ( .D(n1254), .CLK(clk), .RST(rst), .Q(o[9]) );
  DFF \stack_reg[1][9]  ( .D(n1253), .CLK(clk), .RST(rst), .Q(\stack[1][9] )
         );
  DFF \stack_reg[2][9]  ( .D(n1252), .CLK(clk), .RST(rst), .Q(\stack[2][9] )
         );
  DFF \stack_reg[3][9]  ( .D(n1251), .CLK(clk), .RST(rst), .Q(\stack[3][9] )
         );
  DFF \stack_reg[4][9]  ( .D(n1250), .CLK(clk), .RST(rst), .Q(\stack[4][9] )
         );
  DFF \stack_reg[5][9]  ( .D(n1249), .CLK(clk), .RST(rst), .Q(\stack[5][9] )
         );
  DFF \stack_reg[6][9]  ( .D(n1248), .CLK(clk), .RST(rst), .Q(\stack[6][9] )
         );
  DFF \stack_reg[7][9]  ( .D(n1247), .CLK(clk), .RST(rst), .Q(\stack[7][9] )
         );
  DFF \stack_reg[0][10]  ( .D(n1246), .CLK(clk), .RST(rst), .Q(o[10]) );
  DFF \stack_reg[1][10]  ( .D(n1245), .CLK(clk), .RST(rst), .Q(\stack[1][10] )
         );
  DFF \stack_reg[2][10]  ( .D(n1244), .CLK(clk), .RST(rst), .Q(\stack[2][10] )
         );
  DFF \stack_reg[3][10]  ( .D(n1243), .CLK(clk), .RST(rst), .Q(\stack[3][10] )
         );
  DFF \stack_reg[4][10]  ( .D(n1242), .CLK(clk), .RST(rst), .Q(\stack[4][10] )
         );
  DFF \stack_reg[5][10]  ( .D(n1241), .CLK(clk), .RST(rst), .Q(\stack[5][10] )
         );
  DFF \stack_reg[6][10]  ( .D(n1240), .CLK(clk), .RST(rst), .Q(\stack[6][10] )
         );
  DFF \stack_reg[7][10]  ( .D(n1239), .CLK(clk), .RST(rst), .Q(\stack[7][10] )
         );
  DFF \stack_reg[0][11]  ( .D(n1238), .CLK(clk), .RST(rst), .Q(o[11]) );
  DFF \stack_reg[1][11]  ( .D(n1237), .CLK(clk), .RST(rst), .Q(\stack[1][11] )
         );
  DFF \stack_reg[2][11]  ( .D(n1236), .CLK(clk), .RST(rst), .Q(\stack[2][11] )
         );
  DFF \stack_reg[3][11]  ( .D(n1235), .CLK(clk), .RST(rst), .Q(\stack[3][11] )
         );
  DFF \stack_reg[4][11]  ( .D(n1234), .CLK(clk), .RST(rst), .Q(\stack[4][11] )
         );
  DFF \stack_reg[5][11]  ( .D(n1233), .CLK(clk), .RST(rst), .Q(\stack[5][11] )
         );
  DFF \stack_reg[6][11]  ( .D(n1232), .CLK(clk), .RST(rst), .Q(\stack[6][11] )
         );
  DFF \stack_reg[7][11]  ( .D(n1231), .CLK(clk), .RST(rst), .Q(\stack[7][11] )
         );
  DFF \stack_reg[0][12]  ( .D(n1230), .CLK(clk), .RST(rst), .Q(o[12]) );
  DFF \stack_reg[1][12]  ( .D(n1229), .CLK(clk), .RST(rst), .Q(\stack[1][12] )
         );
  DFF \stack_reg[2][12]  ( .D(n1228), .CLK(clk), .RST(rst), .Q(\stack[2][12] )
         );
  DFF \stack_reg[3][12]  ( .D(n1227), .CLK(clk), .RST(rst), .Q(\stack[3][12] )
         );
  DFF \stack_reg[4][12]  ( .D(n1226), .CLK(clk), .RST(rst), .Q(\stack[4][12] )
         );
  DFF \stack_reg[5][12]  ( .D(n1225), .CLK(clk), .RST(rst), .Q(\stack[5][12] )
         );
  DFF \stack_reg[6][12]  ( .D(n1224), .CLK(clk), .RST(rst), .Q(\stack[6][12] )
         );
  DFF \stack_reg[7][12]  ( .D(n1223), .CLK(clk), .RST(rst), .Q(\stack[7][12] )
         );
  DFF \stack_reg[0][13]  ( .D(n1222), .CLK(clk), .RST(rst), .Q(o[13]) );
  DFF \stack_reg[1][13]  ( .D(n1221), .CLK(clk), .RST(rst), .Q(\stack[1][13] )
         );
  DFF \stack_reg[2][13]  ( .D(n1220), .CLK(clk), .RST(rst), .Q(\stack[2][13] )
         );
  DFF \stack_reg[3][13]  ( .D(n1219), .CLK(clk), .RST(rst), .Q(\stack[3][13] )
         );
  DFF \stack_reg[4][13]  ( .D(n1218), .CLK(clk), .RST(rst), .Q(\stack[4][13] )
         );
  DFF \stack_reg[5][13]  ( .D(n1217), .CLK(clk), .RST(rst), .Q(\stack[5][13] )
         );
  DFF \stack_reg[6][13]  ( .D(n1216), .CLK(clk), .RST(rst), .Q(\stack[6][13] )
         );
  DFF \stack_reg[7][13]  ( .D(n1215), .CLK(clk), .RST(rst), .Q(\stack[7][13] )
         );
  DFF \stack_reg[0][14]  ( .D(n1214), .CLK(clk), .RST(rst), .Q(o[14]) );
  DFF \stack_reg[1][14]  ( .D(n1213), .CLK(clk), .RST(rst), .Q(\stack[1][14] )
         );
  DFF \stack_reg[2][14]  ( .D(n1212), .CLK(clk), .RST(rst), .Q(\stack[2][14] )
         );
  DFF \stack_reg[3][14]  ( .D(n1211), .CLK(clk), .RST(rst), .Q(\stack[3][14] )
         );
  DFF \stack_reg[4][14]  ( .D(n1210), .CLK(clk), .RST(rst), .Q(\stack[4][14] )
         );
  DFF \stack_reg[5][14]  ( .D(n1209), .CLK(clk), .RST(rst), .Q(\stack[5][14] )
         );
  DFF \stack_reg[6][14]  ( .D(n1208), .CLK(clk), .RST(rst), .Q(\stack[6][14] )
         );
  DFF \stack_reg[7][14]  ( .D(n1207), .CLK(clk), .RST(rst), .Q(\stack[7][14] )
         );
  DFF \stack_reg[0][15]  ( .D(n1206), .CLK(clk), .RST(rst), .Q(o[15]) );
  DFF \stack_reg[1][15]  ( .D(n1205), .CLK(clk), .RST(rst), .Q(\stack[1][15] )
         );
  DFF \stack_reg[2][15]  ( .D(n1204), .CLK(clk), .RST(rst), .Q(\stack[2][15] )
         );
  DFF \stack_reg[3][15]  ( .D(n1203), .CLK(clk), .RST(rst), .Q(\stack[3][15] )
         );
  DFF \stack_reg[4][15]  ( .D(n1202), .CLK(clk), .RST(rst), .Q(\stack[4][15] )
         );
  DFF \stack_reg[5][15]  ( .D(n1201), .CLK(clk), .RST(rst), .Q(\stack[5][15] )
         );
  DFF \stack_reg[6][15]  ( .D(n1200), .CLK(clk), .RST(rst), .Q(\stack[6][15] )
         );
  DFF \stack_reg[7][15]  ( .D(n1199), .CLK(clk), .RST(rst), .Q(\stack[7][15] )
         );
  DFF \stack_reg[0][16]  ( .D(n1198), .CLK(clk), .RST(rst), .Q(o[16]) );
  DFF \stack_reg[1][16]  ( .D(n1197), .CLK(clk), .RST(rst), .Q(\stack[1][16] )
         );
  DFF \stack_reg[2][16]  ( .D(n1196), .CLK(clk), .RST(rst), .Q(\stack[2][16] )
         );
  DFF \stack_reg[3][16]  ( .D(n1195), .CLK(clk), .RST(rst), .Q(\stack[3][16] )
         );
  DFF \stack_reg[4][16]  ( .D(n1194), .CLK(clk), .RST(rst), .Q(\stack[4][16] )
         );
  DFF \stack_reg[5][16]  ( .D(n1193), .CLK(clk), .RST(rst), .Q(\stack[5][16] )
         );
  DFF \stack_reg[6][16]  ( .D(n1192), .CLK(clk), .RST(rst), .Q(\stack[6][16] )
         );
  DFF \stack_reg[7][16]  ( .D(n1191), .CLK(clk), .RST(rst), .Q(\stack[7][16] )
         );
  DFF \stack_reg[0][17]  ( .D(n1190), .CLK(clk), .RST(rst), .Q(o[17]) );
  DFF \stack_reg[1][17]  ( .D(n1189), .CLK(clk), .RST(rst), .Q(\stack[1][17] )
         );
  DFF \stack_reg[2][17]  ( .D(n1188), .CLK(clk), .RST(rst), .Q(\stack[2][17] )
         );
  DFF \stack_reg[3][17]  ( .D(n1187), .CLK(clk), .RST(rst), .Q(\stack[3][17] )
         );
  DFF \stack_reg[4][17]  ( .D(n1186), .CLK(clk), .RST(rst), .Q(\stack[4][17] )
         );
  DFF \stack_reg[5][17]  ( .D(n1185), .CLK(clk), .RST(rst), .Q(\stack[5][17] )
         );
  DFF \stack_reg[6][17]  ( .D(n1184), .CLK(clk), .RST(rst), .Q(\stack[6][17] )
         );
  DFF \stack_reg[7][17]  ( .D(n1183), .CLK(clk), .RST(rst), .Q(\stack[7][17] )
         );
  DFF \stack_reg[0][18]  ( .D(n1182), .CLK(clk), .RST(rst), .Q(o[18]) );
  DFF \stack_reg[1][18]  ( .D(n1181), .CLK(clk), .RST(rst), .Q(\stack[1][18] )
         );
  DFF \stack_reg[2][18]  ( .D(n1180), .CLK(clk), .RST(rst), .Q(\stack[2][18] )
         );
  DFF \stack_reg[3][18]  ( .D(n1179), .CLK(clk), .RST(rst), .Q(\stack[3][18] )
         );
  DFF \stack_reg[4][18]  ( .D(n1178), .CLK(clk), .RST(rst), .Q(\stack[4][18] )
         );
  DFF \stack_reg[5][18]  ( .D(n1177), .CLK(clk), .RST(rst), .Q(\stack[5][18] )
         );
  DFF \stack_reg[6][18]  ( .D(n1176), .CLK(clk), .RST(rst), .Q(\stack[6][18] )
         );
  DFF \stack_reg[7][18]  ( .D(n1175), .CLK(clk), .RST(rst), .Q(\stack[7][18] )
         );
  DFF \stack_reg[0][19]  ( .D(n1174), .CLK(clk), .RST(rst), .Q(o[19]) );
  DFF \stack_reg[1][19]  ( .D(n1173), .CLK(clk), .RST(rst), .Q(\stack[1][19] )
         );
  DFF \stack_reg[2][19]  ( .D(n1172), .CLK(clk), .RST(rst), .Q(\stack[2][19] )
         );
  DFF \stack_reg[3][19]  ( .D(n1171), .CLK(clk), .RST(rst), .Q(\stack[3][19] )
         );
  DFF \stack_reg[4][19]  ( .D(n1170), .CLK(clk), .RST(rst), .Q(\stack[4][19] )
         );
  DFF \stack_reg[5][19]  ( .D(n1169), .CLK(clk), .RST(rst), .Q(\stack[5][19] )
         );
  DFF \stack_reg[6][19]  ( .D(n1168), .CLK(clk), .RST(rst), .Q(\stack[6][19] )
         );
  DFF \stack_reg[7][19]  ( .D(n1167), .CLK(clk), .RST(rst), .Q(\stack[7][19] )
         );
  DFF \stack_reg[0][20]  ( .D(n1166), .CLK(clk), .RST(rst), .Q(o[20]) );
  DFF \stack_reg[1][20]  ( .D(n1165), .CLK(clk), .RST(rst), .Q(\stack[1][20] )
         );
  DFF \stack_reg[2][20]  ( .D(n1164), .CLK(clk), .RST(rst), .Q(\stack[2][20] )
         );
  DFF \stack_reg[3][20]  ( .D(n1163), .CLK(clk), .RST(rst), .Q(\stack[3][20] )
         );
  DFF \stack_reg[4][20]  ( .D(n1162), .CLK(clk), .RST(rst), .Q(\stack[4][20] )
         );
  DFF \stack_reg[5][20]  ( .D(n1161), .CLK(clk), .RST(rst), .Q(\stack[5][20] )
         );
  DFF \stack_reg[6][20]  ( .D(n1160), .CLK(clk), .RST(rst), .Q(\stack[6][20] )
         );
  DFF \stack_reg[7][20]  ( .D(n1159), .CLK(clk), .RST(rst), .Q(\stack[7][20] )
         );
  DFF \stack_reg[0][21]  ( .D(n1158), .CLK(clk), .RST(rst), .Q(o[21]) );
  DFF \stack_reg[1][21]  ( .D(n1157), .CLK(clk), .RST(rst), .Q(\stack[1][21] )
         );
  DFF \stack_reg[2][21]  ( .D(n1156), .CLK(clk), .RST(rst), .Q(\stack[2][21] )
         );
  DFF \stack_reg[3][21]  ( .D(n1155), .CLK(clk), .RST(rst), .Q(\stack[3][21] )
         );
  DFF \stack_reg[4][21]  ( .D(n1154), .CLK(clk), .RST(rst), .Q(\stack[4][21] )
         );
  DFF \stack_reg[5][21]  ( .D(n1153), .CLK(clk), .RST(rst), .Q(\stack[5][21] )
         );
  DFF \stack_reg[6][21]  ( .D(n1152), .CLK(clk), .RST(rst), .Q(\stack[6][21] )
         );
  DFF \stack_reg[7][21]  ( .D(n1151), .CLK(clk), .RST(rst), .Q(\stack[7][21] )
         );
  DFF \stack_reg[0][22]  ( .D(n1150), .CLK(clk), .RST(rst), .Q(o[22]) );
  DFF \stack_reg[1][22]  ( .D(n1149), .CLK(clk), .RST(rst), .Q(\stack[1][22] )
         );
  DFF \stack_reg[2][22]  ( .D(n1148), .CLK(clk), .RST(rst), .Q(\stack[2][22] )
         );
  DFF \stack_reg[3][22]  ( .D(n1147), .CLK(clk), .RST(rst), .Q(\stack[3][22] )
         );
  DFF \stack_reg[4][22]  ( .D(n1146), .CLK(clk), .RST(rst), .Q(\stack[4][22] )
         );
  DFF \stack_reg[5][22]  ( .D(n1145), .CLK(clk), .RST(rst), .Q(\stack[5][22] )
         );
  DFF \stack_reg[6][22]  ( .D(n1144), .CLK(clk), .RST(rst), .Q(\stack[6][22] )
         );
  DFF \stack_reg[7][22]  ( .D(n1143), .CLK(clk), .RST(rst), .Q(\stack[7][22] )
         );
  DFF \stack_reg[0][23]  ( .D(n1142), .CLK(clk), .RST(rst), .Q(o[23]) );
  DFF \stack_reg[1][23]  ( .D(n1141), .CLK(clk), .RST(rst), .Q(\stack[1][23] )
         );
  DFF \stack_reg[2][23]  ( .D(n1140), .CLK(clk), .RST(rst), .Q(\stack[2][23] )
         );
  DFF \stack_reg[3][23]  ( .D(n1139), .CLK(clk), .RST(rst), .Q(\stack[3][23] )
         );
  DFF \stack_reg[4][23]  ( .D(n1138), .CLK(clk), .RST(rst), .Q(\stack[4][23] )
         );
  DFF \stack_reg[5][23]  ( .D(n1137), .CLK(clk), .RST(rst), .Q(\stack[5][23] )
         );
  DFF \stack_reg[6][23]  ( .D(n1136), .CLK(clk), .RST(rst), .Q(\stack[6][23] )
         );
  DFF \stack_reg[7][23]  ( .D(n1135), .CLK(clk), .RST(rst), .Q(\stack[7][23] )
         );
  DFF \stack_reg[0][24]  ( .D(n1134), .CLK(clk), .RST(rst), .Q(o[24]) );
  DFF \stack_reg[1][24]  ( .D(n1133), .CLK(clk), .RST(rst), .Q(\stack[1][24] )
         );
  DFF \stack_reg[2][24]  ( .D(n1132), .CLK(clk), .RST(rst), .Q(\stack[2][24] )
         );
  DFF \stack_reg[3][24]  ( .D(n1131), .CLK(clk), .RST(rst), .Q(\stack[3][24] )
         );
  DFF \stack_reg[4][24]  ( .D(n1130), .CLK(clk), .RST(rst), .Q(\stack[4][24] )
         );
  DFF \stack_reg[5][24]  ( .D(n1129), .CLK(clk), .RST(rst), .Q(\stack[5][24] )
         );
  DFF \stack_reg[6][24]  ( .D(n1128), .CLK(clk), .RST(rst), .Q(\stack[6][24] )
         );
  DFF \stack_reg[7][24]  ( .D(n1127), .CLK(clk), .RST(rst), .Q(\stack[7][24] )
         );
  DFF \stack_reg[0][25]  ( .D(n1126), .CLK(clk), .RST(rst), .Q(o[25]) );
  DFF \stack_reg[1][25]  ( .D(n1125), .CLK(clk), .RST(rst), .Q(\stack[1][25] )
         );
  DFF \stack_reg[2][25]  ( .D(n1124), .CLK(clk), .RST(rst), .Q(\stack[2][25] )
         );
  DFF \stack_reg[3][25]  ( .D(n1123), .CLK(clk), .RST(rst), .Q(\stack[3][25] )
         );
  DFF \stack_reg[4][25]  ( .D(n1122), .CLK(clk), .RST(rst), .Q(\stack[4][25] )
         );
  DFF \stack_reg[5][25]  ( .D(n1121), .CLK(clk), .RST(rst), .Q(\stack[5][25] )
         );
  DFF \stack_reg[6][25]  ( .D(n1120), .CLK(clk), .RST(rst), .Q(\stack[6][25] )
         );
  DFF \stack_reg[7][25]  ( .D(n1119), .CLK(clk), .RST(rst), .Q(\stack[7][25] )
         );
  DFF \stack_reg[0][26]  ( .D(n1118), .CLK(clk), .RST(rst), .Q(o[26]) );
  DFF \stack_reg[1][26]  ( .D(n1117), .CLK(clk), .RST(rst), .Q(\stack[1][26] )
         );
  DFF \stack_reg[2][26]  ( .D(n1116), .CLK(clk), .RST(rst), .Q(\stack[2][26] )
         );
  DFF \stack_reg[3][26]  ( .D(n1115), .CLK(clk), .RST(rst), .Q(\stack[3][26] )
         );
  DFF \stack_reg[4][26]  ( .D(n1114), .CLK(clk), .RST(rst), .Q(\stack[4][26] )
         );
  DFF \stack_reg[5][26]  ( .D(n1113), .CLK(clk), .RST(rst), .Q(\stack[5][26] )
         );
  DFF \stack_reg[6][26]  ( .D(n1112), .CLK(clk), .RST(rst), .Q(\stack[6][26] )
         );
  DFF \stack_reg[7][26]  ( .D(n1111), .CLK(clk), .RST(rst), .Q(\stack[7][26] )
         );
  DFF \stack_reg[0][27]  ( .D(n1110), .CLK(clk), .RST(rst), .Q(o[27]) );
  DFF \stack_reg[1][27]  ( .D(n1109), .CLK(clk), .RST(rst), .Q(\stack[1][27] )
         );
  DFF \stack_reg[2][27]  ( .D(n1108), .CLK(clk), .RST(rst), .Q(\stack[2][27] )
         );
  DFF \stack_reg[3][27]  ( .D(n1107), .CLK(clk), .RST(rst), .Q(\stack[3][27] )
         );
  DFF \stack_reg[4][27]  ( .D(n1106), .CLK(clk), .RST(rst), .Q(\stack[4][27] )
         );
  DFF \stack_reg[5][27]  ( .D(n1105), .CLK(clk), .RST(rst), .Q(\stack[5][27] )
         );
  DFF \stack_reg[6][27]  ( .D(n1104), .CLK(clk), .RST(rst), .Q(\stack[6][27] )
         );
  DFF \stack_reg[7][27]  ( .D(n1103), .CLK(clk), .RST(rst), .Q(\stack[7][27] )
         );
  DFF \stack_reg[0][28]  ( .D(n1102), .CLK(clk), .RST(rst), .Q(o[28]) );
  DFF \stack_reg[1][28]  ( .D(n1101), .CLK(clk), .RST(rst), .Q(\stack[1][28] )
         );
  DFF \stack_reg[2][28]  ( .D(n1100), .CLK(clk), .RST(rst), .Q(\stack[2][28] )
         );
  DFF \stack_reg[3][28]  ( .D(n1099), .CLK(clk), .RST(rst), .Q(\stack[3][28] )
         );
  DFF \stack_reg[4][28]  ( .D(n1098), .CLK(clk), .RST(rst), .Q(\stack[4][28] )
         );
  DFF \stack_reg[5][28]  ( .D(n1097), .CLK(clk), .RST(rst), .Q(\stack[5][28] )
         );
  DFF \stack_reg[6][28]  ( .D(n1096), .CLK(clk), .RST(rst), .Q(\stack[6][28] )
         );
  DFF \stack_reg[7][28]  ( .D(n1095), .CLK(clk), .RST(rst), .Q(\stack[7][28] )
         );
  DFF \stack_reg[0][29]  ( .D(n1094), .CLK(clk), .RST(rst), .Q(o[29]) );
  DFF \stack_reg[1][29]  ( .D(n1093), .CLK(clk), .RST(rst), .Q(\stack[1][29] )
         );
  DFF \stack_reg[2][29]  ( .D(n1092), .CLK(clk), .RST(rst), .Q(\stack[2][29] )
         );
  DFF \stack_reg[3][29]  ( .D(n1091), .CLK(clk), .RST(rst), .Q(\stack[3][29] )
         );
  DFF \stack_reg[4][29]  ( .D(n1090), .CLK(clk), .RST(rst), .Q(\stack[4][29] )
         );
  DFF \stack_reg[5][29]  ( .D(n1089), .CLK(clk), .RST(rst), .Q(\stack[5][29] )
         );
  DFF \stack_reg[6][29]  ( .D(n1088), .CLK(clk), .RST(rst), .Q(\stack[6][29] )
         );
  DFF \stack_reg[7][29]  ( .D(n1087), .CLK(clk), .RST(rst), .Q(\stack[7][29] )
         );
  DFF \stack_reg[0][30]  ( .D(n1086), .CLK(clk), .RST(rst), .Q(o[30]) );
  DFF \stack_reg[1][30]  ( .D(n1085), .CLK(clk), .RST(rst), .Q(\stack[1][30] )
         );
  DFF \stack_reg[2][30]  ( .D(n1084), .CLK(clk), .RST(rst), .Q(\stack[2][30] )
         );
  DFF \stack_reg[3][30]  ( .D(n1083), .CLK(clk), .RST(rst), .Q(\stack[3][30] )
         );
  DFF \stack_reg[4][30]  ( .D(n1082), .CLK(clk), .RST(rst), .Q(\stack[4][30] )
         );
  DFF \stack_reg[5][30]  ( .D(n1081), .CLK(clk), .RST(rst), .Q(\stack[5][30] )
         );
  DFF \stack_reg[6][30]  ( .D(n1080), .CLK(clk), .RST(rst), .Q(\stack[6][30] )
         );
  DFF \stack_reg[7][30]  ( .D(n1079), .CLK(clk), .RST(rst), .Q(\stack[7][30] )
         );
  DFF \stack_reg[0][31]  ( .D(n1078), .CLK(clk), .RST(rst), .Q(o[31]) );
  DFF \stack_reg[1][31]  ( .D(n1077), .CLK(clk), .RST(rst), .Q(\stack[1][31] )
         );
  DFF \stack_reg[2][31]  ( .D(n1076), .CLK(clk), .RST(rst), .Q(\stack[2][31] )
         );
  DFF \stack_reg[3][31]  ( .D(n1075), .CLK(clk), .RST(rst), .Q(\stack[3][31] )
         );
  DFF \stack_reg[4][31]  ( .D(n1074), .CLK(clk), .RST(rst), .Q(\stack[4][31] )
         );
  DFF \stack_reg[5][31]  ( .D(n1073), .CLK(clk), .RST(rst), .Q(\stack[5][31] )
         );
  DFF \stack_reg[6][31]  ( .D(n1072), .CLK(clk), .RST(rst), .Q(\stack[6][31] )
         );
  DFF \stack_reg[7][31]  ( .D(n1071), .CLK(clk), .RST(rst), .Q(\stack[7][31] )
         );
  DFF \stack_reg[2][0]  ( .D(n1070), .CLK(clk), .RST(rst), .Q(\stack[2][0] )
         );
  DFF \stack_reg[3][0]  ( .D(n1069), .CLK(clk), .RST(rst), .Q(\stack[3][0] )
         );
  DFF \stack_reg[4][0]  ( .D(n1068), .CLK(clk), .RST(rst), .Q(\stack[4][0] )
         );
  DFF \stack_reg[5][0]  ( .D(n1067), .CLK(clk), .RST(rst), .Q(\stack[5][0] )
         );
  DFF \stack_reg[6][0]  ( .D(n1066), .CLK(clk), .RST(rst), .Q(\stack[6][0] )
         );
  DFF \stack_reg[7][0]  ( .D(n1065), .CLK(clk), .RST(rst), .Q(\stack[7][0] )
         );
  XOR \DP_OP_25_64_5665/U149  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_0 ), .Z(
        \DP_OP_25_64_5665/n336 ) );
  XOR \DP_OP_25_64_5665/U148  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_1 ), .Z(
        \DP_OP_25_64_5665/n335 ) );
  XOR \DP_OP_25_64_5665/U147  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_2 ), .Z(
        \DP_OP_25_64_5665/n334 ) );
  XOR \DP_OP_25_64_5665/U146  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_3 ), .Z(
        \DP_OP_25_64_5665/n333 ) );
  XOR \DP_OP_25_64_5665/U145  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_4 ), .Z(
        \DP_OP_25_64_5665/n332 ) );
  XOR \DP_OP_25_64_5665/U144  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_5 ), .Z(
        \DP_OP_25_64_5665/n331 ) );
  XOR \DP_OP_25_64_5665/U143  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_6 ), .Z(
        \DP_OP_25_64_5665/n330 ) );
  XOR \DP_OP_25_64_5665/U142  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_7 ), .Z(
        \DP_OP_25_64_5665/n329 ) );
  XOR \DP_OP_25_64_5665/U141  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_8 ), .Z(
        \DP_OP_25_64_5665/n328 ) );
  XOR \DP_OP_25_64_5665/U140  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_9 ), .Z(
        \DP_OP_25_64_5665/n327 ) );
  XOR \DP_OP_25_64_5665/U139  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_10 ), .Z(
        \DP_OP_25_64_5665/n326 ) );
  XOR \DP_OP_25_64_5665/U138  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_11 ), .Z(
        \DP_OP_25_64_5665/n325 ) );
  XOR \DP_OP_25_64_5665/U137  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_12 ), .Z(
        \DP_OP_25_64_5665/n324 ) );
  XOR \DP_OP_25_64_5665/U136  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_13 ), .Z(
        \DP_OP_25_64_5665/n323 ) );
  XOR \DP_OP_25_64_5665/U135  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_14 ), .Z(
        \DP_OP_25_64_5665/n322 ) );
  XOR \DP_OP_25_64_5665/U134  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_15 ), .Z(
        \DP_OP_25_64_5665/n321 ) );
  XOR \DP_OP_25_64_5665/U133  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_16 ), .Z(
        \DP_OP_25_64_5665/n320 ) );
  XOR \DP_OP_25_64_5665/U132  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_17 ), .Z(
        \DP_OP_25_64_5665/n319 ) );
  XOR \DP_OP_25_64_5665/U131  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_18 ), .Z(
        \DP_OP_25_64_5665/n318 ) );
  XOR \DP_OP_25_64_5665/U109  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_19 ), .Z(
        \DP_OP_25_64_5665/n317 ) );
  XOR \DP_OP_25_64_5665/U108  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_20 ), .Z(
        \DP_OP_25_64_5665/n316 ) );
  XOR \DP_OP_25_64_5665/U107  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_21 ), .Z(
        \DP_OP_25_64_5665/n315 ) );
  XOR \DP_OP_25_64_5665/U106  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_22 ), .Z(
        \DP_OP_25_64_5665/n314 ) );
  XOR \DP_OP_25_64_5665/U105  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_23 ), .Z(
        \DP_OP_25_64_5665/n313 ) );
  XOR \DP_OP_25_64_5665/U104  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_24 ), .Z(
        \DP_OP_25_64_5665/n312 ) );
  XOR \DP_OP_25_64_5665/U103  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_25 ), .Z(
        \DP_OP_25_64_5665/n311 ) );
  XOR \DP_OP_25_64_5665/U102  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_26 ), .Z(
        \DP_OP_25_64_5665/n310 ) );
  XOR \DP_OP_25_64_5665/U101  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_27 ), .Z(
        \DP_OP_25_64_5665/n309 ) );
  XOR \DP_OP_25_64_5665/U100  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_28 ), .Z(
        \DP_OP_25_64_5665/n308 ) );
  XOR \DP_OP_25_64_5665/U99  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_29 ), .Z(
        \DP_OP_25_64_5665/n307 ) );
  XOR \DP_OP_25_64_5665/U98  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_30 ), .Z(
        \DP_OP_25_64_5665/n306 ) );
  XOR \DP_OP_25_64_5665/U97  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_31 ), .Z(
        \DP_OP_25_64_5665/n305 ) );
  XOR \DP_OP_25_64_5665/U94  ( .A(\U1/RSOP_16/C2/Z_0 ), .B(\C1/Z_0 ), .Z(
        \DP_OP_25_64_5665/n269 ) );
  XOR \DP_OP_25_64_5665/U93  ( .A(\DP_OP_25_64_5665/n269 ), .B(
        \DP_OP_25_64_5665/n336 ), .Z(\C3/DATA5_0 ) );
  XOR \DP_OP_25_64_5665/U92  ( .A(\DP_OP_25_64_5665/n335 ), .B(
        \U1/RSOP_16/C2/Z_1 ), .Z(\DP_OP_25_64_5665/n268 ) );
  XOR \DP_OP_25_64_5665/U91  ( .A(\DP_OP_25_64_5665/n300 ), .B(
        \DP_OP_25_64_5665/n268 ), .Z(\C3/DATA5_1 ) );
  XOR \DP_OP_25_64_5665/U90  ( .A(\DP_OP_25_64_5665/n334 ), .B(
        \U1/RSOP_16/C2/Z_2 ), .Z(\DP_OP_25_64_5665/n267 ) );
  XOR \DP_OP_25_64_5665/U89  ( .A(\DP_OP_25_64_5665/n299 ), .B(
        \DP_OP_25_64_5665/n267 ), .Z(\C3/DATA5_2 ) );
  XOR \DP_OP_25_64_5665/U88  ( .A(\DP_OP_25_64_5665/n333 ), .B(
        \U1/RSOP_16/C2/Z_3 ), .Z(\DP_OP_25_64_5665/n266 ) );
  XOR \DP_OP_25_64_5665/U87  ( .A(\DP_OP_25_64_5665/n298 ), .B(
        \DP_OP_25_64_5665/n266 ), .Z(\C3/DATA5_3 ) );
  XOR \DP_OP_25_64_5665/U86  ( .A(\DP_OP_25_64_5665/n332 ), .B(
        \U1/RSOP_16/C2/Z_4 ), .Z(\DP_OP_25_64_5665/n265 ) );
  XOR \DP_OP_25_64_5665/U85  ( .A(\DP_OP_25_64_5665/n297 ), .B(
        \DP_OP_25_64_5665/n265 ), .Z(\C3/DATA5_4 ) );
  XOR \DP_OP_25_64_5665/U84  ( .A(\DP_OP_25_64_5665/n331 ), .B(
        \U1/RSOP_16/C2/Z_5 ), .Z(\DP_OP_25_64_5665/n264 ) );
  XOR \DP_OP_25_64_5665/U83  ( .A(\DP_OP_25_64_5665/n296 ), .B(
        \DP_OP_25_64_5665/n264 ), .Z(\C3/DATA5_5 ) );
  XOR \DP_OP_25_64_5665/U82  ( .A(\DP_OP_25_64_5665/n330 ), .B(
        \U1/RSOP_16/C2/Z_6 ), .Z(\DP_OP_25_64_5665/n263 ) );
  XOR \DP_OP_25_64_5665/U81  ( .A(\DP_OP_25_64_5665/n295 ), .B(
        \DP_OP_25_64_5665/n263 ), .Z(\C3/DATA5_6 ) );
  XOR \DP_OP_25_64_5665/U80  ( .A(\DP_OP_25_64_5665/n329 ), .B(
        \U1/RSOP_16/C2/Z_7 ), .Z(\DP_OP_25_64_5665/n262 ) );
  XOR \DP_OP_25_64_5665/U79  ( .A(\DP_OP_25_64_5665/n294 ), .B(
        \DP_OP_25_64_5665/n262 ), .Z(\C3/DATA5_7 ) );
  XOR \DP_OP_25_64_5665/U78  ( .A(\DP_OP_25_64_5665/n328 ), .B(
        \U1/RSOP_16/C2/Z_8 ), .Z(\DP_OP_25_64_5665/n261 ) );
  XOR \DP_OP_25_64_5665/U77  ( .A(\DP_OP_25_64_5665/n293 ), .B(
        \DP_OP_25_64_5665/n261 ), .Z(\C3/DATA5_8 ) );
  XOR \DP_OP_25_64_5665/U76  ( .A(\DP_OP_25_64_5665/n327 ), .B(
        \U1/RSOP_16/C2/Z_9 ), .Z(\DP_OP_25_64_5665/n260 ) );
  XOR \DP_OP_25_64_5665/U75  ( .A(\DP_OP_25_64_5665/n292 ), .B(
        \DP_OP_25_64_5665/n260 ), .Z(\C3/DATA5_9 ) );
  XOR \DP_OP_25_64_5665/U74  ( .A(\DP_OP_25_64_5665/n326 ), .B(
        \U1/RSOP_16/C2/Z_10 ), .Z(\DP_OP_25_64_5665/n259 ) );
  XOR \DP_OP_25_64_5665/U73  ( .A(\DP_OP_25_64_5665/n291 ), .B(
        \DP_OP_25_64_5665/n259 ), .Z(\C3/DATA5_10 ) );
  XOR \DP_OP_25_64_5665/U72  ( .A(\DP_OP_25_64_5665/n325 ), .B(
        \U1/RSOP_16/C2/Z_11 ), .Z(\DP_OP_25_64_5665/n258 ) );
  XOR \DP_OP_25_64_5665/U71  ( .A(\DP_OP_25_64_5665/n290 ), .B(
        \DP_OP_25_64_5665/n258 ), .Z(\C3/DATA5_11 ) );
  XOR \DP_OP_25_64_5665/U70  ( .A(\DP_OP_25_64_5665/n324 ), .B(
        \U1/RSOP_16/C2/Z_12 ), .Z(\DP_OP_25_64_5665/n257 ) );
  XOR \DP_OP_25_64_5665/U69  ( .A(\DP_OP_25_64_5665/n289 ), .B(
        \DP_OP_25_64_5665/n257 ), .Z(\C3/DATA5_12 ) );
  XOR \DP_OP_25_64_5665/U68  ( .A(\DP_OP_25_64_5665/n323 ), .B(
        \U1/RSOP_16/C2/Z_13 ), .Z(\DP_OP_25_64_5665/n256 ) );
  XOR \DP_OP_25_64_5665/U67  ( .A(\DP_OP_25_64_5665/n288 ), .B(
        \DP_OP_25_64_5665/n256 ), .Z(\C3/DATA5_13 ) );
  XOR \DP_OP_25_64_5665/U66  ( .A(\DP_OP_25_64_5665/n322 ), .B(
        \U1/RSOP_16/C2/Z_14 ), .Z(\DP_OP_25_64_5665/n255 ) );
  XOR \DP_OP_25_64_5665/U65  ( .A(\DP_OP_25_64_5665/n287 ), .B(
        \DP_OP_25_64_5665/n255 ), .Z(\C3/DATA5_14 ) );
  XOR \DP_OP_25_64_5665/U64  ( .A(\DP_OP_25_64_5665/n321 ), .B(
        \U1/RSOP_16/C2/Z_15 ), .Z(\DP_OP_25_64_5665/n254 ) );
  XOR \DP_OP_25_64_5665/U63  ( .A(\DP_OP_25_64_5665/n286 ), .B(
        \DP_OP_25_64_5665/n254 ), .Z(\C3/DATA5_15 ) );
  XOR \DP_OP_25_64_5665/U62  ( .A(\DP_OP_25_64_5665/n320 ), .B(
        \U1/RSOP_16/C2/Z_16 ), .Z(\DP_OP_25_64_5665/n253 ) );
  XOR \DP_OP_25_64_5665/U61  ( .A(\DP_OP_25_64_5665/n285 ), .B(
        \DP_OP_25_64_5665/n253 ), .Z(\C3/DATA5_16 ) );
  XOR \DP_OP_25_64_5665/U60  ( .A(\DP_OP_25_64_5665/n319 ), .B(
        \U1/RSOP_16/C2/Z_17 ), .Z(\DP_OP_25_64_5665/n252 ) );
  XOR \DP_OP_25_64_5665/U59  ( .A(\DP_OP_25_64_5665/n284 ), .B(
        \DP_OP_25_64_5665/n252 ), .Z(\C3/DATA5_17 ) );
  XOR \DP_OP_25_64_5665/U58  ( .A(\DP_OP_25_64_5665/n318 ), .B(
        \U1/RSOP_16/C2/Z_18 ), .Z(\DP_OP_25_64_5665/n251 ) );
  XOR \DP_OP_25_64_5665/U57  ( .A(\DP_OP_25_64_5665/n283 ), .B(
        \DP_OP_25_64_5665/n251 ), .Z(\C3/DATA5_18 ) );
  XOR \DP_OP_25_64_5665/U56  ( .A(\DP_OP_25_64_5665/n317 ), .B(
        \U1/RSOP_16/C2/Z_19 ), .Z(\DP_OP_25_64_5665/n250 ) );
  XOR \DP_OP_25_64_5665/U55  ( .A(\DP_OP_25_64_5665/n282 ), .B(
        \DP_OP_25_64_5665/n250 ), .Z(\C3/DATA5_19 ) );
  XOR \DP_OP_25_64_5665/U54  ( .A(\DP_OP_25_64_5665/n316 ), .B(
        \U1/RSOP_16/C2/Z_20 ), .Z(\DP_OP_25_64_5665/n249 ) );
  XOR \DP_OP_25_64_5665/U53  ( .A(\DP_OP_25_64_5665/n281 ), .B(
        \DP_OP_25_64_5665/n249 ), .Z(\C3/DATA5_20 ) );
  XOR \DP_OP_25_64_5665/U52  ( .A(\DP_OP_25_64_5665/n315 ), .B(
        \U1/RSOP_16/C2/Z_21 ), .Z(\DP_OP_25_64_5665/n248 ) );
  XOR \DP_OP_25_64_5665/U51  ( .A(\DP_OP_25_64_5665/n280 ), .B(
        \DP_OP_25_64_5665/n248 ), .Z(\C3/DATA5_21 ) );
  XOR \DP_OP_25_64_5665/U50  ( .A(\DP_OP_25_64_5665/n314 ), .B(
        \U1/RSOP_16/C2/Z_22 ), .Z(\DP_OP_25_64_5665/n247 ) );
  XOR \DP_OP_25_64_5665/U49  ( .A(\DP_OP_25_64_5665/n279 ), .B(
        \DP_OP_25_64_5665/n247 ), .Z(\C3/DATA5_22 ) );
  XOR \DP_OP_25_64_5665/U48  ( .A(\DP_OP_25_64_5665/n313 ), .B(
        \U1/RSOP_16/C2/Z_23 ), .Z(\DP_OP_25_64_5665/n246 ) );
  XOR \DP_OP_25_64_5665/U47  ( .A(\DP_OP_25_64_5665/n278 ), .B(
        \DP_OP_25_64_5665/n246 ), .Z(\C3/DATA5_23 ) );
  XOR \DP_OP_25_64_5665/U46  ( .A(\DP_OP_25_64_5665/n312 ), .B(
        \U1/RSOP_16/C2/Z_24 ), .Z(\DP_OP_25_64_5665/n245 ) );
  XOR \DP_OP_25_64_5665/U45  ( .A(\DP_OP_25_64_5665/n277 ), .B(
        \DP_OP_25_64_5665/n245 ), .Z(\C3/DATA5_24 ) );
  XOR \DP_OP_25_64_5665/U44  ( .A(\DP_OP_25_64_5665/n311 ), .B(
        \U1/RSOP_16/C2/Z_25 ), .Z(\DP_OP_25_64_5665/n244 ) );
  XOR \DP_OP_25_64_5665/U43  ( .A(\DP_OP_25_64_5665/n276 ), .B(
        \DP_OP_25_64_5665/n244 ), .Z(\C3/DATA5_25 ) );
  XOR \DP_OP_25_64_5665/U42  ( .A(\DP_OP_25_64_5665/n310 ), .B(
        \U1/RSOP_16/C2/Z_26 ), .Z(\DP_OP_25_64_5665/n243 ) );
  XOR \DP_OP_25_64_5665/U41  ( .A(\DP_OP_25_64_5665/n275 ), .B(
        \DP_OP_25_64_5665/n243 ), .Z(\C3/DATA5_26 ) );
  XOR \DP_OP_25_64_5665/U40  ( .A(\DP_OP_25_64_5665/n309 ), .B(
        \U1/RSOP_16/C2/Z_27 ), .Z(\DP_OP_25_64_5665/n242 ) );
  XOR \DP_OP_25_64_5665/U30  ( .A(\DP_OP_25_64_5665/n274 ), .B(
        \DP_OP_25_64_5665/n242 ), .Z(\C3/DATA5_27 ) );
  XOR \DP_OP_25_64_5665/U20  ( .A(\DP_OP_25_64_5665/n308 ), .B(
        \U1/RSOP_16/C2/Z_28 ), .Z(\DP_OP_25_64_5665/n241 ) );
  XOR \DP_OP_25_64_5665/U10  ( .A(\DP_OP_25_64_5665/n273 ), .B(
        \DP_OP_25_64_5665/n241 ), .Z(\C3/DATA5_28 ) );
  XOR \DP_OP_25_64_5665/U9  ( .A(\DP_OP_25_64_5665/n307 ), .B(
        \U1/RSOP_16/C2/Z_29 ), .Z(\DP_OP_25_64_5665/n240 ) );
  XOR \DP_OP_25_64_5665/U8  ( .A(\DP_OP_25_64_5665/n272 ), .B(
        \DP_OP_25_64_5665/n240 ), .Z(\C3/DATA5_29 ) );
  XOR \DP_OP_25_64_5665/U7  ( .A(\DP_OP_25_64_5665/n306 ), .B(
        \U1/RSOP_16/C2/Z_30 ), .Z(\DP_OP_25_64_5665/n239 ) );
  XOR \DP_OP_25_64_5665/U6  ( .A(\DP_OP_25_64_5665/n271 ), .B(
        \DP_OP_25_64_5665/n239 ), .Z(\C3/DATA5_30 ) );
  XOR \DP_OP_25_64_5665/U5  ( .A(\DP_OP_25_64_5665/n305 ), .B(
        \U1/RSOP_16/C2/Z_31 ), .Z(\DP_OP_25_64_5665/n238 ) );
  XOR \DP_OP_25_64_5665/U4  ( .A(\DP_OP_25_64_5665/n270 ), .B(
        \DP_OP_25_64_5665/n238 ), .Z(\C3/DATA5_31 ) );
  NAND \DP_OP_25_64_5665/U130  ( .A(\DP_OP_25_64_5665/n306 ), .B(
        \U1/RSOP_16/C2/Z_30 ), .Z(\DP_OP_25_64_5665/n5 ) );
  NAND \DP_OP_25_64_5665/U230  ( .A(\DP_OP_25_64_5665/n271 ), .B(
        \DP_OP_25_64_5665/n239 ), .Z(\DP_OP_25_64_5665/n8 ) );
  NAND \DP_OP_25_64_5665/U330  ( .A(\DP_OP_25_64_5665/n5 ), .B(
        \DP_OP_25_64_5665/n8 ), .Z(\DP_OP_25_64_5665/n270 ) );
  NAND \DP_OP_25_64_5665/U129  ( .A(\DP_OP_25_64_5665/n307 ), .B(
        \U1/RSOP_16/C2/Z_29 ), .Z(\DP_OP_25_64_5665/n14 ) );
  NAND \DP_OP_25_64_5665/U229  ( .A(\DP_OP_25_64_5665/n272 ), .B(
        \DP_OP_25_64_5665/n240 ), .Z(\DP_OP_25_64_5665/n15 ) );
  NAND \DP_OP_25_64_5665/U329  ( .A(\DP_OP_25_64_5665/n14 ), .B(
        \DP_OP_25_64_5665/n15 ), .Z(\DP_OP_25_64_5665/n271 ) );
  NAND \DP_OP_25_64_5665/U128  ( .A(\DP_OP_25_64_5665/n308 ), .B(
        \U1/RSOP_16/C2/Z_28 ), .Z(\DP_OP_25_64_5665/n21 ) );
  NAND \DP_OP_25_64_5665/U228  ( .A(\DP_OP_25_64_5665/n273 ), .B(
        \DP_OP_25_64_5665/n241 ), .Z(\DP_OP_25_64_5665/n22 ) );
  NAND \DP_OP_25_64_5665/U328  ( .A(\DP_OP_25_64_5665/n21 ), .B(
        \DP_OP_25_64_5665/n22 ), .Z(\DP_OP_25_64_5665/n272 ) );
  NAND \DP_OP_25_64_5665/U127  ( .A(\DP_OP_25_64_5665/n309 ), .B(
        \U1/RSOP_16/C2/Z_27 ), .Z(\DP_OP_25_64_5665/n28 ) );
  NAND \DP_OP_25_64_5665/U227  ( .A(\DP_OP_25_64_5665/n274 ), .B(
        \DP_OP_25_64_5665/n242 ), .Z(\DP_OP_25_64_5665/n29 ) );
  NAND \DP_OP_25_64_5665/U327  ( .A(\DP_OP_25_64_5665/n28 ), .B(
        \DP_OP_25_64_5665/n29 ), .Z(\DP_OP_25_64_5665/n273 ) );
  NAND \DP_OP_25_64_5665/U126  ( .A(\DP_OP_25_64_5665/n310 ), .B(
        \U1/RSOP_16/C2/Z_26 ), .Z(\DP_OP_25_64_5665/n35 ) );
  NAND \DP_OP_25_64_5665/U226  ( .A(\DP_OP_25_64_5665/n275 ), .B(
        \DP_OP_25_64_5665/n243 ), .Z(\DP_OP_25_64_5665/n36 ) );
  NAND \DP_OP_25_64_5665/U326  ( .A(\DP_OP_25_64_5665/n35 ), .B(
        \DP_OP_25_64_5665/n36 ), .Z(\DP_OP_25_64_5665/n274 ) );
  NAND \DP_OP_25_64_5665/U125  ( .A(\DP_OP_25_64_5665/n311 ), .B(
        \U1/RSOP_16/C2/Z_25 ), .Z(\DP_OP_25_64_5665/n42 ) );
  NAND \DP_OP_25_64_5665/U225  ( .A(\DP_OP_25_64_5665/n276 ), .B(
        \DP_OP_25_64_5665/n244 ), .Z(\DP_OP_25_64_5665/n43 ) );
  NAND \DP_OP_25_64_5665/U325  ( .A(\DP_OP_25_64_5665/n42 ), .B(
        \DP_OP_25_64_5665/n43 ), .Z(\DP_OP_25_64_5665/n275 ) );
  NAND \DP_OP_25_64_5665/U124  ( .A(\DP_OP_25_64_5665/n312 ), .B(
        \U1/RSOP_16/C2/Z_24 ), .Z(\DP_OP_25_64_5665/n49 ) );
  NAND \DP_OP_25_64_5665/U224  ( .A(\DP_OP_25_64_5665/n277 ), .B(
        \DP_OP_25_64_5665/n245 ), .Z(\DP_OP_25_64_5665/n50 ) );
  NAND \DP_OP_25_64_5665/U324  ( .A(\DP_OP_25_64_5665/n49 ), .B(
        \DP_OP_25_64_5665/n50 ), .Z(\DP_OP_25_64_5665/n276 ) );
  NAND \DP_OP_25_64_5665/U123  ( .A(\DP_OP_25_64_5665/n313 ), .B(
        \U1/RSOP_16/C2/Z_23 ), .Z(\DP_OP_25_64_5665/n56 ) );
  NAND \DP_OP_25_64_5665/U223  ( .A(\DP_OP_25_64_5665/n278 ), .B(
        \DP_OP_25_64_5665/n246 ), .Z(\DP_OP_25_64_5665/n57 ) );
  NAND \DP_OP_25_64_5665/U323  ( .A(\DP_OP_25_64_5665/n56 ), .B(
        \DP_OP_25_64_5665/n57 ), .Z(\DP_OP_25_64_5665/n277 ) );
  NAND \DP_OP_25_64_5665/U122  ( .A(\DP_OP_25_64_5665/n314 ), .B(
        \U1/RSOP_16/C2/Z_22 ), .Z(\DP_OP_25_64_5665/n81 ) );
  NAND \DP_OP_25_64_5665/U222  ( .A(\DP_OP_25_64_5665/n279 ), .B(
        \DP_OP_25_64_5665/n247 ), .Z(\DP_OP_25_64_5665/n82 ) );
  NAND \DP_OP_25_64_5665/U322  ( .A(\DP_OP_25_64_5665/n81 ), .B(
        \DP_OP_25_64_5665/n82 ), .Z(\DP_OP_25_64_5665/n278 ) );
  NAND \DP_OP_25_64_5665/U121  ( .A(\DP_OP_25_64_5665/n315 ), .B(
        \U1/RSOP_16/C2/Z_21 ), .Z(\DP_OP_25_64_5665/n88 ) );
  NAND \DP_OP_25_64_5665/U221  ( .A(\DP_OP_25_64_5665/n280 ), .B(
        \DP_OP_25_64_5665/n248 ), .Z(\DP_OP_25_64_5665/n89 ) );
  NAND \DP_OP_25_64_5665/U321  ( .A(\DP_OP_25_64_5665/n88 ), .B(
        \DP_OP_25_64_5665/n89 ), .Z(\DP_OP_25_64_5665/n279 ) );
  NAND \DP_OP_25_64_5665/U120  ( .A(\DP_OP_25_64_5665/n316 ), .B(
        \U1/RSOP_16/C2/Z_20 ), .Z(\DP_OP_25_64_5665/n95 ) );
  NAND \DP_OP_25_64_5665/U220  ( .A(\DP_OP_25_64_5665/n281 ), .B(
        \DP_OP_25_64_5665/n249 ), .Z(\DP_OP_25_64_5665/n96 ) );
  NAND \DP_OP_25_64_5665/U320  ( .A(\DP_OP_25_64_5665/n95 ), .B(
        \DP_OP_25_64_5665/n96 ), .Z(\DP_OP_25_64_5665/n280 ) );
  NAND \DP_OP_25_64_5665/U119  ( .A(\DP_OP_25_64_5665/n317 ), .B(
        \U1/RSOP_16/C2/Z_19 ), .Z(\DP_OP_25_64_5665/n102 ) );
  NAND \DP_OP_25_64_5665/U219  ( .A(\DP_OP_25_64_5665/n282 ), .B(
        \DP_OP_25_64_5665/n250 ), .Z(\DP_OP_25_64_5665/n103 ) );
  NAND \DP_OP_25_64_5665/U319  ( .A(\DP_OP_25_64_5665/n102 ), .B(
        \DP_OP_25_64_5665/n103 ), .Z(\DP_OP_25_64_5665/n281 ) );
  NAND \DP_OP_25_64_5665/U118  ( .A(\DP_OP_25_64_5665/n318 ), .B(
        \U1/RSOP_16/C2/Z_18 ), .Z(\DP_OP_25_64_5665/n109 ) );
  NAND \DP_OP_25_64_5665/U218  ( .A(\DP_OP_25_64_5665/n283 ), .B(
        \DP_OP_25_64_5665/n251 ), .Z(\DP_OP_25_64_5665/n110 ) );
  NAND \DP_OP_25_64_5665/U318  ( .A(\DP_OP_25_64_5665/n109 ), .B(
        \DP_OP_25_64_5665/n110 ), .Z(\DP_OP_25_64_5665/n282 ) );
  NAND \DP_OP_25_64_5665/U117  ( .A(\DP_OP_25_64_5665/n319 ), .B(
        \U1/RSOP_16/C2/Z_17 ), .Z(\DP_OP_25_64_5665/n116 ) );
  NAND \DP_OP_25_64_5665/U217  ( .A(\DP_OP_25_64_5665/n284 ), .B(
        \DP_OP_25_64_5665/n252 ), .Z(\DP_OP_25_64_5665/n117 ) );
  NAND \DP_OP_25_64_5665/U317  ( .A(\DP_OP_25_64_5665/n116 ), .B(
        \DP_OP_25_64_5665/n117 ), .Z(\DP_OP_25_64_5665/n283 ) );
  NAND \DP_OP_25_64_5665/U116  ( .A(\DP_OP_25_64_5665/n320 ), .B(
        \U1/RSOP_16/C2/Z_16 ), .Z(\DP_OP_25_64_5665/n123 ) );
  NAND \DP_OP_25_64_5665/U216  ( .A(\DP_OP_25_64_5665/n285 ), .B(
        \DP_OP_25_64_5665/n253 ), .Z(\DP_OP_25_64_5665/n124 ) );
  NAND \DP_OP_25_64_5665/U316  ( .A(\DP_OP_25_64_5665/n123 ), .B(
        \DP_OP_25_64_5665/n124 ), .Z(\DP_OP_25_64_5665/n284 ) );
  NAND \DP_OP_25_64_5665/U115  ( .A(\DP_OP_25_64_5665/n321 ), .B(
        \U1/RSOP_16/C2/Z_15 ), .Z(\DP_OP_25_64_5665/n130 ) );
  NAND \DP_OP_25_64_5665/U215  ( .A(\DP_OP_25_64_5665/n286 ), .B(
        \DP_OP_25_64_5665/n254 ), .Z(\DP_OP_25_64_5665/n131 ) );
  NAND \DP_OP_25_64_5665/U315  ( .A(\DP_OP_25_64_5665/n130 ), .B(
        \DP_OP_25_64_5665/n131 ), .Z(\DP_OP_25_64_5665/n285 ) );
  NAND \DP_OP_25_64_5665/U114  ( .A(\DP_OP_25_64_5665/n322 ), .B(
        \U1/RSOP_16/C2/Z_14 ), .Z(\DP_OP_25_64_5665/n137 ) );
  NAND \DP_OP_25_64_5665/U214  ( .A(\DP_OP_25_64_5665/n287 ), .B(
        \DP_OP_25_64_5665/n255 ), .Z(\DP_OP_25_64_5665/n138 ) );
  NAND \DP_OP_25_64_5665/U314  ( .A(\DP_OP_25_64_5665/n137 ), .B(
        \DP_OP_25_64_5665/n138 ), .Z(\DP_OP_25_64_5665/n286 ) );
  NAND \DP_OP_25_64_5665/U113  ( .A(\DP_OP_25_64_5665/n323 ), .B(
        \U1/RSOP_16/C2/Z_13 ), .Z(\DP_OP_25_64_5665/n144 ) );
  NAND \DP_OP_25_64_5665/U213  ( .A(\DP_OP_25_64_5665/n288 ), .B(
        \DP_OP_25_64_5665/n256 ), .Z(\DP_OP_25_64_5665/n145 ) );
  NAND \DP_OP_25_64_5665/U313  ( .A(\DP_OP_25_64_5665/n144 ), .B(
        \DP_OP_25_64_5665/n145 ), .Z(\DP_OP_25_64_5665/n287 ) );
  NAND \DP_OP_25_64_5665/U112  ( .A(\DP_OP_25_64_5665/n324 ), .B(
        \U1/RSOP_16/C2/Z_12 ), .Z(\DP_OP_25_64_5665/n151 ) );
  NAND \DP_OP_25_64_5665/U212  ( .A(\DP_OP_25_64_5665/n289 ), .B(
        \DP_OP_25_64_5665/n257 ), .Z(\DP_OP_25_64_5665/n152 ) );
  NAND \DP_OP_25_64_5665/U312  ( .A(\DP_OP_25_64_5665/n151 ), .B(
        \DP_OP_25_64_5665/n152 ), .Z(\DP_OP_25_64_5665/n288 ) );
  NAND \DP_OP_25_64_5665/U111  ( .A(\DP_OP_25_64_5665/n325 ), .B(
        \U1/RSOP_16/C2/Z_11 ), .Z(\DP_OP_25_64_5665/n158 ) );
  NAND \DP_OP_25_64_5665/U211  ( .A(\DP_OP_25_64_5665/n290 ), .B(
        \DP_OP_25_64_5665/n258 ), .Z(\DP_OP_25_64_5665/n159 ) );
  NAND \DP_OP_25_64_5665/U311  ( .A(\DP_OP_25_64_5665/n158 ), .B(
        \DP_OP_25_64_5665/n159 ), .Z(\DP_OP_25_64_5665/n289 ) );
  NAND \DP_OP_25_64_5665/U110  ( .A(\DP_OP_25_64_5665/n326 ), .B(
        \U1/RSOP_16/C2/Z_10 ), .Z(\DP_OP_25_64_5665/n165 ) );
  NAND \DP_OP_25_64_5665/U210  ( .A(\DP_OP_25_64_5665/n291 ), .B(
        \DP_OP_25_64_5665/n259 ), .Z(\DP_OP_25_64_5665/n166 ) );
  NAND \DP_OP_25_64_5665/U310  ( .A(\DP_OP_25_64_5665/n165 ), .B(
        \DP_OP_25_64_5665/n166 ), .Z(\DP_OP_25_64_5665/n290 ) );
  NAND \DP_OP_25_64_5665/U19  ( .A(\DP_OP_25_64_5665/n327 ), .B(
        \U1/RSOP_16/C2/Z_9 ), .Z(\DP_OP_25_64_5665/n172 ) );
  NAND \DP_OP_25_64_5665/U29  ( .A(\DP_OP_25_64_5665/n292 ), .B(
        \DP_OP_25_64_5665/n260 ), .Z(\DP_OP_25_64_5665/n173 ) );
  NAND \DP_OP_25_64_5665/U39  ( .A(\DP_OP_25_64_5665/n172 ), .B(
        \DP_OP_25_64_5665/n173 ), .Z(\DP_OP_25_64_5665/n291 ) );
  NAND \DP_OP_25_64_5665/U18  ( .A(\DP_OP_25_64_5665/n328 ), .B(
        \U1/RSOP_16/C2/Z_8 ), .Z(\DP_OP_25_64_5665/n179 ) );
  NAND \DP_OP_25_64_5665/U28  ( .A(\DP_OP_25_64_5665/n293 ), .B(
        \DP_OP_25_64_5665/n261 ), .Z(\DP_OP_25_64_5665/n180 ) );
  NAND \DP_OP_25_64_5665/U38  ( .A(\DP_OP_25_64_5665/n179 ), .B(
        \DP_OP_25_64_5665/n180 ), .Z(\DP_OP_25_64_5665/n292 ) );
  NAND \DP_OP_25_64_5665/U17  ( .A(\DP_OP_25_64_5665/n329 ), .B(
        \U1/RSOP_16/C2/Z_7 ), .Z(\DP_OP_25_64_5665/n186 ) );
  NAND \DP_OP_25_64_5665/U27  ( .A(\DP_OP_25_64_5665/n294 ), .B(
        \DP_OP_25_64_5665/n262 ), .Z(\DP_OP_25_64_5665/n187 ) );
  NAND \DP_OP_25_64_5665/U37  ( .A(\DP_OP_25_64_5665/n186 ), .B(
        \DP_OP_25_64_5665/n187 ), .Z(\DP_OP_25_64_5665/n293 ) );
  NAND \DP_OP_25_64_5665/U16  ( .A(\DP_OP_25_64_5665/n330 ), .B(
        \U1/RSOP_16/C2/Z_6 ), .Z(\DP_OP_25_64_5665/n193 ) );
  NAND \DP_OP_25_64_5665/U26  ( .A(\DP_OP_25_64_5665/n295 ), .B(
        \DP_OP_25_64_5665/n263 ), .Z(\DP_OP_25_64_5665/n194 ) );
  NAND \DP_OP_25_64_5665/U36  ( .A(\DP_OP_25_64_5665/n193 ), .B(
        \DP_OP_25_64_5665/n194 ), .Z(\DP_OP_25_64_5665/n294 ) );
  NAND \DP_OP_25_64_5665/U15  ( .A(\DP_OP_25_64_5665/n331 ), .B(
        \U1/RSOP_16/C2/Z_5 ), .Z(\DP_OP_25_64_5665/n200 ) );
  NAND \DP_OP_25_64_5665/U25  ( .A(\DP_OP_25_64_5665/n296 ), .B(
        \DP_OP_25_64_5665/n264 ), .Z(\DP_OP_25_64_5665/n201 ) );
  NAND \DP_OP_25_64_5665/U35  ( .A(\DP_OP_25_64_5665/n200 ), .B(
        \DP_OP_25_64_5665/n201 ), .Z(\DP_OP_25_64_5665/n295 ) );
  NAND \DP_OP_25_64_5665/U14  ( .A(\DP_OP_25_64_5665/n332 ), .B(
        \U1/RSOP_16/C2/Z_4 ), .Z(\DP_OP_25_64_5665/n207 ) );
  NAND \DP_OP_25_64_5665/U24  ( .A(\DP_OP_25_64_5665/n297 ), .B(
        \DP_OP_25_64_5665/n265 ), .Z(\DP_OP_25_64_5665/n208 ) );
  NAND \DP_OP_25_64_5665/U34  ( .A(\DP_OP_25_64_5665/n207 ), .B(
        \DP_OP_25_64_5665/n208 ), .Z(\DP_OP_25_64_5665/n296 ) );
  NAND \DP_OP_25_64_5665/U13  ( .A(\DP_OP_25_64_5665/n333 ), .B(
        \U1/RSOP_16/C2/Z_3 ), .Z(\DP_OP_25_64_5665/n214 ) );
  NAND \DP_OP_25_64_5665/U23  ( .A(\DP_OP_25_64_5665/n298 ), .B(
        \DP_OP_25_64_5665/n266 ), .Z(\DP_OP_25_64_5665/n215 ) );
  NAND \DP_OP_25_64_5665/U33  ( .A(\DP_OP_25_64_5665/n214 ), .B(
        \DP_OP_25_64_5665/n215 ), .Z(\DP_OP_25_64_5665/n297 ) );
  NAND \DP_OP_25_64_5665/U12  ( .A(\DP_OP_25_64_5665/n334 ), .B(
        \U1/RSOP_16/C2/Z_2 ), .Z(\DP_OP_25_64_5665/n221 ) );
  NAND \DP_OP_25_64_5665/U22  ( .A(\DP_OP_25_64_5665/n299 ), .B(
        \DP_OP_25_64_5665/n267 ), .Z(\DP_OP_25_64_5665/n222 ) );
  NAND \DP_OP_25_64_5665/U32  ( .A(\DP_OP_25_64_5665/n221 ), .B(
        \DP_OP_25_64_5665/n222 ), .Z(\DP_OP_25_64_5665/n298 ) );
  NAND \DP_OP_25_64_5665/U11  ( .A(\DP_OP_25_64_5665/n335 ), .B(
        \U1/RSOP_16/C2/Z_1 ), .Z(\DP_OP_25_64_5665/n228 ) );
  NAND \DP_OP_25_64_5665/U21  ( .A(\DP_OP_25_64_5665/n300 ), .B(
        \DP_OP_25_64_5665/n268 ), .Z(\DP_OP_25_64_5665/n229 ) );
  NAND \DP_OP_25_64_5665/U31  ( .A(\DP_OP_25_64_5665/n228 ), .B(
        \DP_OP_25_64_5665/n229 ), .Z(\DP_OP_25_64_5665/n299 ) );
  NAND \DP_OP_25_64_5665/U1  ( .A(\U1/RSOP_16/C2/Z_0 ), .B(\C1/Z_0 ), .Z(
        \DP_OP_25_64_5665/n235 ) );
  NAND \DP_OP_25_64_5665/U2  ( .A(\DP_OP_25_64_5665/n269 ), .B(
        \DP_OP_25_64_5665/n336 ), .Z(\DP_OP_25_64_5665/n236 ) );
  NAND \DP_OP_25_64_5665/U3  ( .A(\DP_OP_25_64_5665/n235 ), .B(
        \DP_OP_25_64_5665/n236 ), .Z(\DP_OP_25_64_5665/n300 ) );
  XOR U1496 ( .A(n2863), .B(n2864), .Z(n2857) );
  NAND U1497 ( .A(n3108), .B(o[0]), .Z(n1495) );
  XNOR U1498 ( .A(o[2]), .B(n1495), .Z(n1496) );
  AND U1499 ( .A(\stack[1][20] ), .B(n1496), .Z(n3106) );
  NAND U1500 ( .A(n3366), .B(o[0]), .Z(n1497) );
  XNOR U1501 ( .A(o[2]), .B(n1497), .Z(n1498) );
  AND U1502 ( .A(\stack[1][22] ), .B(n1498), .Z(n3364) );
  NAND U1503 ( .A(n2990), .B(o[0]), .Z(n1499) );
  XNOR U1504 ( .A(o[2]), .B(n1499), .Z(n1500) );
  AND U1505 ( .A(\stack[1][19] ), .B(n1500), .Z(n2988) );
  XOR U1506 ( .A(n3090), .B(n3091), .Z(n3084) );
  NAND U1507 ( .A(n3229), .B(o[0]), .Z(n1501) );
  XNOR U1508 ( .A(o[2]), .B(n1501), .Z(n1502) );
  AND U1509 ( .A(\stack[1][21] ), .B(n1502), .Z(n3227) );
  NAND U1510 ( .A(n3505), .B(o[0]), .Z(n1503) );
  XNOR U1511 ( .A(o[2]), .B(n1503), .Z(n1504) );
  AND U1512 ( .A(\stack[1][23] ), .B(n1504), .Z(n3503) );
  NAND U1513 ( .A(n3806), .B(o[0]), .Z(n1505) );
  XNOR U1514 ( .A(o[2]), .B(n1505), .Z(n1506) );
  AND U1515 ( .A(\stack[1][25] ), .B(n1506), .Z(n3804) );
  NAND U1516 ( .A(n4126), .B(o[0]), .Z(n1507) );
  XNOR U1517 ( .A(o[2]), .B(n1507), .Z(n1508) );
  AND U1518 ( .A(\stack[1][27] ), .B(n1508), .Z(n4124) );
  NAND U1519 ( .A(n2768), .B(o[0]), .Z(n1509) );
  XNOR U1520 ( .A(o[2]), .B(n1509), .Z(n1510) );
  AND U1521 ( .A(\stack[1][17] ), .B(n1510), .Z(n2766) );
  NAND U1522 ( .A(o[0]), .B(n2990), .Z(n1511) );
  NANDN U1523 ( .A(o[2]), .B(n1511), .Z(n1512) );
  AND U1524 ( .A(\stack[1][19] ), .B(n1512), .Z(n1513) );
  NANDN U1525 ( .A(n2989), .B(n2988), .Z(n1514) );
  AND U1526 ( .A(n1513), .B(n1514), .Z(n3100) );
  XOR U1527 ( .A(n2297), .B(n2298), .Z(n2291) );
  NAND U1528 ( .A(o[0]), .B(n3229), .Z(n1515) );
  NANDN U1529 ( .A(o[2]), .B(n1515), .Z(n1516) );
  AND U1530 ( .A(\stack[1][21] ), .B(n1516), .Z(n1517) );
  NANDN U1531 ( .A(n3228), .B(n3227), .Z(n1518) );
  AND U1532 ( .A(n1517), .B(n1518), .Z(n3358) );
  NAND U1533 ( .A(o[0]), .B(n3505), .Z(n1519) );
  NANDN U1534 ( .A(o[2]), .B(n1519), .Z(n1520) );
  AND U1535 ( .A(\stack[1][23] ), .B(n1520), .Z(n1521) );
  NANDN U1536 ( .A(n3504), .B(n3503), .Z(n1522) );
  AND U1537 ( .A(n1521), .B(n1522), .Z(n3646) );
  NAND U1538 ( .A(o[0]), .B(n3806), .Z(n1523) );
  NANDN U1539 ( .A(o[2]), .B(n1523), .Z(n1524) );
  AND U1540 ( .A(\stack[1][25] ), .B(n1524), .Z(n1525) );
  NANDN U1541 ( .A(n3805), .B(n3804), .Z(n1526) );
  AND U1542 ( .A(n1525), .B(n1526), .Z(n3960) );
  NAND U1543 ( .A(o[0]), .B(n4126), .Z(n1527) );
  NANDN U1544 ( .A(o[2]), .B(n1527), .Z(n1528) );
  AND U1545 ( .A(\stack[1][27] ), .B(n1528), .Z(n1529) );
  NANDN U1546 ( .A(n4125), .B(n4124), .Z(n1530) );
  AND U1547 ( .A(n1529), .B(n1530), .Z(n4285) );
  NAND U1548 ( .A(n2665), .B(o[0]), .Z(n1531) );
  XNOR U1549 ( .A(o[2]), .B(n1531), .Z(n1532) );
  AND U1550 ( .A(\stack[1][16] ), .B(n1532), .Z(n2663) );
  NAND U1551 ( .A(n2881), .B(o[0]), .Z(n1533) );
  XNOR U1552 ( .A(o[2]), .B(n1533), .Z(n1534) );
  AND U1553 ( .A(\stack[1][18] ), .B(n1534), .Z(n2879) );
  NAND U1554 ( .A(o[0]), .B(n3366), .Z(n1535) );
  NANDN U1555 ( .A(o[2]), .B(n1535), .Z(n1536) );
  AND U1556 ( .A(\stack[1][22] ), .B(n1536), .Z(n1537) );
  NANDN U1557 ( .A(n3365), .B(n3364), .Z(n1538) );
  AND U1558 ( .A(n1537), .B(n1538), .Z(n3497) );
  NAND U1559 ( .A(n3654), .B(o[0]), .Z(n1539) );
  XNOR U1560 ( .A(o[2]), .B(n1539), .Z(n1540) );
  AND U1561 ( .A(\stack[1][24] ), .B(n1540), .Z(n3652) );
  XOR U1562 ( .A(n3636), .B(n3637), .Z(n3630) );
  NAND U1563 ( .A(n3968), .B(o[0]), .Z(n1541) );
  XNOR U1564 ( .A(o[2]), .B(n1541), .Z(n1542) );
  AND U1565 ( .A(\stack[1][26] ), .B(n1542), .Z(n3966) );
  XNOR U1566 ( .A(n2350), .B(n2351), .Z(n2410) );
  NAND U1567 ( .A(n4266), .B(o[0]), .Z(n1543) );
  XNOR U1568 ( .A(o[2]), .B(n1543), .Z(n1544) );
  AND U1569 ( .A(\stack[1][28] ), .B(n1544), .Z(n4264) );
  XOR U1570 ( .A(n4160), .B(n4161), .Z(n4078) );
  XNOR U1571 ( .A(n4026), .B(n4027), .Z(n3871) );
  XNOR U1572 ( .A(n3708), .B(n3709), .Z(n3570) );
  XNOR U1573 ( .A(n3419), .B(n3420), .Z(n3294) );
  XNOR U1574 ( .A(n3155), .B(n3156), .Z(n3043) );
  XNOR U1575 ( .A(n2916), .B(n2917), .Z(n2815) );
  NAND U1576 ( .A(o[0]), .B(n2315), .Z(n1545) );
  NANDN U1577 ( .A(o[2]), .B(n1545), .Z(n1546) );
  AND U1578 ( .A(\stack[1][12] ), .B(n1546), .Z(n1547) );
  NANDN U1579 ( .A(n2314), .B(n2313), .Z(n1548) );
  AND U1580 ( .A(n1547), .B(n1548), .Z(n2378) );
  NAND U1581 ( .A(o[0]), .B(n2239), .Z(n1549) );
  NANDN U1582 ( .A(o[2]), .B(n1549), .Z(n1550) );
  AND U1583 ( .A(\stack[1][11] ), .B(n1550), .Z(n1551) );
  NANDN U1584 ( .A(n2238), .B(n2237), .Z(n1552) );
  AND U1585 ( .A(n1551), .B(n1552), .Z(n2307) );
  NAND U1586 ( .A(o[0]), .B(n2386), .Z(n1553) );
  NANDN U1587 ( .A(o[2]), .B(n1553), .Z(n1554) );
  AND U1588 ( .A(\stack[1][13] ), .B(n1554), .Z(n1555) );
  NANDN U1589 ( .A(n2385), .B(n2384), .Z(n1556) );
  AND U1590 ( .A(n1555), .B(n1556), .Z(n2470) );
  NAND U1591 ( .A(o[0]), .B(n2170), .Z(n1557) );
  NANDN U1592 ( .A(o[2]), .B(n1557), .Z(n1558) );
  AND U1593 ( .A(\stack[1][10] ), .B(n1558), .Z(n1559) );
  NANDN U1594 ( .A(n2169), .B(n2168), .Z(n1560) );
  AND U1595 ( .A(n1559), .B(n1560), .Z(n2231) );
  NAND U1596 ( .A(o[0]), .B(n2478), .Z(n1561) );
  NANDN U1597 ( .A(o[2]), .B(n1561), .Z(n1562) );
  AND U1598 ( .A(\stack[1][14] ), .B(n1562), .Z(n1563) );
  NANDN U1599 ( .A(n2477), .B(n2476), .Z(n1564) );
  AND U1600 ( .A(n1563), .B(n1564), .Z(n2557) );
  NAND U1601 ( .A(o[0]), .B(n2565), .Z(n1565) );
  NANDN U1602 ( .A(o[2]), .B(n1565), .Z(n1566) );
  AND U1603 ( .A(\stack[1][15] ), .B(n1566), .Z(n1567) );
  NANDN U1604 ( .A(n2564), .B(n2563), .Z(n1568) );
  AND U1605 ( .A(n1567), .B(n1568), .Z(n2657) );
  NAND U1606 ( .A(o[0]), .B(n2104), .Z(n1569) );
  NANDN U1607 ( .A(o[2]), .B(n1569), .Z(n1570) );
  AND U1608 ( .A(\stack[1][9] ), .B(n1570), .Z(n1571) );
  NANDN U1609 ( .A(n2103), .B(n2102), .Z(n1572) );
  AND U1610 ( .A(n1571), .B(n1572), .Z(n2162) );
  NAND U1611 ( .A(o[0]), .B(n2665), .Z(n1573) );
  NANDN U1612 ( .A(o[2]), .B(n1573), .Z(n1574) );
  AND U1613 ( .A(\stack[1][16] ), .B(n1574), .Z(n1575) );
  NANDN U1614 ( .A(n2664), .B(n2663), .Z(n1576) );
  AND U1615 ( .A(n1575), .B(n1576), .Z(n2760) );
  NAND U1616 ( .A(o[0]), .B(n2053), .Z(n1577) );
  NANDN U1617 ( .A(o[2]), .B(n1577), .Z(n1578) );
  AND U1618 ( .A(\stack[1][8] ), .B(n1578), .Z(n1579) );
  NANDN U1619 ( .A(n2052), .B(n2051), .Z(n1580) );
  AND U1620 ( .A(n1579), .B(n1580), .Z(n2096) );
  NAND U1621 ( .A(o[0]), .B(n2768), .Z(n1581) );
  NANDN U1622 ( .A(o[2]), .B(n1581), .Z(n1582) );
  AND U1623 ( .A(\stack[1][17] ), .B(n1582), .Z(n1583) );
  NANDN U1624 ( .A(n2767), .B(n2766), .Z(n1584) );
  AND U1625 ( .A(n1583), .B(n1584), .Z(n2873) );
  NAND U1626 ( .A(o[0]), .B(n2881), .Z(n1585) );
  NANDN U1627 ( .A(o[2]), .B(n1585), .Z(n1586) );
  AND U1628 ( .A(\stack[1][18] ), .B(n1586), .Z(n1587) );
  NANDN U1629 ( .A(n2880), .B(n2879), .Z(n1588) );
  AND U1630 ( .A(n1587), .B(n1588), .Z(n2982) );
  XNOR U1631 ( .A(n2948), .B(n2949), .Z(n3005) );
  NAND U1632 ( .A(o[0]), .B(n3108), .Z(n1589) );
  NANDN U1633 ( .A(o[2]), .B(n1589), .Z(n1590) );
  AND U1634 ( .A(\stack[1][20] ), .B(n1590), .Z(n1591) );
  NANDN U1635 ( .A(n3107), .B(n3106), .Z(n1592) );
  AND U1636 ( .A(n1591), .B(n1592), .Z(n3221) );
  XOR U1637 ( .A(n3618), .B(n3619), .Z(n3671) );
  NAND U1638 ( .A(o[0]), .B(n3654), .Z(n1593) );
  NANDN U1639 ( .A(o[2]), .B(n1593), .Z(n1594) );
  AND U1640 ( .A(\stack[1][24] ), .B(n1594), .Z(n1595) );
  NANDN U1641 ( .A(n3653), .B(n3652), .Z(n1596) );
  AND U1642 ( .A(n1595), .B(n1596), .Z(n3798) );
  XNOR U1643 ( .A(n2442), .B(n2443), .Z(n2502) );
  XOR U1644 ( .A(n2147), .B(n2148), .Z(n2181) );
  XNOR U1645 ( .A(n1937), .B(n1938), .Z(n1953) );
  XNOR U1646 ( .A(n3764), .B(n3765), .Z(n3756) );
  XOR U1647 ( .A(n3950), .B(n3951), .Z(n3944) );
  XNOR U1648 ( .A(n3926), .B(n3927), .Z(n3919) );
  XOR U1649 ( .A(n2280), .B(n2281), .Z(n2334) );
  XNOR U1650 ( .A(n5570), .B(n1857), .Z(n1858) );
  NAND U1651 ( .A(o[0]), .B(n3968), .Z(n1597) );
  NANDN U1652 ( .A(o[2]), .B(n1597), .Z(n1598) );
  AND U1653 ( .A(\stack[1][26] ), .B(n1598), .Z(n1599) );
  NANDN U1654 ( .A(n3967), .B(n3966), .Z(n1600) );
  AND U1655 ( .A(n1599), .B(n1600), .Z(n4118) );
  XNOR U1656 ( .A(n4089), .B(n4090), .Z(n4151) );
  XOR U1657 ( .A(n4234), .B(n4235), .Z(n4419) );
  NAND U1658 ( .A(n4266), .B(o[0]), .Z(n1601) );
  NANDN U1659 ( .A(o[2]), .B(n1601), .Z(n1602) );
  NAND U1660 ( .A(n1602), .B(\stack[1][28] ), .Z(n4267) );
  XNOR U1661 ( .A(n4377), .B(n4378), .Z(n4248) );
  XNOR U1662 ( .A(n2203), .B(n2204), .Z(n2198) );
  XNOR U1663 ( .A(n2117), .B(n2118), .Z(n2075) );
  XNOR U1664 ( .A(n2700), .B(n2701), .Z(n2612) );
  XNOR U1665 ( .A(n2509), .B(n2510), .Z(n2430) );
  XNOR U1666 ( .A(n2344), .B(n2345), .Z(n2416) );
  XNOR U1667 ( .A(n2066), .B(n2067), .Z(n2023) );
  XOR U1668 ( .A(n1931), .B(n1932), .Z(n1925) );
  AND U1669 ( .A(\stack[1][0] ), .B(o[29]), .Z(n3867) );
  XNOR U1670 ( .A(n2268), .B(n2269), .Z(n2262) );
  XNOR U1671 ( .A(n1853), .B(n1854), .Z(n1845) );
  AND U1672 ( .A(\stack[1][0] ), .B(o[28]), .Z(n4609) );
  AND U1673 ( .A(\stack[1][0] ), .B(o[26]), .Z(n4685) );
  AND U1674 ( .A(\stack[1][0] ), .B(o[24]), .Z(n4761) );
  AND U1675 ( .A(\stack[1][0] ), .B(o[22]), .Z(n4837) );
  AND U1676 ( .A(\stack[1][0] ), .B(o[20]), .Z(n4913) );
  AND U1677 ( .A(\stack[1][0] ), .B(o[18]), .Z(n4989) );
  AND U1678 ( .A(\stack[1][0] ), .B(o[16]), .Z(n5065) );
  ANDN U1679 ( .B(opcode[2]), .A(opcode[0]), .Z(n1603) );
  AND U1680 ( .A(n1724), .B(n1603), .Z(n5672) );
  IV U1681 ( .A(n5663), .Z(n1604) );
  IV U1682 ( .A(n5672), .Z(n1605) );
  IV U1683 ( .A(\stack[1][0] ), .Z(n1606) );
  IV U1684 ( .A(\stack[1][2] ), .Z(n1607) );
  IV U1685 ( .A(\stack[1][3] ), .Z(n1608) );
  IV U1686 ( .A(\stack[1][4] ), .Z(n1609) );
  IV U1687 ( .A(\stack[1][5] ), .Z(n1610) );
  IV U1688 ( .A(\stack[1][6] ), .Z(n1611) );
  IV U1689 ( .A(\stack[1][7] ), .Z(n1612) );
  IV U1690 ( .A(\stack[1][8] ), .Z(n1613) );
  IV U1691 ( .A(\stack[1][9] ), .Z(n1614) );
  IV U1692 ( .A(\stack[1][10] ), .Z(n1615) );
  IV U1693 ( .A(\stack[1][11] ), .Z(n1616) );
  IV U1694 ( .A(\stack[1][12] ), .Z(n1617) );
  IV U1695 ( .A(\stack[1][14] ), .Z(n1618) );
  IV U1696 ( .A(o[1]), .Z(n1619) );
  IV U1697 ( .A(o[8]), .Z(n1620) );
  IV U1698 ( .A(o[10]), .Z(n1621) );
  IV U1699 ( .A(opcode[1]), .Z(n1724) );
  ANDN U1700 ( .B(opcode[0]), .A(opcode[1]), .Z(n1689) );
  ANDN U1701 ( .B(n1689), .A(opcode[2]), .Z(n1723) );
  NANDN U1702 ( .A(opcode[0]), .B(opcode[1]), .Z(n4499) );
  OR U1703 ( .A(opcode[2]), .B(n4499), .Z(n1688) );
  NANDN U1704 ( .A(n1723), .B(n1688), .Z(n1684) );
  AND U1705 ( .A(o[31]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_31 ) );
  AND U1706 ( .A(o[30]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_30 ) );
  AND U1707 ( .A(o[29]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_29 ) );
  AND U1708 ( .A(o[28]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_28 ) );
  AND U1709 ( .A(o[27]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_27 ) );
  AND U1710 ( .A(o[26]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_26 ) );
  AND U1711 ( .A(o[25]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_25 ) );
  AND U1712 ( .A(o[24]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_24 ) );
  AND U1713 ( .A(o[23]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_23 ) );
  AND U1714 ( .A(o[22]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_22 ) );
  AND U1715 ( .A(o[21]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_21 ) );
  AND U1716 ( .A(o[20]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_20 ) );
  AND U1717 ( .A(o[19]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_19 ) );
  AND U1718 ( .A(o[18]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_18 ) );
  AND U1719 ( .A(o[17]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_17 ) );
  AND U1720 ( .A(o[16]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_16 ) );
  AND U1721 ( .A(o[15]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_15 ) );
  AND U1722 ( .A(o[14]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_14 ) );
  AND U1723 ( .A(o[13]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_13 ) );
  AND U1724 ( .A(o[12]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_12 ) );
  AND U1725 ( .A(o[11]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_11 ) );
  AND U1726 ( .A(o[10]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_10 ) );
  AND U1727 ( .A(o[9]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_9 ) );
  AND U1728 ( .A(o[8]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_8 ) );
  AND U1729 ( .A(o[7]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_7 ) );
  AND U1730 ( .A(o[6]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_6 ) );
  AND U1731 ( .A(o[5]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_5 ) );
  AND U1732 ( .A(o[4]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_4 ) );
  AND U1733 ( .A(o[3]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_3 ) );
  AND U1734 ( .A(o[2]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_2 ) );
  AND U1735 ( .A(o[1]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_1 ) );
  AND U1736 ( .A(o[0]), .B(n1684), .Z(\U1/RSOP_16/C2/Z_0 ) );
  AND U1737 ( .A(n1689), .B(opcode[2]), .Z(n1687) );
  NAND U1738 ( .A(n1687), .B(o[31]), .Z(n1623) );
  NAND U1739 ( .A(\stack[1][31] ), .B(n1684), .Z(n1622) );
  NAND U1740 ( .A(n1623), .B(n1622), .Z(\U1/RSOP_16/C3/Z_31 ) );
  NAND U1741 ( .A(n1687), .B(o[30]), .Z(n1625) );
  NAND U1742 ( .A(\stack[1][30] ), .B(n1684), .Z(n1624) );
  NAND U1743 ( .A(n1625), .B(n1624), .Z(\U1/RSOP_16/C3/Z_30 ) );
  NAND U1744 ( .A(n1687), .B(o[29]), .Z(n1627) );
  NAND U1745 ( .A(\stack[1][29] ), .B(n1684), .Z(n1626) );
  NAND U1746 ( .A(n1627), .B(n1626), .Z(\U1/RSOP_16/C3/Z_29 ) );
  NAND U1747 ( .A(n1687), .B(o[28]), .Z(n1629) );
  NAND U1748 ( .A(\stack[1][28] ), .B(n1684), .Z(n1628) );
  NAND U1749 ( .A(n1629), .B(n1628), .Z(\U1/RSOP_16/C3/Z_28 ) );
  NAND U1750 ( .A(n1687), .B(o[27]), .Z(n1631) );
  NAND U1751 ( .A(\stack[1][27] ), .B(n1684), .Z(n1630) );
  NAND U1752 ( .A(n1631), .B(n1630), .Z(\U1/RSOP_16/C3/Z_27 ) );
  NAND U1753 ( .A(n1687), .B(o[26]), .Z(n1633) );
  NAND U1754 ( .A(\stack[1][26] ), .B(n1684), .Z(n1632) );
  NAND U1755 ( .A(n1633), .B(n1632), .Z(\U1/RSOP_16/C3/Z_26 ) );
  NAND U1756 ( .A(n1687), .B(o[25]), .Z(n1635) );
  NAND U1757 ( .A(\stack[1][25] ), .B(n1684), .Z(n1634) );
  NAND U1758 ( .A(n1635), .B(n1634), .Z(\U1/RSOP_16/C3/Z_25 ) );
  NAND U1759 ( .A(n1687), .B(o[24]), .Z(n1637) );
  NAND U1760 ( .A(\stack[1][24] ), .B(n1684), .Z(n1636) );
  NAND U1761 ( .A(n1637), .B(n1636), .Z(\U1/RSOP_16/C3/Z_24 ) );
  NAND U1762 ( .A(n1687), .B(o[23]), .Z(n1639) );
  NAND U1763 ( .A(\stack[1][23] ), .B(n1684), .Z(n1638) );
  NAND U1764 ( .A(n1639), .B(n1638), .Z(\U1/RSOP_16/C3/Z_23 ) );
  NAND U1765 ( .A(n1687), .B(o[22]), .Z(n1641) );
  NAND U1766 ( .A(\stack[1][22] ), .B(n1684), .Z(n1640) );
  NAND U1767 ( .A(n1641), .B(n1640), .Z(\U1/RSOP_16/C3/Z_22 ) );
  NAND U1768 ( .A(n1687), .B(o[21]), .Z(n1643) );
  NAND U1769 ( .A(\stack[1][21] ), .B(n1684), .Z(n1642) );
  NAND U1770 ( .A(n1643), .B(n1642), .Z(\U1/RSOP_16/C3/Z_21 ) );
  NAND U1771 ( .A(n1687), .B(o[20]), .Z(n1645) );
  NAND U1772 ( .A(\stack[1][20] ), .B(n1684), .Z(n1644) );
  NAND U1773 ( .A(n1645), .B(n1644), .Z(\U1/RSOP_16/C3/Z_20 ) );
  NAND U1774 ( .A(n1687), .B(o[19]), .Z(n1647) );
  NAND U1775 ( .A(\stack[1][19] ), .B(n1684), .Z(n1646) );
  NAND U1776 ( .A(n1647), .B(n1646), .Z(\U1/RSOP_16/C3/Z_19 ) );
  NAND U1777 ( .A(n1687), .B(o[18]), .Z(n1649) );
  NAND U1778 ( .A(\stack[1][18] ), .B(n1684), .Z(n1648) );
  NAND U1779 ( .A(n1649), .B(n1648), .Z(\U1/RSOP_16/C3/Z_18 ) );
  NAND U1780 ( .A(n1687), .B(o[17]), .Z(n1651) );
  NAND U1781 ( .A(\stack[1][17] ), .B(n1684), .Z(n1650) );
  NAND U1782 ( .A(n1651), .B(n1650), .Z(\U1/RSOP_16/C3/Z_17 ) );
  NAND U1783 ( .A(n1687), .B(o[16]), .Z(n1653) );
  NAND U1784 ( .A(\stack[1][16] ), .B(n1684), .Z(n1652) );
  NAND U1785 ( .A(n1653), .B(n1652), .Z(\U1/RSOP_16/C3/Z_16 ) );
  NAND U1786 ( .A(n1687), .B(o[15]), .Z(n1655) );
  NAND U1787 ( .A(\stack[1][15] ), .B(n1684), .Z(n1654) );
  NAND U1788 ( .A(n1655), .B(n1654), .Z(\U1/RSOP_16/C3/Z_15 ) );
  NAND U1789 ( .A(n1687), .B(o[14]), .Z(n1657) );
  NAND U1790 ( .A(\stack[1][14] ), .B(n1684), .Z(n1656) );
  NAND U1791 ( .A(n1657), .B(n1656), .Z(\U1/RSOP_16/C3/Z_14 ) );
  NAND U1792 ( .A(n1687), .B(o[13]), .Z(n1659) );
  NAND U1793 ( .A(\stack[1][13] ), .B(n1684), .Z(n1658) );
  NAND U1794 ( .A(n1659), .B(n1658), .Z(\U1/RSOP_16/C3/Z_13 ) );
  NAND U1795 ( .A(n1687), .B(o[12]), .Z(n1661) );
  NAND U1796 ( .A(\stack[1][12] ), .B(n1684), .Z(n1660) );
  NAND U1797 ( .A(n1661), .B(n1660), .Z(\U1/RSOP_16/C3/Z_12 ) );
  NAND U1798 ( .A(n1687), .B(o[11]), .Z(n1663) );
  NAND U1799 ( .A(\stack[1][11] ), .B(n1684), .Z(n1662) );
  NAND U1800 ( .A(n1663), .B(n1662), .Z(\U1/RSOP_16/C3/Z_11 ) );
  NAND U1801 ( .A(n1687), .B(o[10]), .Z(n1665) );
  NAND U1802 ( .A(\stack[1][10] ), .B(n1684), .Z(n1664) );
  NAND U1803 ( .A(n1665), .B(n1664), .Z(\U1/RSOP_16/C3/Z_10 ) );
  NAND U1804 ( .A(n1687), .B(o[9]), .Z(n1667) );
  NAND U1805 ( .A(\stack[1][9] ), .B(n1684), .Z(n1666) );
  NAND U1806 ( .A(n1667), .B(n1666), .Z(\U1/RSOP_16/C3/Z_9 ) );
  NAND U1807 ( .A(n1687), .B(o[8]), .Z(n1669) );
  NAND U1808 ( .A(\stack[1][8] ), .B(n1684), .Z(n1668) );
  NAND U1809 ( .A(n1669), .B(n1668), .Z(\U1/RSOP_16/C3/Z_8 ) );
  NAND U1810 ( .A(n1687), .B(o[7]), .Z(n1671) );
  NAND U1811 ( .A(\stack[1][7] ), .B(n1684), .Z(n1670) );
  NAND U1812 ( .A(n1671), .B(n1670), .Z(\U1/RSOP_16/C3/Z_7 ) );
  NAND U1813 ( .A(n1687), .B(o[6]), .Z(n1673) );
  NAND U1814 ( .A(\stack[1][6] ), .B(n1684), .Z(n1672) );
  NAND U1815 ( .A(n1673), .B(n1672), .Z(\U1/RSOP_16/C3/Z_6 ) );
  NAND U1816 ( .A(n1687), .B(o[5]), .Z(n1675) );
  NAND U1817 ( .A(\stack[1][5] ), .B(n1684), .Z(n1674) );
  NAND U1818 ( .A(n1675), .B(n1674), .Z(\U1/RSOP_16/C3/Z_5 ) );
  NAND U1819 ( .A(n1687), .B(o[4]), .Z(n1677) );
  NAND U1820 ( .A(\stack[1][4] ), .B(n1684), .Z(n1676) );
  NAND U1821 ( .A(n1677), .B(n1676), .Z(\U1/RSOP_16/C3/Z_4 ) );
  NAND U1822 ( .A(n1687), .B(o[3]), .Z(n1679) );
  NAND U1823 ( .A(\stack[1][3] ), .B(n1684), .Z(n1678) );
  NAND U1824 ( .A(n1679), .B(n1678), .Z(\U1/RSOP_16/C3/Z_3 ) );
  NAND U1825 ( .A(n1687), .B(o[2]), .Z(n1681) );
  NAND U1826 ( .A(\stack[1][2] ), .B(n1684), .Z(n1680) );
  NAND U1827 ( .A(n1681), .B(n1680), .Z(\U1/RSOP_16/C3/Z_2 ) );
  NAND U1828 ( .A(n1687), .B(o[1]), .Z(n1683) );
  NAND U1829 ( .A(\stack[1][1] ), .B(n1684), .Z(n1682) );
  NAND U1830 ( .A(n1683), .B(n1682), .Z(\U1/RSOP_16/C3/Z_1 ) );
  NAND U1831 ( .A(n1687), .B(o[0]), .Z(n1686) );
  NAND U1832 ( .A(\stack[1][0] ), .B(n1684), .Z(n1685) );
  NAND U1833 ( .A(n1686), .B(n1685), .Z(\U1/RSOP_16/C3/Z_0 ) );
  NANDN U1834 ( .A(n1687), .B(n1688), .Z(\C1/Z_0 ) );
  NANDN U1835 ( .A(n1689), .B(n1688), .Z(n1721) );
  NAND U1836 ( .A(\C3/DATA5_31 ), .B(n1721), .Z(n1690) );
  NAND U1837 ( .A(n1773), .B(n1690), .Z(n4496) );
  NAND U1838 ( .A(\C3/DATA5_30 ), .B(n1721), .Z(n1691) );
  AND U1839 ( .A(n4535), .B(n1691), .Z(n4536) );
  NAND U1840 ( .A(\C3/DATA5_29 ), .B(n1721), .Z(n1692) );
  ANDN U1841 ( .B(n1692), .A(n4579), .Z(n4580) );
  NAND U1842 ( .A(\C3/DATA5_28 ), .B(n1721), .Z(n1693) );
  AND U1843 ( .A(n4611), .B(n1693), .Z(n4612) );
  NAND U1844 ( .A(\C3/DATA5_27 ), .B(n1721), .Z(n1694) );
  ANDN U1845 ( .B(n1694), .A(n4655), .Z(n4656) );
  NAND U1846 ( .A(\C3/DATA5_26 ), .B(n1721), .Z(n1695) );
  AND U1847 ( .A(n4687), .B(n1695), .Z(n4688) );
  NAND U1848 ( .A(\C3/DATA5_25 ), .B(n1721), .Z(n1696) );
  ANDN U1849 ( .B(n1696), .A(n4731), .Z(n4732) );
  NAND U1850 ( .A(\C3/DATA5_24 ), .B(n1721), .Z(n1697) );
  AND U1851 ( .A(n4763), .B(n1697), .Z(n4764) );
  NAND U1852 ( .A(\C3/DATA5_23 ), .B(n1721), .Z(n1698) );
  ANDN U1853 ( .B(n1698), .A(n4807), .Z(n4808) );
  NAND U1854 ( .A(\C3/DATA5_22 ), .B(n1721), .Z(n1699) );
  AND U1855 ( .A(n4839), .B(n1699), .Z(n4840) );
  NAND U1856 ( .A(\C3/DATA5_21 ), .B(n1721), .Z(n1700) );
  ANDN U1857 ( .B(n1700), .A(n4883), .Z(n4884) );
  NAND U1858 ( .A(\C3/DATA5_20 ), .B(n1721), .Z(n1701) );
  AND U1859 ( .A(n4915), .B(n1701), .Z(n4916) );
  NAND U1860 ( .A(\C3/DATA5_19 ), .B(n1721), .Z(n1702) );
  ANDN U1861 ( .B(n1702), .A(n4959), .Z(n4960) );
  NAND U1862 ( .A(\C3/DATA5_18 ), .B(n1721), .Z(n1703) );
  AND U1863 ( .A(n4991), .B(n1703), .Z(n4992) );
  NAND U1864 ( .A(\C3/DATA5_17 ), .B(n1721), .Z(n1704) );
  ANDN U1865 ( .B(n1704), .A(n5035), .Z(n5036) );
  NAND U1866 ( .A(\C3/DATA5_16 ), .B(n1721), .Z(n1705) );
  AND U1867 ( .A(n5067), .B(n1705), .Z(n5068) );
  NAND U1868 ( .A(\C3/DATA5_15 ), .B(n1721), .Z(n1706) );
  NAND U1869 ( .A(n5103), .B(n1706), .Z(n5108) );
  NAND U1870 ( .A(\C3/DATA5_14 ), .B(n1721), .Z(n1707) );
  AND U1871 ( .A(n5144), .B(n1707), .Z(n5145) );
  NAND U1872 ( .A(\C3/DATA5_13 ), .B(n1721), .Z(n1708) );
  AND U1873 ( .A(n5183), .B(n1708), .Z(n5184) );
  NAND U1874 ( .A(\C3/DATA5_12 ), .B(n1721), .Z(n1709) );
  AND U1875 ( .A(n5221), .B(n1709), .Z(n5222) );
  NAND U1876 ( .A(\C3/DATA5_11 ), .B(n1721), .Z(n1710) );
  AND U1877 ( .A(n5260), .B(n1710), .Z(n5261) );
  NAND U1878 ( .A(\C3/DATA5_10 ), .B(n1721), .Z(n1711) );
  AND U1879 ( .A(n5298), .B(n1711), .Z(n5299) );
  NAND U1880 ( .A(\C3/DATA5_9 ), .B(n1721), .Z(n1712) );
  AND U1881 ( .A(n5337), .B(n1712), .Z(n5338) );
  NAND U1882 ( .A(\C3/DATA5_8 ), .B(n1721), .Z(n1713) );
  AND U1883 ( .A(n5375), .B(n1713), .Z(n5376) );
  NAND U1884 ( .A(\C3/DATA5_7 ), .B(n1721), .Z(n1714) );
  AND U1885 ( .A(n5413), .B(n1714), .Z(n5414) );
  NAND U1886 ( .A(\C3/DATA5_6 ), .B(n1721), .Z(n1715) );
  AND U1887 ( .A(n5453), .B(n1715), .Z(n5454) );
  NAND U1888 ( .A(\C3/DATA5_5 ), .B(n1721), .Z(n1716) );
  AND U1889 ( .A(n5491), .B(n1716), .Z(n5492) );
  NAND U1890 ( .A(\C3/DATA5_4 ), .B(n1721), .Z(n1717) );
  AND U1891 ( .A(n5529), .B(n1717), .Z(n5530) );
  NAND U1892 ( .A(\C3/DATA5_3 ), .B(n1721), .Z(n1718) );
  NAND U1893 ( .A(n5564), .B(n1718), .Z(n5569) );
  NAND U1894 ( .A(\C3/DATA5_2 ), .B(n1721), .Z(n1719) );
  NAND U1895 ( .A(n5607), .B(n1719), .Z(n5611) );
  NAND U1896 ( .A(\C3/DATA5_1 ), .B(n1721), .Z(n1720) );
  AND U1897 ( .A(n5654), .B(n1720), .Z(n5655) );
  NAND U1898 ( .A(\C3/DATA5_0 ), .B(n1721), .Z(n1722) );
  AND U1899 ( .A(n5673), .B(n1722), .Z(n5674) );
  NAND U1900 ( .A(n5672), .B(\stack[6][0] ), .Z(n1726) );
  NAND U1901 ( .A(n1605), .B(\stack[7][0] ), .Z(n1725) );
  NAND U1902 ( .A(n1726), .B(n1725), .Z(n1065) );
  NAND U1903 ( .A(n5672), .B(\stack[5][0] ), .Z(n1728) );
  ANDN U1904 ( .B(n1724), .A(n1723), .Z(n5657) );
  NANDN U1905 ( .A(n5657), .B(\stack[7][0] ), .Z(n1727) );
  AND U1906 ( .A(n1728), .B(n1727), .Z(n1730) );
  XNOR U1907 ( .A(opcode[2]), .B(opcode[0]), .Z(n4498) );
  NAND U1908 ( .A(n1724), .B(n4498), .Z(n5660) );
  NANDN U1909 ( .A(n5660), .B(\stack[6][0] ), .Z(n1729) );
  NAND U1910 ( .A(n1730), .B(n1729), .Z(n1066) );
  NAND U1911 ( .A(n5672), .B(\stack[4][0] ), .Z(n1732) );
  NANDN U1912 ( .A(n5657), .B(\stack[6][0] ), .Z(n1731) );
  AND U1913 ( .A(n1732), .B(n1731), .Z(n1734) );
  NANDN U1914 ( .A(n5660), .B(\stack[5][0] ), .Z(n1733) );
  NAND U1915 ( .A(n1734), .B(n1733), .Z(n1067) );
  NAND U1916 ( .A(n5672), .B(\stack[3][0] ), .Z(n1736) );
  NANDN U1917 ( .A(n5657), .B(\stack[5][0] ), .Z(n1735) );
  AND U1918 ( .A(n1736), .B(n1735), .Z(n1738) );
  NANDN U1919 ( .A(n5660), .B(\stack[4][0] ), .Z(n1737) );
  NAND U1920 ( .A(n1738), .B(n1737), .Z(n1068) );
  NAND U1921 ( .A(n5672), .B(\stack[2][0] ), .Z(n1740) );
  NANDN U1922 ( .A(n5657), .B(\stack[4][0] ), .Z(n1739) );
  AND U1923 ( .A(n1740), .B(n1739), .Z(n1742) );
  NANDN U1924 ( .A(n5660), .B(\stack[3][0] ), .Z(n1741) );
  NAND U1925 ( .A(n1742), .B(n1741), .Z(n1069) );
  NAND U1926 ( .A(\stack[1][0] ), .B(n5672), .Z(n1744) );
  NANDN U1927 ( .A(n5657), .B(\stack[3][0] ), .Z(n1743) );
  AND U1928 ( .A(n1744), .B(n1743), .Z(n1746) );
  NANDN U1929 ( .A(n5660), .B(\stack[2][0] ), .Z(n1745) );
  NAND U1930 ( .A(n1746), .B(n1745), .Z(n1070) );
  NAND U1931 ( .A(n5672), .B(\stack[6][31] ), .Z(n1748) );
  NAND U1932 ( .A(n1605), .B(\stack[7][31] ), .Z(n1747) );
  NAND U1933 ( .A(n1748), .B(n1747), .Z(n1071) );
  NAND U1934 ( .A(n5672), .B(\stack[5][31] ), .Z(n1750) );
  NANDN U1935 ( .A(n5657), .B(\stack[7][31] ), .Z(n1749) );
  AND U1936 ( .A(n1750), .B(n1749), .Z(n1752) );
  NANDN U1937 ( .A(n5660), .B(\stack[6][31] ), .Z(n1751) );
  NAND U1938 ( .A(n1752), .B(n1751), .Z(n1072) );
  NAND U1939 ( .A(n5672), .B(\stack[4][31] ), .Z(n1754) );
  NANDN U1940 ( .A(n5657), .B(\stack[6][31] ), .Z(n1753) );
  AND U1941 ( .A(n1754), .B(n1753), .Z(n1756) );
  NANDN U1942 ( .A(n5660), .B(\stack[5][31] ), .Z(n1755) );
  NAND U1943 ( .A(n1756), .B(n1755), .Z(n1073) );
  NAND U1944 ( .A(n5672), .B(\stack[3][31] ), .Z(n1758) );
  NANDN U1945 ( .A(n5657), .B(\stack[5][31] ), .Z(n1757) );
  AND U1946 ( .A(n1758), .B(n1757), .Z(n1760) );
  NANDN U1947 ( .A(n5660), .B(\stack[4][31] ), .Z(n1759) );
  NAND U1948 ( .A(n1760), .B(n1759), .Z(n1074) );
  NAND U1949 ( .A(n5672), .B(\stack[2][31] ), .Z(n1762) );
  NANDN U1950 ( .A(n5657), .B(\stack[4][31] ), .Z(n1761) );
  AND U1951 ( .A(n1762), .B(n1761), .Z(n1764) );
  NANDN U1952 ( .A(n5660), .B(\stack[3][31] ), .Z(n1763) );
  NAND U1953 ( .A(n1764), .B(n1763), .Z(n1075) );
  NAND U1954 ( .A(n5672), .B(\stack[1][31] ), .Z(n1766) );
  NANDN U1955 ( .A(n5657), .B(\stack[3][31] ), .Z(n1765) );
  AND U1956 ( .A(n1766), .B(n1765), .Z(n1768) );
  NANDN U1957 ( .A(n5660), .B(\stack[2][31] ), .Z(n1767) );
  NAND U1958 ( .A(n1768), .B(n1767), .Z(n1076) );
  NAND U1959 ( .A(n5672), .B(o[31]), .Z(n1770) );
  NANDN U1960 ( .A(n5657), .B(\stack[2][31] ), .Z(n1769) );
  AND U1961 ( .A(n1770), .B(n1769), .Z(n1772) );
  NANDN U1962 ( .A(n5660), .B(\stack[1][31] ), .Z(n1771) );
  NAND U1963 ( .A(n1772), .B(n1771), .Z(n1077) );
  NAND U1964 ( .A(n5672), .B(x[31]), .Z(n1773) );
  IV U1965 ( .A(o[27]), .Z(n4023) );
  ANDN U1966 ( .B(\stack[1][0] ), .A(n4023), .Z(n3566) );
  IV U1967 ( .A(o[25]), .Z(n4016) );
  ANDN U1968 ( .B(\stack[1][0] ), .A(n4016), .Z(n3290) );
  IV U1969 ( .A(o[23]), .Z(n3699) );
  ANDN U1970 ( .B(\stack[1][0] ), .A(n3699), .Z(n3039) );
  IV U1971 ( .A(o[21]), .Z(n4170) );
  ANDN U1972 ( .B(\stack[1][0] ), .A(n4170), .Z(n2811) );
  IV U1973 ( .A(o[19]), .Z(n4068) );
  ANDN U1974 ( .B(\stack[1][0] ), .A(n4068), .Z(n2608) );
  IV U1975 ( .A(o[17]), .Z(n3911) );
  ANDN U1976 ( .B(\stack[1][0] ), .A(n3911), .Z(n2426) );
  ANDN U1977 ( .B(o[15]), .A(n1606), .Z(n2338) );
  IV U1978 ( .A(o[13]), .Z(n3923) );
  ANDN U1979 ( .B(\stack[1][0] ), .A(n3923), .Z(n2131) );
  IV U1980 ( .A(o[11]), .Z(n4144) );
  ANDN U1981 ( .B(\stack[1][0] ), .A(n4144), .Z(n2019) );
  IV U1982 ( .A(o[9]), .Z(n3977) );
  ANDN U1983 ( .B(\stack[1][0] ), .A(n3977), .Z(n1921) );
  IV U1984 ( .A(o[7]), .Z(n4111) );
  ANDN U1985 ( .B(\stack[1][0] ), .A(n4111), .Z(n1849) );
  IV U1986 ( .A(o[5]), .Z(n4130) );
  ANDN U1987 ( .B(\stack[1][0] ), .A(n4130), .Z(n1802) );
  IV U1988 ( .A(o[3]), .Z(n4127) );
  ANDN U1989 ( .B(\stack[1][0] ), .A(n4127), .Z(n1781) );
  IV U1990 ( .A(\stack[1][1] ), .Z(n4195) );
  ANDN U1991 ( .B(o[0]), .A(n4195), .Z(n5643) );
  NAND U1992 ( .A(o[1]), .B(n5643), .Z(n1774) );
  XNOR U1993 ( .A(o[2]), .B(n1774), .Z(n1775) );
  NAND U1994 ( .A(\stack[1][0] ), .B(n1775), .Z(n5603) );
  AND U1995 ( .A(o[0]), .B(\stack[1][2] ), .Z(n1810) );
  AND U1996 ( .A(\stack[1][1] ), .B(o[1]), .Z(n1776) );
  XOR U1997 ( .A(n1810), .B(n1776), .Z(n5604) );
  OR U1998 ( .A(n5603), .B(n5604), .Z(n1780) );
  NAND U1999 ( .A(o[1]), .B(\stack[1][0] ), .Z(n5642) );
  NANDN U2000 ( .A(n5642), .B(n5643), .Z(n1778) );
  NAND U2001 ( .A(\stack[1][0] ), .B(o[2]), .Z(n1777) );
  AND U2002 ( .A(n1778), .B(n1777), .Z(n1779) );
  ANDN U2003 ( .B(n1780), .A(n1779), .Z(n1782) );
  OR U2004 ( .A(n1781), .B(n1782), .Z(n1787) );
  XNOR U2005 ( .A(n1782), .B(n1781), .Z(n5565) );
  AND U2006 ( .A(\stack[1][2] ), .B(o[1]), .Z(n1783) );
  AND U2007 ( .A(o[0]), .B(\stack[1][3] ), .Z(n1831) );
  XOR U2008 ( .A(n1783), .B(n1831), .Z(n1788) );
  NAND U2009 ( .A(o[1]), .B(\stack[1][2] ), .Z(n1790) );
  NANDN U2010 ( .A(n1790), .B(o[0]), .Z(n1784) );
  XNOR U2011 ( .A(o[2]), .B(n1784), .Z(n1785) );
  NAND U2012 ( .A(\stack[1][1] ), .B(n1785), .Z(n1789) );
  XNOR U2013 ( .A(n1788), .B(n1789), .Z(n5566) );
  OR U2014 ( .A(n5565), .B(n5566), .Z(n1786) );
  AND U2015 ( .A(n1787), .B(n1786), .Z(n1799) );
  OR U2016 ( .A(n1789), .B(n1788), .Z(n1794) );
  NANDN U2017 ( .A(n1790), .B(n5643), .Z(n1792) );
  NAND U2018 ( .A(\stack[1][1] ), .B(o[2]), .Z(n1791) );
  AND U2019 ( .A(n1792), .B(n1791), .Z(n1793) );
  ANDN U2020 ( .B(n1794), .A(n1793), .Z(n1804) );
  ANDN U2021 ( .B(o[3]), .A(n4195), .Z(n1805) );
  XNOR U2022 ( .A(n1804), .B(n1805), .Z(n1807) );
  AND U2023 ( .A(\stack[1][3] ), .B(o[1]), .Z(n1795) );
  AND U2024 ( .A(o[0]), .B(\stack[1][4] ), .Z(n1864) );
  XOR U2025 ( .A(n1795), .B(n1864), .Z(n1813) );
  NAND U2026 ( .A(o[1]), .B(\stack[1][3] ), .Z(n1811) );
  NANDN U2027 ( .A(n1811), .B(o[0]), .Z(n1796) );
  XNOR U2028 ( .A(o[2]), .B(n1796), .Z(n1797) );
  NAND U2029 ( .A(\stack[1][2] ), .B(n1797), .Z(n1814) );
  XNOR U2030 ( .A(n1813), .B(n1814), .Z(n1806) );
  XOR U2031 ( .A(n1807), .B(n1806), .Z(n1798) );
  NANDN U2032 ( .A(n1799), .B(n1798), .Z(n1801) );
  XOR U2033 ( .A(n1799), .B(n1798), .Z(n5526) );
  IV U2034 ( .A(o[4]), .Z(n4129) );
  ANDN U2035 ( .B(\stack[1][0] ), .A(n4129), .Z(n5527) );
  OR U2036 ( .A(n5526), .B(n5527), .Z(n1800) );
  AND U2037 ( .A(n1801), .B(n1800), .Z(n1803) );
  OR U2038 ( .A(n1802), .B(n1803), .Z(n1821) );
  XNOR U2039 ( .A(n1803), .B(n1802), .Z(n5488) );
  OR U2040 ( .A(n1805), .B(n1804), .Z(n1809) );
  OR U2041 ( .A(n1807), .B(n1806), .Z(n1808) );
  NAND U2042 ( .A(n1809), .B(n1808), .Z(n1823) );
  NANDN U2043 ( .A(n1811), .B(n1810), .Z(n1812) );
  NAND U2044 ( .A(\stack[1][2] ), .B(o[2]), .Z(n5606) );
  NAND U2045 ( .A(n1812), .B(n5606), .Z(n1816) );
  OR U2046 ( .A(n1814), .B(n1813), .Z(n1815) );
  AND U2047 ( .A(n1816), .B(n1815), .Z(n1839) );
  ANDN U2048 ( .B(o[3]), .A(n1607), .Z(n1840) );
  XNOR U2049 ( .A(n1839), .B(n1840), .Z(n1842) );
  AND U2050 ( .A(\stack[1][4] ), .B(o[1]), .Z(n1817) );
  AND U2051 ( .A(o[0]), .B(\stack[1][5] ), .Z(n1901) );
  XOR U2052 ( .A(n1817), .B(n1901), .Z(n1835) );
  NAND U2053 ( .A(o[1]), .B(\stack[1][4] ), .Z(n1832) );
  NANDN U2054 ( .A(n1832), .B(o[0]), .Z(n1818) );
  XNOR U2055 ( .A(o[2]), .B(n1818), .Z(n1819) );
  NAND U2056 ( .A(\stack[1][3] ), .B(n1819), .Z(n1836) );
  XNOR U2057 ( .A(n1835), .B(n1836), .Z(n1841) );
  XOR U2058 ( .A(n1842), .B(n1841), .Z(n1822) );
  XOR U2059 ( .A(n1823), .B(n1822), .Z(n1824) );
  NAND U2060 ( .A(\stack[1][1] ), .B(o[4]), .Z(n1825) );
  XNOR U2061 ( .A(n1824), .B(n1825), .Z(n5489) );
  OR U2062 ( .A(n5488), .B(n5489), .Z(n1820) );
  AND U2063 ( .A(n1821), .B(n1820), .Z(n1846) );
  ANDN U2064 ( .B(o[5]), .A(n4195), .Z(n1851) );
  OR U2065 ( .A(n1823), .B(n1822), .Z(n1827) );
  NANDN U2066 ( .A(n1825), .B(n1824), .Z(n1826) );
  NAND U2067 ( .A(n1827), .B(n1826), .Z(n1852) );
  XNOR U2068 ( .A(n1851), .B(n1852), .Z(n1854) );
  AND U2069 ( .A(\stack[1][5] ), .B(o[1]), .Z(n1828) );
  AND U2070 ( .A(o[0]), .B(\stack[1][6] ), .Z(n1943) );
  XNOR U2071 ( .A(n1828), .B(n1943), .Z(n1863) );
  NAND U2072 ( .A(o[1]), .B(\stack[1][5] ), .Z(n1865) );
  NANDN U2073 ( .A(n1865), .B(o[0]), .Z(n1829) );
  XNOR U2074 ( .A(o[2]), .B(n1829), .Z(n1830) );
  ANDN U2075 ( .B(n1830), .A(n1609), .Z(n1862) );
  XOR U2076 ( .A(n1863), .B(n1862), .Z(n1859) );
  ANDN U2077 ( .B(o[3]), .A(n1608), .Z(n5570) );
  NANDN U2078 ( .A(n1832), .B(n1831), .Z(n1834) );
  NAND U2079 ( .A(\stack[1][3] ), .B(o[2]), .Z(n1833) );
  AND U2080 ( .A(n1834), .B(n1833), .Z(n1838) );
  OR U2081 ( .A(n1836), .B(n1835), .Z(n1837) );
  NANDN U2082 ( .A(n1838), .B(n1837), .Z(n1857) );
  XNOR U2083 ( .A(n1859), .B(n1858), .Z(n1873) );
  OR U2084 ( .A(n1840), .B(n1839), .Z(n1844) );
  OR U2085 ( .A(n1842), .B(n1841), .Z(n1843) );
  AND U2086 ( .A(n1844), .B(n1843), .Z(n1874) );
  XNOR U2087 ( .A(n1873), .B(n1874), .Z(n1876) );
  ANDN U2088 ( .B(o[4]), .A(n1607), .Z(n1875) );
  XOR U2089 ( .A(n1876), .B(n1875), .Z(n1853) );
  NANDN U2090 ( .A(n1846), .B(n1845), .Z(n1848) );
  XOR U2091 ( .A(n1846), .B(n1845), .Z(n5449) );
  IV U2092 ( .A(o[6]), .Z(n4137) );
  ANDN U2093 ( .B(\stack[1][0] ), .A(n4137), .Z(n5450) );
  OR U2094 ( .A(n5449), .B(n5450), .Z(n1847) );
  AND U2095 ( .A(n1848), .B(n1847), .Z(n1850) );
  OR U2096 ( .A(n1849), .B(n1850), .Z(n1880) );
  XNOR U2097 ( .A(n1850), .B(n1849), .Z(n5410) );
  NAND U2098 ( .A(\stack[1][1] ), .B(o[6]), .Z(n1884) );
  OR U2099 ( .A(n1852), .B(n1851), .Z(n1856) );
  NANDN U2100 ( .A(n1854), .B(n1853), .Z(n1855) );
  NAND U2101 ( .A(n1856), .B(n1855), .Z(n1882) );
  NANDN U2102 ( .A(n1857), .B(n5570), .Z(n1861) );
  NANDN U2103 ( .A(n1859), .B(n1858), .Z(n1860) );
  AND U2104 ( .A(n1861), .B(n1860), .Z(n1887) );
  NAND U2105 ( .A(n1863), .B(n1862), .Z(n1869) );
  NANDN U2106 ( .A(n1865), .B(n1864), .Z(n1867) );
  NAND U2107 ( .A(\stack[1][4] ), .B(o[2]), .Z(n1866) );
  AND U2108 ( .A(n1867), .B(n1866), .Z(n1868) );
  ANDN U2109 ( .B(n1869), .A(n1868), .Z(n1893) );
  ANDN U2110 ( .B(\stack[1][4] ), .A(n4127), .Z(n1894) );
  XNOR U2111 ( .A(n1893), .B(n1894), .Z(n1896) );
  AND U2112 ( .A(\stack[1][6] ), .B(o[1]), .Z(n1870) );
  AND U2113 ( .A(o[0]), .B(\stack[1][7] ), .Z(n1994) );
  XOR U2114 ( .A(n1870), .B(n1994), .Z(n1899) );
  NAND U2115 ( .A(o[1]), .B(\stack[1][6] ), .Z(n1902) );
  NANDN U2116 ( .A(n1902), .B(o[0]), .Z(n1871) );
  XNOR U2117 ( .A(o[2]), .B(n1871), .Z(n1872) );
  NAND U2118 ( .A(\stack[1][5] ), .B(n1872), .Z(n1900) );
  XNOR U2119 ( .A(n1899), .B(n1900), .Z(n1895) );
  XOR U2120 ( .A(n1896), .B(n1895), .Z(n1888) );
  XNOR U2121 ( .A(n1887), .B(n1888), .Z(n1890) );
  NAND U2122 ( .A(\stack[1][3] ), .B(o[4]), .Z(n1889) );
  XOR U2123 ( .A(n1890), .B(n1889), .Z(n1914) );
  OR U2124 ( .A(n1874), .B(n1873), .Z(n1878) );
  OR U2125 ( .A(n1876), .B(n1875), .Z(n1877) );
  AND U2126 ( .A(n1878), .B(n1877), .Z(n1911) );
  ANDN U2127 ( .B(\stack[1][2] ), .A(n4130), .Z(n1912) );
  XOR U2128 ( .A(n1911), .B(n1912), .Z(n1913) );
  XNOR U2129 ( .A(n1914), .B(n1913), .Z(n1881) );
  XNOR U2130 ( .A(n1882), .B(n1881), .Z(n1883) );
  XOR U2131 ( .A(n1884), .B(n1883), .Z(n5411) );
  OR U2132 ( .A(n5410), .B(n5411), .Z(n1879) );
  AND U2133 ( .A(n1880), .B(n1879), .Z(n1918) );
  ANDN U2134 ( .B(o[7]), .A(n4195), .Z(n1923) );
  OR U2135 ( .A(n1882), .B(n1881), .Z(n1886) );
  OR U2136 ( .A(n1884), .B(n1883), .Z(n1885) );
  NAND U2137 ( .A(n1886), .B(n1885), .Z(n1924) );
  XNOR U2138 ( .A(n1923), .B(n1924), .Z(n1926) );
  NAND U2139 ( .A(o[5]), .B(\stack[1][3] ), .Z(n1960) );
  OR U2140 ( .A(n1888), .B(n1887), .Z(n1892) );
  OR U2141 ( .A(n1890), .B(n1889), .Z(n1891) );
  AND U2142 ( .A(n1892), .B(n1891), .Z(n1959) );
  XNOR U2143 ( .A(n1960), .B(n1959), .Z(n1962) );
  OR U2144 ( .A(n1894), .B(n1893), .Z(n1898) );
  OR U2145 ( .A(n1896), .B(n1895), .Z(n1897) );
  NAND U2146 ( .A(n1898), .B(n1897), .Z(n1954) );
  OR U2147 ( .A(n1900), .B(n1899), .Z(n1906) );
  NANDN U2148 ( .A(n1902), .B(n1901), .Z(n1904) );
  NAND U2149 ( .A(\stack[1][5] ), .B(o[2]), .Z(n1903) );
  AND U2150 ( .A(n1904), .B(n1903), .Z(n1905) );
  ANDN U2151 ( .B(n1906), .A(n1905), .Z(n1935) );
  ANDN U2152 ( .B(\stack[1][5] ), .A(n4127), .Z(n1936) );
  XNOR U2153 ( .A(n1935), .B(n1936), .Z(n1938) );
  AND U2154 ( .A(o[1]), .B(\stack[1][7] ), .Z(n1908) );
  NAND U2155 ( .A(\stack[1][8] ), .B(o[0]), .Z(n1907) );
  XNOR U2156 ( .A(n1908), .B(n1907), .Z(n1941) );
  NAND U2157 ( .A(o[1]), .B(\stack[1][7] ), .Z(n1944) );
  NANDN U2158 ( .A(n1944), .B(o[0]), .Z(n1909) );
  XNOR U2159 ( .A(o[2]), .B(n1909), .Z(n1910) );
  NAND U2160 ( .A(\stack[1][6] ), .B(n1910), .Z(n1942) );
  XOR U2161 ( .A(n1941), .B(n1942), .Z(n1937) );
  XNOR U2162 ( .A(n1954), .B(n1953), .Z(n1956) );
  AND U2163 ( .A(\stack[1][4] ), .B(o[4]), .Z(n1955) );
  XOR U2164 ( .A(n1956), .B(n1955), .Z(n1961) );
  XOR U2165 ( .A(n1962), .B(n1961), .Z(n1929) );
  OR U2166 ( .A(n1912), .B(n1911), .Z(n1916) );
  NANDN U2167 ( .A(n1914), .B(n1913), .Z(n1915) );
  AND U2168 ( .A(n1916), .B(n1915), .Z(n1930) );
  XOR U2169 ( .A(n1929), .B(n1930), .Z(n1931) );
  ANDN U2170 ( .B(o[6]), .A(n1607), .Z(n1932) );
  XOR U2171 ( .A(n1926), .B(n1925), .Z(n1917) );
  NANDN U2172 ( .A(n1918), .B(n1917), .Z(n1920) );
  XOR U2173 ( .A(n1918), .B(n1917), .Z(n5372) );
  ANDN U2174 ( .B(\stack[1][0] ), .A(n1620), .Z(n5373) );
  OR U2175 ( .A(n5372), .B(n5373), .Z(n1919) );
  AND U2176 ( .A(n1920), .B(n1919), .Z(n1922) );
  OR U2177 ( .A(n1921), .B(n1922), .Z(n1966) );
  XNOR U2178 ( .A(n1922), .B(n1921), .Z(n5333) );
  NAND U2179 ( .A(\stack[1][1] ), .B(o[8]), .Z(n2012) );
  OR U2180 ( .A(n1924), .B(n1923), .Z(n1928) );
  OR U2181 ( .A(n1926), .B(n1925), .Z(n1927) );
  NAND U2182 ( .A(n1928), .B(n1927), .Z(n2010) );
  OR U2183 ( .A(n1930), .B(n1929), .Z(n1934) );
  NANDN U2184 ( .A(n1932), .B(n1931), .Z(n1933) );
  AND U2185 ( .A(n1934), .B(n1933), .Z(n1967) );
  ANDN U2186 ( .B(\stack[1][2] ), .A(n4111), .Z(n1968) );
  XNOR U2187 ( .A(n1967), .B(n1968), .Z(n1970) );
  OR U2188 ( .A(n1936), .B(n1935), .Z(n1940) );
  NANDN U2189 ( .A(n1938), .B(n1937), .Z(n1939) );
  NAND U2190 ( .A(n1940), .B(n1939), .Z(n2004) );
  OR U2191 ( .A(n1942), .B(n1941), .Z(n1948) );
  NANDN U2192 ( .A(n1944), .B(n1943), .Z(n1946) );
  NAND U2193 ( .A(\stack[1][6] ), .B(o[2]), .Z(n1945) );
  AND U2194 ( .A(n1946), .B(n1945), .Z(n1947) );
  ANDN U2195 ( .B(n1948), .A(n1947), .Z(n1985) );
  ANDN U2196 ( .B(\stack[1][6] ), .A(n4127), .Z(n1986) );
  XNOR U2197 ( .A(n1985), .B(n1986), .Z(n1988) );
  AND U2198 ( .A(o[1]), .B(\stack[1][8] ), .Z(n1950) );
  NAND U2199 ( .A(\stack[1][9] ), .B(o[0]), .Z(n1949) );
  XNOR U2200 ( .A(n1950), .B(n1949), .Z(n1992) );
  ANDN U2201 ( .B(\stack[1][8] ), .A(n1619), .Z(n1993) );
  NAND U2202 ( .A(o[0]), .B(n1993), .Z(n1951) );
  XNOR U2203 ( .A(o[2]), .B(n1951), .Z(n1952) );
  ANDN U2204 ( .B(n1952), .A(n1612), .Z(n1991) );
  XOR U2205 ( .A(n1992), .B(n1991), .Z(n1987) );
  XOR U2206 ( .A(n1988), .B(n1987), .Z(n2003) );
  XNOR U2207 ( .A(n2004), .B(n2003), .Z(n2006) );
  ANDN U2208 ( .B(o[4]), .A(n1610), .Z(n2005) );
  XNOR U2209 ( .A(n2006), .B(n2005), .Z(n1981) );
  ANDN U2210 ( .B(\stack[1][4] ), .A(n4130), .Z(n1979) );
  OR U2211 ( .A(n1954), .B(n1953), .Z(n1958) );
  NANDN U2212 ( .A(n1956), .B(n1955), .Z(n1957) );
  NAND U2213 ( .A(n1958), .B(n1957), .Z(n1980) );
  XNOR U2214 ( .A(n1979), .B(n1980), .Z(n1982) );
  XNOR U2215 ( .A(n1981), .B(n1982), .Z(n1974) );
  OR U2216 ( .A(n1960), .B(n1959), .Z(n1964) );
  OR U2217 ( .A(n1962), .B(n1961), .Z(n1963) );
  NAND U2218 ( .A(n1964), .B(n1963), .Z(n1973) );
  XNOR U2219 ( .A(n1974), .B(n1973), .Z(n1976) );
  ANDN U2220 ( .B(o[6]), .A(n1608), .Z(n1975) );
  XNOR U2221 ( .A(n1976), .B(n1975), .Z(n1969) );
  XOR U2222 ( .A(n1970), .B(n1969), .Z(n2009) );
  XOR U2223 ( .A(n2010), .B(n2009), .Z(n2011) );
  XNOR U2224 ( .A(n2012), .B(n2011), .Z(n5334) );
  OR U2225 ( .A(n5333), .B(n5334), .Z(n1965) );
  AND U2226 ( .A(n1966), .B(n1965), .Z(n2016) );
  OR U2227 ( .A(n1968), .B(n1967), .Z(n1972) );
  OR U2228 ( .A(n1970), .B(n1969), .Z(n1971) );
  NAND U2229 ( .A(n1972), .B(n1971), .Z(n2065) );
  OR U2230 ( .A(n1974), .B(n1973), .Z(n1978) );
  OR U2231 ( .A(n1976), .B(n1975), .Z(n1977) );
  AND U2232 ( .A(n1978), .B(n1977), .Z(n2027) );
  ANDN U2233 ( .B(\stack[1][3] ), .A(n4111), .Z(n2028) );
  XNOR U2234 ( .A(n2027), .B(n2028), .Z(n2030) );
  OR U2235 ( .A(n1980), .B(n1979), .Z(n1984) );
  OR U2236 ( .A(n1982), .B(n1981), .Z(n1983) );
  AND U2237 ( .A(n1984), .B(n1983), .Z(n2033) );
  OR U2238 ( .A(n1986), .B(n1985), .Z(n1990) );
  OR U2239 ( .A(n1988), .B(n1987), .Z(n1989) );
  NAND U2240 ( .A(n1990), .B(n1989), .Z(n2059) );
  NANDN U2241 ( .A(n1992), .B(n1991), .Z(n1998) );
  NAND U2242 ( .A(n1994), .B(n1993), .Z(n1996) );
  NAND U2243 ( .A(\stack[1][7] ), .B(o[2]), .Z(n1995) );
  AND U2244 ( .A(n1996), .B(n1995), .Z(n1997) );
  ANDN U2245 ( .B(n1998), .A(n1997), .Z(n2045) );
  ANDN U2246 ( .B(\stack[1][7] ), .A(n4127), .Z(n2046) );
  XNOR U2247 ( .A(n2045), .B(n2046), .Z(n2048) );
  AND U2248 ( .A(o[1]), .B(\stack[1][9] ), .Z(n2000) );
  NAND U2249 ( .A(\stack[1][10] ), .B(o[0]), .Z(n1999) );
  XNOR U2250 ( .A(n2000), .B(n1999), .Z(n2052) );
  ANDN U2251 ( .B(\stack[1][9] ), .A(n1619), .Z(n2053) );
  NAND U2252 ( .A(o[0]), .B(n2053), .Z(n2001) );
  XNOR U2253 ( .A(o[2]), .B(n2001), .Z(n2002) );
  ANDN U2254 ( .B(n2002), .A(n1613), .Z(n2051) );
  XOR U2255 ( .A(n2052), .B(n2051), .Z(n2047) );
  XOR U2256 ( .A(n2048), .B(n2047), .Z(n2058) );
  XNOR U2257 ( .A(n2059), .B(n2058), .Z(n2061) );
  ANDN U2258 ( .B(\stack[1][6] ), .A(n4129), .Z(n2060) );
  XNOR U2259 ( .A(n2061), .B(n2060), .Z(n2041) );
  ANDN U2260 ( .B(\stack[1][5] ), .A(n4130), .Z(n2039) );
  OR U2261 ( .A(n2004), .B(n2003), .Z(n2008) );
  NANDN U2262 ( .A(n2006), .B(n2005), .Z(n2007) );
  NAND U2263 ( .A(n2008), .B(n2007), .Z(n2040) );
  XNOR U2264 ( .A(n2039), .B(n2040), .Z(n2042) );
  XNOR U2265 ( .A(n2041), .B(n2042), .Z(n2034) );
  XOR U2266 ( .A(n2033), .B(n2034), .Z(n2035) );
  ANDN U2267 ( .B(o[6]), .A(n1609), .Z(n2036) );
  XOR U2268 ( .A(n2035), .B(n2036), .Z(n2029) );
  XOR U2269 ( .A(n2030), .B(n2029), .Z(n2064) );
  XOR U2270 ( .A(n2065), .B(n2064), .Z(n2066) );
  NAND U2271 ( .A(\stack[1][2] ), .B(o[8]), .Z(n2067) );
  ANDN U2272 ( .B(o[9]), .A(n4195), .Z(n2021) );
  OR U2273 ( .A(n2010), .B(n2009), .Z(n2014) );
  NANDN U2274 ( .A(n2012), .B(n2011), .Z(n2013) );
  NAND U2275 ( .A(n2014), .B(n2013), .Z(n2022) );
  XNOR U2276 ( .A(n2021), .B(n2022), .Z(n2024) );
  XOR U2277 ( .A(n2023), .B(n2024), .Z(n2015) );
  NANDN U2278 ( .A(n2016), .B(n2015), .Z(n2018) );
  XOR U2279 ( .A(n2016), .B(n2015), .Z(n5295) );
  ANDN U2280 ( .B(\stack[1][0] ), .A(n1621), .Z(n5296) );
  OR U2281 ( .A(n5295), .B(n5296), .Z(n2017) );
  AND U2282 ( .A(n2018), .B(n2017), .Z(n2020) );
  OR U2283 ( .A(n2019), .B(n2020), .Z(n2071) );
  XNOR U2284 ( .A(n2020), .B(n2019), .Z(n5256) );
  NAND U2285 ( .A(\stack[1][1] ), .B(o[10]), .Z(n2124) );
  OR U2286 ( .A(n2022), .B(n2021), .Z(n2026) );
  OR U2287 ( .A(n2024), .B(n2023), .Z(n2025) );
  NAND U2288 ( .A(n2026), .B(n2025), .Z(n2122) );
  NAND U2289 ( .A(\stack[1][3] ), .B(o[8]), .Z(n2118) );
  OR U2290 ( .A(n2028), .B(n2027), .Z(n2032) );
  OR U2291 ( .A(n2030), .B(n2029), .Z(n2031) );
  NAND U2292 ( .A(n2032), .B(n2031), .Z(n2116) );
  OR U2293 ( .A(n2034), .B(n2033), .Z(n2038) );
  NANDN U2294 ( .A(n2036), .B(n2035), .Z(n2037) );
  AND U2295 ( .A(n2038), .B(n2037), .Z(n2078) );
  ANDN U2296 ( .B(\stack[1][4] ), .A(n4111), .Z(n2079) );
  XNOR U2297 ( .A(n2078), .B(n2079), .Z(n2081) );
  OR U2298 ( .A(n2040), .B(n2039), .Z(n2044) );
  OR U2299 ( .A(n2042), .B(n2041), .Z(n2043) );
  AND U2300 ( .A(n2044), .B(n2043), .Z(n2084) );
  OR U2301 ( .A(n2046), .B(n2045), .Z(n2050) );
  OR U2302 ( .A(n2048), .B(n2047), .Z(n2049) );
  NAND U2303 ( .A(n2050), .B(n2049), .Z(n2110) );
  ANDN U2304 ( .B(\stack[1][8] ), .A(n4127), .Z(n2097) );
  XNOR U2305 ( .A(n2096), .B(n2097), .Z(n2099) );
  AND U2306 ( .A(o[1]), .B(\stack[1][10] ), .Z(n2055) );
  NAND U2307 ( .A(\stack[1][11] ), .B(o[0]), .Z(n2054) );
  XNOR U2308 ( .A(n2055), .B(n2054), .Z(n2103) );
  ANDN U2309 ( .B(\stack[1][10] ), .A(n1619), .Z(n2104) );
  NAND U2310 ( .A(o[0]), .B(n2104), .Z(n2056) );
  XNOR U2311 ( .A(o[2]), .B(n2056), .Z(n2057) );
  ANDN U2312 ( .B(n2057), .A(n1614), .Z(n2102) );
  XOR U2313 ( .A(n2103), .B(n2102), .Z(n2098) );
  XOR U2314 ( .A(n2099), .B(n2098), .Z(n2109) );
  XNOR U2315 ( .A(n2110), .B(n2109), .Z(n2112) );
  ANDN U2316 ( .B(\stack[1][7] ), .A(n4129), .Z(n2111) );
  XNOR U2317 ( .A(n2112), .B(n2111), .Z(n2092) );
  ANDN U2318 ( .B(\stack[1][6] ), .A(n4130), .Z(n2090) );
  OR U2319 ( .A(n2059), .B(n2058), .Z(n2063) );
  NANDN U2320 ( .A(n2061), .B(n2060), .Z(n2062) );
  NAND U2321 ( .A(n2063), .B(n2062), .Z(n2091) );
  XNOR U2322 ( .A(n2090), .B(n2091), .Z(n2093) );
  XNOR U2323 ( .A(n2092), .B(n2093), .Z(n2085) );
  XOR U2324 ( .A(n2084), .B(n2085), .Z(n2086) );
  ANDN U2325 ( .B(o[6]), .A(n1610), .Z(n2087) );
  XOR U2326 ( .A(n2086), .B(n2087), .Z(n2080) );
  XOR U2327 ( .A(n2081), .B(n2080), .Z(n2115) );
  XOR U2328 ( .A(n2116), .B(n2115), .Z(n2117) );
  ANDN U2329 ( .B(\stack[1][2] ), .A(n3977), .Z(n2072) );
  OR U2330 ( .A(n2065), .B(n2064), .Z(n2069) );
  NANDN U2331 ( .A(n2067), .B(n2066), .Z(n2068) );
  NAND U2332 ( .A(n2069), .B(n2068), .Z(n2073) );
  XOR U2333 ( .A(n2072), .B(n2073), .Z(n2074) );
  XNOR U2334 ( .A(n2075), .B(n2074), .Z(n2121) );
  XNOR U2335 ( .A(n2122), .B(n2121), .Z(n2123) );
  XOR U2336 ( .A(n2124), .B(n2123), .Z(n5257) );
  OR U2337 ( .A(n5256), .B(n5257), .Z(n2070) );
  AND U2338 ( .A(n2071), .B(n2070), .Z(n2128) );
  NAND U2339 ( .A(\stack[1][2] ), .B(o[10]), .Z(n2190) );
  OR U2340 ( .A(n2073), .B(n2072), .Z(n2077) );
  NANDN U2341 ( .A(n2075), .B(n2074), .Z(n2076) );
  NAND U2342 ( .A(n2077), .B(n2076), .Z(n2188) );
  NAND U2343 ( .A(\stack[1][4] ), .B(o[8]), .Z(n2184) );
  OR U2344 ( .A(n2079), .B(n2078), .Z(n2083) );
  OR U2345 ( .A(n2081), .B(n2080), .Z(n2082) );
  NAND U2346 ( .A(n2083), .B(n2082), .Z(n2182) );
  OR U2347 ( .A(n2085), .B(n2084), .Z(n2089) );
  NANDN U2348 ( .A(n2087), .B(n2086), .Z(n2088) );
  AND U2349 ( .A(n2089), .B(n2088), .Z(n2145) );
  ANDN U2350 ( .B(\stack[1][5] ), .A(n4111), .Z(n2146) );
  XNOR U2351 ( .A(n2145), .B(n2146), .Z(n2148) );
  ANDN U2352 ( .B(o[6]), .A(n1611), .Z(n5452) );
  OR U2353 ( .A(n2091), .B(n2090), .Z(n2095) );
  OR U2354 ( .A(n2093), .B(n2092), .Z(n2094) );
  AND U2355 ( .A(n2095), .B(n2094), .Z(n2152) );
  OR U2356 ( .A(n2097), .B(n2096), .Z(n2101) );
  OR U2357 ( .A(n2099), .B(n2098), .Z(n2100) );
  NAND U2358 ( .A(n2101), .B(n2100), .Z(n2176) );
  ANDN U2359 ( .B(\stack[1][9] ), .A(n4127), .Z(n2163) );
  XNOR U2360 ( .A(n2162), .B(n2163), .Z(n2165) );
  AND U2361 ( .A(o[1]), .B(\stack[1][11] ), .Z(n2106) );
  NAND U2362 ( .A(\stack[1][12] ), .B(o[0]), .Z(n2105) );
  XNOR U2363 ( .A(n2106), .B(n2105), .Z(n2169) );
  ANDN U2364 ( .B(\stack[1][11] ), .A(n1619), .Z(n2170) );
  NAND U2365 ( .A(o[0]), .B(n2170), .Z(n2107) );
  XNOR U2366 ( .A(o[2]), .B(n2107), .Z(n2108) );
  ANDN U2367 ( .B(n2108), .A(n1615), .Z(n2168) );
  XOR U2368 ( .A(n2169), .B(n2168), .Z(n2164) );
  XOR U2369 ( .A(n2165), .B(n2164), .Z(n2175) );
  XNOR U2370 ( .A(n2176), .B(n2175), .Z(n2178) );
  AND U2371 ( .A(o[4]), .B(\stack[1][8] ), .Z(n2177) );
  XNOR U2372 ( .A(n2178), .B(n2177), .Z(n2159) );
  NAND U2373 ( .A(\stack[1][7] ), .B(o[5]), .Z(n2156) );
  OR U2374 ( .A(n2110), .B(n2109), .Z(n2114) );
  NANDN U2375 ( .A(n2112), .B(n2111), .Z(n2113) );
  NAND U2376 ( .A(n2114), .B(n2113), .Z(n2157) );
  XOR U2377 ( .A(n2156), .B(n2157), .Z(n2158) );
  XOR U2378 ( .A(n2159), .B(n2158), .Z(n2151) );
  XOR U2379 ( .A(n2152), .B(n2151), .Z(n2153) );
  XOR U2380 ( .A(n5452), .B(n2153), .Z(n2147) );
  XOR U2381 ( .A(n2182), .B(n2181), .Z(n2183) );
  XOR U2382 ( .A(n2184), .B(n2183), .Z(n2142) );
  ANDN U2383 ( .B(\stack[1][3] ), .A(n3977), .Z(n2139) );
  OR U2384 ( .A(n2116), .B(n2115), .Z(n2120) );
  NANDN U2385 ( .A(n2118), .B(n2117), .Z(n2119) );
  NAND U2386 ( .A(n2120), .B(n2119), .Z(n2140) );
  XOR U2387 ( .A(n2139), .B(n2140), .Z(n2141) );
  XNOR U2388 ( .A(n2142), .B(n2141), .Z(n2187) );
  XNOR U2389 ( .A(n2188), .B(n2187), .Z(n2189) );
  XOR U2390 ( .A(n2190), .B(n2189), .Z(n2135) );
  ANDN U2391 ( .B(o[11]), .A(n4195), .Z(n2133) );
  OR U2392 ( .A(n2122), .B(n2121), .Z(n2126) );
  OR U2393 ( .A(n2124), .B(n2123), .Z(n2125) );
  NAND U2394 ( .A(n2126), .B(n2125), .Z(n2134) );
  XNOR U2395 ( .A(n2133), .B(n2134), .Z(n2136) );
  XOR U2396 ( .A(n2135), .B(n2136), .Z(n2127) );
  NANDN U2397 ( .A(n2128), .B(n2127), .Z(n2130) );
  XOR U2398 ( .A(n2128), .B(n2127), .Z(n5218) );
  IV U2399 ( .A(o[12]), .Z(n3990) );
  ANDN U2400 ( .B(\stack[1][0] ), .A(n3990), .Z(n5219) );
  OR U2401 ( .A(n5218), .B(n5219), .Z(n2129) );
  AND U2402 ( .A(n2130), .B(n2129), .Z(n2132) );
  OR U2403 ( .A(n2131), .B(n2132), .Z(n2194) );
  XNOR U2404 ( .A(n2132), .B(n2131), .Z(n5180) );
  NAND U2405 ( .A(\stack[1][1] ), .B(o[12]), .Z(n2259) );
  OR U2406 ( .A(n2134), .B(n2133), .Z(n2138) );
  OR U2407 ( .A(n2136), .B(n2135), .Z(n2137) );
  NAND U2408 ( .A(n2138), .B(n2137), .Z(n2257) );
  NAND U2409 ( .A(\stack[1][3] ), .B(o[10]), .Z(n2204) );
  OR U2410 ( .A(n2140), .B(n2139), .Z(n2144) );
  NANDN U2411 ( .A(n2142), .B(n2141), .Z(n2143) );
  NAND U2412 ( .A(n2144), .B(n2143), .Z(n2202) );
  NAND U2413 ( .A(\stack[1][5] ), .B(o[8]), .Z(n2253) );
  OR U2414 ( .A(n2146), .B(n2145), .Z(n2150) );
  NANDN U2415 ( .A(n2148), .B(n2147), .Z(n2149) );
  NAND U2416 ( .A(n2150), .B(n2149), .Z(n2251) );
  NANDN U2417 ( .A(n2152), .B(n2151), .Z(n2155) );
  OR U2418 ( .A(n5452), .B(n2153), .Z(n2154) );
  AND U2419 ( .A(n2155), .B(n2154), .Z(n2213) );
  ANDN U2420 ( .B(\stack[1][6] ), .A(n4111), .Z(n2214) );
  XNOR U2421 ( .A(n2213), .B(n2214), .Z(n2216) );
  NANDN U2422 ( .A(n2157), .B(n2156), .Z(n2161) );
  OR U2423 ( .A(n2159), .B(n2158), .Z(n2160) );
  AND U2424 ( .A(n2161), .B(n2160), .Z(n2219) );
  OR U2425 ( .A(n2163), .B(n2162), .Z(n2167) );
  OR U2426 ( .A(n2165), .B(n2164), .Z(n2166) );
  NAND U2427 ( .A(n2167), .B(n2166), .Z(n2245) );
  ANDN U2428 ( .B(\stack[1][10] ), .A(n4127), .Z(n2232) );
  XNOR U2429 ( .A(n2231), .B(n2232), .Z(n2234) );
  AND U2430 ( .A(o[1]), .B(\stack[1][12] ), .Z(n2172) );
  NAND U2431 ( .A(\stack[1][13] ), .B(o[0]), .Z(n2171) );
  XNOR U2432 ( .A(n2172), .B(n2171), .Z(n2238) );
  ANDN U2433 ( .B(\stack[1][12] ), .A(n1619), .Z(n2239) );
  NAND U2434 ( .A(o[0]), .B(n2239), .Z(n2173) );
  XNOR U2435 ( .A(o[2]), .B(n2173), .Z(n2174) );
  ANDN U2436 ( .B(n2174), .A(n1616), .Z(n2237) );
  XOR U2437 ( .A(n2238), .B(n2237), .Z(n2233) );
  XOR U2438 ( .A(n2234), .B(n2233), .Z(n2244) );
  XNOR U2439 ( .A(n2245), .B(n2244), .Z(n2247) );
  ANDN U2440 ( .B(\stack[1][9] ), .A(n4129), .Z(n2246) );
  XNOR U2441 ( .A(n2247), .B(n2246), .Z(n2227) );
  ANDN U2442 ( .B(\stack[1][8] ), .A(n4130), .Z(n2225) );
  OR U2443 ( .A(n2176), .B(n2175), .Z(n2180) );
  NANDN U2444 ( .A(n2178), .B(n2177), .Z(n2179) );
  NAND U2445 ( .A(n2180), .B(n2179), .Z(n2226) );
  XNOR U2446 ( .A(n2225), .B(n2226), .Z(n2228) );
  XNOR U2447 ( .A(n2227), .B(n2228), .Z(n2220) );
  XOR U2448 ( .A(n2219), .B(n2220), .Z(n2221) );
  ANDN U2449 ( .B(o[6]), .A(n1612), .Z(n2222) );
  XOR U2450 ( .A(n2221), .B(n2222), .Z(n2215) );
  XOR U2451 ( .A(n2216), .B(n2215), .Z(n2250) );
  XNOR U2452 ( .A(n2251), .B(n2250), .Z(n2252) );
  XNOR U2453 ( .A(n2253), .B(n2252), .Z(n2209) );
  NAND U2454 ( .A(\stack[1][4] ), .B(o[9]), .Z(n2207) );
  NANDN U2455 ( .A(n2182), .B(n2181), .Z(n2186) );
  OR U2456 ( .A(n2184), .B(n2183), .Z(n2185) );
  NAND U2457 ( .A(n2186), .B(n2185), .Z(n2208) );
  XOR U2458 ( .A(n2207), .B(n2208), .Z(n2210) );
  XNOR U2459 ( .A(n2209), .B(n2210), .Z(n2201) );
  XOR U2460 ( .A(n2202), .B(n2201), .Z(n2203) );
  ANDN U2461 ( .B(\stack[1][2] ), .A(n4144), .Z(n2195) );
  OR U2462 ( .A(n2188), .B(n2187), .Z(n2192) );
  OR U2463 ( .A(n2190), .B(n2189), .Z(n2191) );
  NAND U2464 ( .A(n2192), .B(n2191), .Z(n2196) );
  XOR U2465 ( .A(n2195), .B(n2196), .Z(n2197) );
  XNOR U2466 ( .A(n2198), .B(n2197), .Z(n2256) );
  XNOR U2467 ( .A(n2257), .B(n2256), .Z(n2258) );
  XOR U2468 ( .A(n2259), .B(n2258), .Z(n5181) );
  OR U2469 ( .A(n5180), .B(n5181), .Z(n2193) );
  AND U2470 ( .A(n2194), .B(n2193), .Z(n2263) );
  ANDN U2471 ( .B(o[12]), .A(n1607), .Z(n2274) );
  OR U2472 ( .A(n2196), .B(n2195), .Z(n2200) );
  NANDN U2473 ( .A(n2198), .B(n2197), .Z(n2199) );
  AND U2474 ( .A(n2200), .B(n2199), .Z(n2272) );
  ANDN U2475 ( .B(\stack[1][3] ), .A(n4144), .Z(n2332) );
  OR U2476 ( .A(n2202), .B(n2201), .Z(n2206) );
  NANDN U2477 ( .A(n2204), .B(n2203), .Z(n2205) );
  NAND U2478 ( .A(n2206), .B(n2205), .Z(n2333) );
  XNOR U2479 ( .A(n2332), .B(n2333), .Z(n2335) );
  NANDN U2480 ( .A(n2208), .B(n2207), .Z(n2212) );
  NANDN U2481 ( .A(n2210), .B(n2209), .Z(n2211) );
  AND U2482 ( .A(n2212), .B(n2211), .Z(n2278) );
  OR U2483 ( .A(n2214), .B(n2213), .Z(n2218) );
  OR U2484 ( .A(n2216), .B(n2215), .Z(n2217) );
  NAND U2485 ( .A(n2218), .B(n2217), .Z(n2327) );
  ANDN U2486 ( .B(\stack[1][7] ), .A(n4111), .Z(n5416) );
  OR U2487 ( .A(n2220), .B(n2219), .Z(n2224) );
  NANDN U2488 ( .A(n2222), .B(n2221), .Z(n2223) );
  AND U2489 ( .A(n2224), .B(n2223), .Z(n2290) );
  XNOR U2490 ( .A(n5416), .B(n2290), .Z(n2292) );
  OR U2491 ( .A(n2226), .B(n2225), .Z(n2230) );
  OR U2492 ( .A(n2228), .B(n2227), .Z(n2229) );
  AND U2493 ( .A(n2230), .B(n2229), .Z(n2295) );
  OR U2494 ( .A(n2232), .B(n2231), .Z(n2236) );
  OR U2495 ( .A(n2234), .B(n2233), .Z(n2235) );
  NAND U2496 ( .A(n2236), .B(n2235), .Z(n2321) );
  ANDN U2497 ( .B(\stack[1][11] ), .A(n4127), .Z(n2308) );
  XNOR U2498 ( .A(n2307), .B(n2308), .Z(n2310) );
  AND U2499 ( .A(o[1]), .B(\stack[1][13] ), .Z(n2241) );
  NAND U2500 ( .A(\stack[1][14] ), .B(o[0]), .Z(n2240) );
  XNOR U2501 ( .A(n2241), .B(n2240), .Z(n2314) );
  ANDN U2502 ( .B(\stack[1][13] ), .A(n1619), .Z(n2315) );
  NAND U2503 ( .A(o[0]), .B(n2315), .Z(n2242) );
  XNOR U2504 ( .A(o[2]), .B(n2242), .Z(n2243) );
  ANDN U2505 ( .B(n2243), .A(n1617), .Z(n2313) );
  XOR U2506 ( .A(n2314), .B(n2313), .Z(n2309) );
  XOR U2507 ( .A(n2310), .B(n2309), .Z(n2320) );
  XNOR U2508 ( .A(n2321), .B(n2320), .Z(n2323) );
  ANDN U2509 ( .B(\stack[1][10] ), .A(n4129), .Z(n2322) );
  XNOR U2510 ( .A(n2323), .B(n2322), .Z(n2303) );
  ANDN U2511 ( .B(\stack[1][9] ), .A(n4130), .Z(n2301) );
  OR U2512 ( .A(n2245), .B(n2244), .Z(n2249) );
  NANDN U2513 ( .A(n2247), .B(n2246), .Z(n2248) );
  NAND U2514 ( .A(n2249), .B(n2248), .Z(n2302) );
  XNOR U2515 ( .A(n2301), .B(n2302), .Z(n2304) );
  XNOR U2516 ( .A(n2303), .B(n2304), .Z(n2296) );
  XOR U2517 ( .A(n2295), .B(n2296), .Z(n2297) );
  ANDN U2518 ( .B(\stack[1][8] ), .A(n4137), .Z(n2298) );
  XOR U2519 ( .A(n2292), .B(n2291), .Z(n2326) );
  XNOR U2520 ( .A(n2327), .B(n2326), .Z(n2329) );
  ANDN U2521 ( .B(o[8]), .A(n1611), .Z(n2328) );
  XNOR U2522 ( .A(n2329), .B(n2328), .Z(n2286) );
  ANDN U2523 ( .B(\stack[1][5] ), .A(n3977), .Z(n2284) );
  OR U2524 ( .A(n2251), .B(n2250), .Z(n2255) );
  OR U2525 ( .A(n2253), .B(n2252), .Z(n2254) );
  NAND U2526 ( .A(n2255), .B(n2254), .Z(n2285) );
  XNOR U2527 ( .A(n2284), .B(n2285), .Z(n2287) );
  XNOR U2528 ( .A(n2286), .B(n2287), .Z(n2279) );
  XOR U2529 ( .A(n2278), .B(n2279), .Z(n2280) );
  ANDN U2530 ( .B(o[10]), .A(n1609), .Z(n2281) );
  XNOR U2531 ( .A(n2335), .B(n2334), .Z(n2273) );
  XNOR U2532 ( .A(n2272), .B(n2273), .Z(n2275) );
  XNOR U2533 ( .A(n2274), .B(n2275), .Z(n2269) );
  ANDN U2534 ( .B(o[13]), .A(n4195), .Z(n2266) );
  OR U2535 ( .A(n2257), .B(n2256), .Z(n2261) );
  OR U2536 ( .A(n2259), .B(n2258), .Z(n2260) );
  NAND U2537 ( .A(n2261), .B(n2260), .Z(n2267) );
  XOR U2538 ( .A(n2266), .B(n2267), .Z(n2268) );
  NANDN U2539 ( .A(n2263), .B(n2262), .Z(n2265) );
  XOR U2540 ( .A(n2263), .B(n2262), .Z(n5141) );
  ANDN U2541 ( .B(o[14]), .A(n1606), .Z(n5142) );
  OR U2542 ( .A(n5141), .B(n5142), .Z(n2264) );
  AND U2543 ( .A(n2265), .B(n2264), .Z(n2339) );
  OR U2544 ( .A(n2338), .B(n2339), .Z(n2341) );
  ANDN U2545 ( .B(o[14]), .A(n4195), .Z(n2418) );
  OR U2546 ( .A(n2267), .B(n2266), .Z(n2271) );
  NANDN U2547 ( .A(n2269), .B(n2268), .Z(n2270) );
  AND U2548 ( .A(n2271), .B(n2270), .Z(n2417) );
  OR U2549 ( .A(n2273), .B(n2272), .Z(n2277) );
  OR U2550 ( .A(n2275), .B(n2274), .Z(n2276) );
  AND U2551 ( .A(n2277), .B(n2276), .Z(n2342) );
  ANDN U2552 ( .B(\stack[1][2] ), .A(n3923), .Z(n2343) );
  XNOR U2553 ( .A(n2342), .B(n2343), .Z(n2345) );
  OR U2554 ( .A(n2279), .B(n2278), .Z(n2283) );
  NANDN U2555 ( .A(n2281), .B(n2280), .Z(n2282) );
  NAND U2556 ( .A(n2283), .B(n2282), .Z(n2349) );
  AND U2557 ( .A(o[11]), .B(\stack[1][4] ), .Z(n2348) );
  XNOR U2558 ( .A(n2349), .B(n2348), .Z(n2350) );
  NAND U2559 ( .A(\stack[1][5] ), .B(o[10]), .Z(n2407) );
  OR U2560 ( .A(n2285), .B(n2284), .Z(n2289) );
  OR U2561 ( .A(n2287), .B(n2286), .Z(n2288) );
  NAND U2562 ( .A(n2289), .B(n2288), .Z(n2405) );
  NAND U2563 ( .A(\stack[1][7] ), .B(o[8]), .Z(n2401) );
  OR U2564 ( .A(n2290), .B(n5416), .Z(n2294) );
  OR U2565 ( .A(n2292), .B(n2291), .Z(n2293) );
  NAND U2566 ( .A(n2294), .B(n2293), .Z(n2399) );
  OR U2567 ( .A(n2296), .B(n2295), .Z(n2300) );
  NANDN U2568 ( .A(n2298), .B(n2297), .Z(n2299) );
  AND U2569 ( .A(n2300), .B(n2299), .Z(n2360) );
  ANDN U2570 ( .B(\stack[1][8] ), .A(n4111), .Z(n2361) );
  XNOR U2571 ( .A(n2360), .B(n2361), .Z(n2363) );
  OR U2572 ( .A(n2302), .B(n2301), .Z(n2306) );
  OR U2573 ( .A(n2304), .B(n2303), .Z(n2305) );
  AND U2574 ( .A(n2306), .B(n2305), .Z(n2366) );
  OR U2575 ( .A(n2308), .B(n2307), .Z(n2312) );
  OR U2576 ( .A(n2310), .B(n2309), .Z(n2311) );
  NAND U2577 ( .A(n2312), .B(n2311), .Z(n2392) );
  ANDN U2578 ( .B(\stack[1][12] ), .A(n4127), .Z(n2379) );
  XNOR U2579 ( .A(n2378), .B(n2379), .Z(n2381) );
  AND U2580 ( .A(o[1]), .B(\stack[1][14] ), .Z(n2317) );
  NAND U2581 ( .A(\stack[1][15] ), .B(o[0]), .Z(n2316) );
  XNOR U2582 ( .A(n2317), .B(n2316), .Z(n2385) );
  ANDN U2583 ( .B(\stack[1][14] ), .A(n1619), .Z(n2386) );
  NAND U2584 ( .A(o[0]), .B(n2386), .Z(n2318) );
  XNOR U2585 ( .A(o[2]), .B(n2318), .Z(n2319) );
  IV U2586 ( .A(\stack[1][13] ), .Z(n3997) );
  ANDN U2587 ( .B(n2319), .A(n3997), .Z(n2384) );
  XOR U2588 ( .A(n2385), .B(n2384), .Z(n2380) );
  XOR U2589 ( .A(n2381), .B(n2380), .Z(n2391) );
  XNOR U2590 ( .A(n2392), .B(n2391), .Z(n2394) );
  ANDN U2591 ( .B(\stack[1][11] ), .A(n4129), .Z(n2393) );
  XNOR U2592 ( .A(n2394), .B(n2393), .Z(n2374) );
  ANDN U2593 ( .B(\stack[1][10] ), .A(n4130), .Z(n2372) );
  OR U2594 ( .A(n2321), .B(n2320), .Z(n2325) );
  NANDN U2595 ( .A(n2323), .B(n2322), .Z(n2324) );
  NAND U2596 ( .A(n2325), .B(n2324), .Z(n2373) );
  XNOR U2597 ( .A(n2372), .B(n2373), .Z(n2375) );
  XNOR U2598 ( .A(n2374), .B(n2375), .Z(n2367) );
  XOR U2599 ( .A(n2366), .B(n2367), .Z(n2368) );
  ANDN U2600 ( .B(\stack[1][9] ), .A(n4137), .Z(n2369) );
  XOR U2601 ( .A(n2368), .B(n2369), .Z(n2362) );
  XOR U2602 ( .A(n2363), .B(n2362), .Z(n2398) );
  XNOR U2603 ( .A(n2399), .B(n2398), .Z(n2400) );
  XNOR U2604 ( .A(n2401), .B(n2400), .Z(n2356) );
  ANDN U2605 ( .B(\stack[1][6] ), .A(n3977), .Z(n2354) );
  OR U2606 ( .A(n2327), .B(n2326), .Z(n2331) );
  NANDN U2607 ( .A(n2329), .B(n2328), .Z(n2330) );
  NAND U2608 ( .A(n2331), .B(n2330), .Z(n2355) );
  XNOR U2609 ( .A(n2354), .B(n2355), .Z(n2357) );
  XNOR U2610 ( .A(n2356), .B(n2357), .Z(n2404) );
  XNOR U2611 ( .A(n2405), .B(n2404), .Z(n2406) );
  XNOR U2612 ( .A(n2407), .B(n2406), .Z(n2351) );
  OR U2613 ( .A(n2333), .B(n2332), .Z(n2337) );
  OR U2614 ( .A(n2335), .B(n2334), .Z(n2336) );
  AND U2615 ( .A(n2337), .B(n2336), .Z(n2411) );
  XNOR U2616 ( .A(n2410), .B(n2411), .Z(n2413) );
  ANDN U2617 ( .B(o[12]), .A(n1608), .Z(n2412) );
  XOR U2618 ( .A(n2413), .B(n2412), .Z(n2344) );
  XOR U2619 ( .A(n2417), .B(n2416), .Z(n2419) );
  XNOR U2620 ( .A(n2418), .B(n2419), .Z(n5104) );
  XNOR U2621 ( .A(n2339), .B(n2338), .Z(n5105) );
  OR U2622 ( .A(n5104), .B(n5105), .Z(n2340) );
  AND U2623 ( .A(n2341), .B(n2340), .Z(n2423) );
  NAND U2624 ( .A(\stack[1][2] ), .B(o[14]), .Z(n2510) );
  OR U2625 ( .A(n2343), .B(n2342), .Z(n2347) );
  NANDN U2626 ( .A(n2345), .B(n2344), .Z(n2346) );
  NAND U2627 ( .A(n2347), .B(n2346), .Z(n2508) );
  NAND U2628 ( .A(\stack[1][4] ), .B(o[12]), .Z(n2504) );
  NANDN U2629 ( .A(n2349), .B(n2348), .Z(n2353) );
  NANDN U2630 ( .A(n2351), .B(n2350), .Z(n2352) );
  AND U2631 ( .A(n2353), .B(n2352), .Z(n2501) );
  NAND U2632 ( .A(\stack[1][6] ), .B(o[10]), .Z(n2498) );
  OR U2633 ( .A(n2355), .B(n2354), .Z(n2359) );
  NANDN U2634 ( .A(n2357), .B(n2356), .Z(n2358) );
  NAND U2635 ( .A(n2359), .B(n2358), .Z(n2496) );
  OR U2636 ( .A(n2361), .B(n2360), .Z(n2365) );
  OR U2637 ( .A(n2363), .B(n2362), .Z(n2364) );
  NAND U2638 ( .A(n2365), .B(n2364), .Z(n2490) );
  OR U2639 ( .A(n2367), .B(n2366), .Z(n2371) );
  NANDN U2640 ( .A(n2369), .B(n2368), .Z(n2370) );
  AND U2641 ( .A(n2371), .B(n2370), .Z(n2452) );
  ANDN U2642 ( .B(\stack[1][9] ), .A(n4111), .Z(n2453) );
  XNOR U2643 ( .A(n2452), .B(n2453), .Z(n2455) );
  OR U2644 ( .A(n2373), .B(n2372), .Z(n2377) );
  OR U2645 ( .A(n2375), .B(n2374), .Z(n2376) );
  AND U2646 ( .A(n2377), .B(n2376), .Z(n2458) );
  OR U2647 ( .A(n2379), .B(n2378), .Z(n2383) );
  OR U2648 ( .A(n2381), .B(n2380), .Z(n2382) );
  NAND U2649 ( .A(n2383), .B(n2382), .Z(n2484) );
  ANDN U2650 ( .B(\stack[1][13] ), .A(n4127), .Z(n2471) );
  XNOR U2651 ( .A(n2470), .B(n2471), .Z(n2473) );
  AND U2652 ( .A(o[1]), .B(\stack[1][15] ), .Z(n2388) );
  NAND U2653 ( .A(\stack[1][16] ), .B(o[0]), .Z(n2387) );
  XNOR U2654 ( .A(n2388), .B(n2387), .Z(n2477) );
  ANDN U2655 ( .B(\stack[1][15] ), .A(n1619), .Z(n2478) );
  NAND U2656 ( .A(o[0]), .B(n2478), .Z(n2389) );
  XNOR U2657 ( .A(o[2]), .B(n2389), .Z(n2390) );
  ANDN U2658 ( .B(n2390), .A(n1618), .Z(n2476) );
  XOR U2659 ( .A(n2477), .B(n2476), .Z(n2472) );
  XOR U2660 ( .A(n2473), .B(n2472), .Z(n2483) );
  XNOR U2661 ( .A(n2484), .B(n2483), .Z(n2486) );
  ANDN U2662 ( .B(\stack[1][12] ), .A(n4129), .Z(n2485) );
  XNOR U2663 ( .A(n2486), .B(n2485), .Z(n2466) );
  ANDN U2664 ( .B(\stack[1][11] ), .A(n4130), .Z(n2464) );
  OR U2665 ( .A(n2392), .B(n2391), .Z(n2396) );
  NANDN U2666 ( .A(n2394), .B(n2393), .Z(n2395) );
  NAND U2667 ( .A(n2396), .B(n2395), .Z(n2465) );
  XNOR U2668 ( .A(n2464), .B(n2465), .Z(n2467) );
  XNOR U2669 ( .A(n2466), .B(n2467), .Z(n2459) );
  XOR U2670 ( .A(n2458), .B(n2459), .Z(n2460) );
  IV U2671 ( .A(n2460), .Z(n2397) );
  ANDN U2672 ( .B(\stack[1][10] ), .A(n4137), .Z(n2461) );
  XNOR U2673 ( .A(n2397), .B(n2461), .Z(n2454) );
  XNOR U2674 ( .A(n2455), .B(n2454), .Z(n2489) );
  XOR U2675 ( .A(n2490), .B(n2489), .Z(n2492) );
  AND U2676 ( .A(\stack[1][8] ), .B(o[8]), .Z(n2491) );
  XNOR U2677 ( .A(n2492), .B(n2491), .Z(n2449) );
  NAND U2678 ( .A(\stack[1][7] ), .B(o[9]), .Z(n2446) );
  OR U2679 ( .A(n2399), .B(n2398), .Z(n2403) );
  OR U2680 ( .A(n2401), .B(n2400), .Z(n2402) );
  NAND U2681 ( .A(n2403), .B(n2402), .Z(n2447) );
  XOR U2682 ( .A(n2446), .B(n2447), .Z(n2448) );
  XOR U2683 ( .A(n2449), .B(n2448), .Z(n2495) );
  XNOR U2684 ( .A(n2496), .B(n2495), .Z(n2497) );
  XNOR U2685 ( .A(n2498), .B(n2497), .Z(n2442) );
  ANDN U2686 ( .B(\stack[1][5] ), .A(n4144), .Z(n2440) );
  OR U2687 ( .A(n2405), .B(n2404), .Z(n2409) );
  OR U2688 ( .A(n2407), .B(n2406), .Z(n2408) );
  NAND U2689 ( .A(n2409), .B(n2408), .Z(n2441) );
  XNOR U2690 ( .A(n2440), .B(n2441), .Z(n2443) );
  XNOR U2691 ( .A(n2501), .B(n2502), .Z(n2503) );
  XNOR U2692 ( .A(n2504), .B(n2503), .Z(n2436) );
  OR U2693 ( .A(n2411), .B(n2410), .Z(n2415) );
  OR U2694 ( .A(n2413), .B(n2412), .Z(n2414) );
  AND U2695 ( .A(n2415), .B(n2414), .Z(n2435) );
  NAND U2696 ( .A(\stack[1][3] ), .B(o[13]), .Z(n2434) );
  XOR U2697 ( .A(n2435), .B(n2434), .Z(n2437) );
  XNOR U2698 ( .A(n2436), .B(n2437), .Z(n2507) );
  XOR U2699 ( .A(n2508), .B(n2507), .Z(n2509) );
  NANDN U2700 ( .A(n2417), .B(n2416), .Z(n2421) );
  OR U2701 ( .A(n2419), .B(n2418), .Z(n2420) );
  AND U2702 ( .A(n2421), .B(n2420), .Z(n2428) );
  ANDN U2703 ( .B(o[15]), .A(n4195), .Z(n2429) );
  XNOR U2704 ( .A(n2428), .B(n2429), .Z(n2431) );
  XOR U2705 ( .A(n2430), .B(n2431), .Z(n2422) );
  NANDN U2706 ( .A(n2423), .B(n2422), .Z(n2425) );
  XOR U2707 ( .A(n2423), .B(n2422), .Z(n5064) );
  OR U2708 ( .A(n5064), .B(n5065), .Z(n2424) );
  AND U2709 ( .A(n2425), .B(n2424), .Z(n2427) );
  OR U2710 ( .A(n2426), .B(n2427), .Z(n2514) );
  XNOR U2711 ( .A(n2427), .B(n2426), .Z(n5026) );
  NAND U2712 ( .A(\stack[1][1] ), .B(o[16]), .Z(n2601) );
  OR U2713 ( .A(n2429), .B(n2428), .Z(n2433) );
  OR U2714 ( .A(n2431), .B(n2430), .Z(n2432) );
  NAND U2715 ( .A(n2433), .B(n2432), .Z(n2599) );
  NAND U2716 ( .A(\stack[1][3] ), .B(o[14]), .Z(n2595) );
  NANDN U2717 ( .A(n2435), .B(n2434), .Z(n2439) );
  NANDN U2718 ( .A(n2437), .B(n2436), .Z(n2438) );
  NAND U2719 ( .A(n2439), .B(n2438), .Z(n2593) );
  NAND U2720 ( .A(\stack[1][5] ), .B(o[12]), .Z(n2589) );
  OR U2721 ( .A(n2441), .B(n2440), .Z(n2445) );
  NANDN U2722 ( .A(n2443), .B(n2442), .Z(n2444) );
  NAND U2723 ( .A(n2445), .B(n2444), .Z(n2587) );
  NAND U2724 ( .A(\stack[1][7] ), .B(o[10]), .Z(n2583) );
  NANDN U2725 ( .A(n2447), .B(n2446), .Z(n2451) );
  OR U2726 ( .A(n2449), .B(n2448), .Z(n2450) );
  NAND U2727 ( .A(n2451), .B(n2450), .Z(n2581) );
  NAND U2728 ( .A(\stack[1][9] ), .B(o[8]), .Z(n2577) );
  OR U2729 ( .A(n2453), .B(n2452), .Z(n2457) );
  OR U2730 ( .A(n2455), .B(n2454), .Z(n2456) );
  NAND U2731 ( .A(n2457), .B(n2456), .Z(n2575) );
  OR U2732 ( .A(n2459), .B(n2458), .Z(n2463) );
  NANDN U2733 ( .A(n2461), .B(n2460), .Z(n2462) );
  AND U2734 ( .A(n2463), .B(n2462), .Z(n2539) );
  ANDN U2735 ( .B(\stack[1][10] ), .A(n4111), .Z(n2540) );
  XNOR U2736 ( .A(n2539), .B(n2540), .Z(n2542) );
  OR U2737 ( .A(n2465), .B(n2464), .Z(n2469) );
  OR U2738 ( .A(n2467), .B(n2466), .Z(n2468) );
  AND U2739 ( .A(n2469), .B(n2468), .Z(n2545) );
  OR U2740 ( .A(n2471), .B(n2470), .Z(n2475) );
  OR U2741 ( .A(n2473), .B(n2472), .Z(n2474) );
  NAND U2742 ( .A(n2475), .B(n2474), .Z(n2569) );
  ANDN U2743 ( .B(\stack[1][14] ), .A(n4127), .Z(n2558) );
  XNOR U2744 ( .A(n2557), .B(n2558), .Z(n2560) );
  AND U2745 ( .A(o[1]), .B(\stack[1][16] ), .Z(n2480) );
  NAND U2746 ( .A(\stack[1][17] ), .B(o[0]), .Z(n2479) );
  XNOR U2747 ( .A(n2480), .B(n2479), .Z(n2564) );
  ANDN U2748 ( .B(\stack[1][16] ), .A(n1619), .Z(n2565) );
  NAND U2749 ( .A(o[0]), .B(n2565), .Z(n2481) );
  XNOR U2750 ( .A(o[2]), .B(n2481), .Z(n2482) );
  IV U2751 ( .A(\stack[1][15] ), .Z(n4157) );
  ANDN U2752 ( .B(n2482), .A(n4157), .Z(n2563) );
  XOR U2753 ( .A(n2564), .B(n2563), .Z(n2559) );
  XOR U2754 ( .A(n2560), .B(n2559), .Z(n2568) );
  XNOR U2755 ( .A(n2569), .B(n2568), .Z(n2571) );
  ANDN U2756 ( .B(\stack[1][13] ), .A(n4129), .Z(n2570) );
  XNOR U2757 ( .A(n2571), .B(n2570), .Z(n2553) );
  ANDN U2758 ( .B(\stack[1][12] ), .A(n4130), .Z(n2551) );
  OR U2759 ( .A(n2484), .B(n2483), .Z(n2488) );
  NANDN U2760 ( .A(n2486), .B(n2485), .Z(n2487) );
  NAND U2761 ( .A(n2488), .B(n2487), .Z(n2552) );
  XNOR U2762 ( .A(n2551), .B(n2552), .Z(n2554) );
  XNOR U2763 ( .A(n2553), .B(n2554), .Z(n2546) );
  XOR U2764 ( .A(n2545), .B(n2546), .Z(n2547) );
  ANDN U2765 ( .B(\stack[1][11] ), .A(n4137), .Z(n2548) );
  XOR U2766 ( .A(n2547), .B(n2548), .Z(n2541) );
  XOR U2767 ( .A(n2542), .B(n2541), .Z(n2574) );
  XNOR U2768 ( .A(n2575), .B(n2574), .Z(n2576) );
  XNOR U2769 ( .A(n2577), .B(n2576), .Z(n2535) );
  NAND U2770 ( .A(\stack[1][8] ), .B(o[9]), .Z(n2533) );
  NANDN U2771 ( .A(n2490), .B(n2489), .Z(n2494) );
  NANDN U2772 ( .A(n2492), .B(n2491), .Z(n2493) );
  NAND U2773 ( .A(n2494), .B(n2493), .Z(n2534) );
  XOR U2774 ( .A(n2533), .B(n2534), .Z(n2536) );
  XNOR U2775 ( .A(n2535), .B(n2536), .Z(n2580) );
  XNOR U2776 ( .A(n2581), .B(n2580), .Z(n2582) );
  XNOR U2777 ( .A(n2583), .B(n2582), .Z(n2529) );
  NAND U2778 ( .A(\stack[1][6] ), .B(o[11]), .Z(n2527) );
  OR U2779 ( .A(n2496), .B(n2495), .Z(n2500) );
  OR U2780 ( .A(n2498), .B(n2497), .Z(n2499) );
  NAND U2781 ( .A(n2500), .B(n2499), .Z(n2528) );
  XOR U2782 ( .A(n2527), .B(n2528), .Z(n2530) );
  XNOR U2783 ( .A(n2529), .B(n2530), .Z(n2586) );
  XNOR U2784 ( .A(n2587), .B(n2586), .Z(n2588) );
  XNOR U2785 ( .A(n2589), .B(n2588), .Z(n2523) );
  ANDN U2786 ( .B(\stack[1][4] ), .A(n3923), .Z(n2521) );
  OR U2787 ( .A(n2502), .B(n2501), .Z(n2506) );
  OR U2788 ( .A(n2504), .B(n2503), .Z(n2505) );
  NAND U2789 ( .A(n2506), .B(n2505), .Z(n2522) );
  XNOR U2790 ( .A(n2521), .B(n2522), .Z(n2524) );
  XNOR U2791 ( .A(n2523), .B(n2524), .Z(n2592) );
  XNOR U2792 ( .A(n2593), .B(n2592), .Z(n2594) );
  XOR U2793 ( .A(n2595), .B(n2594), .Z(n2518) );
  ANDN U2794 ( .B(o[15]), .A(n1607), .Z(n2515) );
  OR U2795 ( .A(n2508), .B(n2507), .Z(n2512) );
  NANDN U2796 ( .A(n2510), .B(n2509), .Z(n2511) );
  NAND U2797 ( .A(n2512), .B(n2511), .Z(n2516) );
  XOR U2798 ( .A(n2515), .B(n2516), .Z(n2517) );
  XNOR U2799 ( .A(n2518), .B(n2517), .Z(n2598) );
  XNOR U2800 ( .A(n2599), .B(n2598), .Z(n2600) );
  XOR U2801 ( .A(n2601), .B(n2600), .Z(n5027) );
  OR U2802 ( .A(n5026), .B(n5027), .Z(n2513) );
  AND U2803 ( .A(n2514), .B(n2513), .Z(n2605) );
  NAND U2804 ( .A(\stack[1][2] ), .B(o[16]), .Z(n2701) );
  OR U2805 ( .A(n2516), .B(n2515), .Z(n2520) );
  NANDN U2806 ( .A(n2518), .B(n2517), .Z(n2519) );
  NAND U2807 ( .A(n2520), .B(n2519), .Z(n2699) );
  NAND U2808 ( .A(\stack[1][4] ), .B(o[14]), .Z(n2695) );
  OR U2809 ( .A(n2522), .B(n2521), .Z(n2526) );
  NANDN U2810 ( .A(n2524), .B(n2523), .Z(n2525) );
  NAND U2811 ( .A(n2526), .B(n2525), .Z(n2693) );
  NAND U2812 ( .A(\stack[1][6] ), .B(o[12]), .Z(n2689) );
  NANDN U2813 ( .A(n2528), .B(n2527), .Z(n2532) );
  NANDN U2814 ( .A(n2530), .B(n2529), .Z(n2531) );
  NAND U2815 ( .A(n2532), .B(n2531), .Z(n2687) );
  NAND U2816 ( .A(\stack[1][8] ), .B(o[10]), .Z(n2683) );
  NANDN U2817 ( .A(n2534), .B(n2533), .Z(n2538) );
  NANDN U2818 ( .A(n2536), .B(n2535), .Z(n2537) );
  NAND U2819 ( .A(n2538), .B(n2537), .Z(n2681) );
  NAND U2820 ( .A(o[8]), .B(\stack[1][10] ), .Z(n2677) );
  OR U2821 ( .A(n2540), .B(n2539), .Z(n2544) );
  OR U2822 ( .A(n2542), .B(n2541), .Z(n2543) );
  NAND U2823 ( .A(n2544), .B(n2543), .Z(n2675) );
  OR U2824 ( .A(n2546), .B(n2545), .Z(n2550) );
  NANDN U2825 ( .A(n2548), .B(n2547), .Z(n2549) );
  AND U2826 ( .A(n2550), .B(n2549), .Z(n2639) );
  ANDN U2827 ( .B(\stack[1][11] ), .A(n4111), .Z(n2640) );
  XNOR U2828 ( .A(n2639), .B(n2640), .Z(n2642) );
  OR U2829 ( .A(n2552), .B(n2551), .Z(n2556) );
  OR U2830 ( .A(n2554), .B(n2553), .Z(n2555) );
  AND U2831 ( .A(n2556), .B(n2555), .Z(n2645) );
  OR U2832 ( .A(n2558), .B(n2557), .Z(n2562) );
  OR U2833 ( .A(n2560), .B(n2559), .Z(n2561) );
  NAND U2834 ( .A(n2562), .B(n2561), .Z(n2669) );
  ANDN U2835 ( .B(\stack[1][15] ), .A(n4127), .Z(n2658) );
  XNOR U2836 ( .A(n2657), .B(n2658), .Z(n2660) );
  AND U2837 ( .A(o[1]), .B(\stack[1][17] ), .Z(n2567) );
  NAND U2838 ( .A(\stack[1][18] ), .B(o[0]), .Z(n2566) );
  XNOR U2839 ( .A(n2567), .B(n2566), .Z(n2664) );
  ANDN U2840 ( .B(\stack[1][17] ), .A(n1619), .Z(n2665) );
  XOR U2841 ( .A(n2664), .B(n2663), .Z(n2659) );
  XOR U2842 ( .A(n2660), .B(n2659), .Z(n2668) );
  XNOR U2843 ( .A(n2669), .B(n2668), .Z(n2671) );
  ANDN U2844 ( .B(\stack[1][14] ), .A(n4129), .Z(n2670) );
  XNOR U2845 ( .A(n2671), .B(n2670), .Z(n2653) );
  ANDN U2846 ( .B(\stack[1][13] ), .A(n4130), .Z(n2651) );
  OR U2847 ( .A(n2569), .B(n2568), .Z(n2573) );
  NANDN U2848 ( .A(n2571), .B(n2570), .Z(n2572) );
  NAND U2849 ( .A(n2573), .B(n2572), .Z(n2652) );
  XNOR U2850 ( .A(n2651), .B(n2652), .Z(n2654) );
  XNOR U2851 ( .A(n2653), .B(n2654), .Z(n2646) );
  XOR U2852 ( .A(n2645), .B(n2646), .Z(n2647) );
  ANDN U2853 ( .B(\stack[1][12] ), .A(n4137), .Z(n2648) );
  XOR U2854 ( .A(n2647), .B(n2648), .Z(n2641) );
  XOR U2855 ( .A(n2642), .B(n2641), .Z(n2674) );
  XNOR U2856 ( .A(n2675), .B(n2674), .Z(n2676) );
  XNOR U2857 ( .A(n2677), .B(n2676), .Z(n2635) );
  ANDN U2858 ( .B(o[9]), .A(n1614), .Z(n5336) );
  OR U2859 ( .A(n2575), .B(n2574), .Z(n2579) );
  OR U2860 ( .A(n2577), .B(n2576), .Z(n2578) );
  NAND U2861 ( .A(n2579), .B(n2578), .Z(n2634) );
  XNOR U2862 ( .A(n5336), .B(n2634), .Z(n2636) );
  XNOR U2863 ( .A(n2635), .B(n2636), .Z(n2680) );
  XNOR U2864 ( .A(n2681), .B(n2680), .Z(n2682) );
  XNOR U2865 ( .A(n2683), .B(n2682), .Z(n2630) );
  NAND U2866 ( .A(\stack[1][7] ), .B(o[11]), .Z(n2628) );
  OR U2867 ( .A(n2581), .B(n2580), .Z(n2585) );
  OR U2868 ( .A(n2583), .B(n2582), .Z(n2584) );
  NAND U2869 ( .A(n2585), .B(n2584), .Z(n2629) );
  XOR U2870 ( .A(n2628), .B(n2629), .Z(n2631) );
  XNOR U2871 ( .A(n2630), .B(n2631), .Z(n2686) );
  XNOR U2872 ( .A(n2687), .B(n2686), .Z(n2688) );
  XNOR U2873 ( .A(n2689), .B(n2688), .Z(n2624) );
  NAND U2874 ( .A(\stack[1][5] ), .B(o[13]), .Z(n2622) );
  OR U2875 ( .A(n2587), .B(n2586), .Z(n2591) );
  OR U2876 ( .A(n2589), .B(n2588), .Z(n2590) );
  NAND U2877 ( .A(n2591), .B(n2590), .Z(n2623) );
  XOR U2878 ( .A(n2622), .B(n2623), .Z(n2625) );
  XNOR U2879 ( .A(n2624), .B(n2625), .Z(n2692) );
  XNOR U2880 ( .A(n2693), .B(n2692), .Z(n2694) );
  XNOR U2881 ( .A(n2695), .B(n2694), .Z(n2618) );
  NAND U2882 ( .A(\stack[1][3] ), .B(o[15]), .Z(n2616) );
  OR U2883 ( .A(n2593), .B(n2592), .Z(n2597) );
  OR U2884 ( .A(n2595), .B(n2594), .Z(n2596) );
  NAND U2885 ( .A(n2597), .B(n2596), .Z(n2617) );
  XOR U2886 ( .A(n2616), .B(n2617), .Z(n2619) );
  XNOR U2887 ( .A(n2618), .B(n2619), .Z(n2698) );
  XOR U2888 ( .A(n2699), .B(n2698), .Z(n2700) );
  ANDN U2889 ( .B(o[17]), .A(n4195), .Z(n2610) );
  OR U2890 ( .A(n2599), .B(n2598), .Z(n2603) );
  OR U2891 ( .A(n2601), .B(n2600), .Z(n2602) );
  NAND U2892 ( .A(n2603), .B(n2602), .Z(n2611) );
  XNOR U2893 ( .A(n2610), .B(n2611), .Z(n2613) );
  XOR U2894 ( .A(n2612), .B(n2613), .Z(n2604) );
  NANDN U2895 ( .A(n2605), .B(n2604), .Z(n2607) );
  XOR U2896 ( .A(n2605), .B(n2604), .Z(n4988) );
  OR U2897 ( .A(n4988), .B(n4989), .Z(n2606) );
  AND U2898 ( .A(n2607), .B(n2606), .Z(n2609) );
  OR U2899 ( .A(n2608), .B(n2609), .Z(n2705) );
  XNOR U2900 ( .A(n2609), .B(n2608), .Z(n4950) );
  NAND U2901 ( .A(\stack[1][1] ), .B(o[18]), .Z(n2804) );
  OR U2902 ( .A(n2611), .B(n2610), .Z(n2615) );
  OR U2903 ( .A(n2613), .B(n2612), .Z(n2614) );
  NAND U2904 ( .A(n2615), .B(n2614), .Z(n2802) );
  NAND U2905 ( .A(\stack[1][3] ), .B(o[16]), .Z(n2798) );
  NANDN U2906 ( .A(n2617), .B(n2616), .Z(n2621) );
  NANDN U2907 ( .A(n2619), .B(n2618), .Z(n2620) );
  NAND U2908 ( .A(n2621), .B(n2620), .Z(n2796) );
  NAND U2909 ( .A(\stack[1][5] ), .B(o[14]), .Z(n2792) );
  NANDN U2910 ( .A(n2623), .B(n2622), .Z(n2627) );
  NANDN U2911 ( .A(n2625), .B(n2624), .Z(n2626) );
  NAND U2912 ( .A(n2627), .B(n2626), .Z(n2790) );
  NAND U2913 ( .A(\stack[1][7] ), .B(o[12]), .Z(n2786) );
  NANDN U2914 ( .A(n2629), .B(n2628), .Z(n2633) );
  NANDN U2915 ( .A(n2631), .B(n2630), .Z(n2632) );
  NAND U2916 ( .A(n2633), .B(n2632), .Z(n2784) );
  NAND U2917 ( .A(\stack[1][9] ), .B(o[10]), .Z(n2733) );
  OR U2918 ( .A(n2634), .B(n5336), .Z(n2638) );
  NANDN U2919 ( .A(n2636), .B(n2635), .Z(n2637) );
  NAND U2920 ( .A(n2638), .B(n2637), .Z(n2731) );
  NAND U2921 ( .A(o[8]), .B(\stack[1][11] ), .Z(n2780) );
  OR U2922 ( .A(n2640), .B(n2639), .Z(n2644) );
  OR U2923 ( .A(n2642), .B(n2641), .Z(n2643) );
  NAND U2924 ( .A(n2644), .B(n2643), .Z(n2778) );
  OR U2925 ( .A(n2646), .B(n2645), .Z(n2650) );
  NANDN U2926 ( .A(n2648), .B(n2647), .Z(n2649) );
  AND U2927 ( .A(n2650), .B(n2649), .Z(n2742) );
  ANDN U2928 ( .B(\stack[1][12] ), .A(n4111), .Z(n2743) );
  XNOR U2929 ( .A(n2742), .B(n2743), .Z(n2745) );
  OR U2930 ( .A(n2652), .B(n2651), .Z(n2656) );
  OR U2931 ( .A(n2654), .B(n2653), .Z(n2655) );
  AND U2932 ( .A(n2656), .B(n2655), .Z(n2748) );
  OR U2933 ( .A(n2658), .B(n2657), .Z(n2662) );
  OR U2934 ( .A(n2660), .B(n2659), .Z(n2661) );
  NAND U2935 ( .A(n2662), .B(n2661), .Z(n2772) );
  ANDN U2936 ( .B(\stack[1][16] ), .A(n4127), .Z(n2761) );
  XNOR U2937 ( .A(n2760), .B(n2761), .Z(n2763) );
  AND U2938 ( .A(o[1]), .B(\stack[1][18] ), .Z(n2667) );
  NAND U2939 ( .A(\stack[1][19] ), .B(o[0]), .Z(n2666) );
  XNOR U2940 ( .A(n2667), .B(n2666), .Z(n2767) );
  ANDN U2941 ( .B(\stack[1][18] ), .A(n1619), .Z(n2768) );
  XOR U2942 ( .A(n2767), .B(n2766), .Z(n2762) );
  XOR U2943 ( .A(n2763), .B(n2762), .Z(n2771) );
  XNOR U2944 ( .A(n2772), .B(n2771), .Z(n2774) );
  ANDN U2945 ( .B(\stack[1][15] ), .A(n4129), .Z(n2773) );
  XNOR U2946 ( .A(n2774), .B(n2773), .Z(n2756) );
  ANDN U2947 ( .B(\stack[1][14] ), .A(n4130), .Z(n2754) );
  OR U2948 ( .A(n2669), .B(n2668), .Z(n2673) );
  NANDN U2949 ( .A(n2671), .B(n2670), .Z(n2672) );
  NAND U2950 ( .A(n2673), .B(n2672), .Z(n2755) );
  XNOR U2951 ( .A(n2754), .B(n2755), .Z(n2757) );
  XNOR U2952 ( .A(n2756), .B(n2757), .Z(n2749) );
  XOR U2953 ( .A(n2748), .B(n2749), .Z(n2750) );
  ANDN U2954 ( .B(\stack[1][13] ), .A(n4137), .Z(n2751) );
  XOR U2955 ( .A(n2750), .B(n2751), .Z(n2744) );
  XOR U2956 ( .A(n2745), .B(n2744), .Z(n2777) );
  XNOR U2957 ( .A(n2778), .B(n2777), .Z(n2779) );
  XNOR U2958 ( .A(n2780), .B(n2779), .Z(n2738) );
  NAND U2959 ( .A(\stack[1][10] ), .B(o[9]), .Z(n2736) );
  OR U2960 ( .A(n2675), .B(n2674), .Z(n2679) );
  OR U2961 ( .A(n2677), .B(n2676), .Z(n2678) );
  NAND U2962 ( .A(n2679), .B(n2678), .Z(n2737) );
  XOR U2963 ( .A(n2736), .B(n2737), .Z(n2739) );
  XNOR U2964 ( .A(n2738), .B(n2739), .Z(n2730) );
  XNOR U2965 ( .A(n2731), .B(n2730), .Z(n2732) );
  XNOR U2966 ( .A(n2733), .B(n2732), .Z(n2726) );
  NAND U2967 ( .A(\stack[1][8] ), .B(o[11]), .Z(n2724) );
  OR U2968 ( .A(n2681), .B(n2680), .Z(n2685) );
  OR U2969 ( .A(n2683), .B(n2682), .Z(n2684) );
  NAND U2970 ( .A(n2685), .B(n2684), .Z(n2725) );
  XOR U2971 ( .A(n2724), .B(n2725), .Z(n2727) );
  XNOR U2972 ( .A(n2726), .B(n2727), .Z(n2783) );
  XNOR U2973 ( .A(n2784), .B(n2783), .Z(n2785) );
  XNOR U2974 ( .A(n2786), .B(n2785), .Z(n2720) );
  NAND U2975 ( .A(\stack[1][6] ), .B(o[13]), .Z(n2718) );
  OR U2976 ( .A(n2687), .B(n2686), .Z(n2691) );
  OR U2977 ( .A(n2689), .B(n2688), .Z(n2690) );
  NAND U2978 ( .A(n2691), .B(n2690), .Z(n2719) );
  XOR U2979 ( .A(n2718), .B(n2719), .Z(n2721) );
  XNOR U2980 ( .A(n2720), .B(n2721), .Z(n2789) );
  XNOR U2981 ( .A(n2790), .B(n2789), .Z(n2791) );
  XNOR U2982 ( .A(n2792), .B(n2791), .Z(n2714) );
  ANDN U2983 ( .B(o[15]), .A(n1609), .Z(n2712) );
  OR U2984 ( .A(n2693), .B(n2692), .Z(n2697) );
  OR U2985 ( .A(n2695), .B(n2694), .Z(n2696) );
  NAND U2986 ( .A(n2697), .B(n2696), .Z(n2713) );
  XNOR U2987 ( .A(n2712), .B(n2713), .Z(n2715) );
  XNOR U2988 ( .A(n2714), .B(n2715), .Z(n2795) );
  XNOR U2989 ( .A(n2796), .B(n2795), .Z(n2797) );
  XOR U2990 ( .A(n2798), .B(n2797), .Z(n2709) );
  ANDN U2991 ( .B(\stack[1][2] ), .A(n3911), .Z(n2706) );
  OR U2992 ( .A(n2699), .B(n2698), .Z(n2703) );
  NANDN U2993 ( .A(n2701), .B(n2700), .Z(n2702) );
  NAND U2994 ( .A(n2703), .B(n2702), .Z(n2707) );
  XOR U2995 ( .A(n2706), .B(n2707), .Z(n2708) );
  XNOR U2996 ( .A(n2709), .B(n2708), .Z(n2801) );
  XNOR U2997 ( .A(n2802), .B(n2801), .Z(n2803) );
  XOR U2998 ( .A(n2804), .B(n2803), .Z(n4951) );
  OR U2999 ( .A(n4950), .B(n4951), .Z(n2704) );
  AND U3000 ( .A(n2705), .B(n2704), .Z(n2808) );
  NAND U3001 ( .A(\stack[1][2] ), .B(o[18]), .Z(n2917) );
  OR U3002 ( .A(n2707), .B(n2706), .Z(n2711) );
  NANDN U3003 ( .A(n2709), .B(n2708), .Z(n2710) );
  NAND U3004 ( .A(n2711), .B(n2710), .Z(n2915) );
  NAND U3005 ( .A(\stack[1][4] ), .B(o[16]), .Z(n2911) );
  OR U3006 ( .A(n2713), .B(n2712), .Z(n2717) );
  NANDN U3007 ( .A(n2715), .B(n2714), .Z(n2716) );
  NAND U3008 ( .A(n2717), .B(n2716), .Z(n2909) );
  NAND U3009 ( .A(\stack[1][6] ), .B(o[14]), .Z(n2905) );
  NANDN U3010 ( .A(n2719), .B(n2718), .Z(n2723) );
  NANDN U3011 ( .A(n2721), .B(n2720), .Z(n2722) );
  NAND U3012 ( .A(n2723), .B(n2722), .Z(n2903) );
  ANDN U3013 ( .B(o[12]), .A(n1613), .Z(n2840) );
  NANDN U3014 ( .A(n2725), .B(n2724), .Z(n2729) );
  NANDN U3015 ( .A(n2727), .B(n2726), .Z(n2728) );
  AND U3016 ( .A(n2729), .B(n2728), .Z(n2837) );
  ANDN U3017 ( .B(\stack[1][9] ), .A(n4144), .Z(n2896) );
  OR U3018 ( .A(n2731), .B(n2730), .Z(n2735) );
  OR U3019 ( .A(n2733), .B(n2732), .Z(n2734) );
  NAND U3020 ( .A(n2735), .B(n2734), .Z(n2897) );
  XNOR U3021 ( .A(n2896), .B(n2897), .Z(n2899) );
  NAND U3022 ( .A(o[10]), .B(\stack[1][10] ), .Z(n2845) );
  NANDN U3023 ( .A(n2737), .B(n2736), .Z(n2741) );
  NANDN U3024 ( .A(n2739), .B(n2738), .Z(n2740) );
  AND U3025 ( .A(n2741), .B(n2740), .Z(n2844) );
  OR U3026 ( .A(n2743), .B(n2742), .Z(n2747) );
  OR U3027 ( .A(n2745), .B(n2744), .Z(n2746) );
  NAND U3028 ( .A(n2747), .B(n2746), .Z(n2891) );
  OR U3029 ( .A(n2749), .B(n2748), .Z(n2753) );
  NANDN U3030 ( .A(n2751), .B(n2750), .Z(n2752) );
  AND U3031 ( .A(n2753), .B(n2752), .Z(n2855) );
  ANDN U3032 ( .B(\stack[1][13] ), .A(n4111), .Z(n2856) );
  XNOR U3033 ( .A(n2855), .B(n2856), .Z(n2858) );
  OR U3034 ( .A(n2755), .B(n2754), .Z(n2759) );
  OR U3035 ( .A(n2757), .B(n2756), .Z(n2758) );
  AND U3036 ( .A(n2759), .B(n2758), .Z(n2861) );
  OR U3037 ( .A(n2761), .B(n2760), .Z(n2765) );
  OR U3038 ( .A(n2763), .B(n2762), .Z(n2764) );
  NAND U3039 ( .A(n2765), .B(n2764), .Z(n2885) );
  ANDN U3040 ( .B(\stack[1][17] ), .A(n4127), .Z(n2874) );
  XNOR U3041 ( .A(n2873), .B(n2874), .Z(n2876) );
  AND U3042 ( .A(o[1]), .B(\stack[1][19] ), .Z(n2770) );
  NAND U3043 ( .A(\stack[1][20] ), .B(o[0]), .Z(n2769) );
  XNOR U3044 ( .A(n2770), .B(n2769), .Z(n2880) );
  ANDN U3045 ( .B(\stack[1][19] ), .A(n1619), .Z(n2881) );
  XOR U3046 ( .A(n2880), .B(n2879), .Z(n2875) );
  XOR U3047 ( .A(n2876), .B(n2875), .Z(n2884) );
  XNOR U3048 ( .A(n2885), .B(n2884), .Z(n2887) );
  ANDN U3049 ( .B(\stack[1][16] ), .A(n4129), .Z(n2886) );
  XNOR U3050 ( .A(n2887), .B(n2886), .Z(n2869) );
  ANDN U3051 ( .B(\stack[1][15] ), .A(n4130), .Z(n2867) );
  OR U3052 ( .A(n2772), .B(n2771), .Z(n2776) );
  NANDN U3053 ( .A(n2774), .B(n2773), .Z(n2775) );
  NAND U3054 ( .A(n2776), .B(n2775), .Z(n2868) );
  XNOR U3055 ( .A(n2867), .B(n2868), .Z(n2870) );
  XNOR U3056 ( .A(n2869), .B(n2870), .Z(n2862) );
  XOR U3057 ( .A(n2861), .B(n2862), .Z(n2863) );
  ANDN U3058 ( .B(\stack[1][14] ), .A(n4137), .Z(n2864) );
  XNOR U3059 ( .A(n2858), .B(n2857), .Z(n2890) );
  XOR U3060 ( .A(n2891), .B(n2890), .Z(n2893) );
  AND U3061 ( .A(o[8]), .B(\stack[1][12] ), .Z(n2892) );
  XNOR U3062 ( .A(n2893), .B(n2892), .Z(n2852) );
  NAND U3063 ( .A(\stack[1][11] ), .B(o[9]), .Z(n2849) );
  OR U3064 ( .A(n2778), .B(n2777), .Z(n2782) );
  OR U3065 ( .A(n2780), .B(n2779), .Z(n2781) );
  NAND U3066 ( .A(n2782), .B(n2781), .Z(n2850) );
  XOR U3067 ( .A(n2849), .B(n2850), .Z(n2851) );
  XOR U3068 ( .A(n2852), .B(n2851), .Z(n2843) );
  XOR U3069 ( .A(n2844), .B(n2843), .Z(n2846) );
  XNOR U3070 ( .A(n2845), .B(n2846), .Z(n2898) );
  XOR U3071 ( .A(n2899), .B(n2898), .Z(n2838) );
  XOR U3072 ( .A(n2837), .B(n2838), .Z(n2839) );
  XOR U3073 ( .A(n2840), .B(n2839), .Z(n2834) );
  ANDN U3074 ( .B(\stack[1][7] ), .A(n3923), .Z(n2831) );
  OR U3075 ( .A(n2784), .B(n2783), .Z(n2788) );
  OR U3076 ( .A(n2786), .B(n2785), .Z(n2787) );
  NAND U3077 ( .A(n2788), .B(n2787), .Z(n2832) );
  XNOR U3078 ( .A(n2831), .B(n2832), .Z(n2833) );
  XOR U3079 ( .A(n2834), .B(n2833), .Z(n2902) );
  XNOR U3080 ( .A(n2903), .B(n2902), .Z(n2904) );
  XNOR U3081 ( .A(n2905), .B(n2904), .Z(n2827) );
  NAND U3082 ( .A(\stack[1][5] ), .B(o[15]), .Z(n2825) );
  OR U3083 ( .A(n2790), .B(n2789), .Z(n2794) );
  OR U3084 ( .A(n2792), .B(n2791), .Z(n2793) );
  NAND U3085 ( .A(n2794), .B(n2793), .Z(n2826) );
  XOR U3086 ( .A(n2825), .B(n2826), .Z(n2828) );
  XNOR U3087 ( .A(n2827), .B(n2828), .Z(n2908) );
  XNOR U3088 ( .A(n2909), .B(n2908), .Z(n2910) );
  XNOR U3089 ( .A(n2911), .B(n2910), .Z(n2821) );
  NAND U3090 ( .A(\stack[1][3] ), .B(o[17]), .Z(n2819) );
  OR U3091 ( .A(n2796), .B(n2795), .Z(n2800) );
  OR U3092 ( .A(n2798), .B(n2797), .Z(n2799) );
  NAND U3093 ( .A(n2800), .B(n2799), .Z(n2820) );
  XOR U3094 ( .A(n2819), .B(n2820), .Z(n2822) );
  XNOR U3095 ( .A(n2821), .B(n2822), .Z(n2914) );
  XOR U3096 ( .A(n2915), .B(n2914), .Z(n2916) );
  ANDN U3097 ( .B(o[19]), .A(n4195), .Z(n2813) );
  OR U3098 ( .A(n2802), .B(n2801), .Z(n2806) );
  OR U3099 ( .A(n2804), .B(n2803), .Z(n2805) );
  NAND U3100 ( .A(n2806), .B(n2805), .Z(n2814) );
  XNOR U3101 ( .A(n2813), .B(n2814), .Z(n2816) );
  XOR U3102 ( .A(n2815), .B(n2816), .Z(n2807) );
  NANDN U3103 ( .A(n2808), .B(n2807), .Z(n2810) );
  XOR U3104 ( .A(n2808), .B(n2807), .Z(n4912) );
  OR U3105 ( .A(n4912), .B(n4913), .Z(n2809) );
  AND U3106 ( .A(n2810), .B(n2809), .Z(n2812) );
  OR U3107 ( .A(n2811), .B(n2812), .Z(n2921) );
  XNOR U3108 ( .A(n2812), .B(n2811), .Z(n4874) );
  NAND U3109 ( .A(\stack[1][1] ), .B(o[20]), .Z(n3032) );
  OR U3110 ( .A(n2814), .B(n2813), .Z(n2818) );
  OR U3111 ( .A(n2816), .B(n2815), .Z(n2817) );
  NAND U3112 ( .A(n2818), .B(n2817), .Z(n3030) );
  NAND U3113 ( .A(\stack[1][3] ), .B(o[18]), .Z(n3026) );
  NANDN U3114 ( .A(n2820), .B(n2819), .Z(n2824) );
  NANDN U3115 ( .A(n2822), .B(n2821), .Z(n2823) );
  NAND U3116 ( .A(n2824), .B(n2823), .Z(n3024) );
  NAND U3117 ( .A(\stack[1][5] ), .B(o[16]), .Z(n3020) );
  NANDN U3118 ( .A(n2826), .B(n2825), .Z(n2830) );
  NANDN U3119 ( .A(n2828), .B(n2827), .Z(n2829) );
  NAND U3120 ( .A(n2830), .B(n2829), .Z(n3018) );
  ANDN U3121 ( .B(o[14]), .A(n1612), .Z(n3014) );
  OR U3122 ( .A(n2832), .B(n2831), .Z(n2836) );
  OR U3123 ( .A(n2834), .B(n2833), .Z(n2835) );
  AND U3124 ( .A(n2836), .B(n2835), .Z(n3011) );
  OR U3125 ( .A(n2838), .B(n2837), .Z(n2842) );
  NANDN U3126 ( .A(n2840), .B(n2839), .Z(n2841) );
  AND U3127 ( .A(n2842), .B(n2841), .Z(n2940) );
  ANDN U3128 ( .B(\stack[1][8] ), .A(n3923), .Z(n2941) );
  XNOR U3129 ( .A(n2940), .B(n2941), .Z(n2943) );
  NANDN U3130 ( .A(n2844), .B(n2843), .Z(n2848) );
  NANDN U3131 ( .A(n2846), .B(n2845), .Z(n2847) );
  NAND U3132 ( .A(n2848), .B(n2847), .Z(n2947) );
  AND U3133 ( .A(o[11]), .B(\stack[1][10] ), .Z(n2946) );
  XNOR U3134 ( .A(n2947), .B(n2946), .Z(n2948) );
  NAND U3135 ( .A(\stack[1][11] ), .B(o[10]), .Z(n2955) );
  NANDN U3136 ( .A(n2850), .B(n2849), .Z(n2854) );
  OR U3137 ( .A(n2852), .B(n2851), .Z(n2853) );
  NAND U3138 ( .A(n2854), .B(n2853), .Z(n2953) );
  NAND U3139 ( .A(o[8]), .B(\stack[1][13] ), .Z(n3002) );
  OR U3140 ( .A(n2856), .B(n2855), .Z(n2860) );
  OR U3141 ( .A(n2858), .B(n2857), .Z(n2859) );
  NAND U3142 ( .A(n2860), .B(n2859), .Z(n3000) );
  OR U3143 ( .A(n2862), .B(n2861), .Z(n2866) );
  NANDN U3144 ( .A(n2864), .B(n2863), .Z(n2865) );
  AND U3145 ( .A(n2866), .B(n2865), .Z(n2964) );
  ANDN U3146 ( .B(\stack[1][14] ), .A(n4111), .Z(n2965) );
  XNOR U3147 ( .A(n2964), .B(n2965), .Z(n2967) );
  OR U3148 ( .A(n2868), .B(n2867), .Z(n2872) );
  OR U3149 ( .A(n2870), .B(n2869), .Z(n2871) );
  AND U3150 ( .A(n2872), .B(n2871), .Z(n2970) );
  OR U3151 ( .A(n2874), .B(n2873), .Z(n2878) );
  OR U3152 ( .A(n2876), .B(n2875), .Z(n2877) );
  NAND U3153 ( .A(n2878), .B(n2877), .Z(n2994) );
  ANDN U3154 ( .B(\stack[1][18] ), .A(n4127), .Z(n2983) );
  XNOR U3155 ( .A(n2982), .B(n2983), .Z(n2985) );
  AND U3156 ( .A(o[1]), .B(\stack[1][20] ), .Z(n2883) );
  NAND U3157 ( .A(\stack[1][21] ), .B(o[0]), .Z(n2882) );
  XNOR U3158 ( .A(n2883), .B(n2882), .Z(n2989) );
  ANDN U3159 ( .B(\stack[1][20] ), .A(n1619), .Z(n2990) );
  XOR U3160 ( .A(n2989), .B(n2988), .Z(n2984) );
  XOR U3161 ( .A(n2985), .B(n2984), .Z(n2993) );
  XNOR U3162 ( .A(n2994), .B(n2993), .Z(n2996) );
  ANDN U3163 ( .B(\stack[1][17] ), .A(n4129), .Z(n2995) );
  XNOR U3164 ( .A(n2996), .B(n2995), .Z(n2978) );
  ANDN U3165 ( .B(\stack[1][16] ), .A(n4130), .Z(n2976) );
  OR U3166 ( .A(n2885), .B(n2884), .Z(n2889) );
  NANDN U3167 ( .A(n2887), .B(n2886), .Z(n2888) );
  NAND U3168 ( .A(n2889), .B(n2888), .Z(n2977) );
  XNOR U3169 ( .A(n2976), .B(n2977), .Z(n2979) );
  XNOR U3170 ( .A(n2978), .B(n2979), .Z(n2971) );
  XOR U3171 ( .A(n2970), .B(n2971), .Z(n2972) );
  ANDN U3172 ( .B(\stack[1][15] ), .A(n4137), .Z(n2973) );
  XOR U3173 ( .A(n2972), .B(n2973), .Z(n2966) );
  XOR U3174 ( .A(n2967), .B(n2966), .Z(n2999) );
  XNOR U3175 ( .A(n3000), .B(n2999), .Z(n3001) );
  XNOR U3176 ( .A(n3002), .B(n3001), .Z(n2960) );
  ANDN U3177 ( .B(\stack[1][12] ), .A(n3977), .Z(n2958) );
  NANDN U3178 ( .A(n2891), .B(n2890), .Z(n2895) );
  NANDN U3179 ( .A(n2893), .B(n2892), .Z(n2894) );
  NAND U3180 ( .A(n2895), .B(n2894), .Z(n2959) );
  XNOR U3181 ( .A(n2958), .B(n2959), .Z(n2961) );
  XNOR U3182 ( .A(n2960), .B(n2961), .Z(n2952) );
  XNOR U3183 ( .A(n2953), .B(n2952), .Z(n2954) );
  XNOR U3184 ( .A(n2955), .B(n2954), .Z(n2949) );
  OR U3185 ( .A(n2897), .B(n2896), .Z(n2901) );
  NANDN U3186 ( .A(n2899), .B(n2898), .Z(n2900) );
  AND U3187 ( .A(n2901), .B(n2900), .Z(n3006) );
  XNOR U3188 ( .A(n3005), .B(n3006), .Z(n3008) );
  ANDN U3189 ( .B(o[12]), .A(n1614), .Z(n3007) );
  XOR U3190 ( .A(n3008), .B(n3007), .Z(n2942) );
  XOR U3191 ( .A(n2943), .B(n2942), .Z(n3012) );
  XOR U3192 ( .A(n3011), .B(n3012), .Z(n3013) );
  XOR U3193 ( .A(n3014), .B(n3013), .Z(n2937) );
  ANDN U3194 ( .B(o[15]), .A(n1611), .Z(n2934) );
  OR U3195 ( .A(n2903), .B(n2902), .Z(n2907) );
  OR U3196 ( .A(n2905), .B(n2904), .Z(n2906) );
  NAND U3197 ( .A(n2907), .B(n2906), .Z(n2935) );
  XNOR U3198 ( .A(n2934), .B(n2935), .Z(n2936) );
  XOR U3199 ( .A(n2937), .B(n2936), .Z(n3017) );
  XNOR U3200 ( .A(n3018), .B(n3017), .Z(n3019) );
  XNOR U3201 ( .A(n3020), .B(n3019), .Z(n2930) );
  ANDN U3202 ( .B(\stack[1][4] ), .A(n3911), .Z(n2928) );
  OR U3203 ( .A(n2909), .B(n2908), .Z(n2913) );
  OR U3204 ( .A(n2911), .B(n2910), .Z(n2912) );
  NAND U3205 ( .A(n2913), .B(n2912), .Z(n2929) );
  XNOR U3206 ( .A(n2928), .B(n2929), .Z(n2931) );
  XNOR U3207 ( .A(n2930), .B(n2931), .Z(n3023) );
  XNOR U3208 ( .A(n3024), .B(n3023), .Z(n3025) );
  XOR U3209 ( .A(n3026), .B(n3025), .Z(n2925) );
  ANDN U3210 ( .B(\stack[1][2] ), .A(n4068), .Z(n2922) );
  OR U3211 ( .A(n2915), .B(n2914), .Z(n2919) );
  NANDN U3212 ( .A(n2917), .B(n2916), .Z(n2918) );
  NAND U3213 ( .A(n2919), .B(n2918), .Z(n2923) );
  XOR U3214 ( .A(n2922), .B(n2923), .Z(n2924) );
  XNOR U3215 ( .A(n2925), .B(n2924), .Z(n3029) );
  XNOR U3216 ( .A(n3030), .B(n3029), .Z(n3031) );
  XOR U3217 ( .A(n3032), .B(n3031), .Z(n4875) );
  OR U3218 ( .A(n4874), .B(n4875), .Z(n2920) );
  AND U3219 ( .A(n2921), .B(n2920), .Z(n3036) );
  NAND U3220 ( .A(\stack[1][2] ), .B(o[20]), .Z(n3156) );
  OR U3221 ( .A(n2923), .B(n2922), .Z(n2927) );
  NANDN U3222 ( .A(n2925), .B(n2924), .Z(n2926) );
  NAND U3223 ( .A(n2927), .B(n2926), .Z(n3154) );
  NAND U3224 ( .A(\stack[1][4] ), .B(o[18]), .Z(n3150) );
  OR U3225 ( .A(n2929), .B(n2928), .Z(n2933) );
  NANDN U3226 ( .A(n2931), .B(n2930), .Z(n2932) );
  NAND U3227 ( .A(n2933), .B(n2932), .Z(n3148) );
  NAND U3228 ( .A(\stack[1][6] ), .B(o[16]), .Z(n3144) );
  OR U3229 ( .A(n2935), .B(n2934), .Z(n2939) );
  OR U3230 ( .A(n2937), .B(n2936), .Z(n2938) );
  NAND U3231 ( .A(n2939), .B(n2938), .Z(n3142) );
  NAND U3232 ( .A(\stack[1][8] ), .B(o[14]), .Z(n3138) );
  OR U3233 ( .A(n2941), .B(n2940), .Z(n2945) );
  NANDN U3234 ( .A(n2943), .B(n2942), .Z(n2944) );
  NAND U3235 ( .A(n2945), .B(n2944), .Z(n3136) );
  NANDN U3236 ( .A(n2947), .B(n2946), .Z(n2951) );
  NANDN U3237 ( .A(n2949), .B(n2948), .Z(n2950) );
  AND U3238 ( .A(n2951), .B(n2950), .Z(n3129) );
  ANDN U3239 ( .B(\stack[1][11] ), .A(n4144), .Z(n5259) );
  OR U3240 ( .A(n2953), .B(n2952), .Z(n2957) );
  OR U3241 ( .A(n2955), .B(n2954), .Z(n2956) );
  NAND U3242 ( .A(n2957), .B(n2956), .Z(n3071) );
  XNOR U3243 ( .A(n5259), .B(n3071), .Z(n3073) );
  OR U3244 ( .A(n2959), .B(n2958), .Z(n2963) );
  NANDN U3245 ( .A(n2961), .B(n2960), .Z(n2962) );
  AND U3246 ( .A(n2963), .B(n2962), .Z(n3123) );
  OR U3247 ( .A(n2965), .B(n2964), .Z(n2969) );
  OR U3248 ( .A(n2967), .B(n2966), .Z(n2968) );
  NAND U3249 ( .A(n2969), .B(n2968), .Z(n3118) );
  OR U3250 ( .A(n2971), .B(n2970), .Z(n2975) );
  NANDN U3251 ( .A(n2973), .B(n2972), .Z(n2974) );
  AND U3252 ( .A(n2975), .B(n2974), .Z(n3082) );
  ANDN U3253 ( .B(\stack[1][15] ), .A(n4111), .Z(n3083) );
  XNOR U3254 ( .A(n3082), .B(n3083), .Z(n3085) );
  OR U3255 ( .A(n2977), .B(n2976), .Z(n2981) );
  OR U3256 ( .A(n2979), .B(n2978), .Z(n2980) );
  AND U3257 ( .A(n2981), .B(n2980), .Z(n3088) );
  OR U3258 ( .A(n2983), .B(n2982), .Z(n2987) );
  OR U3259 ( .A(n2985), .B(n2984), .Z(n2986) );
  NAND U3260 ( .A(n2987), .B(n2986), .Z(n3112) );
  ANDN U3261 ( .B(\stack[1][19] ), .A(n4127), .Z(n3101) );
  XNOR U3262 ( .A(n3100), .B(n3101), .Z(n3103) );
  AND U3263 ( .A(o[1]), .B(\stack[1][21] ), .Z(n2992) );
  NAND U3264 ( .A(\stack[1][22] ), .B(o[0]), .Z(n2991) );
  XNOR U3265 ( .A(n2992), .B(n2991), .Z(n3107) );
  ANDN U3266 ( .B(\stack[1][21] ), .A(n1619), .Z(n3108) );
  XOR U3267 ( .A(n3107), .B(n3106), .Z(n3102) );
  XOR U3268 ( .A(n3103), .B(n3102), .Z(n3111) );
  XNOR U3269 ( .A(n3112), .B(n3111), .Z(n3114) );
  ANDN U3270 ( .B(\stack[1][18] ), .A(n4129), .Z(n3113) );
  XNOR U3271 ( .A(n3114), .B(n3113), .Z(n3096) );
  ANDN U3272 ( .B(\stack[1][17] ), .A(n4130), .Z(n3094) );
  OR U3273 ( .A(n2994), .B(n2993), .Z(n2998) );
  NANDN U3274 ( .A(n2996), .B(n2995), .Z(n2997) );
  NAND U3275 ( .A(n2998), .B(n2997), .Z(n3095) );
  XNOR U3276 ( .A(n3094), .B(n3095), .Z(n3097) );
  XNOR U3277 ( .A(n3096), .B(n3097), .Z(n3089) );
  XOR U3278 ( .A(n3088), .B(n3089), .Z(n3090) );
  ANDN U3279 ( .B(\stack[1][16] ), .A(n4137), .Z(n3091) );
  XNOR U3280 ( .A(n3085), .B(n3084), .Z(n3117) );
  XOR U3281 ( .A(n3118), .B(n3117), .Z(n3120) );
  ANDN U3282 ( .B(\stack[1][14] ), .A(n1620), .Z(n3119) );
  XNOR U3283 ( .A(n3120), .B(n3119), .Z(n3078) );
  ANDN U3284 ( .B(\stack[1][13] ), .A(n3977), .Z(n3076) );
  OR U3285 ( .A(n3000), .B(n2999), .Z(n3004) );
  OR U3286 ( .A(n3002), .B(n3001), .Z(n3003) );
  NAND U3287 ( .A(n3004), .B(n3003), .Z(n3077) );
  XNOR U3288 ( .A(n3076), .B(n3077), .Z(n3079) );
  XNOR U3289 ( .A(n3078), .B(n3079), .Z(n3124) );
  XOR U3290 ( .A(n3123), .B(n3124), .Z(n3125) );
  ANDN U3291 ( .B(\stack[1][12] ), .A(n1621), .Z(n3126) );
  XOR U3292 ( .A(n3125), .B(n3126), .Z(n3072) );
  XOR U3293 ( .A(n3073), .B(n3072), .Z(n3130) );
  XNOR U3294 ( .A(n3129), .B(n3130), .Z(n3132) );
  AND U3295 ( .A(\stack[1][10] ), .B(o[12]), .Z(n3131) );
  XOR U3296 ( .A(n3132), .B(n3131), .Z(n3067) );
  OR U3297 ( .A(n3006), .B(n3005), .Z(n3010) );
  OR U3298 ( .A(n3008), .B(n3007), .Z(n3009) );
  AND U3299 ( .A(n3010), .B(n3009), .Z(n3066) );
  NAND U3300 ( .A(\stack[1][9] ), .B(o[13]), .Z(n3065) );
  XOR U3301 ( .A(n3066), .B(n3065), .Z(n3068) );
  XNOR U3302 ( .A(n3067), .B(n3068), .Z(n3135) );
  XNOR U3303 ( .A(n3136), .B(n3135), .Z(n3137) );
  XNOR U3304 ( .A(n3138), .B(n3137), .Z(n3061) );
  OR U3305 ( .A(n3012), .B(n3011), .Z(n3016) );
  NANDN U3306 ( .A(n3014), .B(n3013), .Z(n3015) );
  AND U3307 ( .A(n3016), .B(n3015), .Z(n3060) );
  NAND U3308 ( .A(\stack[1][7] ), .B(o[15]), .Z(n3059) );
  XOR U3309 ( .A(n3060), .B(n3059), .Z(n3062) );
  XNOR U3310 ( .A(n3061), .B(n3062), .Z(n3141) );
  XNOR U3311 ( .A(n3142), .B(n3141), .Z(n3143) );
  XNOR U3312 ( .A(n3144), .B(n3143), .Z(n3055) );
  NAND U3313 ( .A(\stack[1][5] ), .B(o[17]), .Z(n3053) );
  OR U3314 ( .A(n3018), .B(n3017), .Z(n3022) );
  OR U3315 ( .A(n3020), .B(n3019), .Z(n3021) );
  NAND U3316 ( .A(n3022), .B(n3021), .Z(n3054) );
  XOR U3317 ( .A(n3053), .B(n3054), .Z(n3056) );
  XNOR U3318 ( .A(n3055), .B(n3056), .Z(n3147) );
  XNOR U3319 ( .A(n3148), .B(n3147), .Z(n3149) );
  XNOR U3320 ( .A(n3150), .B(n3149), .Z(n3049) );
  NAND U3321 ( .A(\stack[1][3] ), .B(o[19]), .Z(n3047) );
  OR U3322 ( .A(n3024), .B(n3023), .Z(n3028) );
  OR U3323 ( .A(n3026), .B(n3025), .Z(n3027) );
  NAND U3324 ( .A(n3028), .B(n3027), .Z(n3048) );
  XOR U3325 ( .A(n3047), .B(n3048), .Z(n3050) );
  XNOR U3326 ( .A(n3049), .B(n3050), .Z(n3153) );
  XOR U3327 ( .A(n3154), .B(n3153), .Z(n3155) );
  ANDN U3328 ( .B(o[21]), .A(n4195), .Z(n3041) );
  OR U3329 ( .A(n3030), .B(n3029), .Z(n3034) );
  OR U3330 ( .A(n3032), .B(n3031), .Z(n3033) );
  NAND U3331 ( .A(n3034), .B(n3033), .Z(n3042) );
  XNOR U3332 ( .A(n3041), .B(n3042), .Z(n3044) );
  XOR U3333 ( .A(n3043), .B(n3044), .Z(n3035) );
  NANDN U3334 ( .A(n3036), .B(n3035), .Z(n3038) );
  XOR U3335 ( .A(n3036), .B(n3035), .Z(n4836) );
  OR U3336 ( .A(n4836), .B(n4837), .Z(n3037) );
  AND U3337 ( .A(n3038), .B(n3037), .Z(n3040) );
  OR U3338 ( .A(n3039), .B(n3040), .Z(n3160) );
  XNOR U3339 ( .A(n3040), .B(n3039), .Z(n4798) );
  NAND U3340 ( .A(\stack[1][1] ), .B(o[22]), .Z(n3283) );
  OR U3341 ( .A(n3042), .B(n3041), .Z(n3046) );
  OR U3342 ( .A(n3044), .B(n3043), .Z(n3045) );
  NAND U3343 ( .A(n3046), .B(n3045), .Z(n3281) );
  NAND U3344 ( .A(\stack[1][3] ), .B(o[20]), .Z(n3277) );
  NANDN U3345 ( .A(n3048), .B(n3047), .Z(n3052) );
  NANDN U3346 ( .A(n3050), .B(n3049), .Z(n3051) );
  NAND U3347 ( .A(n3052), .B(n3051), .Z(n3275) );
  NAND U3348 ( .A(\stack[1][5] ), .B(o[18]), .Z(n3271) );
  NANDN U3349 ( .A(n3054), .B(n3053), .Z(n3058) );
  NANDN U3350 ( .A(n3056), .B(n3055), .Z(n3057) );
  NAND U3351 ( .A(n3058), .B(n3057), .Z(n3269) );
  NAND U3352 ( .A(\stack[1][7] ), .B(o[16]), .Z(n3265) );
  NANDN U3353 ( .A(n3060), .B(n3059), .Z(n3064) );
  NANDN U3354 ( .A(n3062), .B(n3061), .Z(n3063) );
  NAND U3355 ( .A(n3064), .B(n3063), .Z(n3263) );
  NAND U3356 ( .A(\stack[1][9] ), .B(o[14]), .Z(n3259) );
  NANDN U3357 ( .A(n3066), .B(n3065), .Z(n3070) );
  NANDN U3358 ( .A(n3068), .B(n3067), .Z(n3069) );
  NAND U3359 ( .A(n3070), .B(n3069), .Z(n3257) );
  NAND U3360 ( .A(\stack[1][11] ), .B(o[12]), .Z(n3253) );
  OR U3361 ( .A(n3071), .B(n5259), .Z(n3075) );
  OR U3362 ( .A(n3073), .B(n3072), .Z(n3074) );
  NAND U3363 ( .A(n3075), .B(n3074), .Z(n3251) );
  NAND U3364 ( .A(o[10]), .B(\stack[1][13] ), .Z(n3247) );
  OR U3365 ( .A(n3077), .B(n3076), .Z(n3081) );
  OR U3366 ( .A(n3079), .B(n3078), .Z(n3080) );
  NAND U3367 ( .A(n3081), .B(n3080), .Z(n3245) );
  NAND U3368 ( .A(o[8]), .B(\stack[1][15] ), .Z(n3241) );
  OR U3369 ( .A(n3083), .B(n3082), .Z(n3087) );
  OR U3370 ( .A(n3085), .B(n3084), .Z(n3086) );
  NAND U3371 ( .A(n3087), .B(n3086), .Z(n3239) );
  OR U3372 ( .A(n3089), .B(n3088), .Z(n3093) );
  NANDN U3373 ( .A(n3091), .B(n3090), .Z(n3092) );
  AND U3374 ( .A(n3093), .B(n3092), .Z(n3203) );
  ANDN U3375 ( .B(\stack[1][16] ), .A(n4111), .Z(n3204) );
  XNOR U3376 ( .A(n3203), .B(n3204), .Z(n3206) );
  OR U3377 ( .A(n3095), .B(n3094), .Z(n3099) );
  OR U3378 ( .A(n3097), .B(n3096), .Z(n3098) );
  AND U3379 ( .A(n3099), .B(n3098), .Z(n3209) );
  OR U3380 ( .A(n3101), .B(n3100), .Z(n3105) );
  OR U3381 ( .A(n3103), .B(n3102), .Z(n3104) );
  NAND U3382 ( .A(n3105), .B(n3104), .Z(n3233) );
  ANDN U3383 ( .B(\stack[1][20] ), .A(n4127), .Z(n3222) );
  XNOR U3384 ( .A(n3221), .B(n3222), .Z(n3224) );
  AND U3385 ( .A(o[1]), .B(\stack[1][22] ), .Z(n3110) );
  NAND U3386 ( .A(\stack[1][23] ), .B(o[0]), .Z(n3109) );
  XNOR U3387 ( .A(n3110), .B(n3109), .Z(n3228) );
  ANDN U3388 ( .B(\stack[1][22] ), .A(n1619), .Z(n3229) );
  XOR U3389 ( .A(n3228), .B(n3227), .Z(n3223) );
  XOR U3390 ( .A(n3224), .B(n3223), .Z(n3232) );
  XNOR U3391 ( .A(n3233), .B(n3232), .Z(n3235) );
  ANDN U3392 ( .B(\stack[1][19] ), .A(n4129), .Z(n3234) );
  XNOR U3393 ( .A(n3235), .B(n3234), .Z(n3217) );
  ANDN U3394 ( .B(\stack[1][18] ), .A(n4130), .Z(n3215) );
  OR U3395 ( .A(n3112), .B(n3111), .Z(n3116) );
  NANDN U3396 ( .A(n3114), .B(n3113), .Z(n3115) );
  NAND U3397 ( .A(n3116), .B(n3115), .Z(n3216) );
  XNOR U3398 ( .A(n3215), .B(n3216), .Z(n3218) );
  XNOR U3399 ( .A(n3217), .B(n3218), .Z(n3210) );
  XOR U3400 ( .A(n3209), .B(n3210), .Z(n3211) );
  ANDN U3401 ( .B(\stack[1][17] ), .A(n4137), .Z(n3212) );
  XOR U3402 ( .A(n3211), .B(n3212), .Z(n3205) );
  XOR U3403 ( .A(n3206), .B(n3205), .Z(n3238) );
  XNOR U3404 ( .A(n3239), .B(n3238), .Z(n3240) );
  XNOR U3405 ( .A(n3241), .B(n3240), .Z(n3199) );
  NAND U3406 ( .A(\stack[1][14] ), .B(o[9]), .Z(n3197) );
  NANDN U3407 ( .A(n3118), .B(n3117), .Z(n3122) );
  NANDN U3408 ( .A(n3120), .B(n3119), .Z(n3121) );
  NAND U3409 ( .A(n3122), .B(n3121), .Z(n3198) );
  XOR U3410 ( .A(n3197), .B(n3198), .Z(n3200) );
  XNOR U3411 ( .A(n3199), .B(n3200), .Z(n3244) );
  XNOR U3412 ( .A(n3245), .B(n3244), .Z(n3246) );
  XNOR U3413 ( .A(n3247), .B(n3246), .Z(n3193) );
  OR U3414 ( .A(n3124), .B(n3123), .Z(n3128) );
  NANDN U3415 ( .A(n3126), .B(n3125), .Z(n3127) );
  AND U3416 ( .A(n3128), .B(n3127), .Z(n3192) );
  NAND U3417 ( .A(\stack[1][12] ), .B(o[11]), .Z(n3191) );
  XOR U3418 ( .A(n3192), .B(n3191), .Z(n3194) );
  XNOR U3419 ( .A(n3193), .B(n3194), .Z(n3250) );
  XNOR U3420 ( .A(n3251), .B(n3250), .Z(n3252) );
  XNOR U3421 ( .A(n3253), .B(n3252), .Z(n3187) );
  NAND U3422 ( .A(\stack[1][10] ), .B(o[13]), .Z(n3185) );
  OR U3423 ( .A(n3130), .B(n3129), .Z(n3134) );
  NANDN U3424 ( .A(n3132), .B(n3131), .Z(n3133) );
  NAND U3425 ( .A(n3134), .B(n3133), .Z(n3186) );
  XOR U3426 ( .A(n3185), .B(n3186), .Z(n3188) );
  XNOR U3427 ( .A(n3187), .B(n3188), .Z(n3256) );
  XNOR U3428 ( .A(n3257), .B(n3256), .Z(n3258) );
  XNOR U3429 ( .A(n3259), .B(n3258), .Z(n3181) );
  NAND U3430 ( .A(\stack[1][8] ), .B(o[15]), .Z(n3179) );
  OR U3431 ( .A(n3136), .B(n3135), .Z(n3140) );
  OR U3432 ( .A(n3138), .B(n3137), .Z(n3139) );
  NAND U3433 ( .A(n3140), .B(n3139), .Z(n3180) );
  XOR U3434 ( .A(n3179), .B(n3180), .Z(n3182) );
  XNOR U3435 ( .A(n3181), .B(n3182), .Z(n3262) );
  XNOR U3436 ( .A(n3263), .B(n3262), .Z(n3264) );
  XNOR U3437 ( .A(n3265), .B(n3264), .Z(n3175) );
  NAND U3438 ( .A(\stack[1][6] ), .B(o[17]), .Z(n3173) );
  OR U3439 ( .A(n3142), .B(n3141), .Z(n3146) );
  OR U3440 ( .A(n3144), .B(n3143), .Z(n3145) );
  NAND U3441 ( .A(n3146), .B(n3145), .Z(n3174) );
  XOR U3442 ( .A(n3173), .B(n3174), .Z(n3176) );
  XNOR U3443 ( .A(n3175), .B(n3176), .Z(n3268) );
  XNOR U3444 ( .A(n3269), .B(n3268), .Z(n3270) );
  XNOR U3445 ( .A(n3271), .B(n3270), .Z(n3169) );
  ANDN U3446 ( .B(\stack[1][4] ), .A(n4068), .Z(n3167) );
  OR U3447 ( .A(n3148), .B(n3147), .Z(n3152) );
  OR U3448 ( .A(n3150), .B(n3149), .Z(n3151) );
  NAND U3449 ( .A(n3152), .B(n3151), .Z(n3168) );
  XNOR U3450 ( .A(n3167), .B(n3168), .Z(n3170) );
  XNOR U3451 ( .A(n3169), .B(n3170), .Z(n3274) );
  XNOR U3452 ( .A(n3275), .B(n3274), .Z(n3276) );
  XOR U3453 ( .A(n3277), .B(n3276), .Z(n3164) );
  ANDN U3454 ( .B(\stack[1][2] ), .A(n4170), .Z(n3161) );
  OR U3455 ( .A(n3154), .B(n3153), .Z(n3158) );
  NANDN U3456 ( .A(n3156), .B(n3155), .Z(n3157) );
  NAND U3457 ( .A(n3158), .B(n3157), .Z(n3162) );
  XOR U3458 ( .A(n3161), .B(n3162), .Z(n3163) );
  XNOR U3459 ( .A(n3164), .B(n3163), .Z(n3280) );
  XNOR U3460 ( .A(n3281), .B(n3280), .Z(n3282) );
  XOR U3461 ( .A(n3283), .B(n3282), .Z(n4799) );
  OR U3462 ( .A(n4798), .B(n4799), .Z(n3159) );
  AND U3463 ( .A(n3160), .B(n3159), .Z(n3287) );
  NAND U3464 ( .A(\stack[1][2] ), .B(o[22]), .Z(n3420) );
  OR U3465 ( .A(n3162), .B(n3161), .Z(n3166) );
  NANDN U3466 ( .A(n3164), .B(n3163), .Z(n3165) );
  NAND U3467 ( .A(n3166), .B(n3165), .Z(n3418) );
  NAND U3468 ( .A(\stack[1][4] ), .B(o[20]), .Z(n3414) );
  OR U3469 ( .A(n3168), .B(n3167), .Z(n3172) );
  NANDN U3470 ( .A(n3170), .B(n3169), .Z(n3171) );
  NAND U3471 ( .A(n3172), .B(n3171), .Z(n3412) );
  NAND U3472 ( .A(\stack[1][6] ), .B(o[18]), .Z(n3408) );
  NANDN U3473 ( .A(n3174), .B(n3173), .Z(n3178) );
  NANDN U3474 ( .A(n3176), .B(n3175), .Z(n3177) );
  NAND U3475 ( .A(n3178), .B(n3177), .Z(n3406) );
  NAND U3476 ( .A(\stack[1][8] ), .B(o[16]), .Z(n3402) );
  NANDN U3477 ( .A(n3180), .B(n3179), .Z(n3184) );
  NANDN U3478 ( .A(n3182), .B(n3181), .Z(n3183) );
  NAND U3479 ( .A(n3184), .B(n3183), .Z(n3400) );
  NAND U3480 ( .A(\stack[1][10] ), .B(o[14]), .Z(n3396) );
  NANDN U3481 ( .A(n3186), .B(n3185), .Z(n3190) );
  NANDN U3482 ( .A(n3188), .B(n3187), .Z(n3189) );
  NAND U3483 ( .A(n3190), .B(n3189), .Z(n3394) );
  NAND U3484 ( .A(\stack[1][12] ), .B(o[12]), .Z(n3390) );
  NANDN U3485 ( .A(n3192), .B(n3191), .Z(n3196) );
  NANDN U3486 ( .A(n3194), .B(n3193), .Z(n3195) );
  NAND U3487 ( .A(n3196), .B(n3195), .Z(n3388) );
  NAND U3488 ( .A(o[10]), .B(\stack[1][14] ), .Z(n3384) );
  NANDN U3489 ( .A(n3198), .B(n3197), .Z(n3202) );
  NANDN U3490 ( .A(n3200), .B(n3199), .Z(n3201) );
  NAND U3491 ( .A(n3202), .B(n3201), .Z(n3382) );
  NAND U3492 ( .A(o[8]), .B(\stack[1][16] ), .Z(n3378) );
  OR U3493 ( .A(n3204), .B(n3203), .Z(n3208) );
  OR U3494 ( .A(n3206), .B(n3205), .Z(n3207) );
  NAND U3495 ( .A(n3208), .B(n3207), .Z(n3376) );
  OR U3496 ( .A(n3210), .B(n3209), .Z(n3214) );
  NANDN U3497 ( .A(n3212), .B(n3211), .Z(n3213) );
  AND U3498 ( .A(n3214), .B(n3213), .Z(n3340) );
  ANDN U3499 ( .B(\stack[1][17] ), .A(n4111), .Z(n3341) );
  XNOR U3500 ( .A(n3340), .B(n3341), .Z(n3343) );
  OR U3501 ( .A(n3216), .B(n3215), .Z(n3220) );
  OR U3502 ( .A(n3218), .B(n3217), .Z(n3219) );
  AND U3503 ( .A(n3220), .B(n3219), .Z(n3346) );
  OR U3504 ( .A(n3222), .B(n3221), .Z(n3226) );
  OR U3505 ( .A(n3224), .B(n3223), .Z(n3225) );
  NAND U3506 ( .A(n3226), .B(n3225), .Z(n3370) );
  ANDN U3507 ( .B(\stack[1][21] ), .A(n4127), .Z(n3359) );
  XNOR U3508 ( .A(n3358), .B(n3359), .Z(n3361) );
  AND U3509 ( .A(o[1]), .B(\stack[1][23] ), .Z(n3231) );
  NAND U3510 ( .A(\stack[1][24] ), .B(o[0]), .Z(n3230) );
  XNOR U3511 ( .A(n3231), .B(n3230), .Z(n3365) );
  ANDN U3512 ( .B(\stack[1][23] ), .A(n1619), .Z(n3366) );
  XOR U3513 ( .A(n3365), .B(n3364), .Z(n3360) );
  XOR U3514 ( .A(n3361), .B(n3360), .Z(n3369) );
  XNOR U3515 ( .A(n3370), .B(n3369), .Z(n3372) );
  ANDN U3516 ( .B(\stack[1][20] ), .A(n4129), .Z(n3371) );
  XNOR U3517 ( .A(n3372), .B(n3371), .Z(n3354) );
  ANDN U3518 ( .B(\stack[1][19] ), .A(n4130), .Z(n3352) );
  OR U3519 ( .A(n3233), .B(n3232), .Z(n3237) );
  NANDN U3520 ( .A(n3235), .B(n3234), .Z(n3236) );
  NAND U3521 ( .A(n3237), .B(n3236), .Z(n3353) );
  XNOR U3522 ( .A(n3352), .B(n3353), .Z(n3355) );
  XNOR U3523 ( .A(n3354), .B(n3355), .Z(n3347) );
  XOR U3524 ( .A(n3346), .B(n3347), .Z(n3348) );
  ANDN U3525 ( .B(\stack[1][18] ), .A(n4137), .Z(n3349) );
  XOR U3526 ( .A(n3348), .B(n3349), .Z(n3342) );
  XOR U3527 ( .A(n3343), .B(n3342), .Z(n3375) );
  XNOR U3528 ( .A(n3376), .B(n3375), .Z(n3377) );
  XNOR U3529 ( .A(n3378), .B(n3377), .Z(n3336) );
  NAND U3530 ( .A(\stack[1][15] ), .B(o[9]), .Z(n3334) );
  OR U3531 ( .A(n3239), .B(n3238), .Z(n3243) );
  OR U3532 ( .A(n3241), .B(n3240), .Z(n3242) );
  NAND U3533 ( .A(n3243), .B(n3242), .Z(n3335) );
  XOR U3534 ( .A(n3334), .B(n3335), .Z(n3337) );
  XNOR U3535 ( .A(n3336), .B(n3337), .Z(n3381) );
  XNOR U3536 ( .A(n3382), .B(n3381), .Z(n3383) );
  XNOR U3537 ( .A(n3384), .B(n3383), .Z(n3330) );
  NAND U3538 ( .A(\stack[1][13] ), .B(o[11]), .Z(n3328) );
  OR U3539 ( .A(n3245), .B(n3244), .Z(n3249) );
  OR U3540 ( .A(n3247), .B(n3246), .Z(n3248) );
  NAND U3541 ( .A(n3249), .B(n3248), .Z(n3329) );
  XOR U3542 ( .A(n3328), .B(n3329), .Z(n3331) );
  XNOR U3543 ( .A(n3330), .B(n3331), .Z(n3387) );
  XNOR U3544 ( .A(n3388), .B(n3387), .Z(n3389) );
  XNOR U3545 ( .A(n3390), .B(n3389), .Z(n3324) );
  NAND U3546 ( .A(\stack[1][11] ), .B(o[13]), .Z(n3322) );
  OR U3547 ( .A(n3251), .B(n3250), .Z(n3255) );
  OR U3548 ( .A(n3253), .B(n3252), .Z(n3254) );
  NAND U3549 ( .A(n3255), .B(n3254), .Z(n3323) );
  XOR U3550 ( .A(n3322), .B(n3323), .Z(n3325) );
  XNOR U3551 ( .A(n3324), .B(n3325), .Z(n3393) );
  XNOR U3552 ( .A(n3394), .B(n3393), .Z(n3395) );
  XNOR U3553 ( .A(n3396), .B(n3395), .Z(n3318) );
  NAND U3554 ( .A(\stack[1][9] ), .B(o[15]), .Z(n3316) );
  OR U3555 ( .A(n3257), .B(n3256), .Z(n3261) );
  OR U3556 ( .A(n3259), .B(n3258), .Z(n3260) );
  NAND U3557 ( .A(n3261), .B(n3260), .Z(n3317) );
  XOR U3558 ( .A(n3316), .B(n3317), .Z(n3319) );
  XNOR U3559 ( .A(n3318), .B(n3319), .Z(n3399) );
  XNOR U3560 ( .A(n3400), .B(n3399), .Z(n3401) );
  XNOR U3561 ( .A(n3402), .B(n3401), .Z(n3312) );
  NAND U3562 ( .A(\stack[1][7] ), .B(o[17]), .Z(n3310) );
  OR U3563 ( .A(n3263), .B(n3262), .Z(n3267) );
  OR U3564 ( .A(n3265), .B(n3264), .Z(n3266) );
  NAND U3565 ( .A(n3267), .B(n3266), .Z(n3311) );
  XOR U3566 ( .A(n3310), .B(n3311), .Z(n3313) );
  XNOR U3567 ( .A(n3312), .B(n3313), .Z(n3405) );
  XNOR U3568 ( .A(n3406), .B(n3405), .Z(n3407) );
  XNOR U3569 ( .A(n3408), .B(n3407), .Z(n3306) );
  NAND U3570 ( .A(\stack[1][5] ), .B(o[19]), .Z(n3304) );
  OR U3571 ( .A(n3269), .B(n3268), .Z(n3273) );
  OR U3572 ( .A(n3271), .B(n3270), .Z(n3272) );
  NAND U3573 ( .A(n3273), .B(n3272), .Z(n3305) );
  XOR U3574 ( .A(n3304), .B(n3305), .Z(n3307) );
  XNOR U3575 ( .A(n3306), .B(n3307), .Z(n3411) );
  XNOR U3576 ( .A(n3412), .B(n3411), .Z(n3413) );
  XNOR U3577 ( .A(n3414), .B(n3413), .Z(n3300) );
  NAND U3578 ( .A(\stack[1][3] ), .B(o[21]), .Z(n3298) );
  OR U3579 ( .A(n3275), .B(n3274), .Z(n3279) );
  OR U3580 ( .A(n3277), .B(n3276), .Z(n3278) );
  NAND U3581 ( .A(n3279), .B(n3278), .Z(n3299) );
  XOR U3582 ( .A(n3298), .B(n3299), .Z(n3301) );
  XNOR U3583 ( .A(n3300), .B(n3301), .Z(n3417) );
  XOR U3584 ( .A(n3418), .B(n3417), .Z(n3419) );
  ANDN U3585 ( .B(o[23]), .A(n4195), .Z(n3292) );
  OR U3586 ( .A(n3281), .B(n3280), .Z(n3285) );
  OR U3587 ( .A(n3283), .B(n3282), .Z(n3284) );
  NAND U3588 ( .A(n3285), .B(n3284), .Z(n3293) );
  XNOR U3589 ( .A(n3292), .B(n3293), .Z(n3295) );
  XOR U3590 ( .A(n3294), .B(n3295), .Z(n3286) );
  NANDN U3591 ( .A(n3287), .B(n3286), .Z(n3289) );
  XOR U3592 ( .A(n3287), .B(n3286), .Z(n4760) );
  OR U3593 ( .A(n4760), .B(n4761), .Z(n3288) );
  AND U3594 ( .A(n3289), .B(n3288), .Z(n3291) );
  OR U3595 ( .A(n3290), .B(n3291), .Z(n3424) );
  XNOR U3596 ( .A(n3291), .B(n3290), .Z(n4722) );
  NAND U3597 ( .A(\stack[1][1] ), .B(o[24]), .Z(n3559) );
  OR U3598 ( .A(n3293), .B(n3292), .Z(n3297) );
  OR U3599 ( .A(n3295), .B(n3294), .Z(n3296) );
  NAND U3600 ( .A(n3297), .B(n3296), .Z(n3557) );
  NAND U3601 ( .A(\stack[1][3] ), .B(o[22]), .Z(n3553) );
  NANDN U3602 ( .A(n3299), .B(n3298), .Z(n3303) );
  NANDN U3603 ( .A(n3301), .B(n3300), .Z(n3302) );
  NAND U3604 ( .A(n3303), .B(n3302), .Z(n3551) );
  NAND U3605 ( .A(\stack[1][5] ), .B(o[20]), .Z(n3547) );
  NANDN U3606 ( .A(n3305), .B(n3304), .Z(n3309) );
  NANDN U3607 ( .A(n3307), .B(n3306), .Z(n3308) );
  NAND U3608 ( .A(n3309), .B(n3308), .Z(n3545) );
  NAND U3609 ( .A(\stack[1][7] ), .B(o[18]), .Z(n3541) );
  NANDN U3610 ( .A(n3311), .B(n3310), .Z(n3315) );
  NANDN U3611 ( .A(n3313), .B(n3312), .Z(n3314) );
  NAND U3612 ( .A(n3315), .B(n3314), .Z(n3539) );
  NAND U3613 ( .A(\stack[1][9] ), .B(o[16]), .Z(n3535) );
  NANDN U3614 ( .A(n3317), .B(n3316), .Z(n3321) );
  NANDN U3615 ( .A(n3319), .B(n3318), .Z(n3320) );
  NAND U3616 ( .A(n3321), .B(n3320), .Z(n3533) );
  NAND U3617 ( .A(\stack[1][11] ), .B(o[14]), .Z(n3529) );
  NANDN U3618 ( .A(n3323), .B(n3322), .Z(n3327) );
  NANDN U3619 ( .A(n3325), .B(n3324), .Z(n3326) );
  NAND U3620 ( .A(n3327), .B(n3326), .Z(n3527) );
  NAND U3621 ( .A(\stack[1][13] ), .B(o[12]), .Z(n3523) );
  NANDN U3622 ( .A(n3329), .B(n3328), .Z(n3333) );
  NANDN U3623 ( .A(n3331), .B(n3330), .Z(n3332) );
  NAND U3624 ( .A(n3333), .B(n3332), .Z(n3521) );
  NAND U3625 ( .A(o[10]), .B(\stack[1][15] ), .Z(n3470) );
  NANDN U3626 ( .A(n3335), .B(n3334), .Z(n3339) );
  NANDN U3627 ( .A(n3337), .B(n3336), .Z(n3338) );
  NAND U3628 ( .A(n3339), .B(n3338), .Z(n3468) );
  NAND U3629 ( .A(o[8]), .B(\stack[1][17] ), .Z(n3517) );
  OR U3630 ( .A(n3341), .B(n3340), .Z(n3345) );
  OR U3631 ( .A(n3343), .B(n3342), .Z(n3344) );
  NAND U3632 ( .A(n3345), .B(n3344), .Z(n3515) );
  OR U3633 ( .A(n3347), .B(n3346), .Z(n3351) );
  NANDN U3634 ( .A(n3349), .B(n3348), .Z(n3350) );
  AND U3635 ( .A(n3351), .B(n3350), .Z(n3479) );
  ANDN U3636 ( .B(\stack[1][18] ), .A(n4111), .Z(n3480) );
  XNOR U3637 ( .A(n3479), .B(n3480), .Z(n3482) );
  OR U3638 ( .A(n3353), .B(n3352), .Z(n3357) );
  OR U3639 ( .A(n3355), .B(n3354), .Z(n3356) );
  AND U3640 ( .A(n3357), .B(n3356), .Z(n3485) );
  OR U3641 ( .A(n3359), .B(n3358), .Z(n3363) );
  OR U3642 ( .A(n3361), .B(n3360), .Z(n3362) );
  NAND U3643 ( .A(n3363), .B(n3362), .Z(n3509) );
  ANDN U3644 ( .B(\stack[1][22] ), .A(n4127), .Z(n3498) );
  XNOR U3645 ( .A(n3497), .B(n3498), .Z(n3500) );
  AND U3646 ( .A(o[1]), .B(\stack[1][24] ), .Z(n3368) );
  NAND U3647 ( .A(\stack[1][25] ), .B(o[0]), .Z(n3367) );
  XNOR U3648 ( .A(n3368), .B(n3367), .Z(n3504) );
  ANDN U3649 ( .B(\stack[1][24] ), .A(n1619), .Z(n3505) );
  XOR U3650 ( .A(n3504), .B(n3503), .Z(n3499) );
  XOR U3651 ( .A(n3500), .B(n3499), .Z(n3508) );
  XNOR U3652 ( .A(n3509), .B(n3508), .Z(n3511) );
  ANDN U3653 ( .B(\stack[1][21] ), .A(n4129), .Z(n3510) );
  XNOR U3654 ( .A(n3511), .B(n3510), .Z(n3493) );
  ANDN U3655 ( .B(\stack[1][20] ), .A(n4130), .Z(n3491) );
  OR U3656 ( .A(n3370), .B(n3369), .Z(n3374) );
  NANDN U3657 ( .A(n3372), .B(n3371), .Z(n3373) );
  NAND U3658 ( .A(n3374), .B(n3373), .Z(n3492) );
  XNOR U3659 ( .A(n3491), .B(n3492), .Z(n3494) );
  XNOR U3660 ( .A(n3493), .B(n3494), .Z(n3486) );
  XOR U3661 ( .A(n3485), .B(n3486), .Z(n3487) );
  ANDN U3662 ( .B(\stack[1][19] ), .A(n4137), .Z(n3488) );
  XOR U3663 ( .A(n3487), .B(n3488), .Z(n3481) );
  XOR U3664 ( .A(n3482), .B(n3481), .Z(n3514) );
  XNOR U3665 ( .A(n3515), .B(n3514), .Z(n3516) );
  XNOR U3666 ( .A(n3517), .B(n3516), .Z(n3475) );
  NAND U3667 ( .A(\stack[1][16] ), .B(o[9]), .Z(n3473) );
  OR U3668 ( .A(n3376), .B(n3375), .Z(n3380) );
  OR U3669 ( .A(n3378), .B(n3377), .Z(n3379) );
  NAND U3670 ( .A(n3380), .B(n3379), .Z(n3474) );
  XOR U3671 ( .A(n3473), .B(n3474), .Z(n3476) );
  XNOR U3672 ( .A(n3475), .B(n3476), .Z(n3467) );
  XNOR U3673 ( .A(n3468), .B(n3467), .Z(n3469) );
  XNOR U3674 ( .A(n3470), .B(n3469), .Z(n3463) );
  NAND U3675 ( .A(\stack[1][14] ), .B(o[11]), .Z(n3461) );
  OR U3676 ( .A(n3382), .B(n3381), .Z(n3386) );
  OR U3677 ( .A(n3384), .B(n3383), .Z(n3385) );
  NAND U3678 ( .A(n3386), .B(n3385), .Z(n3462) );
  XOR U3679 ( .A(n3461), .B(n3462), .Z(n3464) );
  XNOR U3680 ( .A(n3463), .B(n3464), .Z(n3520) );
  XNOR U3681 ( .A(n3521), .B(n3520), .Z(n3522) );
  XNOR U3682 ( .A(n3523), .B(n3522), .Z(n3457) );
  NAND U3683 ( .A(\stack[1][12] ), .B(o[13]), .Z(n3455) );
  OR U3684 ( .A(n3388), .B(n3387), .Z(n3392) );
  OR U3685 ( .A(n3390), .B(n3389), .Z(n3391) );
  NAND U3686 ( .A(n3392), .B(n3391), .Z(n3456) );
  XOR U3687 ( .A(n3455), .B(n3456), .Z(n3458) );
  XNOR U3688 ( .A(n3457), .B(n3458), .Z(n3526) );
  XNOR U3689 ( .A(n3527), .B(n3526), .Z(n3528) );
  XNOR U3690 ( .A(n3529), .B(n3528), .Z(n3451) );
  NAND U3691 ( .A(\stack[1][10] ), .B(o[15]), .Z(n3449) );
  OR U3692 ( .A(n3394), .B(n3393), .Z(n3398) );
  OR U3693 ( .A(n3396), .B(n3395), .Z(n3397) );
  NAND U3694 ( .A(n3398), .B(n3397), .Z(n3450) );
  XOR U3695 ( .A(n3449), .B(n3450), .Z(n3452) );
  XNOR U3696 ( .A(n3451), .B(n3452), .Z(n3532) );
  XNOR U3697 ( .A(n3533), .B(n3532), .Z(n3534) );
  XNOR U3698 ( .A(n3535), .B(n3534), .Z(n3445) );
  NAND U3699 ( .A(\stack[1][8] ), .B(o[17]), .Z(n3443) );
  OR U3700 ( .A(n3400), .B(n3399), .Z(n3404) );
  OR U3701 ( .A(n3402), .B(n3401), .Z(n3403) );
  NAND U3702 ( .A(n3404), .B(n3403), .Z(n3444) );
  XOR U3703 ( .A(n3443), .B(n3444), .Z(n3446) );
  XNOR U3704 ( .A(n3445), .B(n3446), .Z(n3538) );
  XNOR U3705 ( .A(n3539), .B(n3538), .Z(n3540) );
  XNOR U3706 ( .A(n3541), .B(n3540), .Z(n3439) );
  NAND U3707 ( .A(\stack[1][6] ), .B(o[19]), .Z(n3437) );
  OR U3708 ( .A(n3406), .B(n3405), .Z(n3410) );
  OR U3709 ( .A(n3408), .B(n3407), .Z(n3409) );
  NAND U3710 ( .A(n3410), .B(n3409), .Z(n3438) );
  XOR U3711 ( .A(n3437), .B(n3438), .Z(n3440) );
  XNOR U3712 ( .A(n3439), .B(n3440), .Z(n3544) );
  XNOR U3713 ( .A(n3545), .B(n3544), .Z(n3546) );
  XNOR U3714 ( .A(n3547), .B(n3546), .Z(n3433) );
  ANDN U3715 ( .B(\stack[1][4] ), .A(n4170), .Z(n3431) );
  OR U3716 ( .A(n3412), .B(n3411), .Z(n3416) );
  OR U3717 ( .A(n3414), .B(n3413), .Z(n3415) );
  NAND U3718 ( .A(n3416), .B(n3415), .Z(n3432) );
  XNOR U3719 ( .A(n3431), .B(n3432), .Z(n3434) );
  XNOR U3720 ( .A(n3433), .B(n3434), .Z(n3550) );
  XNOR U3721 ( .A(n3551), .B(n3550), .Z(n3552) );
  XOR U3722 ( .A(n3553), .B(n3552), .Z(n3428) );
  ANDN U3723 ( .B(\stack[1][2] ), .A(n3699), .Z(n3425) );
  OR U3724 ( .A(n3418), .B(n3417), .Z(n3422) );
  NANDN U3725 ( .A(n3420), .B(n3419), .Z(n3421) );
  NAND U3726 ( .A(n3422), .B(n3421), .Z(n3426) );
  XOR U3727 ( .A(n3425), .B(n3426), .Z(n3427) );
  XNOR U3728 ( .A(n3428), .B(n3427), .Z(n3556) );
  XNOR U3729 ( .A(n3557), .B(n3556), .Z(n3558) );
  XOR U3730 ( .A(n3559), .B(n3558), .Z(n4723) );
  OR U3731 ( .A(n4722), .B(n4723), .Z(n3423) );
  AND U3732 ( .A(n3424), .B(n3423), .Z(n3563) );
  NAND U3733 ( .A(\stack[1][2] ), .B(o[24]), .Z(n3709) );
  OR U3734 ( .A(n3426), .B(n3425), .Z(n3430) );
  NANDN U3735 ( .A(n3428), .B(n3427), .Z(n3429) );
  NAND U3736 ( .A(n3430), .B(n3429), .Z(n3707) );
  NAND U3737 ( .A(\stack[1][4] ), .B(o[22]), .Z(n3703) );
  OR U3738 ( .A(n3432), .B(n3431), .Z(n3436) );
  NANDN U3739 ( .A(n3434), .B(n3433), .Z(n3435) );
  NAND U3740 ( .A(n3436), .B(n3435), .Z(n3701) );
  NAND U3741 ( .A(\stack[1][6] ), .B(o[20]), .Z(n3696) );
  NANDN U3742 ( .A(n3438), .B(n3437), .Z(n3442) );
  NANDN U3743 ( .A(n3440), .B(n3439), .Z(n3441) );
  NAND U3744 ( .A(n3442), .B(n3441), .Z(n3694) );
  NAND U3745 ( .A(\stack[1][8] ), .B(o[18]), .Z(n3690) );
  NANDN U3746 ( .A(n3444), .B(n3443), .Z(n3448) );
  NANDN U3747 ( .A(n3446), .B(n3445), .Z(n3447) );
  NAND U3748 ( .A(n3448), .B(n3447), .Z(n3688) );
  NAND U3749 ( .A(\stack[1][10] ), .B(o[16]), .Z(n3684) );
  NANDN U3750 ( .A(n3450), .B(n3449), .Z(n3454) );
  NANDN U3751 ( .A(n3452), .B(n3451), .Z(n3453) );
  NAND U3752 ( .A(n3454), .B(n3453), .Z(n3682) );
  NAND U3753 ( .A(\stack[1][12] ), .B(o[14]), .Z(n3678) );
  NANDN U3754 ( .A(n3456), .B(n3455), .Z(n3460) );
  NANDN U3755 ( .A(n3458), .B(n3457), .Z(n3459) );
  NAND U3756 ( .A(n3460), .B(n3459), .Z(n3676) );
  ANDN U3757 ( .B(\stack[1][14] ), .A(n3990), .Z(n3613) );
  NANDN U3758 ( .A(n3462), .B(n3461), .Z(n3466) );
  NANDN U3759 ( .A(n3464), .B(n3463), .Z(n3465) );
  AND U3760 ( .A(n3466), .B(n3465), .Z(n3610) );
  ANDN U3761 ( .B(\stack[1][15] ), .A(n4144), .Z(n3669) );
  OR U3762 ( .A(n3468), .B(n3467), .Z(n3472) );
  OR U3763 ( .A(n3470), .B(n3469), .Z(n3471) );
  NAND U3764 ( .A(n3472), .B(n3471), .Z(n3670) );
  XNOR U3765 ( .A(n3669), .B(n3670), .Z(n3672) );
  NANDN U3766 ( .A(n3474), .B(n3473), .Z(n3478) );
  NANDN U3767 ( .A(n3476), .B(n3475), .Z(n3477) );
  AND U3768 ( .A(n3478), .B(n3477), .Z(n3616) );
  OR U3769 ( .A(n3480), .B(n3479), .Z(n3484) );
  OR U3770 ( .A(n3482), .B(n3481), .Z(n3483) );
  NAND U3771 ( .A(n3484), .B(n3483), .Z(n3664) );
  OR U3772 ( .A(n3486), .B(n3485), .Z(n3490) );
  NANDN U3773 ( .A(n3488), .B(n3487), .Z(n3489) );
  AND U3774 ( .A(n3490), .B(n3489), .Z(n3628) );
  ANDN U3775 ( .B(\stack[1][19] ), .A(n4111), .Z(n3629) );
  XNOR U3776 ( .A(n3628), .B(n3629), .Z(n3631) );
  OR U3777 ( .A(n3492), .B(n3491), .Z(n3496) );
  OR U3778 ( .A(n3494), .B(n3493), .Z(n3495) );
  AND U3779 ( .A(n3496), .B(n3495), .Z(n3634) );
  OR U3780 ( .A(n3498), .B(n3497), .Z(n3502) );
  OR U3781 ( .A(n3500), .B(n3499), .Z(n3501) );
  NAND U3782 ( .A(n3502), .B(n3501), .Z(n3658) );
  ANDN U3783 ( .B(\stack[1][23] ), .A(n4127), .Z(n3647) );
  XNOR U3784 ( .A(n3646), .B(n3647), .Z(n3649) );
  AND U3785 ( .A(o[1]), .B(\stack[1][25] ), .Z(n3507) );
  NAND U3786 ( .A(\stack[1][26] ), .B(o[0]), .Z(n3506) );
  XNOR U3787 ( .A(n3507), .B(n3506), .Z(n3653) );
  ANDN U3788 ( .B(\stack[1][25] ), .A(n1619), .Z(n3654) );
  XOR U3789 ( .A(n3653), .B(n3652), .Z(n3648) );
  XOR U3790 ( .A(n3649), .B(n3648), .Z(n3657) );
  XNOR U3791 ( .A(n3658), .B(n3657), .Z(n3660) );
  ANDN U3792 ( .B(\stack[1][22] ), .A(n4129), .Z(n3659) );
  XNOR U3793 ( .A(n3660), .B(n3659), .Z(n3642) );
  ANDN U3794 ( .B(\stack[1][21] ), .A(n4130), .Z(n3640) );
  OR U3795 ( .A(n3509), .B(n3508), .Z(n3513) );
  NANDN U3796 ( .A(n3511), .B(n3510), .Z(n3512) );
  NAND U3797 ( .A(n3513), .B(n3512), .Z(n3641) );
  XNOR U3798 ( .A(n3640), .B(n3641), .Z(n3643) );
  XNOR U3799 ( .A(n3642), .B(n3643), .Z(n3635) );
  XOR U3800 ( .A(n3634), .B(n3635), .Z(n3636) );
  ANDN U3801 ( .B(\stack[1][20] ), .A(n4137), .Z(n3637) );
  XNOR U3802 ( .A(n3631), .B(n3630), .Z(n3663) );
  XOR U3803 ( .A(n3664), .B(n3663), .Z(n3666) );
  ANDN U3804 ( .B(\stack[1][18] ), .A(n1620), .Z(n3665) );
  XNOR U3805 ( .A(n3666), .B(n3665), .Z(n3624) );
  ANDN U3806 ( .B(\stack[1][17] ), .A(n3977), .Z(n3622) );
  OR U3807 ( .A(n3515), .B(n3514), .Z(n3519) );
  OR U3808 ( .A(n3517), .B(n3516), .Z(n3518) );
  NAND U3809 ( .A(n3519), .B(n3518), .Z(n3623) );
  XNOR U3810 ( .A(n3622), .B(n3623), .Z(n3625) );
  XNOR U3811 ( .A(n3624), .B(n3625), .Z(n3617) );
  XOR U3812 ( .A(n3616), .B(n3617), .Z(n3618) );
  ANDN U3813 ( .B(\stack[1][16] ), .A(n1621), .Z(n3619) );
  XNOR U3814 ( .A(n3672), .B(n3671), .Z(n3611) );
  XOR U3815 ( .A(n3610), .B(n3611), .Z(n3612) );
  XOR U3816 ( .A(n3613), .B(n3612), .Z(n3607) );
  ANDN U3817 ( .B(\stack[1][13] ), .A(n3923), .Z(n3604) );
  OR U3818 ( .A(n3521), .B(n3520), .Z(n3525) );
  OR U3819 ( .A(n3523), .B(n3522), .Z(n3524) );
  NAND U3820 ( .A(n3525), .B(n3524), .Z(n3605) );
  XNOR U3821 ( .A(n3604), .B(n3605), .Z(n3606) );
  XOR U3822 ( .A(n3607), .B(n3606), .Z(n3675) );
  XNOR U3823 ( .A(n3676), .B(n3675), .Z(n3677) );
  XNOR U3824 ( .A(n3678), .B(n3677), .Z(n3600) );
  NAND U3825 ( .A(\stack[1][11] ), .B(o[15]), .Z(n3598) );
  OR U3826 ( .A(n3527), .B(n3526), .Z(n3531) );
  OR U3827 ( .A(n3529), .B(n3528), .Z(n3530) );
  NAND U3828 ( .A(n3531), .B(n3530), .Z(n3599) );
  XOR U3829 ( .A(n3598), .B(n3599), .Z(n3601) );
  XNOR U3830 ( .A(n3600), .B(n3601), .Z(n3681) );
  XNOR U3831 ( .A(n3682), .B(n3681), .Z(n3683) );
  XNOR U3832 ( .A(n3684), .B(n3683), .Z(n3594) );
  NAND U3833 ( .A(\stack[1][9] ), .B(o[17]), .Z(n3592) );
  OR U3834 ( .A(n3533), .B(n3532), .Z(n3537) );
  OR U3835 ( .A(n3535), .B(n3534), .Z(n3536) );
  NAND U3836 ( .A(n3537), .B(n3536), .Z(n3593) );
  XOR U3837 ( .A(n3592), .B(n3593), .Z(n3595) );
  XNOR U3838 ( .A(n3594), .B(n3595), .Z(n3687) );
  XNOR U3839 ( .A(n3688), .B(n3687), .Z(n3689) );
  XNOR U3840 ( .A(n3690), .B(n3689), .Z(n3588) );
  NAND U3841 ( .A(\stack[1][7] ), .B(o[19]), .Z(n3586) );
  OR U3842 ( .A(n3539), .B(n3538), .Z(n3543) );
  OR U3843 ( .A(n3541), .B(n3540), .Z(n3542) );
  NAND U3844 ( .A(n3543), .B(n3542), .Z(n3587) );
  XOR U3845 ( .A(n3586), .B(n3587), .Z(n3589) );
  XNOR U3846 ( .A(n3588), .B(n3589), .Z(n3693) );
  XNOR U3847 ( .A(n3694), .B(n3693), .Z(n3695) );
  XNOR U3848 ( .A(n3696), .B(n3695), .Z(n3582) );
  NAND U3849 ( .A(\stack[1][5] ), .B(o[21]), .Z(n3580) );
  OR U3850 ( .A(n3545), .B(n3544), .Z(n3549) );
  OR U3851 ( .A(n3547), .B(n3546), .Z(n3548) );
  NAND U3852 ( .A(n3549), .B(n3548), .Z(n3581) );
  XOR U3853 ( .A(n3580), .B(n3581), .Z(n3583) );
  XNOR U3854 ( .A(n3582), .B(n3583), .Z(n3700) );
  XNOR U3855 ( .A(n3701), .B(n3700), .Z(n3702) );
  XNOR U3856 ( .A(n3703), .B(n3702), .Z(n3576) );
  NAND U3857 ( .A(\stack[1][3] ), .B(o[23]), .Z(n3574) );
  OR U3858 ( .A(n3551), .B(n3550), .Z(n3555) );
  OR U3859 ( .A(n3553), .B(n3552), .Z(n3554) );
  NAND U3860 ( .A(n3555), .B(n3554), .Z(n3575) );
  XOR U3861 ( .A(n3574), .B(n3575), .Z(n3577) );
  XNOR U3862 ( .A(n3576), .B(n3577), .Z(n3706) );
  XOR U3863 ( .A(n3707), .B(n3706), .Z(n3708) );
  ANDN U3864 ( .B(o[25]), .A(n4195), .Z(n3568) );
  OR U3865 ( .A(n3557), .B(n3556), .Z(n3561) );
  OR U3866 ( .A(n3559), .B(n3558), .Z(n3560) );
  NAND U3867 ( .A(n3561), .B(n3560), .Z(n3569) );
  XNOR U3868 ( .A(n3568), .B(n3569), .Z(n3571) );
  XOR U3869 ( .A(n3570), .B(n3571), .Z(n3562) );
  NANDN U3870 ( .A(n3563), .B(n3562), .Z(n3565) );
  XOR U3871 ( .A(n3563), .B(n3562), .Z(n4684) );
  OR U3872 ( .A(n4684), .B(n4685), .Z(n3564) );
  AND U3873 ( .A(n3565), .B(n3564), .Z(n3567) );
  OR U3874 ( .A(n3566), .B(n3567), .Z(n3713) );
  XNOR U3875 ( .A(n3567), .B(n3566), .Z(n4646) );
  NAND U3876 ( .A(\stack[1][1] ), .B(o[26]), .Z(n3860) );
  OR U3877 ( .A(n3569), .B(n3568), .Z(n3573) );
  OR U3878 ( .A(n3571), .B(n3570), .Z(n3572) );
  NAND U3879 ( .A(n3573), .B(n3572), .Z(n3858) );
  NAND U3880 ( .A(\stack[1][3] ), .B(o[24]), .Z(n3854) );
  NANDN U3881 ( .A(n3575), .B(n3574), .Z(n3579) );
  NANDN U3882 ( .A(n3577), .B(n3576), .Z(n3578) );
  NAND U3883 ( .A(n3579), .B(n3578), .Z(n3852) );
  NAND U3884 ( .A(\stack[1][5] ), .B(o[22]), .Z(n3848) );
  NANDN U3885 ( .A(n3581), .B(n3580), .Z(n3585) );
  NANDN U3886 ( .A(n3583), .B(n3582), .Z(n3584) );
  NAND U3887 ( .A(n3585), .B(n3584), .Z(n3846) );
  NAND U3888 ( .A(\stack[1][7] ), .B(o[20]), .Z(n3842) );
  NANDN U3889 ( .A(n3587), .B(n3586), .Z(n3591) );
  NANDN U3890 ( .A(n3589), .B(n3588), .Z(n3590) );
  NAND U3891 ( .A(n3591), .B(n3590), .Z(n3840) );
  NAND U3892 ( .A(\stack[1][9] ), .B(o[18]), .Z(n3836) );
  NANDN U3893 ( .A(n3593), .B(n3592), .Z(n3597) );
  NANDN U3894 ( .A(n3595), .B(n3594), .Z(n3596) );
  NAND U3895 ( .A(n3597), .B(n3596), .Z(n3834) );
  NAND U3896 ( .A(\stack[1][11] ), .B(o[16]), .Z(n3830) );
  NANDN U3897 ( .A(n3599), .B(n3598), .Z(n3603) );
  NANDN U3898 ( .A(n3601), .B(n3600), .Z(n3602) );
  NAND U3899 ( .A(n3603), .B(n3602), .Z(n3828) );
  ANDN U3900 ( .B(o[14]), .A(n3997), .Z(n3753) );
  OR U3901 ( .A(n3605), .B(n3604), .Z(n3609) );
  OR U3902 ( .A(n3607), .B(n3606), .Z(n3608) );
  AND U3903 ( .A(n3609), .B(n3608), .Z(n3750) );
  OR U3904 ( .A(n3611), .B(n3610), .Z(n3615) );
  NANDN U3905 ( .A(n3613), .B(n3612), .Z(n3614) );
  AND U3906 ( .A(n3615), .B(n3614), .Z(n3821) );
  ANDN U3907 ( .B(\stack[1][14] ), .A(n3923), .Z(n3822) );
  XNOR U3908 ( .A(n3821), .B(n3822), .Z(n3824) );
  OR U3909 ( .A(n3617), .B(n3616), .Z(n3621) );
  NANDN U3910 ( .A(n3619), .B(n3618), .Z(n3620) );
  NAND U3911 ( .A(n3621), .B(n3620), .Z(n3763) );
  AND U3912 ( .A(o[11]), .B(\stack[1][16] ), .Z(n3762) );
  XNOR U3913 ( .A(n3763), .B(n3762), .Z(n3764) );
  NAND U3914 ( .A(o[10]), .B(\stack[1][17] ), .Z(n3771) );
  OR U3915 ( .A(n3623), .B(n3622), .Z(n3627) );
  OR U3916 ( .A(n3625), .B(n3624), .Z(n3626) );
  NAND U3917 ( .A(n3627), .B(n3626), .Z(n3769) );
  NAND U3918 ( .A(o[8]), .B(\stack[1][19] ), .Z(n3818) );
  OR U3919 ( .A(n3629), .B(n3628), .Z(n3633) );
  OR U3920 ( .A(n3631), .B(n3630), .Z(n3632) );
  NAND U3921 ( .A(n3633), .B(n3632), .Z(n3816) );
  OR U3922 ( .A(n3635), .B(n3634), .Z(n3639) );
  NANDN U3923 ( .A(n3637), .B(n3636), .Z(n3638) );
  AND U3924 ( .A(n3639), .B(n3638), .Z(n3780) );
  ANDN U3925 ( .B(\stack[1][20] ), .A(n4111), .Z(n3781) );
  XNOR U3926 ( .A(n3780), .B(n3781), .Z(n3783) );
  OR U3927 ( .A(n3641), .B(n3640), .Z(n3645) );
  OR U3928 ( .A(n3643), .B(n3642), .Z(n3644) );
  AND U3929 ( .A(n3645), .B(n3644), .Z(n3786) );
  OR U3930 ( .A(n3647), .B(n3646), .Z(n3651) );
  OR U3931 ( .A(n3649), .B(n3648), .Z(n3650) );
  NAND U3932 ( .A(n3651), .B(n3650), .Z(n3810) );
  ANDN U3933 ( .B(\stack[1][24] ), .A(n4127), .Z(n3799) );
  XNOR U3934 ( .A(n3798), .B(n3799), .Z(n3801) );
  AND U3935 ( .A(o[1]), .B(\stack[1][26] ), .Z(n3656) );
  NAND U3936 ( .A(\stack[1][27] ), .B(o[0]), .Z(n3655) );
  XNOR U3937 ( .A(n3656), .B(n3655), .Z(n3805) );
  ANDN U3938 ( .B(\stack[1][26] ), .A(n1619), .Z(n3806) );
  XOR U3939 ( .A(n3805), .B(n3804), .Z(n3800) );
  XOR U3940 ( .A(n3801), .B(n3800), .Z(n3809) );
  XNOR U3941 ( .A(n3810), .B(n3809), .Z(n3812) );
  ANDN U3942 ( .B(\stack[1][23] ), .A(n4129), .Z(n3811) );
  XNOR U3943 ( .A(n3812), .B(n3811), .Z(n3794) );
  ANDN U3944 ( .B(\stack[1][22] ), .A(n4130), .Z(n3792) );
  OR U3945 ( .A(n3658), .B(n3657), .Z(n3662) );
  NANDN U3946 ( .A(n3660), .B(n3659), .Z(n3661) );
  NAND U3947 ( .A(n3662), .B(n3661), .Z(n3793) );
  XNOR U3948 ( .A(n3792), .B(n3793), .Z(n3795) );
  XNOR U3949 ( .A(n3794), .B(n3795), .Z(n3787) );
  XOR U3950 ( .A(n3786), .B(n3787), .Z(n3788) );
  ANDN U3951 ( .B(\stack[1][21] ), .A(n4137), .Z(n3789) );
  XOR U3952 ( .A(n3788), .B(n3789), .Z(n3782) );
  XOR U3953 ( .A(n3783), .B(n3782), .Z(n3815) );
  XNOR U3954 ( .A(n3816), .B(n3815), .Z(n3817) );
  XNOR U3955 ( .A(n3818), .B(n3817), .Z(n3776) );
  ANDN U3956 ( .B(\stack[1][18] ), .A(n3977), .Z(n3774) );
  NANDN U3957 ( .A(n3664), .B(n3663), .Z(n3668) );
  NANDN U3958 ( .A(n3666), .B(n3665), .Z(n3667) );
  NAND U3959 ( .A(n3668), .B(n3667), .Z(n3775) );
  XNOR U3960 ( .A(n3774), .B(n3775), .Z(n3777) );
  XNOR U3961 ( .A(n3776), .B(n3777), .Z(n3768) );
  XNOR U3962 ( .A(n3769), .B(n3768), .Z(n3770) );
  XNOR U3963 ( .A(n3771), .B(n3770), .Z(n3765) );
  OR U3964 ( .A(n3670), .B(n3669), .Z(n3674) );
  OR U3965 ( .A(n3672), .B(n3671), .Z(n3673) );
  AND U3966 ( .A(n3674), .B(n3673), .Z(n3757) );
  XNOR U3967 ( .A(n3756), .B(n3757), .Z(n3759) );
  ANDN U3968 ( .B(\stack[1][15] ), .A(n3990), .Z(n3758) );
  XOR U3969 ( .A(n3759), .B(n3758), .Z(n3823) );
  XOR U3970 ( .A(n3824), .B(n3823), .Z(n3751) );
  XOR U3971 ( .A(n3750), .B(n3751), .Z(n3752) );
  XOR U3972 ( .A(n3753), .B(n3752), .Z(n3747) );
  ANDN U3973 ( .B(o[15]), .A(n1617), .Z(n3744) );
  OR U3974 ( .A(n3676), .B(n3675), .Z(n3680) );
  OR U3975 ( .A(n3678), .B(n3677), .Z(n3679) );
  NAND U3976 ( .A(n3680), .B(n3679), .Z(n3745) );
  XNOR U3977 ( .A(n3744), .B(n3745), .Z(n3746) );
  XOR U3978 ( .A(n3747), .B(n3746), .Z(n3827) );
  XNOR U3979 ( .A(n3828), .B(n3827), .Z(n3829) );
  XNOR U3980 ( .A(n3830), .B(n3829), .Z(n3740) );
  NAND U3981 ( .A(\stack[1][10] ), .B(o[17]), .Z(n3738) );
  OR U3982 ( .A(n3682), .B(n3681), .Z(n3686) );
  OR U3983 ( .A(n3684), .B(n3683), .Z(n3685) );
  NAND U3984 ( .A(n3686), .B(n3685), .Z(n3739) );
  XOR U3985 ( .A(n3738), .B(n3739), .Z(n3741) );
  XNOR U3986 ( .A(n3740), .B(n3741), .Z(n3833) );
  XNOR U3987 ( .A(n3834), .B(n3833), .Z(n3835) );
  XNOR U3988 ( .A(n3836), .B(n3835), .Z(n3734) );
  NAND U3989 ( .A(\stack[1][8] ), .B(o[19]), .Z(n3732) );
  OR U3990 ( .A(n3688), .B(n3687), .Z(n3692) );
  OR U3991 ( .A(n3690), .B(n3689), .Z(n3691) );
  NAND U3992 ( .A(n3692), .B(n3691), .Z(n3733) );
  XOR U3993 ( .A(n3732), .B(n3733), .Z(n3735) );
  XNOR U3994 ( .A(n3734), .B(n3735), .Z(n3839) );
  XNOR U3995 ( .A(n3840), .B(n3839), .Z(n3841) );
  XNOR U3996 ( .A(n3842), .B(n3841), .Z(n3728) );
  NAND U3997 ( .A(\stack[1][6] ), .B(o[21]), .Z(n3726) );
  OR U3998 ( .A(n3694), .B(n3693), .Z(n3698) );
  OR U3999 ( .A(n3696), .B(n3695), .Z(n3697) );
  NAND U4000 ( .A(n3698), .B(n3697), .Z(n3727) );
  XOR U4001 ( .A(n3726), .B(n3727), .Z(n3729) );
  XNOR U4002 ( .A(n3728), .B(n3729), .Z(n3845) );
  XNOR U4003 ( .A(n3846), .B(n3845), .Z(n3847) );
  XNOR U4004 ( .A(n3848), .B(n3847), .Z(n3722) );
  ANDN U4005 ( .B(\stack[1][4] ), .A(n3699), .Z(n3720) );
  OR U4006 ( .A(n3701), .B(n3700), .Z(n3705) );
  OR U4007 ( .A(n3703), .B(n3702), .Z(n3704) );
  NAND U4008 ( .A(n3705), .B(n3704), .Z(n3721) );
  XNOR U4009 ( .A(n3720), .B(n3721), .Z(n3723) );
  XNOR U4010 ( .A(n3722), .B(n3723), .Z(n3851) );
  XNOR U4011 ( .A(n3852), .B(n3851), .Z(n3853) );
  XOR U4012 ( .A(n3854), .B(n3853), .Z(n3717) );
  ANDN U4013 ( .B(\stack[1][2] ), .A(n4016), .Z(n3714) );
  OR U4014 ( .A(n3707), .B(n3706), .Z(n3711) );
  NANDN U4015 ( .A(n3709), .B(n3708), .Z(n3710) );
  NAND U4016 ( .A(n3711), .B(n3710), .Z(n3715) );
  XOR U4017 ( .A(n3714), .B(n3715), .Z(n3716) );
  XNOR U4018 ( .A(n3717), .B(n3716), .Z(n3857) );
  XNOR U4019 ( .A(n3858), .B(n3857), .Z(n3859) );
  XOR U4020 ( .A(n3860), .B(n3859), .Z(n4647) );
  OR U4021 ( .A(n4646), .B(n4647), .Z(n3712) );
  AND U4022 ( .A(n3713), .B(n3712), .Z(n3864) );
  NAND U4023 ( .A(\stack[1][2] ), .B(o[26]), .Z(n4027) );
  OR U4024 ( .A(n3715), .B(n3714), .Z(n3719) );
  NANDN U4025 ( .A(n3717), .B(n3716), .Z(n3718) );
  NAND U4026 ( .A(n3719), .B(n3718), .Z(n4025) );
  NAND U4027 ( .A(\stack[1][4] ), .B(o[24]), .Z(n4020) );
  OR U4028 ( .A(n3721), .B(n3720), .Z(n3725) );
  NANDN U4029 ( .A(n3723), .B(n3722), .Z(n3724) );
  NAND U4030 ( .A(n3725), .B(n3724), .Z(n4018) );
  NAND U4031 ( .A(\stack[1][6] ), .B(o[22]), .Z(n4013) );
  NANDN U4032 ( .A(n3727), .B(n3726), .Z(n3731) );
  NANDN U4033 ( .A(n3729), .B(n3728), .Z(n3730) );
  NAND U4034 ( .A(n3731), .B(n3730), .Z(n4011) );
  NAND U4035 ( .A(\stack[1][8] ), .B(o[20]), .Z(n4007) );
  NANDN U4036 ( .A(n3733), .B(n3732), .Z(n3737) );
  NANDN U4037 ( .A(n3735), .B(n3734), .Z(n3736) );
  NAND U4038 ( .A(n3737), .B(n3736), .Z(n4005) );
  NAND U4039 ( .A(\stack[1][10] ), .B(o[18]), .Z(n4001) );
  NANDN U4040 ( .A(n3739), .B(n3738), .Z(n3743) );
  NANDN U4041 ( .A(n3741), .B(n3740), .Z(n3742) );
  NAND U4042 ( .A(n3743), .B(n3742), .Z(n3999) );
  ANDN U4043 ( .B(o[16]), .A(n1617), .Z(n3908) );
  OR U4044 ( .A(n3745), .B(n3744), .Z(n3749) );
  OR U4045 ( .A(n3747), .B(n3746), .Z(n3748) );
  AND U4046 ( .A(n3749), .B(n3748), .Z(n3905) );
  OR U4047 ( .A(n3751), .B(n3750), .Z(n3755) );
  NANDN U4048 ( .A(n3753), .B(n3752), .Z(n3754) );
  AND U4049 ( .A(n3755), .B(n3754), .Z(n3991) );
  ANDN U4050 ( .B(o[15]), .A(n3997), .Z(n3992) );
  XNOR U4051 ( .A(n3991), .B(n3992), .Z(n3994) );
  ANDN U4052 ( .B(o[14]), .A(n1618), .Z(n5147) );
  OR U4053 ( .A(n3757), .B(n3756), .Z(n3761) );
  OR U4054 ( .A(n3759), .B(n3758), .Z(n3760) );
  NAND U4055 ( .A(n3761), .B(n3760), .Z(n3918) );
  AND U4056 ( .A(o[13]), .B(\stack[1][15] ), .Z(n3917) );
  XNOR U4057 ( .A(n3918), .B(n3917), .Z(n3920) );
  NAND U4058 ( .A(o[12]), .B(\stack[1][16] ), .Z(n3927) );
  NANDN U4059 ( .A(n3763), .B(n3762), .Z(n3767) );
  NANDN U4060 ( .A(n3765), .B(n3764), .Z(n3766) );
  AND U4061 ( .A(n3767), .B(n3766), .Z(n3924) );
  ANDN U4062 ( .B(\stack[1][17] ), .A(n4144), .Z(n3984) );
  OR U4063 ( .A(n3769), .B(n3768), .Z(n3773) );
  OR U4064 ( .A(n3771), .B(n3770), .Z(n3772) );
  NAND U4065 ( .A(n3773), .B(n3772), .Z(n3985) );
  XNOR U4066 ( .A(n3984), .B(n3985), .Z(n3987) );
  OR U4067 ( .A(n3775), .B(n3774), .Z(n3779) );
  NANDN U4068 ( .A(n3777), .B(n3776), .Z(n3778) );
  AND U4069 ( .A(n3779), .B(n3778), .Z(n3930) );
  OR U4070 ( .A(n3781), .B(n3780), .Z(n3785) );
  OR U4071 ( .A(n3783), .B(n3782), .Z(n3784) );
  NAND U4072 ( .A(n3785), .B(n3784), .Z(n3979) );
  OR U4073 ( .A(n3787), .B(n3786), .Z(n3791) );
  NANDN U4074 ( .A(n3789), .B(n3788), .Z(n3790) );
  AND U4075 ( .A(n3791), .B(n3790), .Z(n3942) );
  ANDN U4076 ( .B(\stack[1][21] ), .A(n4111), .Z(n3943) );
  XNOR U4077 ( .A(n3942), .B(n3943), .Z(n3945) );
  OR U4078 ( .A(n3793), .B(n3792), .Z(n3797) );
  OR U4079 ( .A(n3795), .B(n3794), .Z(n3796) );
  AND U4080 ( .A(n3797), .B(n3796), .Z(n3948) );
  OR U4081 ( .A(n3799), .B(n3798), .Z(n3803) );
  OR U4082 ( .A(n3801), .B(n3800), .Z(n3802) );
  NAND U4083 ( .A(n3803), .B(n3802), .Z(n3972) );
  ANDN U4084 ( .B(\stack[1][25] ), .A(n4127), .Z(n3961) );
  XNOR U4085 ( .A(n3960), .B(n3961), .Z(n3963) );
  AND U4086 ( .A(o[1]), .B(\stack[1][27] ), .Z(n3808) );
  NAND U4087 ( .A(\stack[1][28] ), .B(o[0]), .Z(n3807) );
  XNOR U4088 ( .A(n3808), .B(n3807), .Z(n3967) );
  ANDN U4089 ( .B(\stack[1][27] ), .A(n1619), .Z(n3968) );
  XOR U4090 ( .A(n3967), .B(n3966), .Z(n3962) );
  XOR U4091 ( .A(n3963), .B(n3962), .Z(n3971) );
  XNOR U4092 ( .A(n3972), .B(n3971), .Z(n3974) );
  ANDN U4093 ( .B(\stack[1][24] ), .A(n4129), .Z(n3973) );
  XNOR U4094 ( .A(n3974), .B(n3973), .Z(n3956) );
  ANDN U4095 ( .B(\stack[1][23] ), .A(n4130), .Z(n3954) );
  OR U4096 ( .A(n3810), .B(n3809), .Z(n3814) );
  NANDN U4097 ( .A(n3812), .B(n3811), .Z(n3813) );
  NAND U4098 ( .A(n3814), .B(n3813), .Z(n3955) );
  XNOR U4099 ( .A(n3954), .B(n3955), .Z(n3957) );
  XNOR U4100 ( .A(n3956), .B(n3957), .Z(n3949) );
  XOR U4101 ( .A(n3948), .B(n3949), .Z(n3950) );
  ANDN U4102 ( .B(\stack[1][22] ), .A(n4137), .Z(n3951) );
  XNOR U4103 ( .A(n3945), .B(n3944), .Z(n3978) );
  XOR U4104 ( .A(n3979), .B(n3978), .Z(n3981) );
  ANDN U4105 ( .B(\stack[1][20] ), .A(n1620), .Z(n3980) );
  XNOR U4106 ( .A(n3981), .B(n3980), .Z(n3938) );
  ANDN U4107 ( .B(\stack[1][19] ), .A(n3977), .Z(n3936) );
  OR U4108 ( .A(n3816), .B(n3815), .Z(n3820) );
  OR U4109 ( .A(n3818), .B(n3817), .Z(n3819) );
  NAND U4110 ( .A(n3820), .B(n3819), .Z(n3937) );
  XNOR U4111 ( .A(n3936), .B(n3937), .Z(n3939) );
  XNOR U4112 ( .A(n3938), .B(n3939), .Z(n3931) );
  XOR U4113 ( .A(n3930), .B(n3931), .Z(n3932) );
  ANDN U4114 ( .B(\stack[1][18] ), .A(n1621), .Z(n3933) );
  XOR U4115 ( .A(n3932), .B(n3933), .Z(n3986) );
  XOR U4116 ( .A(n3987), .B(n3986), .Z(n3925) );
  XOR U4117 ( .A(n3924), .B(n3925), .Z(n3926) );
  XNOR U4118 ( .A(n3920), .B(n3919), .Z(n3912) );
  OR U4119 ( .A(n3822), .B(n3821), .Z(n3826) );
  NANDN U4120 ( .A(n3824), .B(n3823), .Z(n3825) );
  AND U4121 ( .A(n3826), .B(n3825), .Z(n3913) );
  XOR U4122 ( .A(n3912), .B(n3913), .Z(n3914) );
  XNOR U4123 ( .A(n5147), .B(n3914), .Z(n3993) );
  XNOR U4124 ( .A(n3994), .B(n3993), .Z(n3906) );
  XOR U4125 ( .A(n3905), .B(n3906), .Z(n3907) );
  XOR U4126 ( .A(n3908), .B(n3907), .Z(n3902) );
  ANDN U4127 ( .B(\stack[1][11] ), .A(n3911), .Z(n3899) );
  OR U4128 ( .A(n3828), .B(n3827), .Z(n3832) );
  OR U4129 ( .A(n3830), .B(n3829), .Z(n3831) );
  NAND U4130 ( .A(n3832), .B(n3831), .Z(n3900) );
  XNOR U4131 ( .A(n3899), .B(n3900), .Z(n3901) );
  XOR U4132 ( .A(n3902), .B(n3901), .Z(n3998) );
  XNOR U4133 ( .A(n3999), .B(n3998), .Z(n4000) );
  XNOR U4134 ( .A(n4001), .B(n4000), .Z(n3895) );
  NAND U4135 ( .A(\stack[1][9] ), .B(o[19]), .Z(n3893) );
  OR U4136 ( .A(n3834), .B(n3833), .Z(n3838) );
  OR U4137 ( .A(n3836), .B(n3835), .Z(n3837) );
  NAND U4138 ( .A(n3838), .B(n3837), .Z(n3894) );
  XOR U4139 ( .A(n3893), .B(n3894), .Z(n3896) );
  XNOR U4140 ( .A(n3895), .B(n3896), .Z(n4004) );
  XNOR U4141 ( .A(n4005), .B(n4004), .Z(n4006) );
  XNOR U4142 ( .A(n4007), .B(n4006), .Z(n3889) );
  NAND U4143 ( .A(\stack[1][7] ), .B(o[21]), .Z(n3887) );
  OR U4144 ( .A(n3840), .B(n3839), .Z(n3844) );
  OR U4145 ( .A(n3842), .B(n3841), .Z(n3843) );
  NAND U4146 ( .A(n3844), .B(n3843), .Z(n3888) );
  XOR U4147 ( .A(n3887), .B(n3888), .Z(n3890) );
  XNOR U4148 ( .A(n3889), .B(n3890), .Z(n4010) );
  XNOR U4149 ( .A(n4011), .B(n4010), .Z(n4012) );
  XNOR U4150 ( .A(n4013), .B(n4012), .Z(n3883) );
  NAND U4151 ( .A(\stack[1][5] ), .B(o[23]), .Z(n3881) );
  OR U4152 ( .A(n3846), .B(n3845), .Z(n3850) );
  OR U4153 ( .A(n3848), .B(n3847), .Z(n3849) );
  NAND U4154 ( .A(n3850), .B(n3849), .Z(n3882) );
  XOR U4155 ( .A(n3881), .B(n3882), .Z(n3884) );
  XNOR U4156 ( .A(n3883), .B(n3884), .Z(n4017) );
  XNOR U4157 ( .A(n4018), .B(n4017), .Z(n4019) );
  XNOR U4158 ( .A(n4020), .B(n4019), .Z(n3877) );
  NAND U4159 ( .A(\stack[1][3] ), .B(o[25]), .Z(n3875) );
  OR U4160 ( .A(n3852), .B(n3851), .Z(n3856) );
  OR U4161 ( .A(n3854), .B(n3853), .Z(n3855) );
  NAND U4162 ( .A(n3856), .B(n3855), .Z(n3876) );
  XOR U4163 ( .A(n3875), .B(n3876), .Z(n3878) );
  XNOR U4164 ( .A(n3877), .B(n3878), .Z(n4024) );
  XOR U4165 ( .A(n4025), .B(n4024), .Z(n4026) );
  ANDN U4166 ( .B(o[27]), .A(n4195), .Z(n3869) );
  OR U4167 ( .A(n3858), .B(n3857), .Z(n3862) );
  OR U4168 ( .A(n3860), .B(n3859), .Z(n3861) );
  NAND U4169 ( .A(n3862), .B(n3861), .Z(n3870) );
  XNOR U4170 ( .A(n3869), .B(n3870), .Z(n3872) );
  XOR U4171 ( .A(n3871), .B(n3872), .Z(n3863) );
  NANDN U4172 ( .A(n3864), .B(n3863), .Z(n3866) );
  XOR U4173 ( .A(n3864), .B(n3863), .Z(n4608) );
  OR U4174 ( .A(n4608), .B(n4609), .Z(n3865) );
  AND U4175 ( .A(n3866), .B(n3865), .Z(n3868) );
  OR U4176 ( .A(n3867), .B(n3868), .Z(n4031) );
  XNOR U4177 ( .A(n3868), .B(n3867), .Z(n4570) );
  NAND U4178 ( .A(\stack[1][1] ), .B(o[28]), .Z(n4199) );
  OR U4179 ( .A(n3870), .B(n3869), .Z(n3874) );
  OR U4180 ( .A(n3872), .B(n3871), .Z(n3873) );
  NAND U4181 ( .A(n3874), .B(n3873), .Z(n4197) );
  NAND U4182 ( .A(\stack[1][3] ), .B(o[26]), .Z(n4192) );
  NANDN U4183 ( .A(n3876), .B(n3875), .Z(n3880) );
  NANDN U4184 ( .A(n3878), .B(n3877), .Z(n3879) );
  NAND U4185 ( .A(n3880), .B(n3879), .Z(n4190) );
  NAND U4186 ( .A(\stack[1][5] ), .B(o[24]), .Z(n4186) );
  NANDN U4187 ( .A(n3882), .B(n3881), .Z(n3886) );
  NANDN U4188 ( .A(n3884), .B(n3883), .Z(n3885) );
  NAND U4189 ( .A(n3886), .B(n3885), .Z(n4184) );
  NAND U4190 ( .A(\stack[1][7] ), .B(o[22]), .Z(n4180) );
  NANDN U4191 ( .A(n3888), .B(n3887), .Z(n3892) );
  NANDN U4192 ( .A(n3890), .B(n3889), .Z(n3891) );
  NAND U4193 ( .A(n3892), .B(n3891), .Z(n4178) );
  NAND U4194 ( .A(\stack[1][9] ), .B(o[20]), .Z(n4174) );
  NANDN U4195 ( .A(n3894), .B(n3893), .Z(n3898) );
  NANDN U4196 ( .A(n3896), .B(n3895), .Z(n3897) );
  NAND U4197 ( .A(n3898), .B(n3897), .Z(n4172) );
  ANDN U4198 ( .B(o[18]), .A(n1616), .Z(n4065) );
  OR U4199 ( .A(n3900), .B(n3899), .Z(n3904) );
  OR U4200 ( .A(n3902), .B(n3901), .Z(n3903) );
  AND U4201 ( .A(n3904), .B(n3903), .Z(n4062) );
  OR U4202 ( .A(n3906), .B(n3905), .Z(n3910) );
  NANDN U4203 ( .A(n3908), .B(n3907), .Z(n3909) );
  AND U4204 ( .A(n3910), .B(n3909), .Z(n4164) );
  ANDN U4205 ( .B(\stack[1][12] ), .A(n3911), .Z(n4165) );
  XNOR U4206 ( .A(n4164), .B(n4165), .Z(n4167) );
  NANDN U4207 ( .A(n3913), .B(n3912), .Z(n3916) );
  OR U4208 ( .A(n3914), .B(n5147), .Z(n3915) );
  NAND U4209 ( .A(n3916), .B(n3915), .Z(n4076) );
  AND U4210 ( .A(o[15]), .B(\stack[1][14] ), .Z(n4075) );
  XNOR U4211 ( .A(n4076), .B(n4075), .Z(n4077) );
  NAND U4212 ( .A(\stack[1][15] ), .B(o[14]), .Z(n4161) );
  NANDN U4213 ( .A(n3918), .B(n3917), .Z(n3922) );
  NAND U4214 ( .A(n3920), .B(n3919), .Z(n3921) );
  AND U4215 ( .A(n3922), .B(n3921), .Z(n4158) );
  ANDN U4216 ( .B(\stack[1][16] ), .A(n3923), .Z(n4081) );
  OR U4217 ( .A(n3925), .B(n3924), .Z(n3929) );
  NANDN U4218 ( .A(n3927), .B(n3926), .Z(n3928) );
  NAND U4219 ( .A(n3929), .B(n3928), .Z(n4082) );
  XNOR U4220 ( .A(n4081), .B(n4082), .Z(n4084) );
  OR U4221 ( .A(n3931), .B(n3930), .Z(n3935) );
  NANDN U4222 ( .A(n3933), .B(n3932), .Z(n3934) );
  NAND U4223 ( .A(n3935), .B(n3934), .Z(n4088) );
  AND U4224 ( .A(o[11]), .B(\stack[1][18] ), .Z(n4087) );
  XNOR U4225 ( .A(n4088), .B(n4087), .Z(n4089) );
  NAND U4226 ( .A(o[10]), .B(\stack[1][19] ), .Z(n4148) );
  OR U4227 ( .A(n3937), .B(n3936), .Z(n3941) );
  OR U4228 ( .A(n3939), .B(n3938), .Z(n3940) );
  NAND U4229 ( .A(n3941), .B(n3940), .Z(n4146) );
  NAND U4230 ( .A(o[8]), .B(\stack[1][21] ), .Z(n4141) );
  OR U4231 ( .A(n3943), .B(n3942), .Z(n3947) );
  OR U4232 ( .A(n3945), .B(n3944), .Z(n3946) );
  NAND U4233 ( .A(n3947), .B(n3946), .Z(n4139) );
  OR U4234 ( .A(n3949), .B(n3948), .Z(n3953) );
  NANDN U4235 ( .A(n3951), .B(n3950), .Z(n3952) );
  AND U4236 ( .A(n3953), .B(n3952), .Z(n4099) );
  ANDN U4237 ( .B(\stack[1][22] ), .A(n4111), .Z(n4100) );
  XNOR U4238 ( .A(n4099), .B(n4100), .Z(n4102) );
  OR U4239 ( .A(n3955), .B(n3954), .Z(n3959) );
  OR U4240 ( .A(n3957), .B(n3956), .Z(n3958) );
  AND U4241 ( .A(n3959), .B(n3958), .Z(n4105) );
  OR U4242 ( .A(n3961), .B(n3960), .Z(n3965) );
  OR U4243 ( .A(n3963), .B(n3962), .Z(n3964) );
  NAND U4244 ( .A(n3965), .B(n3964), .Z(n4132) );
  ANDN U4245 ( .B(\stack[1][26] ), .A(n4127), .Z(n4119) );
  XNOR U4246 ( .A(n4118), .B(n4119), .Z(n4121) );
  AND U4247 ( .A(o[1]), .B(\stack[1][28] ), .Z(n3970) );
  NAND U4248 ( .A(o[0]), .B(\stack[1][29] ), .Z(n3969) );
  XNOR U4249 ( .A(n3970), .B(n3969), .Z(n4125) );
  ANDN U4250 ( .B(\stack[1][28] ), .A(n1619), .Z(n4126) );
  XOR U4251 ( .A(n4125), .B(n4124), .Z(n4120) );
  XOR U4252 ( .A(n4121), .B(n4120), .Z(n4131) );
  XNOR U4253 ( .A(n4132), .B(n4131), .Z(n4134) );
  ANDN U4254 ( .B(\stack[1][25] ), .A(n4129), .Z(n4133) );
  XNOR U4255 ( .A(n4134), .B(n4133), .Z(n4114) );
  ANDN U4256 ( .B(\stack[1][24] ), .A(n4130), .Z(n4112) );
  OR U4257 ( .A(n3972), .B(n3971), .Z(n3976) );
  NANDN U4258 ( .A(n3974), .B(n3973), .Z(n3975) );
  NAND U4259 ( .A(n3976), .B(n3975), .Z(n4113) );
  XNOR U4260 ( .A(n4112), .B(n4113), .Z(n4115) );
  XNOR U4261 ( .A(n4114), .B(n4115), .Z(n4106) );
  XOR U4262 ( .A(n4105), .B(n4106), .Z(n4107) );
  ANDN U4263 ( .B(\stack[1][23] ), .A(n4137), .Z(n4108) );
  XOR U4264 ( .A(n4107), .B(n4108), .Z(n4101) );
  XOR U4265 ( .A(n4102), .B(n4101), .Z(n4138) );
  XNOR U4266 ( .A(n4139), .B(n4138), .Z(n4140) );
  XNOR U4267 ( .A(n4141), .B(n4140), .Z(n4095) );
  ANDN U4268 ( .B(\stack[1][20] ), .A(n3977), .Z(n4093) );
  NANDN U4269 ( .A(n3979), .B(n3978), .Z(n3983) );
  NANDN U4270 ( .A(n3981), .B(n3980), .Z(n3982) );
  NAND U4271 ( .A(n3983), .B(n3982), .Z(n4094) );
  XNOR U4272 ( .A(n4093), .B(n4094), .Z(n4096) );
  XNOR U4273 ( .A(n4095), .B(n4096), .Z(n4145) );
  XNOR U4274 ( .A(n4146), .B(n4145), .Z(n4147) );
  XNOR U4275 ( .A(n4148), .B(n4147), .Z(n4090) );
  OR U4276 ( .A(n3985), .B(n3984), .Z(n3989) );
  OR U4277 ( .A(n3987), .B(n3986), .Z(n3988) );
  AND U4278 ( .A(n3989), .B(n3988), .Z(n4152) );
  XNOR U4279 ( .A(n4151), .B(n4152), .Z(n4154) );
  ANDN U4280 ( .B(\stack[1][17] ), .A(n3990), .Z(n4153) );
  XNOR U4281 ( .A(n4154), .B(n4153), .Z(n4083) );
  XOR U4282 ( .A(n4084), .B(n4083), .Z(n4159) );
  XOR U4283 ( .A(n4158), .B(n4159), .Z(n4160) );
  XOR U4284 ( .A(n4077), .B(n4078), .Z(n4069) );
  OR U4285 ( .A(n3992), .B(n3991), .Z(n3996) );
  OR U4286 ( .A(n3994), .B(n3993), .Z(n3995) );
  AND U4287 ( .A(n3996), .B(n3995), .Z(n4070) );
  XOR U4288 ( .A(n4069), .B(n4070), .Z(n4072) );
  ANDN U4289 ( .B(o[16]), .A(n3997), .Z(n4071) );
  XOR U4290 ( .A(n4072), .B(n4071), .Z(n4166) );
  XOR U4291 ( .A(n4167), .B(n4166), .Z(n4063) );
  XOR U4292 ( .A(n4062), .B(n4063), .Z(n4064) );
  XOR U4293 ( .A(n4065), .B(n4064), .Z(n4059) );
  ANDN U4294 ( .B(\stack[1][10] ), .A(n4068), .Z(n4056) );
  OR U4295 ( .A(n3999), .B(n3998), .Z(n4003) );
  OR U4296 ( .A(n4001), .B(n4000), .Z(n4002) );
  NAND U4297 ( .A(n4003), .B(n4002), .Z(n4057) );
  XNOR U4298 ( .A(n4056), .B(n4057), .Z(n4058) );
  XOR U4299 ( .A(n4059), .B(n4058), .Z(n4171) );
  XNOR U4300 ( .A(n4172), .B(n4171), .Z(n4173) );
  XNOR U4301 ( .A(n4174), .B(n4173), .Z(n4052) );
  NAND U4302 ( .A(\stack[1][8] ), .B(o[21]), .Z(n4050) );
  OR U4303 ( .A(n4005), .B(n4004), .Z(n4009) );
  OR U4304 ( .A(n4007), .B(n4006), .Z(n4008) );
  NAND U4305 ( .A(n4009), .B(n4008), .Z(n4051) );
  XOR U4306 ( .A(n4050), .B(n4051), .Z(n4053) );
  XNOR U4307 ( .A(n4052), .B(n4053), .Z(n4177) );
  XNOR U4308 ( .A(n4178), .B(n4177), .Z(n4179) );
  XNOR U4309 ( .A(n4180), .B(n4179), .Z(n4046) );
  NAND U4310 ( .A(\stack[1][6] ), .B(o[23]), .Z(n4044) );
  OR U4311 ( .A(n4011), .B(n4010), .Z(n4015) );
  OR U4312 ( .A(n4013), .B(n4012), .Z(n4014) );
  NAND U4313 ( .A(n4015), .B(n4014), .Z(n4045) );
  XOR U4314 ( .A(n4044), .B(n4045), .Z(n4047) );
  XNOR U4315 ( .A(n4046), .B(n4047), .Z(n4183) );
  XNOR U4316 ( .A(n4184), .B(n4183), .Z(n4185) );
  XNOR U4317 ( .A(n4186), .B(n4185), .Z(n4040) );
  ANDN U4318 ( .B(\stack[1][4] ), .A(n4016), .Z(n4038) );
  OR U4319 ( .A(n4018), .B(n4017), .Z(n4022) );
  OR U4320 ( .A(n4020), .B(n4019), .Z(n4021) );
  NAND U4321 ( .A(n4022), .B(n4021), .Z(n4039) );
  XNOR U4322 ( .A(n4038), .B(n4039), .Z(n4041) );
  XNOR U4323 ( .A(n4040), .B(n4041), .Z(n4189) );
  XNOR U4324 ( .A(n4190), .B(n4189), .Z(n4191) );
  XOR U4325 ( .A(n4192), .B(n4191), .Z(n4035) );
  ANDN U4326 ( .B(\stack[1][2] ), .A(n4023), .Z(n4032) );
  OR U4327 ( .A(n4025), .B(n4024), .Z(n4029) );
  NANDN U4328 ( .A(n4027), .B(n4026), .Z(n4028) );
  NAND U4329 ( .A(n4029), .B(n4028), .Z(n4033) );
  XOR U4330 ( .A(n4032), .B(n4033), .Z(n4034) );
  XNOR U4331 ( .A(n4035), .B(n4034), .Z(n4196) );
  XNOR U4332 ( .A(n4197), .B(n4196), .Z(n4198) );
  XOR U4333 ( .A(n4199), .B(n4198), .Z(n4571) );
  OR U4334 ( .A(n4570), .B(n4571), .Z(n4030) );
  AND U4335 ( .A(n4031), .B(n4030), .Z(n4202) );
  NAND U4336 ( .A(\stack[1][2] ), .B(o[28]), .Z(n4215) );
  OR U4337 ( .A(n4033), .B(n4032), .Z(n4037) );
  NANDN U4338 ( .A(n4035), .B(n4034), .Z(n4036) );
  NAND U4339 ( .A(n4037), .B(n4036), .Z(n4217) );
  NAND U4340 ( .A(\stack[1][4] ), .B(o[26]), .Z(n4475) );
  OR U4341 ( .A(n4039), .B(n4038), .Z(n4043) );
  NANDN U4342 ( .A(n4041), .B(n4040), .Z(n4042) );
  NAND U4343 ( .A(n4043), .B(n4042), .Z(n4477) );
  NAND U4344 ( .A(\stack[1][6] ), .B(o[24]), .Z(n4467) );
  NANDN U4345 ( .A(n4045), .B(n4044), .Z(n4049) );
  NANDN U4346 ( .A(n4047), .B(n4046), .Z(n4048) );
  NAND U4347 ( .A(n4049), .B(n4048), .Z(n4469) );
  NAND U4348 ( .A(\stack[1][8] ), .B(o[22]), .Z(n4455) );
  NANDN U4349 ( .A(n4051), .B(n4050), .Z(n4055) );
  NANDN U4350 ( .A(n4053), .B(n4052), .Z(n4054) );
  NAND U4351 ( .A(n4055), .B(n4054), .Z(n4457) );
  ANDN U4352 ( .B(o[20]), .A(n1615), .Z(n4437) );
  OR U4353 ( .A(n4057), .B(n4056), .Z(n4061) );
  OR U4354 ( .A(n4059), .B(n4058), .Z(n4060) );
  AND U4355 ( .A(n4061), .B(n4060), .Z(n4438) );
  OR U4356 ( .A(n4063), .B(n4062), .Z(n4067) );
  NANDN U4357 ( .A(n4065), .B(n4064), .Z(n4066) );
  AND U4358 ( .A(n4067), .B(n4066), .Z(n4230) );
  ANDN U4359 ( .B(\stack[1][11] ), .A(n4068), .Z(n4231) );
  XNOR U4360 ( .A(n4230), .B(n4231), .Z(n4229) );
  NANDN U4361 ( .A(n4070), .B(n4069), .Z(n4074) );
  OR U4362 ( .A(n4072), .B(n4071), .Z(n4073) );
  NAND U4363 ( .A(n4074), .B(n4073), .Z(n4421) );
  AND U4364 ( .A(o[17]), .B(\stack[1][13] ), .Z(n4420) );
  XNOR U4365 ( .A(n4421), .B(n4420), .Z(n4418) );
  NAND U4366 ( .A(\stack[1][14] ), .B(o[16]), .Z(n4235) );
  NANDN U4367 ( .A(n4076), .B(n4075), .Z(n4080) );
  NANDN U4368 ( .A(n4078), .B(n4077), .Z(n4079) );
  AND U4369 ( .A(n4080), .B(n4079), .Z(n4236) );
  NAND U4370 ( .A(\stack[1][16] ), .B(o[14]), .Z(n4401) );
  OR U4371 ( .A(n4082), .B(n4081), .Z(n4086) );
  OR U4372 ( .A(n4084), .B(n4083), .Z(n4085) );
  NAND U4373 ( .A(n4086), .B(n4085), .Z(n4403) );
  NAND U4374 ( .A(o[12]), .B(\stack[1][18] ), .Z(n4247) );
  NANDN U4375 ( .A(n4088), .B(n4087), .Z(n4092) );
  NANDN U4376 ( .A(n4090), .B(n4089), .Z(n4091) );
  AND U4377 ( .A(n4092), .B(n4091), .Z(n4249) );
  NAND U4378 ( .A(o[10]), .B(\stack[1][20] ), .Z(n4384) );
  OR U4379 ( .A(n4094), .B(n4093), .Z(n4098) );
  NANDN U4380 ( .A(n4096), .B(n4095), .Z(n4097) );
  NAND U4381 ( .A(n4098), .B(n4097), .Z(n4386) );
  NAND U4382 ( .A(o[8]), .B(\stack[1][22] ), .Z(n4253) );
  OR U4383 ( .A(n4100), .B(n4099), .Z(n4104) );
  OR U4384 ( .A(n4102), .B(n4101), .Z(n4103) );
  NAND U4385 ( .A(n4104), .B(n4103), .Z(n4255) );
  OR U4386 ( .A(n4106), .B(n4105), .Z(n4110) );
  NANDN U4387 ( .A(n4108), .B(n4107), .Z(n4109) );
  AND U4388 ( .A(n4110), .B(n4109), .Z(n4367) );
  ANDN U4389 ( .B(\stack[1][23] ), .A(n4111), .Z(n4368) );
  XNOR U4390 ( .A(n4367), .B(n4368), .Z(n4366) );
  OR U4391 ( .A(n4113), .B(n4112), .Z(n4117) );
  OR U4392 ( .A(n4115), .B(n4114), .Z(n4116) );
  AND U4393 ( .A(n4117), .B(n4116), .Z(n4343) );
  OR U4394 ( .A(n4119), .B(n4118), .Z(n4123) );
  OR U4395 ( .A(n4121), .B(n4120), .Z(n4122) );
  NAND U4396 ( .A(n4123), .B(n4122), .Z(n4261) );
  ANDN U4397 ( .B(\stack[1][27] ), .A(n4127), .Z(n4286) );
  XNOR U4398 ( .A(n4285), .B(n4286), .Z(n4284) );
  AND U4399 ( .A(\stack[1][29] ), .B(o[1]), .Z(n4266) );
  NAND U4400 ( .A(o[0]), .B(\stack[1][30] ), .Z(n4128) );
  XNOR U4401 ( .A(n4266), .B(n4128), .Z(n4265) );
  XOR U4402 ( .A(n4265), .B(n4264), .Z(n4283) );
  XOR U4403 ( .A(n4284), .B(n4283), .Z(n4260) );
  XNOR U4404 ( .A(n4261), .B(n4260), .Z(n4259) );
  ANDN U4405 ( .B(\stack[1][26] ), .A(n4129), .Z(n4258) );
  XNOR U4406 ( .A(n4259), .B(n4258), .Z(n4347) );
  ANDN U4407 ( .B(\stack[1][25] ), .A(n4130), .Z(n4349) );
  OR U4408 ( .A(n4132), .B(n4131), .Z(n4136) );
  NANDN U4409 ( .A(n4134), .B(n4133), .Z(n4135) );
  NAND U4410 ( .A(n4136), .B(n4135), .Z(n4350) );
  XNOR U4411 ( .A(n4349), .B(n4350), .Z(n4348) );
  XNOR U4412 ( .A(n4347), .B(n4348), .Z(n4344) );
  XOR U4413 ( .A(n4343), .B(n4344), .Z(n4341) );
  ANDN U4414 ( .B(\stack[1][24] ), .A(n4137), .Z(n4342) );
  XOR U4415 ( .A(n4341), .B(n4342), .Z(n4365) );
  XOR U4416 ( .A(n4366), .B(n4365), .Z(n4254) );
  XNOR U4417 ( .A(n4255), .B(n4254), .Z(n4252) );
  XNOR U4418 ( .A(n4253), .B(n4252), .Z(n4359) );
  NAND U4419 ( .A(\stack[1][21] ), .B(o[9]), .Z(n4361) );
  OR U4420 ( .A(n4139), .B(n4138), .Z(n4143) );
  OR U4421 ( .A(n4141), .B(n4140), .Z(n4142) );
  NAND U4422 ( .A(n4143), .B(n4142), .Z(n4362) );
  XOR U4423 ( .A(n4361), .B(n4362), .Z(n4360) );
  XNOR U4424 ( .A(n4359), .B(n4360), .Z(n4385) );
  XNOR U4425 ( .A(n4386), .B(n4385), .Z(n4383) );
  XNOR U4426 ( .A(n4384), .B(n4383), .Z(n4377) );
  ANDN U4427 ( .B(\stack[1][19] ), .A(n4144), .Z(n4379) );
  OR U4428 ( .A(n4146), .B(n4145), .Z(n4150) );
  OR U4429 ( .A(n4148), .B(n4147), .Z(n4149) );
  NAND U4430 ( .A(n4150), .B(n4149), .Z(n4380) );
  XNOR U4431 ( .A(n4379), .B(n4380), .Z(n4378) );
  XNOR U4432 ( .A(n4249), .B(n4248), .Z(n4246) );
  XNOR U4433 ( .A(n4247), .B(n4246), .Z(n4240) );
  OR U4434 ( .A(n4152), .B(n4151), .Z(n4156) );
  OR U4435 ( .A(n4154), .B(n4153), .Z(n4155) );
  AND U4436 ( .A(n4156), .B(n4155), .Z(n4242) );
  NAND U4437 ( .A(\stack[1][17] ), .B(o[13]), .Z(n4243) );
  XOR U4438 ( .A(n4242), .B(n4243), .Z(n4241) );
  XNOR U4439 ( .A(n4240), .B(n4241), .Z(n4402) );
  XNOR U4440 ( .A(n4403), .B(n4402), .Z(n4400) );
  XNOR U4441 ( .A(n4401), .B(n4400), .Z(n4395) );
  ANDN U4442 ( .B(o[15]), .A(n4157), .Z(n5102) );
  OR U4443 ( .A(n4159), .B(n4158), .Z(n4163) );
  NANDN U4444 ( .A(n4161), .B(n4160), .Z(n4162) );
  NAND U4445 ( .A(n4163), .B(n4162), .Z(n4397) );
  XNOR U4446 ( .A(n5102), .B(n4397), .Z(n4396) );
  XNOR U4447 ( .A(n4395), .B(n4396), .Z(n4237) );
  XOR U4448 ( .A(n4236), .B(n4237), .Z(n4234) );
  XOR U4449 ( .A(n4418), .B(n4419), .Z(n4414) );
  OR U4450 ( .A(n4165), .B(n4164), .Z(n4169) );
  NANDN U4451 ( .A(n4167), .B(n4166), .Z(n4168) );
  AND U4452 ( .A(n4169), .B(n4168), .Z(n4415) );
  XOR U4453 ( .A(n4414), .B(n4415), .Z(n4413) );
  ANDN U4454 ( .B(o[18]), .A(n1617), .Z(n4412) );
  XOR U4455 ( .A(n4413), .B(n4412), .Z(n4228) );
  XOR U4456 ( .A(n4229), .B(n4228), .Z(n4439) );
  XOR U4457 ( .A(n4438), .B(n4439), .Z(n4436) );
  XOR U4458 ( .A(n4437), .B(n4436), .Z(n4431) );
  ANDN U4459 ( .B(\stack[1][9] ), .A(n4170), .Z(n4432) );
  OR U4460 ( .A(n4172), .B(n4171), .Z(n4176) );
  OR U4461 ( .A(n4174), .B(n4173), .Z(n4175) );
  NAND U4462 ( .A(n4176), .B(n4175), .Z(n4433) );
  XNOR U4463 ( .A(n4432), .B(n4433), .Z(n4430) );
  XOR U4464 ( .A(n4431), .B(n4430), .Z(n4456) );
  XNOR U4465 ( .A(n4457), .B(n4456), .Z(n4454) );
  XNOR U4466 ( .A(n4455), .B(n4454), .Z(n4448) );
  NAND U4467 ( .A(\stack[1][7] ), .B(o[23]), .Z(n4450) );
  OR U4468 ( .A(n4178), .B(n4177), .Z(n4182) );
  OR U4469 ( .A(n4180), .B(n4179), .Z(n4181) );
  NAND U4470 ( .A(n4182), .B(n4181), .Z(n4451) );
  XOR U4471 ( .A(n4450), .B(n4451), .Z(n4449) );
  XNOR U4472 ( .A(n4448), .B(n4449), .Z(n4468) );
  XNOR U4473 ( .A(n4469), .B(n4468), .Z(n4466) );
  XNOR U4474 ( .A(n4467), .B(n4466), .Z(n4483) );
  NAND U4475 ( .A(\stack[1][5] ), .B(o[25]), .Z(n4481) );
  OR U4476 ( .A(n4184), .B(n4183), .Z(n4188) );
  OR U4477 ( .A(n4186), .B(n4185), .Z(n4187) );
  NAND U4478 ( .A(n4188), .B(n4187), .Z(n4480) );
  XOR U4479 ( .A(n4481), .B(n4480), .Z(n4482) );
  XNOR U4480 ( .A(n4483), .B(n4482), .Z(n4476) );
  XNOR U4481 ( .A(n4477), .B(n4476), .Z(n4474) );
  XNOR U4482 ( .A(n4475), .B(n4474), .Z(n4222) );
  NAND U4483 ( .A(\stack[1][3] ), .B(o[27]), .Z(n4225) );
  OR U4484 ( .A(n4190), .B(n4189), .Z(n4194) );
  OR U4485 ( .A(n4192), .B(n4191), .Z(n4193) );
  NAND U4486 ( .A(n4194), .B(n4193), .Z(n4224) );
  XOR U4487 ( .A(n4225), .B(n4224), .Z(n4223) );
  XNOR U4488 ( .A(n4222), .B(n4223), .Z(n4216) );
  XOR U4489 ( .A(n4217), .B(n4216), .Z(n4214) );
  XNOR U4490 ( .A(n4215), .B(n4214), .Z(n4206) );
  ANDN U4491 ( .B(o[29]), .A(n4195), .Z(n4208) );
  OR U4492 ( .A(n4197), .B(n4196), .Z(n4201) );
  OR U4493 ( .A(n4199), .B(n4198), .Z(n4200) );
  NAND U4494 ( .A(n4201), .B(n4200), .Z(n4209) );
  XNOR U4495 ( .A(n4208), .B(n4209), .Z(n4207) );
  XNOR U4496 ( .A(n4206), .B(n4207), .Z(n4203) );
  XNOR U4497 ( .A(n4202), .B(n4203), .Z(n4532) );
  ANDN U4498 ( .B(o[30]), .A(n1606), .Z(n4533) );
  OR U4499 ( .A(n4532), .B(n4533), .Z(n4205) );
  OR U4500 ( .A(n4203), .B(n4202), .Z(n4204) );
  AND U4501 ( .A(n4205), .B(n4204), .Z(n4213) );
  OR U4502 ( .A(n4207), .B(n4206), .Z(n4211) );
  OR U4503 ( .A(n4209), .B(n4208), .Z(n4210) );
  NAND U4504 ( .A(n4211), .B(n4210), .Z(n4212) );
  XNOR U4505 ( .A(n4213), .B(n4212), .Z(n4221) );
  NANDN U4506 ( .A(n4215), .B(n4214), .Z(n4219) );
  OR U4507 ( .A(n4217), .B(n4216), .Z(n4218) );
  NAND U4508 ( .A(n4219), .B(n4218), .Z(n4220) );
  XNOR U4509 ( .A(n4221), .B(n4220), .Z(n4493) );
  NANDN U4510 ( .A(n4223), .B(n4222), .Z(n4227) );
  ANDN U4511 ( .B(n4225), .A(n4224), .Z(n4226) );
  ANDN U4512 ( .B(n4227), .A(n4226), .Z(n4491) );
  NANDN U4513 ( .A(n4229), .B(n4228), .Z(n4233) );
  OR U4514 ( .A(n4231), .B(n4230), .Z(n4232) );
  AND U4515 ( .A(n4233), .B(n4232), .Z(n4465) );
  NANDN U4516 ( .A(n4235), .B(n4234), .Z(n4239) );
  OR U4517 ( .A(n4237), .B(n4236), .Z(n4238) );
  AND U4518 ( .A(n4239), .B(n4238), .Z(n4447) );
  NANDN U4519 ( .A(n4241), .B(n4240), .Z(n4245) );
  ANDN U4520 ( .B(n4243), .A(n4242), .Z(n4244) );
  ANDN U4521 ( .B(n4245), .A(n4244), .Z(n4429) );
  OR U4522 ( .A(n4247), .B(n4246), .Z(n4251) );
  NOR U4523 ( .A(n4249), .B(n4248), .Z(n4250) );
  ANDN U4524 ( .B(n4251), .A(n4250), .Z(n4411) );
  OR U4525 ( .A(n4253), .B(n4252), .Z(n4257) );
  OR U4526 ( .A(n4255), .B(n4254), .Z(n4256) );
  AND U4527 ( .A(n4257), .B(n4256), .Z(n4394) );
  NANDN U4528 ( .A(n4259), .B(n4258), .Z(n4263) );
  OR U4529 ( .A(n4261), .B(n4260), .Z(n4262) );
  AND U4530 ( .A(n4263), .B(n4262), .Z(n4376) );
  NANDN U4531 ( .A(n4265), .B(n4264), .Z(n4268) );
  ANDN U4532 ( .B(n4268), .A(n4267), .Z(n4358) );
  AND U4533 ( .A(o[29]), .B(\stack[1][2] ), .Z(n4270) );
  NAND U4534 ( .A(\stack[1][1] ), .B(o[30]), .Z(n4269) );
  XNOR U4535 ( .A(n4270), .B(n4269), .Z(n4274) );
  AND U4536 ( .A(\stack[1][7] ), .B(o[24]), .Z(n4272) );
  NAND U4537 ( .A(\stack[1][3] ), .B(o[28]), .Z(n4271) );
  XNOR U4538 ( .A(n4272), .B(n4271), .Z(n4273) );
  XOR U4539 ( .A(n4274), .B(n4273), .Z(n4282) );
  AND U4540 ( .A(\stack[1][9] ), .B(o[22]), .Z(n4276) );
  NAND U4541 ( .A(\stack[1][5] ), .B(o[26]), .Z(n4275) );
  XNOR U4542 ( .A(n4276), .B(n4275), .Z(n4280) );
  AND U4543 ( .A(o[19]), .B(\stack[1][12] ), .Z(n4278) );
  NAND U4544 ( .A(o[25]), .B(\stack[1][6] ), .Z(n4277) );
  XNOR U4545 ( .A(n4278), .B(n4277), .Z(n4279) );
  XNOR U4546 ( .A(n4280), .B(n4279), .Z(n4281) );
  XNOR U4547 ( .A(n4282), .B(n4281), .Z(n4322) );
  OR U4548 ( .A(n4284), .B(n4283), .Z(n4288) );
  OR U4549 ( .A(n4286), .B(n4285), .Z(n4287) );
  AND U4550 ( .A(n4288), .B(n4287), .Z(n4320) );
  AND U4551 ( .A(\stack[1][13] ), .B(o[18]), .Z(n4290) );
  NAND U4552 ( .A(o[21]), .B(\stack[1][10] ), .Z(n4289) );
  XNOR U4553 ( .A(n4290), .B(n4289), .Z(n4294) );
  AND U4554 ( .A(\stack[1][11] ), .B(o[20]), .Z(n4292) );
  NAND U4555 ( .A(o[8]), .B(\stack[1][23] ), .Z(n4291) );
  XNOR U4556 ( .A(n4292), .B(n4291), .Z(n4293) );
  XOR U4557 ( .A(n4294), .B(n4293), .Z(n4302) );
  AND U4558 ( .A(o[4]), .B(\stack[1][27] ), .Z(n4296) );
  NAND U4559 ( .A(o[3]), .B(\stack[1][28] ), .Z(n4295) );
  XNOR U4560 ( .A(n4296), .B(n4295), .Z(n4300) );
  AND U4561 ( .A(o[5]), .B(\stack[1][26] ), .Z(n4298) );
  NAND U4562 ( .A(\stack[1][31] ), .B(o[0]), .Z(n4297) );
  XNOR U4563 ( .A(n4298), .B(n4297), .Z(n4299) );
  XNOR U4564 ( .A(n4300), .B(n4299), .Z(n4301) );
  XNOR U4565 ( .A(n4302), .B(n4301), .Z(n4318) );
  AND U4566 ( .A(o[10]), .B(\stack[1][21] ), .Z(n4304) );
  NAND U4567 ( .A(o[7]), .B(\stack[1][24] ), .Z(n4303) );
  XNOR U4568 ( .A(n4304), .B(n4303), .Z(n4308) );
  AND U4569 ( .A(o[12]), .B(\stack[1][19] ), .Z(n4306) );
  NAND U4570 ( .A(o[6]), .B(\stack[1][25] ), .Z(n4305) );
  XNOR U4571 ( .A(n4306), .B(n4305), .Z(n4307) );
  XOR U4572 ( .A(n4308), .B(n4307), .Z(n4316) );
  AND U4573 ( .A(o[14]), .B(\stack[1][17] ), .Z(n4310) );
  NAND U4574 ( .A(o[11]), .B(\stack[1][20] ), .Z(n4309) );
  XNOR U4575 ( .A(n4310), .B(n4309), .Z(n4314) );
  AND U4576 ( .A(o[9]), .B(\stack[1][22] ), .Z(n4312) );
  NAND U4577 ( .A(o[17]), .B(\stack[1][14] ), .Z(n4311) );
  XNOR U4578 ( .A(n4312), .B(n4311), .Z(n4313) );
  XNOR U4579 ( .A(n4314), .B(n4313), .Z(n4315) );
  XNOR U4580 ( .A(n4316), .B(n4315), .Z(n4317) );
  XNOR U4581 ( .A(n4318), .B(n4317), .Z(n4319) );
  XNOR U4582 ( .A(n4320), .B(n4319), .Z(n4321) );
  XOR U4583 ( .A(n4322), .B(n4321), .Z(n4340) );
  AND U4584 ( .A(\stack[1][30] ), .B(o[1]), .Z(n4330) );
  NAND U4585 ( .A(o[0]), .B(n4330), .Z(n4323) );
  XNOR U4586 ( .A(o[2]), .B(n4323), .Z(n4324) );
  NAND U4587 ( .A(n4324), .B(\stack[1][29] ), .Z(n4338) );
  AND U4588 ( .A(o[31]), .B(\stack[1][0] ), .Z(n4336) );
  AND U4589 ( .A(o[15]), .B(\stack[1][16] ), .Z(n4326) );
  NAND U4590 ( .A(o[23]), .B(\stack[1][8] ), .Z(n4325) );
  XNOR U4591 ( .A(n4326), .B(n4325), .Z(n4334) );
  AND U4592 ( .A(o[27]), .B(\stack[1][4] ), .Z(n4332) );
  AND U4593 ( .A(\stack[1][15] ), .B(o[16]), .Z(n4328) );
  NAND U4594 ( .A(o[13]), .B(\stack[1][18] ), .Z(n4327) );
  XNOR U4595 ( .A(n4328), .B(n4327), .Z(n4329) );
  XNOR U4596 ( .A(n4330), .B(n4329), .Z(n4331) );
  XNOR U4597 ( .A(n4332), .B(n4331), .Z(n4333) );
  XNOR U4598 ( .A(n4334), .B(n4333), .Z(n4335) );
  XNOR U4599 ( .A(n4336), .B(n4335), .Z(n4337) );
  XNOR U4600 ( .A(n4338), .B(n4337), .Z(n4339) );
  XNOR U4601 ( .A(n4340), .B(n4339), .Z(n4356) );
  NANDN U4602 ( .A(n4342), .B(n4341), .Z(n4346) );
  OR U4603 ( .A(n4344), .B(n4343), .Z(n4345) );
  AND U4604 ( .A(n4346), .B(n4345), .Z(n4354) );
  OR U4605 ( .A(n4348), .B(n4347), .Z(n4352) );
  OR U4606 ( .A(n4350), .B(n4349), .Z(n4351) );
  NAND U4607 ( .A(n4352), .B(n4351), .Z(n4353) );
  XNOR U4608 ( .A(n4354), .B(n4353), .Z(n4355) );
  XNOR U4609 ( .A(n4356), .B(n4355), .Z(n4357) );
  XNOR U4610 ( .A(n4358), .B(n4357), .Z(n4374) );
  NANDN U4611 ( .A(n4360), .B(n4359), .Z(n4364) );
  NANDN U4612 ( .A(n4362), .B(n4361), .Z(n4363) );
  AND U4613 ( .A(n4364), .B(n4363), .Z(n4372) );
  OR U4614 ( .A(n4366), .B(n4365), .Z(n4370) );
  OR U4615 ( .A(n4368), .B(n4367), .Z(n4369) );
  NAND U4616 ( .A(n4370), .B(n4369), .Z(n4371) );
  XNOR U4617 ( .A(n4372), .B(n4371), .Z(n4373) );
  XNOR U4618 ( .A(n4374), .B(n4373), .Z(n4375) );
  XNOR U4619 ( .A(n4376), .B(n4375), .Z(n4392) );
  NANDN U4620 ( .A(n4378), .B(n4377), .Z(n4382) );
  OR U4621 ( .A(n4380), .B(n4379), .Z(n4381) );
  AND U4622 ( .A(n4382), .B(n4381), .Z(n4390) );
  OR U4623 ( .A(n4384), .B(n4383), .Z(n4388) );
  OR U4624 ( .A(n4386), .B(n4385), .Z(n4387) );
  NAND U4625 ( .A(n4388), .B(n4387), .Z(n4389) );
  XNOR U4626 ( .A(n4390), .B(n4389), .Z(n4391) );
  XNOR U4627 ( .A(n4392), .B(n4391), .Z(n4393) );
  XNOR U4628 ( .A(n4394), .B(n4393), .Z(n4409) );
  NANDN U4629 ( .A(n4396), .B(n4395), .Z(n4399) );
  OR U4630 ( .A(n4397), .B(n5102), .Z(n4398) );
  AND U4631 ( .A(n4399), .B(n4398), .Z(n4407) );
  OR U4632 ( .A(n4401), .B(n4400), .Z(n4405) );
  OR U4633 ( .A(n4403), .B(n4402), .Z(n4404) );
  NAND U4634 ( .A(n4405), .B(n4404), .Z(n4406) );
  XNOR U4635 ( .A(n4407), .B(n4406), .Z(n4408) );
  XNOR U4636 ( .A(n4409), .B(n4408), .Z(n4410) );
  XNOR U4637 ( .A(n4411), .B(n4410), .Z(n4427) );
  OR U4638 ( .A(n4413), .B(n4412), .Z(n4417) );
  NANDN U4639 ( .A(n4415), .B(n4414), .Z(n4416) );
  AND U4640 ( .A(n4417), .B(n4416), .Z(n4425) );
  NANDN U4641 ( .A(n4419), .B(n4418), .Z(n4423) );
  NANDN U4642 ( .A(n4421), .B(n4420), .Z(n4422) );
  NAND U4643 ( .A(n4423), .B(n4422), .Z(n4424) );
  XNOR U4644 ( .A(n4425), .B(n4424), .Z(n4426) );
  XNOR U4645 ( .A(n4427), .B(n4426), .Z(n4428) );
  XNOR U4646 ( .A(n4429), .B(n4428), .Z(n4445) );
  OR U4647 ( .A(n4431), .B(n4430), .Z(n4435) );
  OR U4648 ( .A(n4433), .B(n4432), .Z(n4434) );
  AND U4649 ( .A(n4435), .B(n4434), .Z(n4443) );
  NANDN U4650 ( .A(n4437), .B(n4436), .Z(n4441) );
  OR U4651 ( .A(n4439), .B(n4438), .Z(n4440) );
  NAND U4652 ( .A(n4441), .B(n4440), .Z(n4442) );
  XNOR U4653 ( .A(n4443), .B(n4442), .Z(n4444) );
  XNOR U4654 ( .A(n4445), .B(n4444), .Z(n4446) );
  XNOR U4655 ( .A(n4447), .B(n4446), .Z(n4463) );
  NANDN U4656 ( .A(n4449), .B(n4448), .Z(n4453) );
  NANDN U4657 ( .A(n4451), .B(n4450), .Z(n4452) );
  AND U4658 ( .A(n4453), .B(n4452), .Z(n4461) );
  OR U4659 ( .A(n4455), .B(n4454), .Z(n4459) );
  OR U4660 ( .A(n4457), .B(n4456), .Z(n4458) );
  NAND U4661 ( .A(n4459), .B(n4458), .Z(n4460) );
  XNOR U4662 ( .A(n4461), .B(n4460), .Z(n4462) );
  XNOR U4663 ( .A(n4463), .B(n4462), .Z(n4464) );
  XNOR U4664 ( .A(n4465), .B(n4464), .Z(n4473) );
  OR U4665 ( .A(n4467), .B(n4466), .Z(n4471) );
  OR U4666 ( .A(n4469), .B(n4468), .Z(n4470) );
  NAND U4667 ( .A(n4471), .B(n4470), .Z(n4472) );
  XNOR U4668 ( .A(n4473), .B(n4472), .Z(n4489) );
  OR U4669 ( .A(n4475), .B(n4474), .Z(n4479) );
  NOR U4670 ( .A(n4477), .B(n4476), .Z(n4478) );
  ANDN U4671 ( .B(n4479), .A(n4478), .Z(n4487) );
  ANDN U4672 ( .B(n4481), .A(n4480), .Z(n4485) );
  ANDN U4673 ( .B(n4483), .A(n4482), .Z(n4484) );
  OR U4674 ( .A(n4485), .B(n4484), .Z(n4486) );
  XNOR U4675 ( .A(n4487), .B(n4486), .Z(n4488) );
  XNOR U4676 ( .A(n4489), .B(n4488), .Z(n4490) );
  XNOR U4677 ( .A(n4491), .B(n4490), .Z(n4492) );
  XOR U4678 ( .A(n4493), .B(n4492), .Z(n4494) );
  AND U4679 ( .A(opcode[1]), .B(opcode[0]), .Z(n5664) );
  ANDN U4680 ( .B(n5664), .A(opcode[2]), .Z(n5644) );
  NAND U4681 ( .A(n4494), .B(n5644), .Z(n4495) );
  NANDN U4682 ( .A(n4496), .B(n4495), .Z(n4505) );
  XNOR U4683 ( .A(opcode[2]), .B(opcode[1]), .Z(n4497) );
  AND U4684 ( .A(n4498), .B(n4497), .Z(n5663) );
  NAND U4685 ( .A(n5663), .B(o[31]), .Z(n4503) );
  NAND U4686 ( .A(opcode[2]), .B(n5664), .Z(n5667) );
  ANDN U4687 ( .B(opcode[2]), .A(n4499), .Z(n5665) );
  NAND U4688 ( .A(o[31]), .B(n5665), .Z(n4500) );
  NAND U4689 ( .A(n5667), .B(n4500), .Z(n4501) );
  AND U4690 ( .A(\stack[1][31] ), .B(n4501), .Z(n4502) );
  ANDN U4691 ( .B(n4503), .A(n4502), .Z(n4504) );
  NANDN U4692 ( .A(n4505), .B(n4504), .Z(n1078) );
  NAND U4693 ( .A(n5672), .B(\stack[6][30] ), .Z(n4507) );
  NAND U4694 ( .A(n1605), .B(\stack[7][30] ), .Z(n4506) );
  NAND U4695 ( .A(n4507), .B(n4506), .Z(n1079) );
  NAND U4696 ( .A(n5672), .B(\stack[5][30] ), .Z(n4509) );
  NANDN U4697 ( .A(n5657), .B(\stack[7][30] ), .Z(n4508) );
  AND U4698 ( .A(n4509), .B(n4508), .Z(n4511) );
  NANDN U4699 ( .A(n5660), .B(\stack[6][30] ), .Z(n4510) );
  NAND U4700 ( .A(n4511), .B(n4510), .Z(n1080) );
  NAND U4701 ( .A(n5672), .B(\stack[4][30] ), .Z(n4513) );
  NANDN U4702 ( .A(n5657), .B(\stack[6][30] ), .Z(n4512) );
  AND U4703 ( .A(n4513), .B(n4512), .Z(n4515) );
  NANDN U4704 ( .A(n5660), .B(\stack[5][30] ), .Z(n4514) );
  NAND U4705 ( .A(n4515), .B(n4514), .Z(n1081) );
  NAND U4706 ( .A(n5672), .B(\stack[3][30] ), .Z(n4517) );
  NANDN U4707 ( .A(n5657), .B(\stack[5][30] ), .Z(n4516) );
  AND U4708 ( .A(n4517), .B(n4516), .Z(n4519) );
  NANDN U4709 ( .A(n5660), .B(\stack[4][30] ), .Z(n4518) );
  NAND U4710 ( .A(n4519), .B(n4518), .Z(n1082) );
  NAND U4711 ( .A(n5672), .B(\stack[2][30] ), .Z(n4521) );
  NANDN U4712 ( .A(n5657), .B(\stack[4][30] ), .Z(n4520) );
  AND U4713 ( .A(n4521), .B(n4520), .Z(n4523) );
  NANDN U4714 ( .A(n5660), .B(\stack[3][30] ), .Z(n4522) );
  NAND U4715 ( .A(n4523), .B(n4522), .Z(n1083) );
  NAND U4716 ( .A(n5672), .B(\stack[1][30] ), .Z(n4525) );
  NANDN U4717 ( .A(n5657), .B(\stack[3][30] ), .Z(n4524) );
  AND U4718 ( .A(n4525), .B(n4524), .Z(n4527) );
  NANDN U4719 ( .A(n5660), .B(\stack[2][30] ), .Z(n4526) );
  NAND U4720 ( .A(n4527), .B(n4526), .Z(n1084) );
  NAND U4721 ( .A(n5672), .B(o[30]), .Z(n4529) );
  NANDN U4722 ( .A(n5657), .B(\stack[2][30] ), .Z(n4528) );
  AND U4723 ( .A(n4529), .B(n4528), .Z(n4531) );
  NANDN U4724 ( .A(n5660), .B(\stack[1][30] ), .Z(n4530) );
  NAND U4725 ( .A(n4531), .B(n4530), .Z(n1085) );
  XNOR U4726 ( .A(n4533), .B(n4532), .Z(n4534) );
  NAND U4727 ( .A(n4534), .B(n5644), .Z(n4537) );
  NAND U4728 ( .A(n5672), .B(x[30]), .Z(n4535) );
  NAND U4729 ( .A(n4537), .B(n4536), .Z(n4543) );
  NAND U4730 ( .A(n5663), .B(o[30]), .Z(n4541) );
  NAND U4731 ( .A(o[30]), .B(n5665), .Z(n4538) );
  NAND U4732 ( .A(n5667), .B(n4538), .Z(n4539) );
  AND U4733 ( .A(\stack[1][30] ), .B(n4539), .Z(n4540) );
  ANDN U4734 ( .B(n4541), .A(n4540), .Z(n4542) );
  NANDN U4735 ( .A(n4543), .B(n4542), .Z(n1086) );
  NAND U4736 ( .A(n5672), .B(\stack[6][29] ), .Z(n4545) );
  NAND U4737 ( .A(n1605), .B(\stack[7][29] ), .Z(n4544) );
  NAND U4738 ( .A(n4545), .B(n4544), .Z(n1087) );
  NAND U4739 ( .A(n5672), .B(\stack[5][29] ), .Z(n4547) );
  NANDN U4740 ( .A(n5657), .B(\stack[7][29] ), .Z(n4546) );
  AND U4741 ( .A(n4547), .B(n4546), .Z(n4549) );
  NANDN U4742 ( .A(n5660), .B(\stack[6][29] ), .Z(n4548) );
  NAND U4743 ( .A(n4549), .B(n4548), .Z(n1088) );
  NAND U4744 ( .A(n5672), .B(\stack[4][29] ), .Z(n4551) );
  NANDN U4745 ( .A(n5657), .B(\stack[6][29] ), .Z(n4550) );
  AND U4746 ( .A(n4551), .B(n4550), .Z(n4553) );
  NANDN U4747 ( .A(n5660), .B(\stack[5][29] ), .Z(n4552) );
  NAND U4748 ( .A(n4553), .B(n4552), .Z(n1089) );
  NAND U4749 ( .A(n5672), .B(\stack[3][29] ), .Z(n4555) );
  NANDN U4750 ( .A(n5657), .B(\stack[5][29] ), .Z(n4554) );
  AND U4751 ( .A(n4555), .B(n4554), .Z(n4557) );
  NANDN U4752 ( .A(n5660), .B(\stack[4][29] ), .Z(n4556) );
  NAND U4753 ( .A(n4557), .B(n4556), .Z(n1090) );
  NAND U4754 ( .A(n5672), .B(\stack[2][29] ), .Z(n4559) );
  NANDN U4755 ( .A(n5657), .B(\stack[4][29] ), .Z(n4558) );
  AND U4756 ( .A(n4559), .B(n4558), .Z(n4561) );
  NANDN U4757 ( .A(n5660), .B(\stack[3][29] ), .Z(n4560) );
  NAND U4758 ( .A(n4561), .B(n4560), .Z(n1091) );
  NAND U4759 ( .A(n5672), .B(\stack[1][29] ), .Z(n4563) );
  NANDN U4760 ( .A(n5657), .B(\stack[3][29] ), .Z(n4562) );
  AND U4761 ( .A(n4563), .B(n4562), .Z(n4565) );
  NANDN U4762 ( .A(n5660), .B(\stack[2][29] ), .Z(n4564) );
  NAND U4763 ( .A(n4565), .B(n4564), .Z(n1092) );
  NAND U4764 ( .A(o[29]), .B(n5672), .Z(n4567) );
  NANDN U4765 ( .A(n5657), .B(\stack[2][29] ), .Z(n4566) );
  AND U4766 ( .A(n4567), .B(n4566), .Z(n4569) );
  NANDN U4767 ( .A(n5660), .B(\stack[1][29] ), .Z(n4568) );
  NAND U4768 ( .A(n4569), .B(n4568), .Z(n1093) );
  XNOR U4769 ( .A(n4571), .B(n4570), .Z(n4572) );
  NAND U4770 ( .A(n4572), .B(n5644), .Z(n4576) );
  NAND U4771 ( .A(n5672), .B(x[29]), .Z(n4574) );
  IV U4772 ( .A(n5667), .Z(n5651) );
  NAND U4773 ( .A(n5651), .B(\stack[1][29] ), .Z(n4573) );
  AND U4774 ( .A(n4574), .B(n4573), .Z(n4575) );
  NAND U4775 ( .A(n4576), .B(n4575), .Z(n4581) );
  NAND U4776 ( .A(\stack[1][29] ), .B(n5665), .Z(n4577) );
  NAND U4777 ( .A(n1604), .B(n4577), .Z(n4578) );
  AND U4778 ( .A(n4578), .B(o[29]), .Z(n4579) );
  NANDN U4779 ( .A(n4581), .B(n4580), .Z(n1094) );
  NAND U4780 ( .A(n5672), .B(\stack[6][28] ), .Z(n4583) );
  NAND U4781 ( .A(n1605), .B(\stack[7][28] ), .Z(n4582) );
  NAND U4782 ( .A(n4583), .B(n4582), .Z(n1095) );
  NAND U4783 ( .A(n5672), .B(\stack[5][28] ), .Z(n4585) );
  NANDN U4784 ( .A(n5657), .B(\stack[7][28] ), .Z(n4584) );
  AND U4785 ( .A(n4585), .B(n4584), .Z(n4587) );
  NANDN U4786 ( .A(n5660), .B(\stack[6][28] ), .Z(n4586) );
  NAND U4787 ( .A(n4587), .B(n4586), .Z(n1096) );
  NAND U4788 ( .A(n5672), .B(\stack[4][28] ), .Z(n4589) );
  NANDN U4789 ( .A(n5657), .B(\stack[6][28] ), .Z(n4588) );
  AND U4790 ( .A(n4589), .B(n4588), .Z(n4591) );
  NANDN U4791 ( .A(n5660), .B(\stack[5][28] ), .Z(n4590) );
  NAND U4792 ( .A(n4591), .B(n4590), .Z(n1097) );
  NAND U4793 ( .A(n5672), .B(\stack[3][28] ), .Z(n4593) );
  NANDN U4794 ( .A(n5657), .B(\stack[5][28] ), .Z(n4592) );
  AND U4795 ( .A(n4593), .B(n4592), .Z(n4595) );
  NANDN U4796 ( .A(n5660), .B(\stack[4][28] ), .Z(n4594) );
  NAND U4797 ( .A(n4595), .B(n4594), .Z(n1098) );
  NAND U4798 ( .A(n5672), .B(\stack[2][28] ), .Z(n4597) );
  NANDN U4799 ( .A(n5657), .B(\stack[4][28] ), .Z(n4596) );
  AND U4800 ( .A(n4597), .B(n4596), .Z(n4599) );
  NANDN U4801 ( .A(n5660), .B(\stack[3][28] ), .Z(n4598) );
  NAND U4802 ( .A(n4599), .B(n4598), .Z(n1099) );
  NAND U4803 ( .A(\stack[1][28] ), .B(n5672), .Z(n4601) );
  NANDN U4804 ( .A(n5657), .B(\stack[3][28] ), .Z(n4600) );
  AND U4805 ( .A(n4601), .B(n4600), .Z(n4603) );
  NANDN U4806 ( .A(n5660), .B(\stack[2][28] ), .Z(n4602) );
  NAND U4807 ( .A(n4603), .B(n4602), .Z(n1100) );
  NAND U4808 ( .A(o[28]), .B(n5672), .Z(n4605) );
  NANDN U4809 ( .A(n5657), .B(\stack[2][28] ), .Z(n4604) );
  AND U4810 ( .A(n4605), .B(n4604), .Z(n4607) );
  NANDN U4811 ( .A(n5660), .B(\stack[1][28] ), .Z(n4606) );
  NAND U4812 ( .A(n4607), .B(n4606), .Z(n1101) );
  XNOR U4813 ( .A(n4609), .B(n4608), .Z(n4610) );
  NAND U4814 ( .A(n4610), .B(n5644), .Z(n4613) );
  NAND U4815 ( .A(n5672), .B(x[28]), .Z(n4611) );
  NAND U4816 ( .A(n4613), .B(n4612), .Z(n4619) );
  NAND U4817 ( .A(n5663), .B(o[28]), .Z(n4617) );
  NAND U4818 ( .A(o[28]), .B(n5665), .Z(n4614) );
  NAND U4819 ( .A(n5667), .B(n4614), .Z(n4615) );
  AND U4820 ( .A(n4615), .B(\stack[1][28] ), .Z(n4616) );
  ANDN U4821 ( .B(n4617), .A(n4616), .Z(n4618) );
  NANDN U4822 ( .A(n4619), .B(n4618), .Z(n1102) );
  NAND U4823 ( .A(n5672), .B(\stack[6][27] ), .Z(n4621) );
  NAND U4824 ( .A(n1605), .B(\stack[7][27] ), .Z(n4620) );
  NAND U4825 ( .A(n4621), .B(n4620), .Z(n1103) );
  NAND U4826 ( .A(n5672), .B(\stack[5][27] ), .Z(n4623) );
  NANDN U4827 ( .A(n5657), .B(\stack[7][27] ), .Z(n4622) );
  AND U4828 ( .A(n4623), .B(n4622), .Z(n4625) );
  NANDN U4829 ( .A(n5660), .B(\stack[6][27] ), .Z(n4624) );
  NAND U4830 ( .A(n4625), .B(n4624), .Z(n1104) );
  NAND U4831 ( .A(n5672), .B(\stack[4][27] ), .Z(n4627) );
  NANDN U4832 ( .A(n5657), .B(\stack[6][27] ), .Z(n4626) );
  AND U4833 ( .A(n4627), .B(n4626), .Z(n4629) );
  NANDN U4834 ( .A(n5660), .B(\stack[5][27] ), .Z(n4628) );
  NAND U4835 ( .A(n4629), .B(n4628), .Z(n1105) );
  NAND U4836 ( .A(n5672), .B(\stack[3][27] ), .Z(n4631) );
  NANDN U4837 ( .A(n5657), .B(\stack[5][27] ), .Z(n4630) );
  AND U4838 ( .A(n4631), .B(n4630), .Z(n4633) );
  NANDN U4839 ( .A(n5660), .B(\stack[4][27] ), .Z(n4632) );
  NAND U4840 ( .A(n4633), .B(n4632), .Z(n1106) );
  NAND U4841 ( .A(n5672), .B(\stack[2][27] ), .Z(n4635) );
  NANDN U4842 ( .A(n5657), .B(\stack[4][27] ), .Z(n4634) );
  AND U4843 ( .A(n4635), .B(n4634), .Z(n4637) );
  NANDN U4844 ( .A(n5660), .B(\stack[3][27] ), .Z(n4636) );
  NAND U4845 ( .A(n4637), .B(n4636), .Z(n1107) );
  NAND U4846 ( .A(\stack[1][27] ), .B(n5672), .Z(n4639) );
  NANDN U4847 ( .A(n5657), .B(\stack[3][27] ), .Z(n4638) );
  AND U4848 ( .A(n4639), .B(n4638), .Z(n4641) );
  NANDN U4849 ( .A(n5660), .B(\stack[2][27] ), .Z(n4640) );
  NAND U4850 ( .A(n4641), .B(n4640), .Z(n1108) );
  NAND U4851 ( .A(o[27]), .B(n5672), .Z(n4643) );
  NANDN U4852 ( .A(n5657), .B(\stack[2][27] ), .Z(n4642) );
  AND U4853 ( .A(n4643), .B(n4642), .Z(n4645) );
  NANDN U4854 ( .A(n5660), .B(\stack[1][27] ), .Z(n4644) );
  NAND U4855 ( .A(n4645), .B(n4644), .Z(n1109) );
  XNOR U4856 ( .A(n4647), .B(n4646), .Z(n4648) );
  NAND U4857 ( .A(n4648), .B(n5644), .Z(n4652) );
  NAND U4858 ( .A(n5672), .B(x[27]), .Z(n4650) );
  NAND U4859 ( .A(n5651), .B(\stack[1][27] ), .Z(n4649) );
  AND U4860 ( .A(n4650), .B(n4649), .Z(n4651) );
  NAND U4861 ( .A(n4652), .B(n4651), .Z(n4657) );
  NAND U4862 ( .A(\stack[1][27] ), .B(n5665), .Z(n4653) );
  NAND U4863 ( .A(n1604), .B(n4653), .Z(n4654) );
  AND U4864 ( .A(n4654), .B(o[27]), .Z(n4655) );
  NANDN U4865 ( .A(n4657), .B(n4656), .Z(n1110) );
  NAND U4866 ( .A(n5672), .B(\stack[6][26] ), .Z(n4659) );
  NAND U4867 ( .A(n1605), .B(\stack[7][26] ), .Z(n4658) );
  NAND U4868 ( .A(n4659), .B(n4658), .Z(n1111) );
  NAND U4869 ( .A(n5672), .B(\stack[5][26] ), .Z(n4661) );
  NANDN U4870 ( .A(n5657), .B(\stack[7][26] ), .Z(n4660) );
  AND U4871 ( .A(n4661), .B(n4660), .Z(n4663) );
  NANDN U4872 ( .A(n5660), .B(\stack[6][26] ), .Z(n4662) );
  NAND U4873 ( .A(n4663), .B(n4662), .Z(n1112) );
  NAND U4874 ( .A(n5672), .B(\stack[4][26] ), .Z(n4665) );
  NANDN U4875 ( .A(n5657), .B(\stack[6][26] ), .Z(n4664) );
  AND U4876 ( .A(n4665), .B(n4664), .Z(n4667) );
  NANDN U4877 ( .A(n5660), .B(\stack[5][26] ), .Z(n4666) );
  NAND U4878 ( .A(n4667), .B(n4666), .Z(n1113) );
  NAND U4879 ( .A(n5672), .B(\stack[3][26] ), .Z(n4669) );
  NANDN U4880 ( .A(n5657), .B(\stack[5][26] ), .Z(n4668) );
  AND U4881 ( .A(n4669), .B(n4668), .Z(n4671) );
  NANDN U4882 ( .A(n5660), .B(\stack[4][26] ), .Z(n4670) );
  NAND U4883 ( .A(n4671), .B(n4670), .Z(n1114) );
  NAND U4884 ( .A(n5672), .B(\stack[2][26] ), .Z(n4673) );
  NANDN U4885 ( .A(n5657), .B(\stack[4][26] ), .Z(n4672) );
  AND U4886 ( .A(n4673), .B(n4672), .Z(n4675) );
  NANDN U4887 ( .A(n5660), .B(\stack[3][26] ), .Z(n4674) );
  NAND U4888 ( .A(n4675), .B(n4674), .Z(n1115) );
  NAND U4889 ( .A(\stack[1][26] ), .B(n5672), .Z(n4677) );
  NANDN U4890 ( .A(n5657), .B(\stack[3][26] ), .Z(n4676) );
  AND U4891 ( .A(n4677), .B(n4676), .Z(n4679) );
  NANDN U4892 ( .A(n5660), .B(\stack[2][26] ), .Z(n4678) );
  NAND U4893 ( .A(n4679), .B(n4678), .Z(n1116) );
  NAND U4894 ( .A(o[26]), .B(n5672), .Z(n4681) );
  NANDN U4895 ( .A(n5657), .B(\stack[2][26] ), .Z(n4680) );
  AND U4896 ( .A(n4681), .B(n4680), .Z(n4683) );
  NANDN U4897 ( .A(n5660), .B(\stack[1][26] ), .Z(n4682) );
  NAND U4898 ( .A(n4683), .B(n4682), .Z(n1117) );
  XNOR U4899 ( .A(n4685), .B(n4684), .Z(n4686) );
  NAND U4900 ( .A(n4686), .B(n5644), .Z(n4689) );
  NAND U4901 ( .A(n5672), .B(x[26]), .Z(n4687) );
  NAND U4902 ( .A(n4689), .B(n4688), .Z(n4695) );
  NAND U4903 ( .A(n5663), .B(o[26]), .Z(n4693) );
  NAND U4904 ( .A(o[26]), .B(n5665), .Z(n4690) );
  NAND U4905 ( .A(n5667), .B(n4690), .Z(n4691) );
  AND U4906 ( .A(n4691), .B(\stack[1][26] ), .Z(n4692) );
  ANDN U4907 ( .B(n4693), .A(n4692), .Z(n4694) );
  NANDN U4908 ( .A(n4695), .B(n4694), .Z(n1118) );
  NAND U4909 ( .A(n5672), .B(\stack[6][25] ), .Z(n4697) );
  NAND U4910 ( .A(n1605), .B(\stack[7][25] ), .Z(n4696) );
  NAND U4911 ( .A(n4697), .B(n4696), .Z(n1119) );
  NAND U4912 ( .A(n5672), .B(\stack[5][25] ), .Z(n4699) );
  NANDN U4913 ( .A(n5657), .B(\stack[7][25] ), .Z(n4698) );
  AND U4914 ( .A(n4699), .B(n4698), .Z(n4701) );
  NANDN U4915 ( .A(n5660), .B(\stack[6][25] ), .Z(n4700) );
  NAND U4916 ( .A(n4701), .B(n4700), .Z(n1120) );
  NAND U4917 ( .A(n5672), .B(\stack[4][25] ), .Z(n4703) );
  NANDN U4918 ( .A(n5657), .B(\stack[6][25] ), .Z(n4702) );
  AND U4919 ( .A(n4703), .B(n4702), .Z(n4705) );
  NANDN U4920 ( .A(n5660), .B(\stack[5][25] ), .Z(n4704) );
  NAND U4921 ( .A(n4705), .B(n4704), .Z(n1121) );
  NAND U4922 ( .A(n5672), .B(\stack[3][25] ), .Z(n4707) );
  NANDN U4923 ( .A(n5657), .B(\stack[5][25] ), .Z(n4706) );
  AND U4924 ( .A(n4707), .B(n4706), .Z(n4709) );
  NANDN U4925 ( .A(n5660), .B(\stack[4][25] ), .Z(n4708) );
  NAND U4926 ( .A(n4709), .B(n4708), .Z(n1122) );
  NAND U4927 ( .A(n5672), .B(\stack[2][25] ), .Z(n4711) );
  NANDN U4928 ( .A(n5657), .B(\stack[4][25] ), .Z(n4710) );
  AND U4929 ( .A(n4711), .B(n4710), .Z(n4713) );
  NANDN U4930 ( .A(n5660), .B(\stack[3][25] ), .Z(n4712) );
  NAND U4931 ( .A(n4713), .B(n4712), .Z(n1123) );
  NAND U4932 ( .A(\stack[1][25] ), .B(n5672), .Z(n4715) );
  NANDN U4933 ( .A(n5657), .B(\stack[3][25] ), .Z(n4714) );
  AND U4934 ( .A(n4715), .B(n4714), .Z(n4717) );
  NANDN U4935 ( .A(n5660), .B(\stack[2][25] ), .Z(n4716) );
  NAND U4936 ( .A(n4717), .B(n4716), .Z(n1124) );
  NAND U4937 ( .A(o[25]), .B(n5672), .Z(n4719) );
  NANDN U4938 ( .A(n5657), .B(\stack[2][25] ), .Z(n4718) );
  AND U4939 ( .A(n4719), .B(n4718), .Z(n4721) );
  NANDN U4940 ( .A(n5660), .B(\stack[1][25] ), .Z(n4720) );
  NAND U4941 ( .A(n4721), .B(n4720), .Z(n1125) );
  XNOR U4942 ( .A(n4723), .B(n4722), .Z(n4724) );
  NAND U4943 ( .A(n4724), .B(n5644), .Z(n4728) );
  NAND U4944 ( .A(n5672), .B(x[25]), .Z(n4726) );
  NAND U4945 ( .A(n5651), .B(\stack[1][25] ), .Z(n4725) );
  AND U4946 ( .A(n4726), .B(n4725), .Z(n4727) );
  NAND U4947 ( .A(n4728), .B(n4727), .Z(n4733) );
  NAND U4948 ( .A(\stack[1][25] ), .B(n5665), .Z(n4729) );
  NAND U4949 ( .A(n1604), .B(n4729), .Z(n4730) );
  AND U4950 ( .A(n4730), .B(o[25]), .Z(n4731) );
  NANDN U4951 ( .A(n4733), .B(n4732), .Z(n1126) );
  NAND U4952 ( .A(n5672), .B(\stack[6][24] ), .Z(n4735) );
  NAND U4953 ( .A(n1605), .B(\stack[7][24] ), .Z(n4734) );
  NAND U4954 ( .A(n4735), .B(n4734), .Z(n1127) );
  NAND U4955 ( .A(n5672), .B(\stack[5][24] ), .Z(n4737) );
  NANDN U4956 ( .A(n5657), .B(\stack[7][24] ), .Z(n4736) );
  AND U4957 ( .A(n4737), .B(n4736), .Z(n4739) );
  NANDN U4958 ( .A(n5660), .B(\stack[6][24] ), .Z(n4738) );
  NAND U4959 ( .A(n4739), .B(n4738), .Z(n1128) );
  NAND U4960 ( .A(n5672), .B(\stack[4][24] ), .Z(n4741) );
  NANDN U4961 ( .A(n5657), .B(\stack[6][24] ), .Z(n4740) );
  AND U4962 ( .A(n4741), .B(n4740), .Z(n4743) );
  NANDN U4963 ( .A(n5660), .B(\stack[5][24] ), .Z(n4742) );
  NAND U4964 ( .A(n4743), .B(n4742), .Z(n1129) );
  NAND U4965 ( .A(n5672), .B(\stack[3][24] ), .Z(n4745) );
  NANDN U4966 ( .A(n5657), .B(\stack[5][24] ), .Z(n4744) );
  AND U4967 ( .A(n4745), .B(n4744), .Z(n4747) );
  NANDN U4968 ( .A(n5660), .B(\stack[4][24] ), .Z(n4746) );
  NAND U4969 ( .A(n4747), .B(n4746), .Z(n1130) );
  NAND U4970 ( .A(n5672), .B(\stack[2][24] ), .Z(n4749) );
  NANDN U4971 ( .A(n5657), .B(\stack[4][24] ), .Z(n4748) );
  AND U4972 ( .A(n4749), .B(n4748), .Z(n4751) );
  NANDN U4973 ( .A(n5660), .B(\stack[3][24] ), .Z(n4750) );
  NAND U4974 ( .A(n4751), .B(n4750), .Z(n1131) );
  NAND U4975 ( .A(\stack[1][24] ), .B(n5672), .Z(n4753) );
  NANDN U4976 ( .A(n5657), .B(\stack[3][24] ), .Z(n4752) );
  AND U4977 ( .A(n4753), .B(n4752), .Z(n4755) );
  NANDN U4978 ( .A(n5660), .B(\stack[2][24] ), .Z(n4754) );
  NAND U4979 ( .A(n4755), .B(n4754), .Z(n1132) );
  NAND U4980 ( .A(o[24]), .B(n5672), .Z(n4757) );
  NANDN U4981 ( .A(n5657), .B(\stack[2][24] ), .Z(n4756) );
  AND U4982 ( .A(n4757), .B(n4756), .Z(n4759) );
  NANDN U4983 ( .A(n5660), .B(\stack[1][24] ), .Z(n4758) );
  NAND U4984 ( .A(n4759), .B(n4758), .Z(n1133) );
  XNOR U4985 ( .A(n4761), .B(n4760), .Z(n4762) );
  NAND U4986 ( .A(n4762), .B(n5644), .Z(n4765) );
  NAND U4987 ( .A(n5672), .B(x[24]), .Z(n4763) );
  NAND U4988 ( .A(n4765), .B(n4764), .Z(n4771) );
  NAND U4989 ( .A(n5663), .B(o[24]), .Z(n4769) );
  NAND U4990 ( .A(o[24]), .B(n5665), .Z(n4766) );
  NAND U4991 ( .A(n5667), .B(n4766), .Z(n4767) );
  AND U4992 ( .A(n4767), .B(\stack[1][24] ), .Z(n4768) );
  ANDN U4993 ( .B(n4769), .A(n4768), .Z(n4770) );
  NANDN U4994 ( .A(n4771), .B(n4770), .Z(n1134) );
  NAND U4995 ( .A(n5672), .B(\stack[6][23] ), .Z(n4773) );
  NAND U4996 ( .A(n1605), .B(\stack[7][23] ), .Z(n4772) );
  NAND U4997 ( .A(n4773), .B(n4772), .Z(n1135) );
  NAND U4998 ( .A(n5672), .B(\stack[5][23] ), .Z(n4775) );
  NANDN U4999 ( .A(n5657), .B(\stack[7][23] ), .Z(n4774) );
  AND U5000 ( .A(n4775), .B(n4774), .Z(n4777) );
  NANDN U5001 ( .A(n5660), .B(\stack[6][23] ), .Z(n4776) );
  NAND U5002 ( .A(n4777), .B(n4776), .Z(n1136) );
  NAND U5003 ( .A(n5672), .B(\stack[4][23] ), .Z(n4779) );
  NANDN U5004 ( .A(n5657), .B(\stack[6][23] ), .Z(n4778) );
  AND U5005 ( .A(n4779), .B(n4778), .Z(n4781) );
  NANDN U5006 ( .A(n5660), .B(\stack[5][23] ), .Z(n4780) );
  NAND U5007 ( .A(n4781), .B(n4780), .Z(n1137) );
  NAND U5008 ( .A(n5672), .B(\stack[3][23] ), .Z(n4783) );
  NANDN U5009 ( .A(n5657), .B(\stack[5][23] ), .Z(n4782) );
  AND U5010 ( .A(n4783), .B(n4782), .Z(n4785) );
  NANDN U5011 ( .A(n5660), .B(\stack[4][23] ), .Z(n4784) );
  NAND U5012 ( .A(n4785), .B(n4784), .Z(n1138) );
  NAND U5013 ( .A(n5672), .B(\stack[2][23] ), .Z(n4787) );
  NANDN U5014 ( .A(n5657), .B(\stack[4][23] ), .Z(n4786) );
  AND U5015 ( .A(n4787), .B(n4786), .Z(n4789) );
  NANDN U5016 ( .A(n5660), .B(\stack[3][23] ), .Z(n4788) );
  NAND U5017 ( .A(n4789), .B(n4788), .Z(n1139) );
  NAND U5018 ( .A(\stack[1][23] ), .B(n5672), .Z(n4791) );
  NANDN U5019 ( .A(n5657), .B(\stack[3][23] ), .Z(n4790) );
  AND U5020 ( .A(n4791), .B(n4790), .Z(n4793) );
  NANDN U5021 ( .A(n5660), .B(\stack[2][23] ), .Z(n4792) );
  NAND U5022 ( .A(n4793), .B(n4792), .Z(n1140) );
  NAND U5023 ( .A(o[23]), .B(n5672), .Z(n4795) );
  NANDN U5024 ( .A(n5657), .B(\stack[2][23] ), .Z(n4794) );
  AND U5025 ( .A(n4795), .B(n4794), .Z(n4797) );
  NANDN U5026 ( .A(n5660), .B(\stack[1][23] ), .Z(n4796) );
  NAND U5027 ( .A(n4797), .B(n4796), .Z(n1141) );
  XNOR U5028 ( .A(n4799), .B(n4798), .Z(n4800) );
  NAND U5029 ( .A(n4800), .B(n5644), .Z(n4804) );
  NAND U5030 ( .A(n5672), .B(x[23]), .Z(n4802) );
  NAND U5031 ( .A(n5651), .B(\stack[1][23] ), .Z(n4801) );
  AND U5032 ( .A(n4802), .B(n4801), .Z(n4803) );
  NAND U5033 ( .A(n4804), .B(n4803), .Z(n4809) );
  NAND U5034 ( .A(\stack[1][23] ), .B(n5665), .Z(n4805) );
  NAND U5035 ( .A(n1604), .B(n4805), .Z(n4806) );
  AND U5036 ( .A(n4806), .B(o[23]), .Z(n4807) );
  NANDN U5037 ( .A(n4809), .B(n4808), .Z(n1142) );
  NAND U5038 ( .A(n5672), .B(\stack[6][22] ), .Z(n4811) );
  NAND U5039 ( .A(n1605), .B(\stack[7][22] ), .Z(n4810) );
  NAND U5040 ( .A(n4811), .B(n4810), .Z(n1143) );
  NAND U5041 ( .A(n5672), .B(\stack[5][22] ), .Z(n4813) );
  NANDN U5042 ( .A(n5657), .B(\stack[7][22] ), .Z(n4812) );
  AND U5043 ( .A(n4813), .B(n4812), .Z(n4815) );
  NANDN U5044 ( .A(n5660), .B(\stack[6][22] ), .Z(n4814) );
  NAND U5045 ( .A(n4815), .B(n4814), .Z(n1144) );
  NAND U5046 ( .A(n5672), .B(\stack[4][22] ), .Z(n4817) );
  NANDN U5047 ( .A(n5657), .B(\stack[6][22] ), .Z(n4816) );
  AND U5048 ( .A(n4817), .B(n4816), .Z(n4819) );
  NANDN U5049 ( .A(n5660), .B(\stack[5][22] ), .Z(n4818) );
  NAND U5050 ( .A(n4819), .B(n4818), .Z(n1145) );
  NAND U5051 ( .A(n5672), .B(\stack[3][22] ), .Z(n4821) );
  NANDN U5052 ( .A(n5657), .B(\stack[5][22] ), .Z(n4820) );
  AND U5053 ( .A(n4821), .B(n4820), .Z(n4823) );
  NANDN U5054 ( .A(n5660), .B(\stack[4][22] ), .Z(n4822) );
  NAND U5055 ( .A(n4823), .B(n4822), .Z(n1146) );
  NAND U5056 ( .A(n5672), .B(\stack[2][22] ), .Z(n4825) );
  NANDN U5057 ( .A(n5657), .B(\stack[4][22] ), .Z(n4824) );
  AND U5058 ( .A(n4825), .B(n4824), .Z(n4827) );
  NANDN U5059 ( .A(n5660), .B(\stack[3][22] ), .Z(n4826) );
  NAND U5060 ( .A(n4827), .B(n4826), .Z(n1147) );
  NAND U5061 ( .A(\stack[1][22] ), .B(n5672), .Z(n4829) );
  NANDN U5062 ( .A(n5657), .B(\stack[3][22] ), .Z(n4828) );
  AND U5063 ( .A(n4829), .B(n4828), .Z(n4831) );
  NANDN U5064 ( .A(n5660), .B(\stack[2][22] ), .Z(n4830) );
  NAND U5065 ( .A(n4831), .B(n4830), .Z(n1148) );
  NAND U5066 ( .A(o[22]), .B(n5672), .Z(n4833) );
  NANDN U5067 ( .A(n5657), .B(\stack[2][22] ), .Z(n4832) );
  AND U5068 ( .A(n4833), .B(n4832), .Z(n4835) );
  NANDN U5069 ( .A(n5660), .B(\stack[1][22] ), .Z(n4834) );
  NAND U5070 ( .A(n4835), .B(n4834), .Z(n1149) );
  XNOR U5071 ( .A(n4837), .B(n4836), .Z(n4838) );
  NAND U5072 ( .A(n4838), .B(n5644), .Z(n4841) );
  NAND U5073 ( .A(n5672), .B(x[22]), .Z(n4839) );
  NAND U5074 ( .A(n4841), .B(n4840), .Z(n4847) );
  NAND U5075 ( .A(n5663), .B(o[22]), .Z(n4845) );
  NAND U5076 ( .A(o[22]), .B(n5665), .Z(n4842) );
  NAND U5077 ( .A(n5667), .B(n4842), .Z(n4843) );
  AND U5078 ( .A(n4843), .B(\stack[1][22] ), .Z(n4844) );
  ANDN U5079 ( .B(n4845), .A(n4844), .Z(n4846) );
  NANDN U5080 ( .A(n4847), .B(n4846), .Z(n1150) );
  NAND U5081 ( .A(n5672), .B(\stack[6][21] ), .Z(n4849) );
  NAND U5082 ( .A(n1605), .B(\stack[7][21] ), .Z(n4848) );
  NAND U5083 ( .A(n4849), .B(n4848), .Z(n1151) );
  NAND U5084 ( .A(n5672), .B(\stack[5][21] ), .Z(n4851) );
  NANDN U5085 ( .A(n5657), .B(\stack[7][21] ), .Z(n4850) );
  AND U5086 ( .A(n4851), .B(n4850), .Z(n4853) );
  NANDN U5087 ( .A(n5660), .B(\stack[6][21] ), .Z(n4852) );
  NAND U5088 ( .A(n4853), .B(n4852), .Z(n1152) );
  NAND U5089 ( .A(n5672), .B(\stack[4][21] ), .Z(n4855) );
  NANDN U5090 ( .A(n5657), .B(\stack[6][21] ), .Z(n4854) );
  AND U5091 ( .A(n4855), .B(n4854), .Z(n4857) );
  NANDN U5092 ( .A(n5660), .B(\stack[5][21] ), .Z(n4856) );
  NAND U5093 ( .A(n4857), .B(n4856), .Z(n1153) );
  NAND U5094 ( .A(n5672), .B(\stack[3][21] ), .Z(n4859) );
  NANDN U5095 ( .A(n5657), .B(\stack[5][21] ), .Z(n4858) );
  AND U5096 ( .A(n4859), .B(n4858), .Z(n4861) );
  NANDN U5097 ( .A(n5660), .B(\stack[4][21] ), .Z(n4860) );
  NAND U5098 ( .A(n4861), .B(n4860), .Z(n1154) );
  NAND U5099 ( .A(n5672), .B(\stack[2][21] ), .Z(n4863) );
  NANDN U5100 ( .A(n5657), .B(\stack[4][21] ), .Z(n4862) );
  AND U5101 ( .A(n4863), .B(n4862), .Z(n4865) );
  NANDN U5102 ( .A(n5660), .B(\stack[3][21] ), .Z(n4864) );
  NAND U5103 ( .A(n4865), .B(n4864), .Z(n1155) );
  NAND U5104 ( .A(\stack[1][21] ), .B(n5672), .Z(n4867) );
  NANDN U5105 ( .A(n5657), .B(\stack[3][21] ), .Z(n4866) );
  AND U5106 ( .A(n4867), .B(n4866), .Z(n4869) );
  NANDN U5107 ( .A(n5660), .B(\stack[2][21] ), .Z(n4868) );
  NAND U5108 ( .A(n4869), .B(n4868), .Z(n1156) );
  NAND U5109 ( .A(o[21]), .B(n5672), .Z(n4871) );
  NANDN U5110 ( .A(n5657), .B(\stack[2][21] ), .Z(n4870) );
  AND U5111 ( .A(n4871), .B(n4870), .Z(n4873) );
  NANDN U5112 ( .A(n5660), .B(\stack[1][21] ), .Z(n4872) );
  NAND U5113 ( .A(n4873), .B(n4872), .Z(n1157) );
  XNOR U5114 ( .A(n4875), .B(n4874), .Z(n4876) );
  NAND U5115 ( .A(n4876), .B(n5644), .Z(n4880) );
  NAND U5116 ( .A(n5672), .B(x[21]), .Z(n4878) );
  NAND U5117 ( .A(n5651), .B(\stack[1][21] ), .Z(n4877) );
  AND U5118 ( .A(n4878), .B(n4877), .Z(n4879) );
  NAND U5119 ( .A(n4880), .B(n4879), .Z(n4885) );
  NAND U5120 ( .A(\stack[1][21] ), .B(n5665), .Z(n4881) );
  NAND U5121 ( .A(n1604), .B(n4881), .Z(n4882) );
  AND U5122 ( .A(n4882), .B(o[21]), .Z(n4883) );
  NANDN U5123 ( .A(n4885), .B(n4884), .Z(n1158) );
  NAND U5124 ( .A(n5672), .B(\stack[6][20] ), .Z(n4887) );
  NAND U5125 ( .A(n1605), .B(\stack[7][20] ), .Z(n4886) );
  NAND U5126 ( .A(n4887), .B(n4886), .Z(n1159) );
  NAND U5127 ( .A(n5672), .B(\stack[5][20] ), .Z(n4889) );
  NANDN U5128 ( .A(n5657), .B(\stack[7][20] ), .Z(n4888) );
  AND U5129 ( .A(n4889), .B(n4888), .Z(n4891) );
  NANDN U5130 ( .A(n5660), .B(\stack[6][20] ), .Z(n4890) );
  NAND U5131 ( .A(n4891), .B(n4890), .Z(n1160) );
  NAND U5132 ( .A(n5672), .B(\stack[4][20] ), .Z(n4893) );
  NANDN U5133 ( .A(n5657), .B(\stack[6][20] ), .Z(n4892) );
  AND U5134 ( .A(n4893), .B(n4892), .Z(n4895) );
  NANDN U5135 ( .A(n5660), .B(\stack[5][20] ), .Z(n4894) );
  NAND U5136 ( .A(n4895), .B(n4894), .Z(n1161) );
  NAND U5137 ( .A(n5672), .B(\stack[3][20] ), .Z(n4897) );
  NANDN U5138 ( .A(n5657), .B(\stack[5][20] ), .Z(n4896) );
  AND U5139 ( .A(n4897), .B(n4896), .Z(n4899) );
  NANDN U5140 ( .A(n5660), .B(\stack[4][20] ), .Z(n4898) );
  NAND U5141 ( .A(n4899), .B(n4898), .Z(n1162) );
  NAND U5142 ( .A(n5672), .B(\stack[2][20] ), .Z(n4901) );
  NANDN U5143 ( .A(n5657), .B(\stack[4][20] ), .Z(n4900) );
  AND U5144 ( .A(n4901), .B(n4900), .Z(n4903) );
  NANDN U5145 ( .A(n5660), .B(\stack[3][20] ), .Z(n4902) );
  NAND U5146 ( .A(n4903), .B(n4902), .Z(n1163) );
  NAND U5147 ( .A(\stack[1][20] ), .B(n5672), .Z(n4905) );
  NANDN U5148 ( .A(n5657), .B(\stack[3][20] ), .Z(n4904) );
  AND U5149 ( .A(n4905), .B(n4904), .Z(n4907) );
  NANDN U5150 ( .A(n5660), .B(\stack[2][20] ), .Z(n4906) );
  NAND U5151 ( .A(n4907), .B(n4906), .Z(n1164) );
  NAND U5152 ( .A(o[20]), .B(n5672), .Z(n4909) );
  NANDN U5153 ( .A(n5657), .B(\stack[2][20] ), .Z(n4908) );
  AND U5154 ( .A(n4909), .B(n4908), .Z(n4911) );
  NANDN U5155 ( .A(n5660), .B(\stack[1][20] ), .Z(n4910) );
  NAND U5156 ( .A(n4911), .B(n4910), .Z(n1165) );
  XNOR U5157 ( .A(n4913), .B(n4912), .Z(n4914) );
  NAND U5158 ( .A(n4914), .B(n5644), .Z(n4917) );
  NAND U5159 ( .A(n5672), .B(x[20]), .Z(n4915) );
  NAND U5160 ( .A(n4917), .B(n4916), .Z(n4923) );
  NAND U5161 ( .A(n5663), .B(o[20]), .Z(n4921) );
  NAND U5162 ( .A(o[20]), .B(n5665), .Z(n4918) );
  NAND U5163 ( .A(n5667), .B(n4918), .Z(n4919) );
  AND U5164 ( .A(n4919), .B(\stack[1][20] ), .Z(n4920) );
  ANDN U5165 ( .B(n4921), .A(n4920), .Z(n4922) );
  NANDN U5166 ( .A(n4923), .B(n4922), .Z(n1166) );
  NAND U5167 ( .A(n5672), .B(\stack[6][19] ), .Z(n4925) );
  NAND U5168 ( .A(n1605), .B(\stack[7][19] ), .Z(n4924) );
  NAND U5169 ( .A(n4925), .B(n4924), .Z(n1167) );
  NAND U5170 ( .A(n5672), .B(\stack[5][19] ), .Z(n4927) );
  NANDN U5171 ( .A(n5657), .B(\stack[7][19] ), .Z(n4926) );
  AND U5172 ( .A(n4927), .B(n4926), .Z(n4929) );
  NANDN U5173 ( .A(n5660), .B(\stack[6][19] ), .Z(n4928) );
  NAND U5174 ( .A(n4929), .B(n4928), .Z(n1168) );
  NAND U5175 ( .A(n5672), .B(\stack[4][19] ), .Z(n4931) );
  NANDN U5176 ( .A(n5657), .B(\stack[6][19] ), .Z(n4930) );
  AND U5177 ( .A(n4931), .B(n4930), .Z(n4933) );
  NANDN U5178 ( .A(n5660), .B(\stack[5][19] ), .Z(n4932) );
  NAND U5179 ( .A(n4933), .B(n4932), .Z(n1169) );
  NAND U5180 ( .A(n5672), .B(\stack[3][19] ), .Z(n4935) );
  NANDN U5181 ( .A(n5657), .B(\stack[5][19] ), .Z(n4934) );
  AND U5182 ( .A(n4935), .B(n4934), .Z(n4937) );
  NANDN U5183 ( .A(n5660), .B(\stack[4][19] ), .Z(n4936) );
  NAND U5184 ( .A(n4937), .B(n4936), .Z(n1170) );
  NAND U5185 ( .A(n5672), .B(\stack[2][19] ), .Z(n4939) );
  NANDN U5186 ( .A(n5657), .B(\stack[4][19] ), .Z(n4938) );
  AND U5187 ( .A(n4939), .B(n4938), .Z(n4941) );
  NANDN U5188 ( .A(n5660), .B(\stack[3][19] ), .Z(n4940) );
  NAND U5189 ( .A(n4941), .B(n4940), .Z(n1171) );
  NAND U5190 ( .A(\stack[1][19] ), .B(n5672), .Z(n4943) );
  NANDN U5191 ( .A(n5657), .B(\stack[3][19] ), .Z(n4942) );
  AND U5192 ( .A(n4943), .B(n4942), .Z(n4945) );
  NANDN U5193 ( .A(n5660), .B(\stack[2][19] ), .Z(n4944) );
  NAND U5194 ( .A(n4945), .B(n4944), .Z(n1172) );
  NAND U5195 ( .A(o[19]), .B(n5672), .Z(n4947) );
  NANDN U5196 ( .A(n5657), .B(\stack[2][19] ), .Z(n4946) );
  AND U5197 ( .A(n4947), .B(n4946), .Z(n4949) );
  NANDN U5198 ( .A(n5660), .B(\stack[1][19] ), .Z(n4948) );
  NAND U5199 ( .A(n4949), .B(n4948), .Z(n1173) );
  XNOR U5200 ( .A(n4951), .B(n4950), .Z(n4952) );
  NAND U5201 ( .A(n4952), .B(n5644), .Z(n4956) );
  NAND U5202 ( .A(n5672), .B(x[19]), .Z(n4954) );
  NAND U5203 ( .A(n5651), .B(\stack[1][19] ), .Z(n4953) );
  AND U5204 ( .A(n4954), .B(n4953), .Z(n4955) );
  NAND U5205 ( .A(n4956), .B(n4955), .Z(n4961) );
  NAND U5206 ( .A(\stack[1][19] ), .B(n5665), .Z(n4957) );
  NAND U5207 ( .A(n1604), .B(n4957), .Z(n4958) );
  AND U5208 ( .A(n4958), .B(o[19]), .Z(n4959) );
  NANDN U5209 ( .A(n4961), .B(n4960), .Z(n1174) );
  NAND U5210 ( .A(n5672), .B(\stack[6][18] ), .Z(n4963) );
  NAND U5211 ( .A(n1605), .B(\stack[7][18] ), .Z(n4962) );
  NAND U5212 ( .A(n4963), .B(n4962), .Z(n1175) );
  NAND U5213 ( .A(n5672), .B(\stack[5][18] ), .Z(n4965) );
  NANDN U5214 ( .A(n5657), .B(\stack[7][18] ), .Z(n4964) );
  AND U5215 ( .A(n4965), .B(n4964), .Z(n4967) );
  NANDN U5216 ( .A(n5660), .B(\stack[6][18] ), .Z(n4966) );
  NAND U5217 ( .A(n4967), .B(n4966), .Z(n1176) );
  NAND U5218 ( .A(n5672), .B(\stack[4][18] ), .Z(n4969) );
  NANDN U5219 ( .A(n5657), .B(\stack[6][18] ), .Z(n4968) );
  AND U5220 ( .A(n4969), .B(n4968), .Z(n4971) );
  NANDN U5221 ( .A(n5660), .B(\stack[5][18] ), .Z(n4970) );
  NAND U5222 ( .A(n4971), .B(n4970), .Z(n1177) );
  NAND U5223 ( .A(n5672), .B(\stack[3][18] ), .Z(n4973) );
  NANDN U5224 ( .A(n5657), .B(\stack[5][18] ), .Z(n4972) );
  AND U5225 ( .A(n4973), .B(n4972), .Z(n4975) );
  NANDN U5226 ( .A(n5660), .B(\stack[4][18] ), .Z(n4974) );
  NAND U5227 ( .A(n4975), .B(n4974), .Z(n1178) );
  NAND U5228 ( .A(n5672), .B(\stack[2][18] ), .Z(n4977) );
  NANDN U5229 ( .A(n5657), .B(\stack[4][18] ), .Z(n4976) );
  AND U5230 ( .A(n4977), .B(n4976), .Z(n4979) );
  NANDN U5231 ( .A(n5660), .B(\stack[3][18] ), .Z(n4978) );
  NAND U5232 ( .A(n4979), .B(n4978), .Z(n1179) );
  NAND U5233 ( .A(\stack[1][18] ), .B(n5672), .Z(n4981) );
  NANDN U5234 ( .A(n5657), .B(\stack[3][18] ), .Z(n4980) );
  AND U5235 ( .A(n4981), .B(n4980), .Z(n4983) );
  NANDN U5236 ( .A(n5660), .B(\stack[2][18] ), .Z(n4982) );
  NAND U5237 ( .A(n4983), .B(n4982), .Z(n1180) );
  NAND U5238 ( .A(o[18]), .B(n5672), .Z(n4985) );
  NANDN U5239 ( .A(n5657), .B(\stack[2][18] ), .Z(n4984) );
  AND U5240 ( .A(n4985), .B(n4984), .Z(n4987) );
  NANDN U5241 ( .A(n5660), .B(\stack[1][18] ), .Z(n4986) );
  NAND U5242 ( .A(n4987), .B(n4986), .Z(n1181) );
  XNOR U5243 ( .A(n4989), .B(n4988), .Z(n4990) );
  NAND U5244 ( .A(n4990), .B(n5644), .Z(n4993) );
  NAND U5245 ( .A(n5672), .B(x[18]), .Z(n4991) );
  NAND U5246 ( .A(n4993), .B(n4992), .Z(n4999) );
  NAND U5247 ( .A(n5663), .B(o[18]), .Z(n4997) );
  NAND U5248 ( .A(o[18]), .B(n5665), .Z(n4994) );
  NAND U5249 ( .A(n5667), .B(n4994), .Z(n4995) );
  AND U5250 ( .A(n4995), .B(\stack[1][18] ), .Z(n4996) );
  ANDN U5251 ( .B(n4997), .A(n4996), .Z(n4998) );
  NANDN U5252 ( .A(n4999), .B(n4998), .Z(n1182) );
  NAND U5253 ( .A(n5672), .B(\stack[6][17] ), .Z(n5001) );
  NAND U5254 ( .A(n1605), .B(\stack[7][17] ), .Z(n5000) );
  NAND U5255 ( .A(n5001), .B(n5000), .Z(n1183) );
  NAND U5256 ( .A(n5672), .B(\stack[5][17] ), .Z(n5003) );
  NANDN U5257 ( .A(n5657), .B(\stack[7][17] ), .Z(n5002) );
  AND U5258 ( .A(n5003), .B(n5002), .Z(n5005) );
  NANDN U5259 ( .A(n5660), .B(\stack[6][17] ), .Z(n5004) );
  NAND U5260 ( .A(n5005), .B(n5004), .Z(n1184) );
  NAND U5261 ( .A(n5672), .B(\stack[4][17] ), .Z(n5007) );
  NANDN U5262 ( .A(n5657), .B(\stack[6][17] ), .Z(n5006) );
  AND U5263 ( .A(n5007), .B(n5006), .Z(n5009) );
  NANDN U5264 ( .A(n5660), .B(\stack[5][17] ), .Z(n5008) );
  NAND U5265 ( .A(n5009), .B(n5008), .Z(n1185) );
  NAND U5266 ( .A(n5672), .B(\stack[3][17] ), .Z(n5011) );
  NANDN U5267 ( .A(n5657), .B(\stack[5][17] ), .Z(n5010) );
  AND U5268 ( .A(n5011), .B(n5010), .Z(n5013) );
  NANDN U5269 ( .A(n5660), .B(\stack[4][17] ), .Z(n5012) );
  NAND U5270 ( .A(n5013), .B(n5012), .Z(n1186) );
  NAND U5271 ( .A(n5672), .B(\stack[2][17] ), .Z(n5015) );
  NANDN U5272 ( .A(n5657), .B(\stack[4][17] ), .Z(n5014) );
  AND U5273 ( .A(n5015), .B(n5014), .Z(n5017) );
  NANDN U5274 ( .A(n5660), .B(\stack[3][17] ), .Z(n5016) );
  NAND U5275 ( .A(n5017), .B(n5016), .Z(n1187) );
  NAND U5276 ( .A(\stack[1][17] ), .B(n5672), .Z(n5019) );
  NANDN U5277 ( .A(n5657), .B(\stack[3][17] ), .Z(n5018) );
  AND U5278 ( .A(n5019), .B(n5018), .Z(n5021) );
  NANDN U5279 ( .A(n5660), .B(\stack[2][17] ), .Z(n5020) );
  NAND U5280 ( .A(n5021), .B(n5020), .Z(n1188) );
  NAND U5281 ( .A(o[17]), .B(n5672), .Z(n5023) );
  NANDN U5282 ( .A(n5657), .B(\stack[2][17] ), .Z(n5022) );
  AND U5283 ( .A(n5023), .B(n5022), .Z(n5025) );
  NANDN U5284 ( .A(n5660), .B(\stack[1][17] ), .Z(n5024) );
  NAND U5285 ( .A(n5025), .B(n5024), .Z(n1189) );
  XNOR U5286 ( .A(n5027), .B(n5026), .Z(n5028) );
  NAND U5287 ( .A(n5028), .B(n5644), .Z(n5032) );
  NAND U5288 ( .A(n5672), .B(x[17]), .Z(n5030) );
  NAND U5289 ( .A(n5651), .B(\stack[1][17] ), .Z(n5029) );
  AND U5290 ( .A(n5030), .B(n5029), .Z(n5031) );
  NAND U5291 ( .A(n5032), .B(n5031), .Z(n5037) );
  NAND U5292 ( .A(\stack[1][17] ), .B(n5665), .Z(n5033) );
  NAND U5293 ( .A(n1604), .B(n5033), .Z(n5034) );
  AND U5294 ( .A(n5034), .B(o[17]), .Z(n5035) );
  NANDN U5295 ( .A(n5037), .B(n5036), .Z(n1190) );
  NAND U5296 ( .A(n5672), .B(\stack[6][16] ), .Z(n5039) );
  NAND U5297 ( .A(n1605), .B(\stack[7][16] ), .Z(n5038) );
  NAND U5298 ( .A(n5039), .B(n5038), .Z(n1191) );
  NAND U5299 ( .A(n5672), .B(\stack[5][16] ), .Z(n5041) );
  NANDN U5300 ( .A(n5657), .B(\stack[7][16] ), .Z(n5040) );
  AND U5301 ( .A(n5041), .B(n5040), .Z(n5043) );
  NANDN U5302 ( .A(n5660), .B(\stack[6][16] ), .Z(n5042) );
  NAND U5303 ( .A(n5043), .B(n5042), .Z(n1192) );
  NAND U5304 ( .A(n5672), .B(\stack[4][16] ), .Z(n5045) );
  NANDN U5305 ( .A(n5657), .B(\stack[6][16] ), .Z(n5044) );
  AND U5306 ( .A(n5045), .B(n5044), .Z(n5047) );
  NANDN U5307 ( .A(n5660), .B(\stack[5][16] ), .Z(n5046) );
  NAND U5308 ( .A(n5047), .B(n5046), .Z(n1193) );
  NAND U5309 ( .A(n5672), .B(\stack[3][16] ), .Z(n5049) );
  NANDN U5310 ( .A(n5657), .B(\stack[5][16] ), .Z(n5048) );
  AND U5311 ( .A(n5049), .B(n5048), .Z(n5051) );
  NANDN U5312 ( .A(n5660), .B(\stack[4][16] ), .Z(n5050) );
  NAND U5313 ( .A(n5051), .B(n5050), .Z(n1194) );
  NAND U5314 ( .A(n5672), .B(\stack[2][16] ), .Z(n5053) );
  NANDN U5315 ( .A(n5657), .B(\stack[4][16] ), .Z(n5052) );
  AND U5316 ( .A(n5053), .B(n5052), .Z(n5055) );
  NANDN U5317 ( .A(n5660), .B(\stack[3][16] ), .Z(n5054) );
  NAND U5318 ( .A(n5055), .B(n5054), .Z(n1195) );
  NAND U5319 ( .A(\stack[1][16] ), .B(n5672), .Z(n5057) );
  NANDN U5320 ( .A(n5657), .B(\stack[3][16] ), .Z(n5056) );
  AND U5321 ( .A(n5057), .B(n5056), .Z(n5059) );
  NANDN U5322 ( .A(n5660), .B(\stack[2][16] ), .Z(n5058) );
  NAND U5323 ( .A(n5059), .B(n5058), .Z(n1196) );
  NAND U5324 ( .A(o[16]), .B(n5672), .Z(n5061) );
  NANDN U5325 ( .A(n5657), .B(\stack[2][16] ), .Z(n5060) );
  AND U5326 ( .A(n5061), .B(n5060), .Z(n5063) );
  NANDN U5327 ( .A(n5660), .B(\stack[1][16] ), .Z(n5062) );
  NAND U5328 ( .A(n5063), .B(n5062), .Z(n1197) );
  XNOR U5329 ( .A(n5065), .B(n5064), .Z(n5066) );
  NAND U5330 ( .A(n5066), .B(n5644), .Z(n5069) );
  NAND U5331 ( .A(n5672), .B(x[16]), .Z(n5067) );
  NAND U5332 ( .A(n5069), .B(n5068), .Z(n5075) );
  NAND U5333 ( .A(n5663), .B(o[16]), .Z(n5073) );
  NAND U5334 ( .A(o[16]), .B(n5665), .Z(n5070) );
  NAND U5335 ( .A(n5667), .B(n5070), .Z(n5071) );
  AND U5336 ( .A(n5071), .B(\stack[1][16] ), .Z(n5072) );
  ANDN U5337 ( .B(n5073), .A(n5072), .Z(n5074) );
  NANDN U5338 ( .A(n5075), .B(n5074), .Z(n1198) );
  NAND U5339 ( .A(n5672), .B(\stack[6][15] ), .Z(n5077) );
  NAND U5340 ( .A(n1605), .B(\stack[7][15] ), .Z(n5076) );
  NAND U5341 ( .A(n5077), .B(n5076), .Z(n1199) );
  NAND U5342 ( .A(n5672), .B(\stack[5][15] ), .Z(n5079) );
  NANDN U5343 ( .A(n5657), .B(\stack[7][15] ), .Z(n5078) );
  AND U5344 ( .A(n5079), .B(n5078), .Z(n5081) );
  NANDN U5345 ( .A(n5660), .B(\stack[6][15] ), .Z(n5080) );
  NAND U5346 ( .A(n5081), .B(n5080), .Z(n1200) );
  NAND U5347 ( .A(n5672), .B(\stack[4][15] ), .Z(n5083) );
  NANDN U5348 ( .A(n5657), .B(\stack[6][15] ), .Z(n5082) );
  AND U5349 ( .A(n5083), .B(n5082), .Z(n5085) );
  NANDN U5350 ( .A(n5660), .B(\stack[5][15] ), .Z(n5084) );
  NAND U5351 ( .A(n5085), .B(n5084), .Z(n1201) );
  NAND U5352 ( .A(n5672), .B(\stack[3][15] ), .Z(n5087) );
  NANDN U5353 ( .A(n5657), .B(\stack[5][15] ), .Z(n5086) );
  AND U5354 ( .A(n5087), .B(n5086), .Z(n5089) );
  NANDN U5355 ( .A(n5660), .B(\stack[4][15] ), .Z(n5088) );
  NAND U5356 ( .A(n5089), .B(n5088), .Z(n1202) );
  NAND U5357 ( .A(n5672), .B(\stack[2][15] ), .Z(n5091) );
  NANDN U5358 ( .A(n5657), .B(\stack[4][15] ), .Z(n5090) );
  AND U5359 ( .A(n5091), .B(n5090), .Z(n5093) );
  NANDN U5360 ( .A(n5660), .B(\stack[3][15] ), .Z(n5092) );
  NAND U5361 ( .A(n5093), .B(n5092), .Z(n1203) );
  NAND U5362 ( .A(\stack[1][15] ), .B(n5672), .Z(n5095) );
  NANDN U5363 ( .A(n5657), .B(\stack[3][15] ), .Z(n5094) );
  AND U5364 ( .A(n5095), .B(n5094), .Z(n5097) );
  NANDN U5365 ( .A(n5660), .B(\stack[2][15] ), .Z(n5096) );
  NAND U5366 ( .A(n5097), .B(n5096), .Z(n1204) );
  NAND U5367 ( .A(n5672), .B(o[15]), .Z(n5099) );
  NANDN U5368 ( .A(n5657), .B(\stack[2][15] ), .Z(n5098) );
  AND U5369 ( .A(n5099), .B(n5098), .Z(n5101) );
  NANDN U5370 ( .A(n5660), .B(\stack[1][15] ), .Z(n5100) );
  NAND U5371 ( .A(n5101), .B(n5100), .Z(n1205) );
  NAND U5372 ( .A(n5102), .B(n5665), .Z(n5103) );
  XNOR U5373 ( .A(n5105), .B(n5104), .Z(n5106) );
  NAND U5374 ( .A(n5106), .B(n5644), .Z(n5107) );
  NANDN U5375 ( .A(n5108), .B(n5107), .Z(n5114) );
  NAND U5376 ( .A(n5663), .B(o[15]), .Z(n5112) );
  NAND U5377 ( .A(n5672), .B(x[15]), .Z(n5110) );
  NAND U5378 ( .A(n5651), .B(\stack[1][15] ), .Z(n5109) );
  NAND U5379 ( .A(n5110), .B(n5109), .Z(n5111) );
  ANDN U5380 ( .B(n5112), .A(n5111), .Z(n5113) );
  NANDN U5381 ( .A(n5114), .B(n5113), .Z(n1206) );
  NAND U5382 ( .A(n5672), .B(\stack[6][14] ), .Z(n5116) );
  NAND U5383 ( .A(n1605), .B(\stack[7][14] ), .Z(n5115) );
  NAND U5384 ( .A(n5116), .B(n5115), .Z(n1207) );
  NAND U5385 ( .A(n5672), .B(\stack[5][14] ), .Z(n5118) );
  NANDN U5386 ( .A(n5657), .B(\stack[7][14] ), .Z(n5117) );
  AND U5387 ( .A(n5118), .B(n5117), .Z(n5120) );
  NANDN U5388 ( .A(n5660), .B(\stack[6][14] ), .Z(n5119) );
  NAND U5389 ( .A(n5120), .B(n5119), .Z(n1208) );
  NAND U5390 ( .A(n5672), .B(\stack[4][14] ), .Z(n5122) );
  NANDN U5391 ( .A(n5657), .B(\stack[6][14] ), .Z(n5121) );
  AND U5392 ( .A(n5122), .B(n5121), .Z(n5124) );
  NANDN U5393 ( .A(n5660), .B(\stack[5][14] ), .Z(n5123) );
  NAND U5394 ( .A(n5124), .B(n5123), .Z(n1209) );
  NAND U5395 ( .A(n5672), .B(\stack[3][14] ), .Z(n5126) );
  NANDN U5396 ( .A(n5657), .B(\stack[5][14] ), .Z(n5125) );
  AND U5397 ( .A(n5126), .B(n5125), .Z(n5128) );
  NANDN U5398 ( .A(n5660), .B(\stack[4][14] ), .Z(n5127) );
  NAND U5399 ( .A(n5128), .B(n5127), .Z(n1210) );
  NAND U5400 ( .A(n5672), .B(\stack[2][14] ), .Z(n5130) );
  NANDN U5401 ( .A(n5657), .B(\stack[4][14] ), .Z(n5129) );
  AND U5402 ( .A(n5130), .B(n5129), .Z(n5132) );
  NANDN U5403 ( .A(n5660), .B(\stack[3][14] ), .Z(n5131) );
  NAND U5404 ( .A(n5132), .B(n5131), .Z(n1211) );
  NAND U5405 ( .A(\stack[1][14] ), .B(n5672), .Z(n5134) );
  NANDN U5406 ( .A(n5657), .B(\stack[3][14] ), .Z(n5133) );
  AND U5407 ( .A(n5134), .B(n5133), .Z(n5136) );
  NANDN U5408 ( .A(n5660), .B(\stack[2][14] ), .Z(n5135) );
  NAND U5409 ( .A(n5136), .B(n5135), .Z(n1212) );
  NAND U5410 ( .A(n5672), .B(o[14]), .Z(n5138) );
  NANDN U5411 ( .A(n5657), .B(\stack[2][14] ), .Z(n5137) );
  AND U5412 ( .A(n5138), .B(n5137), .Z(n5140) );
  NANDN U5413 ( .A(n5660), .B(\stack[1][14] ), .Z(n5139) );
  NAND U5414 ( .A(n5140), .B(n5139), .Z(n1213) );
  XNOR U5415 ( .A(n5142), .B(n5141), .Z(n5143) );
  NAND U5416 ( .A(n5143), .B(n5644), .Z(n5146) );
  NAND U5417 ( .A(\stack[1][14] ), .B(n5651), .Z(n5144) );
  NAND U5418 ( .A(n5146), .B(n5145), .Z(n5153) );
  NAND U5419 ( .A(n5663), .B(o[14]), .Z(n5151) );
  NAND U5420 ( .A(n5672), .B(x[14]), .Z(n5149) );
  NAND U5421 ( .A(n5147), .B(n5665), .Z(n5148) );
  NAND U5422 ( .A(n5149), .B(n5148), .Z(n5150) );
  ANDN U5423 ( .B(n5151), .A(n5150), .Z(n5152) );
  NANDN U5424 ( .A(n5153), .B(n5152), .Z(n1214) );
  NAND U5425 ( .A(n5672), .B(\stack[6][13] ), .Z(n5155) );
  NAND U5426 ( .A(n1605), .B(\stack[7][13] ), .Z(n5154) );
  NAND U5427 ( .A(n5155), .B(n5154), .Z(n1215) );
  NAND U5428 ( .A(n5672), .B(\stack[5][13] ), .Z(n5157) );
  NANDN U5429 ( .A(n5657), .B(\stack[7][13] ), .Z(n5156) );
  AND U5430 ( .A(n5157), .B(n5156), .Z(n5159) );
  NANDN U5431 ( .A(n5660), .B(\stack[6][13] ), .Z(n5158) );
  NAND U5432 ( .A(n5159), .B(n5158), .Z(n1216) );
  NAND U5433 ( .A(n5672), .B(\stack[4][13] ), .Z(n5161) );
  NANDN U5434 ( .A(n5657), .B(\stack[6][13] ), .Z(n5160) );
  AND U5435 ( .A(n5161), .B(n5160), .Z(n5163) );
  NANDN U5436 ( .A(n5660), .B(\stack[5][13] ), .Z(n5162) );
  NAND U5437 ( .A(n5163), .B(n5162), .Z(n1217) );
  NAND U5438 ( .A(n5672), .B(\stack[3][13] ), .Z(n5165) );
  NANDN U5439 ( .A(n5657), .B(\stack[5][13] ), .Z(n5164) );
  AND U5440 ( .A(n5165), .B(n5164), .Z(n5167) );
  NANDN U5441 ( .A(n5660), .B(\stack[4][13] ), .Z(n5166) );
  NAND U5442 ( .A(n5167), .B(n5166), .Z(n1218) );
  NAND U5443 ( .A(n5672), .B(\stack[2][13] ), .Z(n5169) );
  NANDN U5444 ( .A(n5657), .B(\stack[4][13] ), .Z(n5168) );
  AND U5445 ( .A(n5169), .B(n5168), .Z(n5171) );
  NANDN U5446 ( .A(n5660), .B(\stack[3][13] ), .Z(n5170) );
  NAND U5447 ( .A(n5171), .B(n5170), .Z(n1219) );
  NAND U5448 ( .A(\stack[1][13] ), .B(n5672), .Z(n5173) );
  NANDN U5449 ( .A(n5657), .B(\stack[3][13] ), .Z(n5172) );
  AND U5450 ( .A(n5173), .B(n5172), .Z(n5175) );
  NANDN U5451 ( .A(n5660), .B(\stack[2][13] ), .Z(n5174) );
  NAND U5452 ( .A(n5175), .B(n5174), .Z(n1220) );
  NAND U5453 ( .A(o[13]), .B(n5672), .Z(n5177) );
  NANDN U5454 ( .A(n5657), .B(\stack[2][13] ), .Z(n5176) );
  AND U5455 ( .A(n5177), .B(n5176), .Z(n5179) );
  NANDN U5456 ( .A(n5660), .B(\stack[1][13] ), .Z(n5178) );
  NAND U5457 ( .A(n5179), .B(n5178), .Z(n1221) );
  XNOR U5458 ( .A(n5181), .B(n5180), .Z(n5182) );
  NAND U5459 ( .A(n5182), .B(n5644), .Z(n5185) );
  NAND U5460 ( .A(n5672), .B(x[13]), .Z(n5183) );
  NAND U5461 ( .A(n5185), .B(n5184), .Z(n5191) );
  NAND U5462 ( .A(n5663), .B(o[13]), .Z(n5189) );
  NAND U5463 ( .A(o[13]), .B(n5665), .Z(n5186) );
  NAND U5464 ( .A(n5667), .B(n5186), .Z(n5187) );
  AND U5465 ( .A(n5187), .B(\stack[1][13] ), .Z(n5188) );
  ANDN U5466 ( .B(n5189), .A(n5188), .Z(n5190) );
  NANDN U5467 ( .A(n5191), .B(n5190), .Z(n1222) );
  NAND U5468 ( .A(n5672), .B(\stack[6][12] ), .Z(n5193) );
  NAND U5469 ( .A(n1605), .B(\stack[7][12] ), .Z(n5192) );
  NAND U5470 ( .A(n5193), .B(n5192), .Z(n1223) );
  NAND U5471 ( .A(n5672), .B(\stack[5][12] ), .Z(n5195) );
  NANDN U5472 ( .A(n5657), .B(\stack[7][12] ), .Z(n5194) );
  AND U5473 ( .A(n5195), .B(n5194), .Z(n5197) );
  NANDN U5474 ( .A(n5660), .B(\stack[6][12] ), .Z(n5196) );
  NAND U5475 ( .A(n5197), .B(n5196), .Z(n1224) );
  NAND U5476 ( .A(n5672), .B(\stack[4][12] ), .Z(n5199) );
  NANDN U5477 ( .A(n5657), .B(\stack[6][12] ), .Z(n5198) );
  AND U5478 ( .A(n5199), .B(n5198), .Z(n5201) );
  NANDN U5479 ( .A(n5660), .B(\stack[5][12] ), .Z(n5200) );
  NAND U5480 ( .A(n5201), .B(n5200), .Z(n1225) );
  NAND U5481 ( .A(n5672), .B(\stack[3][12] ), .Z(n5203) );
  NANDN U5482 ( .A(n5657), .B(\stack[5][12] ), .Z(n5202) );
  AND U5483 ( .A(n5203), .B(n5202), .Z(n5205) );
  NANDN U5484 ( .A(n5660), .B(\stack[4][12] ), .Z(n5204) );
  NAND U5485 ( .A(n5205), .B(n5204), .Z(n1226) );
  NAND U5486 ( .A(n5672), .B(\stack[2][12] ), .Z(n5207) );
  NANDN U5487 ( .A(n5657), .B(\stack[4][12] ), .Z(n5206) );
  AND U5488 ( .A(n5207), .B(n5206), .Z(n5209) );
  NANDN U5489 ( .A(n5660), .B(\stack[3][12] ), .Z(n5208) );
  NAND U5490 ( .A(n5209), .B(n5208), .Z(n1227) );
  NAND U5491 ( .A(\stack[1][12] ), .B(n5672), .Z(n5211) );
  NANDN U5492 ( .A(n5657), .B(\stack[3][12] ), .Z(n5210) );
  AND U5493 ( .A(n5211), .B(n5210), .Z(n5213) );
  NANDN U5494 ( .A(n5660), .B(\stack[2][12] ), .Z(n5212) );
  NAND U5495 ( .A(n5213), .B(n5212), .Z(n1228) );
  NAND U5496 ( .A(o[12]), .B(n5672), .Z(n5215) );
  NANDN U5497 ( .A(n5657), .B(\stack[2][12] ), .Z(n5214) );
  AND U5498 ( .A(n5215), .B(n5214), .Z(n5217) );
  NANDN U5499 ( .A(n5660), .B(\stack[1][12] ), .Z(n5216) );
  NAND U5500 ( .A(n5217), .B(n5216), .Z(n1229) );
  XNOR U5501 ( .A(n5219), .B(n5218), .Z(n5220) );
  NAND U5502 ( .A(n5220), .B(n5644), .Z(n5223) );
  NAND U5503 ( .A(n5672), .B(x[12]), .Z(n5221) );
  NAND U5504 ( .A(n5223), .B(n5222), .Z(n5229) );
  NAND U5505 ( .A(n5663), .B(o[12]), .Z(n5227) );
  NAND U5506 ( .A(o[12]), .B(n5665), .Z(n5224) );
  NAND U5507 ( .A(n5667), .B(n5224), .Z(n5225) );
  AND U5508 ( .A(n5225), .B(\stack[1][12] ), .Z(n5226) );
  ANDN U5509 ( .B(n5227), .A(n5226), .Z(n5228) );
  NANDN U5510 ( .A(n5229), .B(n5228), .Z(n1230) );
  NAND U5511 ( .A(n5672), .B(\stack[6][11] ), .Z(n5231) );
  NAND U5512 ( .A(n1605), .B(\stack[7][11] ), .Z(n5230) );
  NAND U5513 ( .A(n5231), .B(n5230), .Z(n1231) );
  NAND U5514 ( .A(n5672), .B(\stack[5][11] ), .Z(n5233) );
  NANDN U5515 ( .A(n5657), .B(\stack[7][11] ), .Z(n5232) );
  AND U5516 ( .A(n5233), .B(n5232), .Z(n5235) );
  NANDN U5517 ( .A(n5660), .B(\stack[6][11] ), .Z(n5234) );
  NAND U5518 ( .A(n5235), .B(n5234), .Z(n1232) );
  NAND U5519 ( .A(n5672), .B(\stack[4][11] ), .Z(n5237) );
  NANDN U5520 ( .A(n5657), .B(\stack[6][11] ), .Z(n5236) );
  AND U5521 ( .A(n5237), .B(n5236), .Z(n5239) );
  NANDN U5522 ( .A(n5660), .B(\stack[5][11] ), .Z(n5238) );
  NAND U5523 ( .A(n5239), .B(n5238), .Z(n1233) );
  NAND U5524 ( .A(n5672), .B(\stack[3][11] ), .Z(n5241) );
  NANDN U5525 ( .A(n5657), .B(\stack[5][11] ), .Z(n5240) );
  AND U5526 ( .A(n5241), .B(n5240), .Z(n5243) );
  NANDN U5527 ( .A(n5660), .B(\stack[4][11] ), .Z(n5242) );
  NAND U5528 ( .A(n5243), .B(n5242), .Z(n1234) );
  NAND U5529 ( .A(n5672), .B(\stack[2][11] ), .Z(n5245) );
  NANDN U5530 ( .A(n5657), .B(\stack[4][11] ), .Z(n5244) );
  AND U5531 ( .A(n5245), .B(n5244), .Z(n5247) );
  NANDN U5532 ( .A(n5660), .B(\stack[3][11] ), .Z(n5246) );
  NAND U5533 ( .A(n5247), .B(n5246), .Z(n1235) );
  NAND U5534 ( .A(\stack[1][11] ), .B(n5672), .Z(n5249) );
  NANDN U5535 ( .A(n5657), .B(\stack[3][11] ), .Z(n5248) );
  AND U5536 ( .A(n5249), .B(n5248), .Z(n5251) );
  NANDN U5537 ( .A(n5660), .B(\stack[2][11] ), .Z(n5250) );
  NAND U5538 ( .A(n5251), .B(n5250), .Z(n1236) );
  NAND U5539 ( .A(o[11]), .B(n5672), .Z(n5253) );
  NANDN U5540 ( .A(n5657), .B(\stack[2][11] ), .Z(n5252) );
  AND U5541 ( .A(n5253), .B(n5252), .Z(n5255) );
  NANDN U5542 ( .A(n5660), .B(\stack[1][11] ), .Z(n5254) );
  NAND U5543 ( .A(n5255), .B(n5254), .Z(n1237) );
  XNOR U5544 ( .A(n5257), .B(n5256), .Z(n5258) );
  NAND U5545 ( .A(n5258), .B(n5644), .Z(n5262) );
  NAND U5546 ( .A(n5259), .B(n5665), .Z(n5260) );
  NAND U5547 ( .A(n5262), .B(n5261), .Z(n5268) );
  NAND U5548 ( .A(n5663), .B(o[11]), .Z(n5266) );
  NAND U5549 ( .A(n5672), .B(x[11]), .Z(n5264) );
  NAND U5550 ( .A(n5651), .B(\stack[1][11] ), .Z(n5263) );
  NAND U5551 ( .A(n5264), .B(n5263), .Z(n5265) );
  ANDN U5552 ( .B(n5266), .A(n5265), .Z(n5267) );
  NANDN U5553 ( .A(n5268), .B(n5267), .Z(n1238) );
  NAND U5554 ( .A(n5672), .B(\stack[6][10] ), .Z(n5270) );
  NAND U5555 ( .A(n1605), .B(\stack[7][10] ), .Z(n5269) );
  NAND U5556 ( .A(n5270), .B(n5269), .Z(n1239) );
  NAND U5557 ( .A(n5672), .B(\stack[5][10] ), .Z(n5272) );
  NANDN U5558 ( .A(n5657), .B(\stack[7][10] ), .Z(n5271) );
  AND U5559 ( .A(n5272), .B(n5271), .Z(n5274) );
  NANDN U5560 ( .A(n5660), .B(\stack[6][10] ), .Z(n5273) );
  NAND U5561 ( .A(n5274), .B(n5273), .Z(n1240) );
  NAND U5562 ( .A(n5672), .B(\stack[4][10] ), .Z(n5276) );
  NANDN U5563 ( .A(n5657), .B(\stack[6][10] ), .Z(n5275) );
  AND U5564 ( .A(n5276), .B(n5275), .Z(n5278) );
  NANDN U5565 ( .A(n5660), .B(\stack[5][10] ), .Z(n5277) );
  NAND U5566 ( .A(n5278), .B(n5277), .Z(n1241) );
  NAND U5567 ( .A(n5672), .B(\stack[3][10] ), .Z(n5280) );
  NANDN U5568 ( .A(n5657), .B(\stack[5][10] ), .Z(n5279) );
  AND U5569 ( .A(n5280), .B(n5279), .Z(n5282) );
  NANDN U5570 ( .A(n5660), .B(\stack[4][10] ), .Z(n5281) );
  NAND U5571 ( .A(n5282), .B(n5281), .Z(n1242) );
  NAND U5572 ( .A(n5672), .B(\stack[2][10] ), .Z(n5284) );
  NANDN U5573 ( .A(n5657), .B(\stack[4][10] ), .Z(n5283) );
  AND U5574 ( .A(n5284), .B(n5283), .Z(n5286) );
  NANDN U5575 ( .A(n5660), .B(\stack[3][10] ), .Z(n5285) );
  NAND U5576 ( .A(n5286), .B(n5285), .Z(n1243) );
  NAND U5577 ( .A(\stack[1][10] ), .B(n5672), .Z(n5288) );
  NANDN U5578 ( .A(n5657), .B(\stack[3][10] ), .Z(n5287) );
  AND U5579 ( .A(n5288), .B(n5287), .Z(n5290) );
  NANDN U5580 ( .A(n5660), .B(\stack[2][10] ), .Z(n5289) );
  NAND U5581 ( .A(n5290), .B(n5289), .Z(n1244) );
  NAND U5582 ( .A(o[10]), .B(n5672), .Z(n5292) );
  NANDN U5583 ( .A(n5657), .B(\stack[2][10] ), .Z(n5291) );
  AND U5584 ( .A(n5292), .B(n5291), .Z(n5294) );
  NANDN U5585 ( .A(n5660), .B(\stack[1][10] ), .Z(n5293) );
  NAND U5586 ( .A(n5294), .B(n5293), .Z(n1245) );
  XNOR U5587 ( .A(n5296), .B(n5295), .Z(n5297) );
  NAND U5588 ( .A(n5297), .B(n5644), .Z(n5300) );
  NAND U5589 ( .A(n5672), .B(x[10]), .Z(n5298) );
  NAND U5590 ( .A(n5300), .B(n5299), .Z(n5306) );
  NAND U5591 ( .A(n5663), .B(o[10]), .Z(n5304) );
  NAND U5592 ( .A(o[10]), .B(n5665), .Z(n5301) );
  NAND U5593 ( .A(n5667), .B(n5301), .Z(n5302) );
  AND U5594 ( .A(n5302), .B(\stack[1][10] ), .Z(n5303) );
  ANDN U5595 ( .B(n5304), .A(n5303), .Z(n5305) );
  NANDN U5596 ( .A(n5306), .B(n5305), .Z(n1246) );
  NAND U5597 ( .A(n5672), .B(\stack[6][9] ), .Z(n5308) );
  NAND U5598 ( .A(n1605), .B(\stack[7][9] ), .Z(n5307) );
  NAND U5599 ( .A(n5308), .B(n5307), .Z(n1247) );
  NAND U5600 ( .A(n5672), .B(\stack[5][9] ), .Z(n5310) );
  NANDN U5601 ( .A(n5657), .B(\stack[7][9] ), .Z(n5309) );
  AND U5602 ( .A(n5310), .B(n5309), .Z(n5312) );
  NANDN U5603 ( .A(n5660), .B(\stack[6][9] ), .Z(n5311) );
  NAND U5604 ( .A(n5312), .B(n5311), .Z(n1248) );
  NAND U5605 ( .A(n5672), .B(\stack[4][9] ), .Z(n5314) );
  NANDN U5606 ( .A(n5657), .B(\stack[6][9] ), .Z(n5313) );
  AND U5607 ( .A(n5314), .B(n5313), .Z(n5316) );
  NANDN U5608 ( .A(n5660), .B(\stack[5][9] ), .Z(n5315) );
  NAND U5609 ( .A(n5316), .B(n5315), .Z(n1249) );
  NAND U5610 ( .A(n5672), .B(\stack[3][9] ), .Z(n5318) );
  NANDN U5611 ( .A(n5657), .B(\stack[5][9] ), .Z(n5317) );
  AND U5612 ( .A(n5318), .B(n5317), .Z(n5320) );
  NANDN U5613 ( .A(n5660), .B(\stack[4][9] ), .Z(n5319) );
  NAND U5614 ( .A(n5320), .B(n5319), .Z(n1250) );
  NAND U5615 ( .A(n5672), .B(\stack[2][9] ), .Z(n5322) );
  NANDN U5616 ( .A(n5657), .B(\stack[4][9] ), .Z(n5321) );
  AND U5617 ( .A(n5322), .B(n5321), .Z(n5324) );
  NANDN U5618 ( .A(n5660), .B(\stack[3][9] ), .Z(n5323) );
  NAND U5619 ( .A(n5324), .B(n5323), .Z(n1251) );
  NAND U5620 ( .A(\stack[1][9] ), .B(n5672), .Z(n5326) );
  NANDN U5621 ( .A(n5657), .B(\stack[3][9] ), .Z(n5325) );
  AND U5622 ( .A(n5326), .B(n5325), .Z(n5328) );
  NANDN U5623 ( .A(n5660), .B(\stack[2][9] ), .Z(n5327) );
  NAND U5624 ( .A(n5328), .B(n5327), .Z(n1252) );
  NAND U5625 ( .A(o[9]), .B(n5672), .Z(n5330) );
  NANDN U5626 ( .A(n5657), .B(\stack[2][9] ), .Z(n5329) );
  AND U5627 ( .A(n5330), .B(n5329), .Z(n5332) );
  NANDN U5628 ( .A(n5660), .B(\stack[1][9] ), .Z(n5331) );
  NAND U5629 ( .A(n5332), .B(n5331), .Z(n1253) );
  XNOR U5630 ( .A(n5334), .B(n5333), .Z(n5335) );
  NAND U5631 ( .A(n5335), .B(n5644), .Z(n5339) );
  NAND U5632 ( .A(n5336), .B(n5665), .Z(n5337) );
  NAND U5633 ( .A(n5339), .B(n5338), .Z(n5345) );
  NAND U5634 ( .A(n5663), .B(o[9]), .Z(n5343) );
  NAND U5635 ( .A(n5672), .B(x[9]), .Z(n5341) );
  NAND U5636 ( .A(n5651), .B(\stack[1][9] ), .Z(n5340) );
  NAND U5637 ( .A(n5341), .B(n5340), .Z(n5342) );
  ANDN U5638 ( .B(n5343), .A(n5342), .Z(n5344) );
  NANDN U5639 ( .A(n5345), .B(n5344), .Z(n1254) );
  NAND U5640 ( .A(n5672), .B(\stack[6][8] ), .Z(n5347) );
  NAND U5641 ( .A(n1605), .B(\stack[7][8] ), .Z(n5346) );
  NAND U5642 ( .A(n5347), .B(n5346), .Z(n1255) );
  NAND U5643 ( .A(n5672), .B(\stack[5][8] ), .Z(n5349) );
  NANDN U5644 ( .A(n5657), .B(\stack[7][8] ), .Z(n5348) );
  AND U5645 ( .A(n5349), .B(n5348), .Z(n5351) );
  NANDN U5646 ( .A(n5660), .B(\stack[6][8] ), .Z(n5350) );
  NAND U5647 ( .A(n5351), .B(n5350), .Z(n1256) );
  NAND U5648 ( .A(n5672), .B(\stack[4][8] ), .Z(n5353) );
  NANDN U5649 ( .A(n5657), .B(\stack[6][8] ), .Z(n5352) );
  AND U5650 ( .A(n5353), .B(n5352), .Z(n5355) );
  NANDN U5651 ( .A(n5660), .B(\stack[5][8] ), .Z(n5354) );
  NAND U5652 ( .A(n5355), .B(n5354), .Z(n1257) );
  NAND U5653 ( .A(n5672), .B(\stack[3][8] ), .Z(n5357) );
  NANDN U5654 ( .A(n5657), .B(\stack[5][8] ), .Z(n5356) );
  AND U5655 ( .A(n5357), .B(n5356), .Z(n5359) );
  NANDN U5656 ( .A(n5660), .B(\stack[4][8] ), .Z(n5358) );
  NAND U5657 ( .A(n5359), .B(n5358), .Z(n1258) );
  NAND U5658 ( .A(n5672), .B(\stack[2][8] ), .Z(n5361) );
  NANDN U5659 ( .A(n5657), .B(\stack[4][8] ), .Z(n5360) );
  AND U5660 ( .A(n5361), .B(n5360), .Z(n5363) );
  NANDN U5661 ( .A(n5660), .B(\stack[3][8] ), .Z(n5362) );
  NAND U5662 ( .A(n5363), .B(n5362), .Z(n1259) );
  NAND U5663 ( .A(\stack[1][8] ), .B(n5672), .Z(n5365) );
  NANDN U5664 ( .A(n5657), .B(\stack[3][8] ), .Z(n5364) );
  AND U5665 ( .A(n5365), .B(n5364), .Z(n5367) );
  NANDN U5666 ( .A(n5660), .B(\stack[2][8] ), .Z(n5366) );
  NAND U5667 ( .A(n5367), .B(n5366), .Z(n1260) );
  NAND U5668 ( .A(o[8]), .B(n5672), .Z(n5369) );
  NANDN U5669 ( .A(n5657), .B(\stack[2][8] ), .Z(n5368) );
  AND U5670 ( .A(n5369), .B(n5368), .Z(n5371) );
  NANDN U5671 ( .A(n5660), .B(\stack[1][8] ), .Z(n5370) );
  NAND U5672 ( .A(n5371), .B(n5370), .Z(n1261) );
  XNOR U5673 ( .A(n5373), .B(n5372), .Z(n5374) );
  NAND U5674 ( .A(n5374), .B(n5644), .Z(n5377) );
  NAND U5675 ( .A(n5672), .B(x[8]), .Z(n5375) );
  NAND U5676 ( .A(n5377), .B(n5376), .Z(n5383) );
  NAND U5677 ( .A(n5663), .B(o[8]), .Z(n5381) );
  NAND U5678 ( .A(o[8]), .B(n5665), .Z(n5378) );
  NAND U5679 ( .A(n5667), .B(n5378), .Z(n5379) );
  AND U5680 ( .A(n5379), .B(\stack[1][8] ), .Z(n5380) );
  ANDN U5681 ( .B(n5381), .A(n5380), .Z(n5382) );
  NANDN U5682 ( .A(n5383), .B(n5382), .Z(n1262) );
  NAND U5683 ( .A(n5672), .B(\stack[6][7] ), .Z(n5385) );
  NAND U5684 ( .A(n1605), .B(\stack[7][7] ), .Z(n5384) );
  NAND U5685 ( .A(n5385), .B(n5384), .Z(n1263) );
  NAND U5686 ( .A(n5672), .B(\stack[5][7] ), .Z(n5387) );
  NANDN U5687 ( .A(n5657), .B(\stack[7][7] ), .Z(n5386) );
  AND U5688 ( .A(n5387), .B(n5386), .Z(n5389) );
  NANDN U5689 ( .A(n5660), .B(\stack[6][7] ), .Z(n5388) );
  NAND U5690 ( .A(n5389), .B(n5388), .Z(n1264) );
  NAND U5691 ( .A(n5672), .B(\stack[4][7] ), .Z(n5391) );
  NANDN U5692 ( .A(n5657), .B(\stack[6][7] ), .Z(n5390) );
  AND U5693 ( .A(n5391), .B(n5390), .Z(n5393) );
  NANDN U5694 ( .A(n5660), .B(\stack[5][7] ), .Z(n5392) );
  NAND U5695 ( .A(n5393), .B(n5392), .Z(n1265) );
  NAND U5696 ( .A(n5672), .B(\stack[3][7] ), .Z(n5395) );
  NANDN U5697 ( .A(n5657), .B(\stack[5][7] ), .Z(n5394) );
  AND U5698 ( .A(n5395), .B(n5394), .Z(n5397) );
  NANDN U5699 ( .A(n5660), .B(\stack[4][7] ), .Z(n5396) );
  NAND U5700 ( .A(n5397), .B(n5396), .Z(n1266) );
  NAND U5701 ( .A(n5672), .B(\stack[2][7] ), .Z(n5399) );
  NANDN U5702 ( .A(n5657), .B(\stack[4][7] ), .Z(n5398) );
  AND U5703 ( .A(n5399), .B(n5398), .Z(n5401) );
  NANDN U5704 ( .A(n5660), .B(\stack[3][7] ), .Z(n5400) );
  NAND U5705 ( .A(n5401), .B(n5400), .Z(n1267) );
  NAND U5706 ( .A(\stack[1][7] ), .B(n5672), .Z(n5403) );
  NANDN U5707 ( .A(n5657), .B(\stack[3][7] ), .Z(n5402) );
  AND U5708 ( .A(n5403), .B(n5402), .Z(n5405) );
  NANDN U5709 ( .A(n5660), .B(\stack[2][7] ), .Z(n5404) );
  NAND U5710 ( .A(n5405), .B(n5404), .Z(n1268) );
  NAND U5711 ( .A(o[7]), .B(n5672), .Z(n5407) );
  NANDN U5712 ( .A(n5657), .B(\stack[2][7] ), .Z(n5406) );
  AND U5713 ( .A(n5407), .B(n5406), .Z(n5409) );
  NANDN U5714 ( .A(n5660), .B(\stack[1][7] ), .Z(n5408) );
  NAND U5715 ( .A(n5409), .B(n5408), .Z(n1269) );
  XNOR U5716 ( .A(n5411), .B(n5410), .Z(n5412) );
  NAND U5717 ( .A(n5412), .B(n5644), .Z(n5415) );
  NAND U5718 ( .A(\stack[1][7] ), .B(n5651), .Z(n5413) );
  NAND U5719 ( .A(n5415), .B(n5414), .Z(n5422) );
  NAND U5720 ( .A(n5663), .B(o[7]), .Z(n5420) );
  NAND U5721 ( .A(n5672), .B(x[7]), .Z(n5418) );
  NAND U5722 ( .A(n5665), .B(n5416), .Z(n5417) );
  NAND U5723 ( .A(n5418), .B(n5417), .Z(n5419) );
  ANDN U5724 ( .B(n5420), .A(n5419), .Z(n5421) );
  NANDN U5725 ( .A(n5422), .B(n5421), .Z(n1270) );
  NAND U5726 ( .A(n5672), .B(\stack[6][6] ), .Z(n5424) );
  NAND U5727 ( .A(n1605), .B(\stack[7][6] ), .Z(n5423) );
  NAND U5728 ( .A(n5424), .B(n5423), .Z(n1271) );
  NAND U5729 ( .A(n5672), .B(\stack[5][6] ), .Z(n5426) );
  NANDN U5730 ( .A(n5657), .B(\stack[7][6] ), .Z(n5425) );
  AND U5731 ( .A(n5426), .B(n5425), .Z(n5428) );
  NANDN U5732 ( .A(n5660), .B(\stack[6][6] ), .Z(n5427) );
  NAND U5733 ( .A(n5428), .B(n5427), .Z(n1272) );
  NAND U5734 ( .A(n5672), .B(\stack[4][6] ), .Z(n5430) );
  NANDN U5735 ( .A(n5657), .B(\stack[6][6] ), .Z(n5429) );
  AND U5736 ( .A(n5430), .B(n5429), .Z(n5432) );
  NANDN U5737 ( .A(n5660), .B(\stack[5][6] ), .Z(n5431) );
  NAND U5738 ( .A(n5432), .B(n5431), .Z(n1273) );
  NAND U5739 ( .A(n5672), .B(\stack[3][6] ), .Z(n5434) );
  NANDN U5740 ( .A(n5657), .B(\stack[5][6] ), .Z(n5433) );
  AND U5741 ( .A(n5434), .B(n5433), .Z(n5436) );
  NANDN U5742 ( .A(n5660), .B(\stack[4][6] ), .Z(n5435) );
  NAND U5743 ( .A(n5436), .B(n5435), .Z(n1274) );
  NAND U5744 ( .A(n5672), .B(\stack[2][6] ), .Z(n5438) );
  NANDN U5745 ( .A(n5657), .B(\stack[4][6] ), .Z(n5437) );
  AND U5746 ( .A(n5438), .B(n5437), .Z(n5440) );
  NANDN U5747 ( .A(n5660), .B(\stack[3][6] ), .Z(n5439) );
  NAND U5748 ( .A(n5440), .B(n5439), .Z(n1275) );
  NAND U5749 ( .A(\stack[1][6] ), .B(n5672), .Z(n5442) );
  NANDN U5750 ( .A(n5657), .B(\stack[3][6] ), .Z(n5441) );
  AND U5751 ( .A(n5442), .B(n5441), .Z(n5444) );
  NANDN U5752 ( .A(n5660), .B(\stack[2][6] ), .Z(n5443) );
  NAND U5753 ( .A(n5444), .B(n5443), .Z(n1276) );
  NAND U5754 ( .A(o[6]), .B(n5672), .Z(n5446) );
  NANDN U5755 ( .A(n5657), .B(\stack[2][6] ), .Z(n5445) );
  AND U5756 ( .A(n5446), .B(n5445), .Z(n5448) );
  NANDN U5757 ( .A(n5660), .B(\stack[1][6] ), .Z(n5447) );
  NAND U5758 ( .A(n5448), .B(n5447), .Z(n1277) );
  XNOR U5759 ( .A(n5450), .B(n5449), .Z(n5451) );
  NAND U5760 ( .A(n5451), .B(n5644), .Z(n5455) );
  NAND U5761 ( .A(n5452), .B(n5665), .Z(n5453) );
  NAND U5762 ( .A(n5455), .B(n5454), .Z(n5461) );
  NAND U5763 ( .A(n5663), .B(o[6]), .Z(n5459) );
  NAND U5764 ( .A(n5672), .B(x[6]), .Z(n5457) );
  NAND U5765 ( .A(n5651), .B(\stack[1][6] ), .Z(n5456) );
  NAND U5766 ( .A(n5457), .B(n5456), .Z(n5458) );
  ANDN U5767 ( .B(n5459), .A(n5458), .Z(n5460) );
  NANDN U5768 ( .A(n5461), .B(n5460), .Z(n1278) );
  NAND U5769 ( .A(n5672), .B(\stack[6][5] ), .Z(n5463) );
  NAND U5770 ( .A(n1605), .B(\stack[7][5] ), .Z(n5462) );
  NAND U5771 ( .A(n5463), .B(n5462), .Z(n1279) );
  NAND U5772 ( .A(n5672), .B(\stack[5][5] ), .Z(n5465) );
  NANDN U5773 ( .A(n5657), .B(\stack[7][5] ), .Z(n5464) );
  AND U5774 ( .A(n5465), .B(n5464), .Z(n5467) );
  NANDN U5775 ( .A(n5660), .B(\stack[6][5] ), .Z(n5466) );
  NAND U5776 ( .A(n5467), .B(n5466), .Z(n1280) );
  NAND U5777 ( .A(n5672), .B(\stack[4][5] ), .Z(n5469) );
  NANDN U5778 ( .A(n5657), .B(\stack[6][5] ), .Z(n5468) );
  AND U5779 ( .A(n5469), .B(n5468), .Z(n5471) );
  NANDN U5780 ( .A(n5660), .B(\stack[5][5] ), .Z(n5470) );
  NAND U5781 ( .A(n5471), .B(n5470), .Z(n1281) );
  NAND U5782 ( .A(n5672), .B(\stack[3][5] ), .Z(n5473) );
  NANDN U5783 ( .A(n5657), .B(\stack[5][5] ), .Z(n5472) );
  AND U5784 ( .A(n5473), .B(n5472), .Z(n5475) );
  NANDN U5785 ( .A(n5660), .B(\stack[4][5] ), .Z(n5474) );
  NAND U5786 ( .A(n5475), .B(n5474), .Z(n1282) );
  NAND U5787 ( .A(n5672), .B(\stack[2][5] ), .Z(n5477) );
  NANDN U5788 ( .A(n5657), .B(\stack[4][5] ), .Z(n5476) );
  AND U5789 ( .A(n5477), .B(n5476), .Z(n5479) );
  NANDN U5790 ( .A(n5660), .B(\stack[3][5] ), .Z(n5478) );
  NAND U5791 ( .A(n5479), .B(n5478), .Z(n1283) );
  NAND U5792 ( .A(\stack[1][5] ), .B(n5672), .Z(n5481) );
  NANDN U5793 ( .A(n5657), .B(\stack[3][5] ), .Z(n5480) );
  AND U5794 ( .A(n5481), .B(n5480), .Z(n5483) );
  NANDN U5795 ( .A(n5660), .B(\stack[2][5] ), .Z(n5482) );
  NAND U5796 ( .A(n5483), .B(n5482), .Z(n1284) );
  NAND U5797 ( .A(o[5]), .B(n5672), .Z(n5485) );
  NANDN U5798 ( .A(n5657), .B(\stack[2][5] ), .Z(n5484) );
  AND U5799 ( .A(n5485), .B(n5484), .Z(n5487) );
  NANDN U5800 ( .A(n5660), .B(\stack[1][5] ), .Z(n5486) );
  NAND U5801 ( .A(n5487), .B(n5486), .Z(n1285) );
  XNOR U5802 ( .A(n5489), .B(n5488), .Z(n5490) );
  NAND U5803 ( .A(n5490), .B(n5644), .Z(n5493) );
  NAND U5804 ( .A(n5672), .B(x[5]), .Z(n5491) );
  NAND U5805 ( .A(n5493), .B(n5492), .Z(n5499) );
  NAND U5806 ( .A(n5663), .B(o[5]), .Z(n5497) );
  NAND U5807 ( .A(o[5]), .B(n5665), .Z(n5494) );
  NAND U5808 ( .A(n5667), .B(n5494), .Z(n5495) );
  AND U5809 ( .A(n5495), .B(\stack[1][5] ), .Z(n5496) );
  ANDN U5810 ( .B(n5497), .A(n5496), .Z(n5498) );
  NANDN U5811 ( .A(n5499), .B(n5498), .Z(n1286) );
  NAND U5812 ( .A(n5672), .B(\stack[6][4] ), .Z(n5501) );
  NAND U5813 ( .A(n1605), .B(\stack[7][4] ), .Z(n5500) );
  NAND U5814 ( .A(n5501), .B(n5500), .Z(n1287) );
  NAND U5815 ( .A(n5672), .B(\stack[5][4] ), .Z(n5503) );
  NANDN U5816 ( .A(n5657), .B(\stack[7][4] ), .Z(n5502) );
  AND U5817 ( .A(n5503), .B(n5502), .Z(n5505) );
  NANDN U5818 ( .A(n5660), .B(\stack[6][4] ), .Z(n5504) );
  NAND U5819 ( .A(n5505), .B(n5504), .Z(n1288) );
  NAND U5820 ( .A(n5672), .B(\stack[4][4] ), .Z(n5507) );
  NANDN U5821 ( .A(n5657), .B(\stack[6][4] ), .Z(n5506) );
  AND U5822 ( .A(n5507), .B(n5506), .Z(n5509) );
  NANDN U5823 ( .A(n5660), .B(\stack[5][4] ), .Z(n5508) );
  NAND U5824 ( .A(n5509), .B(n5508), .Z(n1289) );
  NAND U5825 ( .A(n5672), .B(\stack[3][4] ), .Z(n5511) );
  NANDN U5826 ( .A(n5657), .B(\stack[5][4] ), .Z(n5510) );
  AND U5827 ( .A(n5511), .B(n5510), .Z(n5513) );
  NANDN U5828 ( .A(n5660), .B(\stack[4][4] ), .Z(n5512) );
  NAND U5829 ( .A(n5513), .B(n5512), .Z(n1290) );
  NAND U5830 ( .A(n5672), .B(\stack[2][4] ), .Z(n5515) );
  NANDN U5831 ( .A(n5657), .B(\stack[4][4] ), .Z(n5514) );
  AND U5832 ( .A(n5515), .B(n5514), .Z(n5517) );
  NANDN U5833 ( .A(n5660), .B(\stack[3][4] ), .Z(n5516) );
  NAND U5834 ( .A(n5517), .B(n5516), .Z(n1291) );
  NAND U5835 ( .A(\stack[1][4] ), .B(n5672), .Z(n5519) );
  NANDN U5836 ( .A(n5657), .B(\stack[3][4] ), .Z(n5518) );
  AND U5837 ( .A(n5519), .B(n5518), .Z(n5521) );
  NANDN U5838 ( .A(n5660), .B(\stack[2][4] ), .Z(n5520) );
  NAND U5839 ( .A(n5521), .B(n5520), .Z(n1292) );
  NAND U5840 ( .A(o[4]), .B(n5672), .Z(n5523) );
  NANDN U5841 ( .A(n5657), .B(\stack[2][4] ), .Z(n5522) );
  AND U5842 ( .A(n5523), .B(n5522), .Z(n5525) );
  NANDN U5843 ( .A(n5660), .B(\stack[1][4] ), .Z(n5524) );
  NAND U5844 ( .A(n5525), .B(n5524), .Z(n1293) );
  XNOR U5845 ( .A(n5527), .B(n5526), .Z(n5528) );
  NAND U5846 ( .A(n5528), .B(n5644), .Z(n5531) );
  NAND U5847 ( .A(n5672), .B(x[4]), .Z(n5529) );
  NAND U5848 ( .A(n5531), .B(n5530), .Z(n5537) );
  NAND U5849 ( .A(n5663), .B(o[4]), .Z(n5535) );
  NAND U5850 ( .A(o[4]), .B(n5665), .Z(n5532) );
  NAND U5851 ( .A(n5667), .B(n5532), .Z(n5533) );
  AND U5852 ( .A(n5533), .B(\stack[1][4] ), .Z(n5534) );
  ANDN U5853 ( .B(n5535), .A(n5534), .Z(n5536) );
  NANDN U5854 ( .A(n5537), .B(n5536), .Z(n1294) );
  NAND U5855 ( .A(n5672), .B(\stack[6][3] ), .Z(n5539) );
  NAND U5856 ( .A(n1605), .B(\stack[7][3] ), .Z(n5538) );
  NAND U5857 ( .A(n5539), .B(n5538), .Z(n1295) );
  NAND U5858 ( .A(n5672), .B(\stack[5][3] ), .Z(n5541) );
  NANDN U5859 ( .A(n5657), .B(\stack[7][3] ), .Z(n5540) );
  AND U5860 ( .A(n5541), .B(n5540), .Z(n5543) );
  NANDN U5861 ( .A(n5660), .B(\stack[6][3] ), .Z(n5542) );
  NAND U5862 ( .A(n5543), .B(n5542), .Z(n1296) );
  NAND U5863 ( .A(n5672), .B(\stack[4][3] ), .Z(n5545) );
  NANDN U5864 ( .A(n5657), .B(\stack[6][3] ), .Z(n5544) );
  AND U5865 ( .A(n5545), .B(n5544), .Z(n5547) );
  NANDN U5866 ( .A(n5660), .B(\stack[5][3] ), .Z(n5546) );
  NAND U5867 ( .A(n5547), .B(n5546), .Z(n1297) );
  NAND U5868 ( .A(n5672), .B(\stack[3][3] ), .Z(n5549) );
  NANDN U5869 ( .A(n5657), .B(\stack[5][3] ), .Z(n5548) );
  AND U5870 ( .A(n5549), .B(n5548), .Z(n5551) );
  NANDN U5871 ( .A(n5660), .B(\stack[4][3] ), .Z(n5550) );
  NAND U5872 ( .A(n5551), .B(n5550), .Z(n1298) );
  NAND U5873 ( .A(n5672), .B(\stack[2][3] ), .Z(n5553) );
  NANDN U5874 ( .A(n5657), .B(\stack[4][3] ), .Z(n5552) );
  AND U5875 ( .A(n5553), .B(n5552), .Z(n5555) );
  NANDN U5876 ( .A(n5660), .B(\stack[3][3] ), .Z(n5554) );
  NAND U5877 ( .A(n5555), .B(n5554), .Z(n1299) );
  NAND U5878 ( .A(\stack[1][3] ), .B(n5672), .Z(n5557) );
  NANDN U5879 ( .A(n5657), .B(\stack[3][3] ), .Z(n5556) );
  AND U5880 ( .A(n5557), .B(n5556), .Z(n5559) );
  NANDN U5881 ( .A(n5660), .B(\stack[2][3] ), .Z(n5558) );
  NAND U5882 ( .A(n5559), .B(n5558), .Z(n1300) );
  NAND U5883 ( .A(o[3]), .B(n5672), .Z(n5561) );
  NANDN U5884 ( .A(n5657), .B(\stack[2][3] ), .Z(n5560) );
  AND U5885 ( .A(n5561), .B(n5560), .Z(n5563) );
  NANDN U5886 ( .A(n5660), .B(\stack[1][3] ), .Z(n5562) );
  NAND U5887 ( .A(n5563), .B(n5562), .Z(n1301) );
  NAND U5888 ( .A(\stack[1][3] ), .B(n5651), .Z(n5564) );
  XNOR U5889 ( .A(n5566), .B(n5565), .Z(n5567) );
  NAND U5890 ( .A(n5567), .B(n5644), .Z(n5568) );
  NANDN U5891 ( .A(n5569), .B(n5568), .Z(n5576) );
  NAND U5892 ( .A(n5663), .B(o[3]), .Z(n5574) );
  NAND U5893 ( .A(n5672), .B(x[3]), .Z(n5572) );
  NAND U5894 ( .A(n5570), .B(n5665), .Z(n5571) );
  NAND U5895 ( .A(n5572), .B(n5571), .Z(n5573) );
  ANDN U5896 ( .B(n5574), .A(n5573), .Z(n5575) );
  NANDN U5897 ( .A(n5576), .B(n5575), .Z(n1302) );
  NAND U5898 ( .A(n5672), .B(\stack[6][2] ), .Z(n5578) );
  NAND U5899 ( .A(n1605), .B(\stack[7][2] ), .Z(n5577) );
  NAND U5900 ( .A(n5578), .B(n5577), .Z(n1303) );
  NAND U5901 ( .A(n5672), .B(\stack[5][2] ), .Z(n5580) );
  NANDN U5902 ( .A(n5657), .B(\stack[7][2] ), .Z(n5579) );
  AND U5903 ( .A(n5580), .B(n5579), .Z(n5582) );
  NANDN U5904 ( .A(n5660), .B(\stack[6][2] ), .Z(n5581) );
  NAND U5905 ( .A(n5582), .B(n5581), .Z(n1304) );
  NAND U5906 ( .A(n5672), .B(\stack[4][2] ), .Z(n5584) );
  NANDN U5907 ( .A(n5657), .B(\stack[6][2] ), .Z(n5583) );
  AND U5908 ( .A(n5584), .B(n5583), .Z(n5586) );
  NANDN U5909 ( .A(n5660), .B(\stack[5][2] ), .Z(n5585) );
  NAND U5910 ( .A(n5586), .B(n5585), .Z(n1305) );
  NAND U5911 ( .A(n5672), .B(\stack[3][2] ), .Z(n5588) );
  NANDN U5912 ( .A(n5657), .B(\stack[5][2] ), .Z(n5587) );
  AND U5913 ( .A(n5588), .B(n5587), .Z(n5590) );
  NANDN U5914 ( .A(n5660), .B(\stack[4][2] ), .Z(n5589) );
  NAND U5915 ( .A(n5590), .B(n5589), .Z(n1306) );
  NAND U5916 ( .A(n5672), .B(\stack[2][2] ), .Z(n5592) );
  NANDN U5917 ( .A(n5657), .B(\stack[4][2] ), .Z(n5591) );
  AND U5918 ( .A(n5592), .B(n5591), .Z(n5594) );
  NANDN U5919 ( .A(n5660), .B(\stack[3][2] ), .Z(n5593) );
  NAND U5920 ( .A(n5594), .B(n5593), .Z(n1307) );
  NAND U5921 ( .A(\stack[1][2] ), .B(n5672), .Z(n5596) );
  NANDN U5922 ( .A(n5657), .B(\stack[3][2] ), .Z(n5595) );
  AND U5923 ( .A(n5596), .B(n5595), .Z(n5598) );
  NANDN U5924 ( .A(n5660), .B(\stack[2][2] ), .Z(n5597) );
  NAND U5925 ( .A(n5598), .B(n5597), .Z(n1308) );
  NAND U5926 ( .A(n5672), .B(o[2]), .Z(n5600) );
  NANDN U5927 ( .A(n5657), .B(\stack[2][2] ), .Z(n5599) );
  AND U5928 ( .A(n5600), .B(n5599), .Z(n5602) );
  NANDN U5929 ( .A(n5660), .B(\stack[1][2] ), .Z(n5601) );
  NAND U5930 ( .A(n5602), .B(n5601), .Z(n1309) );
  XNOR U5931 ( .A(n5604), .B(n5603), .Z(n5605) );
  NAND U5932 ( .A(n5605), .B(n5644), .Z(n5615) );
  NANDN U5933 ( .A(n5606), .B(n5665), .Z(n5607) );
  NAND U5934 ( .A(n5672), .B(x[2]), .Z(n5609) );
  NAND U5935 ( .A(n5651), .B(\stack[1][2] ), .Z(n5608) );
  NAND U5936 ( .A(n5609), .B(n5608), .Z(n5610) );
  NOR U5937 ( .A(n5611), .B(n5610), .Z(n5613) );
  NAND U5938 ( .A(n5663), .B(o[2]), .Z(n5612) );
  AND U5939 ( .A(n5613), .B(n5612), .Z(n5614) );
  NAND U5940 ( .A(n5615), .B(n5614), .Z(n1310) );
  NAND U5941 ( .A(n5672), .B(\stack[6][1] ), .Z(n5617) );
  NAND U5942 ( .A(n1605), .B(\stack[7][1] ), .Z(n5616) );
  NAND U5943 ( .A(n5617), .B(n5616), .Z(n1311) );
  NAND U5944 ( .A(n5672), .B(\stack[5][1] ), .Z(n5619) );
  NANDN U5945 ( .A(n5657), .B(\stack[7][1] ), .Z(n5618) );
  AND U5946 ( .A(n5619), .B(n5618), .Z(n5621) );
  NANDN U5947 ( .A(n5660), .B(\stack[6][1] ), .Z(n5620) );
  NAND U5948 ( .A(n5621), .B(n5620), .Z(n1312) );
  NAND U5949 ( .A(n5672), .B(\stack[4][1] ), .Z(n5623) );
  NANDN U5950 ( .A(n5657), .B(\stack[6][1] ), .Z(n5622) );
  AND U5951 ( .A(n5623), .B(n5622), .Z(n5625) );
  NANDN U5952 ( .A(n5660), .B(\stack[5][1] ), .Z(n5624) );
  NAND U5953 ( .A(n5625), .B(n5624), .Z(n1313) );
  NAND U5954 ( .A(n5672), .B(\stack[3][1] ), .Z(n5627) );
  NANDN U5955 ( .A(n5657), .B(\stack[5][1] ), .Z(n5626) );
  AND U5956 ( .A(n5627), .B(n5626), .Z(n5629) );
  NANDN U5957 ( .A(n5660), .B(\stack[4][1] ), .Z(n5628) );
  NAND U5958 ( .A(n5629), .B(n5628), .Z(n1314) );
  NAND U5959 ( .A(n5672), .B(\stack[2][1] ), .Z(n5631) );
  NANDN U5960 ( .A(n5657), .B(\stack[4][1] ), .Z(n5630) );
  AND U5961 ( .A(n5631), .B(n5630), .Z(n5633) );
  NANDN U5962 ( .A(n5660), .B(\stack[3][1] ), .Z(n5632) );
  NAND U5963 ( .A(n5633), .B(n5632), .Z(n1315) );
  NAND U5964 ( .A(\stack[1][1] ), .B(n5672), .Z(n5635) );
  NANDN U5965 ( .A(n5657), .B(\stack[3][1] ), .Z(n5634) );
  AND U5966 ( .A(n5635), .B(n5634), .Z(n5637) );
  NANDN U5967 ( .A(n5660), .B(\stack[2][1] ), .Z(n5636) );
  NAND U5968 ( .A(n5637), .B(n5636), .Z(n1316) );
  NAND U5969 ( .A(o[1]), .B(n5672), .Z(n5639) );
  NANDN U5970 ( .A(n5657), .B(\stack[2][1] ), .Z(n5638) );
  AND U5971 ( .A(n5639), .B(n5638), .Z(n5641) );
  NANDN U5972 ( .A(n5660), .B(\stack[1][1] ), .Z(n5640) );
  NAND U5973 ( .A(n5641), .B(n5640), .Z(n1317) );
  XNOR U5974 ( .A(n5643), .B(n5642), .Z(n5645) );
  NAND U5975 ( .A(n5645), .B(n5644), .Z(n5650) );
  NAND U5976 ( .A(n5672), .B(x[1]), .Z(n5648) );
  NAND U5977 ( .A(o[1]), .B(\stack[1][1] ), .Z(n5646) );
  NANDN U5978 ( .A(n5646), .B(n5665), .Z(n5647) );
  AND U5979 ( .A(n5648), .B(n5647), .Z(n5649) );
  AND U5980 ( .A(n5650), .B(n5649), .Z(n5653) );
  NAND U5981 ( .A(n5651), .B(\stack[1][1] ), .Z(n5652) );
  AND U5982 ( .A(n5653), .B(n5652), .Z(n5656) );
  NAND U5983 ( .A(o[1]), .B(n5663), .Z(n5654) );
  NAND U5984 ( .A(n5656), .B(n5655), .Z(n1318) );
  NAND U5985 ( .A(n5672), .B(o[0]), .Z(n5659) );
  NANDN U5986 ( .A(n5657), .B(\stack[2][0] ), .Z(n5658) );
  AND U5987 ( .A(n5659), .B(n5658), .Z(n5662) );
  NANDN U5988 ( .A(n5660), .B(\stack[1][0] ), .Z(n5661) );
  NAND U5989 ( .A(n5662), .B(n5661), .Z(n1319) );
  NAND U5990 ( .A(n5663), .B(o[0]), .Z(n5671) );
  OR U5991 ( .A(n5665), .B(n5664), .Z(n5666) );
  NAND U5992 ( .A(n5666), .B(o[0]), .Z(n5668) );
  AND U5993 ( .A(n5668), .B(n5667), .Z(n5669) );
  NANDN U5994 ( .A(n5669), .B(\stack[1][0] ), .Z(n5670) );
  AND U5995 ( .A(n5671), .B(n5670), .Z(n5675) );
  NAND U5996 ( .A(n5672), .B(x[0]), .Z(n5673) );
  NAND U5997 ( .A(n5675), .B(n5674), .Z(n1320) );
endmodule

